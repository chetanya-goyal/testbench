* NGSPICE file created from diffpair568.ext - technology: sky130A

.subckt diffpair568 minus drain_right drain_left source plus
X0 source.t39 minus.t0 drain_right.t13 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X1 drain_right.t12 minus.t1 source.t38 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 source.t13 plus.t0 drain_left.t19 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 drain_right.t7 minus.t2 source.t37 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X4 source.t36 minus.t3 drain_right.t6 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X5 source.t11 plus.t1 drain_left.t18 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X6 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X7 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X8 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X9 drain_left.t17 plus.t2 source.t15 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X10 drain_left.t16 plus.t3 source.t1 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source.t6 plus.t4 drain_left.t15 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 source.t35 minus.t4 drain_right.t17 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X13 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X14 source.t2 plus.t5 drain_left.t14 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 drain_right.t16 minus.t5 source.t34 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X16 drain_right.t15 minus.t6 source.t33 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_left.t13 plus.t6 source.t5 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X18 source.t32 minus.t7 drain_right.t14 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 source.t31 minus.t8 drain_right.t3 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X20 drain_right.t2 minus.t9 source.t30 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 source.t29 minus.t10 drain_right.t19 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 drain_left.t12 plus.t7 source.t17 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X23 drain_left.t11 plus.t8 source.t16 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X24 source.t8 plus.t9 drain_left.t10 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X25 drain_right.t18 minus.t11 source.t28 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X26 drain_right.t9 minus.t12 source.t27 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 source.t26 minus.t13 drain_right.t8 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X28 drain_right.t1 minus.t14 source.t25 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X29 drain_left.t9 plus.t10 source.t7 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X30 drain_left.t8 plus.t11 source.t18 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X31 source.t24 minus.t15 drain_right.t0 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X32 drain_right.t11 minus.t16 source.t23 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X33 drain_left.t7 plus.t12 source.t19 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X34 source.t3 plus.t13 drain_left.t6 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X35 source.t14 plus.t14 drain_left.t5 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X36 drain_right.t10 minus.t17 source.t22 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X37 source.t0 plus.t15 drain_left.t4 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X38 source.t21 minus.t18 drain_right.t5 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X39 source.t10 plus.t16 drain_left.t3 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X40 drain_left.t2 plus.t17 source.t12 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X41 drain_left.t1 plus.t18 source.t4 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X42 source.t20 minus.t19 drain_right.t4 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X43 source.t9 plus.t19 drain_left.t0 a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n27 minus.t18 3484.28
R1 minus.n7 minus.t5 3484.28
R2 minus.n56 minus.t17 3484.28
R3 minus.n35 minus.t3 3484.28
R4 minus.n26 minus.t9 3422.2
R5 minus.n24 minus.t13 3422.2
R6 minus.n3 minus.t12 3422.2
R7 minus.n18 minus.t15 3422.2
R8 minus.n16 minus.t6 3422.2
R9 minus.n4 minus.t8 3422.2
R10 minus.n10 minus.t11 3422.2
R11 minus.n6 minus.t4 3422.2
R12 minus.n55 minus.t10 3422.2
R13 minus.n53 minus.t2 3422.2
R14 minus.n47 minus.t0 3422.2
R15 minus.n46 minus.t16 3422.2
R16 minus.n44 minus.t7 3422.2
R17 minus.n32 minus.t1 3422.2
R18 minus.n38 minus.t19 3422.2
R19 minus.n34 minus.t14 3422.2
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 69.3793
R47 minus.n15 minus.n4 69.3793
R48 minus.n43 minus.n32 69.3793
R49 minus.n48 minus.n47 69.3793
R50 minus.n25 minus.n24 54.7732
R51 minus.n10 minus.n9 54.7732
R52 minus.n38 minus.n37 54.7732
R53 minus.n54 minus.n53 54.7732
R54 minus.n18 minus.n17 47.4702
R55 minus.n17 minus.n16 47.4702
R56 minus.n45 minus.n44 47.4702
R57 minus.n46 minus.n45 47.4702
R58 minus.n58 minus.n28 43.3717
R59 minus.n26 minus.n25 40.1672
R60 minus.n9 minus.n6 40.1672
R61 minus.n37 minus.n34 40.1672
R62 minus.n55 minus.n54 40.1672
R63 minus.n27 minus.n26 32.8641
R64 minus.n7 minus.n6 32.8641
R65 minus.n35 minus.n34 32.8641
R66 minus.n56 minus.n55 32.8641
R67 minus.n19 minus.n18 25.5611
R68 minus.n16 minus.n15 25.5611
R69 minus.n44 minus.n43 25.5611
R70 minus.n48 minus.n46 25.5611
R71 minus.n24 minus.n23 18.2581
R72 minus.n11 minus.n10 18.2581
R73 minus.n39 minus.n38 18.2581
R74 minus.n53 minus.n52 18.2581
R75 minus.n58 minus.n57 6.56111
R76 minus.n3 minus.n1 3.65202
R77 minus.n12 minus.n4 3.65202
R78 minus.n40 minus.n32 3.65202
R79 minus.n47 minus.n30 3.65202
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 drain_right.n10 drain_right.n8 60.3788
R100 drain_right.n6 drain_right.n4 60.3788
R101 drain_right.n2 drain_right.n0 60.3788
R102 drain_right.n10 drain_right.n9 59.8185
R103 drain_right.n12 drain_right.n11 59.8185
R104 drain_right.n14 drain_right.n13 59.8185
R105 drain_right.n16 drain_right.n15 59.8185
R106 drain_right.n7 drain_right.n3 59.8184
R107 drain_right.n6 drain_right.n5 59.8184
R108 drain_right.n2 drain_right.n1 59.8184
R109 drain_right drain_right.n7 37.3572
R110 drain_right drain_right.n16 6.21356
R111 drain_right.n3 drain_right.t14 1.5005
R112 drain_right.n3 drain_right.t11 1.5005
R113 drain_right.n4 drain_right.t19 1.5005
R114 drain_right.n4 drain_right.t10 1.5005
R115 drain_right.n5 drain_right.t13 1.5005
R116 drain_right.n5 drain_right.t7 1.5005
R117 drain_right.n1 drain_right.t4 1.5005
R118 drain_right.n1 drain_right.t12 1.5005
R119 drain_right.n0 drain_right.t6 1.5005
R120 drain_right.n0 drain_right.t1 1.5005
R121 drain_right.n8 drain_right.t17 1.5005
R122 drain_right.n8 drain_right.t16 1.5005
R123 drain_right.n9 drain_right.t3 1.5005
R124 drain_right.n9 drain_right.t18 1.5005
R125 drain_right.n11 drain_right.t0 1.5005
R126 drain_right.n11 drain_right.t15 1.5005
R127 drain_right.n13 drain_right.t8 1.5005
R128 drain_right.n13 drain_right.t9 1.5005
R129 drain_right.n15 drain_right.t5 1.5005
R130 drain_right.n15 drain_right.t2 1.5005
R131 drain_right.n16 drain_right.n14 0.560845
R132 drain_right.n14 drain_right.n12 0.560845
R133 drain_right.n12 drain_right.n10 0.560845
R134 drain_right.n7 drain_right.n6 0.505499
R135 drain_right.n7 drain_right.n2 0.505499
R136 source.n0 source.t19 44.6397
R137 source.n9 source.t8 44.6396
R138 source.n10 source.t34 44.6396
R139 source.n19 source.t21 44.6396
R140 source.n39 source.t22 44.6395
R141 source.n30 source.t36 44.6395
R142 source.n29 source.t17 44.6395
R143 source.n20 source.t13 44.6395
R144 source.n2 source.n1 43.1397
R145 source.n4 source.n3 43.1397
R146 source.n6 source.n5 43.1397
R147 source.n8 source.n7 43.1397
R148 source.n12 source.n11 43.1397
R149 source.n14 source.n13 43.1397
R150 source.n16 source.n15 43.1397
R151 source.n18 source.n17 43.1397
R152 source.n38 source.n37 43.1396
R153 source.n36 source.n35 43.1396
R154 source.n34 source.n33 43.1396
R155 source.n32 source.n31 43.1396
R156 source.n28 source.n27 43.1396
R157 source.n26 source.n25 43.1396
R158 source.n24 source.n23 43.1396
R159 source.n22 source.n21 43.1396
R160 source.n20 source.n19 27.9087
R161 source.n40 source.n0 22.3656
R162 source.n40 source.n39 5.5436
R163 source.n37 source.t37 1.5005
R164 source.n37 source.t29 1.5005
R165 source.n35 source.t23 1.5005
R166 source.n35 source.t39 1.5005
R167 source.n33 source.t38 1.5005
R168 source.n33 source.t32 1.5005
R169 source.n31 source.t25 1.5005
R170 source.n31 source.t20 1.5005
R171 source.n27 source.t15 1.5005
R172 source.n27 source.t0 1.5005
R173 source.n25 source.t7 1.5005
R174 source.n25 source.t2 1.5005
R175 source.n23 source.t1 1.5005
R176 source.n23 source.t11 1.5005
R177 source.n21 source.t5 1.5005
R178 source.n21 source.t6 1.5005
R179 source.n1 source.t16 1.5005
R180 source.n1 source.t10 1.5005
R181 source.n3 source.t12 1.5005
R182 source.n3 source.t3 1.5005
R183 source.n5 source.t18 1.5005
R184 source.n5 source.t9 1.5005
R185 source.n7 source.t4 1.5005
R186 source.n7 source.t14 1.5005
R187 source.n11 source.t28 1.5005
R188 source.n11 source.t35 1.5005
R189 source.n13 source.t33 1.5005
R190 source.n13 source.t31 1.5005
R191 source.n15 source.t27 1.5005
R192 source.n15 source.t24 1.5005
R193 source.n17 source.t30 1.5005
R194 source.n17 source.t26 1.5005
R195 source.n19 source.n18 0.560845
R196 source.n18 source.n16 0.560845
R197 source.n16 source.n14 0.560845
R198 source.n14 source.n12 0.560845
R199 source.n12 source.n10 0.560845
R200 source.n9 source.n8 0.560845
R201 source.n8 source.n6 0.560845
R202 source.n6 source.n4 0.560845
R203 source.n4 source.n2 0.560845
R204 source.n2 source.n0 0.560845
R205 source.n22 source.n20 0.560845
R206 source.n24 source.n22 0.560845
R207 source.n26 source.n24 0.560845
R208 source.n28 source.n26 0.560845
R209 source.n29 source.n28 0.560845
R210 source.n32 source.n30 0.560845
R211 source.n34 source.n32 0.560845
R212 source.n36 source.n34 0.560845
R213 source.n38 source.n36 0.560845
R214 source.n39 source.n38 0.560845
R215 source.n10 source.n9 0.470328
R216 source.n30 source.n29 0.470328
R217 source source.n40 0.188
R218 plus.n6 plus.t9 3484.28
R219 plus.n27 plus.t12 3484.28
R220 plus.n36 plus.t7 3484.28
R221 plus.n56 plus.t0 3484.28
R222 plus.n5 plus.t18 3422.2
R223 plus.n9 plus.t14 3422.2
R224 plus.n3 plus.t11 3422.2
R225 plus.n15 plus.t19 3422.2
R226 plus.n17 plus.t17 3422.2
R227 plus.n18 plus.t13 3422.2
R228 plus.n24 plus.t8 3422.2
R229 plus.n26 plus.t16 3422.2
R230 plus.n35 plus.t15 3422.2
R231 plus.n39 plus.t2 3422.2
R232 plus.n33 plus.t5 3422.2
R233 plus.n45 plus.t10 3422.2
R234 plus.n47 plus.t1 3422.2
R235 plus.n32 plus.t3 3422.2
R236 plus.n53 plus.t4 3422.2
R237 plus.n55 plus.t6 3422.2
R238 plus.n7 plus.n6 161.489
R239 plus.n37 plus.n36 161.489
R240 plus.n8 plus.n7 161.3
R241 plus.n10 plus.n4 161.3
R242 plus.n12 plus.n11 161.3
R243 plus.n14 plus.n13 161.3
R244 plus.n16 plus.n2 161.3
R245 plus.n20 plus.n19 161.3
R246 plus.n21 plus.n1 161.3
R247 plus.n23 plus.n22 161.3
R248 plus.n25 plus.n0 161.3
R249 plus.n28 plus.n27 161.3
R250 plus.n38 plus.n37 161.3
R251 plus.n40 plus.n34 161.3
R252 plus.n42 plus.n41 161.3
R253 plus.n44 plus.n43 161.3
R254 plus.n46 plus.n31 161.3
R255 plus.n49 plus.n48 161.3
R256 plus.n50 plus.n30 161.3
R257 plus.n52 plus.n51 161.3
R258 plus.n54 plus.n29 161.3
R259 plus.n57 plus.n56 161.3
R260 plus.n11 plus.n10 73.0308
R261 plus.n23 plus.n1 73.0308
R262 plus.n52 plus.n30 73.0308
R263 plus.n41 plus.n40 73.0308
R264 plus.n14 plus.n3 69.3793
R265 plus.n19 plus.n18 69.3793
R266 plus.n48 plus.n32 69.3793
R267 plus.n44 plus.n33 69.3793
R268 plus.n9 plus.n8 54.7732
R269 plus.n25 plus.n24 54.7732
R270 plus.n54 plus.n53 54.7732
R271 plus.n39 plus.n38 54.7732
R272 plus.n16 plus.n15 47.4702
R273 plus.n17 plus.n16 47.4702
R274 plus.n47 plus.n46 47.4702
R275 plus.n46 plus.n45 47.4702
R276 plus.n8 plus.n5 40.1672
R277 plus.n26 plus.n25 40.1672
R278 plus.n55 plus.n54 40.1672
R279 plus.n38 plus.n35 40.1672
R280 plus plus.n57 34.2225
R281 plus.n6 plus.n5 32.8641
R282 plus.n27 plus.n26 32.8641
R283 plus.n56 plus.n55 32.8641
R284 plus.n36 plus.n35 32.8641
R285 plus.n15 plus.n14 25.5611
R286 plus.n19 plus.n17 25.5611
R287 plus.n48 plus.n47 25.5611
R288 plus.n45 plus.n44 25.5611
R289 plus.n10 plus.n9 18.2581
R290 plus.n24 plus.n23 18.2581
R291 plus.n53 plus.n52 18.2581
R292 plus.n40 plus.n39 18.2581
R293 plus plus.n28 15.2353
R294 plus.n11 plus.n3 3.65202
R295 plus.n18 plus.n1 3.65202
R296 plus.n32 plus.n30 3.65202
R297 plus.n41 plus.n33 3.65202
R298 plus.n7 plus.n4 0.189894
R299 plus.n12 plus.n4 0.189894
R300 plus.n13 plus.n12 0.189894
R301 plus.n13 plus.n2 0.189894
R302 plus.n20 plus.n2 0.189894
R303 plus.n21 plus.n20 0.189894
R304 plus.n22 plus.n21 0.189894
R305 plus.n22 plus.n0 0.189894
R306 plus.n28 plus.n0 0.189894
R307 plus.n57 plus.n29 0.189894
R308 plus.n51 plus.n29 0.189894
R309 plus.n51 plus.n50 0.189894
R310 plus.n50 plus.n49 0.189894
R311 plus.n49 plus.n31 0.189894
R312 plus.n43 plus.n31 0.189894
R313 plus.n43 plus.n42 0.189894
R314 plus.n42 plus.n34 0.189894
R315 plus.n37 plus.n34 0.189894
R316 drain_left.n10 drain_left.n8 60.3788
R317 drain_left.n6 drain_left.n4 60.3788
R318 drain_left.n2 drain_left.n0 60.3788
R319 drain_left.n16 drain_left.n15 59.8185
R320 drain_left.n14 drain_left.n13 59.8185
R321 drain_left.n12 drain_left.n11 59.8185
R322 drain_left.n10 drain_left.n9 59.8185
R323 drain_left.n7 drain_left.n3 59.8184
R324 drain_left.n6 drain_left.n5 59.8184
R325 drain_left.n2 drain_left.n1 59.8184
R326 drain_left drain_left.n7 37.9104
R327 drain_left drain_left.n16 6.21356
R328 drain_left.n3 drain_left.t18 1.5005
R329 drain_left.n3 drain_left.t9 1.5005
R330 drain_left.n4 drain_left.t4 1.5005
R331 drain_left.n4 drain_left.t12 1.5005
R332 drain_left.n5 drain_left.t14 1.5005
R333 drain_left.n5 drain_left.t17 1.5005
R334 drain_left.n1 drain_left.t15 1.5005
R335 drain_left.n1 drain_left.t16 1.5005
R336 drain_left.n0 drain_left.t19 1.5005
R337 drain_left.n0 drain_left.t13 1.5005
R338 drain_left.n15 drain_left.t3 1.5005
R339 drain_left.n15 drain_left.t7 1.5005
R340 drain_left.n13 drain_left.t6 1.5005
R341 drain_left.n13 drain_left.t11 1.5005
R342 drain_left.n11 drain_left.t0 1.5005
R343 drain_left.n11 drain_left.t2 1.5005
R344 drain_left.n9 drain_left.t5 1.5005
R345 drain_left.n9 drain_left.t8 1.5005
R346 drain_left.n8 drain_left.t10 1.5005
R347 drain_left.n8 drain_left.t1 1.5005
R348 drain_left.n12 drain_left.n10 0.560845
R349 drain_left.n14 drain_left.n12 0.560845
R350 drain_left.n16 drain_left.n14 0.560845
R351 drain_left.n7 drain_left.n6 0.505499
R352 drain_left.n7 drain_left.n2 0.505499
C0 plus drain_right 0.364841f
C1 drain_left source 61.494003f
C2 drain_left drain_right 1.13563f
C3 plus minus 7.294351f
C4 source drain_right 61.494495f
C5 drain_left minus 0.171338f
C6 source minus 5.79447f
C7 plus drain_left 6.84392f
C8 drain_right minus 6.63324f
C9 plus source 5.80851f
C10 drain_right a_n2146_n4888# 7.92161f
C11 drain_left a_n2146_n4888# 8.234641f
C12 source a_n2146_n4888# 13.193032f
C13 minus a_n2146_n4888# 8.467093f
C14 plus a_n2146_n4888# 11.20389f
C15 drain_left.t19 a_n2146_n4888# 0.676065f
C16 drain_left.t13 a_n2146_n4888# 0.676065f
C17 drain_left.n0 a_n2146_n4888# 4.54227f
C18 drain_left.t15 a_n2146_n4888# 0.676065f
C19 drain_left.t16 a_n2146_n4888# 0.676065f
C20 drain_left.n1 a_n2146_n4888# 4.53901f
C21 drain_left.n2 a_n2146_n4888# 0.684754f
C22 drain_left.t18 a_n2146_n4888# 0.676065f
C23 drain_left.t9 a_n2146_n4888# 0.676065f
C24 drain_left.n3 a_n2146_n4888# 4.53901f
C25 drain_left.t4 a_n2146_n4888# 0.676065f
C26 drain_left.t12 a_n2146_n4888# 0.676065f
C27 drain_left.n4 a_n2146_n4888# 4.54227f
C28 drain_left.t14 a_n2146_n4888# 0.676065f
C29 drain_left.t17 a_n2146_n4888# 0.676065f
C30 drain_left.n5 a_n2146_n4888# 4.53901f
C31 drain_left.n6 a_n2146_n4888# 0.684754f
C32 drain_left.n7 a_n2146_n4888# 2.31928f
C33 drain_left.t10 a_n2146_n4888# 0.676065f
C34 drain_left.t1 a_n2146_n4888# 0.676065f
C35 drain_left.n8 a_n2146_n4888# 4.54227f
C36 drain_left.t5 a_n2146_n4888# 0.676065f
C37 drain_left.t8 a_n2146_n4888# 0.676065f
C38 drain_left.n9 a_n2146_n4888# 4.53901f
C39 drain_left.n10 a_n2146_n4888# 0.688504f
C40 drain_left.t0 a_n2146_n4888# 0.676065f
C41 drain_left.t2 a_n2146_n4888# 0.676065f
C42 drain_left.n11 a_n2146_n4888# 4.53901f
C43 drain_left.n12 a_n2146_n4888# 0.340198f
C44 drain_left.t6 a_n2146_n4888# 0.676065f
C45 drain_left.t11 a_n2146_n4888# 0.676065f
C46 drain_left.n13 a_n2146_n4888# 4.53901f
C47 drain_left.n14 a_n2146_n4888# 0.340198f
C48 drain_left.t3 a_n2146_n4888# 0.676065f
C49 drain_left.t7 a_n2146_n4888# 0.676065f
C50 drain_left.n15 a_n2146_n4888# 4.53901f
C51 drain_left.n16 a_n2146_n4888# 0.575969f
C52 plus.n0 a_n2146_n4888# 0.053549f
C53 plus.t16 a_n2146_n4888# 0.452463f
C54 plus.t8 a_n2146_n4888# 0.452463f
C55 plus.n1 a_n2146_n4888# 0.01859f
C56 plus.n2 a_n2146_n4888# 0.053549f
C57 plus.t17 a_n2146_n4888# 0.452463f
C58 plus.t19 a_n2146_n4888# 0.452463f
C59 plus.t11 a_n2146_n4888# 0.452463f
C60 plus.n3 a_n2146_n4888# 0.176333f
C61 plus.n4 a_n2146_n4888# 0.053549f
C62 plus.t14 a_n2146_n4888# 0.452463f
C63 plus.t18 a_n2146_n4888# 0.452463f
C64 plus.n5 a_n2146_n4888# 0.176333f
C65 plus.t9 a_n2146_n4888# 0.455648f
C66 plus.n6 a_n2146_n4888# 0.198422f
C67 plus.n7 a_n2146_n4888# 0.123524f
C68 plus.n8 a_n2146_n4888# 0.022716f
C69 plus.n9 a_n2146_n4888# 0.176333f
C70 plus.n10 a_n2146_n4888# 0.021891f
C71 plus.n11 a_n2146_n4888# 0.01859f
C72 plus.n12 a_n2146_n4888# 0.053549f
C73 plus.n13 a_n2146_n4888# 0.053549f
C74 plus.n14 a_n2146_n4888# 0.022716f
C75 plus.n15 a_n2146_n4888# 0.176333f
C76 plus.n16 a_n2146_n4888# 0.022716f
C77 plus.n17 a_n2146_n4888# 0.176333f
C78 plus.t13 a_n2146_n4888# 0.452463f
C79 plus.n18 a_n2146_n4888# 0.176333f
C80 plus.n19 a_n2146_n4888# 0.022716f
C81 plus.n20 a_n2146_n4888# 0.053549f
C82 plus.n21 a_n2146_n4888# 0.053549f
C83 plus.n22 a_n2146_n4888# 0.053549f
C84 plus.n23 a_n2146_n4888# 0.021891f
C85 plus.n24 a_n2146_n4888# 0.176333f
C86 plus.n25 a_n2146_n4888# 0.022716f
C87 plus.n26 a_n2146_n4888# 0.176333f
C88 plus.t12 a_n2146_n4888# 0.455648f
C89 plus.n27 a_n2146_n4888# 0.19834f
C90 plus.n28 a_n2146_n4888# 0.82063f
C91 plus.n29 a_n2146_n4888# 0.053549f
C92 plus.t0 a_n2146_n4888# 0.455648f
C93 plus.t6 a_n2146_n4888# 0.452463f
C94 plus.t4 a_n2146_n4888# 0.452463f
C95 plus.n30 a_n2146_n4888# 0.01859f
C96 plus.n31 a_n2146_n4888# 0.053549f
C97 plus.t3 a_n2146_n4888# 0.452463f
C98 plus.n32 a_n2146_n4888# 0.176333f
C99 plus.t1 a_n2146_n4888# 0.452463f
C100 plus.t10 a_n2146_n4888# 0.452463f
C101 plus.t5 a_n2146_n4888# 0.452463f
C102 plus.n33 a_n2146_n4888# 0.176333f
C103 plus.n34 a_n2146_n4888# 0.053549f
C104 plus.t2 a_n2146_n4888# 0.452463f
C105 plus.t15 a_n2146_n4888# 0.452463f
C106 plus.n35 a_n2146_n4888# 0.176333f
C107 plus.t7 a_n2146_n4888# 0.455648f
C108 plus.n36 a_n2146_n4888# 0.198422f
C109 plus.n37 a_n2146_n4888# 0.123524f
C110 plus.n38 a_n2146_n4888# 0.022716f
C111 plus.n39 a_n2146_n4888# 0.176333f
C112 plus.n40 a_n2146_n4888# 0.021891f
C113 plus.n41 a_n2146_n4888# 0.01859f
C114 plus.n42 a_n2146_n4888# 0.053549f
C115 plus.n43 a_n2146_n4888# 0.053549f
C116 plus.n44 a_n2146_n4888# 0.022716f
C117 plus.n45 a_n2146_n4888# 0.176333f
C118 plus.n46 a_n2146_n4888# 0.022716f
C119 plus.n47 a_n2146_n4888# 0.176333f
C120 plus.n48 a_n2146_n4888# 0.022716f
C121 plus.n49 a_n2146_n4888# 0.053549f
C122 plus.n50 a_n2146_n4888# 0.053549f
C123 plus.n51 a_n2146_n4888# 0.053549f
C124 plus.n52 a_n2146_n4888# 0.021891f
C125 plus.n53 a_n2146_n4888# 0.176333f
C126 plus.n54 a_n2146_n4888# 0.022716f
C127 plus.n55 a_n2146_n4888# 0.176333f
C128 plus.n56 a_n2146_n4888# 0.19834f
C129 plus.n57 a_n2146_n4888# 1.97792f
C130 source.t19 a_n2146_n4888# 4.7355f
C131 source.n0 a_n2146_n4888# 1.92263f
C132 source.t16 a_n2146_n4888# 0.582281f
C133 source.t10 a_n2146_n4888# 0.582281f
C134 source.n1 a_n2146_n4888# 3.83181f
C135 source.n2 a_n2146_n4888# 0.3375f
C136 source.t12 a_n2146_n4888# 0.582281f
C137 source.t3 a_n2146_n4888# 0.582281f
C138 source.n3 a_n2146_n4888# 3.83181f
C139 source.n4 a_n2146_n4888# 0.3375f
C140 source.t18 a_n2146_n4888# 0.582281f
C141 source.t9 a_n2146_n4888# 0.582281f
C142 source.n5 a_n2146_n4888# 3.83181f
C143 source.n6 a_n2146_n4888# 0.3375f
C144 source.t4 a_n2146_n4888# 0.582281f
C145 source.t14 a_n2146_n4888# 0.582281f
C146 source.n7 a_n2146_n4888# 3.83181f
C147 source.n8 a_n2146_n4888# 0.3375f
C148 source.t8 a_n2146_n4888# 4.73551f
C149 source.n9 a_n2146_n4888# 0.474811f
C150 source.t34 a_n2146_n4888# 4.73551f
C151 source.n10 a_n2146_n4888# 0.474811f
C152 source.t28 a_n2146_n4888# 0.582281f
C153 source.t35 a_n2146_n4888# 0.582281f
C154 source.n11 a_n2146_n4888# 3.83181f
C155 source.n12 a_n2146_n4888# 0.3375f
C156 source.t33 a_n2146_n4888# 0.582281f
C157 source.t31 a_n2146_n4888# 0.582281f
C158 source.n13 a_n2146_n4888# 3.83181f
C159 source.n14 a_n2146_n4888# 0.3375f
C160 source.t27 a_n2146_n4888# 0.582281f
C161 source.t24 a_n2146_n4888# 0.582281f
C162 source.n15 a_n2146_n4888# 3.83181f
C163 source.n16 a_n2146_n4888# 0.3375f
C164 source.t30 a_n2146_n4888# 0.582281f
C165 source.t26 a_n2146_n4888# 0.582281f
C166 source.n17 a_n2146_n4888# 3.83181f
C167 source.n18 a_n2146_n4888# 0.3375f
C168 source.t21 a_n2146_n4888# 4.73551f
C169 source.n19 a_n2146_n4888# 2.35411f
C170 source.t13 a_n2146_n4888# 4.73549f
C171 source.n20 a_n2146_n4888# 2.35414f
C172 source.t5 a_n2146_n4888# 0.582281f
C173 source.t6 a_n2146_n4888# 0.582281f
C174 source.n21 a_n2146_n4888# 3.83182f
C175 source.n22 a_n2146_n4888# 0.337494f
C176 source.t1 a_n2146_n4888# 0.582281f
C177 source.t11 a_n2146_n4888# 0.582281f
C178 source.n23 a_n2146_n4888# 3.83182f
C179 source.n24 a_n2146_n4888# 0.337494f
C180 source.t7 a_n2146_n4888# 0.582281f
C181 source.t2 a_n2146_n4888# 0.582281f
C182 source.n25 a_n2146_n4888# 3.83182f
C183 source.n26 a_n2146_n4888# 0.337494f
C184 source.t15 a_n2146_n4888# 0.582281f
C185 source.t0 a_n2146_n4888# 0.582281f
C186 source.n27 a_n2146_n4888# 3.83182f
C187 source.n28 a_n2146_n4888# 0.337494f
C188 source.t17 a_n2146_n4888# 4.73549f
C189 source.n29 a_n2146_n4888# 0.474836f
C190 source.t36 a_n2146_n4888# 4.73549f
C191 source.n30 a_n2146_n4888# 0.474836f
C192 source.t25 a_n2146_n4888# 0.582281f
C193 source.t20 a_n2146_n4888# 0.582281f
C194 source.n31 a_n2146_n4888# 3.83182f
C195 source.n32 a_n2146_n4888# 0.337494f
C196 source.t38 a_n2146_n4888# 0.582281f
C197 source.t32 a_n2146_n4888# 0.582281f
C198 source.n33 a_n2146_n4888# 3.83182f
C199 source.n34 a_n2146_n4888# 0.337494f
C200 source.t23 a_n2146_n4888# 0.582281f
C201 source.t39 a_n2146_n4888# 0.582281f
C202 source.n35 a_n2146_n4888# 3.83182f
C203 source.n36 a_n2146_n4888# 0.337494f
C204 source.t37 a_n2146_n4888# 0.582281f
C205 source.t29 a_n2146_n4888# 0.582281f
C206 source.n37 a_n2146_n4888# 3.83182f
C207 source.n38 a_n2146_n4888# 0.337494f
C208 source.t22 a_n2146_n4888# 4.73549f
C209 source.n39 a_n2146_n4888# 0.613179f
C210 source.n40 a_n2146_n4888# 2.18975f
C211 drain_right.t6 a_n2146_n4888# 0.675177f
C212 drain_right.t1 a_n2146_n4888# 0.675177f
C213 drain_right.n0 a_n2146_n4888# 4.53631f
C214 drain_right.t4 a_n2146_n4888# 0.675177f
C215 drain_right.t12 a_n2146_n4888# 0.675177f
C216 drain_right.n1 a_n2146_n4888# 4.53305f
C217 drain_right.n2 a_n2146_n4888# 0.683855f
C218 drain_right.t14 a_n2146_n4888# 0.675177f
C219 drain_right.t11 a_n2146_n4888# 0.675177f
C220 drain_right.n3 a_n2146_n4888# 4.53305f
C221 drain_right.t19 a_n2146_n4888# 0.675177f
C222 drain_right.t10 a_n2146_n4888# 0.675177f
C223 drain_right.n4 a_n2146_n4888# 4.53631f
C224 drain_right.t13 a_n2146_n4888# 0.675177f
C225 drain_right.t7 a_n2146_n4888# 0.675177f
C226 drain_right.n5 a_n2146_n4888# 4.53305f
C227 drain_right.n6 a_n2146_n4888# 0.683855f
C228 drain_right.n7 a_n2146_n4888# 2.25781f
C229 drain_right.t17 a_n2146_n4888# 0.675177f
C230 drain_right.t16 a_n2146_n4888# 0.675177f
C231 drain_right.n8 a_n2146_n4888# 4.5363f
C232 drain_right.t3 a_n2146_n4888# 0.675177f
C233 drain_right.t18 a_n2146_n4888# 0.675177f
C234 drain_right.n9 a_n2146_n4888# 4.53304f
C235 drain_right.n10 a_n2146_n4888# 0.6876f
C236 drain_right.t0 a_n2146_n4888# 0.675177f
C237 drain_right.t15 a_n2146_n4888# 0.675177f
C238 drain_right.n11 a_n2146_n4888# 4.53304f
C239 drain_right.n12 a_n2146_n4888# 0.339751f
C240 drain_right.t8 a_n2146_n4888# 0.675177f
C241 drain_right.t9 a_n2146_n4888# 0.675177f
C242 drain_right.n13 a_n2146_n4888# 4.53304f
C243 drain_right.n14 a_n2146_n4888# 0.339751f
C244 drain_right.t5 a_n2146_n4888# 0.675177f
C245 drain_right.t2 a_n2146_n4888# 0.675177f
C246 drain_right.n15 a_n2146_n4888# 4.53304f
C247 drain_right.n16 a_n2146_n4888# 0.575212f
C248 minus.n0 a_n2146_n4888# 0.052724f
C249 minus.t18 a_n2146_n4888# 0.448628f
C250 minus.t9 a_n2146_n4888# 0.445491f
C251 minus.t13 a_n2146_n4888# 0.445491f
C252 minus.n1 a_n2146_n4888# 0.018303f
C253 minus.n2 a_n2146_n4888# 0.052724f
C254 minus.t12 a_n2146_n4888# 0.445491f
C255 minus.n3 a_n2146_n4888# 0.173616f
C256 minus.t15 a_n2146_n4888# 0.445491f
C257 minus.t6 a_n2146_n4888# 0.445491f
C258 minus.t8 a_n2146_n4888# 0.445491f
C259 minus.n4 a_n2146_n4888# 0.173616f
C260 minus.n5 a_n2146_n4888# 0.052724f
C261 minus.t11 a_n2146_n4888# 0.445491f
C262 minus.t4 a_n2146_n4888# 0.445491f
C263 minus.n6 a_n2146_n4888# 0.173616f
C264 minus.t5 a_n2146_n4888# 0.448628f
C265 minus.n7 a_n2146_n4888# 0.195365f
C266 minus.n8 a_n2146_n4888# 0.121621f
C267 minus.n9 a_n2146_n4888# 0.022366f
C268 minus.n10 a_n2146_n4888# 0.173616f
C269 minus.n11 a_n2146_n4888# 0.021554f
C270 minus.n12 a_n2146_n4888# 0.018303f
C271 minus.n13 a_n2146_n4888# 0.052724f
C272 minus.n14 a_n2146_n4888# 0.052724f
C273 minus.n15 a_n2146_n4888# 0.022366f
C274 minus.n16 a_n2146_n4888# 0.173616f
C275 minus.n17 a_n2146_n4888# 0.022366f
C276 minus.n18 a_n2146_n4888# 0.173616f
C277 minus.n19 a_n2146_n4888# 0.022366f
C278 minus.n20 a_n2146_n4888# 0.052724f
C279 minus.n21 a_n2146_n4888# 0.052724f
C280 minus.n22 a_n2146_n4888# 0.052724f
C281 minus.n23 a_n2146_n4888# 0.021554f
C282 minus.n24 a_n2146_n4888# 0.173616f
C283 minus.n25 a_n2146_n4888# 0.022366f
C284 minus.n26 a_n2146_n4888# 0.173616f
C285 minus.n27 a_n2146_n4888# 0.195284f
C286 minus.n28 a_n2146_n4888# 2.44951f
C287 minus.n29 a_n2146_n4888# 0.052724f
C288 minus.t10 a_n2146_n4888# 0.445491f
C289 minus.t2 a_n2146_n4888# 0.445491f
C290 minus.n30 a_n2146_n4888# 0.018303f
C291 minus.n31 a_n2146_n4888# 0.052724f
C292 minus.t16 a_n2146_n4888# 0.445491f
C293 minus.t7 a_n2146_n4888# 0.445491f
C294 minus.t1 a_n2146_n4888# 0.445491f
C295 minus.n32 a_n2146_n4888# 0.173616f
C296 minus.n33 a_n2146_n4888# 0.052724f
C297 minus.t19 a_n2146_n4888# 0.445491f
C298 minus.t14 a_n2146_n4888# 0.445491f
C299 minus.n34 a_n2146_n4888# 0.173616f
C300 minus.t3 a_n2146_n4888# 0.448628f
C301 minus.n35 a_n2146_n4888# 0.195365f
C302 minus.n36 a_n2146_n4888# 0.121621f
C303 minus.n37 a_n2146_n4888# 0.022366f
C304 minus.n38 a_n2146_n4888# 0.173616f
C305 minus.n39 a_n2146_n4888# 0.021554f
C306 minus.n40 a_n2146_n4888# 0.018303f
C307 minus.n41 a_n2146_n4888# 0.052724f
C308 minus.n42 a_n2146_n4888# 0.052724f
C309 minus.n43 a_n2146_n4888# 0.022366f
C310 minus.n44 a_n2146_n4888# 0.173616f
C311 minus.n45 a_n2146_n4888# 0.022366f
C312 minus.n46 a_n2146_n4888# 0.173616f
C313 minus.t0 a_n2146_n4888# 0.445491f
C314 minus.n47 a_n2146_n4888# 0.173616f
C315 minus.n48 a_n2146_n4888# 0.022366f
C316 minus.n49 a_n2146_n4888# 0.052724f
C317 minus.n50 a_n2146_n4888# 0.052724f
C318 minus.n51 a_n2146_n4888# 0.052724f
C319 minus.n52 a_n2146_n4888# 0.021554f
C320 minus.n53 a_n2146_n4888# 0.173616f
C321 minus.n54 a_n2146_n4888# 0.022366f
C322 minus.n55 a_n2146_n4888# 0.173616f
C323 minus.t17 a_n2146_n4888# 0.448628f
C324 minus.n56 a_n2146_n4888# 0.195284f
C325 minus.n57 a_n2146_n4888# 0.352266f
C326 minus.n58 a_n2146_n4888# 2.91215f
.ends

