* NGSPICE file created from diffpair567.ext - technology: sky130A

.subckt diffpair567 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t7 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X1 drain_right.t6 minus.t1 source.t30 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 drain_right.t1 minus.t2 source.t29 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X3 source.t28 minus.t3 drain_right.t0 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X4 source.t7 plus.t0 drain_left.t15 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X5 drain_left.t14 plus.t1 source.t10 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X6 a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X7 drain_left.t13 plus.t2 source.t0 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X8 source.t13 plus.t3 drain_left.t12 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X9 a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X10 source.t27 minus.t4 drain_right.t5 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source.t2 plus.t4 drain_left.t11 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 drain_right.t4 minus.t5 source.t26 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X13 drain_right.t3 minus.t6 source.t25 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X14 a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X15 source.t24 minus.t7 drain_right.t2 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X16 source.t23 minus.t8 drain_right.t9 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_left.t10 plus.t5 source.t1 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X18 drain_left.t9 plus.t6 source.t15 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X19 source.t4 plus.t7 drain_left.t8 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X20 drain_right.t8 minus.t9 source.t22 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 drain_right.t11 minus.t10 source.t21 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 source.t20 minus.t11 drain_right.t10 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X23 drain_right.t13 minus.t12 source.t19 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X24 drain_left.t7 plus.t8 source.t14 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X25 drain_left.t6 plus.t9 source.t5 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X26 source.t18 minus.t13 drain_right.t12 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 drain_right.t15 minus.t14 source.t17 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X28 source.t8 plus.t10 drain_left.t5 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X29 source.t11 plus.t11 drain_left.t4 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X30 source.t3 plus.t12 drain_left.t3 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X31 a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X32 drain_left.t2 plus.t13 source.t12 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X33 drain_left.t1 plus.t14 source.t6 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X34 source.t16 minus.t15 drain_right.t14 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X35 source.t9 plus.t15 drain_left.t0 a_n1886_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n21 minus.t11 3462.37
R1 minus.n5 minus.t5 3462.37
R2 minus.n44 minus.t2 3462.37
R3 minus.n28 minus.t3 3462.37
R4 minus.n20 minus.t10 3422.2
R5 minus.n1 minus.t13 3422.2
R6 minus.n14 minus.t6 3422.2
R7 minus.n12 minus.t8 3422.2
R8 minus.n3 minus.t9 3422.2
R9 minus.n6 minus.t4 3422.2
R10 minus.n43 minus.t0 3422.2
R11 minus.n24 minus.t14 3422.2
R12 minus.n37 minus.t7 3422.2
R13 minus.n35 minus.t1 3422.2
R14 minus.n26 minus.t15 3422.2
R15 minus.n29 minus.t12 3422.2
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 69.3793
R39 minus.n11 minus.n3 69.3793
R40 minus.n34 minus.n26 69.3793
R41 minus.n38 minus.n24 69.3793
R42 minus.n21 minus.n20 54.7732
R43 minus.n6 minus.n5 54.7732
R44 minus.n29 minus.n28 54.7732
R45 minus.n44 minus.n43 54.7732
R46 minus.n14 minus.n13 47.4702
R47 minus.n13 minus.n12 47.4702
R48 minus.n36 minus.n35 47.4702
R49 minus.n37 minus.n36 47.4702
R50 minus.n46 minus.n22 42.33
R51 minus.n15 minus.n14 25.5611
R52 minus.n12 minus.n11 25.5611
R53 minus.n35 minus.n34 25.5611
R54 minus.n38 minus.n37 25.5611
R55 minus.n20 minus.n19 18.2581
R56 minus.n7 minus.n6 18.2581
R57 minus.n30 minus.n29 18.2581
R58 minus.n43 minus.n42 18.2581
R59 minus.n46 minus.n45 6.50429
R60 minus.n18 minus.n1 3.65202
R61 minus.n8 minus.n3 3.65202
R62 minus.n31 minus.n26 3.65202
R63 minus.n41 minus.n24 3.65202
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 drain_right.n9 drain_right.n7 60.3788
R80 drain_right.n5 drain_right.n3 60.3788
R81 drain_right.n2 drain_right.n0 60.3788
R82 drain_right.n9 drain_right.n8 59.8185
R83 drain_right.n11 drain_right.n10 59.8185
R84 drain_right.n13 drain_right.n12 59.8185
R85 drain_right.n5 drain_right.n4 59.8184
R86 drain_right.n2 drain_right.n1 59.8184
R87 drain_right drain_right.n6 36.5167
R88 drain_right drain_right.n13 6.21356
R89 drain_right.n3 drain_right.t7 1.5005
R90 drain_right.n3 drain_right.t1 1.5005
R91 drain_right.n4 drain_right.t2 1.5005
R92 drain_right.n4 drain_right.t15 1.5005
R93 drain_right.n1 drain_right.t14 1.5005
R94 drain_right.n1 drain_right.t6 1.5005
R95 drain_right.n0 drain_right.t0 1.5005
R96 drain_right.n0 drain_right.t13 1.5005
R97 drain_right.n7 drain_right.t5 1.5005
R98 drain_right.n7 drain_right.t4 1.5005
R99 drain_right.n8 drain_right.t9 1.5005
R100 drain_right.n8 drain_right.t8 1.5005
R101 drain_right.n10 drain_right.t12 1.5005
R102 drain_right.n10 drain_right.t3 1.5005
R103 drain_right.n12 drain_right.t10 1.5005
R104 drain_right.n12 drain_right.t11 1.5005
R105 drain_right.n13 drain_right.n11 0.560845
R106 drain_right.n11 drain_right.n9 0.560845
R107 drain_right.n6 drain_right.n5 0.225326
R108 drain_right.n6 drain_right.n2 0.225326
R109 source.n0 source.t15 44.6397
R110 source.n7 source.t4 44.6396
R111 source.n8 source.t26 44.6396
R112 source.n15 source.t20 44.6396
R113 source.n31 source.t29 44.6395
R114 source.n24 source.t28 44.6395
R115 source.n23 source.t1 44.6395
R116 source.n16 source.t13 44.6395
R117 source.n2 source.n1 43.1397
R118 source.n4 source.n3 43.1397
R119 source.n6 source.n5 43.1397
R120 source.n10 source.n9 43.1397
R121 source.n12 source.n11 43.1397
R122 source.n14 source.n13 43.1397
R123 source.n30 source.n29 43.1396
R124 source.n28 source.n27 43.1396
R125 source.n26 source.n25 43.1396
R126 source.n22 source.n21 43.1396
R127 source.n20 source.n19 43.1396
R128 source.n18 source.n17 43.1396
R129 source.n16 source.n15 27.9087
R130 source.n32 source.n0 22.3656
R131 source.n32 source.n31 5.5436
R132 source.n29 source.t17 1.5005
R133 source.n29 source.t31 1.5005
R134 source.n27 source.t30 1.5005
R135 source.n27 source.t24 1.5005
R136 source.n25 source.t19 1.5005
R137 source.n25 source.t16 1.5005
R138 source.n21 source.t10 1.5005
R139 source.n21 source.t3 1.5005
R140 source.n19 source.t14 1.5005
R141 source.n19 source.t2 1.5005
R142 source.n17 source.t0 1.5005
R143 source.n17 source.t7 1.5005
R144 source.n1 source.t12 1.5005
R145 source.n1 source.t8 1.5005
R146 source.n3 source.t5 1.5005
R147 source.n3 source.t9 1.5005
R148 source.n5 source.t6 1.5005
R149 source.n5 source.t11 1.5005
R150 source.n9 source.t22 1.5005
R151 source.n9 source.t27 1.5005
R152 source.n11 source.t25 1.5005
R153 source.n11 source.t23 1.5005
R154 source.n13 source.t21 1.5005
R155 source.n13 source.t18 1.5005
R156 source.n15 source.n14 0.560845
R157 source.n14 source.n12 0.560845
R158 source.n12 source.n10 0.560845
R159 source.n10 source.n8 0.560845
R160 source.n7 source.n6 0.560845
R161 source.n6 source.n4 0.560845
R162 source.n4 source.n2 0.560845
R163 source.n2 source.n0 0.560845
R164 source.n18 source.n16 0.560845
R165 source.n20 source.n18 0.560845
R166 source.n22 source.n20 0.560845
R167 source.n23 source.n22 0.560845
R168 source.n26 source.n24 0.560845
R169 source.n28 source.n26 0.560845
R170 source.n30 source.n28 0.560845
R171 source.n31 source.n30 0.560845
R172 source.n8 source.n7 0.470328
R173 source.n24 source.n23 0.470328
R174 source source.n32 0.188
R175 plus.n5 plus.t7 3462.37
R176 plus.n21 plus.t6 3462.37
R177 plus.n28 plus.t5 3462.37
R178 plus.n44 plus.t3 3462.37
R179 plus.n6 plus.t14 3422.2
R180 plus.n3 plus.t11 3422.2
R181 plus.n12 plus.t9 3422.2
R182 plus.n14 plus.t15 3422.2
R183 plus.n1 plus.t13 3422.2
R184 plus.n20 plus.t10 3422.2
R185 plus.n29 plus.t12 3422.2
R186 plus.n26 plus.t1 3422.2
R187 plus.n35 plus.t4 3422.2
R188 plus.n37 plus.t8 3422.2
R189 plus.n24 plus.t0 3422.2
R190 plus.n43 plus.t2 3422.2
R191 plus.n5 plus.n4 161.489
R192 plus.n28 plus.n27 161.489
R193 plus.n7 plus.n4 161.3
R194 plus.n9 plus.n8 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n13 plus.n2 161.3
R197 plus.n16 plus.n15 161.3
R198 plus.n18 plus.n17 161.3
R199 plus.n19 plus.n0 161.3
R200 plus.n22 plus.n21 161.3
R201 plus.n30 plus.n27 161.3
R202 plus.n32 plus.n31 161.3
R203 plus.n34 plus.n33 161.3
R204 plus.n36 plus.n25 161.3
R205 plus.n39 plus.n38 161.3
R206 plus.n41 plus.n40 161.3
R207 plus.n42 plus.n23 161.3
R208 plus.n45 plus.n44 161.3
R209 plus.n8 plus.n7 73.0308
R210 plus.n19 plus.n18 73.0308
R211 plus.n42 plus.n41 73.0308
R212 plus.n31 plus.n30 73.0308
R213 plus.n11 plus.n3 69.3793
R214 plus.n15 plus.n1 69.3793
R215 plus.n38 plus.n24 69.3793
R216 plus.n34 plus.n26 69.3793
R217 plus.n6 plus.n5 54.7732
R218 plus.n21 plus.n20 54.7732
R219 plus.n44 plus.n43 54.7732
R220 plus.n29 plus.n28 54.7732
R221 plus.n13 plus.n12 47.4702
R222 plus.n14 plus.n13 47.4702
R223 plus.n37 plus.n36 47.4702
R224 plus.n36 plus.n35 47.4702
R225 plus plus.n45 33.1808
R226 plus.n12 plus.n11 25.5611
R227 plus.n15 plus.n14 25.5611
R228 plus.n38 plus.n37 25.5611
R229 plus.n35 plus.n34 25.5611
R230 plus.n7 plus.n6 18.2581
R231 plus.n20 plus.n19 18.2581
R232 plus.n43 plus.n42 18.2581
R233 plus.n30 plus.n29 18.2581
R234 plus plus.n22 15.1785
R235 plus.n8 plus.n3 3.65202
R236 plus.n18 plus.n1 3.65202
R237 plus.n41 plus.n24 3.65202
R238 plus.n31 plus.n26 3.65202
R239 plus.n9 plus.n4 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n2 0.189894
R242 plus.n16 plus.n2 0.189894
R243 plus.n17 plus.n16 0.189894
R244 plus.n17 plus.n0 0.189894
R245 plus.n22 plus.n0 0.189894
R246 plus.n45 plus.n23 0.189894
R247 plus.n40 plus.n23 0.189894
R248 plus.n40 plus.n39 0.189894
R249 plus.n39 plus.n25 0.189894
R250 plus.n33 plus.n25 0.189894
R251 plus.n33 plus.n32 0.189894
R252 plus.n32 plus.n27 0.189894
R253 drain_left.n9 drain_left.n7 60.3788
R254 drain_left.n5 drain_left.n3 60.3788
R255 drain_left.n2 drain_left.n0 60.3788
R256 drain_left.n13 drain_left.n12 59.8185
R257 drain_left.n11 drain_left.n10 59.8185
R258 drain_left.n9 drain_left.n8 59.8185
R259 drain_left.n5 drain_left.n4 59.8184
R260 drain_left.n2 drain_left.n1 59.8184
R261 drain_left drain_left.n6 37.0699
R262 drain_left drain_left.n13 6.21356
R263 drain_left.n3 drain_left.t3 1.5005
R264 drain_left.n3 drain_left.t10 1.5005
R265 drain_left.n4 drain_left.t11 1.5005
R266 drain_left.n4 drain_left.t14 1.5005
R267 drain_left.n1 drain_left.t15 1.5005
R268 drain_left.n1 drain_left.t7 1.5005
R269 drain_left.n0 drain_left.t12 1.5005
R270 drain_left.n0 drain_left.t13 1.5005
R271 drain_left.n12 drain_left.t5 1.5005
R272 drain_left.n12 drain_left.t9 1.5005
R273 drain_left.n10 drain_left.t0 1.5005
R274 drain_left.n10 drain_left.t2 1.5005
R275 drain_left.n8 drain_left.t4 1.5005
R276 drain_left.n8 drain_left.t6 1.5005
R277 drain_left.n7 drain_left.t8 1.5005
R278 drain_left.n7 drain_left.t1 1.5005
R279 drain_left.n11 drain_left.n9 0.560845
R280 drain_left.n13 drain_left.n11 0.560845
R281 drain_left.n6 drain_left.n5 0.225326
R282 drain_left.n6 drain_left.n2 0.225326
C0 drain_right minus 5.5569f
C1 source drain_left 49.9801f
C2 plus minus 6.97383f
C3 drain_right drain_left 0.96779f
C4 plus drain_left 5.74048f
C5 drain_left minus 0.170952f
C6 source drain_right 49.9805f
C7 plus source 4.69642f
C8 plus drain_right 0.337321f
C9 source minus 4.68238f
C10 drain_right a_n1886_n4888# 7.580821f
C11 drain_left a_n1886_n4888# 7.85589f
C12 source a_n1886_n4888# 13.101635f
C13 minus a_n1886_n4888# 7.506397f
C14 plus a_n1886_n4888# 10.23737f
C15 drain_left.t12 a_n1886_n4888# 0.676254f
C16 drain_left.t13 a_n1886_n4888# 0.676254f
C17 drain_left.n0 a_n1886_n4888# 4.54355f
C18 drain_left.t15 a_n1886_n4888# 0.676254f
C19 drain_left.t7 a_n1886_n4888# 0.676254f
C20 drain_left.n1 a_n1886_n4888# 4.54028f
C21 drain_left.n2 a_n1886_n4888# 0.661067f
C22 drain_left.t3 a_n1886_n4888# 0.676254f
C23 drain_left.t10 a_n1886_n4888# 0.676254f
C24 drain_left.n3 a_n1886_n4888# 4.54355f
C25 drain_left.t11 a_n1886_n4888# 0.676254f
C26 drain_left.t14 a_n1886_n4888# 0.676254f
C27 drain_left.n4 a_n1886_n4888# 4.54028f
C28 drain_left.n5 a_n1886_n4888# 0.661067f
C29 drain_left.n6 a_n1886_n4888# 1.95115f
C30 drain_left.t8 a_n1886_n4888# 0.676254f
C31 drain_left.t1 a_n1886_n4888# 0.676254f
C32 drain_left.n7 a_n1886_n4888# 4.54354f
C33 drain_left.t4 a_n1886_n4888# 0.676254f
C34 drain_left.t6 a_n1886_n4888# 0.676254f
C35 drain_left.n8 a_n1886_n4888# 4.54028f
C36 drain_left.n9 a_n1886_n4888# 0.688697f
C37 drain_left.t0 a_n1886_n4888# 0.676254f
C38 drain_left.t2 a_n1886_n4888# 0.676254f
C39 drain_left.n10 a_n1886_n4888# 4.54028f
C40 drain_left.n11 a_n1886_n4888# 0.340293f
C41 drain_left.t5 a_n1886_n4888# 0.676254f
C42 drain_left.t9 a_n1886_n4888# 0.676254f
C43 drain_left.n12 a_n1886_n4888# 4.54028f
C44 drain_left.n13 a_n1886_n4888# 0.57613f
C45 plus.n0 a_n1886_n4888# 0.055302f
C46 plus.t10 a_n1886_n4888# 0.467269f
C47 plus.t13 a_n1886_n4888# 0.467269f
C48 plus.n1 a_n1886_n4888# 0.182103f
C49 plus.n2 a_n1886_n4888# 0.055302f
C50 plus.t15 a_n1886_n4888# 0.467269f
C51 plus.t9 a_n1886_n4888# 0.467269f
C52 plus.t11 a_n1886_n4888# 0.467269f
C53 plus.n3 a_n1886_n4888# 0.182103f
C54 plus.n4 a_n1886_n4888# 0.11735f
C55 plus.t14 a_n1886_n4888# 0.467269f
C56 plus.t7 a_n1886_n4888# 0.469352f
C57 plus.n5 a_n1886_n4888# 0.200996f
C58 plus.n6 a_n1886_n4888# 0.182103f
C59 plus.n7 a_n1886_n4888# 0.022607f
C60 plus.n8 a_n1886_n4888# 0.019198f
C61 plus.n9 a_n1886_n4888# 0.055302f
C62 plus.n10 a_n1886_n4888# 0.055302f
C63 plus.n11 a_n1886_n4888# 0.02346f
C64 plus.n12 a_n1886_n4888# 0.182103f
C65 plus.n13 a_n1886_n4888# 0.02346f
C66 plus.n14 a_n1886_n4888# 0.182103f
C67 plus.n15 a_n1886_n4888# 0.02346f
C68 plus.n16 a_n1886_n4888# 0.055302f
C69 plus.n17 a_n1886_n4888# 0.055302f
C70 plus.n18 a_n1886_n4888# 0.019198f
C71 plus.n19 a_n1886_n4888# 0.022607f
C72 plus.n20 a_n1886_n4888# 0.182103f
C73 plus.t6 a_n1886_n4888# 0.469352f
C74 plus.n21 a_n1886_n4888# 0.200923f
C75 plus.n22 a_n1886_n4888# 0.840266f
C76 plus.n23 a_n1886_n4888# 0.055302f
C77 plus.t3 a_n1886_n4888# 0.469352f
C78 plus.t2 a_n1886_n4888# 0.467269f
C79 plus.t0 a_n1886_n4888# 0.467269f
C80 plus.n24 a_n1886_n4888# 0.182103f
C81 plus.n25 a_n1886_n4888# 0.055302f
C82 plus.t8 a_n1886_n4888# 0.467269f
C83 plus.t4 a_n1886_n4888# 0.467269f
C84 plus.t1 a_n1886_n4888# 0.467269f
C85 plus.n26 a_n1886_n4888# 0.182103f
C86 plus.n27 a_n1886_n4888# 0.11735f
C87 plus.t12 a_n1886_n4888# 0.467269f
C88 plus.t5 a_n1886_n4888# 0.469352f
C89 plus.n28 a_n1886_n4888# 0.200996f
C90 plus.n29 a_n1886_n4888# 0.182103f
C91 plus.n30 a_n1886_n4888# 0.022607f
C92 plus.n31 a_n1886_n4888# 0.019198f
C93 plus.n32 a_n1886_n4888# 0.055302f
C94 plus.n33 a_n1886_n4888# 0.055302f
C95 plus.n34 a_n1886_n4888# 0.02346f
C96 plus.n35 a_n1886_n4888# 0.182103f
C97 plus.n36 a_n1886_n4888# 0.02346f
C98 plus.n37 a_n1886_n4888# 0.182103f
C99 plus.n38 a_n1886_n4888# 0.02346f
C100 plus.n39 a_n1886_n4888# 0.055302f
C101 plus.n40 a_n1886_n4888# 0.055302f
C102 plus.n41 a_n1886_n4888# 0.019198f
C103 plus.n42 a_n1886_n4888# 0.022607f
C104 plus.n43 a_n1886_n4888# 0.182103f
C105 plus.n44 a_n1886_n4888# 0.200923f
C106 plus.n45 a_n1886_n4888# 1.96092f
C107 source.t15 a_n1886_n4888# 4.57393f
C108 source.n0 a_n1886_n4888# 1.85703f
C109 source.t12 a_n1886_n4888# 0.562414f
C110 source.t8 a_n1886_n4888# 0.562414f
C111 source.n1 a_n1886_n4888# 3.70107f
C112 source.n2 a_n1886_n4888# 0.325985f
C113 source.t5 a_n1886_n4888# 0.562414f
C114 source.t9 a_n1886_n4888# 0.562414f
C115 source.n3 a_n1886_n4888# 3.70107f
C116 source.n4 a_n1886_n4888# 0.325985f
C117 source.t6 a_n1886_n4888# 0.562414f
C118 source.t11 a_n1886_n4888# 0.562414f
C119 source.n5 a_n1886_n4888# 3.70107f
C120 source.n6 a_n1886_n4888# 0.325985f
C121 source.t4 a_n1886_n4888# 4.57394f
C122 source.n7 a_n1886_n4888# 0.458611f
C123 source.t26 a_n1886_n4888# 4.57394f
C124 source.n8 a_n1886_n4888# 0.458611f
C125 source.t22 a_n1886_n4888# 0.562414f
C126 source.t27 a_n1886_n4888# 0.562414f
C127 source.n9 a_n1886_n4888# 3.70107f
C128 source.n10 a_n1886_n4888# 0.325985f
C129 source.t25 a_n1886_n4888# 0.562414f
C130 source.t23 a_n1886_n4888# 0.562414f
C131 source.n11 a_n1886_n4888# 3.70107f
C132 source.n12 a_n1886_n4888# 0.325985f
C133 source.t21 a_n1886_n4888# 0.562414f
C134 source.t18 a_n1886_n4888# 0.562414f
C135 source.n13 a_n1886_n4888# 3.70107f
C136 source.n14 a_n1886_n4888# 0.325985f
C137 source.t20 a_n1886_n4888# 4.57394f
C138 source.n15 a_n1886_n4888# 2.27379f
C139 source.t13 a_n1886_n4888# 4.57392f
C140 source.n16 a_n1886_n4888# 2.27382f
C141 source.t0 a_n1886_n4888# 0.562414f
C142 source.t7 a_n1886_n4888# 0.562414f
C143 source.n17 a_n1886_n4888# 3.70108f
C144 source.n18 a_n1886_n4888# 0.325979f
C145 source.t14 a_n1886_n4888# 0.562414f
C146 source.t2 a_n1886_n4888# 0.562414f
C147 source.n19 a_n1886_n4888# 3.70108f
C148 source.n20 a_n1886_n4888# 0.325979f
C149 source.t10 a_n1886_n4888# 0.562414f
C150 source.t3 a_n1886_n4888# 0.562414f
C151 source.n21 a_n1886_n4888# 3.70108f
C152 source.n22 a_n1886_n4888# 0.325979f
C153 source.t1 a_n1886_n4888# 4.57392f
C154 source.n23 a_n1886_n4888# 0.458635f
C155 source.t28 a_n1886_n4888# 4.57392f
C156 source.n24 a_n1886_n4888# 0.458635f
C157 source.t19 a_n1886_n4888# 0.562414f
C158 source.t16 a_n1886_n4888# 0.562414f
C159 source.n25 a_n1886_n4888# 3.70108f
C160 source.n26 a_n1886_n4888# 0.325979f
C161 source.t30 a_n1886_n4888# 0.562414f
C162 source.t24 a_n1886_n4888# 0.562414f
C163 source.n27 a_n1886_n4888# 3.70108f
C164 source.n28 a_n1886_n4888# 0.325979f
C165 source.t17 a_n1886_n4888# 0.562414f
C166 source.t31 a_n1886_n4888# 0.562414f
C167 source.n29 a_n1886_n4888# 3.70108f
C168 source.n30 a_n1886_n4888# 0.325979f
C169 source.t29 a_n1886_n4888# 4.57392f
C170 source.n31 a_n1886_n4888# 0.592258f
C171 source.n32 a_n1886_n4888# 2.11503f
C172 drain_right.t0 a_n1886_n4888# 0.676382f
C173 drain_right.t13 a_n1886_n4888# 0.676382f
C174 drain_right.n0 a_n1886_n4888# 4.5444f
C175 drain_right.t14 a_n1886_n4888# 0.676382f
C176 drain_right.t6 a_n1886_n4888# 0.676382f
C177 drain_right.n1 a_n1886_n4888# 4.54114f
C178 drain_right.n2 a_n1886_n4888# 0.661191f
C179 drain_right.t7 a_n1886_n4888# 0.676382f
C180 drain_right.t1 a_n1886_n4888# 0.676382f
C181 drain_right.n3 a_n1886_n4888# 4.5444f
C182 drain_right.t2 a_n1886_n4888# 0.676382f
C183 drain_right.t15 a_n1886_n4888# 0.676382f
C184 drain_right.n4 a_n1886_n4888# 4.54114f
C185 drain_right.n5 a_n1886_n4888# 0.661191f
C186 drain_right.n6 a_n1886_n4888# 1.89277f
C187 drain_right.t5 a_n1886_n4888# 0.676382f
C188 drain_right.t4 a_n1886_n4888# 0.676382f
C189 drain_right.n7 a_n1886_n4888# 4.5444f
C190 drain_right.t9 a_n1886_n4888# 0.676382f
C191 drain_right.t8 a_n1886_n4888# 0.676382f
C192 drain_right.n8 a_n1886_n4888# 4.54113f
C193 drain_right.n9 a_n1886_n4888# 0.688827f
C194 drain_right.t12 a_n1886_n4888# 0.676382f
C195 drain_right.t3 a_n1886_n4888# 0.676382f
C196 drain_right.n10 a_n1886_n4888# 4.54113f
C197 drain_right.n11 a_n1886_n4888# 0.340357f
C198 drain_right.t10 a_n1886_n4888# 0.676382f
C199 drain_right.t11 a_n1886_n4888# 0.676382f
C200 drain_right.n12 a_n1886_n4888# 4.54113f
C201 drain_right.n13 a_n1886_n4888# 0.576239f
C202 minus.n0 a_n1886_n4888# 0.054633f
C203 minus.t11 a_n1886_n4888# 0.463674f
C204 minus.t10 a_n1886_n4888# 0.461617f
C205 minus.t13 a_n1886_n4888# 0.461617f
C206 minus.n1 a_n1886_n4888# 0.1799f
C207 minus.n2 a_n1886_n4888# 0.054633f
C208 minus.t6 a_n1886_n4888# 0.461617f
C209 minus.t8 a_n1886_n4888# 0.461617f
C210 minus.t9 a_n1886_n4888# 0.461617f
C211 minus.n3 a_n1886_n4888# 0.1799f
C212 minus.n4 a_n1886_n4888# 0.11593f
C213 minus.t4 a_n1886_n4888# 0.461617f
C214 minus.t5 a_n1886_n4888# 0.463674f
C215 minus.n5 a_n1886_n4888# 0.198564f
C216 minus.n6 a_n1886_n4888# 0.1799f
C217 minus.n7 a_n1886_n4888# 0.022334f
C218 minus.n8 a_n1886_n4888# 0.018966f
C219 minus.n9 a_n1886_n4888# 0.054633f
C220 minus.n10 a_n1886_n4888# 0.054633f
C221 minus.n11 a_n1886_n4888# 0.023176f
C222 minus.n12 a_n1886_n4888# 0.1799f
C223 minus.n13 a_n1886_n4888# 0.023176f
C224 minus.n14 a_n1886_n4888# 0.1799f
C225 minus.n15 a_n1886_n4888# 0.023176f
C226 minus.n16 a_n1886_n4888# 0.054633f
C227 minus.n17 a_n1886_n4888# 0.054633f
C228 minus.n18 a_n1886_n4888# 0.018966f
C229 minus.n19 a_n1886_n4888# 0.022334f
C230 minus.n20 a_n1886_n4888# 0.1799f
C231 minus.n21 a_n1886_n4888# 0.198492f
C232 minus.n22 a_n1886_n4888# 2.44766f
C233 minus.n23 a_n1886_n4888# 0.054633f
C234 minus.t0 a_n1886_n4888# 0.461617f
C235 minus.t14 a_n1886_n4888# 0.461617f
C236 minus.n24 a_n1886_n4888# 0.1799f
C237 minus.n25 a_n1886_n4888# 0.054633f
C238 minus.t7 a_n1886_n4888# 0.461617f
C239 minus.t1 a_n1886_n4888# 0.461617f
C240 minus.t15 a_n1886_n4888# 0.461617f
C241 minus.n26 a_n1886_n4888# 0.1799f
C242 minus.n27 a_n1886_n4888# 0.11593f
C243 minus.t12 a_n1886_n4888# 0.461617f
C244 minus.t3 a_n1886_n4888# 0.463674f
C245 minus.n28 a_n1886_n4888# 0.198564f
C246 minus.n29 a_n1886_n4888# 0.1799f
C247 minus.n30 a_n1886_n4888# 0.022334f
C248 minus.n31 a_n1886_n4888# 0.018966f
C249 minus.n32 a_n1886_n4888# 0.054633f
C250 minus.n33 a_n1886_n4888# 0.054633f
C251 minus.n34 a_n1886_n4888# 0.023176f
C252 minus.n35 a_n1886_n4888# 0.1799f
C253 minus.n36 a_n1886_n4888# 0.023176f
C254 minus.n37 a_n1886_n4888# 0.1799f
C255 minus.n38 a_n1886_n4888# 0.023176f
C256 minus.n39 a_n1886_n4888# 0.054633f
C257 minus.n40 a_n1886_n4888# 0.054633f
C258 minus.n41 a_n1886_n4888# 0.018966f
C259 minus.n42 a_n1886_n4888# 0.022334f
C260 minus.n43 a_n1886_n4888# 0.1799f
C261 minus.t2 a_n1886_n4888# 0.463674f
C262 minus.n44 a_n1886_n4888# 0.198492f
C263 minus.n45 a_n1886_n4888# 0.357727f
C264 minus.n46 a_n1886_n4888# 2.92001f
.ends

