* NGSPICE file created from diffpair203.ext - technology: sky130A

.subckt diffpair203 minus drain_right drain_left source plus
X0 source.t15 minus.t0 drain_right.t0 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X1 source.t14 minus.t1 drain_right.t7 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X2 a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X3 drain_left.t7 plus.t0 source.t6 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X4 a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X5 source.t2 plus.t1 drain_left.t6 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X6 source.t13 minus.t2 drain_right.t6 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 drain_right.t5 minus.t3 source.t12 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X8 drain_left.t5 plus.t2 source.t3 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X9 a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X10 drain_right.t3 minus.t4 source.t11 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X11 drain_left.t4 plus.t3 source.t5 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X12 drain_right.t1 minus.t5 source.t10 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X13 source.t1 plus.t4 drain_left.t3 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X14 source.t4 plus.t5 drain_left.t2 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X15 drain_right.t4 minus.t6 source.t9 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X16 drain_left.t1 plus.t6 source.t0 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X17 source.t8 minus.t7 drain_right.t2 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X18 a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X19 source.t7 plus.t7 drain_left.t0 a_n1546_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
R0 minus.n2 minus.t6 244.149
R1 minus.n10 minus.t2 244.149
R2 minus.n1 minus.t1 223.167
R3 minus.n5 minus.t4 223.167
R4 minus.n6 minus.t7 223.167
R5 minus.n9 minus.t5 223.167
R6 minus.n13 minus.t0 223.167
R7 minus.n14 minus.t3 223.167
R8 minus.n7 minus.n6 161.3
R9 minus.n5 minus.n0 161.3
R10 minus.n4 minus.n3 161.3
R11 minus.n15 minus.n14 161.3
R12 minus.n13 minus.n8 161.3
R13 minus.n12 minus.n11 161.3
R14 minus.n3 minus.n2 70.4033
R15 minus.n11 minus.n10 70.4033
R16 minus.n6 minus.n5 48.2005
R17 minus.n14 minus.n13 48.2005
R18 minus.n16 minus.n7 28.2543
R19 minus.n5 minus.n4 24.1005
R20 minus.n4 minus.n1 24.1005
R21 minus.n12 minus.n9 24.1005
R22 minus.n13 minus.n12 24.1005
R23 minus.n2 minus.n1 20.9576
R24 minus.n10 minus.n9 20.9576
R25 minus.n16 minus.n15 6.5952
R26 minus.n7 minus.n0 0.189894
R27 minus.n3 minus.n0 0.189894
R28 minus.n11 minus.n8 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 drain_right.n5 drain_right.n3 80.4886
R32 drain_right.n2 drain_right.n1 80.0754
R33 drain_right.n2 drain_right.n0 80.0754
R34 drain_right.n5 drain_right.n4 79.7731
R35 drain_right drain_right.n2 22.5
R36 drain_right.n1 drain_right.t0 6.6005
R37 drain_right.n1 drain_right.t5 6.6005
R38 drain_right.n0 drain_right.t6 6.6005
R39 drain_right.n0 drain_right.t1 6.6005
R40 drain_right.n3 drain_right.t7 6.6005
R41 drain_right.n3 drain_right.t4 6.6005
R42 drain_right.n4 drain_right.t2 6.6005
R43 drain_right.n4 drain_right.t3 6.6005
R44 drain_right drain_right.n5 6.36873
R45 source.n0 source.t5 69.6943
R46 source.n3 source.t2 69.6943
R47 source.n4 source.t9 69.6943
R48 source.n7 source.t8 69.6943
R49 source.n15 source.t12 69.6942
R50 source.n12 source.t13 69.6942
R51 source.n11 source.t3 69.6942
R52 source.n8 source.t4 69.6942
R53 source.n2 source.n1 63.0943
R54 source.n6 source.n5 63.0943
R55 source.n14 source.n13 63.0942
R56 source.n10 source.n9 63.0942
R57 source.n8 source.n7 15.1851
R58 source.n16 source.n0 9.56437
R59 source.n13 source.t10 6.6005
R60 source.n13 source.t15 6.6005
R61 source.n9 source.t6 6.6005
R62 source.n9 source.t1 6.6005
R63 source.n1 source.t0 6.6005
R64 source.n1 source.t7 6.6005
R65 source.n5 source.t11 6.6005
R66 source.n5 source.t14 6.6005
R67 source.n16 source.n15 5.62119
R68 source.n7 source.n6 0.716017
R69 source.n6 source.n4 0.716017
R70 source.n3 source.n2 0.716017
R71 source.n2 source.n0 0.716017
R72 source.n10 source.n8 0.716017
R73 source.n11 source.n10 0.716017
R74 source.n14 source.n12 0.716017
R75 source.n15 source.n14 0.716017
R76 source.n4 source.n3 0.470328
R77 source.n12 source.n11 0.470328
R78 source source.n16 0.188
R79 plus.n2 plus.t1 244.149
R80 plus.n10 plus.t2 244.149
R81 plus.n6 plus.t3 223.167
R82 plus.n5 plus.t7 223.167
R83 plus.n1 plus.t6 223.167
R84 plus.n14 plus.t5 223.167
R85 plus.n13 plus.t0 223.167
R86 plus.n9 plus.t4 223.167
R87 plus.n4 plus.n3 161.3
R88 plus.n5 plus.n0 161.3
R89 plus.n7 plus.n6 161.3
R90 plus.n12 plus.n11 161.3
R91 plus.n13 plus.n8 161.3
R92 plus.n15 plus.n14 161.3
R93 plus.n3 plus.n2 70.4033
R94 plus.n11 plus.n10 70.4033
R95 plus.n6 plus.n5 48.2005
R96 plus.n14 plus.n13 48.2005
R97 plus plus.n15 25.5445
R98 plus.n4 plus.n1 24.1005
R99 plus.n5 plus.n4 24.1005
R100 plus.n13 plus.n12 24.1005
R101 plus.n12 plus.n9 24.1005
R102 plus.n2 plus.n1 20.9576
R103 plus.n10 plus.n9 20.9576
R104 plus plus.n7 8.83005
R105 plus.n3 plus.n0 0.189894
R106 plus.n7 plus.n0 0.189894
R107 plus.n15 plus.n8 0.189894
R108 plus.n11 plus.n8 0.189894
R109 drain_left.n5 drain_left.n3 80.4886
R110 drain_left.n2 drain_left.n1 80.0754
R111 drain_left.n2 drain_left.n0 80.0754
R112 drain_left.n5 drain_left.n4 79.7731
R113 drain_left drain_left.n2 23.0532
R114 drain_left.n1 drain_left.t3 6.6005
R115 drain_left.n1 drain_left.t5 6.6005
R116 drain_left.n0 drain_left.t2 6.6005
R117 drain_left.n0 drain_left.t7 6.6005
R118 drain_left.n4 drain_left.t0 6.6005
R119 drain_left.n4 drain_left.t4 6.6005
R120 drain_left.n3 drain_left.t6 6.6005
R121 drain_left.n3 drain_left.t1 6.6005
R122 drain_left drain_left.n5 6.36873
C0 minus plus 3.41149f
C1 source minus 1.54696f
C2 drain_right plus 0.307597f
C3 source drain_right 4.76276f
C4 source plus 1.56095f
C5 minus drain_left 0.176136f
C6 drain_right drain_left 0.727126f
C7 drain_left plus 1.57131f
C8 source drain_left 4.76226f
C9 minus drain_right 1.42329f
C10 drain_right a_n1546_n1488# 3.36561f
C11 drain_left a_n1546_n1488# 3.5638f
C12 source a_n1546_n1488# 3.555765f
C13 minus a_n1546_n1488# 5.237386f
C14 plus a_n1546_n1488# 5.826118f
C15 drain_left.t2 a_n1546_n1488# 0.049444f
C16 drain_left.t7 a_n1546_n1488# 0.049444f
C17 drain_left.n0 a_n1546_n1488# 0.357511f
C18 drain_left.t3 a_n1546_n1488# 0.049444f
C19 drain_left.t5 a_n1546_n1488# 0.049444f
C20 drain_left.n1 a_n1546_n1488# 0.357511f
C21 drain_left.n2 a_n1546_n1488# 1.06798f
C22 drain_left.t6 a_n1546_n1488# 0.049444f
C23 drain_left.t1 a_n1546_n1488# 0.049444f
C24 drain_left.n3 a_n1546_n1488# 0.359f
C25 drain_left.t0 a_n1546_n1488# 0.049444f
C26 drain_left.t4 a_n1546_n1488# 0.049444f
C27 drain_left.n4 a_n1546_n1488# 0.356586f
C28 drain_left.n5 a_n1546_n1488# 0.711414f
C29 plus.n0 a_n1546_n1488# 0.027214f
C30 plus.t3 a_n1546_n1488# 0.122406f
C31 plus.t7 a_n1546_n1488# 0.122406f
C32 plus.t6 a_n1546_n1488# 0.122406f
C33 plus.n1 a_n1546_n1488# 0.076184f
C34 plus.t1 a_n1546_n1488# 0.128719f
C35 plus.n2 a_n1546_n1488# 0.067313f
C36 plus.n3 a_n1546_n1488# 0.089652f
C37 plus.n4 a_n1546_n1488# 0.006175f
C38 plus.n5 a_n1546_n1488# 0.076184f
C39 plus.n6 a_n1546_n1488# 0.073416f
C40 plus.n7 a_n1546_n1488# 0.209682f
C41 plus.n8 a_n1546_n1488# 0.027214f
C42 plus.t5 a_n1546_n1488# 0.122406f
C43 plus.t0 a_n1546_n1488# 0.122406f
C44 plus.t4 a_n1546_n1488# 0.122406f
C45 plus.n9 a_n1546_n1488# 0.076184f
C46 plus.t2 a_n1546_n1488# 0.128719f
C47 plus.n10 a_n1546_n1488# 0.067313f
C48 plus.n11 a_n1546_n1488# 0.089652f
C49 plus.n12 a_n1546_n1488# 0.006175f
C50 plus.n13 a_n1546_n1488# 0.076184f
C51 plus.n14 a_n1546_n1488# 0.073416f
C52 plus.n15 a_n1546_n1488# 0.604239f
C53 source.t5 a_n1546_n1488# 0.375563f
C54 source.n0 a_n1546_n1488# 0.531035f
C55 source.t0 a_n1546_n1488# 0.045228f
C56 source.t7 a_n1546_n1488# 0.045228f
C57 source.n1 a_n1546_n1488# 0.286769f
C58 source.n2 a_n1546_n1488# 0.254163f
C59 source.t2 a_n1546_n1488# 0.375563f
C60 source.n3 a_n1546_n1488# 0.273614f
C61 source.t9 a_n1546_n1488# 0.375563f
C62 source.n4 a_n1546_n1488# 0.273614f
C63 source.t11 a_n1546_n1488# 0.045228f
C64 source.t14 a_n1546_n1488# 0.045228f
C65 source.n5 a_n1546_n1488# 0.286769f
C66 source.n6 a_n1546_n1488# 0.254163f
C67 source.t8 a_n1546_n1488# 0.375563f
C68 source.n7 a_n1546_n1488# 0.732452f
C69 source.t4 a_n1546_n1488# 0.375561f
C70 source.n8 a_n1546_n1488# 0.732453f
C71 source.t6 a_n1546_n1488# 0.045228f
C72 source.t1 a_n1546_n1488# 0.045228f
C73 source.n9 a_n1546_n1488# 0.286767f
C74 source.n10 a_n1546_n1488# 0.254165f
C75 source.t3 a_n1546_n1488# 0.375561f
C76 source.n11 a_n1546_n1488# 0.273616f
C77 source.t13 a_n1546_n1488# 0.375561f
C78 source.n12 a_n1546_n1488# 0.273616f
C79 source.t10 a_n1546_n1488# 0.045228f
C80 source.t15 a_n1546_n1488# 0.045228f
C81 source.n13 a_n1546_n1488# 0.286767f
C82 source.n14 a_n1546_n1488# 0.254165f
C83 source.t12 a_n1546_n1488# 0.375561f
C84 source.n15 a_n1546_n1488# 0.389733f
C85 source.n16 a_n1546_n1488# 0.557706f
C86 drain_right.t6 a_n1546_n1488# 0.050299f
C87 drain_right.t1 a_n1546_n1488# 0.050299f
C88 drain_right.n0 a_n1546_n1488# 0.363693f
C89 drain_right.t0 a_n1546_n1488# 0.050299f
C90 drain_right.t5 a_n1546_n1488# 0.050299f
C91 drain_right.n1 a_n1546_n1488# 0.363693f
C92 drain_right.n2 a_n1546_n1488# 1.04424f
C93 drain_right.t7 a_n1546_n1488# 0.050299f
C94 drain_right.t4 a_n1546_n1488# 0.050299f
C95 drain_right.n3 a_n1546_n1488# 0.365208f
C96 drain_right.t2 a_n1546_n1488# 0.050299f
C97 drain_right.t3 a_n1546_n1488# 0.050299f
C98 drain_right.n4 a_n1546_n1488# 0.362752f
C99 drain_right.n5 a_n1546_n1488# 0.723716f
C100 minus.n0 a_n1546_n1488# 0.02678f
C101 minus.t1 a_n1546_n1488# 0.120456f
C102 minus.n1 a_n1546_n1488# 0.074971f
C103 minus.t6 a_n1546_n1488# 0.126668f
C104 minus.n2 a_n1546_n1488# 0.066241f
C105 minus.n3 a_n1546_n1488# 0.088224f
C106 minus.n4 a_n1546_n1488# 0.006077f
C107 minus.t4 a_n1546_n1488# 0.120456f
C108 minus.n5 a_n1546_n1488# 0.074971f
C109 minus.t7 a_n1546_n1488# 0.120456f
C110 minus.n6 a_n1546_n1488# 0.072246f
C111 minus.n7 a_n1546_n1488# 0.630385f
C112 minus.n8 a_n1546_n1488# 0.02678f
C113 minus.t5 a_n1546_n1488# 0.120456f
C114 minus.n9 a_n1546_n1488# 0.074971f
C115 minus.t2 a_n1546_n1488# 0.126668f
C116 minus.n10 a_n1546_n1488# 0.066241f
C117 minus.n11 a_n1546_n1488# 0.088224f
C118 minus.n12 a_n1546_n1488# 0.006077f
C119 minus.t0 a_n1546_n1488# 0.120456f
C120 minus.n13 a_n1546_n1488# 0.074971f
C121 minus.t3 a_n1546_n1488# 0.120456f
C122 minus.n14 a_n1546_n1488# 0.072246f
C123 minus.n15 a_n1546_n1488# 0.181061f
C124 minus.n16 a_n1546_n1488# 0.775873f
.ends

