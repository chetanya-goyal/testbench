* NGSPICE file created from diffpair272.ext - technology: sky130A

.subckt diffpair272 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t11 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t0 plus.t0 drain_left.t5 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X3 drain_left.t4 plus.t1 source.t4 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X4 a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X5 source.t8 minus.t1 drain_right.t4 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X6 a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X7 a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X8 source.t3 plus.t2 drain_left.t3 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X9 drain_left.t2 plus.t3 source.t2 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X10 drain_left.t1 plus.t4 source.t1 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X11 drain_right.t3 minus.t2 source.t10 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X12 drain_right.t2 minus.t3 source.t9 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X13 drain_right.t1 minus.t4 source.t6 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X14 drain_left.t0 plus.t5 source.t5 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X15 source.t7 minus.t5 drain_right.t0 a_n1220_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n2 minus.t0 641.937
R1 minus.n0 minus.t2 641.937
R2 minus.n6 minus.t3 641.937
R3 minus.n4 minus.t4 641.937
R4 minus.n1 minus.t5 586.433
R5 minus.n5 minus.t1 586.433
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 29.2297
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 source.n130 source.n104 289.615
R18 source.n96 source.n70 289.615
R19 source.n26 source.n0 289.615
R20 source.n60 source.n34 289.615
R21 source.n115 source.n114 185
R22 source.n112 source.n111 185
R23 source.n121 source.n120 185
R24 source.n123 source.n122 185
R25 source.n108 source.n107 185
R26 source.n129 source.n128 185
R27 source.n131 source.n130 185
R28 source.n81 source.n80 185
R29 source.n78 source.n77 185
R30 source.n87 source.n86 185
R31 source.n89 source.n88 185
R32 source.n74 source.n73 185
R33 source.n95 source.n94 185
R34 source.n97 source.n96 185
R35 source.n27 source.n26 185
R36 source.n25 source.n24 185
R37 source.n4 source.n3 185
R38 source.n19 source.n18 185
R39 source.n17 source.n16 185
R40 source.n8 source.n7 185
R41 source.n11 source.n10 185
R42 source.n61 source.n60 185
R43 source.n59 source.n58 185
R44 source.n38 source.n37 185
R45 source.n53 source.n52 185
R46 source.n51 source.n50 185
R47 source.n42 source.n41 185
R48 source.n45 source.n44 185
R49 source.t9 source.n113 147.661
R50 source.t2 source.n79 147.661
R51 source.t5 source.n9 147.661
R52 source.t10 source.n43 147.661
R53 source.n114 source.n111 104.615
R54 source.n121 source.n111 104.615
R55 source.n122 source.n121 104.615
R56 source.n122 source.n107 104.615
R57 source.n129 source.n107 104.615
R58 source.n130 source.n129 104.615
R59 source.n80 source.n77 104.615
R60 source.n87 source.n77 104.615
R61 source.n88 source.n87 104.615
R62 source.n88 source.n73 104.615
R63 source.n95 source.n73 104.615
R64 source.n96 source.n95 104.615
R65 source.n26 source.n25 104.615
R66 source.n25 source.n3 104.615
R67 source.n18 source.n3 104.615
R68 source.n18 source.n17 104.615
R69 source.n17 source.n7 104.615
R70 source.n10 source.n7 104.615
R71 source.n60 source.n59 104.615
R72 source.n59 source.n37 104.615
R73 source.n52 source.n37 104.615
R74 source.n52 source.n51 104.615
R75 source.n51 source.n41 104.615
R76 source.n44 source.n41 104.615
R77 source.n114 source.t9 52.3082
R78 source.n80 source.t2 52.3082
R79 source.n10 source.t5 52.3082
R80 source.n44 source.t10 52.3082
R81 source.n33 source.n32 50.512
R82 source.n67 source.n66 50.512
R83 source.n103 source.n102 50.5119
R84 source.n69 source.n68 50.5119
R85 source.n135 source.n134 32.1853
R86 source.n101 source.n100 32.1853
R87 source.n31 source.n30 32.1853
R88 source.n65 source.n64 32.1853
R89 source.n69 source.n67 17.8285
R90 source.n115 source.n113 15.6674
R91 source.n81 source.n79 15.6674
R92 source.n11 source.n9 15.6674
R93 source.n45 source.n43 15.6674
R94 source.n116 source.n112 12.8005
R95 source.n82 source.n78 12.8005
R96 source.n12 source.n8 12.8005
R97 source.n46 source.n42 12.8005
R98 source.n120 source.n119 12.0247
R99 source.n86 source.n85 12.0247
R100 source.n16 source.n15 12.0247
R101 source.n50 source.n49 12.0247
R102 source.n136 source.n31 11.7509
R103 source.n123 source.n110 11.249
R104 source.n89 source.n76 11.249
R105 source.n19 source.n6 11.249
R106 source.n53 source.n40 11.249
R107 source.n124 source.n108 10.4732
R108 source.n90 source.n74 10.4732
R109 source.n20 source.n4 10.4732
R110 source.n54 source.n38 10.4732
R111 source.n128 source.n127 9.69747
R112 source.n94 source.n93 9.69747
R113 source.n24 source.n23 9.69747
R114 source.n58 source.n57 9.69747
R115 source.n134 source.n133 9.45567
R116 source.n100 source.n99 9.45567
R117 source.n30 source.n29 9.45567
R118 source.n64 source.n63 9.45567
R119 source.n133 source.n132 9.3005
R120 source.n106 source.n105 9.3005
R121 source.n127 source.n126 9.3005
R122 source.n125 source.n124 9.3005
R123 source.n110 source.n109 9.3005
R124 source.n119 source.n118 9.3005
R125 source.n117 source.n116 9.3005
R126 source.n99 source.n98 9.3005
R127 source.n72 source.n71 9.3005
R128 source.n93 source.n92 9.3005
R129 source.n91 source.n90 9.3005
R130 source.n76 source.n75 9.3005
R131 source.n85 source.n84 9.3005
R132 source.n83 source.n82 9.3005
R133 source.n29 source.n28 9.3005
R134 source.n2 source.n1 9.3005
R135 source.n23 source.n22 9.3005
R136 source.n21 source.n20 9.3005
R137 source.n6 source.n5 9.3005
R138 source.n15 source.n14 9.3005
R139 source.n13 source.n12 9.3005
R140 source.n63 source.n62 9.3005
R141 source.n36 source.n35 9.3005
R142 source.n57 source.n56 9.3005
R143 source.n55 source.n54 9.3005
R144 source.n40 source.n39 9.3005
R145 source.n49 source.n48 9.3005
R146 source.n47 source.n46 9.3005
R147 source.n131 source.n106 8.92171
R148 source.n97 source.n72 8.92171
R149 source.n27 source.n2 8.92171
R150 source.n61 source.n36 8.92171
R151 source.n132 source.n104 8.14595
R152 source.n98 source.n70 8.14595
R153 source.n28 source.n0 8.14595
R154 source.n62 source.n34 8.14595
R155 source.n134 source.n104 5.81868
R156 source.n100 source.n70 5.81868
R157 source.n30 source.n0 5.81868
R158 source.n64 source.n34 5.81868
R159 source.n136 source.n135 5.53498
R160 source.n132 source.n131 5.04292
R161 source.n98 source.n97 5.04292
R162 source.n28 source.n27 5.04292
R163 source.n62 source.n61 5.04292
R164 source.n117 source.n113 4.38594
R165 source.n83 source.n79 4.38594
R166 source.n13 source.n9 4.38594
R167 source.n47 source.n43 4.38594
R168 source.n128 source.n106 4.26717
R169 source.n94 source.n72 4.26717
R170 source.n24 source.n2 4.26717
R171 source.n58 source.n36 4.26717
R172 source.n127 source.n108 3.49141
R173 source.n93 source.n74 3.49141
R174 source.n23 source.n4 3.49141
R175 source.n57 source.n38 3.49141
R176 source.n102 source.t6 3.3005
R177 source.n102 source.t8 3.3005
R178 source.n68 source.t1 3.3005
R179 source.n68 source.t0 3.3005
R180 source.n32 source.t4 3.3005
R181 source.n32 source.t3 3.3005
R182 source.n66 source.t11 3.3005
R183 source.n66 source.t7 3.3005
R184 source.n124 source.n123 2.71565
R185 source.n90 source.n89 2.71565
R186 source.n20 source.n19 2.71565
R187 source.n54 source.n53 2.71565
R188 source.n120 source.n110 1.93989
R189 source.n86 source.n76 1.93989
R190 source.n16 source.n6 1.93989
R191 source.n50 source.n40 1.93989
R192 source.n119 source.n112 1.16414
R193 source.n85 source.n78 1.16414
R194 source.n15 source.n8 1.16414
R195 source.n49 source.n42 1.16414
R196 source.n65 source.n33 0.741879
R197 source.n103 source.n101 0.741879
R198 source.n67 source.n65 0.543603
R199 source.n33 source.n31 0.543603
R200 source.n101 source.n69 0.543603
R201 source.n135 source.n103 0.543603
R202 source.n116 source.n115 0.388379
R203 source.n82 source.n81 0.388379
R204 source.n12 source.n11 0.388379
R205 source.n46 source.n45 0.388379
R206 source source.n136 0.188
R207 source.n118 source.n117 0.155672
R208 source.n118 source.n109 0.155672
R209 source.n125 source.n109 0.155672
R210 source.n126 source.n125 0.155672
R211 source.n126 source.n105 0.155672
R212 source.n133 source.n105 0.155672
R213 source.n84 source.n83 0.155672
R214 source.n84 source.n75 0.155672
R215 source.n91 source.n75 0.155672
R216 source.n92 source.n91 0.155672
R217 source.n92 source.n71 0.155672
R218 source.n99 source.n71 0.155672
R219 source.n29 source.n1 0.155672
R220 source.n22 source.n1 0.155672
R221 source.n22 source.n21 0.155672
R222 source.n21 source.n5 0.155672
R223 source.n14 source.n5 0.155672
R224 source.n14 source.n13 0.155672
R225 source.n63 source.n35 0.155672
R226 source.n56 source.n35 0.155672
R227 source.n56 source.n55 0.155672
R228 source.n55 source.n39 0.155672
R229 source.n48 source.n39 0.155672
R230 source.n48 source.n47 0.155672
R231 drain_right.n26 drain_right.n0 289.615
R232 drain_right.n60 drain_right.n34 289.615
R233 drain_right.n11 drain_right.n10 185
R234 drain_right.n8 drain_right.n7 185
R235 drain_right.n17 drain_right.n16 185
R236 drain_right.n19 drain_right.n18 185
R237 drain_right.n4 drain_right.n3 185
R238 drain_right.n25 drain_right.n24 185
R239 drain_right.n27 drain_right.n26 185
R240 drain_right.n61 drain_right.n60 185
R241 drain_right.n59 drain_right.n58 185
R242 drain_right.n38 drain_right.n37 185
R243 drain_right.n53 drain_right.n52 185
R244 drain_right.n51 drain_right.n50 185
R245 drain_right.n42 drain_right.n41 185
R246 drain_right.n45 drain_right.n44 185
R247 drain_right.t1 drain_right.n9 147.661
R248 drain_right.t5 drain_right.n43 147.661
R249 drain_right.n10 drain_right.n7 104.615
R250 drain_right.n17 drain_right.n7 104.615
R251 drain_right.n18 drain_right.n17 104.615
R252 drain_right.n18 drain_right.n3 104.615
R253 drain_right.n25 drain_right.n3 104.615
R254 drain_right.n26 drain_right.n25 104.615
R255 drain_right.n60 drain_right.n59 104.615
R256 drain_right.n59 drain_right.n37 104.615
R257 drain_right.n52 drain_right.n37 104.615
R258 drain_right.n52 drain_right.n51 104.615
R259 drain_right.n51 drain_right.n41 104.615
R260 drain_right.n44 drain_right.n41 104.615
R261 drain_right.n65 drain_right.n33 67.7338
R262 drain_right.n32 drain_right.n31 67.2711
R263 drain_right.n10 drain_right.t1 52.3082
R264 drain_right.n44 drain_right.t5 52.3082
R265 drain_right.n32 drain_right.n30 49.2161
R266 drain_right.n65 drain_right.n64 48.8641
R267 drain_right drain_right.n32 23.7619
R268 drain_right.n11 drain_right.n9 15.6674
R269 drain_right.n45 drain_right.n43 15.6674
R270 drain_right.n12 drain_right.n8 12.8005
R271 drain_right.n46 drain_right.n42 12.8005
R272 drain_right.n16 drain_right.n15 12.0247
R273 drain_right.n50 drain_right.n49 12.0247
R274 drain_right.n19 drain_right.n6 11.249
R275 drain_right.n53 drain_right.n40 11.249
R276 drain_right.n20 drain_right.n4 10.4732
R277 drain_right.n54 drain_right.n38 10.4732
R278 drain_right.n24 drain_right.n23 9.69747
R279 drain_right.n58 drain_right.n57 9.69747
R280 drain_right.n30 drain_right.n29 9.45567
R281 drain_right.n64 drain_right.n63 9.45567
R282 drain_right.n29 drain_right.n28 9.3005
R283 drain_right.n2 drain_right.n1 9.3005
R284 drain_right.n23 drain_right.n22 9.3005
R285 drain_right.n21 drain_right.n20 9.3005
R286 drain_right.n6 drain_right.n5 9.3005
R287 drain_right.n15 drain_right.n14 9.3005
R288 drain_right.n13 drain_right.n12 9.3005
R289 drain_right.n63 drain_right.n62 9.3005
R290 drain_right.n36 drain_right.n35 9.3005
R291 drain_right.n57 drain_right.n56 9.3005
R292 drain_right.n55 drain_right.n54 9.3005
R293 drain_right.n40 drain_right.n39 9.3005
R294 drain_right.n49 drain_right.n48 9.3005
R295 drain_right.n47 drain_right.n46 9.3005
R296 drain_right.n27 drain_right.n2 8.92171
R297 drain_right.n61 drain_right.n36 8.92171
R298 drain_right.n28 drain_right.n0 8.14595
R299 drain_right.n62 drain_right.n34 8.14595
R300 drain_right drain_right.n65 5.92477
R301 drain_right.n30 drain_right.n0 5.81868
R302 drain_right.n64 drain_right.n34 5.81868
R303 drain_right.n28 drain_right.n27 5.04292
R304 drain_right.n62 drain_right.n61 5.04292
R305 drain_right.n13 drain_right.n9 4.38594
R306 drain_right.n47 drain_right.n43 4.38594
R307 drain_right.n24 drain_right.n2 4.26717
R308 drain_right.n58 drain_right.n36 4.26717
R309 drain_right.n23 drain_right.n4 3.49141
R310 drain_right.n57 drain_right.n38 3.49141
R311 drain_right.n31 drain_right.t4 3.3005
R312 drain_right.n31 drain_right.t2 3.3005
R313 drain_right.n33 drain_right.t0 3.3005
R314 drain_right.n33 drain_right.t3 3.3005
R315 drain_right.n20 drain_right.n19 2.71565
R316 drain_right.n54 drain_right.n53 2.71565
R317 drain_right.n16 drain_right.n6 1.93989
R318 drain_right.n50 drain_right.n40 1.93989
R319 drain_right.n15 drain_right.n8 1.16414
R320 drain_right.n49 drain_right.n42 1.16414
R321 drain_right.n12 drain_right.n11 0.388379
R322 drain_right.n46 drain_right.n45 0.388379
R323 drain_right.n14 drain_right.n13 0.155672
R324 drain_right.n14 drain_right.n5 0.155672
R325 drain_right.n21 drain_right.n5 0.155672
R326 drain_right.n22 drain_right.n21 0.155672
R327 drain_right.n22 drain_right.n1 0.155672
R328 drain_right.n29 drain_right.n1 0.155672
R329 drain_right.n63 drain_right.n35 0.155672
R330 drain_right.n56 drain_right.n35 0.155672
R331 drain_right.n56 drain_right.n55 0.155672
R332 drain_right.n55 drain_right.n39 0.155672
R333 drain_right.n48 drain_right.n39 0.155672
R334 drain_right.n48 drain_right.n47 0.155672
R335 plus.n0 plus.t1 641.937
R336 plus.n2 plus.t5 641.937
R337 plus.n4 plus.t3 641.937
R338 plus.n6 plus.t4 641.937
R339 plus.n1 plus.t2 586.433
R340 plus.n5 plus.t0 586.433
R341 plus.n3 plus.n0 161.489
R342 plus.n7 plus.n4 161.489
R343 plus.n3 plus.n2 161.3
R344 plus.n7 plus.n6 161.3
R345 plus.n1 plus.n0 36.5157
R346 plus.n2 plus.n1 36.5157
R347 plus.n6 plus.n5 36.5157
R348 plus.n5 plus.n4 36.5157
R349 plus plus.n7 25.3835
R350 plus plus.n3 9.90391
R351 drain_left.n26 drain_left.n0 289.615
R352 drain_left.n59 drain_left.n33 289.615
R353 drain_left.n11 drain_left.n10 185
R354 drain_left.n8 drain_left.n7 185
R355 drain_left.n17 drain_left.n16 185
R356 drain_left.n19 drain_left.n18 185
R357 drain_left.n4 drain_left.n3 185
R358 drain_left.n25 drain_left.n24 185
R359 drain_left.n27 drain_left.n26 185
R360 drain_left.n60 drain_left.n59 185
R361 drain_left.n58 drain_left.n57 185
R362 drain_left.n37 drain_left.n36 185
R363 drain_left.n52 drain_left.n51 185
R364 drain_left.n50 drain_left.n49 185
R365 drain_left.n41 drain_left.n40 185
R366 drain_left.n44 drain_left.n43 185
R367 drain_left.t1 drain_left.n9 147.661
R368 drain_left.t4 drain_left.n42 147.661
R369 drain_left.n10 drain_left.n7 104.615
R370 drain_left.n17 drain_left.n7 104.615
R371 drain_left.n18 drain_left.n17 104.615
R372 drain_left.n18 drain_left.n3 104.615
R373 drain_left.n25 drain_left.n3 104.615
R374 drain_left.n26 drain_left.n25 104.615
R375 drain_left.n59 drain_left.n58 104.615
R376 drain_left.n58 drain_left.n36 104.615
R377 drain_left.n51 drain_left.n36 104.615
R378 drain_left.n51 drain_left.n50 104.615
R379 drain_left.n50 drain_left.n40 104.615
R380 drain_left.n43 drain_left.n40 104.615
R381 drain_left.n32 drain_left.n31 67.2711
R382 drain_left.n65 drain_left.n64 67.1907
R383 drain_left.n10 drain_left.t1 52.3082
R384 drain_left.n43 drain_left.t4 52.3082
R385 drain_left.n65 drain_left.n63 49.4072
R386 drain_left.n32 drain_left.n30 49.2161
R387 drain_left drain_left.n32 24.3152
R388 drain_left.n11 drain_left.n9 15.6674
R389 drain_left.n44 drain_left.n42 15.6674
R390 drain_left.n12 drain_left.n8 12.8005
R391 drain_left.n45 drain_left.n41 12.8005
R392 drain_left.n16 drain_left.n15 12.0247
R393 drain_left.n49 drain_left.n48 12.0247
R394 drain_left.n19 drain_left.n6 11.249
R395 drain_left.n52 drain_left.n39 11.249
R396 drain_left.n20 drain_left.n4 10.4732
R397 drain_left.n53 drain_left.n37 10.4732
R398 drain_left.n24 drain_left.n23 9.69747
R399 drain_left.n57 drain_left.n56 9.69747
R400 drain_left.n30 drain_left.n29 9.45567
R401 drain_left.n63 drain_left.n62 9.45567
R402 drain_left.n29 drain_left.n28 9.3005
R403 drain_left.n2 drain_left.n1 9.3005
R404 drain_left.n23 drain_left.n22 9.3005
R405 drain_left.n21 drain_left.n20 9.3005
R406 drain_left.n6 drain_left.n5 9.3005
R407 drain_left.n15 drain_left.n14 9.3005
R408 drain_left.n13 drain_left.n12 9.3005
R409 drain_left.n62 drain_left.n61 9.3005
R410 drain_left.n35 drain_left.n34 9.3005
R411 drain_left.n56 drain_left.n55 9.3005
R412 drain_left.n54 drain_left.n53 9.3005
R413 drain_left.n39 drain_left.n38 9.3005
R414 drain_left.n48 drain_left.n47 9.3005
R415 drain_left.n46 drain_left.n45 9.3005
R416 drain_left.n27 drain_left.n2 8.92171
R417 drain_left.n60 drain_left.n35 8.92171
R418 drain_left.n28 drain_left.n0 8.14595
R419 drain_left.n61 drain_left.n33 8.14595
R420 drain_left drain_left.n65 6.19632
R421 drain_left.n30 drain_left.n0 5.81868
R422 drain_left.n63 drain_left.n33 5.81868
R423 drain_left.n28 drain_left.n27 5.04292
R424 drain_left.n61 drain_left.n60 5.04292
R425 drain_left.n13 drain_left.n9 4.38594
R426 drain_left.n46 drain_left.n42 4.38594
R427 drain_left.n24 drain_left.n2 4.26717
R428 drain_left.n57 drain_left.n35 4.26717
R429 drain_left.n23 drain_left.n4 3.49141
R430 drain_left.n56 drain_left.n37 3.49141
R431 drain_left.n31 drain_left.t5 3.3005
R432 drain_left.n31 drain_left.t2 3.3005
R433 drain_left.n64 drain_left.t3 3.3005
R434 drain_left.n64 drain_left.t0 3.3005
R435 drain_left.n20 drain_left.n19 2.71565
R436 drain_left.n53 drain_left.n52 2.71565
R437 drain_left.n16 drain_left.n6 1.93989
R438 drain_left.n49 drain_left.n39 1.93989
R439 drain_left.n15 drain_left.n8 1.16414
R440 drain_left.n48 drain_left.n41 1.16414
R441 drain_left.n12 drain_left.n11 0.388379
R442 drain_left.n45 drain_left.n44 0.388379
R443 drain_left.n14 drain_left.n13 0.155672
R444 drain_left.n14 drain_left.n5 0.155672
R445 drain_left.n21 drain_left.n5 0.155672
R446 drain_left.n22 drain_left.n21 0.155672
R447 drain_left.n22 drain_left.n1 0.155672
R448 drain_left.n29 drain_left.n1 0.155672
R449 drain_left.n62 drain_left.n34 0.155672
R450 drain_left.n55 drain_left.n34 0.155672
R451 drain_left.n55 drain_left.n54 0.155672
R452 drain_left.n54 drain_left.n38 0.155672
R453 drain_left.n47 drain_left.n38 0.155672
R454 drain_left.n47 drain_left.n46 0.155672
C0 drain_left plus 1.63569f
C1 source minus 1.35466f
C2 drain_right plus 0.268691f
C3 drain_left minus 0.17071f
C4 drain_left source 7.86778f
C5 drain_right minus 1.52296f
C6 source drain_right 7.86099f
C7 drain_left drain_right 0.566534f
C8 minus plus 3.55718f
C9 source plus 1.369f
C10 drain_right a_n1220_n2088# 4.26199f
C11 drain_left a_n1220_n2088# 4.42282f
C12 source a_n1220_n2088# 3.819627f
C13 minus a_n1220_n2088# 4.186829f
C14 plus a_n1220_n2088# 5.001717f
C15 drain_left.n0 a_n1220_n2088# 0.031709f
C16 drain_left.n1 a_n1220_n2088# 0.022559f
C17 drain_left.n2 a_n1220_n2088# 0.012122f
C18 drain_left.n3 a_n1220_n2088# 0.028653f
C19 drain_left.n4 a_n1220_n2088# 0.012835f
C20 drain_left.n5 a_n1220_n2088# 0.022559f
C21 drain_left.n6 a_n1220_n2088# 0.012122f
C22 drain_left.n7 a_n1220_n2088# 0.028653f
C23 drain_left.n8 a_n1220_n2088# 0.012835f
C24 drain_left.n9 a_n1220_n2088# 0.096538f
C25 drain_left.t1 a_n1220_n2088# 0.0467f
C26 drain_left.n10 a_n1220_n2088# 0.02149f
C27 drain_left.n11 a_n1220_n2088# 0.016925f
C28 drain_left.n12 a_n1220_n2088# 0.012122f
C29 drain_left.n13 a_n1220_n2088# 0.536775f
C30 drain_left.n14 a_n1220_n2088# 0.022559f
C31 drain_left.n15 a_n1220_n2088# 0.012122f
C32 drain_left.n16 a_n1220_n2088# 0.012835f
C33 drain_left.n17 a_n1220_n2088# 0.028653f
C34 drain_left.n18 a_n1220_n2088# 0.028653f
C35 drain_left.n19 a_n1220_n2088# 0.012835f
C36 drain_left.n20 a_n1220_n2088# 0.012122f
C37 drain_left.n21 a_n1220_n2088# 0.022559f
C38 drain_left.n22 a_n1220_n2088# 0.022559f
C39 drain_left.n23 a_n1220_n2088# 0.012122f
C40 drain_left.n24 a_n1220_n2088# 0.012835f
C41 drain_left.n25 a_n1220_n2088# 0.028653f
C42 drain_left.n26 a_n1220_n2088# 0.062029f
C43 drain_left.n27 a_n1220_n2088# 0.012835f
C44 drain_left.n28 a_n1220_n2088# 0.012122f
C45 drain_left.n29 a_n1220_n2088# 0.052145f
C46 drain_left.n30 a_n1220_n2088# 0.050788f
C47 drain_left.t5 a_n1220_n2088# 0.106962f
C48 drain_left.t2 a_n1220_n2088# 0.106962f
C49 drain_left.n31 a_n1220_n2088# 0.892355f
C50 drain_left.n32 a_n1220_n2088# 0.977717f
C51 drain_left.n33 a_n1220_n2088# 0.031709f
C52 drain_left.n34 a_n1220_n2088# 0.022559f
C53 drain_left.n35 a_n1220_n2088# 0.012122f
C54 drain_left.n36 a_n1220_n2088# 0.028653f
C55 drain_left.n37 a_n1220_n2088# 0.012835f
C56 drain_left.n38 a_n1220_n2088# 0.022559f
C57 drain_left.n39 a_n1220_n2088# 0.012122f
C58 drain_left.n40 a_n1220_n2088# 0.028653f
C59 drain_left.n41 a_n1220_n2088# 0.012835f
C60 drain_left.n42 a_n1220_n2088# 0.096538f
C61 drain_left.t4 a_n1220_n2088# 0.0467f
C62 drain_left.n43 a_n1220_n2088# 0.02149f
C63 drain_left.n44 a_n1220_n2088# 0.016925f
C64 drain_left.n45 a_n1220_n2088# 0.012122f
C65 drain_left.n46 a_n1220_n2088# 0.536775f
C66 drain_left.n47 a_n1220_n2088# 0.022559f
C67 drain_left.n48 a_n1220_n2088# 0.012122f
C68 drain_left.n49 a_n1220_n2088# 0.012835f
C69 drain_left.n50 a_n1220_n2088# 0.028653f
C70 drain_left.n51 a_n1220_n2088# 0.028653f
C71 drain_left.n52 a_n1220_n2088# 0.012835f
C72 drain_left.n53 a_n1220_n2088# 0.012122f
C73 drain_left.n54 a_n1220_n2088# 0.022559f
C74 drain_left.n55 a_n1220_n2088# 0.022559f
C75 drain_left.n56 a_n1220_n2088# 0.012122f
C76 drain_left.n57 a_n1220_n2088# 0.012835f
C77 drain_left.n58 a_n1220_n2088# 0.028653f
C78 drain_left.n59 a_n1220_n2088# 0.062029f
C79 drain_left.n60 a_n1220_n2088# 0.012835f
C80 drain_left.n61 a_n1220_n2088# 0.012122f
C81 drain_left.n62 a_n1220_n2088# 0.052145f
C82 drain_left.n63 a_n1220_n2088# 0.051195f
C83 drain_left.t3 a_n1220_n2088# 0.106962f
C84 drain_left.t0 a_n1220_n2088# 0.106962f
C85 drain_left.n64 a_n1220_n2088# 0.892063f
C86 drain_left.n65 a_n1220_n2088# 0.531837f
C87 plus.t1 a_n1220_n2088# 0.173939f
C88 plus.n0 a_n1220_n2088# 0.086792f
C89 plus.t2 a_n1220_n2088# 0.166998f
C90 plus.n1 a_n1220_n2088# 0.076655f
C91 plus.t5 a_n1220_n2088# 0.173939f
C92 plus.n2 a_n1220_n2088# 0.086741f
C93 plus.n3 a_n1220_n2088# 0.325396f
C94 plus.t3 a_n1220_n2088# 0.173939f
C95 plus.n4 a_n1220_n2088# 0.086792f
C96 plus.t4 a_n1220_n2088# 0.173939f
C97 plus.t0 a_n1220_n2088# 0.166998f
C98 plus.n5 a_n1220_n2088# 0.076655f
C99 plus.n6 a_n1220_n2088# 0.086741f
C100 plus.n7 a_n1220_n2088# 0.777961f
C101 drain_right.n0 a_n1220_n2088# 0.032067f
C102 drain_right.n1 a_n1220_n2088# 0.022814f
C103 drain_right.n2 a_n1220_n2088# 0.012259f
C104 drain_right.n3 a_n1220_n2088# 0.028977f
C105 drain_right.n4 a_n1220_n2088# 0.01298f
C106 drain_right.n5 a_n1220_n2088# 0.022814f
C107 drain_right.n6 a_n1220_n2088# 0.012259f
C108 drain_right.n7 a_n1220_n2088# 0.028977f
C109 drain_right.n8 a_n1220_n2088# 0.01298f
C110 drain_right.n9 a_n1220_n2088# 0.097628f
C111 drain_right.t1 a_n1220_n2088# 0.047228f
C112 drain_right.n10 a_n1220_n2088# 0.021732f
C113 drain_right.n11 a_n1220_n2088# 0.017116f
C114 drain_right.n12 a_n1220_n2088# 0.012259f
C115 drain_right.n13 a_n1220_n2088# 0.542839f
C116 drain_right.n14 a_n1220_n2088# 0.022814f
C117 drain_right.n15 a_n1220_n2088# 0.012259f
C118 drain_right.n16 a_n1220_n2088# 0.01298f
C119 drain_right.n17 a_n1220_n2088# 0.028977f
C120 drain_right.n18 a_n1220_n2088# 0.028977f
C121 drain_right.n19 a_n1220_n2088# 0.01298f
C122 drain_right.n20 a_n1220_n2088# 0.012259f
C123 drain_right.n21 a_n1220_n2088# 0.022814f
C124 drain_right.n22 a_n1220_n2088# 0.022814f
C125 drain_right.n23 a_n1220_n2088# 0.012259f
C126 drain_right.n24 a_n1220_n2088# 0.01298f
C127 drain_right.n25 a_n1220_n2088# 0.028977f
C128 drain_right.n26 a_n1220_n2088# 0.062729f
C129 drain_right.n27 a_n1220_n2088# 0.01298f
C130 drain_right.n28 a_n1220_n2088# 0.012259f
C131 drain_right.n29 a_n1220_n2088# 0.052734f
C132 drain_right.n30 a_n1220_n2088# 0.051362f
C133 drain_right.t4 a_n1220_n2088# 0.10817f
C134 drain_right.t2 a_n1220_n2088# 0.10817f
C135 drain_right.n31 a_n1220_n2088# 0.902435f
C136 drain_right.n32 a_n1220_n2088# 0.941939f
C137 drain_right.t0 a_n1220_n2088# 0.10817f
C138 drain_right.t3 a_n1220_n2088# 0.10817f
C139 drain_right.n33 a_n1220_n2088# 0.904339f
C140 drain_right.n34 a_n1220_n2088# 0.032067f
C141 drain_right.n35 a_n1220_n2088# 0.022814f
C142 drain_right.n36 a_n1220_n2088# 0.012259f
C143 drain_right.n37 a_n1220_n2088# 0.028977f
C144 drain_right.n38 a_n1220_n2088# 0.01298f
C145 drain_right.n39 a_n1220_n2088# 0.022814f
C146 drain_right.n40 a_n1220_n2088# 0.012259f
C147 drain_right.n41 a_n1220_n2088# 0.028977f
C148 drain_right.n42 a_n1220_n2088# 0.01298f
C149 drain_right.n43 a_n1220_n2088# 0.097628f
C150 drain_right.t5 a_n1220_n2088# 0.047228f
C151 drain_right.n44 a_n1220_n2088# 0.021732f
C152 drain_right.n45 a_n1220_n2088# 0.017116f
C153 drain_right.n46 a_n1220_n2088# 0.012259f
C154 drain_right.n47 a_n1220_n2088# 0.542839f
C155 drain_right.n48 a_n1220_n2088# 0.022814f
C156 drain_right.n49 a_n1220_n2088# 0.012259f
C157 drain_right.n50 a_n1220_n2088# 0.01298f
C158 drain_right.n51 a_n1220_n2088# 0.028977f
C159 drain_right.n52 a_n1220_n2088# 0.028977f
C160 drain_right.n53 a_n1220_n2088# 0.01298f
C161 drain_right.n54 a_n1220_n2088# 0.012259f
C162 drain_right.n55 a_n1220_n2088# 0.022814f
C163 drain_right.n56 a_n1220_n2088# 0.022814f
C164 drain_right.n57 a_n1220_n2088# 0.012259f
C165 drain_right.n58 a_n1220_n2088# 0.01298f
C166 drain_right.n59 a_n1220_n2088# 0.028977f
C167 drain_right.n60 a_n1220_n2088# 0.062729f
C168 drain_right.n61 a_n1220_n2088# 0.01298f
C169 drain_right.n62 a_n1220_n2088# 0.012259f
C170 drain_right.n63 a_n1220_n2088# 0.052734f
C171 drain_right.n64 a_n1220_n2088# 0.050852f
C172 drain_right.n65 a_n1220_n2088# 0.546187f
C173 source.n0 a_n1220_n2088# 0.035393f
C174 source.n1 a_n1220_n2088# 0.02518f
C175 source.n2 a_n1220_n2088# 0.013531f
C176 source.n3 a_n1220_n2088# 0.031982f
C177 source.n4 a_n1220_n2088# 0.014327f
C178 source.n5 a_n1220_n2088# 0.02518f
C179 source.n6 a_n1220_n2088# 0.013531f
C180 source.n7 a_n1220_n2088# 0.031982f
C181 source.n8 a_n1220_n2088# 0.014327f
C182 source.n9 a_n1220_n2088# 0.107754f
C183 source.t5 a_n1220_n2088# 0.052126f
C184 source.n10 a_n1220_n2088# 0.023986f
C185 source.n11 a_n1220_n2088# 0.018891f
C186 source.n12 a_n1220_n2088# 0.013531f
C187 source.n13 a_n1220_n2088# 0.59914f
C188 source.n14 a_n1220_n2088# 0.02518f
C189 source.n15 a_n1220_n2088# 0.013531f
C190 source.n16 a_n1220_n2088# 0.014327f
C191 source.n17 a_n1220_n2088# 0.031982f
C192 source.n18 a_n1220_n2088# 0.031982f
C193 source.n19 a_n1220_n2088# 0.014327f
C194 source.n20 a_n1220_n2088# 0.013531f
C195 source.n21 a_n1220_n2088# 0.02518f
C196 source.n22 a_n1220_n2088# 0.02518f
C197 source.n23 a_n1220_n2088# 0.013531f
C198 source.n24 a_n1220_n2088# 0.014327f
C199 source.n25 a_n1220_n2088# 0.031982f
C200 source.n26 a_n1220_n2088# 0.069235f
C201 source.n27 a_n1220_n2088# 0.014327f
C202 source.n28 a_n1220_n2088# 0.013531f
C203 source.n29 a_n1220_n2088# 0.058203f
C204 source.n30 a_n1220_n2088# 0.03874f
C205 source.n31 a_n1220_n2088# 0.609916f
C206 source.t4 a_n1220_n2088# 0.119389f
C207 source.t3 a_n1220_n2088# 0.119389f
C208 source.n32 a_n1220_n2088# 0.929813f
C209 source.n33 a_n1220_n2088# 0.340259f
C210 source.n34 a_n1220_n2088# 0.035393f
C211 source.n35 a_n1220_n2088# 0.02518f
C212 source.n36 a_n1220_n2088# 0.013531f
C213 source.n37 a_n1220_n2088# 0.031982f
C214 source.n38 a_n1220_n2088# 0.014327f
C215 source.n39 a_n1220_n2088# 0.02518f
C216 source.n40 a_n1220_n2088# 0.013531f
C217 source.n41 a_n1220_n2088# 0.031982f
C218 source.n42 a_n1220_n2088# 0.014327f
C219 source.n43 a_n1220_n2088# 0.107754f
C220 source.t10 a_n1220_n2088# 0.052126f
C221 source.n44 a_n1220_n2088# 0.023986f
C222 source.n45 a_n1220_n2088# 0.018891f
C223 source.n46 a_n1220_n2088# 0.013531f
C224 source.n47 a_n1220_n2088# 0.59914f
C225 source.n48 a_n1220_n2088# 0.02518f
C226 source.n49 a_n1220_n2088# 0.013531f
C227 source.n50 a_n1220_n2088# 0.014327f
C228 source.n51 a_n1220_n2088# 0.031982f
C229 source.n52 a_n1220_n2088# 0.031982f
C230 source.n53 a_n1220_n2088# 0.014327f
C231 source.n54 a_n1220_n2088# 0.013531f
C232 source.n55 a_n1220_n2088# 0.02518f
C233 source.n56 a_n1220_n2088# 0.02518f
C234 source.n57 a_n1220_n2088# 0.013531f
C235 source.n58 a_n1220_n2088# 0.014327f
C236 source.n59 a_n1220_n2088# 0.031982f
C237 source.n60 a_n1220_n2088# 0.069235f
C238 source.n61 a_n1220_n2088# 0.014327f
C239 source.n62 a_n1220_n2088# 0.013531f
C240 source.n63 a_n1220_n2088# 0.058203f
C241 source.n64 a_n1220_n2088# 0.03874f
C242 source.n65 a_n1220_n2088# 0.125724f
C243 source.t11 a_n1220_n2088# 0.119389f
C244 source.t7 a_n1220_n2088# 0.119389f
C245 source.n66 a_n1220_n2088# 0.929813f
C246 source.n67 a_n1220_n2088# 1.19269f
C247 source.t1 a_n1220_n2088# 0.119389f
C248 source.t0 a_n1220_n2088# 0.119389f
C249 source.n68 a_n1220_n2088# 0.929807f
C250 source.n69 a_n1220_n2088# 1.19269f
C251 source.n70 a_n1220_n2088# 0.035393f
C252 source.n71 a_n1220_n2088# 0.02518f
C253 source.n72 a_n1220_n2088# 0.013531f
C254 source.n73 a_n1220_n2088# 0.031982f
C255 source.n74 a_n1220_n2088# 0.014327f
C256 source.n75 a_n1220_n2088# 0.02518f
C257 source.n76 a_n1220_n2088# 0.013531f
C258 source.n77 a_n1220_n2088# 0.031982f
C259 source.n78 a_n1220_n2088# 0.014327f
C260 source.n79 a_n1220_n2088# 0.107754f
C261 source.t2 a_n1220_n2088# 0.052126f
C262 source.n80 a_n1220_n2088# 0.023986f
C263 source.n81 a_n1220_n2088# 0.018891f
C264 source.n82 a_n1220_n2088# 0.013531f
C265 source.n83 a_n1220_n2088# 0.59914f
C266 source.n84 a_n1220_n2088# 0.02518f
C267 source.n85 a_n1220_n2088# 0.013531f
C268 source.n86 a_n1220_n2088# 0.014327f
C269 source.n87 a_n1220_n2088# 0.031982f
C270 source.n88 a_n1220_n2088# 0.031982f
C271 source.n89 a_n1220_n2088# 0.014327f
C272 source.n90 a_n1220_n2088# 0.013531f
C273 source.n91 a_n1220_n2088# 0.02518f
C274 source.n92 a_n1220_n2088# 0.02518f
C275 source.n93 a_n1220_n2088# 0.013531f
C276 source.n94 a_n1220_n2088# 0.014327f
C277 source.n95 a_n1220_n2088# 0.031982f
C278 source.n96 a_n1220_n2088# 0.069235f
C279 source.n97 a_n1220_n2088# 0.014327f
C280 source.n98 a_n1220_n2088# 0.013531f
C281 source.n99 a_n1220_n2088# 0.058203f
C282 source.n100 a_n1220_n2088# 0.03874f
C283 source.n101 a_n1220_n2088# 0.125724f
C284 source.t6 a_n1220_n2088# 0.119389f
C285 source.t8 a_n1220_n2088# 0.119389f
C286 source.n102 a_n1220_n2088# 0.929807f
C287 source.n103 a_n1220_n2088# 0.340266f
C288 source.n104 a_n1220_n2088# 0.035393f
C289 source.n105 a_n1220_n2088# 0.02518f
C290 source.n106 a_n1220_n2088# 0.013531f
C291 source.n107 a_n1220_n2088# 0.031982f
C292 source.n108 a_n1220_n2088# 0.014327f
C293 source.n109 a_n1220_n2088# 0.02518f
C294 source.n110 a_n1220_n2088# 0.013531f
C295 source.n111 a_n1220_n2088# 0.031982f
C296 source.n112 a_n1220_n2088# 0.014327f
C297 source.n113 a_n1220_n2088# 0.107754f
C298 source.t9 a_n1220_n2088# 0.052126f
C299 source.n114 a_n1220_n2088# 0.023986f
C300 source.n115 a_n1220_n2088# 0.018891f
C301 source.n116 a_n1220_n2088# 0.013531f
C302 source.n117 a_n1220_n2088# 0.59914f
C303 source.n118 a_n1220_n2088# 0.02518f
C304 source.n119 a_n1220_n2088# 0.013531f
C305 source.n120 a_n1220_n2088# 0.014327f
C306 source.n121 a_n1220_n2088# 0.031982f
C307 source.n122 a_n1220_n2088# 0.031982f
C308 source.n123 a_n1220_n2088# 0.014327f
C309 source.n124 a_n1220_n2088# 0.013531f
C310 source.n125 a_n1220_n2088# 0.02518f
C311 source.n126 a_n1220_n2088# 0.02518f
C312 source.n127 a_n1220_n2088# 0.013531f
C313 source.n128 a_n1220_n2088# 0.014327f
C314 source.n129 a_n1220_n2088# 0.031982f
C315 source.n130 a_n1220_n2088# 0.069235f
C316 source.n131 a_n1220_n2088# 0.014327f
C317 source.n132 a_n1220_n2088# 0.013531f
C318 source.n133 a_n1220_n2088# 0.058203f
C319 source.n134 a_n1220_n2088# 0.03874f
C320 source.n135 a_n1220_n2088# 0.245834f
C321 source.n136 a_n1220_n2088# 1.03033f
C322 minus.t2 a_n1220_n2088# 0.170814f
C323 minus.n0 a_n1220_n2088# 0.085233f
C324 minus.t0 a_n1220_n2088# 0.170814f
C325 minus.t5 a_n1220_n2088# 0.163999f
C326 minus.n1 a_n1220_n2088# 0.075278f
C327 minus.n2 a_n1220_n2088# 0.085183f
C328 minus.n3 a_n1220_n2088# 0.839465f
C329 minus.t4 a_n1220_n2088# 0.170814f
C330 minus.n4 a_n1220_n2088# 0.085233f
C331 minus.t1 a_n1220_n2088# 0.163999f
C332 minus.n5 a_n1220_n2088# 0.075278f
C333 minus.t3 a_n1220_n2088# 0.170814f
C334 minus.n6 a_n1220_n2088# 0.085183f
C335 minus.n7 a_n1220_n2088# 0.25449f
C336 minus.n8 a_n1220_n2088# 0.982405f
.ends

