* NGSPICE file created from diffpair570.ext - technology: sky130A

.subckt diffpair570 minus drain_right drain_left source plus
X0 drain_right minus source a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.2
X1 a_n928_n4892# a_n928_n4892# a_n928_n4892# a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X2 a_n928_n4892# a_n928_n4892# a_n928_n4892# a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X3 drain_left plus source a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.2
X4 a_n928_n4892# a_n928_n4892# a_n928_n4892# a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X5 a_n928_n4892# a_n928_n4892# a_n928_n4892# a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X6 drain_right minus source a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.2
X7 drain_left plus source a_n928_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.2
.ends

