* NGSPICE file created from diffpair271.ext - technology: sky130A

.subckt diffpair271 minus drain_right drain_left source plus
X0 drain_right minus source a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X1 a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X2 source minus drain_right a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X3 a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X4 source minus drain_right a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X5 a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X6 source plus drain_left a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X7 a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X8 source plus drain_left a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X9 drain_right minus source a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X10 drain_left plus source a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X11 drain_left plus source a_n1094_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
.ends

