* NGSPICE file created from diffpair414.ext - technology: sky130A

.subckt diffpair414 minus drain_right drain_left source plus
X0 a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X1 drain_right.t9 minus.t0 source.t15 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X2 drain_right.t8 minus.t1 source.t17 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X3 drain_right.t7 minus.t2 source.t13 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X4 source.t6 plus.t0 drain_left.t9 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X5 source.t14 minus.t3 drain_right.t6 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X6 source.t16 minus.t4 drain_right.t5 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X7 source.t9 minus.t5 drain_right.t4 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X8 drain_left.t8 plus.t1 source.t4 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X9 drain_right.t3 minus.t6 source.t11 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X10 a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X11 a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X12 drain_right.t2 minus.t7 source.t10 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X13 drain_right.t1 minus.t8 source.t18 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X14 source.t19 plus.t2 drain_left.t7 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X15 drain_left.t6 plus.t3 source.t1 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X16 source.t5 plus.t4 drain_left.t5 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X17 drain_left.t4 plus.t5 source.t8 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X18 drain_left.t3 plus.t6 source.t7 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X19 source.t12 minus.t9 drain_right.t0 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X20 drain_left.t2 plus.t7 source.t0 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X21 a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X22 drain_left.t1 plus.t8 source.t3 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X23 source.t2 plus.t9 drain_left.t0 a_n1352_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 minus.n8 minus.t8 1647.93
R1 minus.n2 minus.t7 1647.93
R2 minus.n18 minus.t6 1647.93
R3 minus.n12 minus.t2 1647.93
R4 minus.n7 minus.t9 1602.65
R5 minus.n5 minus.t0 1602.65
R6 minus.n1 minus.t5 1602.65
R7 minus.n17 minus.t3 1602.65
R8 minus.n15 minus.t1 1602.65
R9 minus.n11 minus.t4 1602.65
R10 minus.n3 minus.n2 161.489
R11 minus.n13 minus.n12 161.489
R12 minus.n9 minus.n8 161.3
R13 minus.n6 minus.n0 161.3
R14 minus.n4 minus.n3 161.3
R15 minus.n19 minus.n18 161.3
R16 minus.n16 minus.n10 161.3
R17 minus.n14 minus.n13 161.3
R18 minus.n7 minus.n6 40.8975
R19 minus.n4 minus.n1 40.8975
R20 minus.n14 minus.n11 40.8975
R21 minus.n17 minus.n16 40.8975
R22 minus.n6 minus.n5 36.5157
R23 minus.n5 minus.n4 36.5157
R24 minus.n15 minus.n14 36.5157
R25 minus.n16 minus.n15 36.5157
R26 minus.n20 minus.n9 34.1918
R27 minus.n8 minus.n7 32.1338
R28 minus.n2 minus.n1 32.1338
R29 minus.n12 minus.n11 32.1338
R30 minus.n18 minus.n17 32.1338
R31 minus.n20 minus.n19 6.44936
R32 minus.n9 minus.n0 0.189894
R33 minus.n3 minus.n0 0.189894
R34 minus.n13 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n274 source.n214 289.615
R38 source.n204 source.n144 289.615
R39 source.n60 source.n0 289.615
R40 source.n130 source.n70 289.615
R41 source.n234 source.n233 185
R42 source.n239 source.n238 185
R43 source.n241 source.n240 185
R44 source.n230 source.n229 185
R45 source.n247 source.n246 185
R46 source.n249 source.n248 185
R47 source.n226 source.n225 185
R48 source.n256 source.n255 185
R49 source.n257 source.n224 185
R50 source.n259 source.n258 185
R51 source.n222 source.n221 185
R52 source.n265 source.n264 185
R53 source.n267 source.n266 185
R54 source.n218 source.n217 185
R55 source.n273 source.n272 185
R56 source.n275 source.n274 185
R57 source.n164 source.n163 185
R58 source.n169 source.n168 185
R59 source.n171 source.n170 185
R60 source.n160 source.n159 185
R61 source.n177 source.n176 185
R62 source.n179 source.n178 185
R63 source.n156 source.n155 185
R64 source.n186 source.n185 185
R65 source.n187 source.n154 185
R66 source.n189 source.n188 185
R67 source.n152 source.n151 185
R68 source.n195 source.n194 185
R69 source.n197 source.n196 185
R70 source.n148 source.n147 185
R71 source.n203 source.n202 185
R72 source.n205 source.n204 185
R73 source.n61 source.n60 185
R74 source.n59 source.n58 185
R75 source.n4 source.n3 185
R76 source.n53 source.n52 185
R77 source.n51 source.n50 185
R78 source.n8 source.n7 185
R79 source.n45 source.n44 185
R80 source.n43 source.n10 185
R81 source.n42 source.n41 185
R82 source.n13 source.n11 185
R83 source.n36 source.n35 185
R84 source.n34 source.n33 185
R85 source.n17 source.n16 185
R86 source.n28 source.n27 185
R87 source.n26 source.n25 185
R88 source.n21 source.n20 185
R89 source.n131 source.n130 185
R90 source.n129 source.n128 185
R91 source.n74 source.n73 185
R92 source.n123 source.n122 185
R93 source.n121 source.n120 185
R94 source.n78 source.n77 185
R95 source.n115 source.n114 185
R96 source.n113 source.n80 185
R97 source.n112 source.n111 185
R98 source.n83 source.n81 185
R99 source.n106 source.n105 185
R100 source.n104 source.n103 185
R101 source.n87 source.n86 185
R102 source.n98 source.n97 185
R103 source.n96 source.n95 185
R104 source.n91 source.n90 185
R105 source.n235 source.t11 149.524
R106 source.n165 source.t0 149.524
R107 source.n22 source.t1 149.524
R108 source.n92 source.t10 149.524
R109 source.n239 source.n233 104.615
R110 source.n240 source.n239 104.615
R111 source.n240 source.n229 104.615
R112 source.n247 source.n229 104.615
R113 source.n248 source.n247 104.615
R114 source.n248 source.n225 104.615
R115 source.n256 source.n225 104.615
R116 source.n257 source.n256 104.615
R117 source.n258 source.n257 104.615
R118 source.n258 source.n221 104.615
R119 source.n265 source.n221 104.615
R120 source.n266 source.n265 104.615
R121 source.n266 source.n217 104.615
R122 source.n273 source.n217 104.615
R123 source.n274 source.n273 104.615
R124 source.n169 source.n163 104.615
R125 source.n170 source.n169 104.615
R126 source.n170 source.n159 104.615
R127 source.n177 source.n159 104.615
R128 source.n178 source.n177 104.615
R129 source.n178 source.n155 104.615
R130 source.n186 source.n155 104.615
R131 source.n187 source.n186 104.615
R132 source.n188 source.n187 104.615
R133 source.n188 source.n151 104.615
R134 source.n195 source.n151 104.615
R135 source.n196 source.n195 104.615
R136 source.n196 source.n147 104.615
R137 source.n203 source.n147 104.615
R138 source.n204 source.n203 104.615
R139 source.n60 source.n59 104.615
R140 source.n59 source.n3 104.615
R141 source.n52 source.n3 104.615
R142 source.n52 source.n51 104.615
R143 source.n51 source.n7 104.615
R144 source.n44 source.n7 104.615
R145 source.n44 source.n43 104.615
R146 source.n43 source.n42 104.615
R147 source.n42 source.n11 104.615
R148 source.n35 source.n11 104.615
R149 source.n35 source.n34 104.615
R150 source.n34 source.n16 104.615
R151 source.n27 source.n16 104.615
R152 source.n27 source.n26 104.615
R153 source.n26 source.n20 104.615
R154 source.n130 source.n129 104.615
R155 source.n129 source.n73 104.615
R156 source.n122 source.n73 104.615
R157 source.n122 source.n121 104.615
R158 source.n121 source.n77 104.615
R159 source.n114 source.n77 104.615
R160 source.n114 source.n113 104.615
R161 source.n113 source.n112 104.615
R162 source.n112 source.n81 104.615
R163 source.n105 source.n81 104.615
R164 source.n105 source.n104 104.615
R165 source.n104 source.n86 104.615
R166 source.n97 source.n86 104.615
R167 source.n97 source.n96 104.615
R168 source.n96 source.n90 104.615
R169 source.t11 source.n233 52.3082
R170 source.t0 source.n163 52.3082
R171 source.t1 source.n20 52.3082
R172 source.t10 source.n90 52.3082
R173 source.n67 source.n66 42.8739
R174 source.n69 source.n68 42.8739
R175 source.n137 source.n136 42.8739
R176 source.n139 source.n138 42.8739
R177 source.n213 source.n212 42.8737
R178 source.n211 source.n210 42.8737
R179 source.n143 source.n142 42.8737
R180 source.n141 source.n140 42.8737
R181 source.n279 source.n278 29.8581
R182 source.n209 source.n208 29.8581
R183 source.n65 source.n64 29.8581
R184 source.n135 source.n134 29.8581
R185 source.n141 source.n139 22.2015
R186 source.n280 source.n65 16.2532
R187 source.n259 source.n224 13.1884
R188 source.n189 source.n154 13.1884
R189 source.n45 source.n10 13.1884
R190 source.n115 source.n80 13.1884
R191 source.n255 source.n254 12.8005
R192 source.n260 source.n222 12.8005
R193 source.n185 source.n184 12.8005
R194 source.n190 source.n152 12.8005
R195 source.n46 source.n8 12.8005
R196 source.n41 source.n12 12.8005
R197 source.n116 source.n78 12.8005
R198 source.n111 source.n82 12.8005
R199 source.n253 source.n226 12.0247
R200 source.n264 source.n263 12.0247
R201 source.n183 source.n156 12.0247
R202 source.n194 source.n193 12.0247
R203 source.n50 source.n49 12.0247
R204 source.n40 source.n13 12.0247
R205 source.n120 source.n119 12.0247
R206 source.n110 source.n83 12.0247
R207 source.n250 source.n249 11.249
R208 source.n267 source.n220 11.249
R209 source.n180 source.n179 11.249
R210 source.n197 source.n150 11.249
R211 source.n53 source.n6 11.249
R212 source.n37 source.n36 11.249
R213 source.n123 source.n76 11.249
R214 source.n107 source.n106 11.249
R215 source.n246 source.n228 10.4732
R216 source.n268 source.n218 10.4732
R217 source.n176 source.n158 10.4732
R218 source.n198 source.n148 10.4732
R219 source.n54 source.n4 10.4732
R220 source.n33 source.n15 10.4732
R221 source.n124 source.n74 10.4732
R222 source.n103 source.n85 10.4732
R223 source.n235 source.n234 10.2747
R224 source.n165 source.n164 10.2747
R225 source.n22 source.n21 10.2747
R226 source.n92 source.n91 10.2747
R227 source.n245 source.n230 9.69747
R228 source.n272 source.n271 9.69747
R229 source.n175 source.n160 9.69747
R230 source.n202 source.n201 9.69747
R231 source.n58 source.n57 9.69747
R232 source.n32 source.n17 9.69747
R233 source.n128 source.n127 9.69747
R234 source.n102 source.n87 9.69747
R235 source.n278 source.n277 9.45567
R236 source.n208 source.n207 9.45567
R237 source.n64 source.n63 9.45567
R238 source.n134 source.n133 9.45567
R239 source.n277 source.n276 9.3005
R240 source.n216 source.n215 9.3005
R241 source.n271 source.n270 9.3005
R242 source.n269 source.n268 9.3005
R243 source.n220 source.n219 9.3005
R244 source.n263 source.n262 9.3005
R245 source.n261 source.n260 9.3005
R246 source.n237 source.n236 9.3005
R247 source.n232 source.n231 9.3005
R248 source.n243 source.n242 9.3005
R249 source.n245 source.n244 9.3005
R250 source.n228 source.n227 9.3005
R251 source.n251 source.n250 9.3005
R252 source.n253 source.n252 9.3005
R253 source.n254 source.n223 9.3005
R254 source.n207 source.n206 9.3005
R255 source.n146 source.n145 9.3005
R256 source.n201 source.n200 9.3005
R257 source.n199 source.n198 9.3005
R258 source.n150 source.n149 9.3005
R259 source.n193 source.n192 9.3005
R260 source.n191 source.n190 9.3005
R261 source.n167 source.n166 9.3005
R262 source.n162 source.n161 9.3005
R263 source.n173 source.n172 9.3005
R264 source.n175 source.n174 9.3005
R265 source.n158 source.n157 9.3005
R266 source.n181 source.n180 9.3005
R267 source.n183 source.n182 9.3005
R268 source.n184 source.n153 9.3005
R269 source.n24 source.n23 9.3005
R270 source.n19 source.n18 9.3005
R271 source.n30 source.n29 9.3005
R272 source.n32 source.n31 9.3005
R273 source.n15 source.n14 9.3005
R274 source.n38 source.n37 9.3005
R275 source.n40 source.n39 9.3005
R276 source.n12 source.n9 9.3005
R277 source.n63 source.n62 9.3005
R278 source.n2 source.n1 9.3005
R279 source.n57 source.n56 9.3005
R280 source.n55 source.n54 9.3005
R281 source.n6 source.n5 9.3005
R282 source.n49 source.n48 9.3005
R283 source.n47 source.n46 9.3005
R284 source.n94 source.n93 9.3005
R285 source.n89 source.n88 9.3005
R286 source.n100 source.n99 9.3005
R287 source.n102 source.n101 9.3005
R288 source.n85 source.n84 9.3005
R289 source.n108 source.n107 9.3005
R290 source.n110 source.n109 9.3005
R291 source.n82 source.n79 9.3005
R292 source.n133 source.n132 9.3005
R293 source.n72 source.n71 9.3005
R294 source.n127 source.n126 9.3005
R295 source.n125 source.n124 9.3005
R296 source.n76 source.n75 9.3005
R297 source.n119 source.n118 9.3005
R298 source.n117 source.n116 9.3005
R299 source.n242 source.n241 8.92171
R300 source.n275 source.n216 8.92171
R301 source.n172 source.n171 8.92171
R302 source.n205 source.n146 8.92171
R303 source.n61 source.n2 8.92171
R304 source.n29 source.n28 8.92171
R305 source.n131 source.n72 8.92171
R306 source.n99 source.n98 8.92171
R307 source.n238 source.n232 8.14595
R308 source.n276 source.n214 8.14595
R309 source.n168 source.n162 8.14595
R310 source.n206 source.n144 8.14595
R311 source.n62 source.n0 8.14595
R312 source.n25 source.n19 8.14595
R313 source.n132 source.n70 8.14595
R314 source.n95 source.n89 8.14595
R315 source.n237 source.n234 7.3702
R316 source.n167 source.n164 7.3702
R317 source.n24 source.n21 7.3702
R318 source.n94 source.n91 7.3702
R319 source.n238 source.n237 5.81868
R320 source.n278 source.n214 5.81868
R321 source.n168 source.n167 5.81868
R322 source.n208 source.n144 5.81868
R323 source.n64 source.n0 5.81868
R324 source.n25 source.n24 5.81868
R325 source.n134 source.n70 5.81868
R326 source.n95 source.n94 5.81868
R327 source.n280 source.n279 5.49188
R328 source.n241 source.n232 5.04292
R329 source.n276 source.n275 5.04292
R330 source.n171 source.n162 5.04292
R331 source.n206 source.n205 5.04292
R332 source.n62 source.n61 5.04292
R333 source.n28 source.n19 5.04292
R334 source.n132 source.n131 5.04292
R335 source.n98 source.n89 5.04292
R336 source.n242 source.n230 4.26717
R337 source.n272 source.n216 4.26717
R338 source.n172 source.n160 4.26717
R339 source.n202 source.n146 4.26717
R340 source.n58 source.n2 4.26717
R341 source.n29 source.n17 4.26717
R342 source.n128 source.n72 4.26717
R343 source.n99 source.n87 4.26717
R344 source.n246 source.n245 3.49141
R345 source.n271 source.n218 3.49141
R346 source.n176 source.n175 3.49141
R347 source.n201 source.n148 3.49141
R348 source.n57 source.n4 3.49141
R349 source.n33 source.n32 3.49141
R350 source.n127 source.n74 3.49141
R351 source.n103 source.n102 3.49141
R352 source.n236 source.n235 2.84303
R353 source.n166 source.n165 2.84303
R354 source.n23 source.n22 2.84303
R355 source.n93 source.n92 2.84303
R356 source.n249 source.n228 2.71565
R357 source.n268 source.n267 2.71565
R358 source.n179 source.n158 2.71565
R359 source.n198 source.n197 2.71565
R360 source.n54 source.n53 2.71565
R361 source.n36 source.n15 2.71565
R362 source.n124 source.n123 2.71565
R363 source.n106 source.n85 2.71565
R364 source.n250 source.n226 1.93989
R365 source.n264 source.n220 1.93989
R366 source.n180 source.n156 1.93989
R367 source.n194 source.n150 1.93989
R368 source.n50 source.n6 1.93989
R369 source.n37 source.n13 1.93989
R370 source.n120 source.n76 1.93989
R371 source.n107 source.n83 1.93989
R372 source.n212 source.t17 1.6505
R373 source.n212 source.t14 1.6505
R374 source.n210 source.t13 1.6505
R375 source.n210 source.t16 1.6505
R376 source.n142 source.t8 1.6505
R377 source.n142 source.t2 1.6505
R378 source.n140 source.t7 1.6505
R379 source.n140 source.t19 1.6505
R380 source.n66 source.t3 1.6505
R381 source.n66 source.t5 1.6505
R382 source.n68 source.t4 1.6505
R383 source.n68 source.t6 1.6505
R384 source.n136 source.t15 1.6505
R385 source.n136 source.t9 1.6505
R386 source.n138 source.t18 1.6505
R387 source.n138 source.t12 1.6505
R388 source.n255 source.n253 1.16414
R389 source.n263 source.n222 1.16414
R390 source.n185 source.n183 1.16414
R391 source.n193 source.n152 1.16414
R392 source.n49 source.n8 1.16414
R393 source.n41 source.n40 1.16414
R394 source.n119 source.n78 1.16414
R395 source.n111 source.n110 1.16414
R396 source.n135 source.n69 0.698776
R397 source.n211 source.n209 0.698776
R398 source.n139 source.n137 0.457397
R399 source.n137 source.n135 0.457397
R400 source.n69 source.n67 0.457397
R401 source.n67 source.n65 0.457397
R402 source.n143 source.n141 0.457397
R403 source.n209 source.n143 0.457397
R404 source.n213 source.n211 0.457397
R405 source.n279 source.n213 0.457397
R406 source.n254 source.n224 0.388379
R407 source.n260 source.n259 0.388379
R408 source.n184 source.n154 0.388379
R409 source.n190 source.n189 0.388379
R410 source.n46 source.n45 0.388379
R411 source.n12 source.n10 0.388379
R412 source.n116 source.n115 0.388379
R413 source.n82 source.n80 0.388379
R414 source source.n280 0.188
R415 source.n236 source.n231 0.155672
R416 source.n243 source.n231 0.155672
R417 source.n244 source.n243 0.155672
R418 source.n244 source.n227 0.155672
R419 source.n251 source.n227 0.155672
R420 source.n252 source.n251 0.155672
R421 source.n252 source.n223 0.155672
R422 source.n261 source.n223 0.155672
R423 source.n262 source.n261 0.155672
R424 source.n262 source.n219 0.155672
R425 source.n269 source.n219 0.155672
R426 source.n270 source.n269 0.155672
R427 source.n270 source.n215 0.155672
R428 source.n277 source.n215 0.155672
R429 source.n166 source.n161 0.155672
R430 source.n173 source.n161 0.155672
R431 source.n174 source.n173 0.155672
R432 source.n174 source.n157 0.155672
R433 source.n181 source.n157 0.155672
R434 source.n182 source.n181 0.155672
R435 source.n182 source.n153 0.155672
R436 source.n191 source.n153 0.155672
R437 source.n192 source.n191 0.155672
R438 source.n192 source.n149 0.155672
R439 source.n199 source.n149 0.155672
R440 source.n200 source.n199 0.155672
R441 source.n200 source.n145 0.155672
R442 source.n207 source.n145 0.155672
R443 source.n63 source.n1 0.155672
R444 source.n56 source.n1 0.155672
R445 source.n56 source.n55 0.155672
R446 source.n55 source.n5 0.155672
R447 source.n48 source.n5 0.155672
R448 source.n48 source.n47 0.155672
R449 source.n47 source.n9 0.155672
R450 source.n39 source.n9 0.155672
R451 source.n39 source.n38 0.155672
R452 source.n38 source.n14 0.155672
R453 source.n31 source.n14 0.155672
R454 source.n31 source.n30 0.155672
R455 source.n30 source.n18 0.155672
R456 source.n23 source.n18 0.155672
R457 source.n133 source.n71 0.155672
R458 source.n126 source.n71 0.155672
R459 source.n126 source.n125 0.155672
R460 source.n125 source.n75 0.155672
R461 source.n118 source.n75 0.155672
R462 source.n118 source.n117 0.155672
R463 source.n117 source.n79 0.155672
R464 source.n109 source.n79 0.155672
R465 source.n109 source.n108 0.155672
R466 source.n108 source.n84 0.155672
R467 source.n101 source.n84 0.155672
R468 source.n101 source.n100 0.155672
R469 source.n100 source.n88 0.155672
R470 source.n93 source.n88 0.155672
R471 drain_right.n60 drain_right.n0 289.615
R472 drain_right.n132 drain_right.n72 289.615
R473 drain_right.n20 drain_right.n19 185
R474 drain_right.n25 drain_right.n24 185
R475 drain_right.n27 drain_right.n26 185
R476 drain_right.n16 drain_right.n15 185
R477 drain_right.n33 drain_right.n32 185
R478 drain_right.n35 drain_right.n34 185
R479 drain_right.n12 drain_right.n11 185
R480 drain_right.n42 drain_right.n41 185
R481 drain_right.n43 drain_right.n10 185
R482 drain_right.n45 drain_right.n44 185
R483 drain_right.n8 drain_right.n7 185
R484 drain_right.n51 drain_right.n50 185
R485 drain_right.n53 drain_right.n52 185
R486 drain_right.n4 drain_right.n3 185
R487 drain_right.n59 drain_right.n58 185
R488 drain_right.n61 drain_right.n60 185
R489 drain_right.n133 drain_right.n132 185
R490 drain_right.n131 drain_right.n130 185
R491 drain_right.n76 drain_right.n75 185
R492 drain_right.n125 drain_right.n124 185
R493 drain_right.n123 drain_right.n122 185
R494 drain_right.n80 drain_right.n79 185
R495 drain_right.n117 drain_right.n116 185
R496 drain_right.n115 drain_right.n82 185
R497 drain_right.n114 drain_right.n113 185
R498 drain_right.n85 drain_right.n83 185
R499 drain_right.n108 drain_right.n107 185
R500 drain_right.n106 drain_right.n105 185
R501 drain_right.n89 drain_right.n88 185
R502 drain_right.n100 drain_right.n99 185
R503 drain_right.n98 drain_right.n97 185
R504 drain_right.n93 drain_right.n92 185
R505 drain_right.n21 drain_right.t7 149.524
R506 drain_right.n94 drain_right.t1 149.524
R507 drain_right.n25 drain_right.n19 104.615
R508 drain_right.n26 drain_right.n25 104.615
R509 drain_right.n26 drain_right.n15 104.615
R510 drain_right.n33 drain_right.n15 104.615
R511 drain_right.n34 drain_right.n33 104.615
R512 drain_right.n34 drain_right.n11 104.615
R513 drain_right.n42 drain_right.n11 104.615
R514 drain_right.n43 drain_right.n42 104.615
R515 drain_right.n44 drain_right.n43 104.615
R516 drain_right.n44 drain_right.n7 104.615
R517 drain_right.n51 drain_right.n7 104.615
R518 drain_right.n52 drain_right.n51 104.615
R519 drain_right.n52 drain_right.n3 104.615
R520 drain_right.n59 drain_right.n3 104.615
R521 drain_right.n60 drain_right.n59 104.615
R522 drain_right.n132 drain_right.n131 104.615
R523 drain_right.n131 drain_right.n75 104.615
R524 drain_right.n124 drain_right.n75 104.615
R525 drain_right.n124 drain_right.n123 104.615
R526 drain_right.n123 drain_right.n79 104.615
R527 drain_right.n116 drain_right.n79 104.615
R528 drain_right.n116 drain_right.n115 104.615
R529 drain_right.n115 drain_right.n114 104.615
R530 drain_right.n114 drain_right.n83 104.615
R531 drain_right.n107 drain_right.n83 104.615
R532 drain_right.n107 drain_right.n106 104.615
R533 drain_right.n106 drain_right.n88 104.615
R534 drain_right.n99 drain_right.n88 104.615
R535 drain_right.n99 drain_right.n98 104.615
R536 drain_right.n98 drain_right.n92 104.615
R537 drain_right.n71 drain_right.n69 60.0094
R538 drain_right.n68 drain_right.n67 59.8398
R539 drain_right.n71 drain_right.n70 59.5527
R540 drain_right.n66 drain_right.n65 59.5525
R541 drain_right.t7 drain_right.n19 52.3082
R542 drain_right.t1 drain_right.n92 52.3082
R543 drain_right.n66 drain_right.n64 46.9938
R544 drain_right.n137 drain_right.n136 46.5369
R545 drain_right drain_right.n68 28.7557
R546 drain_right.n45 drain_right.n10 13.1884
R547 drain_right.n117 drain_right.n82 13.1884
R548 drain_right.n41 drain_right.n40 12.8005
R549 drain_right.n46 drain_right.n8 12.8005
R550 drain_right.n118 drain_right.n80 12.8005
R551 drain_right.n113 drain_right.n84 12.8005
R552 drain_right.n39 drain_right.n12 12.0247
R553 drain_right.n50 drain_right.n49 12.0247
R554 drain_right.n122 drain_right.n121 12.0247
R555 drain_right.n112 drain_right.n85 12.0247
R556 drain_right.n36 drain_right.n35 11.249
R557 drain_right.n53 drain_right.n6 11.249
R558 drain_right.n125 drain_right.n78 11.249
R559 drain_right.n109 drain_right.n108 11.249
R560 drain_right.n32 drain_right.n14 10.4732
R561 drain_right.n54 drain_right.n4 10.4732
R562 drain_right.n126 drain_right.n76 10.4732
R563 drain_right.n105 drain_right.n87 10.4732
R564 drain_right.n21 drain_right.n20 10.2747
R565 drain_right.n94 drain_right.n93 10.2747
R566 drain_right.n31 drain_right.n16 9.69747
R567 drain_right.n58 drain_right.n57 9.69747
R568 drain_right.n130 drain_right.n129 9.69747
R569 drain_right.n104 drain_right.n89 9.69747
R570 drain_right.n64 drain_right.n63 9.45567
R571 drain_right.n136 drain_right.n135 9.45567
R572 drain_right.n63 drain_right.n62 9.3005
R573 drain_right.n2 drain_right.n1 9.3005
R574 drain_right.n57 drain_right.n56 9.3005
R575 drain_right.n55 drain_right.n54 9.3005
R576 drain_right.n6 drain_right.n5 9.3005
R577 drain_right.n49 drain_right.n48 9.3005
R578 drain_right.n47 drain_right.n46 9.3005
R579 drain_right.n23 drain_right.n22 9.3005
R580 drain_right.n18 drain_right.n17 9.3005
R581 drain_right.n29 drain_right.n28 9.3005
R582 drain_right.n31 drain_right.n30 9.3005
R583 drain_right.n14 drain_right.n13 9.3005
R584 drain_right.n37 drain_right.n36 9.3005
R585 drain_right.n39 drain_right.n38 9.3005
R586 drain_right.n40 drain_right.n9 9.3005
R587 drain_right.n96 drain_right.n95 9.3005
R588 drain_right.n91 drain_right.n90 9.3005
R589 drain_right.n102 drain_right.n101 9.3005
R590 drain_right.n104 drain_right.n103 9.3005
R591 drain_right.n87 drain_right.n86 9.3005
R592 drain_right.n110 drain_right.n109 9.3005
R593 drain_right.n112 drain_right.n111 9.3005
R594 drain_right.n84 drain_right.n81 9.3005
R595 drain_right.n135 drain_right.n134 9.3005
R596 drain_right.n74 drain_right.n73 9.3005
R597 drain_right.n129 drain_right.n128 9.3005
R598 drain_right.n127 drain_right.n126 9.3005
R599 drain_right.n78 drain_right.n77 9.3005
R600 drain_right.n121 drain_right.n120 9.3005
R601 drain_right.n119 drain_right.n118 9.3005
R602 drain_right.n28 drain_right.n27 8.92171
R603 drain_right.n61 drain_right.n2 8.92171
R604 drain_right.n133 drain_right.n74 8.92171
R605 drain_right.n101 drain_right.n100 8.92171
R606 drain_right.n24 drain_right.n18 8.14595
R607 drain_right.n62 drain_right.n0 8.14595
R608 drain_right.n134 drain_right.n72 8.14595
R609 drain_right.n97 drain_right.n91 8.14595
R610 drain_right.n23 drain_right.n20 7.3702
R611 drain_right.n96 drain_right.n93 7.3702
R612 drain_right drain_right.n137 5.88166
R613 drain_right.n24 drain_right.n23 5.81868
R614 drain_right.n64 drain_right.n0 5.81868
R615 drain_right.n136 drain_right.n72 5.81868
R616 drain_right.n97 drain_right.n96 5.81868
R617 drain_right.n27 drain_right.n18 5.04292
R618 drain_right.n62 drain_right.n61 5.04292
R619 drain_right.n134 drain_right.n133 5.04292
R620 drain_right.n100 drain_right.n91 5.04292
R621 drain_right.n28 drain_right.n16 4.26717
R622 drain_right.n58 drain_right.n2 4.26717
R623 drain_right.n130 drain_right.n74 4.26717
R624 drain_right.n101 drain_right.n89 4.26717
R625 drain_right.n32 drain_right.n31 3.49141
R626 drain_right.n57 drain_right.n4 3.49141
R627 drain_right.n129 drain_right.n76 3.49141
R628 drain_right.n105 drain_right.n104 3.49141
R629 drain_right.n22 drain_right.n21 2.84303
R630 drain_right.n95 drain_right.n94 2.84303
R631 drain_right.n35 drain_right.n14 2.71565
R632 drain_right.n54 drain_right.n53 2.71565
R633 drain_right.n126 drain_right.n125 2.71565
R634 drain_right.n108 drain_right.n87 2.71565
R635 drain_right.n36 drain_right.n12 1.93989
R636 drain_right.n50 drain_right.n6 1.93989
R637 drain_right.n122 drain_right.n78 1.93989
R638 drain_right.n109 drain_right.n85 1.93989
R639 drain_right.n67 drain_right.t6 1.6505
R640 drain_right.n67 drain_right.t3 1.6505
R641 drain_right.n65 drain_right.t5 1.6505
R642 drain_right.n65 drain_right.t8 1.6505
R643 drain_right.n69 drain_right.t4 1.6505
R644 drain_right.n69 drain_right.t2 1.6505
R645 drain_right.n70 drain_right.t0 1.6505
R646 drain_right.n70 drain_right.t9 1.6505
R647 drain_right.n41 drain_right.n39 1.16414
R648 drain_right.n49 drain_right.n8 1.16414
R649 drain_right.n121 drain_right.n80 1.16414
R650 drain_right.n113 drain_right.n112 1.16414
R651 drain_right.n137 drain_right.n71 0.457397
R652 drain_right.n40 drain_right.n10 0.388379
R653 drain_right.n46 drain_right.n45 0.388379
R654 drain_right.n118 drain_right.n117 0.388379
R655 drain_right.n84 drain_right.n82 0.388379
R656 drain_right.n22 drain_right.n17 0.155672
R657 drain_right.n29 drain_right.n17 0.155672
R658 drain_right.n30 drain_right.n29 0.155672
R659 drain_right.n30 drain_right.n13 0.155672
R660 drain_right.n37 drain_right.n13 0.155672
R661 drain_right.n38 drain_right.n37 0.155672
R662 drain_right.n38 drain_right.n9 0.155672
R663 drain_right.n47 drain_right.n9 0.155672
R664 drain_right.n48 drain_right.n47 0.155672
R665 drain_right.n48 drain_right.n5 0.155672
R666 drain_right.n55 drain_right.n5 0.155672
R667 drain_right.n56 drain_right.n55 0.155672
R668 drain_right.n56 drain_right.n1 0.155672
R669 drain_right.n63 drain_right.n1 0.155672
R670 drain_right.n135 drain_right.n73 0.155672
R671 drain_right.n128 drain_right.n73 0.155672
R672 drain_right.n128 drain_right.n127 0.155672
R673 drain_right.n127 drain_right.n77 0.155672
R674 drain_right.n120 drain_right.n77 0.155672
R675 drain_right.n120 drain_right.n119 0.155672
R676 drain_right.n119 drain_right.n81 0.155672
R677 drain_right.n111 drain_right.n81 0.155672
R678 drain_right.n111 drain_right.n110 0.155672
R679 drain_right.n110 drain_right.n86 0.155672
R680 drain_right.n103 drain_right.n86 0.155672
R681 drain_right.n103 drain_right.n102 0.155672
R682 drain_right.n102 drain_right.n90 0.155672
R683 drain_right.n95 drain_right.n90 0.155672
R684 drain_right.n68 drain_right.n66 0.0593781
R685 plus.n2 plus.t1 1647.93
R686 plus.n8 plus.t3 1647.93
R687 plus.n12 plus.t7 1647.93
R688 plus.n18 plus.t6 1647.93
R689 plus.n1 plus.t0 1602.65
R690 plus.n5 plus.t8 1602.65
R691 plus.n7 plus.t4 1602.65
R692 plus.n11 plus.t9 1602.65
R693 plus.n15 plus.t5 1602.65
R694 plus.n17 plus.t2 1602.65
R695 plus.n3 plus.n2 161.489
R696 plus.n13 plus.n12 161.489
R697 plus.n4 plus.n3 161.3
R698 plus.n6 plus.n0 161.3
R699 plus.n9 plus.n8 161.3
R700 plus.n14 plus.n13 161.3
R701 plus.n16 plus.n10 161.3
R702 plus.n19 plus.n18 161.3
R703 plus.n4 plus.n1 40.8975
R704 plus.n7 plus.n6 40.8975
R705 plus.n17 plus.n16 40.8975
R706 plus.n14 plus.n11 40.8975
R707 plus.n5 plus.n4 36.5157
R708 plus.n6 plus.n5 36.5157
R709 plus.n16 plus.n15 36.5157
R710 plus.n15 plus.n14 36.5157
R711 plus.n2 plus.n1 32.1338
R712 plus.n8 plus.n7 32.1338
R713 plus.n18 plus.n17 32.1338
R714 plus.n12 plus.n11 32.1338
R715 plus plus.n19 28.0729
R716 plus plus.n9 12.0933
R717 plus.n3 plus.n0 0.189894
R718 plus.n9 plus.n0 0.189894
R719 plus.n19 plus.n10 0.189894
R720 plus.n13 plus.n10 0.189894
R721 drain_left.n60 drain_left.n0 289.615
R722 drain_left.n129 drain_left.n69 289.615
R723 drain_left.n20 drain_left.n19 185
R724 drain_left.n25 drain_left.n24 185
R725 drain_left.n27 drain_left.n26 185
R726 drain_left.n16 drain_left.n15 185
R727 drain_left.n33 drain_left.n32 185
R728 drain_left.n35 drain_left.n34 185
R729 drain_left.n12 drain_left.n11 185
R730 drain_left.n42 drain_left.n41 185
R731 drain_left.n43 drain_left.n10 185
R732 drain_left.n45 drain_left.n44 185
R733 drain_left.n8 drain_left.n7 185
R734 drain_left.n51 drain_left.n50 185
R735 drain_left.n53 drain_left.n52 185
R736 drain_left.n4 drain_left.n3 185
R737 drain_left.n59 drain_left.n58 185
R738 drain_left.n61 drain_left.n60 185
R739 drain_left.n130 drain_left.n129 185
R740 drain_left.n128 drain_left.n127 185
R741 drain_left.n73 drain_left.n72 185
R742 drain_left.n122 drain_left.n121 185
R743 drain_left.n120 drain_left.n119 185
R744 drain_left.n77 drain_left.n76 185
R745 drain_left.n114 drain_left.n113 185
R746 drain_left.n112 drain_left.n79 185
R747 drain_left.n111 drain_left.n110 185
R748 drain_left.n82 drain_left.n80 185
R749 drain_left.n105 drain_left.n104 185
R750 drain_left.n103 drain_left.n102 185
R751 drain_left.n86 drain_left.n85 185
R752 drain_left.n97 drain_left.n96 185
R753 drain_left.n95 drain_left.n94 185
R754 drain_left.n90 drain_left.n89 185
R755 drain_left.n21 drain_left.t3 149.524
R756 drain_left.n91 drain_left.t8 149.524
R757 drain_left.n25 drain_left.n19 104.615
R758 drain_left.n26 drain_left.n25 104.615
R759 drain_left.n26 drain_left.n15 104.615
R760 drain_left.n33 drain_left.n15 104.615
R761 drain_left.n34 drain_left.n33 104.615
R762 drain_left.n34 drain_left.n11 104.615
R763 drain_left.n42 drain_left.n11 104.615
R764 drain_left.n43 drain_left.n42 104.615
R765 drain_left.n44 drain_left.n43 104.615
R766 drain_left.n44 drain_left.n7 104.615
R767 drain_left.n51 drain_left.n7 104.615
R768 drain_left.n52 drain_left.n51 104.615
R769 drain_left.n52 drain_left.n3 104.615
R770 drain_left.n59 drain_left.n3 104.615
R771 drain_left.n60 drain_left.n59 104.615
R772 drain_left.n129 drain_left.n128 104.615
R773 drain_left.n128 drain_left.n72 104.615
R774 drain_left.n121 drain_left.n72 104.615
R775 drain_left.n121 drain_left.n120 104.615
R776 drain_left.n120 drain_left.n76 104.615
R777 drain_left.n113 drain_left.n76 104.615
R778 drain_left.n113 drain_left.n112 104.615
R779 drain_left.n112 drain_left.n111 104.615
R780 drain_left.n111 drain_left.n80 104.615
R781 drain_left.n104 drain_left.n80 104.615
R782 drain_left.n104 drain_left.n103 104.615
R783 drain_left.n103 drain_left.n85 104.615
R784 drain_left.n96 drain_left.n85 104.615
R785 drain_left.n96 drain_left.n95 104.615
R786 drain_left.n95 drain_left.n89 104.615
R787 drain_left.n68 drain_left.n67 59.8398
R788 drain_left.n135 drain_left.n134 59.5527
R789 drain_left.n66 drain_left.n65 59.5525
R790 drain_left.n137 drain_left.n136 59.5525
R791 drain_left.t3 drain_left.n19 52.3082
R792 drain_left.t8 drain_left.n89 52.3082
R793 drain_left.n66 drain_left.n64 46.9938
R794 drain_left.n135 drain_left.n133 46.9938
R795 drain_left drain_left.n68 29.3089
R796 drain_left.n45 drain_left.n10 13.1884
R797 drain_left.n114 drain_left.n79 13.1884
R798 drain_left.n41 drain_left.n40 12.8005
R799 drain_left.n46 drain_left.n8 12.8005
R800 drain_left.n115 drain_left.n77 12.8005
R801 drain_left.n110 drain_left.n81 12.8005
R802 drain_left.n39 drain_left.n12 12.0247
R803 drain_left.n50 drain_left.n49 12.0247
R804 drain_left.n119 drain_left.n118 12.0247
R805 drain_left.n109 drain_left.n82 12.0247
R806 drain_left.n36 drain_left.n35 11.249
R807 drain_left.n53 drain_left.n6 11.249
R808 drain_left.n122 drain_left.n75 11.249
R809 drain_left.n106 drain_left.n105 11.249
R810 drain_left.n32 drain_left.n14 10.4732
R811 drain_left.n54 drain_left.n4 10.4732
R812 drain_left.n123 drain_left.n73 10.4732
R813 drain_left.n102 drain_left.n84 10.4732
R814 drain_left.n21 drain_left.n20 10.2747
R815 drain_left.n91 drain_left.n90 10.2747
R816 drain_left.n31 drain_left.n16 9.69747
R817 drain_left.n58 drain_left.n57 9.69747
R818 drain_left.n127 drain_left.n126 9.69747
R819 drain_left.n101 drain_left.n86 9.69747
R820 drain_left.n64 drain_left.n63 9.45567
R821 drain_left.n133 drain_left.n132 9.45567
R822 drain_left.n63 drain_left.n62 9.3005
R823 drain_left.n2 drain_left.n1 9.3005
R824 drain_left.n57 drain_left.n56 9.3005
R825 drain_left.n55 drain_left.n54 9.3005
R826 drain_left.n6 drain_left.n5 9.3005
R827 drain_left.n49 drain_left.n48 9.3005
R828 drain_left.n47 drain_left.n46 9.3005
R829 drain_left.n23 drain_left.n22 9.3005
R830 drain_left.n18 drain_left.n17 9.3005
R831 drain_left.n29 drain_left.n28 9.3005
R832 drain_left.n31 drain_left.n30 9.3005
R833 drain_left.n14 drain_left.n13 9.3005
R834 drain_left.n37 drain_left.n36 9.3005
R835 drain_left.n39 drain_left.n38 9.3005
R836 drain_left.n40 drain_left.n9 9.3005
R837 drain_left.n93 drain_left.n92 9.3005
R838 drain_left.n88 drain_left.n87 9.3005
R839 drain_left.n99 drain_left.n98 9.3005
R840 drain_left.n101 drain_left.n100 9.3005
R841 drain_left.n84 drain_left.n83 9.3005
R842 drain_left.n107 drain_left.n106 9.3005
R843 drain_left.n109 drain_left.n108 9.3005
R844 drain_left.n81 drain_left.n78 9.3005
R845 drain_left.n132 drain_left.n131 9.3005
R846 drain_left.n71 drain_left.n70 9.3005
R847 drain_left.n126 drain_left.n125 9.3005
R848 drain_left.n124 drain_left.n123 9.3005
R849 drain_left.n75 drain_left.n74 9.3005
R850 drain_left.n118 drain_left.n117 9.3005
R851 drain_left.n116 drain_left.n115 9.3005
R852 drain_left.n28 drain_left.n27 8.92171
R853 drain_left.n61 drain_left.n2 8.92171
R854 drain_left.n130 drain_left.n71 8.92171
R855 drain_left.n98 drain_left.n97 8.92171
R856 drain_left.n24 drain_left.n18 8.14595
R857 drain_left.n62 drain_left.n0 8.14595
R858 drain_left.n131 drain_left.n69 8.14595
R859 drain_left.n94 drain_left.n88 8.14595
R860 drain_left.n23 drain_left.n20 7.3702
R861 drain_left.n93 drain_left.n90 7.3702
R862 drain_left drain_left.n137 6.11011
R863 drain_left.n24 drain_left.n23 5.81868
R864 drain_left.n64 drain_left.n0 5.81868
R865 drain_left.n133 drain_left.n69 5.81868
R866 drain_left.n94 drain_left.n93 5.81868
R867 drain_left.n27 drain_left.n18 5.04292
R868 drain_left.n62 drain_left.n61 5.04292
R869 drain_left.n131 drain_left.n130 5.04292
R870 drain_left.n97 drain_left.n88 5.04292
R871 drain_left.n28 drain_left.n16 4.26717
R872 drain_left.n58 drain_left.n2 4.26717
R873 drain_left.n127 drain_left.n71 4.26717
R874 drain_left.n98 drain_left.n86 4.26717
R875 drain_left.n32 drain_left.n31 3.49141
R876 drain_left.n57 drain_left.n4 3.49141
R877 drain_left.n126 drain_left.n73 3.49141
R878 drain_left.n102 drain_left.n101 3.49141
R879 drain_left.n22 drain_left.n21 2.84303
R880 drain_left.n92 drain_left.n91 2.84303
R881 drain_left.n35 drain_left.n14 2.71565
R882 drain_left.n54 drain_left.n53 2.71565
R883 drain_left.n123 drain_left.n122 2.71565
R884 drain_left.n105 drain_left.n84 2.71565
R885 drain_left.n36 drain_left.n12 1.93989
R886 drain_left.n50 drain_left.n6 1.93989
R887 drain_left.n119 drain_left.n75 1.93989
R888 drain_left.n106 drain_left.n82 1.93989
R889 drain_left.n67 drain_left.t0 1.6505
R890 drain_left.n67 drain_left.t2 1.6505
R891 drain_left.n65 drain_left.t7 1.6505
R892 drain_left.n65 drain_left.t4 1.6505
R893 drain_left.n136 drain_left.t5 1.6505
R894 drain_left.n136 drain_left.t6 1.6505
R895 drain_left.n134 drain_left.t9 1.6505
R896 drain_left.n134 drain_left.t1 1.6505
R897 drain_left.n41 drain_left.n39 1.16414
R898 drain_left.n49 drain_left.n8 1.16414
R899 drain_left.n118 drain_left.n77 1.16414
R900 drain_left.n110 drain_left.n109 1.16414
R901 drain_left.n137 drain_left.n135 0.457397
R902 drain_left.n40 drain_left.n10 0.388379
R903 drain_left.n46 drain_left.n45 0.388379
R904 drain_left.n115 drain_left.n114 0.388379
R905 drain_left.n81 drain_left.n79 0.388379
R906 drain_left.n22 drain_left.n17 0.155672
R907 drain_left.n29 drain_left.n17 0.155672
R908 drain_left.n30 drain_left.n29 0.155672
R909 drain_left.n30 drain_left.n13 0.155672
R910 drain_left.n37 drain_left.n13 0.155672
R911 drain_left.n38 drain_left.n37 0.155672
R912 drain_left.n38 drain_left.n9 0.155672
R913 drain_left.n47 drain_left.n9 0.155672
R914 drain_left.n48 drain_left.n47 0.155672
R915 drain_left.n48 drain_left.n5 0.155672
R916 drain_left.n55 drain_left.n5 0.155672
R917 drain_left.n56 drain_left.n55 0.155672
R918 drain_left.n56 drain_left.n1 0.155672
R919 drain_left.n63 drain_left.n1 0.155672
R920 drain_left.n132 drain_left.n70 0.155672
R921 drain_left.n125 drain_left.n70 0.155672
R922 drain_left.n125 drain_left.n124 0.155672
R923 drain_left.n124 drain_left.n74 0.155672
R924 drain_left.n117 drain_left.n74 0.155672
R925 drain_left.n117 drain_left.n116 0.155672
R926 drain_left.n116 drain_left.n78 0.155672
R927 drain_left.n108 drain_left.n78 0.155672
R928 drain_left.n108 drain_left.n107 0.155672
R929 drain_left.n107 drain_left.n83 0.155672
R930 drain_left.n100 drain_left.n83 0.155672
R931 drain_left.n100 drain_left.n99 0.155672
R932 drain_left.n99 drain_left.n87 0.155672
R933 drain_left.n92 drain_left.n87 0.155672
R934 drain_left.n68 drain_left.n66 0.0593781
C0 source drain_right 24.9094f
C1 drain_left plus 3.19997f
C2 drain_right plus 0.283675f
C3 drain_left drain_right 0.662958f
C4 minus source 2.60852f
C5 minus plus 4.84055f
C6 minus drain_left 0.170748f
C7 source plus 2.62326f
C8 drain_left source 24.9218f
C9 minus drain_right 3.07501f
C10 drain_right a_n1352_n3288# 7.07924f
C11 drain_left a_n1352_n3288# 7.29344f
C12 source a_n1352_n3288# 5.958905f
C13 minus a_n1352_n3288# 5.212883f
C14 plus a_n1352_n3288# 7.28792f
C15 drain_left.n0 a_n1352_n3288# 0.044116f
C16 drain_left.n1 a_n1352_n3288# 0.033305f
C17 drain_left.n2 a_n1352_n3288# 0.017897f
C18 drain_left.n3 a_n1352_n3288# 0.042301f
C19 drain_left.n4 a_n1352_n3288# 0.018949f
C20 drain_left.n5 a_n1352_n3288# 0.033305f
C21 drain_left.n6 a_n1352_n3288# 0.017897f
C22 drain_left.n7 a_n1352_n3288# 0.042301f
C23 drain_left.n8 a_n1352_n3288# 0.018949f
C24 drain_left.n9 a_n1352_n3288# 0.033305f
C25 drain_left.n10 a_n1352_n3288# 0.018423f
C26 drain_left.n11 a_n1352_n3288# 0.042301f
C27 drain_left.n12 a_n1352_n3288# 0.018949f
C28 drain_left.n13 a_n1352_n3288# 0.033305f
C29 drain_left.n14 a_n1352_n3288# 0.017897f
C30 drain_left.n15 a_n1352_n3288# 0.042301f
C31 drain_left.n16 a_n1352_n3288# 0.018949f
C32 drain_left.n17 a_n1352_n3288# 0.033305f
C33 drain_left.n18 a_n1352_n3288# 0.017897f
C34 drain_left.n19 a_n1352_n3288# 0.031726f
C35 drain_left.n20 a_n1352_n3288# 0.029903f
C36 drain_left.t3 a_n1352_n3288# 0.071444f
C37 drain_left.n21 a_n1352_n3288# 0.240124f
C38 drain_left.n22 a_n1352_n3288# 1.68017f
C39 drain_left.n23 a_n1352_n3288# 0.017897f
C40 drain_left.n24 a_n1352_n3288# 0.018949f
C41 drain_left.n25 a_n1352_n3288# 0.042301f
C42 drain_left.n26 a_n1352_n3288# 0.042301f
C43 drain_left.n27 a_n1352_n3288# 0.018949f
C44 drain_left.n28 a_n1352_n3288# 0.017897f
C45 drain_left.n29 a_n1352_n3288# 0.033305f
C46 drain_left.n30 a_n1352_n3288# 0.033305f
C47 drain_left.n31 a_n1352_n3288# 0.017897f
C48 drain_left.n32 a_n1352_n3288# 0.018949f
C49 drain_left.n33 a_n1352_n3288# 0.042301f
C50 drain_left.n34 a_n1352_n3288# 0.042301f
C51 drain_left.n35 a_n1352_n3288# 0.018949f
C52 drain_left.n36 a_n1352_n3288# 0.017897f
C53 drain_left.n37 a_n1352_n3288# 0.033305f
C54 drain_left.n38 a_n1352_n3288# 0.033305f
C55 drain_left.n39 a_n1352_n3288# 0.017897f
C56 drain_left.n40 a_n1352_n3288# 0.017897f
C57 drain_left.n41 a_n1352_n3288# 0.018949f
C58 drain_left.n42 a_n1352_n3288# 0.042301f
C59 drain_left.n43 a_n1352_n3288# 0.042301f
C60 drain_left.n44 a_n1352_n3288# 0.042301f
C61 drain_left.n45 a_n1352_n3288# 0.018423f
C62 drain_left.n46 a_n1352_n3288# 0.017897f
C63 drain_left.n47 a_n1352_n3288# 0.033305f
C64 drain_left.n48 a_n1352_n3288# 0.033305f
C65 drain_left.n49 a_n1352_n3288# 0.017897f
C66 drain_left.n50 a_n1352_n3288# 0.018949f
C67 drain_left.n51 a_n1352_n3288# 0.042301f
C68 drain_left.n52 a_n1352_n3288# 0.042301f
C69 drain_left.n53 a_n1352_n3288# 0.018949f
C70 drain_left.n54 a_n1352_n3288# 0.017897f
C71 drain_left.n55 a_n1352_n3288# 0.033305f
C72 drain_left.n56 a_n1352_n3288# 0.033305f
C73 drain_left.n57 a_n1352_n3288# 0.017897f
C74 drain_left.n58 a_n1352_n3288# 0.018949f
C75 drain_left.n59 a_n1352_n3288# 0.042301f
C76 drain_left.n60 a_n1352_n3288# 0.086806f
C77 drain_left.n61 a_n1352_n3288# 0.018949f
C78 drain_left.n62 a_n1352_n3288# 0.017897f
C79 drain_left.n63 a_n1352_n3288# 0.071523f
C80 drain_left.n64 a_n1352_n3288# 0.072021f
C81 drain_left.t7 a_n1352_n3288# 0.315822f
C82 drain_left.t4 a_n1352_n3288# 0.315822f
C83 drain_left.n65 a_n1352_n3288# 2.81033f
C84 drain_left.n66 a_n1352_n3288# 0.456947f
C85 drain_left.t0 a_n1352_n3288# 0.315822f
C86 drain_left.t2 a_n1352_n3288# 0.315822f
C87 drain_left.n67 a_n1352_n3288# 2.81213f
C88 drain_left.n68 a_n1352_n3288# 1.81825f
C89 drain_left.n69 a_n1352_n3288# 0.044116f
C90 drain_left.n70 a_n1352_n3288# 0.033305f
C91 drain_left.n71 a_n1352_n3288# 0.017897f
C92 drain_left.n72 a_n1352_n3288# 0.042301f
C93 drain_left.n73 a_n1352_n3288# 0.018949f
C94 drain_left.n74 a_n1352_n3288# 0.033305f
C95 drain_left.n75 a_n1352_n3288# 0.017897f
C96 drain_left.n76 a_n1352_n3288# 0.042301f
C97 drain_left.n77 a_n1352_n3288# 0.018949f
C98 drain_left.n78 a_n1352_n3288# 0.033305f
C99 drain_left.n79 a_n1352_n3288# 0.018423f
C100 drain_left.n80 a_n1352_n3288# 0.042301f
C101 drain_left.n81 a_n1352_n3288# 0.017897f
C102 drain_left.n82 a_n1352_n3288# 0.018949f
C103 drain_left.n83 a_n1352_n3288# 0.033305f
C104 drain_left.n84 a_n1352_n3288# 0.017897f
C105 drain_left.n85 a_n1352_n3288# 0.042301f
C106 drain_left.n86 a_n1352_n3288# 0.018949f
C107 drain_left.n87 a_n1352_n3288# 0.033305f
C108 drain_left.n88 a_n1352_n3288# 0.017897f
C109 drain_left.n89 a_n1352_n3288# 0.031726f
C110 drain_left.n90 a_n1352_n3288# 0.029903f
C111 drain_left.t8 a_n1352_n3288# 0.071444f
C112 drain_left.n91 a_n1352_n3288# 0.240124f
C113 drain_left.n92 a_n1352_n3288# 1.68017f
C114 drain_left.n93 a_n1352_n3288# 0.017897f
C115 drain_left.n94 a_n1352_n3288# 0.018949f
C116 drain_left.n95 a_n1352_n3288# 0.042301f
C117 drain_left.n96 a_n1352_n3288# 0.042301f
C118 drain_left.n97 a_n1352_n3288# 0.018949f
C119 drain_left.n98 a_n1352_n3288# 0.017897f
C120 drain_left.n99 a_n1352_n3288# 0.033305f
C121 drain_left.n100 a_n1352_n3288# 0.033305f
C122 drain_left.n101 a_n1352_n3288# 0.017897f
C123 drain_left.n102 a_n1352_n3288# 0.018949f
C124 drain_left.n103 a_n1352_n3288# 0.042301f
C125 drain_left.n104 a_n1352_n3288# 0.042301f
C126 drain_left.n105 a_n1352_n3288# 0.018949f
C127 drain_left.n106 a_n1352_n3288# 0.017897f
C128 drain_left.n107 a_n1352_n3288# 0.033305f
C129 drain_left.n108 a_n1352_n3288# 0.033305f
C130 drain_left.n109 a_n1352_n3288# 0.017897f
C131 drain_left.n110 a_n1352_n3288# 0.018949f
C132 drain_left.n111 a_n1352_n3288# 0.042301f
C133 drain_left.n112 a_n1352_n3288# 0.042301f
C134 drain_left.n113 a_n1352_n3288# 0.042301f
C135 drain_left.n114 a_n1352_n3288# 0.018423f
C136 drain_left.n115 a_n1352_n3288# 0.017897f
C137 drain_left.n116 a_n1352_n3288# 0.033305f
C138 drain_left.n117 a_n1352_n3288# 0.033305f
C139 drain_left.n118 a_n1352_n3288# 0.017897f
C140 drain_left.n119 a_n1352_n3288# 0.018949f
C141 drain_left.n120 a_n1352_n3288# 0.042301f
C142 drain_left.n121 a_n1352_n3288# 0.042301f
C143 drain_left.n122 a_n1352_n3288# 0.018949f
C144 drain_left.n123 a_n1352_n3288# 0.017897f
C145 drain_left.n124 a_n1352_n3288# 0.033305f
C146 drain_left.n125 a_n1352_n3288# 0.033305f
C147 drain_left.n126 a_n1352_n3288# 0.017897f
C148 drain_left.n127 a_n1352_n3288# 0.018949f
C149 drain_left.n128 a_n1352_n3288# 0.042301f
C150 drain_left.n129 a_n1352_n3288# 0.086806f
C151 drain_left.n130 a_n1352_n3288# 0.018949f
C152 drain_left.n131 a_n1352_n3288# 0.017897f
C153 drain_left.n132 a_n1352_n3288# 0.071523f
C154 drain_left.n133 a_n1352_n3288# 0.072021f
C155 drain_left.t9 a_n1352_n3288# 0.315822f
C156 drain_left.t1 a_n1352_n3288# 0.315822f
C157 drain_left.n134 a_n1352_n3288# 2.81034f
C158 drain_left.n135 a_n1352_n3288# 0.486535f
C159 drain_left.t5 a_n1352_n3288# 0.315822f
C160 drain_left.t6 a_n1352_n3288# 0.315822f
C161 drain_left.n136 a_n1352_n3288# 2.81033f
C162 drain_left.n137 a_n1352_n3288# 0.650146f
C163 plus.n0 a_n1352_n3288# 0.058327f
C164 plus.t4 a_n1352_n3288# 0.395575f
C165 plus.t8 a_n1352_n3288# 0.395575f
C166 plus.t0 a_n1352_n3288# 0.395575f
C167 plus.n1 a_n1352_n3288# 0.162916f
C168 plus.t1 a_n1352_n3288# 0.400061f
C169 plus.n2 a_n1352_n3288# 0.179299f
C170 plus.n3 a_n1352_n3288# 0.128081f
C171 plus.n4 a_n1352_n3288# 0.020428f
C172 plus.n5 a_n1352_n3288# 0.162916f
C173 plus.n6 a_n1352_n3288# 0.020428f
C174 plus.n7 a_n1352_n3288# 0.162916f
C175 plus.t3 a_n1352_n3288# 0.400061f
C176 plus.n8 a_n1352_n3288# 0.179217f
C177 plus.n9 a_n1352_n3288# 0.645524f
C178 plus.n10 a_n1352_n3288# 0.058327f
C179 plus.t6 a_n1352_n3288# 0.400061f
C180 plus.t2 a_n1352_n3288# 0.395575f
C181 plus.t5 a_n1352_n3288# 0.395575f
C182 plus.t9 a_n1352_n3288# 0.395575f
C183 plus.n11 a_n1352_n3288# 0.162916f
C184 plus.t7 a_n1352_n3288# 0.400061f
C185 plus.n12 a_n1352_n3288# 0.179299f
C186 plus.n13 a_n1352_n3288# 0.128081f
C187 plus.n14 a_n1352_n3288# 0.020428f
C188 plus.n15 a_n1352_n3288# 0.162916f
C189 plus.n16 a_n1352_n3288# 0.020428f
C190 plus.n17 a_n1352_n3288# 0.162916f
C191 plus.n18 a_n1352_n3288# 0.179217f
C192 plus.n19 a_n1352_n3288# 1.58429f
C193 drain_right.n0 a_n1352_n3288# 0.044164f
C194 drain_right.n1 a_n1352_n3288# 0.033341f
C195 drain_right.n2 a_n1352_n3288# 0.017916f
C196 drain_right.n3 a_n1352_n3288# 0.042347f
C197 drain_right.n4 a_n1352_n3288# 0.01897f
C198 drain_right.n5 a_n1352_n3288# 0.033341f
C199 drain_right.n6 a_n1352_n3288# 0.017916f
C200 drain_right.n7 a_n1352_n3288# 0.042347f
C201 drain_right.n8 a_n1352_n3288# 0.01897f
C202 drain_right.n9 a_n1352_n3288# 0.033341f
C203 drain_right.n10 a_n1352_n3288# 0.018443f
C204 drain_right.n11 a_n1352_n3288# 0.042347f
C205 drain_right.n12 a_n1352_n3288# 0.01897f
C206 drain_right.n13 a_n1352_n3288# 0.033341f
C207 drain_right.n14 a_n1352_n3288# 0.017916f
C208 drain_right.n15 a_n1352_n3288# 0.042347f
C209 drain_right.n16 a_n1352_n3288# 0.01897f
C210 drain_right.n17 a_n1352_n3288# 0.033341f
C211 drain_right.n18 a_n1352_n3288# 0.017916f
C212 drain_right.n19 a_n1352_n3288# 0.03176f
C213 drain_right.n20 a_n1352_n3288# 0.029936f
C214 drain_right.t7 a_n1352_n3288# 0.071521f
C215 drain_right.n21 a_n1352_n3288# 0.240384f
C216 drain_right.n22 a_n1352_n3288# 1.68199f
C217 drain_right.n23 a_n1352_n3288# 0.017916f
C218 drain_right.n24 a_n1352_n3288# 0.01897f
C219 drain_right.n25 a_n1352_n3288# 0.042347f
C220 drain_right.n26 a_n1352_n3288# 0.042347f
C221 drain_right.n27 a_n1352_n3288# 0.01897f
C222 drain_right.n28 a_n1352_n3288# 0.017916f
C223 drain_right.n29 a_n1352_n3288# 0.033341f
C224 drain_right.n30 a_n1352_n3288# 0.033341f
C225 drain_right.n31 a_n1352_n3288# 0.017916f
C226 drain_right.n32 a_n1352_n3288# 0.01897f
C227 drain_right.n33 a_n1352_n3288# 0.042347f
C228 drain_right.n34 a_n1352_n3288# 0.042347f
C229 drain_right.n35 a_n1352_n3288# 0.01897f
C230 drain_right.n36 a_n1352_n3288# 0.017916f
C231 drain_right.n37 a_n1352_n3288# 0.033341f
C232 drain_right.n38 a_n1352_n3288# 0.033341f
C233 drain_right.n39 a_n1352_n3288# 0.017916f
C234 drain_right.n40 a_n1352_n3288# 0.017916f
C235 drain_right.n41 a_n1352_n3288# 0.01897f
C236 drain_right.n42 a_n1352_n3288# 0.042347f
C237 drain_right.n43 a_n1352_n3288# 0.042347f
C238 drain_right.n44 a_n1352_n3288# 0.042347f
C239 drain_right.n45 a_n1352_n3288# 0.018443f
C240 drain_right.n46 a_n1352_n3288# 0.017916f
C241 drain_right.n47 a_n1352_n3288# 0.033341f
C242 drain_right.n48 a_n1352_n3288# 0.033341f
C243 drain_right.n49 a_n1352_n3288# 0.017916f
C244 drain_right.n50 a_n1352_n3288# 0.01897f
C245 drain_right.n51 a_n1352_n3288# 0.042347f
C246 drain_right.n52 a_n1352_n3288# 0.042347f
C247 drain_right.n53 a_n1352_n3288# 0.01897f
C248 drain_right.n54 a_n1352_n3288# 0.017916f
C249 drain_right.n55 a_n1352_n3288# 0.033341f
C250 drain_right.n56 a_n1352_n3288# 0.033341f
C251 drain_right.n57 a_n1352_n3288# 0.017916f
C252 drain_right.n58 a_n1352_n3288# 0.01897f
C253 drain_right.n59 a_n1352_n3288# 0.042347f
C254 drain_right.n60 a_n1352_n3288# 0.0869f
C255 drain_right.n61 a_n1352_n3288# 0.01897f
C256 drain_right.n62 a_n1352_n3288# 0.017916f
C257 drain_right.n63 a_n1352_n3288# 0.0716f
C258 drain_right.n64 a_n1352_n3288# 0.072099f
C259 drain_right.t5 a_n1352_n3288# 0.316164f
C260 drain_right.t8 a_n1352_n3288# 0.316164f
C261 drain_right.n65 a_n1352_n3288# 2.81337f
C262 drain_right.n66 a_n1352_n3288# 0.457442f
C263 drain_right.t6 a_n1352_n3288# 0.316164f
C264 drain_right.t3 a_n1352_n3288# 0.316164f
C265 drain_right.n67 a_n1352_n3288# 2.81517f
C266 drain_right.n68 a_n1352_n3288# 1.75043f
C267 drain_right.t4 a_n1352_n3288# 0.316164f
C268 drain_right.t2 a_n1352_n3288# 0.316164f
C269 drain_right.n69 a_n1352_n3288# 2.81635f
C270 drain_right.t0 a_n1352_n3288# 0.316164f
C271 drain_right.t9 a_n1352_n3288# 0.316164f
C272 drain_right.n70 a_n1352_n3288# 2.81338f
C273 drain_right.n71 a_n1352_n3288# 0.766409f
C274 drain_right.n72 a_n1352_n3288# 0.044164f
C275 drain_right.n73 a_n1352_n3288# 0.033341f
C276 drain_right.n74 a_n1352_n3288# 0.017916f
C277 drain_right.n75 a_n1352_n3288# 0.042347f
C278 drain_right.n76 a_n1352_n3288# 0.01897f
C279 drain_right.n77 a_n1352_n3288# 0.033341f
C280 drain_right.n78 a_n1352_n3288# 0.017916f
C281 drain_right.n79 a_n1352_n3288# 0.042347f
C282 drain_right.n80 a_n1352_n3288# 0.01897f
C283 drain_right.n81 a_n1352_n3288# 0.033341f
C284 drain_right.n82 a_n1352_n3288# 0.018443f
C285 drain_right.n83 a_n1352_n3288# 0.042347f
C286 drain_right.n84 a_n1352_n3288# 0.017916f
C287 drain_right.n85 a_n1352_n3288# 0.01897f
C288 drain_right.n86 a_n1352_n3288# 0.033341f
C289 drain_right.n87 a_n1352_n3288# 0.017916f
C290 drain_right.n88 a_n1352_n3288# 0.042347f
C291 drain_right.n89 a_n1352_n3288# 0.01897f
C292 drain_right.n90 a_n1352_n3288# 0.033341f
C293 drain_right.n91 a_n1352_n3288# 0.017916f
C294 drain_right.n92 a_n1352_n3288# 0.03176f
C295 drain_right.n93 a_n1352_n3288# 0.029936f
C296 drain_right.t1 a_n1352_n3288# 0.071521f
C297 drain_right.n94 a_n1352_n3288# 0.240384f
C298 drain_right.n95 a_n1352_n3288# 1.68199f
C299 drain_right.n96 a_n1352_n3288# 0.017916f
C300 drain_right.n97 a_n1352_n3288# 0.01897f
C301 drain_right.n98 a_n1352_n3288# 0.042347f
C302 drain_right.n99 a_n1352_n3288# 0.042347f
C303 drain_right.n100 a_n1352_n3288# 0.01897f
C304 drain_right.n101 a_n1352_n3288# 0.017916f
C305 drain_right.n102 a_n1352_n3288# 0.033341f
C306 drain_right.n103 a_n1352_n3288# 0.033341f
C307 drain_right.n104 a_n1352_n3288# 0.017916f
C308 drain_right.n105 a_n1352_n3288# 0.01897f
C309 drain_right.n106 a_n1352_n3288# 0.042347f
C310 drain_right.n107 a_n1352_n3288# 0.042347f
C311 drain_right.n108 a_n1352_n3288# 0.01897f
C312 drain_right.n109 a_n1352_n3288# 0.017916f
C313 drain_right.n110 a_n1352_n3288# 0.033341f
C314 drain_right.n111 a_n1352_n3288# 0.033341f
C315 drain_right.n112 a_n1352_n3288# 0.017916f
C316 drain_right.n113 a_n1352_n3288# 0.01897f
C317 drain_right.n114 a_n1352_n3288# 0.042347f
C318 drain_right.n115 a_n1352_n3288# 0.042347f
C319 drain_right.n116 a_n1352_n3288# 0.042347f
C320 drain_right.n117 a_n1352_n3288# 0.018443f
C321 drain_right.n118 a_n1352_n3288# 0.017916f
C322 drain_right.n119 a_n1352_n3288# 0.033341f
C323 drain_right.n120 a_n1352_n3288# 0.033341f
C324 drain_right.n121 a_n1352_n3288# 0.017916f
C325 drain_right.n122 a_n1352_n3288# 0.01897f
C326 drain_right.n123 a_n1352_n3288# 0.042347f
C327 drain_right.n124 a_n1352_n3288# 0.042347f
C328 drain_right.n125 a_n1352_n3288# 0.01897f
C329 drain_right.n126 a_n1352_n3288# 0.017916f
C330 drain_right.n127 a_n1352_n3288# 0.033341f
C331 drain_right.n128 a_n1352_n3288# 0.033341f
C332 drain_right.n129 a_n1352_n3288# 0.017916f
C333 drain_right.n130 a_n1352_n3288# 0.01897f
C334 drain_right.n131 a_n1352_n3288# 0.042347f
C335 drain_right.n132 a_n1352_n3288# 0.0869f
C336 drain_right.n133 a_n1352_n3288# 0.01897f
C337 drain_right.n134 a_n1352_n3288# 0.017916f
C338 drain_right.n135 a_n1352_n3288# 0.0716f
C339 drain_right.n136 a_n1352_n3288# 0.071028f
C340 drain_right.n137 a_n1352_n3288# 0.381146f
C341 source.n0 a_n1352_n3288# 0.045455f
C342 source.n1 a_n1352_n3288# 0.034316f
C343 source.n2 a_n1352_n3288# 0.01844f
C344 source.n3 a_n1352_n3288# 0.043585f
C345 source.n4 a_n1352_n3288# 0.019524f
C346 source.n5 a_n1352_n3288# 0.034316f
C347 source.n6 a_n1352_n3288# 0.01844f
C348 source.n7 a_n1352_n3288# 0.043585f
C349 source.n8 a_n1352_n3288# 0.019524f
C350 source.n9 a_n1352_n3288# 0.034316f
C351 source.n10 a_n1352_n3288# 0.018982f
C352 source.n11 a_n1352_n3288# 0.043585f
C353 source.n12 a_n1352_n3288# 0.01844f
C354 source.n13 a_n1352_n3288# 0.019524f
C355 source.n14 a_n1352_n3288# 0.034316f
C356 source.n15 a_n1352_n3288# 0.01844f
C357 source.n16 a_n1352_n3288# 0.043585f
C358 source.n17 a_n1352_n3288# 0.019524f
C359 source.n18 a_n1352_n3288# 0.034316f
C360 source.n19 a_n1352_n3288# 0.01844f
C361 source.n20 a_n1352_n3288# 0.032689f
C362 source.n21 a_n1352_n3288# 0.030811f
C363 source.t1 a_n1352_n3288# 0.073612f
C364 source.n22 a_n1352_n3288# 0.247412f
C365 source.n23 a_n1352_n3288# 1.73116f
C366 source.n24 a_n1352_n3288# 0.01844f
C367 source.n25 a_n1352_n3288# 0.019524f
C368 source.n26 a_n1352_n3288# 0.043585f
C369 source.n27 a_n1352_n3288# 0.043585f
C370 source.n28 a_n1352_n3288# 0.019524f
C371 source.n29 a_n1352_n3288# 0.01844f
C372 source.n30 a_n1352_n3288# 0.034316f
C373 source.n31 a_n1352_n3288# 0.034316f
C374 source.n32 a_n1352_n3288# 0.01844f
C375 source.n33 a_n1352_n3288# 0.019524f
C376 source.n34 a_n1352_n3288# 0.043585f
C377 source.n35 a_n1352_n3288# 0.043585f
C378 source.n36 a_n1352_n3288# 0.019524f
C379 source.n37 a_n1352_n3288# 0.01844f
C380 source.n38 a_n1352_n3288# 0.034316f
C381 source.n39 a_n1352_n3288# 0.034316f
C382 source.n40 a_n1352_n3288# 0.01844f
C383 source.n41 a_n1352_n3288# 0.019524f
C384 source.n42 a_n1352_n3288# 0.043585f
C385 source.n43 a_n1352_n3288# 0.043585f
C386 source.n44 a_n1352_n3288# 0.043585f
C387 source.n45 a_n1352_n3288# 0.018982f
C388 source.n46 a_n1352_n3288# 0.01844f
C389 source.n47 a_n1352_n3288# 0.034316f
C390 source.n48 a_n1352_n3288# 0.034316f
C391 source.n49 a_n1352_n3288# 0.01844f
C392 source.n50 a_n1352_n3288# 0.019524f
C393 source.n51 a_n1352_n3288# 0.043585f
C394 source.n52 a_n1352_n3288# 0.043585f
C395 source.n53 a_n1352_n3288# 0.019524f
C396 source.n54 a_n1352_n3288# 0.01844f
C397 source.n55 a_n1352_n3288# 0.034316f
C398 source.n56 a_n1352_n3288# 0.034316f
C399 source.n57 a_n1352_n3288# 0.01844f
C400 source.n58 a_n1352_n3288# 0.019524f
C401 source.n59 a_n1352_n3288# 0.043585f
C402 source.n60 a_n1352_n3288# 0.089441f
C403 source.n61 a_n1352_n3288# 0.019524f
C404 source.n62 a_n1352_n3288# 0.01844f
C405 source.n63 a_n1352_n3288# 0.073693f
C406 source.n64 a_n1352_n3288# 0.049362f
C407 source.n65 a_n1352_n3288# 1.36539f
C408 source.t3 a_n1352_n3288# 0.325407f
C409 source.t5 a_n1352_n3288# 0.325407f
C410 source.n66 a_n1352_n3288# 2.78614f
C411 source.n67 a_n1352_n3288# 0.451874f
C412 source.t4 a_n1352_n3288# 0.325407f
C413 source.t6 a_n1352_n3288# 0.325407f
C414 source.n68 a_n1352_n3288# 2.78614f
C415 source.n69 a_n1352_n3288# 0.478564f
C416 source.n70 a_n1352_n3288# 0.045455f
C417 source.n71 a_n1352_n3288# 0.034316f
C418 source.n72 a_n1352_n3288# 0.01844f
C419 source.n73 a_n1352_n3288# 0.043585f
C420 source.n74 a_n1352_n3288# 0.019524f
C421 source.n75 a_n1352_n3288# 0.034316f
C422 source.n76 a_n1352_n3288# 0.01844f
C423 source.n77 a_n1352_n3288# 0.043585f
C424 source.n78 a_n1352_n3288# 0.019524f
C425 source.n79 a_n1352_n3288# 0.034316f
C426 source.n80 a_n1352_n3288# 0.018982f
C427 source.n81 a_n1352_n3288# 0.043585f
C428 source.n82 a_n1352_n3288# 0.01844f
C429 source.n83 a_n1352_n3288# 0.019524f
C430 source.n84 a_n1352_n3288# 0.034316f
C431 source.n85 a_n1352_n3288# 0.01844f
C432 source.n86 a_n1352_n3288# 0.043585f
C433 source.n87 a_n1352_n3288# 0.019524f
C434 source.n88 a_n1352_n3288# 0.034316f
C435 source.n89 a_n1352_n3288# 0.01844f
C436 source.n90 a_n1352_n3288# 0.032689f
C437 source.n91 a_n1352_n3288# 0.030811f
C438 source.t10 a_n1352_n3288# 0.073612f
C439 source.n92 a_n1352_n3288# 0.247412f
C440 source.n93 a_n1352_n3288# 1.73116f
C441 source.n94 a_n1352_n3288# 0.01844f
C442 source.n95 a_n1352_n3288# 0.019524f
C443 source.n96 a_n1352_n3288# 0.043585f
C444 source.n97 a_n1352_n3288# 0.043585f
C445 source.n98 a_n1352_n3288# 0.019524f
C446 source.n99 a_n1352_n3288# 0.01844f
C447 source.n100 a_n1352_n3288# 0.034316f
C448 source.n101 a_n1352_n3288# 0.034316f
C449 source.n102 a_n1352_n3288# 0.01844f
C450 source.n103 a_n1352_n3288# 0.019524f
C451 source.n104 a_n1352_n3288# 0.043585f
C452 source.n105 a_n1352_n3288# 0.043585f
C453 source.n106 a_n1352_n3288# 0.019524f
C454 source.n107 a_n1352_n3288# 0.01844f
C455 source.n108 a_n1352_n3288# 0.034316f
C456 source.n109 a_n1352_n3288# 0.034316f
C457 source.n110 a_n1352_n3288# 0.01844f
C458 source.n111 a_n1352_n3288# 0.019524f
C459 source.n112 a_n1352_n3288# 0.043585f
C460 source.n113 a_n1352_n3288# 0.043585f
C461 source.n114 a_n1352_n3288# 0.043585f
C462 source.n115 a_n1352_n3288# 0.018982f
C463 source.n116 a_n1352_n3288# 0.01844f
C464 source.n117 a_n1352_n3288# 0.034316f
C465 source.n118 a_n1352_n3288# 0.034316f
C466 source.n119 a_n1352_n3288# 0.01844f
C467 source.n120 a_n1352_n3288# 0.019524f
C468 source.n121 a_n1352_n3288# 0.043585f
C469 source.n122 a_n1352_n3288# 0.043585f
C470 source.n123 a_n1352_n3288# 0.019524f
C471 source.n124 a_n1352_n3288# 0.01844f
C472 source.n125 a_n1352_n3288# 0.034316f
C473 source.n126 a_n1352_n3288# 0.034316f
C474 source.n127 a_n1352_n3288# 0.01844f
C475 source.n128 a_n1352_n3288# 0.019524f
C476 source.n129 a_n1352_n3288# 0.043585f
C477 source.n130 a_n1352_n3288# 0.089441f
C478 source.n131 a_n1352_n3288# 0.019524f
C479 source.n132 a_n1352_n3288# 0.01844f
C480 source.n133 a_n1352_n3288# 0.073693f
C481 source.n134 a_n1352_n3288# 0.049362f
C482 source.n135 a_n1352_n3288# 0.15387f
C483 source.t15 a_n1352_n3288# 0.325407f
C484 source.t9 a_n1352_n3288# 0.325407f
C485 source.n136 a_n1352_n3288# 2.78614f
C486 source.n137 a_n1352_n3288# 0.451874f
C487 source.t18 a_n1352_n3288# 0.325407f
C488 source.t12 a_n1352_n3288# 0.325407f
C489 source.n138 a_n1352_n3288# 2.78614f
C490 source.n139 a_n1352_n3288# 2.27676f
C491 source.t7 a_n1352_n3288# 0.325407f
C492 source.t19 a_n1352_n3288# 0.325407f
C493 source.n140 a_n1352_n3288# 2.78612f
C494 source.n141 a_n1352_n3288# 2.27678f
C495 source.t8 a_n1352_n3288# 0.325407f
C496 source.t2 a_n1352_n3288# 0.325407f
C497 source.n142 a_n1352_n3288# 2.78612f
C498 source.n143 a_n1352_n3288# 0.451891f
C499 source.n144 a_n1352_n3288# 0.045455f
C500 source.n145 a_n1352_n3288# 0.034316f
C501 source.n146 a_n1352_n3288# 0.01844f
C502 source.n147 a_n1352_n3288# 0.043585f
C503 source.n148 a_n1352_n3288# 0.019524f
C504 source.n149 a_n1352_n3288# 0.034316f
C505 source.n150 a_n1352_n3288# 0.01844f
C506 source.n151 a_n1352_n3288# 0.043585f
C507 source.n152 a_n1352_n3288# 0.019524f
C508 source.n153 a_n1352_n3288# 0.034316f
C509 source.n154 a_n1352_n3288# 0.018982f
C510 source.n155 a_n1352_n3288# 0.043585f
C511 source.n156 a_n1352_n3288# 0.019524f
C512 source.n157 a_n1352_n3288# 0.034316f
C513 source.n158 a_n1352_n3288# 0.01844f
C514 source.n159 a_n1352_n3288# 0.043585f
C515 source.n160 a_n1352_n3288# 0.019524f
C516 source.n161 a_n1352_n3288# 0.034316f
C517 source.n162 a_n1352_n3288# 0.01844f
C518 source.n163 a_n1352_n3288# 0.032689f
C519 source.n164 a_n1352_n3288# 0.030811f
C520 source.t0 a_n1352_n3288# 0.073612f
C521 source.n165 a_n1352_n3288# 0.247412f
C522 source.n166 a_n1352_n3288# 1.73116f
C523 source.n167 a_n1352_n3288# 0.01844f
C524 source.n168 a_n1352_n3288# 0.019524f
C525 source.n169 a_n1352_n3288# 0.043585f
C526 source.n170 a_n1352_n3288# 0.043585f
C527 source.n171 a_n1352_n3288# 0.019524f
C528 source.n172 a_n1352_n3288# 0.01844f
C529 source.n173 a_n1352_n3288# 0.034316f
C530 source.n174 a_n1352_n3288# 0.034316f
C531 source.n175 a_n1352_n3288# 0.01844f
C532 source.n176 a_n1352_n3288# 0.019524f
C533 source.n177 a_n1352_n3288# 0.043585f
C534 source.n178 a_n1352_n3288# 0.043585f
C535 source.n179 a_n1352_n3288# 0.019524f
C536 source.n180 a_n1352_n3288# 0.01844f
C537 source.n181 a_n1352_n3288# 0.034316f
C538 source.n182 a_n1352_n3288# 0.034316f
C539 source.n183 a_n1352_n3288# 0.01844f
C540 source.n184 a_n1352_n3288# 0.01844f
C541 source.n185 a_n1352_n3288# 0.019524f
C542 source.n186 a_n1352_n3288# 0.043585f
C543 source.n187 a_n1352_n3288# 0.043585f
C544 source.n188 a_n1352_n3288# 0.043585f
C545 source.n189 a_n1352_n3288# 0.018982f
C546 source.n190 a_n1352_n3288# 0.01844f
C547 source.n191 a_n1352_n3288# 0.034316f
C548 source.n192 a_n1352_n3288# 0.034316f
C549 source.n193 a_n1352_n3288# 0.01844f
C550 source.n194 a_n1352_n3288# 0.019524f
C551 source.n195 a_n1352_n3288# 0.043585f
C552 source.n196 a_n1352_n3288# 0.043585f
C553 source.n197 a_n1352_n3288# 0.019524f
C554 source.n198 a_n1352_n3288# 0.01844f
C555 source.n199 a_n1352_n3288# 0.034316f
C556 source.n200 a_n1352_n3288# 0.034316f
C557 source.n201 a_n1352_n3288# 0.01844f
C558 source.n202 a_n1352_n3288# 0.019524f
C559 source.n203 a_n1352_n3288# 0.043585f
C560 source.n204 a_n1352_n3288# 0.089441f
C561 source.n205 a_n1352_n3288# 0.019524f
C562 source.n206 a_n1352_n3288# 0.01844f
C563 source.n207 a_n1352_n3288# 0.073693f
C564 source.n208 a_n1352_n3288# 0.049362f
C565 source.n209 a_n1352_n3288# 0.15387f
C566 source.t13 a_n1352_n3288# 0.325407f
C567 source.t16 a_n1352_n3288# 0.325407f
C568 source.n210 a_n1352_n3288# 2.78612f
C569 source.n211 a_n1352_n3288# 0.478581f
C570 source.t17 a_n1352_n3288# 0.325407f
C571 source.t14 a_n1352_n3288# 0.325407f
C572 source.n212 a_n1352_n3288# 2.78612f
C573 source.n213 a_n1352_n3288# 0.451891f
C574 source.n214 a_n1352_n3288# 0.045455f
C575 source.n215 a_n1352_n3288# 0.034316f
C576 source.n216 a_n1352_n3288# 0.01844f
C577 source.n217 a_n1352_n3288# 0.043585f
C578 source.n218 a_n1352_n3288# 0.019524f
C579 source.n219 a_n1352_n3288# 0.034316f
C580 source.n220 a_n1352_n3288# 0.01844f
C581 source.n221 a_n1352_n3288# 0.043585f
C582 source.n222 a_n1352_n3288# 0.019524f
C583 source.n223 a_n1352_n3288# 0.034316f
C584 source.n224 a_n1352_n3288# 0.018982f
C585 source.n225 a_n1352_n3288# 0.043585f
C586 source.n226 a_n1352_n3288# 0.019524f
C587 source.n227 a_n1352_n3288# 0.034316f
C588 source.n228 a_n1352_n3288# 0.01844f
C589 source.n229 a_n1352_n3288# 0.043585f
C590 source.n230 a_n1352_n3288# 0.019524f
C591 source.n231 a_n1352_n3288# 0.034316f
C592 source.n232 a_n1352_n3288# 0.01844f
C593 source.n233 a_n1352_n3288# 0.032689f
C594 source.n234 a_n1352_n3288# 0.030811f
C595 source.t11 a_n1352_n3288# 0.073612f
C596 source.n235 a_n1352_n3288# 0.247412f
C597 source.n236 a_n1352_n3288# 1.73116f
C598 source.n237 a_n1352_n3288# 0.01844f
C599 source.n238 a_n1352_n3288# 0.019524f
C600 source.n239 a_n1352_n3288# 0.043585f
C601 source.n240 a_n1352_n3288# 0.043585f
C602 source.n241 a_n1352_n3288# 0.019524f
C603 source.n242 a_n1352_n3288# 0.01844f
C604 source.n243 a_n1352_n3288# 0.034316f
C605 source.n244 a_n1352_n3288# 0.034316f
C606 source.n245 a_n1352_n3288# 0.01844f
C607 source.n246 a_n1352_n3288# 0.019524f
C608 source.n247 a_n1352_n3288# 0.043585f
C609 source.n248 a_n1352_n3288# 0.043585f
C610 source.n249 a_n1352_n3288# 0.019524f
C611 source.n250 a_n1352_n3288# 0.01844f
C612 source.n251 a_n1352_n3288# 0.034316f
C613 source.n252 a_n1352_n3288# 0.034316f
C614 source.n253 a_n1352_n3288# 0.01844f
C615 source.n254 a_n1352_n3288# 0.01844f
C616 source.n255 a_n1352_n3288# 0.019524f
C617 source.n256 a_n1352_n3288# 0.043585f
C618 source.n257 a_n1352_n3288# 0.043585f
C619 source.n258 a_n1352_n3288# 0.043585f
C620 source.n259 a_n1352_n3288# 0.018982f
C621 source.n260 a_n1352_n3288# 0.01844f
C622 source.n261 a_n1352_n3288# 0.034316f
C623 source.n262 a_n1352_n3288# 0.034316f
C624 source.n263 a_n1352_n3288# 0.01844f
C625 source.n264 a_n1352_n3288# 0.019524f
C626 source.n265 a_n1352_n3288# 0.043585f
C627 source.n266 a_n1352_n3288# 0.043585f
C628 source.n267 a_n1352_n3288# 0.019524f
C629 source.n268 a_n1352_n3288# 0.01844f
C630 source.n269 a_n1352_n3288# 0.034316f
C631 source.n270 a_n1352_n3288# 0.034316f
C632 source.n271 a_n1352_n3288# 0.01844f
C633 source.n272 a_n1352_n3288# 0.019524f
C634 source.n273 a_n1352_n3288# 0.043585f
C635 source.n274 a_n1352_n3288# 0.089441f
C636 source.n275 a_n1352_n3288# 0.019524f
C637 source.n276 a_n1352_n3288# 0.01844f
C638 source.n277 a_n1352_n3288# 0.073693f
C639 source.n278 a_n1352_n3288# 0.049362f
C640 source.n279 a_n1352_n3288# 0.31468f
C641 source.n280 a_n1352_n3288# 2.14744f
C642 minus.n0 a_n1352_n3288# 0.057141f
C643 minus.t8 a_n1352_n3288# 0.391926f
C644 minus.t9 a_n1352_n3288# 0.387531f
C645 minus.t0 a_n1352_n3288# 0.387531f
C646 minus.t5 a_n1352_n3288# 0.387531f
C647 minus.n1 a_n1352_n3288# 0.159603f
C648 minus.t7 a_n1352_n3288# 0.391926f
C649 minus.n2 a_n1352_n3288# 0.175653f
C650 minus.n3 a_n1352_n3288# 0.125476f
C651 minus.n4 a_n1352_n3288# 0.020013f
C652 minus.n5 a_n1352_n3288# 0.159603f
C653 minus.n6 a_n1352_n3288# 0.020013f
C654 minus.n7 a_n1352_n3288# 0.159603f
C655 minus.n8 a_n1352_n3288# 0.175573f
C656 minus.n9 a_n1352_n3288# 1.8431f
C657 minus.n10 a_n1352_n3288# 0.057141f
C658 minus.t3 a_n1352_n3288# 0.387531f
C659 minus.t1 a_n1352_n3288# 0.387531f
C660 minus.t4 a_n1352_n3288# 0.387531f
C661 minus.n11 a_n1352_n3288# 0.159603f
C662 minus.t2 a_n1352_n3288# 0.391926f
C663 minus.n12 a_n1352_n3288# 0.175653f
C664 minus.n13 a_n1352_n3288# 0.125476f
C665 minus.n14 a_n1352_n3288# 0.020013f
C666 minus.n15 a_n1352_n3288# 0.159603f
C667 minus.n16 a_n1352_n3288# 0.020013f
C668 minus.n17 a_n1352_n3288# 0.159603f
C669 minus.t6 a_n1352_n3288# 0.391926f
C670 minus.n18 a_n1352_n3288# 0.175573f
C671 minus.n19 a_n1352_n3288# 0.366742f
C672 minus.n20 a_n1352_n3288# 2.25439f
.ends

