* NGSPICE file created from diffpair307.ext - technology: sky130A

.subckt diffpair307 minus drain_right drain_left source plus
X0 a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X1 source.t31 plus.t0 drain_left.t12 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X2 source.t30 plus.t1 drain_left.t3 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 source.t29 plus.t2 drain_left.t8 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 source.t8 minus.t0 drain_right.t15 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X5 drain_left.t13 plus.t3 source.t28 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X6 source.t27 plus.t4 drain_left.t10 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X7 source.t26 plus.t5 drain_left.t4 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X8 drain_right.t14 minus.t1 source.t0 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X9 a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X10 drain_left.t9 plus.t6 source.t25 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X11 drain_right.t13 minus.t2 source.t11 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 drain_right.t12 minus.t3 source.t2 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 drain_right.t11 minus.t4 source.t6 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X14 source.t3 minus.t5 drain_right.t10 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 source.t24 plus.t7 drain_left.t6 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X16 drain_left.t2 plus.t8 source.t23 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X17 drain_left.t11 plus.t9 source.t22 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X18 drain_right.t9 minus.t6 source.t10 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X19 source.t12 minus.t7 drain_right.t8 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X20 source.t21 plus.t10 drain_left.t7 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X21 drain_left.t5 plus.t11 source.t20 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X22 drain_right.t7 minus.t8 source.t4 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X23 drain_left.t14 plus.t12 source.t19 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X24 drain_right.t6 minus.t9 source.t7 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X25 source.t9 minus.t10 drain_right.t5 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X26 drain_left.t0 plus.t13 source.t18 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X27 a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X28 source.t17 plus.t14 drain_left.t1 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X29 drain_left.t15 plus.t15 source.t16 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X30 source.t1 minus.t11 drain_right.t4 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X31 drain_right.t3 minus.t12 source.t5 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X32 source.t14 minus.t13 drain_right.t2 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X33 a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X34 source.t13 minus.t14 drain_right.t1 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X35 source.t15 minus.t15 drain_right.t0 a_n2570_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n7 plus.t5 287.065
R1 plus.n33 plus.t9 287.065
R2 plus.n24 plus.t8 262.69
R3 plus.n22 plus.t0 262.69
R4 plus.n2 plus.t12 262.69
R5 plus.n16 plus.t4 262.69
R6 plus.n4 plus.t11 262.69
R7 plus.n10 plus.t2 262.69
R8 plus.n6 plus.t13 262.69
R9 plus.n50 plus.t7 262.69
R10 plus.n48 plus.t15 262.69
R11 plus.n28 plus.t14 262.69
R12 plus.n42 plus.t3 262.69
R13 plus.n30 plus.t1 262.69
R14 plus.n36 plus.t6 262.69
R15 plus.n32 plus.t10 262.69
R16 plus.n9 plus.n8 161.3
R17 plus.n10 plus.n5 161.3
R18 plus.n12 plus.n11 161.3
R19 plus.n13 plus.n4 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n16 plus.n3 161.3
R22 plus.n18 plus.n17 161.3
R23 plus.n19 plus.n2 161.3
R24 plus.n21 plus.n20 161.3
R25 plus.n22 plus.n1 161.3
R26 plus.n23 plus.n0 161.3
R27 plus.n25 plus.n24 161.3
R28 plus.n35 plus.n34 161.3
R29 plus.n36 plus.n31 161.3
R30 plus.n38 plus.n37 161.3
R31 plus.n39 plus.n30 161.3
R32 plus.n41 plus.n40 161.3
R33 plus.n42 plus.n29 161.3
R34 plus.n44 plus.n43 161.3
R35 plus.n45 plus.n28 161.3
R36 plus.n47 plus.n46 161.3
R37 plus.n48 plus.n27 161.3
R38 plus.n49 plus.n26 161.3
R39 plus.n51 plus.n50 161.3
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus.n22 plus.n21 32.8641
R45 plus.n9 plus.n6 32.8641
R46 plus.n48 plus.n47 32.8641
R47 plus.n35 plus.n32 32.8641
R48 plus plus.n51 30.6202
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus.n23 plus.n22 10.955
R68 plus.n49 plus.n48 10.955
R69 plus plus.n25 10.027
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 drain_left.n9 drain_left.n7 68.0787
R93 drain_left.n5 drain_left.n3 68.0786
R94 drain_left.n2 drain_left.n0 68.0786
R95 drain_left.n11 drain_left.n10 67.1908
R96 drain_left.n9 drain_left.n8 67.1908
R97 drain_left.n13 drain_left.n12 67.1907
R98 drain_left.n5 drain_left.n4 67.1907
R99 drain_left.n2 drain_left.n1 67.1907
R100 drain_left drain_left.n6 28.5932
R101 drain_left drain_left.n13 6.54115
R102 drain_left.n3 drain_left.t7 3.3005
R103 drain_left.n3 drain_left.t11 3.3005
R104 drain_left.n4 drain_left.t3 3.3005
R105 drain_left.n4 drain_left.t9 3.3005
R106 drain_left.n1 drain_left.t1 3.3005
R107 drain_left.n1 drain_left.t13 3.3005
R108 drain_left.n0 drain_left.t6 3.3005
R109 drain_left.n0 drain_left.t15 3.3005
R110 drain_left.n12 drain_left.t12 3.3005
R111 drain_left.n12 drain_left.t2 3.3005
R112 drain_left.n10 drain_left.t10 3.3005
R113 drain_left.n10 drain_left.t14 3.3005
R114 drain_left.n8 drain_left.t8 3.3005
R115 drain_left.n8 drain_left.t5 3.3005
R116 drain_left.n7 drain_left.t4 3.3005
R117 drain_left.n7 drain_left.t0 3.3005
R118 drain_left.n11 drain_left.n9 0.888431
R119 drain_left.n13 drain_left.n11 0.888431
R120 drain_left.n6 drain_left.n5 0.389119
R121 drain_left.n6 drain_left.n2 0.389119
R122 source.n274 source.n248 289.615
R123 source.n236 source.n210 289.615
R124 source.n204 source.n178 289.615
R125 source.n166 source.n140 289.615
R126 source.n26 source.n0 289.615
R127 source.n64 source.n38 289.615
R128 source.n96 source.n70 289.615
R129 source.n134 source.n108 289.615
R130 source.n259 source.n258 185
R131 source.n256 source.n255 185
R132 source.n265 source.n264 185
R133 source.n267 source.n266 185
R134 source.n252 source.n251 185
R135 source.n273 source.n272 185
R136 source.n275 source.n274 185
R137 source.n221 source.n220 185
R138 source.n218 source.n217 185
R139 source.n227 source.n226 185
R140 source.n229 source.n228 185
R141 source.n214 source.n213 185
R142 source.n235 source.n234 185
R143 source.n237 source.n236 185
R144 source.n189 source.n188 185
R145 source.n186 source.n185 185
R146 source.n195 source.n194 185
R147 source.n197 source.n196 185
R148 source.n182 source.n181 185
R149 source.n203 source.n202 185
R150 source.n205 source.n204 185
R151 source.n151 source.n150 185
R152 source.n148 source.n147 185
R153 source.n157 source.n156 185
R154 source.n159 source.n158 185
R155 source.n144 source.n143 185
R156 source.n165 source.n164 185
R157 source.n167 source.n166 185
R158 source.n27 source.n26 185
R159 source.n25 source.n24 185
R160 source.n4 source.n3 185
R161 source.n19 source.n18 185
R162 source.n17 source.n16 185
R163 source.n8 source.n7 185
R164 source.n11 source.n10 185
R165 source.n65 source.n64 185
R166 source.n63 source.n62 185
R167 source.n42 source.n41 185
R168 source.n57 source.n56 185
R169 source.n55 source.n54 185
R170 source.n46 source.n45 185
R171 source.n49 source.n48 185
R172 source.n97 source.n96 185
R173 source.n95 source.n94 185
R174 source.n74 source.n73 185
R175 source.n89 source.n88 185
R176 source.n87 source.n86 185
R177 source.n78 source.n77 185
R178 source.n81 source.n80 185
R179 source.n135 source.n134 185
R180 source.n133 source.n132 185
R181 source.n112 source.n111 185
R182 source.n127 source.n126 185
R183 source.n125 source.n124 185
R184 source.n116 source.n115 185
R185 source.n119 source.n118 185
R186 source.t0 source.n257 147.661
R187 source.t1 source.n219 147.661
R188 source.t22 source.n187 147.661
R189 source.t24 source.n149 147.661
R190 source.t23 source.n9 147.661
R191 source.t26 source.n47 147.661
R192 source.t7 source.n79 147.661
R193 source.t14 source.n117 147.661
R194 source.n258 source.n255 104.615
R195 source.n265 source.n255 104.615
R196 source.n266 source.n265 104.615
R197 source.n266 source.n251 104.615
R198 source.n273 source.n251 104.615
R199 source.n274 source.n273 104.615
R200 source.n220 source.n217 104.615
R201 source.n227 source.n217 104.615
R202 source.n228 source.n227 104.615
R203 source.n228 source.n213 104.615
R204 source.n235 source.n213 104.615
R205 source.n236 source.n235 104.615
R206 source.n188 source.n185 104.615
R207 source.n195 source.n185 104.615
R208 source.n196 source.n195 104.615
R209 source.n196 source.n181 104.615
R210 source.n203 source.n181 104.615
R211 source.n204 source.n203 104.615
R212 source.n150 source.n147 104.615
R213 source.n157 source.n147 104.615
R214 source.n158 source.n157 104.615
R215 source.n158 source.n143 104.615
R216 source.n165 source.n143 104.615
R217 source.n166 source.n165 104.615
R218 source.n26 source.n25 104.615
R219 source.n25 source.n3 104.615
R220 source.n18 source.n3 104.615
R221 source.n18 source.n17 104.615
R222 source.n17 source.n7 104.615
R223 source.n10 source.n7 104.615
R224 source.n64 source.n63 104.615
R225 source.n63 source.n41 104.615
R226 source.n56 source.n41 104.615
R227 source.n56 source.n55 104.615
R228 source.n55 source.n45 104.615
R229 source.n48 source.n45 104.615
R230 source.n96 source.n95 104.615
R231 source.n95 source.n73 104.615
R232 source.n88 source.n73 104.615
R233 source.n88 source.n87 104.615
R234 source.n87 source.n77 104.615
R235 source.n80 source.n77 104.615
R236 source.n134 source.n133 104.615
R237 source.n133 source.n111 104.615
R238 source.n126 source.n111 104.615
R239 source.n126 source.n125 104.615
R240 source.n125 source.n115 104.615
R241 source.n118 source.n115 104.615
R242 source.n258 source.t0 52.3082
R243 source.n220 source.t1 52.3082
R244 source.n188 source.t22 52.3082
R245 source.n150 source.t24 52.3082
R246 source.n10 source.t23 52.3082
R247 source.n48 source.t26 52.3082
R248 source.n80 source.t7 52.3082
R249 source.n118 source.t14 52.3082
R250 source.n33 source.n32 50.512
R251 source.n35 source.n34 50.512
R252 source.n37 source.n36 50.512
R253 source.n103 source.n102 50.512
R254 source.n105 source.n104 50.512
R255 source.n107 source.n106 50.512
R256 source.n247 source.n246 50.5119
R257 source.n245 source.n244 50.5119
R258 source.n243 source.n242 50.5119
R259 source.n177 source.n176 50.5119
R260 source.n175 source.n174 50.5119
R261 source.n173 source.n172 50.5119
R262 source.n279 source.n278 32.1853
R263 source.n241 source.n240 32.1853
R264 source.n209 source.n208 32.1853
R265 source.n171 source.n170 32.1853
R266 source.n31 source.n30 32.1853
R267 source.n69 source.n68 32.1853
R268 source.n101 source.n100 32.1853
R269 source.n139 source.n138 32.1853
R270 source.n171 source.n139 17.6302
R271 source.n259 source.n257 15.6674
R272 source.n221 source.n219 15.6674
R273 source.n189 source.n187 15.6674
R274 source.n151 source.n149 15.6674
R275 source.n11 source.n9 15.6674
R276 source.n49 source.n47 15.6674
R277 source.n81 source.n79 15.6674
R278 source.n119 source.n117 15.6674
R279 source.n260 source.n256 12.8005
R280 source.n222 source.n218 12.8005
R281 source.n190 source.n186 12.8005
R282 source.n152 source.n148 12.8005
R283 source.n12 source.n8 12.8005
R284 source.n50 source.n46 12.8005
R285 source.n82 source.n78 12.8005
R286 source.n120 source.n116 12.8005
R287 source.n264 source.n263 12.0247
R288 source.n226 source.n225 12.0247
R289 source.n194 source.n193 12.0247
R290 source.n156 source.n155 12.0247
R291 source.n16 source.n15 12.0247
R292 source.n54 source.n53 12.0247
R293 source.n86 source.n85 12.0247
R294 source.n124 source.n123 12.0247
R295 source.n280 source.n31 11.9233
R296 source.n267 source.n254 11.249
R297 source.n229 source.n216 11.249
R298 source.n197 source.n184 11.249
R299 source.n159 source.n146 11.249
R300 source.n19 source.n6 11.249
R301 source.n57 source.n44 11.249
R302 source.n89 source.n76 11.249
R303 source.n127 source.n114 11.249
R304 source.n268 source.n252 10.4732
R305 source.n230 source.n214 10.4732
R306 source.n198 source.n182 10.4732
R307 source.n160 source.n144 10.4732
R308 source.n20 source.n4 10.4732
R309 source.n58 source.n42 10.4732
R310 source.n90 source.n74 10.4732
R311 source.n128 source.n112 10.4732
R312 source.n272 source.n271 9.69747
R313 source.n234 source.n233 9.69747
R314 source.n202 source.n201 9.69747
R315 source.n164 source.n163 9.69747
R316 source.n24 source.n23 9.69747
R317 source.n62 source.n61 9.69747
R318 source.n94 source.n93 9.69747
R319 source.n132 source.n131 9.69747
R320 source.n278 source.n277 9.45567
R321 source.n240 source.n239 9.45567
R322 source.n208 source.n207 9.45567
R323 source.n170 source.n169 9.45567
R324 source.n30 source.n29 9.45567
R325 source.n68 source.n67 9.45567
R326 source.n100 source.n99 9.45567
R327 source.n138 source.n137 9.45567
R328 source.n277 source.n276 9.3005
R329 source.n250 source.n249 9.3005
R330 source.n271 source.n270 9.3005
R331 source.n269 source.n268 9.3005
R332 source.n254 source.n253 9.3005
R333 source.n263 source.n262 9.3005
R334 source.n261 source.n260 9.3005
R335 source.n239 source.n238 9.3005
R336 source.n212 source.n211 9.3005
R337 source.n233 source.n232 9.3005
R338 source.n231 source.n230 9.3005
R339 source.n216 source.n215 9.3005
R340 source.n225 source.n224 9.3005
R341 source.n223 source.n222 9.3005
R342 source.n207 source.n206 9.3005
R343 source.n180 source.n179 9.3005
R344 source.n201 source.n200 9.3005
R345 source.n199 source.n198 9.3005
R346 source.n184 source.n183 9.3005
R347 source.n193 source.n192 9.3005
R348 source.n191 source.n190 9.3005
R349 source.n169 source.n168 9.3005
R350 source.n142 source.n141 9.3005
R351 source.n163 source.n162 9.3005
R352 source.n161 source.n160 9.3005
R353 source.n146 source.n145 9.3005
R354 source.n155 source.n154 9.3005
R355 source.n153 source.n152 9.3005
R356 source.n29 source.n28 9.3005
R357 source.n2 source.n1 9.3005
R358 source.n23 source.n22 9.3005
R359 source.n21 source.n20 9.3005
R360 source.n6 source.n5 9.3005
R361 source.n15 source.n14 9.3005
R362 source.n13 source.n12 9.3005
R363 source.n67 source.n66 9.3005
R364 source.n40 source.n39 9.3005
R365 source.n61 source.n60 9.3005
R366 source.n59 source.n58 9.3005
R367 source.n44 source.n43 9.3005
R368 source.n53 source.n52 9.3005
R369 source.n51 source.n50 9.3005
R370 source.n99 source.n98 9.3005
R371 source.n72 source.n71 9.3005
R372 source.n93 source.n92 9.3005
R373 source.n91 source.n90 9.3005
R374 source.n76 source.n75 9.3005
R375 source.n85 source.n84 9.3005
R376 source.n83 source.n82 9.3005
R377 source.n137 source.n136 9.3005
R378 source.n110 source.n109 9.3005
R379 source.n131 source.n130 9.3005
R380 source.n129 source.n128 9.3005
R381 source.n114 source.n113 9.3005
R382 source.n123 source.n122 9.3005
R383 source.n121 source.n120 9.3005
R384 source.n275 source.n250 8.92171
R385 source.n237 source.n212 8.92171
R386 source.n205 source.n180 8.92171
R387 source.n167 source.n142 8.92171
R388 source.n27 source.n2 8.92171
R389 source.n65 source.n40 8.92171
R390 source.n97 source.n72 8.92171
R391 source.n135 source.n110 8.92171
R392 source.n276 source.n248 8.14595
R393 source.n238 source.n210 8.14595
R394 source.n206 source.n178 8.14595
R395 source.n168 source.n140 8.14595
R396 source.n28 source.n0 8.14595
R397 source.n66 source.n38 8.14595
R398 source.n98 source.n70 8.14595
R399 source.n136 source.n108 8.14595
R400 source.n278 source.n248 5.81868
R401 source.n240 source.n210 5.81868
R402 source.n208 source.n178 5.81868
R403 source.n170 source.n140 5.81868
R404 source.n30 source.n0 5.81868
R405 source.n68 source.n38 5.81868
R406 source.n100 source.n70 5.81868
R407 source.n138 source.n108 5.81868
R408 source.n280 source.n279 5.7074
R409 source.n276 source.n275 5.04292
R410 source.n238 source.n237 5.04292
R411 source.n206 source.n205 5.04292
R412 source.n168 source.n167 5.04292
R413 source.n28 source.n27 5.04292
R414 source.n66 source.n65 5.04292
R415 source.n98 source.n97 5.04292
R416 source.n136 source.n135 5.04292
R417 source.n261 source.n257 4.38594
R418 source.n223 source.n219 4.38594
R419 source.n191 source.n187 4.38594
R420 source.n153 source.n149 4.38594
R421 source.n13 source.n9 4.38594
R422 source.n51 source.n47 4.38594
R423 source.n83 source.n79 4.38594
R424 source.n121 source.n117 4.38594
R425 source.n272 source.n250 4.26717
R426 source.n234 source.n212 4.26717
R427 source.n202 source.n180 4.26717
R428 source.n164 source.n142 4.26717
R429 source.n24 source.n2 4.26717
R430 source.n62 source.n40 4.26717
R431 source.n94 source.n72 4.26717
R432 source.n132 source.n110 4.26717
R433 source.n271 source.n252 3.49141
R434 source.n233 source.n214 3.49141
R435 source.n201 source.n182 3.49141
R436 source.n163 source.n144 3.49141
R437 source.n23 source.n4 3.49141
R438 source.n61 source.n42 3.49141
R439 source.n93 source.n74 3.49141
R440 source.n131 source.n112 3.49141
R441 source.n246 source.t2 3.3005
R442 source.n246 source.t3 3.3005
R443 source.n244 source.t4 3.3005
R444 source.n244 source.t9 3.3005
R445 source.n242 source.t5 3.3005
R446 source.n242 source.t12 3.3005
R447 source.n176 source.t25 3.3005
R448 source.n176 source.t21 3.3005
R449 source.n174 source.t28 3.3005
R450 source.n174 source.t30 3.3005
R451 source.n172 source.t16 3.3005
R452 source.n172 source.t17 3.3005
R453 source.n32 source.t19 3.3005
R454 source.n32 source.t31 3.3005
R455 source.n34 source.t20 3.3005
R456 source.n34 source.t27 3.3005
R457 source.n36 source.t18 3.3005
R458 source.n36 source.t29 3.3005
R459 source.n102 source.t10 3.3005
R460 source.n102 source.t8 3.3005
R461 source.n104 source.t6 3.3005
R462 source.n104 source.t13 3.3005
R463 source.n106 source.t11 3.3005
R464 source.n106 source.t15 3.3005
R465 source.n268 source.n267 2.71565
R466 source.n230 source.n229 2.71565
R467 source.n198 source.n197 2.71565
R468 source.n160 source.n159 2.71565
R469 source.n20 source.n19 2.71565
R470 source.n58 source.n57 2.71565
R471 source.n90 source.n89 2.71565
R472 source.n128 source.n127 2.71565
R473 source.n264 source.n254 1.93989
R474 source.n226 source.n216 1.93989
R475 source.n194 source.n184 1.93989
R476 source.n156 source.n146 1.93989
R477 source.n16 source.n6 1.93989
R478 source.n54 source.n44 1.93989
R479 source.n86 source.n76 1.93989
R480 source.n124 source.n114 1.93989
R481 source.n263 source.n256 1.16414
R482 source.n225 source.n218 1.16414
R483 source.n193 source.n186 1.16414
R484 source.n155 source.n148 1.16414
R485 source.n15 source.n8 1.16414
R486 source.n53 source.n46 1.16414
R487 source.n85 source.n78 1.16414
R488 source.n123 source.n116 1.16414
R489 source.n139 source.n107 0.888431
R490 source.n107 source.n105 0.888431
R491 source.n105 source.n103 0.888431
R492 source.n103 source.n101 0.888431
R493 source.n69 source.n37 0.888431
R494 source.n37 source.n35 0.888431
R495 source.n35 source.n33 0.888431
R496 source.n33 source.n31 0.888431
R497 source.n173 source.n171 0.888431
R498 source.n175 source.n173 0.888431
R499 source.n177 source.n175 0.888431
R500 source.n209 source.n177 0.888431
R501 source.n243 source.n241 0.888431
R502 source.n245 source.n243 0.888431
R503 source.n247 source.n245 0.888431
R504 source.n279 source.n247 0.888431
R505 source.n101 source.n69 0.470328
R506 source.n241 source.n209 0.470328
R507 source.n260 source.n259 0.388379
R508 source.n222 source.n221 0.388379
R509 source.n190 source.n189 0.388379
R510 source.n152 source.n151 0.388379
R511 source.n12 source.n11 0.388379
R512 source.n50 source.n49 0.388379
R513 source.n82 source.n81 0.388379
R514 source.n120 source.n119 0.388379
R515 source source.n280 0.188
R516 source.n262 source.n261 0.155672
R517 source.n262 source.n253 0.155672
R518 source.n269 source.n253 0.155672
R519 source.n270 source.n269 0.155672
R520 source.n270 source.n249 0.155672
R521 source.n277 source.n249 0.155672
R522 source.n224 source.n223 0.155672
R523 source.n224 source.n215 0.155672
R524 source.n231 source.n215 0.155672
R525 source.n232 source.n231 0.155672
R526 source.n232 source.n211 0.155672
R527 source.n239 source.n211 0.155672
R528 source.n192 source.n191 0.155672
R529 source.n192 source.n183 0.155672
R530 source.n199 source.n183 0.155672
R531 source.n200 source.n199 0.155672
R532 source.n200 source.n179 0.155672
R533 source.n207 source.n179 0.155672
R534 source.n154 source.n153 0.155672
R535 source.n154 source.n145 0.155672
R536 source.n161 source.n145 0.155672
R537 source.n162 source.n161 0.155672
R538 source.n162 source.n141 0.155672
R539 source.n169 source.n141 0.155672
R540 source.n29 source.n1 0.155672
R541 source.n22 source.n1 0.155672
R542 source.n22 source.n21 0.155672
R543 source.n21 source.n5 0.155672
R544 source.n14 source.n5 0.155672
R545 source.n14 source.n13 0.155672
R546 source.n67 source.n39 0.155672
R547 source.n60 source.n39 0.155672
R548 source.n60 source.n59 0.155672
R549 source.n59 source.n43 0.155672
R550 source.n52 source.n43 0.155672
R551 source.n52 source.n51 0.155672
R552 source.n99 source.n71 0.155672
R553 source.n92 source.n71 0.155672
R554 source.n92 source.n91 0.155672
R555 source.n91 source.n75 0.155672
R556 source.n84 source.n75 0.155672
R557 source.n84 source.n83 0.155672
R558 source.n137 source.n109 0.155672
R559 source.n130 source.n109 0.155672
R560 source.n130 source.n129 0.155672
R561 source.n129 source.n113 0.155672
R562 source.n122 source.n113 0.155672
R563 source.n122 source.n121 0.155672
R564 minus.n7 minus.t9 287.065
R565 minus.n33 minus.t11 287.065
R566 minus.n6 minus.t0 262.69
R567 minus.n10 minus.t6 262.69
R568 minus.n12 minus.t14 262.69
R569 minus.n16 minus.t4 262.69
R570 minus.n18 minus.t15 262.69
R571 minus.n22 minus.t2 262.69
R572 minus.n24 minus.t13 262.69
R573 minus.n32 minus.t12 262.69
R574 minus.n36 minus.t7 262.69
R575 minus.n38 minus.t8 262.69
R576 minus.n42 minus.t10 262.69
R577 minus.n44 minus.t3 262.69
R578 minus.n48 minus.t5 262.69
R579 minus.n50 minus.t1 262.69
R580 minus.n25 minus.n24 161.3
R581 minus.n23 minus.n0 161.3
R582 minus.n22 minus.n21 161.3
R583 minus.n20 minus.n1 161.3
R584 minus.n19 minus.n18 161.3
R585 minus.n17 minus.n2 161.3
R586 minus.n16 minus.n15 161.3
R587 minus.n14 minus.n3 161.3
R588 minus.n13 minus.n12 161.3
R589 minus.n11 minus.n4 161.3
R590 minus.n10 minus.n9 161.3
R591 minus.n8 minus.n5 161.3
R592 minus.n51 minus.n50 161.3
R593 minus.n49 minus.n26 161.3
R594 minus.n48 minus.n47 161.3
R595 minus.n46 minus.n27 161.3
R596 minus.n45 minus.n44 161.3
R597 minus.n43 minus.n28 161.3
R598 minus.n42 minus.n41 161.3
R599 minus.n40 minus.n29 161.3
R600 minus.n39 minus.n38 161.3
R601 minus.n37 minus.n30 161.3
R602 minus.n36 minus.n35 161.3
R603 minus.n34 minus.n31 161.3
R604 minus.n8 minus.n7 44.9377
R605 minus.n34 minus.n33 44.9377
R606 minus.n24 minus.n23 37.246
R607 minus.n50 minus.n49 37.246
R608 minus.n52 minus.n25 34.4664
R609 minus.n6 minus.n5 32.8641
R610 minus.n22 minus.n1 32.8641
R611 minus.n32 minus.n31 32.8641
R612 minus.n48 minus.n27 32.8641
R613 minus.n11 minus.n10 28.4823
R614 minus.n18 minus.n17 28.4823
R615 minus.n37 minus.n36 28.4823
R616 minus.n44 minus.n43 28.4823
R617 minus.n16 minus.n3 24.1005
R618 minus.n12 minus.n3 24.1005
R619 minus.n38 minus.n29 24.1005
R620 minus.n42 minus.n29 24.1005
R621 minus.n12 minus.n11 19.7187
R622 minus.n17 minus.n16 19.7187
R623 minus.n38 minus.n37 19.7187
R624 minus.n43 minus.n42 19.7187
R625 minus.n7 minus.n6 17.0522
R626 minus.n33 minus.n32 17.0522
R627 minus.n10 minus.n5 15.3369
R628 minus.n18 minus.n1 15.3369
R629 minus.n36 minus.n31 15.3369
R630 minus.n44 minus.n27 15.3369
R631 minus.n23 minus.n22 10.955
R632 minus.n49 minus.n48 10.955
R633 minus.n52 minus.n51 6.6558
R634 minus.n25 minus.n0 0.189894
R635 minus.n21 minus.n0 0.189894
R636 minus.n21 minus.n20 0.189894
R637 minus.n20 minus.n19 0.189894
R638 minus.n19 minus.n2 0.189894
R639 minus.n15 minus.n2 0.189894
R640 minus.n15 minus.n14 0.189894
R641 minus.n14 minus.n13 0.189894
R642 minus.n13 minus.n4 0.189894
R643 minus.n9 minus.n4 0.189894
R644 minus.n9 minus.n8 0.189894
R645 minus.n35 minus.n34 0.189894
R646 minus.n35 minus.n30 0.189894
R647 minus.n39 minus.n30 0.189894
R648 minus.n40 minus.n39 0.189894
R649 minus.n41 minus.n40 0.189894
R650 minus.n41 minus.n28 0.189894
R651 minus.n45 minus.n28 0.189894
R652 minus.n46 minus.n45 0.189894
R653 minus.n47 minus.n46 0.189894
R654 minus.n47 minus.n26 0.189894
R655 minus.n51 minus.n26 0.189894
R656 minus minus.n52 0.188
R657 drain_right.n9 drain_right.n7 68.0786
R658 drain_right.n5 drain_right.n3 68.0786
R659 drain_right.n2 drain_right.n0 68.0786
R660 drain_right.n9 drain_right.n8 67.1908
R661 drain_right.n11 drain_right.n10 67.1908
R662 drain_right.n13 drain_right.n12 67.1908
R663 drain_right.n5 drain_right.n4 67.1907
R664 drain_right.n2 drain_right.n1 67.1907
R665 drain_right drain_right.n6 28.0399
R666 drain_right drain_right.n13 6.54115
R667 drain_right.n3 drain_right.t10 3.3005
R668 drain_right.n3 drain_right.t14 3.3005
R669 drain_right.n4 drain_right.t5 3.3005
R670 drain_right.n4 drain_right.t12 3.3005
R671 drain_right.n1 drain_right.t8 3.3005
R672 drain_right.n1 drain_right.t7 3.3005
R673 drain_right.n0 drain_right.t4 3.3005
R674 drain_right.n0 drain_right.t3 3.3005
R675 drain_right.n7 drain_right.t15 3.3005
R676 drain_right.n7 drain_right.t6 3.3005
R677 drain_right.n8 drain_right.t1 3.3005
R678 drain_right.n8 drain_right.t9 3.3005
R679 drain_right.n10 drain_right.t0 3.3005
R680 drain_right.n10 drain_right.t11 3.3005
R681 drain_right.n12 drain_right.t2 3.3005
R682 drain_right.n12 drain_right.t13 3.3005
R683 drain_right.n13 drain_right.n11 0.888431
R684 drain_right.n11 drain_right.n9 0.888431
R685 drain_right.n6 drain_right.n5 0.389119
R686 drain_right.n6 drain_right.n2 0.389119
C0 minus plus 5.23905f
C1 source drain_right 11.6322f
C2 plus source 5.7896f
C3 drain_left drain_right 1.34352f
C4 plus drain_left 5.67267f
C5 minus source 5.77558f
C6 plus drain_right 0.410755f
C7 minus drain_left 0.172697f
C8 drain_left source 11.6299f
C9 minus drain_right 5.41803f
C10 drain_right a_n2570_n2088# 5.62864f
C11 drain_left a_n2570_n2088# 6.0053f
C12 source a_n2570_n2088# 5.671676f
C13 minus a_n2570_n2088# 9.738084f
C14 plus a_n2570_n2088# 11.21367f
C15 drain_right.t4 a_n2570_n2088# 0.127556f
C16 drain_right.t3 a_n2570_n2088# 0.127556f
C17 drain_right.n0 a_n2570_n2088# 1.06881f
C18 drain_right.t8 a_n2570_n2088# 0.127556f
C19 drain_right.t7 a_n2570_n2088# 0.127556f
C20 drain_right.n1 a_n2570_n2088# 1.06382f
C21 drain_right.n2 a_n2570_n2088# 0.708749f
C22 drain_right.t10 a_n2570_n2088# 0.127556f
C23 drain_right.t14 a_n2570_n2088# 0.127556f
C24 drain_right.n3 a_n2570_n2088# 1.06881f
C25 drain_right.t5 a_n2570_n2088# 0.127556f
C26 drain_right.t12 a_n2570_n2088# 0.127556f
C27 drain_right.n4 a_n2570_n2088# 1.06382f
C28 drain_right.n5 a_n2570_n2088# 0.708748f
C29 drain_right.n6 a_n2570_n2088# 1.13671f
C30 drain_right.t15 a_n2570_n2088# 0.127556f
C31 drain_right.t6 a_n2570_n2088# 0.127556f
C32 drain_right.n7 a_n2570_n2088# 1.06881f
C33 drain_right.t1 a_n2570_n2088# 0.127556f
C34 drain_right.t9 a_n2570_n2088# 0.127556f
C35 drain_right.n8 a_n2570_n2088# 1.06382f
C36 drain_right.n9 a_n2570_n2088# 0.750422f
C37 drain_right.t0 a_n2570_n2088# 0.127556f
C38 drain_right.t11 a_n2570_n2088# 0.127556f
C39 drain_right.n10 a_n2570_n2088# 1.06382f
C40 drain_right.n11 a_n2570_n2088# 0.372289f
C41 drain_right.t2 a_n2570_n2088# 0.127556f
C42 drain_right.t13 a_n2570_n2088# 0.127556f
C43 drain_right.n12 a_n2570_n2088# 1.06382f
C44 drain_right.n13 a_n2570_n2088# 0.610245f
C45 minus.n0 a_n2570_n2088# 0.04132f
C46 minus.n1 a_n2570_n2088# 0.009376f
C47 minus.t2 a_n2570_n2088# 0.503368f
C48 minus.n2 a_n2570_n2088# 0.04132f
C49 minus.n3 a_n2570_n2088# 0.009376f
C50 minus.t4 a_n2570_n2088# 0.503368f
C51 minus.n4 a_n2570_n2088# 0.04132f
C52 minus.n5 a_n2570_n2088# 0.009376f
C53 minus.t6 a_n2570_n2088# 0.503368f
C54 minus.t9 a_n2570_n2088# 0.523132f
C55 minus.t0 a_n2570_n2088# 0.503368f
C56 minus.n6 a_n2570_n2088# 0.238262f
C57 minus.n7 a_n2570_n2088# 0.216275f
C58 minus.n8 a_n2570_n2088# 0.174854f
C59 minus.n9 a_n2570_n2088# 0.04132f
C60 minus.n10 a_n2570_n2088# 0.232601f
C61 minus.n11 a_n2570_n2088# 0.009376f
C62 minus.t14 a_n2570_n2088# 0.503368f
C63 minus.n12 a_n2570_n2088# 0.232601f
C64 minus.n13 a_n2570_n2088# 0.04132f
C65 minus.n14 a_n2570_n2088# 0.04132f
C66 minus.n15 a_n2570_n2088# 0.04132f
C67 minus.n16 a_n2570_n2088# 0.232601f
C68 minus.n17 a_n2570_n2088# 0.009376f
C69 minus.t15 a_n2570_n2088# 0.503368f
C70 minus.n18 a_n2570_n2088# 0.232601f
C71 minus.n19 a_n2570_n2088# 0.04132f
C72 minus.n20 a_n2570_n2088# 0.04132f
C73 minus.n21 a_n2570_n2088# 0.04132f
C74 minus.n22 a_n2570_n2088# 0.232601f
C75 minus.n23 a_n2570_n2088# 0.009376f
C76 minus.t13 a_n2570_n2088# 0.503368f
C77 minus.n24 a_n2570_n2088# 0.231455f
C78 minus.n25 a_n2570_n2088# 1.35689f
C79 minus.n26 a_n2570_n2088# 0.04132f
C80 minus.n27 a_n2570_n2088# 0.009376f
C81 minus.n28 a_n2570_n2088# 0.04132f
C82 minus.n29 a_n2570_n2088# 0.009376f
C83 minus.n30 a_n2570_n2088# 0.04132f
C84 minus.n31 a_n2570_n2088# 0.009376f
C85 minus.t11 a_n2570_n2088# 0.523132f
C86 minus.t12 a_n2570_n2088# 0.503368f
C87 minus.n32 a_n2570_n2088# 0.238262f
C88 minus.n33 a_n2570_n2088# 0.216275f
C89 minus.n34 a_n2570_n2088# 0.174854f
C90 minus.n35 a_n2570_n2088# 0.04132f
C91 minus.t7 a_n2570_n2088# 0.503368f
C92 minus.n36 a_n2570_n2088# 0.232601f
C93 minus.n37 a_n2570_n2088# 0.009376f
C94 minus.t8 a_n2570_n2088# 0.503368f
C95 minus.n38 a_n2570_n2088# 0.232601f
C96 minus.n39 a_n2570_n2088# 0.04132f
C97 minus.n40 a_n2570_n2088# 0.04132f
C98 minus.n41 a_n2570_n2088# 0.04132f
C99 minus.t10 a_n2570_n2088# 0.503368f
C100 minus.n42 a_n2570_n2088# 0.232601f
C101 minus.n43 a_n2570_n2088# 0.009376f
C102 minus.t3 a_n2570_n2088# 0.503368f
C103 minus.n44 a_n2570_n2088# 0.232601f
C104 minus.n45 a_n2570_n2088# 0.04132f
C105 minus.n46 a_n2570_n2088# 0.04132f
C106 minus.n47 a_n2570_n2088# 0.04132f
C107 minus.t5 a_n2570_n2088# 0.503368f
C108 minus.n48 a_n2570_n2088# 0.232601f
C109 minus.n49 a_n2570_n2088# 0.009376f
C110 minus.t1 a_n2570_n2088# 0.503368f
C111 minus.n50 a_n2570_n2088# 0.231455f
C112 minus.n51 a_n2570_n2088# 0.285193f
C113 minus.n52 a_n2570_n2088# 1.65076f
C114 source.n0 a_n2570_n2088# 0.0353f
C115 source.n1 a_n2570_n2088# 0.025114f
C116 source.n2 a_n2570_n2088# 0.013495f
C117 source.n3 a_n2570_n2088# 0.031898f
C118 source.n4 a_n2570_n2088# 0.014289f
C119 source.n5 a_n2570_n2088# 0.025114f
C120 source.n6 a_n2570_n2088# 0.013495f
C121 source.n7 a_n2570_n2088# 0.031898f
C122 source.n8 a_n2570_n2088# 0.014289f
C123 source.n9 a_n2570_n2088# 0.107472f
C124 source.t23 a_n2570_n2088# 0.05199f
C125 source.n10 a_n2570_n2088# 0.023923f
C126 source.n11 a_n2570_n2088# 0.018842f
C127 source.n12 a_n2570_n2088# 0.013495f
C128 source.n13 a_n2570_n2088# 0.59757f
C129 source.n14 a_n2570_n2088# 0.025114f
C130 source.n15 a_n2570_n2088# 0.013495f
C131 source.n16 a_n2570_n2088# 0.014289f
C132 source.n17 a_n2570_n2088# 0.031898f
C133 source.n18 a_n2570_n2088# 0.031898f
C134 source.n19 a_n2570_n2088# 0.014289f
C135 source.n20 a_n2570_n2088# 0.013495f
C136 source.n21 a_n2570_n2088# 0.025114f
C137 source.n22 a_n2570_n2088# 0.025114f
C138 source.n23 a_n2570_n2088# 0.013495f
C139 source.n24 a_n2570_n2088# 0.014289f
C140 source.n25 a_n2570_n2088# 0.031898f
C141 source.n26 a_n2570_n2088# 0.069054f
C142 source.n27 a_n2570_n2088# 0.014289f
C143 source.n28 a_n2570_n2088# 0.013495f
C144 source.n29 a_n2570_n2088# 0.05805f
C145 source.n30 a_n2570_n2088# 0.038638f
C146 source.n31 a_n2570_n2088# 0.656075f
C147 source.t19 a_n2570_n2088# 0.119076f
C148 source.t31 a_n2570_n2088# 0.119076f
C149 source.n32 a_n2570_n2088# 0.927377f
C150 source.n33 a_n2570_n2088# 0.379132f
C151 source.t20 a_n2570_n2088# 0.119076f
C152 source.t27 a_n2570_n2088# 0.119076f
C153 source.n34 a_n2570_n2088# 0.927377f
C154 source.n35 a_n2570_n2088# 0.379132f
C155 source.t18 a_n2570_n2088# 0.119076f
C156 source.t29 a_n2570_n2088# 0.119076f
C157 source.n36 a_n2570_n2088# 0.927377f
C158 source.n37 a_n2570_n2088# 0.379132f
C159 source.n38 a_n2570_n2088# 0.0353f
C160 source.n39 a_n2570_n2088# 0.025114f
C161 source.n40 a_n2570_n2088# 0.013495f
C162 source.n41 a_n2570_n2088# 0.031898f
C163 source.n42 a_n2570_n2088# 0.014289f
C164 source.n43 a_n2570_n2088# 0.025114f
C165 source.n44 a_n2570_n2088# 0.013495f
C166 source.n45 a_n2570_n2088# 0.031898f
C167 source.n46 a_n2570_n2088# 0.014289f
C168 source.n47 a_n2570_n2088# 0.107472f
C169 source.t26 a_n2570_n2088# 0.05199f
C170 source.n48 a_n2570_n2088# 0.023923f
C171 source.n49 a_n2570_n2088# 0.018842f
C172 source.n50 a_n2570_n2088# 0.013495f
C173 source.n51 a_n2570_n2088# 0.59757f
C174 source.n52 a_n2570_n2088# 0.025114f
C175 source.n53 a_n2570_n2088# 0.013495f
C176 source.n54 a_n2570_n2088# 0.014289f
C177 source.n55 a_n2570_n2088# 0.031898f
C178 source.n56 a_n2570_n2088# 0.031898f
C179 source.n57 a_n2570_n2088# 0.014289f
C180 source.n58 a_n2570_n2088# 0.013495f
C181 source.n59 a_n2570_n2088# 0.025114f
C182 source.n60 a_n2570_n2088# 0.025114f
C183 source.n61 a_n2570_n2088# 0.013495f
C184 source.n62 a_n2570_n2088# 0.014289f
C185 source.n63 a_n2570_n2088# 0.031898f
C186 source.n64 a_n2570_n2088# 0.069054f
C187 source.n65 a_n2570_n2088# 0.014289f
C188 source.n66 a_n2570_n2088# 0.013495f
C189 source.n67 a_n2570_n2088# 0.05805f
C190 source.n68 a_n2570_n2088# 0.038638f
C191 source.n69 a_n2570_n2088# 0.131324f
C192 source.n70 a_n2570_n2088# 0.0353f
C193 source.n71 a_n2570_n2088# 0.025114f
C194 source.n72 a_n2570_n2088# 0.013495f
C195 source.n73 a_n2570_n2088# 0.031898f
C196 source.n74 a_n2570_n2088# 0.014289f
C197 source.n75 a_n2570_n2088# 0.025114f
C198 source.n76 a_n2570_n2088# 0.013495f
C199 source.n77 a_n2570_n2088# 0.031898f
C200 source.n78 a_n2570_n2088# 0.014289f
C201 source.n79 a_n2570_n2088# 0.107472f
C202 source.t7 a_n2570_n2088# 0.05199f
C203 source.n80 a_n2570_n2088# 0.023923f
C204 source.n81 a_n2570_n2088# 0.018842f
C205 source.n82 a_n2570_n2088# 0.013495f
C206 source.n83 a_n2570_n2088# 0.59757f
C207 source.n84 a_n2570_n2088# 0.025114f
C208 source.n85 a_n2570_n2088# 0.013495f
C209 source.n86 a_n2570_n2088# 0.014289f
C210 source.n87 a_n2570_n2088# 0.031898f
C211 source.n88 a_n2570_n2088# 0.031898f
C212 source.n89 a_n2570_n2088# 0.014289f
C213 source.n90 a_n2570_n2088# 0.013495f
C214 source.n91 a_n2570_n2088# 0.025114f
C215 source.n92 a_n2570_n2088# 0.025114f
C216 source.n93 a_n2570_n2088# 0.013495f
C217 source.n94 a_n2570_n2088# 0.014289f
C218 source.n95 a_n2570_n2088# 0.031898f
C219 source.n96 a_n2570_n2088# 0.069054f
C220 source.n97 a_n2570_n2088# 0.014289f
C221 source.n98 a_n2570_n2088# 0.013495f
C222 source.n99 a_n2570_n2088# 0.05805f
C223 source.n100 a_n2570_n2088# 0.038638f
C224 source.n101 a_n2570_n2088# 0.131324f
C225 source.t10 a_n2570_n2088# 0.119076f
C226 source.t8 a_n2570_n2088# 0.119076f
C227 source.n102 a_n2570_n2088# 0.927377f
C228 source.n103 a_n2570_n2088# 0.379132f
C229 source.t6 a_n2570_n2088# 0.119076f
C230 source.t13 a_n2570_n2088# 0.119076f
C231 source.n104 a_n2570_n2088# 0.927377f
C232 source.n105 a_n2570_n2088# 0.379132f
C233 source.t11 a_n2570_n2088# 0.119076f
C234 source.t15 a_n2570_n2088# 0.119076f
C235 source.n106 a_n2570_n2088# 0.927377f
C236 source.n107 a_n2570_n2088# 0.379132f
C237 source.n108 a_n2570_n2088# 0.0353f
C238 source.n109 a_n2570_n2088# 0.025114f
C239 source.n110 a_n2570_n2088# 0.013495f
C240 source.n111 a_n2570_n2088# 0.031898f
C241 source.n112 a_n2570_n2088# 0.014289f
C242 source.n113 a_n2570_n2088# 0.025114f
C243 source.n114 a_n2570_n2088# 0.013495f
C244 source.n115 a_n2570_n2088# 0.031898f
C245 source.n116 a_n2570_n2088# 0.014289f
C246 source.n117 a_n2570_n2088# 0.107472f
C247 source.t14 a_n2570_n2088# 0.05199f
C248 source.n118 a_n2570_n2088# 0.023923f
C249 source.n119 a_n2570_n2088# 0.018842f
C250 source.n120 a_n2570_n2088# 0.013495f
C251 source.n121 a_n2570_n2088# 0.59757f
C252 source.n122 a_n2570_n2088# 0.025114f
C253 source.n123 a_n2570_n2088# 0.013495f
C254 source.n124 a_n2570_n2088# 0.014289f
C255 source.n125 a_n2570_n2088# 0.031898f
C256 source.n126 a_n2570_n2088# 0.031898f
C257 source.n127 a_n2570_n2088# 0.014289f
C258 source.n128 a_n2570_n2088# 0.013495f
C259 source.n129 a_n2570_n2088# 0.025114f
C260 source.n130 a_n2570_n2088# 0.025114f
C261 source.n131 a_n2570_n2088# 0.013495f
C262 source.n132 a_n2570_n2088# 0.014289f
C263 source.n133 a_n2570_n2088# 0.031898f
C264 source.n134 a_n2570_n2088# 0.069054f
C265 source.n135 a_n2570_n2088# 0.014289f
C266 source.n136 a_n2570_n2088# 0.013495f
C267 source.n137 a_n2570_n2088# 0.05805f
C268 source.n138 a_n2570_n2088# 0.038638f
C269 source.n139 a_n2570_n2088# 0.987448f
C270 source.n140 a_n2570_n2088# 0.0353f
C271 source.n141 a_n2570_n2088# 0.025114f
C272 source.n142 a_n2570_n2088# 0.013495f
C273 source.n143 a_n2570_n2088# 0.031898f
C274 source.n144 a_n2570_n2088# 0.014289f
C275 source.n145 a_n2570_n2088# 0.025114f
C276 source.n146 a_n2570_n2088# 0.013495f
C277 source.n147 a_n2570_n2088# 0.031898f
C278 source.n148 a_n2570_n2088# 0.014289f
C279 source.n149 a_n2570_n2088# 0.107472f
C280 source.t24 a_n2570_n2088# 0.05199f
C281 source.n150 a_n2570_n2088# 0.023923f
C282 source.n151 a_n2570_n2088# 0.018842f
C283 source.n152 a_n2570_n2088# 0.013495f
C284 source.n153 a_n2570_n2088# 0.59757f
C285 source.n154 a_n2570_n2088# 0.025114f
C286 source.n155 a_n2570_n2088# 0.013495f
C287 source.n156 a_n2570_n2088# 0.014289f
C288 source.n157 a_n2570_n2088# 0.031898f
C289 source.n158 a_n2570_n2088# 0.031898f
C290 source.n159 a_n2570_n2088# 0.014289f
C291 source.n160 a_n2570_n2088# 0.013495f
C292 source.n161 a_n2570_n2088# 0.025114f
C293 source.n162 a_n2570_n2088# 0.025114f
C294 source.n163 a_n2570_n2088# 0.013495f
C295 source.n164 a_n2570_n2088# 0.014289f
C296 source.n165 a_n2570_n2088# 0.031898f
C297 source.n166 a_n2570_n2088# 0.069054f
C298 source.n167 a_n2570_n2088# 0.014289f
C299 source.n168 a_n2570_n2088# 0.013495f
C300 source.n169 a_n2570_n2088# 0.05805f
C301 source.n170 a_n2570_n2088# 0.038638f
C302 source.n171 a_n2570_n2088# 0.987448f
C303 source.t16 a_n2570_n2088# 0.119076f
C304 source.t17 a_n2570_n2088# 0.119076f
C305 source.n172 a_n2570_n2088# 0.927371f
C306 source.n173 a_n2570_n2088# 0.379138f
C307 source.t28 a_n2570_n2088# 0.119076f
C308 source.t30 a_n2570_n2088# 0.119076f
C309 source.n174 a_n2570_n2088# 0.927371f
C310 source.n175 a_n2570_n2088# 0.379138f
C311 source.t25 a_n2570_n2088# 0.119076f
C312 source.t21 a_n2570_n2088# 0.119076f
C313 source.n176 a_n2570_n2088# 0.927371f
C314 source.n177 a_n2570_n2088# 0.379138f
C315 source.n178 a_n2570_n2088# 0.0353f
C316 source.n179 a_n2570_n2088# 0.025114f
C317 source.n180 a_n2570_n2088# 0.013495f
C318 source.n181 a_n2570_n2088# 0.031898f
C319 source.n182 a_n2570_n2088# 0.014289f
C320 source.n183 a_n2570_n2088# 0.025114f
C321 source.n184 a_n2570_n2088# 0.013495f
C322 source.n185 a_n2570_n2088# 0.031898f
C323 source.n186 a_n2570_n2088# 0.014289f
C324 source.n187 a_n2570_n2088# 0.107472f
C325 source.t22 a_n2570_n2088# 0.05199f
C326 source.n188 a_n2570_n2088# 0.023923f
C327 source.n189 a_n2570_n2088# 0.018842f
C328 source.n190 a_n2570_n2088# 0.013495f
C329 source.n191 a_n2570_n2088# 0.59757f
C330 source.n192 a_n2570_n2088# 0.025114f
C331 source.n193 a_n2570_n2088# 0.013495f
C332 source.n194 a_n2570_n2088# 0.014289f
C333 source.n195 a_n2570_n2088# 0.031898f
C334 source.n196 a_n2570_n2088# 0.031898f
C335 source.n197 a_n2570_n2088# 0.014289f
C336 source.n198 a_n2570_n2088# 0.013495f
C337 source.n199 a_n2570_n2088# 0.025114f
C338 source.n200 a_n2570_n2088# 0.025114f
C339 source.n201 a_n2570_n2088# 0.013495f
C340 source.n202 a_n2570_n2088# 0.014289f
C341 source.n203 a_n2570_n2088# 0.031898f
C342 source.n204 a_n2570_n2088# 0.069054f
C343 source.n205 a_n2570_n2088# 0.014289f
C344 source.n206 a_n2570_n2088# 0.013495f
C345 source.n207 a_n2570_n2088# 0.05805f
C346 source.n208 a_n2570_n2088# 0.038638f
C347 source.n209 a_n2570_n2088# 0.131324f
C348 source.n210 a_n2570_n2088# 0.0353f
C349 source.n211 a_n2570_n2088# 0.025114f
C350 source.n212 a_n2570_n2088# 0.013495f
C351 source.n213 a_n2570_n2088# 0.031898f
C352 source.n214 a_n2570_n2088# 0.014289f
C353 source.n215 a_n2570_n2088# 0.025114f
C354 source.n216 a_n2570_n2088# 0.013495f
C355 source.n217 a_n2570_n2088# 0.031898f
C356 source.n218 a_n2570_n2088# 0.014289f
C357 source.n219 a_n2570_n2088# 0.107472f
C358 source.t1 a_n2570_n2088# 0.05199f
C359 source.n220 a_n2570_n2088# 0.023923f
C360 source.n221 a_n2570_n2088# 0.018842f
C361 source.n222 a_n2570_n2088# 0.013495f
C362 source.n223 a_n2570_n2088# 0.59757f
C363 source.n224 a_n2570_n2088# 0.025114f
C364 source.n225 a_n2570_n2088# 0.013495f
C365 source.n226 a_n2570_n2088# 0.014289f
C366 source.n227 a_n2570_n2088# 0.031898f
C367 source.n228 a_n2570_n2088# 0.031898f
C368 source.n229 a_n2570_n2088# 0.014289f
C369 source.n230 a_n2570_n2088# 0.013495f
C370 source.n231 a_n2570_n2088# 0.025114f
C371 source.n232 a_n2570_n2088# 0.025114f
C372 source.n233 a_n2570_n2088# 0.013495f
C373 source.n234 a_n2570_n2088# 0.014289f
C374 source.n235 a_n2570_n2088# 0.031898f
C375 source.n236 a_n2570_n2088# 0.069054f
C376 source.n237 a_n2570_n2088# 0.014289f
C377 source.n238 a_n2570_n2088# 0.013495f
C378 source.n239 a_n2570_n2088# 0.05805f
C379 source.n240 a_n2570_n2088# 0.038638f
C380 source.n241 a_n2570_n2088# 0.131324f
C381 source.t5 a_n2570_n2088# 0.119076f
C382 source.t12 a_n2570_n2088# 0.119076f
C383 source.n242 a_n2570_n2088# 0.927371f
C384 source.n243 a_n2570_n2088# 0.379138f
C385 source.t4 a_n2570_n2088# 0.119076f
C386 source.t9 a_n2570_n2088# 0.119076f
C387 source.n244 a_n2570_n2088# 0.927371f
C388 source.n245 a_n2570_n2088# 0.379138f
C389 source.t2 a_n2570_n2088# 0.119076f
C390 source.t3 a_n2570_n2088# 0.119076f
C391 source.n246 a_n2570_n2088# 0.927371f
C392 source.n247 a_n2570_n2088# 0.379138f
C393 source.n248 a_n2570_n2088# 0.0353f
C394 source.n249 a_n2570_n2088# 0.025114f
C395 source.n250 a_n2570_n2088# 0.013495f
C396 source.n251 a_n2570_n2088# 0.031898f
C397 source.n252 a_n2570_n2088# 0.014289f
C398 source.n253 a_n2570_n2088# 0.025114f
C399 source.n254 a_n2570_n2088# 0.013495f
C400 source.n255 a_n2570_n2088# 0.031898f
C401 source.n256 a_n2570_n2088# 0.014289f
C402 source.n257 a_n2570_n2088# 0.107472f
C403 source.t0 a_n2570_n2088# 0.05199f
C404 source.n258 a_n2570_n2088# 0.023923f
C405 source.n259 a_n2570_n2088# 0.018842f
C406 source.n260 a_n2570_n2088# 0.013495f
C407 source.n261 a_n2570_n2088# 0.59757f
C408 source.n262 a_n2570_n2088# 0.025114f
C409 source.n263 a_n2570_n2088# 0.013495f
C410 source.n264 a_n2570_n2088# 0.014289f
C411 source.n265 a_n2570_n2088# 0.031898f
C412 source.n266 a_n2570_n2088# 0.031898f
C413 source.n267 a_n2570_n2088# 0.014289f
C414 source.n268 a_n2570_n2088# 0.013495f
C415 source.n269 a_n2570_n2088# 0.025114f
C416 source.n270 a_n2570_n2088# 0.025114f
C417 source.n271 a_n2570_n2088# 0.013495f
C418 source.n272 a_n2570_n2088# 0.014289f
C419 source.n273 a_n2570_n2088# 0.031898f
C420 source.n274 a_n2570_n2088# 0.069054f
C421 source.n275 a_n2570_n2088# 0.014289f
C422 source.n276 a_n2570_n2088# 0.013495f
C423 source.n277 a_n2570_n2088# 0.05805f
C424 source.n278 a_n2570_n2088# 0.038638f
C425 source.n279 a_n2570_n2088# 0.295146f
C426 source.n280 a_n2570_n2088# 1.04154f
C427 drain_left.t6 a_n2570_n2088# 0.129008f
C428 drain_left.t15 a_n2570_n2088# 0.129008f
C429 drain_left.n0 a_n2570_n2088# 1.08098f
C430 drain_left.t1 a_n2570_n2088# 0.129008f
C431 drain_left.t13 a_n2570_n2088# 0.129008f
C432 drain_left.n1 a_n2570_n2088# 1.07593f
C433 drain_left.n2 a_n2570_n2088# 0.716818f
C434 drain_left.t7 a_n2570_n2088# 0.129008f
C435 drain_left.t11 a_n2570_n2088# 0.129008f
C436 drain_left.n3 a_n2570_n2088# 1.08098f
C437 drain_left.t3 a_n2570_n2088# 0.129008f
C438 drain_left.t9 a_n2570_n2088# 0.129008f
C439 drain_left.n4 a_n2570_n2088# 1.07593f
C440 drain_left.n5 a_n2570_n2088# 0.716818f
C441 drain_left.n6 a_n2570_n2088# 1.20428f
C442 drain_left.t4 a_n2570_n2088# 0.129008f
C443 drain_left.t0 a_n2570_n2088# 0.129008f
C444 drain_left.n7 a_n2570_n2088# 1.08099f
C445 drain_left.t8 a_n2570_n2088# 0.129008f
C446 drain_left.t5 a_n2570_n2088# 0.129008f
C447 drain_left.n8 a_n2570_n2088# 1.07593f
C448 drain_left.n9 a_n2570_n2088# 0.758961f
C449 drain_left.t10 a_n2570_n2088# 0.129008f
C450 drain_left.t14 a_n2570_n2088# 0.129008f
C451 drain_left.n10 a_n2570_n2088# 1.07593f
C452 drain_left.n11 a_n2570_n2088# 0.376528f
C453 drain_left.t12 a_n2570_n2088# 0.129008f
C454 drain_left.t2 a_n2570_n2088# 0.129008f
C455 drain_left.n12 a_n2570_n2088# 1.07593f
C456 drain_left.n13 a_n2570_n2088# 0.617198f
C457 plus.n0 a_n2570_n2088# 0.042291f
C458 plus.t8 a_n2570_n2088# 0.515201f
C459 plus.t0 a_n2570_n2088# 0.515201f
C460 plus.n1 a_n2570_n2088# 0.042291f
C461 plus.t12 a_n2570_n2088# 0.515201f
C462 plus.n2 a_n2570_n2088# 0.238069f
C463 plus.n3 a_n2570_n2088# 0.042291f
C464 plus.t4 a_n2570_n2088# 0.515201f
C465 plus.t11 a_n2570_n2088# 0.515201f
C466 plus.n4 a_n2570_n2088# 0.238069f
C467 plus.n5 a_n2570_n2088# 0.042291f
C468 plus.t2 a_n2570_n2088# 0.515201f
C469 plus.t13 a_n2570_n2088# 0.515201f
C470 plus.n6 a_n2570_n2088# 0.243863f
C471 plus.t5 a_n2570_n2088# 0.53543f
C472 plus.n7 a_n2570_n2088# 0.221359f
C473 plus.n8 a_n2570_n2088# 0.178965f
C474 plus.n9 a_n2570_n2088# 0.009597f
C475 plus.n10 a_n2570_n2088# 0.238069f
C476 plus.n11 a_n2570_n2088# 0.009597f
C477 plus.n12 a_n2570_n2088# 0.042291f
C478 plus.n13 a_n2570_n2088# 0.042291f
C479 plus.n14 a_n2570_n2088# 0.042291f
C480 plus.n15 a_n2570_n2088# 0.009597f
C481 plus.n16 a_n2570_n2088# 0.238069f
C482 plus.n17 a_n2570_n2088# 0.009597f
C483 plus.n18 a_n2570_n2088# 0.042291f
C484 plus.n19 a_n2570_n2088# 0.042291f
C485 plus.n20 a_n2570_n2088# 0.042291f
C486 plus.n21 a_n2570_n2088# 0.009597f
C487 plus.n22 a_n2570_n2088# 0.238069f
C488 plus.n23 a_n2570_n2088# 0.009597f
C489 plus.n24 a_n2570_n2088# 0.236896f
C490 plus.n25 a_n2570_n2088# 0.378494f
C491 plus.n26 a_n2570_n2088# 0.042291f
C492 plus.t7 a_n2570_n2088# 0.515201f
C493 plus.n27 a_n2570_n2088# 0.042291f
C494 plus.t15 a_n2570_n2088# 0.515201f
C495 plus.t14 a_n2570_n2088# 0.515201f
C496 plus.n28 a_n2570_n2088# 0.238069f
C497 plus.n29 a_n2570_n2088# 0.042291f
C498 plus.t3 a_n2570_n2088# 0.515201f
C499 plus.t1 a_n2570_n2088# 0.515201f
C500 plus.n30 a_n2570_n2088# 0.238069f
C501 plus.n31 a_n2570_n2088# 0.042291f
C502 plus.t6 a_n2570_n2088# 0.515201f
C503 plus.t10 a_n2570_n2088# 0.515201f
C504 plus.n32 a_n2570_n2088# 0.243863f
C505 plus.t9 a_n2570_n2088# 0.53543f
C506 plus.n33 a_n2570_n2088# 0.221359f
C507 plus.n34 a_n2570_n2088# 0.178965f
C508 plus.n35 a_n2570_n2088# 0.009597f
C509 plus.n36 a_n2570_n2088# 0.238069f
C510 plus.n37 a_n2570_n2088# 0.009597f
C511 plus.n38 a_n2570_n2088# 0.042291f
C512 plus.n39 a_n2570_n2088# 0.042291f
C513 plus.n40 a_n2570_n2088# 0.042291f
C514 plus.n41 a_n2570_n2088# 0.009597f
C515 plus.n42 a_n2570_n2088# 0.238069f
C516 plus.n43 a_n2570_n2088# 0.009597f
C517 plus.n44 a_n2570_n2088# 0.042291f
C518 plus.n45 a_n2570_n2088# 0.042291f
C519 plus.n46 a_n2570_n2088# 0.042291f
C520 plus.n47 a_n2570_n2088# 0.009597f
C521 plus.n48 a_n2570_n2088# 0.238069f
C522 plus.n49 a_n2570_n2088# 0.009597f
C523 plus.n50 a_n2570_n2088# 0.236896f
C524 plus.n51 a_n2570_n2088# 1.25761f
.ends

