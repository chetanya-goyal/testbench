* NGSPICE file created from diffpair571.ext - technology: sky130A

.subckt diffpair571 minus drain_right drain_left source plus
X0 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X1 drain_right.t3 minus.t0 source.t5 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X2 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X3 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X4 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X5 drain_left.t3 plus.t0 source.t3 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X6 source.t2 plus.t1 drain_left.t2 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X7 drain_left.t1 plus.t2 source.t1 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X8 source.t6 minus.t1 drain_right.t2 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X9 source.t4 minus.t2 drain_right.t1 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X10 drain_right.t0 minus.t3 source.t7 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X11 source.t0 plus.t3 drain_left.t0 a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
R0 minus.n0 minus.t2 2605.36
R1 minus.n0 minus.t0 2605.36
R2 minus.n1 minus.t3 2605.36
R3 minus.n1 minus.t1 2605.36
R4 minus.n2 minus.n0 200.345
R5 minus.n2 minus.n1 167.732
R6 minus minus.n2 0.188
R7 source.n0 source.t1 44.1297
R8 source.n1 source.t0 44.1296
R9 source.n2 source.t5 44.1296
R10 source.n3 source.t4 44.1296
R11 source.n7 source.t7 44.1295
R12 source.n6 source.t6 44.1295
R13 source.n5 source.t3 44.1295
R14 source.n4 source.t2 44.1295
R15 source.n4 source.n3 27.8204
R16 source.n8 source.n0 22.329
R17 source.n8 source.n7 5.49188
R18 source.n2 source.n1 0.470328
R19 source.n6 source.n5 0.470328
R20 source.n3 source.n2 0.457397
R21 source.n1 source.n0 0.457397
R22 source.n5 source.n4 0.457397
R23 source.n7 source.n6 0.457397
R24 source source.n8 0.188
R25 drain_right drain_right.n0 93.6213
R26 drain_right drain_right.n1 65.9281
R27 drain_right.n0 drain_right.t2 0.9905
R28 drain_right.n0 drain_right.t0 0.9905
R29 drain_right.n1 drain_right.t1 0.9905
R30 drain_right.n1 drain_right.t3 0.9905
R31 plus.n0 plus.t3 2605.36
R32 plus.n0 plus.t2 2605.36
R33 plus.n1 plus.t0 2605.36
R34 plus.n1 plus.t1 2605.36
R35 plus plus.n1 191.196
R36 plus plus.n0 176.406
R37 drain_left drain_left.n0 94.1745
R38 drain_left drain_left.n1 65.9281
R39 drain_left.n0 drain_left.t2 0.9905
R40 drain_left.n0 drain_left.t3 0.9905
R41 drain_left.n1 drain_left.t0 0.9905
R42 drain_left.n1 drain_left.t1 0.9905
C0 drain_left drain_right 0.457115f
C1 drain_left source 17.6864f
C2 drain_left minus 0.171239f
C3 source drain_right 17.6844f
C4 minus drain_right 2.69903f
C5 source minus 1.74355f
C6 plus drain_left 2.79374f
C7 plus drain_right 0.248706f
C8 plus source 1.75758f
C9 plus minus 5.92147f
C10 drain_right a_n1034_n4892# 9.55099f
C11 drain_left a_n1034_n4892# 9.745669f
C12 source a_n1034_n4892# 12.228801f
C13 minus a_n1034_n4892# 4.490845f
C14 plus a_n1034_n4892# 9.17296f
C15 drain_left.t2 a_n1034_n4892# 0.579914f
C16 drain_left.t3 a_n1034_n4892# 0.579914f
C17 drain_left.n0 a_n1034_n4892# 6.17853f
C18 drain_left.t0 a_n1034_n4892# 0.579914f
C19 drain_left.t1 a_n1034_n4892# 0.579914f
C20 drain_left.n1 a_n1034_n4892# 5.3696f
C21 plus.t3 a_n1034_n4892# 0.633371f
C22 plus.t2 a_n1034_n4892# 0.633371f
C23 plus.n0 a_n1034_n4892# 0.562126f
C24 plus.t1 a_n1034_n4892# 0.633371f
C25 plus.t0 a_n1034_n4892# 0.633371f
C26 plus.n1 a_n1034_n4892# 0.761785f
C27 drain_right.t2 a_n1034_n4892# 0.581154f
C28 drain_right.t0 a_n1034_n4892# 0.581154f
C29 drain_right.n0 a_n1034_n4892# 6.15471f
C30 drain_right.t1 a_n1034_n4892# 0.581154f
C31 drain_right.t3 a_n1034_n4892# 0.581154f
C32 drain_right.n1 a_n1034_n4892# 5.38109f
C33 source.t1 a_n1034_n4892# 3.37998f
C34 source.n0 a_n1034_n4892# 1.43054f
C35 source.t0 a_n1034_n4892# 3.37998f
C36 source.n1 a_n1034_n4892# 0.318809f
C37 source.t5 a_n1034_n4892# 3.37998f
C38 source.n2 a_n1034_n4892# 0.318809f
C39 source.t4 a_n1034_n4892# 3.37998f
C40 source.n3 a_n1034_n4892# 1.76002f
C41 source.t2 a_n1034_n4892# 3.37996f
C42 source.n4 a_n1034_n4892# 1.76004f
C43 source.t3 a_n1034_n4892# 3.37996f
C44 source.n5 a_n1034_n4892# 0.318828f
C45 source.t6 a_n1034_n4892# 3.37996f
C46 source.n6 a_n1034_n4892# 0.318828f
C47 source.t7 a_n1034_n4892# 3.37996f
C48 source.n7 a_n1034_n4892# 0.420296f
C49 source.n8 a_n1034_n4892# 1.68255f
C50 minus.t2 a_n1034_n4892# 0.618059f
C51 minus.t0 a_n1034_n4892# 0.618059f
C52 minus.n0 a_n1034_n4892# 0.900872f
C53 minus.t1 a_n1034_n4892# 0.618059f
C54 minus.t3 a_n1034_n4892# 0.618059f
C55 minus.n1 a_n1034_n4892# 0.491306f
C56 minus.n2 a_n1034_n4892# 4.69976f
.ends

