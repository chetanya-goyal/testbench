* NGSPICE file created from diffpair615.ext - technology: sky130A

.subckt diffpair615 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t18 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X1 drain_left.t11 plus.t0 source.t4 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X2 source.t22 plus.t1 drain_left.t10 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X3 drain_left.t9 plus.t2 source.t6 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X4 drain_right.t10 minus.t1 source.t16 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X5 drain_right.t9 minus.t2 source.t10 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X6 drain_left.t8 plus.t3 source.t0 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X7 source.t9 minus.t3 drain_right.t8 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X8 source.t13 minus.t4 drain_right.t7 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X9 drain_right.t6 minus.t5 source.t14 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X10 source.t23 plus.t4 drain_left.t7 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X11 source.t2 plus.t5 drain_left.t6 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X12 source.t15 minus.t6 drain_right.t5 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X13 source.t17 minus.t7 drain_right.t4 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X14 drain_right.t3 minus.t8 source.t8 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X15 source.t1 plus.t6 drain_left.t5 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X16 drain_left.t4 plus.t7 source.t20 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X17 source.t7 minus.t9 drain_right.t2 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X18 a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X19 source.t21 plus.t8 drain_left.t3 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X20 drain_right.t1 minus.t10 source.t12 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X21 a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X22 drain_left.t2 plus.t9 source.t19 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X23 source.t5 plus.t10 drain_left.t1 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X24 source.t11 minus.t11 drain_right.t0 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X25 a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X26 a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X27 drain_left.t0 plus.t11 source.t3 a_n2018_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
R0 minus.n2 minus.t10 893.865
R1 minus.n14 minus.t11 893.865
R2 minus.n3 minus.t9 868.806
R3 minus.n4 minus.t8 868.806
R4 minus.n1 minus.t6 868.806
R5 minus.n8 minus.t2 868.806
R6 minus.n10 minus.t3 868.806
R7 minus.n15 minus.t5 868.806
R8 minus.n16 minus.t7 868.806
R9 minus.n13 minus.t0 868.806
R10 minus.n20 minus.t4 868.806
R11 minus.n22 minus.t1 868.806
R12 minus.n11 minus.n10 161.3
R13 minus.n9 minus.n0 161.3
R14 minus.n8 minus.n7 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n6 minus.n1 80.6037
R19 minus.n5 minus.n4 80.6037
R20 minus.n18 minus.n13 80.6037
R21 minus.n17 minus.n16 80.6037
R22 minus.n4 minus.n3 48.2005
R23 minus.n4 minus.n1 48.2005
R24 minus.n8 minus.n1 48.2005
R25 minus.n16 minus.n15 48.2005
R26 minus.n16 minus.n13 48.2005
R27 minus.n20 minus.n13 48.2005
R28 minus.n5 minus.n2 45.0744
R29 minus.n17 minus.n14 45.0744
R30 minus.n24 minus.n11 42.9134
R31 minus.n10 minus.n9 40.1672
R32 minus.n22 minus.n21 40.1672
R33 minus.n3 minus.n2 16.1124
R34 minus.n15 minus.n14 16.1124
R35 minus.n9 minus.n8 8.03383
R36 minus.n21 minus.n20 8.03383
R37 minus.n24 minus.n23 6.58762
R38 minus.n6 minus.n5 0.380177
R39 minus.n18 minus.n17 0.380177
R40 minus.n7 minus.n6 0.285035
R41 minus.n19 minus.n18 0.285035
R42 minus.n11 minus.n0 0.189894
R43 minus.n7 minus.n0 0.189894
R44 minus.n19 minus.n12 0.189894
R45 minus.n23 minus.n12 0.189894
R46 minus minus.n24 0.188
R47 source.n0 source.t6 44.1297
R48 source.n5 source.t5 44.1296
R49 source.n6 source.t12 44.1296
R50 source.n11 source.t9 44.1296
R51 source.n23 source.t16 44.1295
R52 source.n18 source.t11 44.1295
R53 source.n17 source.t4 44.1295
R54 source.n12 source.t23 44.1295
R55 source.n2 source.n1 43.1397
R56 source.n4 source.n3 43.1397
R57 source.n8 source.n7 43.1397
R58 source.n10 source.n9 43.1397
R59 source.n22 source.n21 43.1396
R60 source.n20 source.n19 43.1396
R61 source.n16 source.n15 43.1396
R62 source.n14 source.n13 43.1396
R63 source.n12 source.n11 28.1501
R64 source.n24 source.n0 22.4863
R65 source.n24 source.n23 5.66429
R66 source.n21 source.t18 0.9905
R67 source.n21 source.t13 0.9905
R68 source.n19 source.t14 0.9905
R69 source.n19 source.t17 0.9905
R70 source.n15 source.t3 0.9905
R71 source.n15 source.t1 0.9905
R72 source.n13 source.t0 0.9905
R73 source.n13 source.t22 0.9905
R74 source.n1 source.t20 0.9905
R75 source.n1 source.t2 0.9905
R76 source.n3 source.t19 0.9905
R77 source.n3 source.t21 0.9905
R78 source.n7 source.t8 0.9905
R79 source.n7 source.t7 0.9905
R80 source.n9 source.t10 0.9905
R81 source.n9 source.t15 0.9905
R82 source.n11 source.n10 0.802224
R83 source.n10 source.n8 0.802224
R84 source.n8 source.n6 0.802224
R85 source.n5 source.n4 0.802224
R86 source.n4 source.n2 0.802224
R87 source.n2 source.n0 0.802224
R88 source.n14 source.n12 0.802224
R89 source.n16 source.n14 0.802224
R90 source.n17 source.n16 0.802224
R91 source.n20 source.n18 0.802224
R92 source.n22 source.n20 0.802224
R93 source.n23 source.n22 0.802224
R94 source.n6 source.n5 0.470328
R95 source.n18 source.n17 0.470328
R96 source source.n24 0.188
R97 drain_right.n6 drain_right.n4 60.6202
R98 drain_right.n3 drain_right.n2 60.5648
R99 drain_right.n3 drain_right.n0 60.5648
R100 drain_right.n6 drain_right.n5 59.8185
R101 drain_right.n8 drain_right.n7 59.8185
R102 drain_right.n3 drain_right.n1 59.8184
R103 drain_right drain_right.n3 36.8831
R104 drain_right drain_right.n8 6.45494
R105 drain_right.n1 drain_right.t4 0.9905
R106 drain_right.n1 drain_right.t11 0.9905
R107 drain_right.n2 drain_right.t7 0.9905
R108 drain_right.n2 drain_right.t10 0.9905
R109 drain_right.n0 drain_right.t0 0.9905
R110 drain_right.n0 drain_right.t6 0.9905
R111 drain_right.n4 drain_right.t2 0.9905
R112 drain_right.n4 drain_right.t1 0.9905
R113 drain_right.n5 drain_right.t5 0.9905
R114 drain_right.n5 drain_right.t3 0.9905
R115 drain_right.n7 drain_right.t8 0.9905
R116 drain_right.n7 drain_right.t9 0.9905
R117 drain_right.n8 drain_right.n6 0.802224
R118 plus.n4 plus.t10 893.865
R119 plus.n16 plus.t0 893.865
R120 plus.n10 plus.t2 868.806
R121 plus.n8 plus.t5 868.806
R122 plus.n7 plus.t7 868.806
R123 plus.n6 plus.t8 868.806
R124 plus.n5 plus.t9 868.806
R125 plus.n22 plus.t4 868.806
R126 plus.n20 plus.t3 868.806
R127 plus.n19 plus.t1 868.806
R128 plus.n18 plus.t11 868.806
R129 plus.n17 plus.t6 868.806
R130 plus.n8 plus.n1 161.3
R131 plus.n9 plus.n0 161.3
R132 plus.n11 plus.n10 161.3
R133 plus.n20 plus.n13 161.3
R134 plus.n21 plus.n12 161.3
R135 plus.n23 plus.n22 161.3
R136 plus.n6 plus.n3 80.6037
R137 plus.n7 plus.n2 80.6037
R138 plus.n18 plus.n15 80.6037
R139 plus.n19 plus.n14 80.6037
R140 plus.n8 plus.n7 48.2005
R141 plus.n7 plus.n6 48.2005
R142 plus.n6 plus.n5 48.2005
R143 plus.n20 plus.n19 48.2005
R144 plus.n19 plus.n18 48.2005
R145 plus.n18 plus.n17 48.2005
R146 plus.n4 plus.n3 45.0744
R147 plus.n16 plus.n15 45.0744
R148 plus.n10 plus.n9 40.1672
R149 plus.n22 plus.n21 40.1672
R150 plus plus.n23 33.7642
R151 plus.n5 plus.n4 16.1124
R152 plus.n17 plus.n16 16.1124
R153 plus plus.n11 15.2619
R154 plus.n9 plus.n8 8.03383
R155 plus.n21 plus.n20 8.03383
R156 plus.n3 plus.n2 0.380177
R157 plus.n15 plus.n14 0.380177
R158 plus.n2 plus.n1 0.285035
R159 plus.n14 plus.n13 0.285035
R160 plus.n1 plus.n0 0.189894
R161 plus.n11 plus.n0 0.189894
R162 plus.n23 plus.n12 0.189894
R163 plus.n13 plus.n12 0.189894
R164 drain_left.n6 drain_left.n4 60.6202
R165 drain_left.n3 drain_left.n2 60.5648
R166 drain_left.n3 drain_left.n0 60.5648
R167 drain_left.n8 drain_left.n7 59.8185
R168 drain_left.n6 drain_left.n5 59.8185
R169 drain_left.n3 drain_left.n1 59.8184
R170 drain_left drain_left.n3 37.4363
R171 drain_left drain_left.n8 6.45494
R172 drain_left.n1 drain_left.t10 0.9905
R173 drain_left.n1 drain_left.t0 0.9905
R174 drain_left.n2 drain_left.t5 0.9905
R175 drain_left.n2 drain_left.t11 0.9905
R176 drain_left.n0 drain_left.t7 0.9905
R177 drain_left.n0 drain_left.t8 0.9905
R178 drain_left.n7 drain_left.t6 0.9905
R179 drain_left.n7 drain_left.t9 0.9905
R180 drain_left.n5 drain_left.t3 0.9905
R181 drain_left.n5 drain_left.t4 0.9905
R182 drain_left.n4 drain_left.t1 0.9905
R183 drain_left.n4 drain_left.t2 0.9905
R184 drain_left.n8 drain_left.n6 0.802224
C0 plus drain_left 11.925f
C1 source plus 11.2725f
C2 minus drain_right 11.727799f
C3 source drain_left 26.0706f
C4 plus drain_right 0.352374f
C5 drain_left drain_right 1.01253f
C6 source drain_right 26.072199f
C7 minus plus 7.1455f
C8 minus drain_left 0.17204f
C9 minus source 11.2585f
C10 drain_right a_n2018_n4888# 7.643939f
C11 drain_left a_n2018_n4888# 7.93838f
C12 source a_n2018_n4888# 13.487007f
C13 minus a_n2018_n4888# 8.470071f
C14 plus a_n2018_n4888# 10.665021f
C15 drain_left.t7 a_n2018_n4888# 0.445533f
C16 drain_left.t8 a_n2018_n4888# 0.445533f
C17 drain_left.n0 a_n2018_n4888# 4.07797f
C18 drain_left.t10 a_n2018_n4888# 0.445533f
C19 drain_left.t0 a_n2018_n4888# 0.445533f
C20 drain_left.n1 a_n2018_n4888# 4.07316f
C21 drain_left.t5 a_n2018_n4888# 0.445533f
C22 drain_left.t11 a_n2018_n4888# 0.445533f
C23 drain_left.n2 a_n2018_n4888# 4.07797f
C24 drain_left.n3 a_n2018_n4888# 3.08939f
C25 drain_left.t1 a_n2018_n4888# 0.445533f
C26 drain_left.t2 a_n2018_n4888# 0.445533f
C27 drain_left.n4 a_n2018_n4888# 4.07838f
C28 drain_left.t3 a_n2018_n4888# 0.445533f
C29 drain_left.t4 a_n2018_n4888# 0.445533f
C30 drain_left.n5 a_n2018_n4888# 4.07315f
C31 drain_left.n6 a_n2018_n4888# 0.773208f
C32 drain_left.t6 a_n2018_n4888# 0.445533f
C33 drain_left.t9 a_n2018_n4888# 0.445533f
C34 drain_left.n7 a_n2018_n4888# 4.07315f
C35 drain_left.n8 a_n2018_n4888# 0.629353f
C36 plus.n0 a_n2018_n4888# 0.044159f
C37 plus.t2 a_n2018_n4888# 1.50063f
C38 plus.t5 a_n2018_n4888# 1.50063f
C39 plus.n1 a_n2018_n4888# 0.058924f
C40 plus.t7 a_n2018_n4888# 1.50063f
C41 plus.n2 a_n2018_n4888# 0.073552f
C42 plus.t8 a_n2018_n4888# 1.50063f
C43 plus.n3 a_n2018_n4888# 0.226319f
C44 plus.t9 a_n2018_n4888# 1.50063f
C45 plus.t10 a_n2018_n4888# 1.51636f
C46 plus.n4 a_n2018_n4888# 0.548871f
C47 plus.n5 a_n2018_n4888# 0.57012f
C48 plus.n6 a_n2018_n4888# 0.571732f
C49 plus.n7 a_n2018_n4888# 0.571732f
C50 plus.n8 a_n2018_n4888# 0.563209f
C51 plus.n9 a_n2018_n4888# 0.010021f
C52 plus.n10 a_n2018_n4888# 0.560215f
C53 plus.n11 a_n2018_n4888# 0.679404f
C54 plus.n12 a_n2018_n4888# 0.044159f
C55 plus.t4 a_n2018_n4888# 1.50063f
C56 plus.n13 a_n2018_n4888# 0.058924f
C57 plus.t3 a_n2018_n4888# 1.50063f
C58 plus.n14 a_n2018_n4888# 0.073552f
C59 plus.t1 a_n2018_n4888# 1.50063f
C60 plus.n15 a_n2018_n4888# 0.226319f
C61 plus.t11 a_n2018_n4888# 1.50063f
C62 plus.t0 a_n2018_n4888# 1.51636f
C63 plus.n16 a_n2018_n4888# 0.548871f
C64 plus.t6 a_n2018_n4888# 1.50063f
C65 plus.n17 a_n2018_n4888# 0.57012f
C66 plus.n18 a_n2018_n4888# 0.571732f
C67 plus.n19 a_n2018_n4888# 0.571732f
C68 plus.n20 a_n2018_n4888# 0.563209f
C69 plus.n21 a_n2018_n4888# 0.010021f
C70 plus.n22 a_n2018_n4888# 0.560215f
C71 plus.n23 a_n2018_n4888# 1.60415f
C72 drain_right.t0 a_n2018_n4888# 0.444478f
C73 drain_right.t6 a_n2018_n4888# 0.444478f
C74 drain_right.n0 a_n2018_n4888# 4.06832f
C75 drain_right.t4 a_n2018_n4888# 0.444478f
C76 drain_right.t11 a_n2018_n4888# 0.444478f
C77 drain_right.n1 a_n2018_n4888# 4.06351f
C78 drain_right.t7 a_n2018_n4888# 0.444478f
C79 drain_right.t10 a_n2018_n4888# 0.444478f
C80 drain_right.n2 a_n2018_n4888# 4.06832f
C81 drain_right.n3 a_n2018_n4888# 3.02367f
C82 drain_right.t2 a_n2018_n4888# 0.444478f
C83 drain_right.t1 a_n2018_n4888# 0.444478f
C84 drain_right.n4 a_n2018_n4888# 4.06872f
C85 drain_right.t5 a_n2018_n4888# 0.444478f
C86 drain_right.t3 a_n2018_n4888# 0.444478f
C87 drain_right.n5 a_n2018_n4888# 4.06351f
C88 drain_right.n6 a_n2018_n4888# 0.771377f
C89 drain_right.t8 a_n2018_n4888# 0.444478f
C90 drain_right.t9 a_n2018_n4888# 0.444478f
C91 drain_right.n7 a_n2018_n4888# 4.06351f
C92 drain_right.n8 a_n2018_n4888# 0.627863f
C93 source.t6 a_n2018_n4888# 3.9602f
C94 source.n0 a_n2018_n4888# 1.7132f
C95 source.t20 a_n2018_n4888# 0.346523f
C96 source.t2 a_n2018_n4888# 0.346523f
C97 source.n1 a_n2018_n4888# 3.09806f
C98 source.n2 a_n2018_n4888# 0.338426f
C99 source.t19 a_n2018_n4888# 0.346523f
C100 source.t21 a_n2018_n4888# 0.346523f
C101 source.n3 a_n2018_n4888# 3.09806f
C102 source.n4 a_n2018_n4888# 0.338426f
C103 source.t5 a_n2018_n4888# 3.96021f
C104 source.n5 a_n2018_n4888# 0.397899f
C105 source.t12 a_n2018_n4888# 3.96021f
C106 source.n6 a_n2018_n4888# 0.397899f
C107 source.t8 a_n2018_n4888# 0.346523f
C108 source.t7 a_n2018_n4888# 0.346523f
C109 source.n7 a_n2018_n4888# 3.09806f
C110 source.n8 a_n2018_n4888# 0.338426f
C111 source.t10 a_n2018_n4888# 0.346523f
C112 source.t15 a_n2018_n4888# 0.346523f
C113 source.n9 a_n2018_n4888# 3.09806f
C114 source.n10 a_n2018_n4888# 0.338426f
C115 source.t9 a_n2018_n4888# 3.96021f
C116 source.n11 a_n2018_n4888# 2.10949f
C117 source.t23 a_n2018_n4888# 3.96018f
C118 source.n12 a_n2018_n4888# 2.10951f
C119 source.t0 a_n2018_n4888# 0.346523f
C120 source.t22 a_n2018_n4888# 0.346523f
C121 source.n13 a_n2018_n4888# 3.09807f
C122 source.n14 a_n2018_n4888# 0.33842f
C123 source.t3 a_n2018_n4888# 0.346523f
C124 source.t1 a_n2018_n4888# 0.346523f
C125 source.n15 a_n2018_n4888# 3.09807f
C126 source.n16 a_n2018_n4888# 0.33842f
C127 source.t4 a_n2018_n4888# 3.96018f
C128 source.n17 a_n2018_n4888# 0.397921f
C129 source.t11 a_n2018_n4888# 3.96018f
C130 source.n18 a_n2018_n4888# 0.397921f
C131 source.t14 a_n2018_n4888# 0.346523f
C132 source.t17 a_n2018_n4888# 0.346523f
C133 source.n19 a_n2018_n4888# 3.09807f
C134 source.n20 a_n2018_n4888# 0.33842f
C135 source.t18 a_n2018_n4888# 0.346523f
C136 source.t13 a_n2018_n4888# 0.346523f
C137 source.n21 a_n2018_n4888# 3.09807f
C138 source.n22 a_n2018_n4888# 0.33842f
C139 source.t16 a_n2018_n4888# 3.96018f
C140 source.n23 a_n2018_n4888# 0.536169f
C141 source.n24 a_n2018_n4888# 1.98524f
C142 minus.n0 a_n2018_n4888# 0.043738f
C143 minus.t6 a_n2018_n4888# 1.48634f
C144 minus.n1 a_n2018_n4888# 0.56629f
C145 minus.t2 a_n2018_n4888# 1.48634f
C146 minus.t10 a_n2018_n4888# 1.50193f
C147 minus.n2 a_n2018_n4888# 0.543645f
C148 minus.t9 a_n2018_n4888# 1.48634f
C149 minus.n3 a_n2018_n4888# 0.564693f
C150 minus.t8 a_n2018_n4888# 1.48634f
C151 minus.n4 a_n2018_n4888# 0.56629f
C152 minus.n5 a_n2018_n4888# 0.224165f
C153 minus.n6 a_n2018_n4888# 0.072852f
C154 minus.n7 a_n2018_n4888# 0.058363f
C155 minus.n8 a_n2018_n4888# 0.557848f
C156 minus.n9 a_n2018_n4888# 0.009925f
C157 minus.t3 a_n2018_n4888# 1.48634f
C158 minus.n10 a_n2018_n4888# 0.554881f
C159 minus.n11 a_n2018_n4888# 2.0016f
C160 minus.n12 a_n2018_n4888# 0.043738f
C161 minus.t0 a_n2018_n4888# 1.48634f
C162 minus.n13 a_n2018_n4888# 0.56629f
C163 minus.t11 a_n2018_n4888# 1.50193f
C164 minus.n14 a_n2018_n4888# 0.543645f
C165 minus.t5 a_n2018_n4888# 1.48634f
C166 minus.n15 a_n2018_n4888# 0.564693f
C167 minus.t7 a_n2018_n4888# 1.48634f
C168 minus.n16 a_n2018_n4888# 0.56629f
C169 minus.n17 a_n2018_n4888# 0.224165f
C170 minus.n18 a_n2018_n4888# 0.072852f
C171 minus.n19 a_n2018_n4888# 0.058363f
C172 minus.t4 a_n2018_n4888# 1.48634f
C173 minus.n20 a_n2018_n4888# 0.557848f
C174 minus.n21 a_n2018_n4888# 0.009925f
C175 minus.t1 a_n2018_n4888# 1.48634f
C176 minus.n22 a_n2018_n4888# 0.554881f
C177 minus.n23 a_n2018_n4888# 0.294941f
C178 minus.n24 a_n2018_n4888# 2.38205f
.ends

