* NGSPICE file created from diffpair315.ext - technology: sky130A

.subckt diffpair315 minus drain_right drain_left source plus
X0 source.t21 plus.t0 drain_left.t3 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X1 drain_right.t11 minus.t0 source.t22 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X3 a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X4 drain_left.t10 plus.t1 source.t20 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X5 drain_left.t4 plus.t2 source.t19 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X6 a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X7 source.t9 minus.t1 drain_right.t10 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X8 a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X9 drain_right.t9 minus.t2 source.t0 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X10 drain_left.t2 plus.t3 source.t18 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X11 source.t6 minus.t3 drain_right.t8 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X12 source.t7 minus.t4 drain_right.t7 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X13 source.t8 minus.t5 drain_right.t6 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X14 source.t17 plus.t4 drain_left.t5 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X15 drain_right.t5 minus.t6 source.t3 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X16 source.t5 minus.t7 drain_right.t4 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X17 source.t4 minus.t8 drain_right.t3 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X18 drain_right.t2 minus.t9 source.t2 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X19 drain_left.t7 plus.t5 source.t16 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X20 drain_left.t8 plus.t6 source.t15 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X21 source.t14 plus.t7 drain_left.t0 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X22 drain_right.t1 minus.t10 source.t23 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X23 source.t13 plus.t8 drain_left.t11 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X24 drain_left.t1 plus.t9 source.t12 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X25 source.t11 plus.t10 drain_left.t6 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X26 drain_right.t0 minus.t11 source.t1 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X27 source.t10 plus.t11 drain_left.t9 a_n2298_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
R0 plus.n4 plus.t10 251.25
R1 plus.n20 plus.t3 251.25
R2 plus.n14 plus.t5 229.855
R3 plus.n12 plus.t8 229.855
R4 plus.n2 plus.t6 229.855
R5 plus.n7 plus.t7 229.855
R6 plus.n5 plus.t9 229.855
R7 plus.n30 plus.t4 229.855
R8 plus.n28 plus.t2 229.855
R9 plus.n18 plus.t11 229.855
R10 plus.n23 plus.t1 229.855
R11 plus.n21 plus.t0 229.855
R12 plus.n6 plus.n3 161.3
R13 plus.n11 plus.n10 161.3
R14 plus.n12 plus.n1 161.3
R15 plus.n13 plus.n0 161.3
R16 plus.n15 plus.n14 161.3
R17 plus.n22 plus.n19 161.3
R18 plus.n27 plus.n26 161.3
R19 plus.n28 plus.n17 161.3
R20 plus.n29 plus.n16 161.3
R21 plus.n31 plus.n30 161.3
R22 plus.n8 plus.n7 80.6037
R23 plus.n9 plus.n2 80.6037
R24 plus.n24 plus.n23 80.6037
R25 plus.n25 plus.n18 80.6037
R26 plus.n7 plus.n2 48.2005
R27 plus.n23 plus.n18 48.2005
R28 plus.n4 plus.n3 44.853
R29 plus.n20 plus.n19 44.853
R30 plus.n11 plus.n2 41.6278
R31 plus.n7 plus.n6 41.6278
R32 plus.n27 plus.n18 41.6278
R33 plus.n23 plus.n22 41.6278
R34 plus plus.n31 29.6354
R35 plus.n14 plus.n13 25.5611
R36 plus.n30 plus.n29 25.5611
R37 plus.n13 plus.n12 22.6399
R38 plus.n29 plus.n28 22.6399
R39 plus.n5 plus.n4 20.5405
R40 plus.n21 plus.n20 20.5405
R41 plus plus.n15 10.0725
R42 plus.n12 plus.n11 6.57323
R43 plus.n6 plus.n5 6.57323
R44 plus.n28 plus.n27 6.57323
R45 plus.n22 plus.n21 6.57323
R46 plus.n9 plus.n8 0.380177
R47 plus.n25 plus.n24 0.380177
R48 plus.n8 plus.n3 0.285035
R49 plus.n10 plus.n9 0.285035
R50 plus.n26 plus.n25 0.285035
R51 plus.n24 plus.n19 0.285035
R52 plus.n10 plus.n1 0.189894
R53 plus.n1 plus.n0 0.189894
R54 plus.n15 plus.n0 0.189894
R55 plus.n31 plus.n16 0.189894
R56 plus.n17 plus.n16 0.189894
R57 plus.n26 plus.n17 0.189894
R58 drain_left.n6 drain_left.n4 68.165
R59 drain_left.n3 drain_left.n2 68.1095
R60 drain_left.n3 drain_left.n0 68.1095
R61 drain_left.n6 drain_left.n5 67.1908
R62 drain_left.n8 drain_left.n7 67.1907
R63 drain_left.n3 drain_left.n1 67.1907
R64 drain_left drain_left.n3 27.6923
R65 drain_left drain_left.n8 6.62735
R66 drain_left.n1 drain_left.t9 3.3005
R67 drain_left.n1 drain_left.t10 3.3005
R68 drain_left.n2 drain_left.t3 3.3005
R69 drain_left.n2 drain_left.t2 3.3005
R70 drain_left.n0 drain_left.t5 3.3005
R71 drain_left.n0 drain_left.t4 3.3005
R72 drain_left.n7 drain_left.t11 3.3005
R73 drain_left.n7 drain_left.t7 3.3005
R74 drain_left.n5 drain_left.t0 3.3005
R75 drain_left.n5 drain_left.t8 3.3005
R76 drain_left.n4 drain_left.t6 3.3005
R77 drain_left.n4 drain_left.t1 3.3005
R78 drain_left.n8 drain_left.n6 0.974638
R79 source.n266 source.n240 289.615
R80 source.n230 source.n204 289.615
R81 source.n198 source.n172 289.615
R82 source.n162 source.n136 289.615
R83 source.n26 source.n0 289.615
R84 source.n62 source.n36 289.615
R85 source.n94 source.n68 289.615
R86 source.n130 source.n104 289.615
R87 source.n251 source.n250 185
R88 source.n248 source.n247 185
R89 source.n257 source.n256 185
R90 source.n259 source.n258 185
R91 source.n244 source.n243 185
R92 source.n265 source.n264 185
R93 source.n267 source.n266 185
R94 source.n215 source.n214 185
R95 source.n212 source.n211 185
R96 source.n221 source.n220 185
R97 source.n223 source.n222 185
R98 source.n208 source.n207 185
R99 source.n229 source.n228 185
R100 source.n231 source.n230 185
R101 source.n183 source.n182 185
R102 source.n180 source.n179 185
R103 source.n189 source.n188 185
R104 source.n191 source.n190 185
R105 source.n176 source.n175 185
R106 source.n197 source.n196 185
R107 source.n199 source.n198 185
R108 source.n147 source.n146 185
R109 source.n144 source.n143 185
R110 source.n153 source.n152 185
R111 source.n155 source.n154 185
R112 source.n140 source.n139 185
R113 source.n161 source.n160 185
R114 source.n163 source.n162 185
R115 source.n27 source.n26 185
R116 source.n25 source.n24 185
R117 source.n4 source.n3 185
R118 source.n19 source.n18 185
R119 source.n17 source.n16 185
R120 source.n8 source.n7 185
R121 source.n11 source.n10 185
R122 source.n63 source.n62 185
R123 source.n61 source.n60 185
R124 source.n40 source.n39 185
R125 source.n55 source.n54 185
R126 source.n53 source.n52 185
R127 source.n44 source.n43 185
R128 source.n47 source.n46 185
R129 source.n95 source.n94 185
R130 source.n93 source.n92 185
R131 source.n72 source.n71 185
R132 source.n87 source.n86 185
R133 source.n85 source.n84 185
R134 source.n76 source.n75 185
R135 source.n79 source.n78 185
R136 source.n131 source.n130 185
R137 source.n129 source.n128 185
R138 source.n108 source.n107 185
R139 source.n123 source.n122 185
R140 source.n121 source.n120 185
R141 source.n112 source.n111 185
R142 source.n115 source.n114 185
R143 source.t23 source.n249 147.661
R144 source.t8 source.n213 147.661
R145 source.t18 source.n181 147.661
R146 source.t17 source.n145 147.661
R147 source.t16 source.n9 147.661
R148 source.t11 source.n45 147.661
R149 source.t3 source.n77 147.661
R150 source.t5 source.n113 147.661
R151 source.n250 source.n247 104.615
R152 source.n257 source.n247 104.615
R153 source.n258 source.n257 104.615
R154 source.n258 source.n243 104.615
R155 source.n265 source.n243 104.615
R156 source.n266 source.n265 104.615
R157 source.n214 source.n211 104.615
R158 source.n221 source.n211 104.615
R159 source.n222 source.n221 104.615
R160 source.n222 source.n207 104.615
R161 source.n229 source.n207 104.615
R162 source.n230 source.n229 104.615
R163 source.n182 source.n179 104.615
R164 source.n189 source.n179 104.615
R165 source.n190 source.n189 104.615
R166 source.n190 source.n175 104.615
R167 source.n197 source.n175 104.615
R168 source.n198 source.n197 104.615
R169 source.n146 source.n143 104.615
R170 source.n153 source.n143 104.615
R171 source.n154 source.n153 104.615
R172 source.n154 source.n139 104.615
R173 source.n161 source.n139 104.615
R174 source.n162 source.n161 104.615
R175 source.n26 source.n25 104.615
R176 source.n25 source.n3 104.615
R177 source.n18 source.n3 104.615
R178 source.n18 source.n17 104.615
R179 source.n17 source.n7 104.615
R180 source.n10 source.n7 104.615
R181 source.n62 source.n61 104.615
R182 source.n61 source.n39 104.615
R183 source.n54 source.n39 104.615
R184 source.n54 source.n53 104.615
R185 source.n53 source.n43 104.615
R186 source.n46 source.n43 104.615
R187 source.n94 source.n93 104.615
R188 source.n93 source.n71 104.615
R189 source.n86 source.n71 104.615
R190 source.n86 source.n85 104.615
R191 source.n85 source.n75 104.615
R192 source.n78 source.n75 104.615
R193 source.n130 source.n129 104.615
R194 source.n129 source.n107 104.615
R195 source.n122 source.n107 104.615
R196 source.n122 source.n121 104.615
R197 source.n121 source.n111 104.615
R198 source.n114 source.n111 104.615
R199 source.n250 source.t23 52.3082
R200 source.n214 source.t8 52.3082
R201 source.n182 source.t18 52.3082
R202 source.n146 source.t17 52.3082
R203 source.n10 source.t16 52.3082
R204 source.n46 source.t11 52.3082
R205 source.n78 source.t3 52.3082
R206 source.n114 source.t5 52.3082
R207 source.n33 source.n32 50.512
R208 source.n35 source.n34 50.512
R209 source.n101 source.n100 50.512
R210 source.n103 source.n102 50.512
R211 source.n239 source.n238 50.5119
R212 source.n237 source.n236 50.5119
R213 source.n171 source.n170 50.5119
R214 source.n169 source.n168 50.5119
R215 source.n271 source.n270 32.1853
R216 source.n235 source.n234 32.1853
R217 source.n203 source.n202 32.1853
R218 source.n167 source.n166 32.1853
R219 source.n31 source.n30 32.1853
R220 source.n67 source.n66 32.1853
R221 source.n99 source.n98 32.1853
R222 source.n135 source.n134 32.1853
R223 source.n167 source.n135 17.7164
R224 source.n251 source.n249 15.6674
R225 source.n215 source.n213 15.6674
R226 source.n183 source.n181 15.6674
R227 source.n147 source.n145 15.6674
R228 source.n11 source.n9 15.6674
R229 source.n47 source.n45 15.6674
R230 source.n79 source.n77 15.6674
R231 source.n115 source.n113 15.6674
R232 source.n252 source.n248 12.8005
R233 source.n216 source.n212 12.8005
R234 source.n184 source.n180 12.8005
R235 source.n148 source.n144 12.8005
R236 source.n12 source.n8 12.8005
R237 source.n48 source.n44 12.8005
R238 source.n80 source.n76 12.8005
R239 source.n116 source.n112 12.8005
R240 source.n256 source.n255 12.0247
R241 source.n220 source.n219 12.0247
R242 source.n188 source.n187 12.0247
R243 source.n152 source.n151 12.0247
R244 source.n16 source.n15 12.0247
R245 source.n52 source.n51 12.0247
R246 source.n84 source.n83 12.0247
R247 source.n120 source.n119 12.0247
R248 source.n272 source.n31 11.9664
R249 source.n259 source.n246 11.249
R250 source.n223 source.n210 11.249
R251 source.n191 source.n178 11.249
R252 source.n155 source.n142 11.249
R253 source.n19 source.n6 11.249
R254 source.n55 source.n42 11.249
R255 source.n87 source.n74 11.249
R256 source.n123 source.n110 11.249
R257 source.n260 source.n244 10.4732
R258 source.n224 source.n208 10.4732
R259 source.n192 source.n176 10.4732
R260 source.n156 source.n140 10.4732
R261 source.n20 source.n4 10.4732
R262 source.n56 source.n40 10.4732
R263 source.n88 source.n72 10.4732
R264 source.n124 source.n108 10.4732
R265 source.n264 source.n263 9.69747
R266 source.n228 source.n227 9.69747
R267 source.n196 source.n195 9.69747
R268 source.n160 source.n159 9.69747
R269 source.n24 source.n23 9.69747
R270 source.n60 source.n59 9.69747
R271 source.n92 source.n91 9.69747
R272 source.n128 source.n127 9.69747
R273 source.n270 source.n269 9.45567
R274 source.n234 source.n233 9.45567
R275 source.n202 source.n201 9.45567
R276 source.n166 source.n165 9.45567
R277 source.n30 source.n29 9.45567
R278 source.n66 source.n65 9.45567
R279 source.n98 source.n97 9.45567
R280 source.n134 source.n133 9.45567
R281 source.n269 source.n268 9.3005
R282 source.n242 source.n241 9.3005
R283 source.n263 source.n262 9.3005
R284 source.n261 source.n260 9.3005
R285 source.n246 source.n245 9.3005
R286 source.n255 source.n254 9.3005
R287 source.n253 source.n252 9.3005
R288 source.n233 source.n232 9.3005
R289 source.n206 source.n205 9.3005
R290 source.n227 source.n226 9.3005
R291 source.n225 source.n224 9.3005
R292 source.n210 source.n209 9.3005
R293 source.n219 source.n218 9.3005
R294 source.n217 source.n216 9.3005
R295 source.n201 source.n200 9.3005
R296 source.n174 source.n173 9.3005
R297 source.n195 source.n194 9.3005
R298 source.n193 source.n192 9.3005
R299 source.n178 source.n177 9.3005
R300 source.n187 source.n186 9.3005
R301 source.n185 source.n184 9.3005
R302 source.n165 source.n164 9.3005
R303 source.n138 source.n137 9.3005
R304 source.n159 source.n158 9.3005
R305 source.n157 source.n156 9.3005
R306 source.n142 source.n141 9.3005
R307 source.n151 source.n150 9.3005
R308 source.n149 source.n148 9.3005
R309 source.n29 source.n28 9.3005
R310 source.n2 source.n1 9.3005
R311 source.n23 source.n22 9.3005
R312 source.n21 source.n20 9.3005
R313 source.n6 source.n5 9.3005
R314 source.n15 source.n14 9.3005
R315 source.n13 source.n12 9.3005
R316 source.n65 source.n64 9.3005
R317 source.n38 source.n37 9.3005
R318 source.n59 source.n58 9.3005
R319 source.n57 source.n56 9.3005
R320 source.n42 source.n41 9.3005
R321 source.n51 source.n50 9.3005
R322 source.n49 source.n48 9.3005
R323 source.n97 source.n96 9.3005
R324 source.n70 source.n69 9.3005
R325 source.n91 source.n90 9.3005
R326 source.n89 source.n88 9.3005
R327 source.n74 source.n73 9.3005
R328 source.n83 source.n82 9.3005
R329 source.n81 source.n80 9.3005
R330 source.n133 source.n132 9.3005
R331 source.n106 source.n105 9.3005
R332 source.n127 source.n126 9.3005
R333 source.n125 source.n124 9.3005
R334 source.n110 source.n109 9.3005
R335 source.n119 source.n118 9.3005
R336 source.n117 source.n116 9.3005
R337 source.n267 source.n242 8.92171
R338 source.n231 source.n206 8.92171
R339 source.n199 source.n174 8.92171
R340 source.n163 source.n138 8.92171
R341 source.n27 source.n2 8.92171
R342 source.n63 source.n38 8.92171
R343 source.n95 source.n70 8.92171
R344 source.n131 source.n106 8.92171
R345 source.n268 source.n240 8.14595
R346 source.n232 source.n204 8.14595
R347 source.n200 source.n172 8.14595
R348 source.n164 source.n136 8.14595
R349 source.n28 source.n0 8.14595
R350 source.n64 source.n36 8.14595
R351 source.n96 source.n68 8.14595
R352 source.n132 source.n104 8.14595
R353 source.n270 source.n240 5.81868
R354 source.n234 source.n204 5.81868
R355 source.n202 source.n172 5.81868
R356 source.n166 source.n136 5.81868
R357 source.n30 source.n0 5.81868
R358 source.n66 source.n36 5.81868
R359 source.n98 source.n68 5.81868
R360 source.n134 source.n104 5.81868
R361 source.n272 source.n271 5.7505
R362 source.n268 source.n267 5.04292
R363 source.n232 source.n231 5.04292
R364 source.n200 source.n199 5.04292
R365 source.n164 source.n163 5.04292
R366 source.n28 source.n27 5.04292
R367 source.n64 source.n63 5.04292
R368 source.n96 source.n95 5.04292
R369 source.n132 source.n131 5.04292
R370 source.n253 source.n249 4.38594
R371 source.n217 source.n213 4.38594
R372 source.n185 source.n181 4.38594
R373 source.n149 source.n145 4.38594
R374 source.n13 source.n9 4.38594
R375 source.n49 source.n45 4.38594
R376 source.n81 source.n77 4.38594
R377 source.n117 source.n113 4.38594
R378 source.n264 source.n242 4.26717
R379 source.n228 source.n206 4.26717
R380 source.n196 source.n174 4.26717
R381 source.n160 source.n138 4.26717
R382 source.n24 source.n2 4.26717
R383 source.n60 source.n38 4.26717
R384 source.n92 source.n70 4.26717
R385 source.n128 source.n106 4.26717
R386 source.n263 source.n244 3.49141
R387 source.n227 source.n208 3.49141
R388 source.n195 source.n176 3.49141
R389 source.n159 source.n140 3.49141
R390 source.n23 source.n4 3.49141
R391 source.n59 source.n40 3.49141
R392 source.n91 source.n72 3.49141
R393 source.n127 source.n108 3.49141
R394 source.n238 source.t1 3.3005
R395 source.n238 source.t6 3.3005
R396 source.n236 source.t22 3.3005
R397 source.n236 source.t9 3.3005
R398 source.n170 source.t20 3.3005
R399 source.n170 source.t21 3.3005
R400 source.n168 source.t19 3.3005
R401 source.n168 source.t10 3.3005
R402 source.n32 source.t15 3.3005
R403 source.n32 source.t13 3.3005
R404 source.n34 source.t12 3.3005
R405 source.n34 source.t14 3.3005
R406 source.n100 source.t0 3.3005
R407 source.n100 source.t7 3.3005
R408 source.n102 source.t2 3.3005
R409 source.n102 source.t4 3.3005
R410 source.n260 source.n259 2.71565
R411 source.n224 source.n223 2.71565
R412 source.n192 source.n191 2.71565
R413 source.n156 source.n155 2.71565
R414 source.n20 source.n19 2.71565
R415 source.n56 source.n55 2.71565
R416 source.n88 source.n87 2.71565
R417 source.n124 source.n123 2.71565
R418 source.n256 source.n246 1.93989
R419 source.n220 source.n210 1.93989
R420 source.n188 source.n178 1.93989
R421 source.n152 source.n142 1.93989
R422 source.n16 source.n6 1.93989
R423 source.n52 source.n42 1.93989
R424 source.n84 source.n74 1.93989
R425 source.n120 source.n110 1.93989
R426 source.n255 source.n248 1.16414
R427 source.n219 source.n212 1.16414
R428 source.n187 source.n180 1.16414
R429 source.n151 source.n144 1.16414
R430 source.n15 source.n8 1.16414
R431 source.n51 source.n44 1.16414
R432 source.n83 source.n76 1.16414
R433 source.n119 source.n112 1.16414
R434 source.n135 source.n103 0.974638
R435 source.n103 source.n101 0.974638
R436 source.n101 source.n99 0.974638
R437 source.n67 source.n35 0.974638
R438 source.n35 source.n33 0.974638
R439 source.n33 source.n31 0.974638
R440 source.n169 source.n167 0.974638
R441 source.n171 source.n169 0.974638
R442 source.n203 source.n171 0.974638
R443 source.n237 source.n235 0.974638
R444 source.n239 source.n237 0.974638
R445 source.n271 source.n239 0.974638
R446 source.n99 source.n67 0.470328
R447 source.n235 source.n203 0.470328
R448 source.n252 source.n251 0.388379
R449 source.n216 source.n215 0.388379
R450 source.n184 source.n183 0.388379
R451 source.n148 source.n147 0.388379
R452 source.n12 source.n11 0.388379
R453 source.n48 source.n47 0.388379
R454 source.n80 source.n79 0.388379
R455 source.n116 source.n115 0.388379
R456 source source.n272 0.188
R457 source.n254 source.n253 0.155672
R458 source.n254 source.n245 0.155672
R459 source.n261 source.n245 0.155672
R460 source.n262 source.n261 0.155672
R461 source.n262 source.n241 0.155672
R462 source.n269 source.n241 0.155672
R463 source.n218 source.n217 0.155672
R464 source.n218 source.n209 0.155672
R465 source.n225 source.n209 0.155672
R466 source.n226 source.n225 0.155672
R467 source.n226 source.n205 0.155672
R468 source.n233 source.n205 0.155672
R469 source.n186 source.n185 0.155672
R470 source.n186 source.n177 0.155672
R471 source.n193 source.n177 0.155672
R472 source.n194 source.n193 0.155672
R473 source.n194 source.n173 0.155672
R474 source.n201 source.n173 0.155672
R475 source.n150 source.n149 0.155672
R476 source.n150 source.n141 0.155672
R477 source.n157 source.n141 0.155672
R478 source.n158 source.n157 0.155672
R479 source.n158 source.n137 0.155672
R480 source.n165 source.n137 0.155672
R481 source.n29 source.n1 0.155672
R482 source.n22 source.n1 0.155672
R483 source.n22 source.n21 0.155672
R484 source.n21 source.n5 0.155672
R485 source.n14 source.n5 0.155672
R486 source.n14 source.n13 0.155672
R487 source.n65 source.n37 0.155672
R488 source.n58 source.n37 0.155672
R489 source.n58 source.n57 0.155672
R490 source.n57 source.n41 0.155672
R491 source.n50 source.n41 0.155672
R492 source.n50 source.n49 0.155672
R493 source.n97 source.n69 0.155672
R494 source.n90 source.n69 0.155672
R495 source.n90 source.n89 0.155672
R496 source.n89 source.n73 0.155672
R497 source.n82 source.n73 0.155672
R498 source.n82 source.n81 0.155672
R499 source.n133 source.n105 0.155672
R500 source.n126 source.n105 0.155672
R501 source.n126 source.n125 0.155672
R502 source.n125 source.n109 0.155672
R503 source.n118 source.n109 0.155672
R504 source.n118 source.n117 0.155672
R505 minus.n4 minus.t6 251.25
R506 minus.n20 minus.t5 251.25
R507 minus.n3 minus.t4 229.855
R508 minus.n7 minus.t2 229.855
R509 minus.n8 minus.t8 229.855
R510 minus.n12 minus.t9 229.855
R511 minus.n14 minus.t7 229.855
R512 minus.n19 minus.t0 229.855
R513 minus.n23 minus.t1 229.855
R514 minus.n24 minus.t11 229.855
R515 minus.n28 minus.t3 229.855
R516 minus.n30 minus.t10 229.855
R517 minus.n15 minus.n14 161.3
R518 minus.n13 minus.n0 161.3
R519 minus.n12 minus.n11 161.3
R520 minus.n10 minus.n1 161.3
R521 minus.n6 minus.n5 161.3
R522 minus.n31 minus.n30 161.3
R523 minus.n29 minus.n16 161.3
R524 minus.n28 minus.n27 161.3
R525 minus.n26 minus.n17 161.3
R526 minus.n22 minus.n21 161.3
R527 minus.n9 minus.n8 80.6037
R528 minus.n7 minus.n2 80.6037
R529 minus.n25 minus.n24 80.6037
R530 minus.n23 minus.n18 80.6037
R531 minus.n8 minus.n7 48.2005
R532 minus.n24 minus.n23 48.2005
R533 minus.n5 minus.n4 44.853
R534 minus.n21 minus.n20 44.853
R535 minus.n7 minus.n6 41.6278
R536 minus.n8 minus.n1 41.6278
R537 minus.n23 minus.n22 41.6278
R538 minus.n24 minus.n17 41.6278
R539 minus.n32 minus.n15 33.4816
R540 minus.n14 minus.n13 25.5611
R541 minus.n30 minus.n29 25.5611
R542 minus.n13 minus.n12 22.6399
R543 minus.n29 minus.n28 22.6399
R544 minus.n4 minus.n3 20.5405
R545 minus.n20 minus.n19 20.5405
R546 minus.n32 minus.n31 6.70126
R547 minus.n6 minus.n3 6.57323
R548 minus.n12 minus.n1 6.57323
R549 minus.n22 minus.n19 6.57323
R550 minus.n28 minus.n17 6.57323
R551 minus.n9 minus.n2 0.380177
R552 minus.n25 minus.n18 0.380177
R553 minus.n10 minus.n9 0.285035
R554 minus.n5 minus.n2 0.285035
R555 minus.n21 minus.n18 0.285035
R556 minus.n26 minus.n25 0.285035
R557 minus.n15 minus.n0 0.189894
R558 minus.n11 minus.n0 0.189894
R559 minus.n11 minus.n10 0.189894
R560 minus.n27 minus.n26 0.189894
R561 minus.n27 minus.n16 0.189894
R562 minus.n31 minus.n16 0.189894
R563 minus minus.n32 0.188
R564 drain_right.n6 drain_right.n4 68.1648
R565 drain_right.n3 drain_right.n2 68.1095
R566 drain_right.n3 drain_right.n0 68.1095
R567 drain_right.n6 drain_right.n5 67.1908
R568 drain_right.n8 drain_right.n7 67.1908
R569 drain_right.n3 drain_right.n1 67.1907
R570 drain_right drain_right.n3 27.1391
R571 drain_right drain_right.n8 6.62735
R572 drain_right.n1 drain_right.t10 3.3005
R573 drain_right.n1 drain_right.t0 3.3005
R574 drain_right.n2 drain_right.t8 3.3005
R575 drain_right.n2 drain_right.t1 3.3005
R576 drain_right.n0 drain_right.t6 3.3005
R577 drain_right.n0 drain_right.t11 3.3005
R578 drain_right.n4 drain_right.t7 3.3005
R579 drain_right.n4 drain_right.t5 3.3005
R580 drain_right.n5 drain_right.t3 3.3005
R581 drain_right.n5 drain_right.t9 3.3005
R582 drain_right.n7 drain_right.t4 3.3005
R583 drain_right.n7 drain_right.t2 3.3005
R584 drain_right.n8 drain_right.n6 0.974638
C0 source drain_right 8.759339f
C1 source plus 4.76062f
C2 source minus 4.7466f
C3 drain_left drain_right 1.16185f
C4 plus drain_left 4.70491f
C5 minus drain_left 0.17224f
C6 plus drain_right 0.381869f
C7 minus drain_right 4.4786f
C8 minus plus 4.89443f
C9 source drain_left 8.75678f
C10 drain_right a_n2298_n2088# 5.17693f
C11 drain_left a_n2298_n2088# 5.50628f
C12 source a_n2298_n2088# 5.613978f
C13 minus a_n2298_n2088# 8.568169f
C14 plus a_n2298_n2088# 9.95917f
C15 drain_right.t6 a_n2298_n2088# 0.125124f
C16 drain_right.t11 a_n2298_n2088# 0.125124f
C17 drain_right.n0 a_n2298_n2088# 1.04874f
C18 drain_right.t10 a_n2298_n2088# 0.125124f
C19 drain_right.t0 a_n2298_n2088# 0.125124f
C20 drain_right.n1 a_n2298_n2088# 1.04353f
C21 drain_right.t8 a_n2298_n2088# 0.125124f
C22 drain_right.t1 a_n2298_n2088# 0.125124f
C23 drain_right.n2 a_n2298_n2088# 1.04874f
C24 drain_right.n3 a_n2298_n2088# 2.10833f
C25 drain_right.t7 a_n2298_n2088# 0.125124f
C26 drain_right.t5 a_n2298_n2088# 0.125124f
C27 drain_right.n4 a_n2298_n2088# 1.04911f
C28 drain_right.t3 a_n2298_n2088# 0.125124f
C29 drain_right.t9 a_n2298_n2088# 0.125124f
C30 drain_right.n5 a_n2298_n2088# 1.04354f
C31 drain_right.n6 a_n2298_n2088# 0.764757f
C32 drain_right.t4 a_n2298_n2088# 0.125124f
C33 drain_right.t2 a_n2298_n2088# 0.125124f
C34 drain_right.n7 a_n2298_n2088# 1.04354f
C35 drain_right.n8 a_n2298_n2088# 0.616486f
C36 minus.n0 a_n2298_n2088# 0.040764f
C37 minus.n1 a_n2298_n2088# 0.00925f
C38 minus.t9 a_n2298_n2088# 0.567543f
C39 minus.n2 a_n2298_n2088# 0.067897f
C40 minus.t4 a_n2298_n2088# 0.567543f
C41 minus.n3 a_n2298_n2088# 0.261705f
C42 minus.t6 a_n2298_n2088# 0.589751f
C43 minus.n4 a_n2298_n2088# 0.242626f
C44 minus.n5 a_n2298_n2088# 0.187138f
C45 minus.n6 a_n2298_n2088# 0.00925f
C46 minus.t2 a_n2298_n2088# 0.567543f
C47 minus.n7 a_n2298_n2088# 0.269915f
C48 minus.t8 a_n2298_n2088# 0.567543f
C49 minus.n8 a_n2298_n2088# 0.269915f
C50 minus.n9 a_n2298_n2088# 0.067897f
C51 minus.n10 a_n2298_n2088# 0.054394f
C52 minus.n11 a_n2298_n2088# 0.040764f
C53 minus.n12 a_n2298_n2088# 0.258529f
C54 minus.n13 a_n2298_n2088# 0.00925f
C55 minus.t7 a_n2298_n2088# 0.567543f
C56 minus.n14 a_n2298_n2088# 0.257901f
C57 minus.n15 a_n2298_n2088# 1.2796f
C58 minus.n16 a_n2298_n2088# 0.040764f
C59 minus.n17 a_n2298_n2088# 0.00925f
C60 minus.n18 a_n2298_n2088# 0.067897f
C61 minus.t0 a_n2298_n2088# 0.567543f
C62 minus.n19 a_n2298_n2088# 0.261705f
C63 minus.t5 a_n2298_n2088# 0.589751f
C64 minus.n20 a_n2298_n2088# 0.242626f
C65 minus.n21 a_n2298_n2088# 0.187138f
C66 minus.n22 a_n2298_n2088# 0.00925f
C67 minus.t1 a_n2298_n2088# 0.567543f
C68 minus.n23 a_n2298_n2088# 0.269915f
C69 minus.t11 a_n2298_n2088# 0.567543f
C70 minus.n24 a_n2298_n2088# 0.269915f
C71 minus.n25 a_n2298_n2088# 0.067897f
C72 minus.n26 a_n2298_n2088# 0.054394f
C73 minus.n27 a_n2298_n2088# 0.040764f
C74 minus.t3 a_n2298_n2088# 0.567543f
C75 minus.n28 a_n2298_n2088# 0.258529f
C76 minus.n29 a_n2298_n2088# 0.00925f
C77 minus.t10 a_n2298_n2088# 0.567543f
C78 minus.n30 a_n2298_n2088# 0.257901f
C79 minus.n31 a_n2298_n2088# 0.285653f
C80 minus.n32 a_n2298_n2088# 1.55866f
C81 source.n0 a_n2298_n2088# 0.033197f
C82 source.n1 a_n2298_n2088# 0.023618f
C83 source.n2 a_n2298_n2088# 0.012691f
C84 source.n3 a_n2298_n2088# 0.029998f
C85 source.n4 a_n2298_n2088# 0.013438f
C86 source.n5 a_n2298_n2088# 0.023618f
C87 source.n6 a_n2298_n2088# 0.012691f
C88 source.n7 a_n2298_n2088# 0.029998f
C89 source.n8 a_n2298_n2088# 0.013438f
C90 source.n9 a_n2298_n2088# 0.101069f
C91 source.t16 a_n2298_n2088# 0.048893f
C92 source.n10 a_n2298_n2088# 0.022498f
C93 source.n11 a_n2298_n2088# 0.017719f
C94 source.n12 a_n2298_n2088# 0.012691f
C95 source.n13 a_n2298_n2088# 0.561971f
C96 source.n14 a_n2298_n2088# 0.023618f
C97 source.n15 a_n2298_n2088# 0.012691f
C98 source.n16 a_n2298_n2088# 0.013438f
C99 source.n17 a_n2298_n2088# 0.029998f
C100 source.n18 a_n2298_n2088# 0.029998f
C101 source.n19 a_n2298_n2088# 0.013438f
C102 source.n20 a_n2298_n2088# 0.012691f
C103 source.n21 a_n2298_n2088# 0.023618f
C104 source.n22 a_n2298_n2088# 0.023618f
C105 source.n23 a_n2298_n2088# 0.012691f
C106 source.n24 a_n2298_n2088# 0.013438f
C107 source.n25 a_n2298_n2088# 0.029998f
C108 source.n26 a_n2298_n2088# 0.06494f
C109 source.n27 a_n2298_n2088# 0.013438f
C110 source.n28 a_n2298_n2088# 0.012691f
C111 source.n29 a_n2298_n2088# 0.054592f
C112 source.n30 a_n2298_n2088# 0.036337f
C113 source.n31 a_n2298_n2088# 0.628194f
C114 source.t15 a_n2298_n2088# 0.111983f
C115 source.t13 a_n2298_n2088# 0.111983f
C116 source.n32 a_n2298_n2088# 0.872131f
C117 source.n33 a_n2298_n2088# 0.369667f
C118 source.t12 a_n2298_n2088# 0.111983f
C119 source.t14 a_n2298_n2088# 0.111983f
C120 source.n34 a_n2298_n2088# 0.872131f
C121 source.n35 a_n2298_n2088# 0.369667f
C122 source.n36 a_n2298_n2088# 0.033197f
C123 source.n37 a_n2298_n2088# 0.023618f
C124 source.n38 a_n2298_n2088# 0.012691f
C125 source.n39 a_n2298_n2088# 0.029998f
C126 source.n40 a_n2298_n2088# 0.013438f
C127 source.n41 a_n2298_n2088# 0.023618f
C128 source.n42 a_n2298_n2088# 0.012691f
C129 source.n43 a_n2298_n2088# 0.029998f
C130 source.n44 a_n2298_n2088# 0.013438f
C131 source.n45 a_n2298_n2088# 0.101069f
C132 source.t11 a_n2298_n2088# 0.048893f
C133 source.n46 a_n2298_n2088# 0.022498f
C134 source.n47 a_n2298_n2088# 0.017719f
C135 source.n48 a_n2298_n2088# 0.012691f
C136 source.n49 a_n2298_n2088# 0.561971f
C137 source.n50 a_n2298_n2088# 0.023618f
C138 source.n51 a_n2298_n2088# 0.012691f
C139 source.n52 a_n2298_n2088# 0.013438f
C140 source.n53 a_n2298_n2088# 0.029998f
C141 source.n54 a_n2298_n2088# 0.029998f
C142 source.n55 a_n2298_n2088# 0.013438f
C143 source.n56 a_n2298_n2088# 0.012691f
C144 source.n57 a_n2298_n2088# 0.023618f
C145 source.n58 a_n2298_n2088# 0.023618f
C146 source.n59 a_n2298_n2088# 0.012691f
C147 source.n60 a_n2298_n2088# 0.013438f
C148 source.n61 a_n2298_n2088# 0.029998f
C149 source.n62 a_n2298_n2088# 0.06494f
C150 source.n63 a_n2298_n2088# 0.013438f
C151 source.n64 a_n2298_n2088# 0.012691f
C152 source.n65 a_n2298_n2088# 0.054592f
C153 source.n66 a_n2298_n2088# 0.036337f
C154 source.n67 a_n2298_n2088# 0.130062f
C155 source.n68 a_n2298_n2088# 0.033197f
C156 source.n69 a_n2298_n2088# 0.023618f
C157 source.n70 a_n2298_n2088# 0.012691f
C158 source.n71 a_n2298_n2088# 0.029998f
C159 source.n72 a_n2298_n2088# 0.013438f
C160 source.n73 a_n2298_n2088# 0.023618f
C161 source.n74 a_n2298_n2088# 0.012691f
C162 source.n75 a_n2298_n2088# 0.029998f
C163 source.n76 a_n2298_n2088# 0.013438f
C164 source.n77 a_n2298_n2088# 0.101069f
C165 source.t3 a_n2298_n2088# 0.048893f
C166 source.n78 a_n2298_n2088# 0.022498f
C167 source.n79 a_n2298_n2088# 0.017719f
C168 source.n80 a_n2298_n2088# 0.012691f
C169 source.n81 a_n2298_n2088# 0.561971f
C170 source.n82 a_n2298_n2088# 0.023618f
C171 source.n83 a_n2298_n2088# 0.012691f
C172 source.n84 a_n2298_n2088# 0.013438f
C173 source.n85 a_n2298_n2088# 0.029998f
C174 source.n86 a_n2298_n2088# 0.029998f
C175 source.n87 a_n2298_n2088# 0.013438f
C176 source.n88 a_n2298_n2088# 0.012691f
C177 source.n89 a_n2298_n2088# 0.023618f
C178 source.n90 a_n2298_n2088# 0.023618f
C179 source.n91 a_n2298_n2088# 0.012691f
C180 source.n92 a_n2298_n2088# 0.013438f
C181 source.n93 a_n2298_n2088# 0.029998f
C182 source.n94 a_n2298_n2088# 0.06494f
C183 source.n95 a_n2298_n2088# 0.013438f
C184 source.n96 a_n2298_n2088# 0.012691f
C185 source.n97 a_n2298_n2088# 0.054592f
C186 source.n98 a_n2298_n2088# 0.036337f
C187 source.n99 a_n2298_n2088# 0.130062f
C188 source.t0 a_n2298_n2088# 0.111983f
C189 source.t7 a_n2298_n2088# 0.111983f
C190 source.n100 a_n2298_n2088# 0.872131f
C191 source.n101 a_n2298_n2088# 0.369667f
C192 source.t2 a_n2298_n2088# 0.111983f
C193 source.t4 a_n2298_n2088# 0.111983f
C194 source.n102 a_n2298_n2088# 0.872131f
C195 source.n103 a_n2298_n2088# 0.369667f
C196 source.n104 a_n2298_n2088# 0.033197f
C197 source.n105 a_n2298_n2088# 0.023618f
C198 source.n106 a_n2298_n2088# 0.012691f
C199 source.n107 a_n2298_n2088# 0.029998f
C200 source.n108 a_n2298_n2088# 0.013438f
C201 source.n109 a_n2298_n2088# 0.023618f
C202 source.n110 a_n2298_n2088# 0.012691f
C203 source.n111 a_n2298_n2088# 0.029998f
C204 source.n112 a_n2298_n2088# 0.013438f
C205 source.n113 a_n2298_n2088# 0.101069f
C206 source.t5 a_n2298_n2088# 0.048893f
C207 source.n114 a_n2298_n2088# 0.022498f
C208 source.n115 a_n2298_n2088# 0.017719f
C209 source.n116 a_n2298_n2088# 0.012691f
C210 source.n117 a_n2298_n2088# 0.561971f
C211 source.n118 a_n2298_n2088# 0.023618f
C212 source.n119 a_n2298_n2088# 0.012691f
C213 source.n120 a_n2298_n2088# 0.013438f
C214 source.n121 a_n2298_n2088# 0.029998f
C215 source.n122 a_n2298_n2088# 0.029998f
C216 source.n123 a_n2298_n2088# 0.013438f
C217 source.n124 a_n2298_n2088# 0.012691f
C218 source.n125 a_n2298_n2088# 0.023618f
C219 source.n126 a_n2298_n2088# 0.023618f
C220 source.n127 a_n2298_n2088# 0.012691f
C221 source.n128 a_n2298_n2088# 0.013438f
C222 source.n129 a_n2298_n2088# 0.029998f
C223 source.n130 a_n2298_n2088# 0.06494f
C224 source.n131 a_n2298_n2088# 0.013438f
C225 source.n132 a_n2298_n2088# 0.012691f
C226 source.n133 a_n2298_n2088# 0.054592f
C227 source.n134 a_n2298_n2088# 0.036337f
C228 source.n135 a_n2298_n2088# 0.941744f
C229 source.n136 a_n2298_n2088# 0.033197f
C230 source.n137 a_n2298_n2088# 0.023618f
C231 source.n138 a_n2298_n2088# 0.012691f
C232 source.n139 a_n2298_n2088# 0.029998f
C233 source.n140 a_n2298_n2088# 0.013438f
C234 source.n141 a_n2298_n2088# 0.023618f
C235 source.n142 a_n2298_n2088# 0.012691f
C236 source.n143 a_n2298_n2088# 0.029998f
C237 source.n144 a_n2298_n2088# 0.013438f
C238 source.n145 a_n2298_n2088# 0.101069f
C239 source.t17 a_n2298_n2088# 0.048893f
C240 source.n146 a_n2298_n2088# 0.022498f
C241 source.n147 a_n2298_n2088# 0.017719f
C242 source.n148 a_n2298_n2088# 0.012691f
C243 source.n149 a_n2298_n2088# 0.561971f
C244 source.n150 a_n2298_n2088# 0.023618f
C245 source.n151 a_n2298_n2088# 0.012691f
C246 source.n152 a_n2298_n2088# 0.013438f
C247 source.n153 a_n2298_n2088# 0.029998f
C248 source.n154 a_n2298_n2088# 0.029998f
C249 source.n155 a_n2298_n2088# 0.013438f
C250 source.n156 a_n2298_n2088# 0.012691f
C251 source.n157 a_n2298_n2088# 0.023618f
C252 source.n158 a_n2298_n2088# 0.023618f
C253 source.n159 a_n2298_n2088# 0.012691f
C254 source.n160 a_n2298_n2088# 0.013438f
C255 source.n161 a_n2298_n2088# 0.029998f
C256 source.n162 a_n2298_n2088# 0.06494f
C257 source.n163 a_n2298_n2088# 0.013438f
C258 source.n164 a_n2298_n2088# 0.012691f
C259 source.n165 a_n2298_n2088# 0.054592f
C260 source.n166 a_n2298_n2088# 0.036337f
C261 source.n167 a_n2298_n2088# 0.941744f
C262 source.t19 a_n2298_n2088# 0.111983f
C263 source.t10 a_n2298_n2088# 0.111983f
C264 source.n168 a_n2298_n2088# 0.872125f
C265 source.n169 a_n2298_n2088# 0.369673f
C266 source.t20 a_n2298_n2088# 0.111983f
C267 source.t21 a_n2298_n2088# 0.111983f
C268 source.n170 a_n2298_n2088# 0.872125f
C269 source.n171 a_n2298_n2088# 0.369673f
C270 source.n172 a_n2298_n2088# 0.033197f
C271 source.n173 a_n2298_n2088# 0.023618f
C272 source.n174 a_n2298_n2088# 0.012691f
C273 source.n175 a_n2298_n2088# 0.029998f
C274 source.n176 a_n2298_n2088# 0.013438f
C275 source.n177 a_n2298_n2088# 0.023618f
C276 source.n178 a_n2298_n2088# 0.012691f
C277 source.n179 a_n2298_n2088# 0.029998f
C278 source.n180 a_n2298_n2088# 0.013438f
C279 source.n181 a_n2298_n2088# 0.101069f
C280 source.t18 a_n2298_n2088# 0.048893f
C281 source.n182 a_n2298_n2088# 0.022498f
C282 source.n183 a_n2298_n2088# 0.017719f
C283 source.n184 a_n2298_n2088# 0.012691f
C284 source.n185 a_n2298_n2088# 0.561971f
C285 source.n186 a_n2298_n2088# 0.023618f
C286 source.n187 a_n2298_n2088# 0.012691f
C287 source.n188 a_n2298_n2088# 0.013438f
C288 source.n189 a_n2298_n2088# 0.029998f
C289 source.n190 a_n2298_n2088# 0.029998f
C290 source.n191 a_n2298_n2088# 0.013438f
C291 source.n192 a_n2298_n2088# 0.012691f
C292 source.n193 a_n2298_n2088# 0.023618f
C293 source.n194 a_n2298_n2088# 0.023618f
C294 source.n195 a_n2298_n2088# 0.012691f
C295 source.n196 a_n2298_n2088# 0.013438f
C296 source.n197 a_n2298_n2088# 0.029998f
C297 source.n198 a_n2298_n2088# 0.06494f
C298 source.n199 a_n2298_n2088# 0.013438f
C299 source.n200 a_n2298_n2088# 0.012691f
C300 source.n201 a_n2298_n2088# 0.054592f
C301 source.n202 a_n2298_n2088# 0.036337f
C302 source.n203 a_n2298_n2088# 0.130062f
C303 source.n204 a_n2298_n2088# 0.033197f
C304 source.n205 a_n2298_n2088# 0.023618f
C305 source.n206 a_n2298_n2088# 0.012691f
C306 source.n207 a_n2298_n2088# 0.029998f
C307 source.n208 a_n2298_n2088# 0.013438f
C308 source.n209 a_n2298_n2088# 0.023618f
C309 source.n210 a_n2298_n2088# 0.012691f
C310 source.n211 a_n2298_n2088# 0.029998f
C311 source.n212 a_n2298_n2088# 0.013438f
C312 source.n213 a_n2298_n2088# 0.101069f
C313 source.t8 a_n2298_n2088# 0.048893f
C314 source.n214 a_n2298_n2088# 0.022498f
C315 source.n215 a_n2298_n2088# 0.017719f
C316 source.n216 a_n2298_n2088# 0.012691f
C317 source.n217 a_n2298_n2088# 0.561971f
C318 source.n218 a_n2298_n2088# 0.023618f
C319 source.n219 a_n2298_n2088# 0.012691f
C320 source.n220 a_n2298_n2088# 0.013438f
C321 source.n221 a_n2298_n2088# 0.029998f
C322 source.n222 a_n2298_n2088# 0.029998f
C323 source.n223 a_n2298_n2088# 0.013438f
C324 source.n224 a_n2298_n2088# 0.012691f
C325 source.n225 a_n2298_n2088# 0.023618f
C326 source.n226 a_n2298_n2088# 0.023618f
C327 source.n227 a_n2298_n2088# 0.012691f
C328 source.n228 a_n2298_n2088# 0.013438f
C329 source.n229 a_n2298_n2088# 0.029998f
C330 source.n230 a_n2298_n2088# 0.06494f
C331 source.n231 a_n2298_n2088# 0.013438f
C332 source.n232 a_n2298_n2088# 0.012691f
C333 source.n233 a_n2298_n2088# 0.054592f
C334 source.n234 a_n2298_n2088# 0.036337f
C335 source.n235 a_n2298_n2088# 0.130062f
C336 source.t22 a_n2298_n2088# 0.111983f
C337 source.t9 a_n2298_n2088# 0.111983f
C338 source.n236 a_n2298_n2088# 0.872125f
C339 source.n237 a_n2298_n2088# 0.369673f
C340 source.t1 a_n2298_n2088# 0.111983f
C341 source.t6 a_n2298_n2088# 0.111983f
C342 source.n238 a_n2298_n2088# 0.872125f
C343 source.n239 a_n2298_n2088# 0.369673f
C344 source.n240 a_n2298_n2088# 0.033197f
C345 source.n241 a_n2298_n2088# 0.023618f
C346 source.n242 a_n2298_n2088# 0.012691f
C347 source.n243 a_n2298_n2088# 0.029998f
C348 source.n244 a_n2298_n2088# 0.013438f
C349 source.n245 a_n2298_n2088# 0.023618f
C350 source.n246 a_n2298_n2088# 0.012691f
C351 source.n247 a_n2298_n2088# 0.029998f
C352 source.n248 a_n2298_n2088# 0.013438f
C353 source.n249 a_n2298_n2088# 0.101069f
C354 source.t23 a_n2298_n2088# 0.048893f
C355 source.n250 a_n2298_n2088# 0.022498f
C356 source.n251 a_n2298_n2088# 0.017719f
C357 source.n252 a_n2298_n2088# 0.012691f
C358 source.n253 a_n2298_n2088# 0.561971f
C359 source.n254 a_n2298_n2088# 0.023618f
C360 source.n255 a_n2298_n2088# 0.012691f
C361 source.n256 a_n2298_n2088# 0.013438f
C362 source.n257 a_n2298_n2088# 0.029998f
C363 source.n258 a_n2298_n2088# 0.029998f
C364 source.n259 a_n2298_n2088# 0.013438f
C365 source.n260 a_n2298_n2088# 0.012691f
C366 source.n261 a_n2298_n2088# 0.023618f
C367 source.n262 a_n2298_n2088# 0.023618f
C368 source.n263 a_n2298_n2088# 0.012691f
C369 source.n264 a_n2298_n2088# 0.013438f
C370 source.n265 a_n2298_n2088# 0.029998f
C371 source.n266 a_n2298_n2088# 0.06494f
C372 source.n267 a_n2298_n2088# 0.013438f
C373 source.n268 a_n2298_n2088# 0.012691f
C374 source.n269 a_n2298_n2088# 0.054592f
C375 source.n270 a_n2298_n2088# 0.036337f
C376 source.n271 a_n2298_n2088# 0.289237f
C377 source.n272 a_n2298_n2088# 0.982857f
C378 drain_left.t5 a_n2298_n2088# 0.126027f
C379 drain_left.t4 a_n2298_n2088# 0.126027f
C380 drain_left.n0 a_n2298_n2088# 1.05632f
C381 drain_left.t9 a_n2298_n2088# 0.126027f
C382 drain_left.t10 a_n2298_n2088# 0.126027f
C383 drain_left.n1 a_n2298_n2088# 1.05107f
C384 drain_left.t3 a_n2298_n2088# 0.126027f
C385 drain_left.t2 a_n2298_n2088# 0.126027f
C386 drain_left.n2 a_n2298_n2088# 1.05632f
C387 drain_left.n3 a_n2298_n2088# 2.17713f
C388 drain_left.t6 a_n2298_n2088# 0.126027f
C389 drain_left.t1 a_n2298_n2088# 0.126027f
C390 drain_left.n4 a_n2298_n2088# 1.05669f
C391 drain_left.t0 a_n2298_n2088# 0.126027f
C392 drain_left.t8 a_n2298_n2088# 0.126027f
C393 drain_left.n5 a_n2298_n2088# 1.05107f
C394 drain_left.n6 a_n2298_n2088# 0.770273f
C395 drain_left.t11 a_n2298_n2088# 0.126027f
C396 drain_left.t7 a_n2298_n2088# 0.126027f
C397 drain_left.n7 a_n2298_n2088# 1.05107f
C398 drain_left.n8 a_n2298_n2088# 0.620942f
C399 plus.n0 a_n2298_n2088# 0.041876f
C400 plus.t5 a_n2298_n2088# 0.583027f
C401 plus.t8 a_n2298_n2088# 0.583027f
C402 plus.n1 a_n2298_n2088# 0.041876f
C403 plus.t6 a_n2298_n2088# 0.583027f
C404 plus.n2 a_n2298_n2088# 0.277279f
C405 plus.n3 a_n2298_n2088# 0.192243f
C406 plus.t7 a_n2298_n2088# 0.583027f
C407 plus.t9 a_n2298_n2088# 0.583027f
C408 plus.t10 a_n2298_n2088# 0.605841f
C409 plus.n4 a_n2298_n2088# 0.249245f
C410 plus.n5 a_n2298_n2088# 0.268845f
C411 plus.n6 a_n2298_n2088# 0.009503f
C412 plus.n7 a_n2298_n2088# 0.277279f
C413 plus.n8 a_n2298_n2088# 0.06975f
C414 plus.n9 a_n2298_n2088# 0.06975f
C415 plus.n10 a_n2298_n2088# 0.055878f
C416 plus.n11 a_n2298_n2088# 0.009503f
C417 plus.n12 a_n2298_n2088# 0.265582f
C418 plus.n13 a_n2298_n2088# 0.009503f
C419 plus.n14 a_n2298_n2088# 0.264937f
C420 plus.n15 a_n2298_n2088# 0.379404f
C421 plus.n16 a_n2298_n2088# 0.041876f
C422 plus.t4 a_n2298_n2088# 0.583027f
C423 plus.n17 a_n2298_n2088# 0.041876f
C424 plus.t2 a_n2298_n2088# 0.583027f
C425 plus.t11 a_n2298_n2088# 0.583027f
C426 plus.n18 a_n2298_n2088# 0.277279f
C427 plus.n19 a_n2298_n2088# 0.192243f
C428 plus.t1 a_n2298_n2088# 0.583027f
C429 plus.t3 a_n2298_n2088# 0.605841f
C430 plus.n20 a_n2298_n2088# 0.249245f
C431 plus.t0 a_n2298_n2088# 0.583027f
C432 plus.n21 a_n2298_n2088# 0.268845f
C433 plus.n22 a_n2298_n2088# 0.009503f
C434 plus.n23 a_n2298_n2088# 0.277279f
C435 plus.n24 a_n2298_n2088# 0.06975f
C436 plus.n25 a_n2298_n2088# 0.06975f
C437 plus.n26 a_n2298_n2088# 0.055878f
C438 plus.n27 a_n2298_n2088# 0.009503f
C439 plus.n28 a_n2298_n2088# 0.265582f
C440 plus.n29 a_n2298_n2088# 0.009503f
C441 plus.n30 a_n2298_n2088# 0.264937f
C442 plus.n31 a_n2298_n2088# 1.18985f
.ends

