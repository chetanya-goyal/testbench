* NGSPICE file created from diffpair328.ext - technology: sky130A

.subckt diffpair328 minus drain_right drain_left source plus
X0 a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X1 drain_left.t19 plus.t0 source.t24 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 drain_left.t18 plus.t1 source.t26 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X3 source.t36 plus.t2 drain_left.t17 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X4 source.t30 plus.t3 drain_left.t16 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X5 drain_left.t15 plus.t4 source.t32 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X6 source.t1 minus.t0 drain_right.t19 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X8 source.t4 minus.t1 drain_right.t18 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 drain_left.t14 plus.t5 source.t20 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X10 drain_right.t17 minus.t2 source.t8 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X11 drain_left.t13 plus.t6 source.t33 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X12 drain_right.t16 minus.t3 source.t10 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X13 source.t14 minus.t4 drain_right.t15 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X14 drain_right.t14 minus.t5 source.t15 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X15 source.t25 plus.t7 drain_left.t12 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X16 a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X17 drain_right.t13 minus.t6 source.t38 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X18 drain_right.t12 minus.t7 source.t39 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t3 minus.t8 drain_right.t11 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X20 source.t0 minus.t9 drain_right.t10 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X21 drain_right.t9 minus.t10 source.t2 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X22 source.t13 minus.t11 drain_right.t8 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X23 drain_left.t11 plus.t8 source.t35 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X24 source.t27 plus.t9 drain_left.t10 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X25 drain_right.t7 minus.t12 source.t11 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X26 drain_right.t6 minus.t13 source.t7 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X27 source.t9 minus.t14 drain_right.t5 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X28 drain_left.t9 plus.t10 source.t23 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X29 source.t12 minus.t15 drain_right.t4 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X30 drain_right.t3 minus.t16 source.t5 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X31 source.t19 plus.t11 drain_left.t8 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X32 drain_left.t7 plus.t12 source.t28 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X33 source.t37 plus.t13 drain_left.t6 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X34 source.t34 plus.t14 drain_left.t5 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X35 drain_right.t2 minus.t17 source.t6 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X36 source.t17 minus.t18 drain_right.t1 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X37 source.t31 plus.t15 drain_left.t4 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X38 drain_left.t3 plus.t16 source.t21 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X39 drain_left.t2 plus.t17 source.t29 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X40 source.t16 minus.t19 drain_right.t0 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X41 source.t22 plus.t18 drain_left.t1 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X42 a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X43 source.t18 plus.t19 drain_left.t0 a_n2146_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n6 plus.t9 1716.94
R1 plus.n27 plus.t12 1716.94
R2 plus.n36 plus.t5 1716.94
R3 plus.n56 plus.t11 1716.94
R4 plus.n5 plus.t17 1654.87
R5 plus.n9 plus.t14 1654.87
R6 plus.n3 plus.t10 1654.87
R7 plus.n15 plus.t19 1654.87
R8 plus.n17 plus.t16 1654.87
R9 plus.n18 plus.t13 1654.87
R10 plus.n24 plus.t8 1654.87
R11 plus.n26 plus.t15 1654.87
R12 plus.n35 plus.t7 1654.87
R13 plus.n39 plus.t0 1654.87
R14 plus.n33 plus.t3 1654.87
R15 plus.n45 plus.t6 1654.87
R16 plus.n47 plus.t18 1654.87
R17 plus.n32 plus.t1 1654.87
R18 plus.n53 plus.t2 1654.87
R19 plus.n55 plus.t4 1654.87
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 69.3793
R47 plus.n19 plus.n18 69.3793
R48 plus.n48 plus.n32 69.3793
R49 plus.n44 plus.n33 69.3793
R50 plus.n9 plus.n8 54.7732
R51 plus.n25 plus.n24 54.7732
R52 plus.n54 plus.n53 54.7732
R53 plus.n39 plus.n38 54.7732
R54 plus.n16 plus.n15 47.4702
R55 plus.n17 plus.n16 47.4702
R56 plus.n47 plus.n46 47.4702
R57 plus.n46 plus.n45 47.4702
R58 plus.n8 plus.n5 40.1672
R59 plus.n26 plus.n25 40.1672
R60 plus.n55 plus.n54 40.1672
R61 plus.n38 plus.n35 40.1672
R62 plus.n6 plus.n5 32.8641
R63 plus.n27 plus.n26 32.8641
R64 plus.n56 plus.n55 32.8641
R65 plus.n36 plus.n35 32.8641
R66 plus plus.n57 30.0558
R67 plus.n15 plus.n14 25.5611
R68 plus.n19 plus.n17 25.5611
R69 plus.n48 plus.n47 25.5611
R70 plus.n45 plus.n44 25.5611
R71 plus.n10 plus.n9 18.2581
R72 plus.n24 plus.n23 18.2581
R73 plus.n53 plus.n52 18.2581
R74 plus.n40 plus.n39 18.2581
R75 plus plus.n28 11.0687
R76 plus.n11 plus.n3 3.65202
R77 plus.n18 plus.n1 3.65202
R78 plus.n32 plus.n30 3.65202
R79 plus.n41 plus.n33 3.65202
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n9 source.t27 52.1921
R99 source.n10 source.t38 52.1921
R100 source.n19 source.t17 52.1921
R101 source.n39 source.t15 52.1919
R102 source.n30 source.t16 52.1919
R103 source.n29 source.t20 52.1919
R104 source.n20 source.t19 52.1919
R105 source.n0 source.t28 52.1919
R106 source.n2 source.n1 48.8588
R107 source.n4 source.n3 48.8588
R108 source.n6 source.n5 48.8588
R109 source.n8 source.n7 48.8588
R110 source.n12 source.n11 48.8588
R111 source.n14 source.n13 48.8588
R112 source.n16 source.n15 48.8588
R113 source.n18 source.n17 48.8588
R114 source.n38 source.n37 48.8586
R115 source.n36 source.n35 48.8586
R116 source.n34 source.n33 48.8586
R117 source.n32 source.n31 48.8586
R118 source.n28 source.n27 48.8586
R119 source.n26 source.n25 48.8586
R120 source.n24 source.n23 48.8586
R121 source.n22 source.n21 48.8586
R122 source.n20 source.n19 19.5753
R123 source.n40 source.n0 14.0322
R124 source.n40 source.n39 5.5436
R125 source.n37 source.t6 3.33383
R126 source.n37 source.t4 3.33383
R127 source.n35 source.t10 3.33383
R128 source.n35 source.t13 3.33383
R129 source.n33 source.t5 3.33383
R130 source.n33 source.t1 3.33383
R131 source.n31 source.t8 3.33383
R132 source.n31 source.t3 3.33383
R133 source.n27 source.t24 3.33383
R134 source.n27 source.t25 3.33383
R135 source.n25 source.t33 3.33383
R136 source.n25 source.t30 3.33383
R137 source.n23 source.t26 3.33383
R138 source.n23 source.t22 3.33383
R139 source.n21 source.t32 3.33383
R140 source.n21 source.t36 3.33383
R141 source.n1 source.t35 3.33383
R142 source.n1 source.t31 3.33383
R143 source.n3 source.t21 3.33383
R144 source.n3 source.t37 3.33383
R145 source.n5 source.t23 3.33383
R146 source.n5 source.t18 3.33383
R147 source.n7 source.t29 3.33383
R148 source.n7 source.t34 3.33383
R149 source.n11 source.t11 3.33383
R150 source.n11 source.t14 3.33383
R151 source.n13 source.t39 3.33383
R152 source.n13 source.t0 3.33383
R153 source.n15 source.t7 3.33383
R154 source.n15 source.t12 3.33383
R155 source.n17 source.t2 3.33383
R156 source.n17 source.t9 3.33383
R157 source.n19 source.n18 0.560845
R158 source.n18 source.n16 0.560845
R159 source.n16 source.n14 0.560845
R160 source.n14 source.n12 0.560845
R161 source.n12 source.n10 0.560845
R162 source.n9 source.n8 0.560845
R163 source.n8 source.n6 0.560845
R164 source.n6 source.n4 0.560845
R165 source.n4 source.n2 0.560845
R166 source.n2 source.n0 0.560845
R167 source.n22 source.n20 0.560845
R168 source.n24 source.n22 0.560845
R169 source.n26 source.n24 0.560845
R170 source.n28 source.n26 0.560845
R171 source.n29 source.n28 0.560845
R172 source.n32 source.n30 0.560845
R173 source.n34 source.n32 0.560845
R174 source.n36 source.n34 0.560845
R175 source.n38 source.n36 0.560845
R176 source.n39 source.n38 0.560845
R177 source.n10 source.n9 0.470328
R178 source.n30 source.n29 0.470328
R179 source source.n40 0.188
R180 drain_left.n10 drain_left.n8 66.0979
R181 drain_left.n6 drain_left.n4 66.0977
R182 drain_left.n2 drain_left.n0 66.0977
R183 drain_left.n14 drain_left.n13 65.5376
R184 drain_left.n12 drain_left.n11 65.5376
R185 drain_left.n10 drain_left.n9 65.5376
R186 drain_left.n16 drain_left.n15 65.5374
R187 drain_left.n7 drain_left.n3 65.5373
R188 drain_left.n6 drain_left.n5 65.5373
R189 drain_left.n2 drain_left.n1 65.5373
R190 drain_left drain_left.n7 29.5771
R191 drain_left drain_left.n16 6.21356
R192 drain_left.n3 drain_left.t1 3.33383
R193 drain_left.n3 drain_left.t13 3.33383
R194 drain_left.n4 drain_left.t12 3.33383
R195 drain_left.n4 drain_left.t14 3.33383
R196 drain_left.n5 drain_left.t16 3.33383
R197 drain_left.n5 drain_left.t19 3.33383
R198 drain_left.n1 drain_left.t17 3.33383
R199 drain_left.n1 drain_left.t18 3.33383
R200 drain_left.n0 drain_left.t8 3.33383
R201 drain_left.n0 drain_left.t15 3.33383
R202 drain_left.n15 drain_left.t4 3.33383
R203 drain_left.n15 drain_left.t7 3.33383
R204 drain_left.n13 drain_left.t6 3.33383
R205 drain_left.n13 drain_left.t11 3.33383
R206 drain_left.n11 drain_left.t0 3.33383
R207 drain_left.n11 drain_left.t3 3.33383
R208 drain_left.n9 drain_left.t5 3.33383
R209 drain_left.n9 drain_left.t9 3.33383
R210 drain_left.n8 drain_left.t10 3.33383
R211 drain_left.n8 drain_left.t2 3.33383
R212 drain_left.n12 drain_left.n10 0.560845
R213 drain_left.n14 drain_left.n12 0.560845
R214 drain_left.n16 drain_left.n14 0.560845
R215 drain_left.n7 drain_left.n6 0.505499
R216 drain_left.n7 drain_left.n2 0.505499
R217 minus.n27 minus.t18 1716.94
R218 minus.n7 minus.t6 1716.94
R219 minus.n56 minus.t5 1716.94
R220 minus.n35 minus.t19 1716.94
R221 minus.n26 minus.t10 1654.87
R222 minus.n24 minus.t14 1654.87
R223 minus.n3 minus.t13 1654.87
R224 minus.n18 minus.t15 1654.87
R225 minus.n16 minus.t7 1654.87
R226 minus.n4 minus.t9 1654.87
R227 minus.n10 minus.t12 1654.87
R228 minus.n6 minus.t4 1654.87
R229 minus.n55 minus.t1 1654.87
R230 minus.n53 minus.t17 1654.87
R231 minus.n47 minus.t11 1654.87
R232 minus.n46 minus.t3 1654.87
R233 minus.n44 minus.t0 1654.87
R234 minus.n32 minus.t16 1654.87
R235 minus.n38 minus.t8 1654.87
R236 minus.n34 minus.t2 1654.87
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 69.3793
R264 minus.n15 minus.n4 69.3793
R265 minus.n43 minus.n32 69.3793
R266 minus.n48 minus.n47 69.3793
R267 minus.n25 minus.n24 54.7732
R268 minus.n10 minus.n9 54.7732
R269 minus.n38 minus.n37 54.7732
R270 minus.n54 minus.n53 54.7732
R271 minus.n18 minus.n17 47.4702
R272 minus.n17 minus.n16 47.4702
R273 minus.n45 minus.n44 47.4702
R274 minus.n46 minus.n45 47.4702
R275 minus.n26 minus.n25 40.1672
R276 minus.n9 minus.n6 40.1672
R277 minus.n37 minus.n34 40.1672
R278 minus.n55 minus.n54 40.1672
R279 minus.n58 minus.n28 35.0384
R280 minus.n27 minus.n26 32.8641
R281 minus.n7 minus.n6 32.8641
R282 minus.n35 minus.n34 32.8641
R283 minus.n56 minus.n55 32.8641
R284 minus.n19 minus.n18 25.5611
R285 minus.n16 minus.n15 25.5611
R286 minus.n44 minus.n43 25.5611
R287 minus.n48 minus.n46 25.5611
R288 minus.n24 minus.n23 18.2581
R289 minus.n11 minus.n10 18.2581
R290 minus.n39 minus.n38 18.2581
R291 minus.n53 minus.n52 18.2581
R292 minus.n58 minus.n57 6.56111
R293 minus.n3 minus.n1 3.65202
R294 minus.n12 minus.n4 3.65202
R295 minus.n40 minus.n32 3.65202
R296 minus.n47 minus.n30 3.65202
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 66.0978
R317 drain_right.n6 drain_right.n4 66.0977
R318 drain_right.n2 drain_right.n0 66.0977
R319 drain_right.n10 drain_right.n9 65.5376
R320 drain_right.n12 drain_right.n11 65.5376
R321 drain_right.n14 drain_right.n13 65.5376
R322 drain_right.n16 drain_right.n15 65.5376
R323 drain_right.n7 drain_right.n3 65.5373
R324 drain_right.n6 drain_right.n5 65.5373
R325 drain_right.n2 drain_right.n1 65.5373
R326 drain_right drain_right.n7 29.0239
R327 drain_right drain_right.n16 6.21356
R328 drain_right.n3 drain_right.t19 3.33383
R329 drain_right.n3 drain_right.t16 3.33383
R330 drain_right.n4 drain_right.t18 3.33383
R331 drain_right.n4 drain_right.t14 3.33383
R332 drain_right.n5 drain_right.t8 3.33383
R333 drain_right.n5 drain_right.t2 3.33383
R334 drain_right.n1 drain_right.t11 3.33383
R335 drain_right.n1 drain_right.t3 3.33383
R336 drain_right.n0 drain_right.t0 3.33383
R337 drain_right.n0 drain_right.t17 3.33383
R338 drain_right.n8 drain_right.t15 3.33383
R339 drain_right.n8 drain_right.t13 3.33383
R340 drain_right.n9 drain_right.t10 3.33383
R341 drain_right.n9 drain_right.t7 3.33383
R342 drain_right.n11 drain_right.t4 3.33383
R343 drain_right.n11 drain_right.t12 3.33383
R344 drain_right.n13 drain_right.t5 3.33383
R345 drain_right.n13 drain_right.t6 3.33383
R346 drain_right.n15 drain_right.t1 3.33383
R347 drain_right.n15 drain_right.t9 3.33383
R348 drain_right.n16 drain_right.n14 0.560845
R349 drain_right.n14 drain_right.n12 0.560845
R350 drain_right.n12 drain_right.n10 0.560845
R351 drain_right.n7 drain_right.n6 0.505499
R352 drain_right.n7 drain_right.n2 0.505499
C0 drain_right plus 0.364841f
C1 drain_right minus 3.31904f
C2 drain_right source 29.545301f
C3 drain_left plus 3.52973f
C4 drain_left minus 0.171338f
C5 plus minus 5.25731f
C6 drain_left source 29.5448f
C7 plus source 3.01175f
C8 minus source 2.99771f
C9 drain_left drain_right 1.13563f
C10 drain_right a_n2146_n2688# 5.87101f
C11 drain_left a_n2146_n2688# 6.1866f
C12 source a_n2146_n2688# 7.297064f
C13 minus a_n2146_n2688# 7.725148f
C14 plus a_n2146_n2688# 9.69234f
C15 drain_right.t0 a_n2146_n2688# 0.303215f
C16 drain_right.t17 a_n2146_n2688# 0.303215f
C17 drain_right.n0 a_n2146_n2688# 1.95945f
C18 drain_right.t11 a_n2146_n2688# 0.303215f
C19 drain_right.t3 a_n2146_n2688# 0.303215f
C20 drain_right.n1 a_n2146_n2688# 1.95658f
C21 drain_right.n2 a_n2146_n2688# 0.658742f
C22 drain_right.t19 a_n2146_n2688# 0.303215f
C23 drain_right.t16 a_n2146_n2688# 0.303215f
C24 drain_right.n3 a_n2146_n2688# 1.95658f
C25 drain_right.t18 a_n2146_n2688# 0.303215f
C26 drain_right.t14 a_n2146_n2688# 0.303215f
C27 drain_right.n4 a_n2146_n2688# 1.95945f
C28 drain_right.t8 a_n2146_n2688# 0.303215f
C29 drain_right.t2 a_n2146_n2688# 0.303215f
C30 drain_right.n5 a_n2146_n2688# 1.95658f
C31 drain_right.n6 a_n2146_n2688# 0.658742f
C32 drain_right.n7 a_n2146_n2688# 1.49839f
C33 drain_right.t15 a_n2146_n2688# 0.303215f
C34 drain_right.t13 a_n2146_n2688# 0.303215f
C35 drain_right.n8 a_n2146_n2688# 1.95945f
C36 drain_right.t10 a_n2146_n2688# 0.303215f
C37 drain_right.t7 a_n2146_n2688# 0.303215f
C38 drain_right.n9 a_n2146_n2688# 1.95658f
C39 drain_right.n10 a_n2146_n2688# 0.662469f
C40 drain_right.t4 a_n2146_n2688# 0.303215f
C41 drain_right.t12 a_n2146_n2688# 0.303215f
C42 drain_right.n11 a_n2146_n2688# 1.95658f
C43 drain_right.n12 a_n2146_n2688# 0.326998f
C44 drain_right.t5 a_n2146_n2688# 0.303215f
C45 drain_right.t6 a_n2146_n2688# 0.303215f
C46 drain_right.n13 a_n2146_n2688# 1.95658f
C47 drain_right.n14 a_n2146_n2688# 0.326998f
C48 drain_right.t1 a_n2146_n2688# 0.303215f
C49 drain_right.t9 a_n2146_n2688# 0.303215f
C50 drain_right.n15 a_n2146_n2688# 1.95658f
C51 drain_right.n16 a_n2146_n2688# 0.561983f
C52 minus.n0 a_n2146_n2688# 0.05197f
C53 minus.t18 a_n2146_n2688# 0.202183f
C54 minus.t10 a_n2146_n2688# 0.198805f
C55 minus.t14 a_n2146_n2688# 0.198805f
C56 minus.n1 a_n2146_n2688# 0.018041f
C57 minus.n2 a_n2146_n2688# 0.05197f
C58 minus.t13 a_n2146_n2688# 0.198805f
C59 minus.n3 a_n2146_n2688# 0.091028f
C60 minus.t15 a_n2146_n2688# 0.198805f
C61 minus.t7 a_n2146_n2688# 0.198805f
C62 minus.t9 a_n2146_n2688# 0.198805f
C63 minus.n4 a_n2146_n2688# 0.091028f
C64 minus.n5 a_n2146_n2688# 0.05197f
C65 minus.t12 a_n2146_n2688# 0.198805f
C66 minus.t4 a_n2146_n2688# 0.198805f
C67 minus.n6 a_n2146_n2688# 0.091028f
C68 minus.t6 a_n2146_n2688# 0.202183f
C69 minus.n7 a_n2146_n2688# 0.112179f
C70 minus.n8 a_n2146_n2688# 0.119881f
C71 minus.n9 a_n2146_n2688# 0.022046f
C72 minus.n10 a_n2146_n2688# 0.091028f
C73 minus.n11 a_n2146_n2688# 0.021245f
C74 minus.n12 a_n2146_n2688# 0.018041f
C75 minus.n13 a_n2146_n2688# 0.05197f
C76 minus.n14 a_n2146_n2688# 0.05197f
C77 minus.n15 a_n2146_n2688# 0.022046f
C78 minus.n16 a_n2146_n2688# 0.091028f
C79 minus.n17 a_n2146_n2688# 0.022046f
C80 minus.n18 a_n2146_n2688# 0.091028f
C81 minus.n19 a_n2146_n2688# 0.022046f
C82 minus.n20 a_n2146_n2688# 0.05197f
C83 minus.n21 a_n2146_n2688# 0.05197f
C84 minus.n22 a_n2146_n2688# 0.05197f
C85 minus.n23 a_n2146_n2688# 0.021245f
C86 minus.n24 a_n2146_n2688# 0.091028f
C87 minus.n25 a_n2146_n2688# 0.022046f
C88 minus.n26 a_n2146_n2688# 0.091028f
C89 minus.n27 a_n2146_n2688# 0.1121f
C90 minus.n28 a_n2146_n2688# 1.74774f
C91 minus.n29 a_n2146_n2688# 0.05197f
C92 minus.t1 a_n2146_n2688# 0.198805f
C93 minus.t17 a_n2146_n2688# 0.198805f
C94 minus.n30 a_n2146_n2688# 0.018041f
C95 minus.n31 a_n2146_n2688# 0.05197f
C96 minus.t3 a_n2146_n2688# 0.198805f
C97 minus.t0 a_n2146_n2688# 0.198805f
C98 minus.t16 a_n2146_n2688# 0.198805f
C99 minus.n32 a_n2146_n2688# 0.091028f
C100 minus.n33 a_n2146_n2688# 0.05197f
C101 minus.t8 a_n2146_n2688# 0.198805f
C102 minus.t2 a_n2146_n2688# 0.198805f
C103 minus.n34 a_n2146_n2688# 0.091028f
C104 minus.t19 a_n2146_n2688# 0.202183f
C105 minus.n35 a_n2146_n2688# 0.112179f
C106 minus.n36 a_n2146_n2688# 0.119881f
C107 minus.n37 a_n2146_n2688# 0.022046f
C108 minus.n38 a_n2146_n2688# 0.091028f
C109 minus.n39 a_n2146_n2688# 0.021245f
C110 minus.n40 a_n2146_n2688# 0.018041f
C111 minus.n41 a_n2146_n2688# 0.05197f
C112 minus.n42 a_n2146_n2688# 0.05197f
C113 minus.n43 a_n2146_n2688# 0.022046f
C114 minus.n44 a_n2146_n2688# 0.091028f
C115 minus.n45 a_n2146_n2688# 0.022046f
C116 minus.n46 a_n2146_n2688# 0.091028f
C117 minus.t11 a_n2146_n2688# 0.198805f
C118 minus.n47 a_n2146_n2688# 0.091028f
C119 minus.n48 a_n2146_n2688# 0.022046f
C120 minus.n49 a_n2146_n2688# 0.05197f
C121 minus.n50 a_n2146_n2688# 0.05197f
C122 minus.n51 a_n2146_n2688# 0.05197f
C123 minus.n52 a_n2146_n2688# 0.021245f
C124 minus.n53 a_n2146_n2688# 0.091028f
C125 minus.n54 a_n2146_n2688# 0.022046f
C126 minus.n55 a_n2146_n2688# 0.091028f
C127 minus.t5 a_n2146_n2688# 0.202183f
C128 minus.n56 a_n2146_n2688# 0.1121f
C129 minus.n57 a_n2146_n2688# 0.347228f
C130 minus.n58 a_n2146_n2688# 2.12739f
C131 drain_left.t8 a_n2146_n2688# 0.304043f
C132 drain_left.t15 a_n2146_n2688# 0.304043f
C133 drain_left.n0 a_n2146_n2688# 1.9648f
C134 drain_left.t17 a_n2146_n2688# 0.304043f
C135 drain_left.t18 a_n2146_n2688# 0.304043f
C136 drain_left.n1 a_n2146_n2688# 1.96193f
C137 drain_left.n2 a_n2146_n2688# 0.660542f
C138 drain_left.t1 a_n2146_n2688# 0.304043f
C139 drain_left.t13 a_n2146_n2688# 0.304043f
C140 drain_left.n3 a_n2146_n2688# 1.96193f
C141 drain_left.t12 a_n2146_n2688# 0.304043f
C142 drain_left.t14 a_n2146_n2688# 0.304043f
C143 drain_left.n4 a_n2146_n2688# 1.9648f
C144 drain_left.t16 a_n2146_n2688# 0.304043f
C145 drain_left.t19 a_n2146_n2688# 0.304043f
C146 drain_left.n5 a_n2146_n2688# 1.96193f
C147 drain_left.n6 a_n2146_n2688# 0.660542f
C148 drain_left.n7 a_n2146_n2688# 1.56025f
C149 drain_left.t10 a_n2146_n2688# 0.304043f
C150 drain_left.t2 a_n2146_n2688# 0.304043f
C151 drain_left.n8 a_n2146_n2688# 1.96481f
C152 drain_left.t5 a_n2146_n2688# 0.304043f
C153 drain_left.t9 a_n2146_n2688# 0.304043f
C154 drain_left.n9 a_n2146_n2688# 1.96193f
C155 drain_left.n10 a_n2146_n2688# 0.664271f
C156 drain_left.t0 a_n2146_n2688# 0.304043f
C157 drain_left.t3 a_n2146_n2688# 0.304043f
C158 drain_left.n11 a_n2146_n2688# 1.96193f
C159 drain_left.n12 a_n2146_n2688# 0.327892f
C160 drain_left.t6 a_n2146_n2688# 0.304043f
C161 drain_left.t11 a_n2146_n2688# 0.304043f
C162 drain_left.n13 a_n2146_n2688# 1.96193f
C163 drain_left.n14 a_n2146_n2688# 0.327892f
C164 drain_left.t4 a_n2146_n2688# 0.304043f
C165 drain_left.t7 a_n2146_n2688# 0.304043f
C166 drain_left.n15 a_n2146_n2688# 1.96192f
C167 drain_left.n16 a_n2146_n2688# 0.563526f
C168 source.t28 a_n2146_n2688# 2.04763f
C169 source.n0 a_n2146_n2688# 1.14221f
C170 source.t35 a_n2146_n2688# 0.270934f
C171 source.t31 a_n2146_n2688# 0.270934f
C172 source.n1 a_n2146_n2688# 1.68117f
C173 source.n2 a_n2146_n2688# 0.325128f
C174 source.t21 a_n2146_n2688# 0.270934f
C175 source.t37 a_n2146_n2688# 0.270934f
C176 source.n3 a_n2146_n2688# 1.68117f
C177 source.n4 a_n2146_n2688# 0.325128f
C178 source.t23 a_n2146_n2688# 0.270934f
C179 source.t18 a_n2146_n2688# 0.270934f
C180 source.n5 a_n2146_n2688# 1.68117f
C181 source.n6 a_n2146_n2688# 0.325128f
C182 source.t29 a_n2146_n2688# 0.270934f
C183 source.t34 a_n2146_n2688# 0.270934f
C184 source.n7 a_n2146_n2688# 1.68117f
C185 source.n8 a_n2146_n2688# 0.325128f
C186 source.t27 a_n2146_n2688# 2.04764f
C187 source.n9 a_n2146_n2688# 0.439009f
C188 source.t38 a_n2146_n2688# 2.04764f
C189 source.n10 a_n2146_n2688# 0.439009f
C190 source.t11 a_n2146_n2688# 0.270934f
C191 source.t14 a_n2146_n2688# 0.270934f
C192 source.n11 a_n2146_n2688# 1.68117f
C193 source.n12 a_n2146_n2688# 0.325128f
C194 source.t39 a_n2146_n2688# 0.270934f
C195 source.t0 a_n2146_n2688# 0.270934f
C196 source.n13 a_n2146_n2688# 1.68117f
C197 source.n14 a_n2146_n2688# 0.325128f
C198 source.t7 a_n2146_n2688# 0.270934f
C199 source.t12 a_n2146_n2688# 0.270934f
C200 source.n15 a_n2146_n2688# 1.68117f
C201 source.n16 a_n2146_n2688# 0.325128f
C202 source.t2 a_n2146_n2688# 0.270934f
C203 source.t9 a_n2146_n2688# 0.270934f
C204 source.n17 a_n2146_n2688# 1.68117f
C205 source.n18 a_n2146_n2688# 0.325128f
C206 source.t17 a_n2146_n2688# 2.04764f
C207 source.n19 a_n2146_n2688# 1.50798f
C208 source.t19 a_n2146_n2688# 2.04763f
C209 source.n20 a_n2146_n2688# 1.50799f
C210 source.t32 a_n2146_n2688# 0.270934f
C211 source.t36 a_n2146_n2688# 0.270934f
C212 source.n21 a_n2146_n2688# 1.68117f
C213 source.n22 a_n2146_n2688# 0.325132f
C214 source.t26 a_n2146_n2688# 0.270934f
C215 source.t22 a_n2146_n2688# 0.270934f
C216 source.n23 a_n2146_n2688# 1.68117f
C217 source.n24 a_n2146_n2688# 0.325132f
C218 source.t33 a_n2146_n2688# 0.270934f
C219 source.t30 a_n2146_n2688# 0.270934f
C220 source.n25 a_n2146_n2688# 1.68117f
C221 source.n26 a_n2146_n2688# 0.325132f
C222 source.t24 a_n2146_n2688# 0.270934f
C223 source.t25 a_n2146_n2688# 0.270934f
C224 source.n27 a_n2146_n2688# 1.68117f
C225 source.n28 a_n2146_n2688# 0.325132f
C226 source.t20 a_n2146_n2688# 2.04763f
C227 source.n29 a_n2146_n2688# 0.439014f
C228 source.t16 a_n2146_n2688# 2.04763f
C229 source.n30 a_n2146_n2688# 0.439014f
C230 source.t8 a_n2146_n2688# 0.270934f
C231 source.t3 a_n2146_n2688# 0.270934f
C232 source.n31 a_n2146_n2688# 1.68117f
C233 source.n32 a_n2146_n2688# 0.325132f
C234 source.t5 a_n2146_n2688# 0.270934f
C235 source.t1 a_n2146_n2688# 0.270934f
C236 source.n33 a_n2146_n2688# 1.68117f
C237 source.n34 a_n2146_n2688# 0.325132f
C238 source.t10 a_n2146_n2688# 0.270934f
C239 source.t13 a_n2146_n2688# 0.270934f
C240 source.n35 a_n2146_n2688# 1.68117f
C241 source.n36 a_n2146_n2688# 0.325132f
C242 source.t6 a_n2146_n2688# 0.270934f
C243 source.t4 a_n2146_n2688# 0.270934f
C244 source.n37 a_n2146_n2688# 1.68117f
C245 source.n38 a_n2146_n2688# 0.325132f
C246 source.t15 a_n2146_n2688# 2.04763f
C247 source.n39 a_n2146_n2688# 0.58206f
C248 source.n40 a_n2146_n2688# 1.30959f
C249 plus.n0 a_n2146_n2688# 0.053349f
C250 plus.t15 a_n2146_n2688# 0.204082f
C251 plus.t8 a_n2146_n2688# 0.204082f
C252 plus.n1 a_n2146_n2688# 0.01852f
C253 plus.n2 a_n2146_n2688# 0.053349f
C254 plus.t16 a_n2146_n2688# 0.204082f
C255 plus.t19 a_n2146_n2688# 0.204082f
C256 plus.t10 a_n2146_n2688# 0.204082f
C257 plus.n3 a_n2146_n2688# 0.093444f
C258 plus.n4 a_n2146_n2688# 0.053349f
C259 plus.t14 a_n2146_n2688# 0.204082f
C260 plus.t17 a_n2146_n2688# 0.204082f
C261 plus.n5 a_n2146_n2688# 0.093444f
C262 plus.t9 a_n2146_n2688# 0.207549f
C263 plus.n6 a_n2146_n2688# 0.115157f
C264 plus.n7 a_n2146_n2688# 0.123063f
C265 plus.n8 a_n2146_n2688# 0.022632f
C266 plus.n9 a_n2146_n2688# 0.093444f
C267 plus.n10 a_n2146_n2688# 0.021809f
C268 plus.n11 a_n2146_n2688# 0.01852f
C269 plus.n12 a_n2146_n2688# 0.053349f
C270 plus.n13 a_n2146_n2688# 0.053349f
C271 plus.n14 a_n2146_n2688# 0.022632f
C272 plus.n15 a_n2146_n2688# 0.093444f
C273 plus.n16 a_n2146_n2688# 0.022632f
C274 plus.n17 a_n2146_n2688# 0.093444f
C275 plus.t13 a_n2146_n2688# 0.204082f
C276 plus.n18 a_n2146_n2688# 0.093444f
C277 plus.n19 a_n2146_n2688# 0.022632f
C278 plus.n20 a_n2146_n2688# 0.053349f
C279 plus.n21 a_n2146_n2688# 0.053349f
C280 plus.n22 a_n2146_n2688# 0.053349f
C281 plus.n23 a_n2146_n2688# 0.021809f
C282 plus.n24 a_n2146_n2688# 0.093444f
C283 plus.n25 a_n2146_n2688# 0.022632f
C284 plus.n26 a_n2146_n2688# 0.093444f
C285 plus.t12 a_n2146_n2688# 0.207549f
C286 plus.n27 a_n2146_n2688# 0.115075f
C287 plus.n28 a_n2146_n2688# 0.531945f
C288 plus.n29 a_n2146_n2688# 0.053349f
C289 plus.t11 a_n2146_n2688# 0.207549f
C290 plus.t4 a_n2146_n2688# 0.204082f
C291 plus.t2 a_n2146_n2688# 0.204082f
C292 plus.n30 a_n2146_n2688# 0.01852f
C293 plus.n31 a_n2146_n2688# 0.053349f
C294 plus.t1 a_n2146_n2688# 0.204082f
C295 plus.n32 a_n2146_n2688# 0.093444f
C296 plus.t18 a_n2146_n2688# 0.204082f
C297 plus.t6 a_n2146_n2688# 0.204082f
C298 plus.t3 a_n2146_n2688# 0.204082f
C299 plus.n33 a_n2146_n2688# 0.093444f
C300 plus.n34 a_n2146_n2688# 0.053349f
C301 plus.t0 a_n2146_n2688# 0.204082f
C302 plus.t7 a_n2146_n2688# 0.204082f
C303 plus.n35 a_n2146_n2688# 0.093444f
C304 plus.t5 a_n2146_n2688# 0.207549f
C305 plus.n36 a_n2146_n2688# 0.115157f
C306 plus.n37 a_n2146_n2688# 0.123063f
C307 plus.n38 a_n2146_n2688# 0.022632f
C308 plus.n39 a_n2146_n2688# 0.093444f
C309 plus.n40 a_n2146_n2688# 0.021809f
C310 plus.n41 a_n2146_n2688# 0.01852f
C311 plus.n42 a_n2146_n2688# 0.053349f
C312 plus.n43 a_n2146_n2688# 0.053349f
C313 plus.n44 a_n2146_n2688# 0.022632f
C314 plus.n45 a_n2146_n2688# 0.093444f
C315 plus.n46 a_n2146_n2688# 0.022632f
C316 plus.n47 a_n2146_n2688# 0.093444f
C317 plus.n48 a_n2146_n2688# 0.022632f
C318 plus.n49 a_n2146_n2688# 0.053349f
C319 plus.n50 a_n2146_n2688# 0.053349f
C320 plus.n51 a_n2146_n2688# 0.053349f
C321 plus.n52 a_n2146_n2688# 0.021809f
C322 plus.n53 a_n2146_n2688# 0.093444f
C323 plus.n54 a_n2146_n2688# 0.022632f
C324 plus.n55 a_n2146_n2688# 0.093444f
C325 plus.n56 a_n2146_n2688# 0.115075f
C326 plus.n57 a_n2146_n2688# 1.56805f
.ends

