* NGSPICE file created from diffpair594.ext - technology: sky130A

.subckt diffpair594 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t9 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 drain_left.t8 plus.t1 source.t14 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X2 a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X3 drain_right.t9 minus.t0 source.t5 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X4 a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X5 drain_right.t8 minus.t1 source.t7 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X6 drain_right.t7 minus.t2 source.t6 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X7 drain_left.t7 plus.t2 source.t13 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X8 drain_left.t6 plus.t3 source.t12 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X9 drain_left.t5 plus.t4 source.t11 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X10 source.t15 plus.t5 drain_left.t4 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X11 drain_right.t6 minus.t3 source.t0 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X12 source.t4 minus.t4 drain_right.t5 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X13 a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X14 drain_right.t4 minus.t5 source.t1 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X15 source.t10 plus.t6 drain_left.t3 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X16 a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X17 drain_left.t2 plus.t7 source.t8 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X18 source.t16 plus.t8 drain_left.t1 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X19 source.t3 minus.t6 drain_right.t3 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X20 source.t2 minus.t7 drain_right.t2 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X21 drain_right.t1 minus.t8 source.t18 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X22 source.t19 minus.t9 drain_right.t0 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X23 source.t17 plus.t9 drain_left.t0 a_n1472_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
R0 plus.n3 plus.t2 1749.08
R1 plus.n9 plus.t4 1749.08
R2 plus.n14 plus.t0 1749.08
R3 plus.n20 plus.t3 1749.08
R4 plus.n6 plus.t7 1711.1
R5 plus.n2 plus.t5 1711.1
R6 plus.n8 plus.t9 1711.1
R7 plus.n17 plus.t1 1711.1
R8 plus.n13 plus.t6 1711.1
R9 plus.n19 plus.t8 1711.1
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 54.0429
R25 plus.n9 plus.n8 54.0429
R26 plus.n20 plus.n19 54.0429
R27 plus.n14 plus.n13 54.0429
R28 plus plus.n21 31.5956
R29 plus.n2 plus.n1 18.9884
R30 plus.n8 plus.n7 18.9884
R31 plus.n19 plus.n18 18.9884
R32 plus.n13 plus.n12 18.9884
R33 plus plus.n10 15.1615
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n0 source.t11 44.1297
R41 source.n5 source.t1 44.1296
R42 source.n19 source.t0 44.1295
R43 source.n14 source.t9 44.1295
R44 source.n2 source.n1 43.1397
R45 source.n4 source.n3 43.1397
R46 source.n7 source.n6 43.1397
R47 source.n9 source.n8 43.1397
R48 source.n18 source.n17 43.1396
R49 source.n16 source.n15 43.1396
R50 source.n13 source.n12 43.1396
R51 source.n11 source.n10 43.1396
R52 source.n11 source.n9 28.4345
R53 source.n20 source.n0 22.357
R54 source.n20 source.n19 5.53498
R55 source.n17 source.t7 0.9905
R56 source.n17 source.t3 0.9905
R57 source.n15 source.t6 0.9905
R58 source.n15 source.t2 0.9905
R59 source.n12 source.t14 0.9905
R60 source.n12 source.t10 0.9905
R61 source.n10 source.t12 0.9905
R62 source.n10 source.t16 0.9905
R63 source.n1 source.t8 0.9905
R64 source.n1 source.t17 0.9905
R65 source.n3 source.t13 0.9905
R66 source.n3 source.t15 0.9905
R67 source.n6 source.t5 0.9905
R68 source.n6 source.t19 0.9905
R69 source.n8 source.t18 0.9905
R70 source.n8 source.t4 0.9905
R71 source.n5 source.n4 0.741879
R72 source.n16 source.n14 0.741879
R73 source.n9 source.n7 0.543603
R74 source.n7 source.n5 0.543603
R75 source.n4 source.n2 0.543603
R76 source.n2 source.n0 0.543603
R77 source.n13 source.n11 0.543603
R78 source.n14 source.n13 0.543603
R79 source.n18 source.n16 0.543603
R80 source.n19 source.n18 0.543603
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t7 61.3515
R83 drain_left.n1 drain_left.t6 61.3514
R84 drain_left.n3 drain_left.n2 60.1704
R85 drain_left.n7 drain_left.n6 59.8185
R86 drain_left.n5 drain_left.n4 59.8185
R87 drain_left.n1 drain_left.n0 59.8184
R88 drain_left drain_left.n3 35.7359
R89 drain_left drain_left.n7 6.19632
R90 drain_left.n2 drain_left.t3 0.9905
R91 drain_left.n2 drain_left.t9 0.9905
R92 drain_left.n0 drain_left.t1 0.9905
R93 drain_left.n0 drain_left.t8 0.9905
R94 drain_left.n6 drain_left.t0 0.9905
R95 drain_left.n6 drain_left.t5 0.9905
R96 drain_left.n4 drain_left.t4 0.9905
R97 drain_left.n4 drain_left.t2 0.9905
R98 drain_left.n7 drain_left.n5 0.543603
R99 drain_left.n3 drain_left.n1 0.0809298
R100 minus.n9 minus.t8 1749.08
R101 minus.n3 minus.t5 1749.08
R102 minus.n20 minus.t3 1749.08
R103 minus.n14 minus.t2 1749.08
R104 minus.n6 minus.t0 1711.1
R105 minus.n8 minus.t4 1711.1
R106 minus.n2 minus.t9 1711.1
R107 minus.n17 minus.t1 1711.1
R108 minus.n19 minus.t6 1711.1
R109 minus.n13 minus.t7 1711.1
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 54.0429
R125 minus.n3 minus.n2 54.0429
R126 minus.n14 minus.n13 54.0429
R127 minus.n20 minus.n19 54.0429
R128 minus.n22 minus.n10 40.7448
R129 minus.n8 minus.n7 18.9884
R130 minus.n2 minus.n1 18.9884
R131 minus.n13 minus.n12 18.9884
R132 minus.n19 minus.n18 18.9884
R133 minus.n22 minus.n21 6.48724
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t7 61.3514
R142 drain_right.n7 drain_right.t1 60.8084
R143 drain_right.n6 drain_right.n4 60.3616
R144 drain_right.n3 drain_right.n2 60.1704
R145 drain_right.n6 drain_right.n5 59.8185
R146 drain_right.n1 drain_right.n0 59.8184
R147 drain_right drain_right.n3 35.1826
R148 drain_right drain_right.n7 5.92477
R149 drain_right.n2 drain_right.t3 0.9905
R150 drain_right.n2 drain_right.t6 0.9905
R151 drain_right.n0 drain_right.t2 0.9905
R152 drain_right.n0 drain_right.t8 0.9905
R153 drain_right.n4 drain_right.t0 0.9905
R154 drain_right.n4 drain_right.t4 0.9905
R155 drain_right.n5 drain_right.t5 0.9905
R156 drain_right.n5 drain_right.t9 0.9905
R157 drain_right.n7 drain_right.n6 0.543603
R158 drain_right.n3 drain_right.n1 0.0809298
C0 source drain_left 33.6492f
C1 minus drain_left 0.171269f
C2 drain_right drain_left 0.728007f
C3 source minus 5.66287f
C4 drain_right source 33.631603f
C5 plus drain_left 6.54084f
C6 drain_right minus 6.40513f
C7 source plus 5.67799f
C8 plus minus 6.46934f
C9 drain_right plus 0.298091f
C10 drain_right a_n1472_n4888# 9.2716f
C11 drain_left a_n1472_n4888# 9.51052f
C12 source a_n1472_n4888# 8.892789f
C13 minus a_n1472_n4888# 6.232105f
C14 plus a_n1472_n4888# 8.77507f
C15 drain_right.t7 a_n1472_n4888# 5.5125f
C16 drain_right.t2 a_n1472_n4888# 0.471154f
C17 drain_right.t8 a_n1472_n4888# 0.471154f
C18 drain_right.n0 a_n1472_n4888# 4.30739f
C19 drain_right.n1 a_n1472_n4888# 0.715655f
C20 drain_right.t3 a_n1472_n4888# 0.471154f
C21 drain_right.t6 a_n1472_n4888# 0.471154f
C22 drain_right.n2 a_n1472_n4888# 4.30945f
C23 drain_right.n3 a_n1472_n4888# 2.21295f
C24 drain_right.t0 a_n1472_n4888# 0.471154f
C25 drain_right.t4 a_n1472_n4888# 0.471154f
C26 drain_right.n4 a_n1472_n4888# 4.3107f
C27 drain_right.t5 a_n1472_n4888# 0.471154f
C28 drain_right.t9 a_n1472_n4888# 0.471154f
C29 drain_right.n5 a_n1472_n4888# 4.30739f
C30 drain_right.n6 a_n1472_n4888# 0.720515f
C31 drain_right.t1 a_n1472_n4888# 5.50899f
C32 drain_right.n7 a_n1472_n4888# 0.647814f
C33 minus.n0 a_n1472_n4888# 0.053991f
C34 minus.t8 a_n1472_n4888# 0.919785f
C35 minus.t4 a_n1472_n4888# 0.912383f
C36 minus.t0 a_n1472_n4888# 0.912383f
C37 minus.n1 a_n1472_n4888# 0.022238f
C38 minus.t9 a_n1472_n4888# 0.912383f
C39 minus.n2 a_n1472_n4888# 0.338928f
C40 minus.t5 a_n1472_n4888# 0.919785f
C41 minus.n3 a_n1472_n4888# 0.355837f
C42 minus.n4 a_n1472_n4888# 0.118558f
C43 minus.n5 a_n1472_n4888# 0.053991f
C44 minus.n6 a_n1472_n4888# 0.356839f
C45 minus.n7 a_n1472_n4888# 0.022238f
C46 minus.n8 a_n1472_n4888# 0.338928f
C47 minus.n9 a_n1472_n4888# 0.355761f
C48 minus.n10 a_n1472_n4888# 2.28552f
C49 minus.n11 a_n1472_n4888# 0.053991f
C50 minus.t6 a_n1472_n4888# 0.912383f
C51 minus.t1 a_n1472_n4888# 0.912383f
C52 minus.n12 a_n1472_n4888# 0.022238f
C53 minus.t2 a_n1472_n4888# 0.919785f
C54 minus.t7 a_n1472_n4888# 0.912383f
C55 minus.n13 a_n1472_n4888# 0.338928f
C56 minus.n14 a_n1472_n4888# 0.355837f
C57 minus.n15 a_n1472_n4888# 0.118558f
C58 minus.n16 a_n1472_n4888# 0.053991f
C59 minus.n17 a_n1472_n4888# 0.356839f
C60 minus.n18 a_n1472_n4888# 0.022238f
C61 minus.n19 a_n1472_n4888# 0.338928f
C62 minus.t3 a_n1472_n4888# 0.919785f
C63 minus.n20 a_n1472_n4888# 0.355761f
C64 minus.n21 a_n1472_n4888# 0.351354f
C65 minus.n22 a_n1472_n4888# 2.73962f
C66 drain_left.t6 a_n1472_n4888# 5.51021f
C67 drain_left.t1 a_n1472_n4888# 0.470959f
C68 drain_left.t8 a_n1472_n4888# 0.470959f
C69 drain_left.n0 a_n1472_n4888# 4.30561f
C70 drain_left.n1 a_n1472_n4888# 0.715359f
C71 drain_left.t3 a_n1472_n4888# 0.470959f
C72 drain_left.t9 a_n1472_n4888# 0.470959f
C73 drain_left.n2 a_n1472_n4888# 4.30767f
C74 drain_left.n3 a_n1472_n4888# 2.27441f
C75 drain_left.t7 a_n1472_n4888# 5.51024f
C76 drain_left.t4 a_n1472_n4888# 0.470959f
C77 drain_left.t2 a_n1472_n4888# 0.470959f
C78 drain_left.n4 a_n1472_n4888# 4.3056f
C79 drain_left.n5 a_n1472_n4888# 0.75118f
C80 drain_left.t0 a_n1472_n4888# 0.470959f
C81 drain_left.t5 a_n1472_n4888# 0.470959f
C82 drain_left.n6 a_n1472_n4888# 4.3056f
C83 drain_left.n7 a_n1472_n4888# 0.603796f
C84 source.t11 a_n1472_n4888# 5.45499f
C85 source.n0 a_n1472_n4888# 2.32019f
C86 source.t8 a_n1472_n4888# 0.477319f
C87 source.t17 a_n1472_n4888# 0.477319f
C88 source.n1 a_n1472_n4888# 4.26744f
C89 source.n2 a_n1472_n4888# 0.41583f
C90 source.t13 a_n1472_n4888# 0.477319f
C91 source.t15 a_n1472_n4888# 0.477319f
C92 source.n3 a_n1472_n4888# 4.26744f
C93 source.n4 a_n1472_n4888# 0.435125f
C94 source.t1 a_n1472_n4888# 5.455f
C95 source.n5 a_n1472_n4888# 0.549346f
C96 source.t5 a_n1472_n4888# 0.477319f
C97 source.t19 a_n1472_n4888# 0.477319f
C98 source.n6 a_n1472_n4888# 4.26744f
C99 source.n7 a_n1472_n4888# 0.41583f
C100 source.t18 a_n1472_n4888# 0.477319f
C101 source.t4 a_n1472_n4888# 0.477319f
C102 source.n8 a_n1472_n4888# 4.26744f
C103 source.n9 a_n1472_n4888# 2.79402f
C104 source.t12 a_n1472_n4888# 0.477319f
C105 source.t16 a_n1472_n4888# 0.477319f
C106 source.n10 a_n1472_n4888# 4.26745f
C107 source.n11 a_n1472_n4888# 2.79401f
C108 source.t14 a_n1472_n4888# 0.477319f
C109 source.t10 a_n1472_n4888# 0.477319f
C110 source.n12 a_n1472_n4888# 4.26745f
C111 source.n13 a_n1472_n4888# 0.415822f
C112 source.t9 a_n1472_n4888# 5.45497f
C113 source.n14 a_n1472_n4888# 0.549376f
C114 source.t6 a_n1472_n4888# 0.477319f
C115 source.t2 a_n1472_n4888# 0.477319f
C116 source.n15 a_n1472_n4888# 4.26745f
C117 source.n16 a_n1472_n4888# 0.435117f
C118 source.t7 a_n1472_n4888# 0.477319f
C119 source.t3 a_n1472_n4888# 0.477319f
C120 source.n17 a_n1472_n4888# 4.26745f
C121 source.n18 a_n1472_n4888# 0.415822f
C122 source.t0 a_n1472_n4888# 5.45497f
C123 source.n19 a_n1472_n4888# 0.693436f
C124 source.n20 a_n1472_n4888# 2.71868f
C125 plus.n0 a_n1472_n4888# 0.054602f
C126 plus.t9 a_n1472_n4888# 0.922704f
C127 plus.t7 a_n1472_n4888# 0.922704f
C128 plus.n1 a_n1472_n4888# 0.02249f
C129 plus.t2 a_n1472_n4888# 0.93019f
C130 plus.t5 a_n1472_n4888# 0.922704f
C131 plus.n2 a_n1472_n4888# 0.342762f
C132 plus.n3 a_n1472_n4888# 0.359863f
C133 plus.n4 a_n1472_n4888# 0.119899f
C134 plus.n5 a_n1472_n4888# 0.054602f
C135 plus.n6 a_n1472_n4888# 0.360876f
C136 plus.n7 a_n1472_n4888# 0.02249f
C137 plus.n8 a_n1472_n4888# 0.342762f
C138 plus.t4 a_n1472_n4888# 0.93019f
C139 plus.n9 a_n1472_n4888# 0.359786f
C140 plus.n10 a_n1472_n4888# 0.827484f
C141 plus.n11 a_n1472_n4888# 0.054602f
C142 plus.t3 a_n1472_n4888# 0.93019f
C143 plus.t8 a_n1472_n4888# 0.922704f
C144 plus.t1 a_n1472_n4888# 0.922704f
C145 plus.n12 a_n1472_n4888# 0.02249f
C146 plus.t6 a_n1472_n4888# 0.922704f
C147 plus.n13 a_n1472_n4888# 0.342762f
C148 plus.t0 a_n1472_n4888# 0.93019f
C149 plus.n14 a_n1472_n4888# 0.359863f
C150 plus.n15 a_n1472_n4888# 0.119899f
C151 plus.n16 a_n1472_n4888# 0.054602f
C152 plus.n17 a_n1472_n4888# 0.360876f
C153 plus.n18 a_n1472_n4888# 0.02249f
C154 plus.n19 a_n1472_n4888# 0.342762f
C155 plus.n20 a_n1472_n4888# 0.359786f
C156 plus.n21 a_n1472_n4888# 1.81816f
.ends

