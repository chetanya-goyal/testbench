* NGSPICE file created from diffpair428.ext - technology: sky130A

.subckt diffpair428 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t24 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 drain_left.t18 plus.t1 source.t28 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 drain_left.t17 plus.t2 source.t34 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X3 source.t15 minus.t0 drain_right.t19 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X4 drain_left.t16 plus.t3 source.t22 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X5 source.t9 minus.t1 drain_right.t18 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 drain_right.t17 minus.t2 source.t8 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X7 a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X8 drain_right.t16 minus.t3 source.t2 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X9 drain_left.t15 plus.t4 source.t25 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 source.t18 plus.t5 drain_left.t14 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X11 source.t6 minus.t4 drain_right.t15 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X12 source.t31 plus.t6 drain_left.t13 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X13 source.t10 minus.t5 drain_right.t14 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X14 source.t11 minus.t6 drain_right.t13 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X15 drain_left.t12 plus.t7 source.t29 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X16 source.t16 minus.t7 drain_right.t12 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X17 source.t36 plus.t8 drain_left.t11 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X18 source.t35 plus.t9 drain_left.t10 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X19 source.t23 plus.t10 drain_left.t9 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X20 a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X21 source.t1 minus.t8 drain_right.t11 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X22 drain_right.t10 minus.t9 source.t3 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X23 source.t26 plus.t11 drain_left.t8 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X24 source.t20 plus.t12 drain_left.t7 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X25 drain_right.t9 minus.t10 source.t39 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X26 drain_right.t8 minus.t11 source.t5 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X27 a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X28 drain_left.t6 plus.t13 source.t19 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X29 drain_right.t7 minus.t12 source.t0 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X30 source.t32 plus.t14 drain_left.t5 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X31 drain_left.t4 plus.t15 source.t30 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X32 source.t4 minus.t13 drain_right.t6 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X33 source.t14 minus.t14 drain_right.t5 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X34 source.t37 plus.t16 drain_left.t3 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X35 drain_right.t4 minus.t15 source.t12 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X36 drain_right.t3 minus.t16 source.t17 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X37 drain_left.t2 plus.t17 source.t27 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X38 drain_right.t2 minus.t17 source.t38 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X39 drain_right.t1 minus.t18 source.t13 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X40 drain_left.t1 plus.t18 source.t33 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X41 source.t7 minus.t19 drain_right.t0 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X42 a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X43 source.t21 plus.t19 drain_left.t0 a_n1992_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n6 plus.t5 1334.7
R1 plus.n25 plus.t2 1334.7
R2 plus.n33 plus.t17 1334.7
R3 plus.n52 plus.t11 1334.7
R4 plus.n5 plus.t1 1282.12
R5 plus.n9 plus.t10 1282.12
R6 plus.n11 plus.t0 1282.12
R7 plus.n3 plus.t9 1282.12
R8 plus.n17 plus.t18 1282.12
R9 plus.n1 plus.t8 1282.12
R10 plus.n22 plus.t3 1282.12
R11 plus.n24 plus.t12 1282.12
R12 plus.n32 plus.t14 1282.12
R13 plus.n36 plus.t7 1282.12
R14 plus.n38 plus.t19 1282.12
R15 plus.n30 plus.t4 1282.12
R16 plus.n44 plus.t16 1282.12
R17 plus.n28 plus.t13 1282.12
R18 plus.n49 plus.t6 1282.12
R19 plus.n51 plus.t15 1282.12
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus plus.n53 30.5445
R63 plus.n10 plus.n9 29.2126
R64 plus.n22 plus.n21 29.2126
R65 plus.n49 plus.n48 29.2126
R66 plus.n37 plus.n36 29.2126
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 12.1407
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n554 source.n494 289.615
R93 source.n480 source.n420 289.615
R94 source.n414 source.n354 289.615
R95 source.n340 source.n280 289.615
R96 source.n60 source.n0 289.615
R97 source.n134 source.n74 289.615
R98 source.n200 source.n140 289.615
R99 source.n274 source.n214 289.615
R100 source.n514 source.n513 185
R101 source.n519 source.n518 185
R102 source.n521 source.n520 185
R103 source.n510 source.n509 185
R104 source.n527 source.n526 185
R105 source.n529 source.n528 185
R106 source.n506 source.n505 185
R107 source.n536 source.n535 185
R108 source.n537 source.n504 185
R109 source.n539 source.n538 185
R110 source.n502 source.n501 185
R111 source.n545 source.n544 185
R112 source.n547 source.n546 185
R113 source.n498 source.n497 185
R114 source.n553 source.n552 185
R115 source.n555 source.n554 185
R116 source.n440 source.n439 185
R117 source.n445 source.n444 185
R118 source.n447 source.n446 185
R119 source.n436 source.n435 185
R120 source.n453 source.n452 185
R121 source.n455 source.n454 185
R122 source.n432 source.n431 185
R123 source.n462 source.n461 185
R124 source.n463 source.n430 185
R125 source.n465 source.n464 185
R126 source.n428 source.n427 185
R127 source.n471 source.n470 185
R128 source.n473 source.n472 185
R129 source.n424 source.n423 185
R130 source.n479 source.n478 185
R131 source.n481 source.n480 185
R132 source.n374 source.n373 185
R133 source.n379 source.n378 185
R134 source.n381 source.n380 185
R135 source.n370 source.n369 185
R136 source.n387 source.n386 185
R137 source.n389 source.n388 185
R138 source.n366 source.n365 185
R139 source.n396 source.n395 185
R140 source.n397 source.n364 185
R141 source.n399 source.n398 185
R142 source.n362 source.n361 185
R143 source.n405 source.n404 185
R144 source.n407 source.n406 185
R145 source.n358 source.n357 185
R146 source.n413 source.n412 185
R147 source.n415 source.n414 185
R148 source.n300 source.n299 185
R149 source.n305 source.n304 185
R150 source.n307 source.n306 185
R151 source.n296 source.n295 185
R152 source.n313 source.n312 185
R153 source.n315 source.n314 185
R154 source.n292 source.n291 185
R155 source.n322 source.n321 185
R156 source.n323 source.n290 185
R157 source.n325 source.n324 185
R158 source.n288 source.n287 185
R159 source.n331 source.n330 185
R160 source.n333 source.n332 185
R161 source.n284 source.n283 185
R162 source.n339 source.n338 185
R163 source.n341 source.n340 185
R164 source.n61 source.n60 185
R165 source.n59 source.n58 185
R166 source.n4 source.n3 185
R167 source.n53 source.n52 185
R168 source.n51 source.n50 185
R169 source.n8 source.n7 185
R170 source.n45 source.n44 185
R171 source.n43 source.n10 185
R172 source.n42 source.n41 185
R173 source.n13 source.n11 185
R174 source.n36 source.n35 185
R175 source.n34 source.n33 185
R176 source.n17 source.n16 185
R177 source.n28 source.n27 185
R178 source.n26 source.n25 185
R179 source.n21 source.n20 185
R180 source.n135 source.n134 185
R181 source.n133 source.n132 185
R182 source.n78 source.n77 185
R183 source.n127 source.n126 185
R184 source.n125 source.n124 185
R185 source.n82 source.n81 185
R186 source.n119 source.n118 185
R187 source.n117 source.n84 185
R188 source.n116 source.n115 185
R189 source.n87 source.n85 185
R190 source.n110 source.n109 185
R191 source.n108 source.n107 185
R192 source.n91 source.n90 185
R193 source.n102 source.n101 185
R194 source.n100 source.n99 185
R195 source.n95 source.n94 185
R196 source.n201 source.n200 185
R197 source.n199 source.n198 185
R198 source.n144 source.n143 185
R199 source.n193 source.n192 185
R200 source.n191 source.n190 185
R201 source.n148 source.n147 185
R202 source.n185 source.n184 185
R203 source.n183 source.n150 185
R204 source.n182 source.n181 185
R205 source.n153 source.n151 185
R206 source.n176 source.n175 185
R207 source.n174 source.n173 185
R208 source.n157 source.n156 185
R209 source.n168 source.n167 185
R210 source.n166 source.n165 185
R211 source.n161 source.n160 185
R212 source.n275 source.n274 185
R213 source.n273 source.n272 185
R214 source.n218 source.n217 185
R215 source.n267 source.n266 185
R216 source.n265 source.n264 185
R217 source.n222 source.n221 185
R218 source.n259 source.n258 185
R219 source.n257 source.n224 185
R220 source.n256 source.n255 185
R221 source.n227 source.n225 185
R222 source.n250 source.n249 185
R223 source.n248 source.n247 185
R224 source.n231 source.n230 185
R225 source.n242 source.n241 185
R226 source.n240 source.n239 185
R227 source.n235 source.n234 185
R228 source.n515 source.t2 149.524
R229 source.n441 source.t7 149.524
R230 source.n375 source.t27 149.524
R231 source.n301 source.t26 149.524
R232 source.n22 source.t34 149.524
R233 source.n96 source.t18 149.524
R234 source.n162 source.t39 149.524
R235 source.n236 source.t16 149.524
R236 source.n519 source.n513 104.615
R237 source.n520 source.n519 104.615
R238 source.n520 source.n509 104.615
R239 source.n527 source.n509 104.615
R240 source.n528 source.n527 104.615
R241 source.n528 source.n505 104.615
R242 source.n536 source.n505 104.615
R243 source.n537 source.n536 104.615
R244 source.n538 source.n537 104.615
R245 source.n538 source.n501 104.615
R246 source.n545 source.n501 104.615
R247 source.n546 source.n545 104.615
R248 source.n546 source.n497 104.615
R249 source.n553 source.n497 104.615
R250 source.n554 source.n553 104.615
R251 source.n445 source.n439 104.615
R252 source.n446 source.n445 104.615
R253 source.n446 source.n435 104.615
R254 source.n453 source.n435 104.615
R255 source.n454 source.n453 104.615
R256 source.n454 source.n431 104.615
R257 source.n462 source.n431 104.615
R258 source.n463 source.n462 104.615
R259 source.n464 source.n463 104.615
R260 source.n464 source.n427 104.615
R261 source.n471 source.n427 104.615
R262 source.n472 source.n471 104.615
R263 source.n472 source.n423 104.615
R264 source.n479 source.n423 104.615
R265 source.n480 source.n479 104.615
R266 source.n379 source.n373 104.615
R267 source.n380 source.n379 104.615
R268 source.n380 source.n369 104.615
R269 source.n387 source.n369 104.615
R270 source.n388 source.n387 104.615
R271 source.n388 source.n365 104.615
R272 source.n396 source.n365 104.615
R273 source.n397 source.n396 104.615
R274 source.n398 source.n397 104.615
R275 source.n398 source.n361 104.615
R276 source.n405 source.n361 104.615
R277 source.n406 source.n405 104.615
R278 source.n406 source.n357 104.615
R279 source.n413 source.n357 104.615
R280 source.n414 source.n413 104.615
R281 source.n305 source.n299 104.615
R282 source.n306 source.n305 104.615
R283 source.n306 source.n295 104.615
R284 source.n313 source.n295 104.615
R285 source.n314 source.n313 104.615
R286 source.n314 source.n291 104.615
R287 source.n322 source.n291 104.615
R288 source.n323 source.n322 104.615
R289 source.n324 source.n323 104.615
R290 source.n324 source.n287 104.615
R291 source.n331 source.n287 104.615
R292 source.n332 source.n331 104.615
R293 source.n332 source.n283 104.615
R294 source.n339 source.n283 104.615
R295 source.n340 source.n339 104.615
R296 source.n60 source.n59 104.615
R297 source.n59 source.n3 104.615
R298 source.n52 source.n3 104.615
R299 source.n52 source.n51 104.615
R300 source.n51 source.n7 104.615
R301 source.n44 source.n7 104.615
R302 source.n44 source.n43 104.615
R303 source.n43 source.n42 104.615
R304 source.n42 source.n11 104.615
R305 source.n35 source.n11 104.615
R306 source.n35 source.n34 104.615
R307 source.n34 source.n16 104.615
R308 source.n27 source.n16 104.615
R309 source.n27 source.n26 104.615
R310 source.n26 source.n20 104.615
R311 source.n134 source.n133 104.615
R312 source.n133 source.n77 104.615
R313 source.n126 source.n77 104.615
R314 source.n126 source.n125 104.615
R315 source.n125 source.n81 104.615
R316 source.n118 source.n81 104.615
R317 source.n118 source.n117 104.615
R318 source.n117 source.n116 104.615
R319 source.n116 source.n85 104.615
R320 source.n109 source.n85 104.615
R321 source.n109 source.n108 104.615
R322 source.n108 source.n90 104.615
R323 source.n101 source.n90 104.615
R324 source.n101 source.n100 104.615
R325 source.n100 source.n94 104.615
R326 source.n200 source.n199 104.615
R327 source.n199 source.n143 104.615
R328 source.n192 source.n143 104.615
R329 source.n192 source.n191 104.615
R330 source.n191 source.n147 104.615
R331 source.n184 source.n147 104.615
R332 source.n184 source.n183 104.615
R333 source.n183 source.n182 104.615
R334 source.n182 source.n151 104.615
R335 source.n175 source.n151 104.615
R336 source.n175 source.n174 104.615
R337 source.n174 source.n156 104.615
R338 source.n167 source.n156 104.615
R339 source.n167 source.n166 104.615
R340 source.n166 source.n160 104.615
R341 source.n274 source.n273 104.615
R342 source.n273 source.n217 104.615
R343 source.n266 source.n217 104.615
R344 source.n266 source.n265 104.615
R345 source.n265 source.n221 104.615
R346 source.n258 source.n221 104.615
R347 source.n258 source.n257 104.615
R348 source.n257 source.n256 104.615
R349 source.n256 source.n225 104.615
R350 source.n249 source.n225 104.615
R351 source.n249 source.n248 104.615
R352 source.n248 source.n230 104.615
R353 source.n241 source.n230 104.615
R354 source.n241 source.n240 104.615
R355 source.n240 source.n234 104.615
R356 source.t2 source.n513 52.3082
R357 source.t7 source.n439 52.3082
R358 source.t27 source.n373 52.3082
R359 source.t26 source.n299 52.3082
R360 source.t34 source.n20 52.3082
R361 source.t18 source.n94 52.3082
R362 source.t39 source.n160 52.3082
R363 source.t16 source.n234 52.3082
R364 source.n67 source.n66 42.8739
R365 source.n69 source.n68 42.8739
R366 source.n71 source.n70 42.8739
R367 source.n73 source.n72 42.8739
R368 source.n207 source.n206 42.8739
R369 source.n209 source.n208 42.8739
R370 source.n211 source.n210 42.8739
R371 source.n213 source.n212 42.8739
R372 source.n493 source.n492 42.8737
R373 source.n491 source.n490 42.8737
R374 source.n489 source.n488 42.8737
R375 source.n487 source.n486 42.8737
R376 source.n353 source.n352 42.8737
R377 source.n351 source.n350 42.8737
R378 source.n349 source.n348 42.8737
R379 source.n347 source.n346 42.8737
R380 source.n559 source.n558 29.8581
R381 source.n485 source.n484 29.8581
R382 source.n419 source.n418 29.8581
R383 source.n345 source.n344 29.8581
R384 source.n65 source.n64 29.8581
R385 source.n139 source.n138 29.8581
R386 source.n205 source.n204 29.8581
R387 source.n279 source.n278 29.8581
R388 source.n345 source.n279 21.7877
R389 source.n560 source.n65 16.2748
R390 source.n539 source.n504 13.1884
R391 source.n465 source.n430 13.1884
R392 source.n399 source.n364 13.1884
R393 source.n325 source.n290 13.1884
R394 source.n45 source.n10 13.1884
R395 source.n119 source.n84 13.1884
R396 source.n185 source.n150 13.1884
R397 source.n259 source.n224 13.1884
R398 source.n535 source.n534 12.8005
R399 source.n540 source.n502 12.8005
R400 source.n461 source.n460 12.8005
R401 source.n466 source.n428 12.8005
R402 source.n395 source.n394 12.8005
R403 source.n400 source.n362 12.8005
R404 source.n321 source.n320 12.8005
R405 source.n326 source.n288 12.8005
R406 source.n46 source.n8 12.8005
R407 source.n41 source.n12 12.8005
R408 source.n120 source.n82 12.8005
R409 source.n115 source.n86 12.8005
R410 source.n186 source.n148 12.8005
R411 source.n181 source.n152 12.8005
R412 source.n260 source.n222 12.8005
R413 source.n255 source.n226 12.8005
R414 source.n533 source.n506 12.0247
R415 source.n544 source.n543 12.0247
R416 source.n459 source.n432 12.0247
R417 source.n470 source.n469 12.0247
R418 source.n393 source.n366 12.0247
R419 source.n404 source.n403 12.0247
R420 source.n319 source.n292 12.0247
R421 source.n330 source.n329 12.0247
R422 source.n50 source.n49 12.0247
R423 source.n40 source.n13 12.0247
R424 source.n124 source.n123 12.0247
R425 source.n114 source.n87 12.0247
R426 source.n190 source.n189 12.0247
R427 source.n180 source.n153 12.0247
R428 source.n264 source.n263 12.0247
R429 source.n254 source.n227 12.0247
R430 source.n530 source.n529 11.249
R431 source.n547 source.n500 11.249
R432 source.n456 source.n455 11.249
R433 source.n473 source.n426 11.249
R434 source.n390 source.n389 11.249
R435 source.n407 source.n360 11.249
R436 source.n316 source.n315 11.249
R437 source.n333 source.n286 11.249
R438 source.n53 source.n6 11.249
R439 source.n37 source.n36 11.249
R440 source.n127 source.n80 11.249
R441 source.n111 source.n110 11.249
R442 source.n193 source.n146 11.249
R443 source.n177 source.n176 11.249
R444 source.n267 source.n220 11.249
R445 source.n251 source.n250 11.249
R446 source.n526 source.n508 10.4732
R447 source.n548 source.n498 10.4732
R448 source.n452 source.n434 10.4732
R449 source.n474 source.n424 10.4732
R450 source.n386 source.n368 10.4732
R451 source.n408 source.n358 10.4732
R452 source.n312 source.n294 10.4732
R453 source.n334 source.n284 10.4732
R454 source.n54 source.n4 10.4732
R455 source.n33 source.n15 10.4732
R456 source.n128 source.n78 10.4732
R457 source.n107 source.n89 10.4732
R458 source.n194 source.n144 10.4732
R459 source.n173 source.n155 10.4732
R460 source.n268 source.n218 10.4732
R461 source.n247 source.n229 10.4732
R462 source.n515 source.n514 10.2747
R463 source.n441 source.n440 10.2747
R464 source.n375 source.n374 10.2747
R465 source.n301 source.n300 10.2747
R466 source.n22 source.n21 10.2747
R467 source.n96 source.n95 10.2747
R468 source.n162 source.n161 10.2747
R469 source.n236 source.n235 10.2747
R470 source.n525 source.n510 9.69747
R471 source.n552 source.n551 9.69747
R472 source.n451 source.n436 9.69747
R473 source.n478 source.n477 9.69747
R474 source.n385 source.n370 9.69747
R475 source.n412 source.n411 9.69747
R476 source.n311 source.n296 9.69747
R477 source.n338 source.n337 9.69747
R478 source.n58 source.n57 9.69747
R479 source.n32 source.n17 9.69747
R480 source.n132 source.n131 9.69747
R481 source.n106 source.n91 9.69747
R482 source.n198 source.n197 9.69747
R483 source.n172 source.n157 9.69747
R484 source.n272 source.n271 9.69747
R485 source.n246 source.n231 9.69747
R486 source.n558 source.n557 9.45567
R487 source.n484 source.n483 9.45567
R488 source.n418 source.n417 9.45567
R489 source.n344 source.n343 9.45567
R490 source.n64 source.n63 9.45567
R491 source.n138 source.n137 9.45567
R492 source.n204 source.n203 9.45567
R493 source.n278 source.n277 9.45567
R494 source.n557 source.n556 9.3005
R495 source.n496 source.n495 9.3005
R496 source.n551 source.n550 9.3005
R497 source.n549 source.n548 9.3005
R498 source.n500 source.n499 9.3005
R499 source.n543 source.n542 9.3005
R500 source.n541 source.n540 9.3005
R501 source.n517 source.n516 9.3005
R502 source.n512 source.n511 9.3005
R503 source.n523 source.n522 9.3005
R504 source.n525 source.n524 9.3005
R505 source.n508 source.n507 9.3005
R506 source.n531 source.n530 9.3005
R507 source.n533 source.n532 9.3005
R508 source.n534 source.n503 9.3005
R509 source.n483 source.n482 9.3005
R510 source.n422 source.n421 9.3005
R511 source.n477 source.n476 9.3005
R512 source.n475 source.n474 9.3005
R513 source.n426 source.n425 9.3005
R514 source.n469 source.n468 9.3005
R515 source.n467 source.n466 9.3005
R516 source.n443 source.n442 9.3005
R517 source.n438 source.n437 9.3005
R518 source.n449 source.n448 9.3005
R519 source.n451 source.n450 9.3005
R520 source.n434 source.n433 9.3005
R521 source.n457 source.n456 9.3005
R522 source.n459 source.n458 9.3005
R523 source.n460 source.n429 9.3005
R524 source.n417 source.n416 9.3005
R525 source.n356 source.n355 9.3005
R526 source.n411 source.n410 9.3005
R527 source.n409 source.n408 9.3005
R528 source.n360 source.n359 9.3005
R529 source.n403 source.n402 9.3005
R530 source.n401 source.n400 9.3005
R531 source.n377 source.n376 9.3005
R532 source.n372 source.n371 9.3005
R533 source.n383 source.n382 9.3005
R534 source.n385 source.n384 9.3005
R535 source.n368 source.n367 9.3005
R536 source.n391 source.n390 9.3005
R537 source.n393 source.n392 9.3005
R538 source.n394 source.n363 9.3005
R539 source.n343 source.n342 9.3005
R540 source.n282 source.n281 9.3005
R541 source.n337 source.n336 9.3005
R542 source.n335 source.n334 9.3005
R543 source.n286 source.n285 9.3005
R544 source.n329 source.n328 9.3005
R545 source.n327 source.n326 9.3005
R546 source.n303 source.n302 9.3005
R547 source.n298 source.n297 9.3005
R548 source.n309 source.n308 9.3005
R549 source.n311 source.n310 9.3005
R550 source.n294 source.n293 9.3005
R551 source.n317 source.n316 9.3005
R552 source.n319 source.n318 9.3005
R553 source.n320 source.n289 9.3005
R554 source.n24 source.n23 9.3005
R555 source.n19 source.n18 9.3005
R556 source.n30 source.n29 9.3005
R557 source.n32 source.n31 9.3005
R558 source.n15 source.n14 9.3005
R559 source.n38 source.n37 9.3005
R560 source.n40 source.n39 9.3005
R561 source.n12 source.n9 9.3005
R562 source.n63 source.n62 9.3005
R563 source.n2 source.n1 9.3005
R564 source.n57 source.n56 9.3005
R565 source.n55 source.n54 9.3005
R566 source.n6 source.n5 9.3005
R567 source.n49 source.n48 9.3005
R568 source.n47 source.n46 9.3005
R569 source.n98 source.n97 9.3005
R570 source.n93 source.n92 9.3005
R571 source.n104 source.n103 9.3005
R572 source.n106 source.n105 9.3005
R573 source.n89 source.n88 9.3005
R574 source.n112 source.n111 9.3005
R575 source.n114 source.n113 9.3005
R576 source.n86 source.n83 9.3005
R577 source.n137 source.n136 9.3005
R578 source.n76 source.n75 9.3005
R579 source.n131 source.n130 9.3005
R580 source.n129 source.n128 9.3005
R581 source.n80 source.n79 9.3005
R582 source.n123 source.n122 9.3005
R583 source.n121 source.n120 9.3005
R584 source.n164 source.n163 9.3005
R585 source.n159 source.n158 9.3005
R586 source.n170 source.n169 9.3005
R587 source.n172 source.n171 9.3005
R588 source.n155 source.n154 9.3005
R589 source.n178 source.n177 9.3005
R590 source.n180 source.n179 9.3005
R591 source.n152 source.n149 9.3005
R592 source.n203 source.n202 9.3005
R593 source.n142 source.n141 9.3005
R594 source.n197 source.n196 9.3005
R595 source.n195 source.n194 9.3005
R596 source.n146 source.n145 9.3005
R597 source.n189 source.n188 9.3005
R598 source.n187 source.n186 9.3005
R599 source.n238 source.n237 9.3005
R600 source.n233 source.n232 9.3005
R601 source.n244 source.n243 9.3005
R602 source.n246 source.n245 9.3005
R603 source.n229 source.n228 9.3005
R604 source.n252 source.n251 9.3005
R605 source.n254 source.n253 9.3005
R606 source.n226 source.n223 9.3005
R607 source.n277 source.n276 9.3005
R608 source.n216 source.n215 9.3005
R609 source.n271 source.n270 9.3005
R610 source.n269 source.n268 9.3005
R611 source.n220 source.n219 9.3005
R612 source.n263 source.n262 9.3005
R613 source.n261 source.n260 9.3005
R614 source.n522 source.n521 8.92171
R615 source.n555 source.n496 8.92171
R616 source.n448 source.n447 8.92171
R617 source.n481 source.n422 8.92171
R618 source.n382 source.n381 8.92171
R619 source.n415 source.n356 8.92171
R620 source.n308 source.n307 8.92171
R621 source.n341 source.n282 8.92171
R622 source.n61 source.n2 8.92171
R623 source.n29 source.n28 8.92171
R624 source.n135 source.n76 8.92171
R625 source.n103 source.n102 8.92171
R626 source.n201 source.n142 8.92171
R627 source.n169 source.n168 8.92171
R628 source.n275 source.n216 8.92171
R629 source.n243 source.n242 8.92171
R630 source.n518 source.n512 8.14595
R631 source.n556 source.n494 8.14595
R632 source.n444 source.n438 8.14595
R633 source.n482 source.n420 8.14595
R634 source.n378 source.n372 8.14595
R635 source.n416 source.n354 8.14595
R636 source.n304 source.n298 8.14595
R637 source.n342 source.n280 8.14595
R638 source.n62 source.n0 8.14595
R639 source.n25 source.n19 8.14595
R640 source.n136 source.n74 8.14595
R641 source.n99 source.n93 8.14595
R642 source.n202 source.n140 8.14595
R643 source.n165 source.n159 8.14595
R644 source.n276 source.n214 8.14595
R645 source.n239 source.n233 8.14595
R646 source.n517 source.n514 7.3702
R647 source.n443 source.n440 7.3702
R648 source.n377 source.n374 7.3702
R649 source.n303 source.n300 7.3702
R650 source.n24 source.n21 7.3702
R651 source.n98 source.n95 7.3702
R652 source.n164 source.n161 7.3702
R653 source.n238 source.n235 7.3702
R654 source.n518 source.n517 5.81868
R655 source.n558 source.n494 5.81868
R656 source.n444 source.n443 5.81868
R657 source.n484 source.n420 5.81868
R658 source.n378 source.n377 5.81868
R659 source.n418 source.n354 5.81868
R660 source.n304 source.n303 5.81868
R661 source.n344 source.n280 5.81868
R662 source.n64 source.n0 5.81868
R663 source.n25 source.n24 5.81868
R664 source.n138 source.n74 5.81868
R665 source.n99 source.n98 5.81868
R666 source.n204 source.n140 5.81868
R667 source.n165 source.n164 5.81868
R668 source.n278 source.n214 5.81868
R669 source.n239 source.n238 5.81868
R670 source.n560 source.n559 5.51343
R671 source.n521 source.n512 5.04292
R672 source.n556 source.n555 5.04292
R673 source.n447 source.n438 5.04292
R674 source.n482 source.n481 5.04292
R675 source.n381 source.n372 5.04292
R676 source.n416 source.n415 5.04292
R677 source.n307 source.n298 5.04292
R678 source.n342 source.n341 5.04292
R679 source.n62 source.n61 5.04292
R680 source.n28 source.n19 5.04292
R681 source.n136 source.n135 5.04292
R682 source.n102 source.n93 5.04292
R683 source.n202 source.n201 5.04292
R684 source.n168 source.n159 5.04292
R685 source.n276 source.n275 5.04292
R686 source.n242 source.n233 5.04292
R687 source.n522 source.n510 4.26717
R688 source.n552 source.n496 4.26717
R689 source.n448 source.n436 4.26717
R690 source.n478 source.n422 4.26717
R691 source.n382 source.n370 4.26717
R692 source.n412 source.n356 4.26717
R693 source.n308 source.n296 4.26717
R694 source.n338 source.n282 4.26717
R695 source.n58 source.n2 4.26717
R696 source.n29 source.n17 4.26717
R697 source.n132 source.n76 4.26717
R698 source.n103 source.n91 4.26717
R699 source.n198 source.n142 4.26717
R700 source.n169 source.n157 4.26717
R701 source.n272 source.n216 4.26717
R702 source.n243 source.n231 4.26717
R703 source.n526 source.n525 3.49141
R704 source.n551 source.n498 3.49141
R705 source.n452 source.n451 3.49141
R706 source.n477 source.n424 3.49141
R707 source.n386 source.n385 3.49141
R708 source.n411 source.n358 3.49141
R709 source.n312 source.n311 3.49141
R710 source.n337 source.n284 3.49141
R711 source.n57 source.n4 3.49141
R712 source.n33 source.n32 3.49141
R713 source.n131 source.n78 3.49141
R714 source.n107 source.n106 3.49141
R715 source.n197 source.n144 3.49141
R716 source.n173 source.n172 3.49141
R717 source.n271 source.n218 3.49141
R718 source.n247 source.n246 3.49141
R719 source.n516 source.n515 2.84303
R720 source.n442 source.n441 2.84303
R721 source.n376 source.n375 2.84303
R722 source.n302 source.n301 2.84303
R723 source.n23 source.n22 2.84303
R724 source.n97 source.n96 2.84303
R725 source.n163 source.n162 2.84303
R726 source.n237 source.n236 2.84303
R727 source.n529 source.n508 2.71565
R728 source.n548 source.n547 2.71565
R729 source.n455 source.n434 2.71565
R730 source.n474 source.n473 2.71565
R731 source.n389 source.n368 2.71565
R732 source.n408 source.n407 2.71565
R733 source.n315 source.n294 2.71565
R734 source.n334 source.n333 2.71565
R735 source.n54 source.n53 2.71565
R736 source.n36 source.n15 2.71565
R737 source.n128 source.n127 2.71565
R738 source.n110 source.n89 2.71565
R739 source.n194 source.n193 2.71565
R740 source.n176 source.n155 2.71565
R741 source.n268 source.n267 2.71565
R742 source.n250 source.n229 2.71565
R743 source.n530 source.n506 1.93989
R744 source.n544 source.n500 1.93989
R745 source.n456 source.n432 1.93989
R746 source.n470 source.n426 1.93989
R747 source.n390 source.n366 1.93989
R748 source.n404 source.n360 1.93989
R749 source.n316 source.n292 1.93989
R750 source.n330 source.n286 1.93989
R751 source.n50 source.n6 1.93989
R752 source.n37 source.n13 1.93989
R753 source.n124 source.n80 1.93989
R754 source.n111 source.n87 1.93989
R755 source.n190 source.n146 1.93989
R756 source.n177 source.n153 1.93989
R757 source.n264 source.n220 1.93989
R758 source.n251 source.n227 1.93989
R759 source.n492 source.t0 1.6505
R760 source.n492 source.t1 1.6505
R761 source.n490 source.t13 1.6505
R762 source.n490 source.t4 1.6505
R763 source.n488 source.t5 1.6505
R764 source.n488 source.t6 1.6505
R765 source.n486 source.t8 1.6505
R766 source.n486 source.t14 1.6505
R767 source.n352 source.t29 1.6505
R768 source.n352 source.t32 1.6505
R769 source.n350 source.t25 1.6505
R770 source.n350 source.t21 1.6505
R771 source.n348 source.t19 1.6505
R772 source.n348 source.t37 1.6505
R773 source.n346 source.t30 1.6505
R774 source.n346 source.t31 1.6505
R775 source.n66 source.t22 1.6505
R776 source.n66 source.t20 1.6505
R777 source.n68 source.t33 1.6505
R778 source.n68 source.t36 1.6505
R779 source.n70 source.t24 1.6505
R780 source.n70 source.t35 1.6505
R781 source.n72 source.t28 1.6505
R782 source.n72 source.t23 1.6505
R783 source.n206 source.t3 1.6505
R784 source.n206 source.t9 1.6505
R785 source.n208 source.t12 1.6505
R786 source.n208 source.t15 1.6505
R787 source.n210 source.t17 1.6505
R788 source.n210 source.t11 1.6505
R789 source.n212 source.t38 1.6505
R790 source.n212 source.t10 1.6505
R791 source.n535 source.n533 1.16414
R792 source.n543 source.n502 1.16414
R793 source.n461 source.n459 1.16414
R794 source.n469 source.n428 1.16414
R795 source.n395 source.n393 1.16414
R796 source.n403 source.n362 1.16414
R797 source.n321 source.n319 1.16414
R798 source.n329 source.n288 1.16414
R799 source.n49 source.n8 1.16414
R800 source.n41 source.n40 1.16414
R801 source.n123 source.n82 1.16414
R802 source.n115 source.n114 1.16414
R803 source.n189 source.n148 1.16414
R804 source.n181 source.n180 1.16414
R805 source.n263 source.n222 1.16414
R806 source.n255 source.n254 1.16414
R807 source.n279 source.n213 0.5005
R808 source.n213 source.n211 0.5005
R809 source.n211 source.n209 0.5005
R810 source.n209 source.n207 0.5005
R811 source.n207 source.n205 0.5005
R812 source.n139 source.n73 0.5005
R813 source.n73 source.n71 0.5005
R814 source.n71 source.n69 0.5005
R815 source.n69 source.n67 0.5005
R816 source.n67 source.n65 0.5005
R817 source.n347 source.n345 0.5005
R818 source.n349 source.n347 0.5005
R819 source.n351 source.n349 0.5005
R820 source.n353 source.n351 0.5005
R821 source.n419 source.n353 0.5005
R822 source.n487 source.n485 0.5005
R823 source.n489 source.n487 0.5005
R824 source.n491 source.n489 0.5005
R825 source.n493 source.n491 0.5005
R826 source.n559 source.n493 0.5005
R827 source.n205 source.n139 0.470328
R828 source.n485 source.n419 0.470328
R829 source.n534 source.n504 0.388379
R830 source.n540 source.n539 0.388379
R831 source.n460 source.n430 0.388379
R832 source.n466 source.n465 0.388379
R833 source.n394 source.n364 0.388379
R834 source.n400 source.n399 0.388379
R835 source.n320 source.n290 0.388379
R836 source.n326 source.n325 0.388379
R837 source.n46 source.n45 0.388379
R838 source.n12 source.n10 0.388379
R839 source.n120 source.n119 0.388379
R840 source.n86 source.n84 0.388379
R841 source.n186 source.n185 0.388379
R842 source.n152 source.n150 0.388379
R843 source.n260 source.n259 0.388379
R844 source.n226 source.n224 0.388379
R845 source source.n560 0.188
R846 source.n516 source.n511 0.155672
R847 source.n523 source.n511 0.155672
R848 source.n524 source.n523 0.155672
R849 source.n524 source.n507 0.155672
R850 source.n531 source.n507 0.155672
R851 source.n532 source.n531 0.155672
R852 source.n532 source.n503 0.155672
R853 source.n541 source.n503 0.155672
R854 source.n542 source.n541 0.155672
R855 source.n542 source.n499 0.155672
R856 source.n549 source.n499 0.155672
R857 source.n550 source.n549 0.155672
R858 source.n550 source.n495 0.155672
R859 source.n557 source.n495 0.155672
R860 source.n442 source.n437 0.155672
R861 source.n449 source.n437 0.155672
R862 source.n450 source.n449 0.155672
R863 source.n450 source.n433 0.155672
R864 source.n457 source.n433 0.155672
R865 source.n458 source.n457 0.155672
R866 source.n458 source.n429 0.155672
R867 source.n467 source.n429 0.155672
R868 source.n468 source.n467 0.155672
R869 source.n468 source.n425 0.155672
R870 source.n475 source.n425 0.155672
R871 source.n476 source.n475 0.155672
R872 source.n476 source.n421 0.155672
R873 source.n483 source.n421 0.155672
R874 source.n376 source.n371 0.155672
R875 source.n383 source.n371 0.155672
R876 source.n384 source.n383 0.155672
R877 source.n384 source.n367 0.155672
R878 source.n391 source.n367 0.155672
R879 source.n392 source.n391 0.155672
R880 source.n392 source.n363 0.155672
R881 source.n401 source.n363 0.155672
R882 source.n402 source.n401 0.155672
R883 source.n402 source.n359 0.155672
R884 source.n409 source.n359 0.155672
R885 source.n410 source.n409 0.155672
R886 source.n410 source.n355 0.155672
R887 source.n417 source.n355 0.155672
R888 source.n302 source.n297 0.155672
R889 source.n309 source.n297 0.155672
R890 source.n310 source.n309 0.155672
R891 source.n310 source.n293 0.155672
R892 source.n317 source.n293 0.155672
R893 source.n318 source.n317 0.155672
R894 source.n318 source.n289 0.155672
R895 source.n327 source.n289 0.155672
R896 source.n328 source.n327 0.155672
R897 source.n328 source.n285 0.155672
R898 source.n335 source.n285 0.155672
R899 source.n336 source.n335 0.155672
R900 source.n336 source.n281 0.155672
R901 source.n343 source.n281 0.155672
R902 source.n63 source.n1 0.155672
R903 source.n56 source.n1 0.155672
R904 source.n56 source.n55 0.155672
R905 source.n55 source.n5 0.155672
R906 source.n48 source.n5 0.155672
R907 source.n48 source.n47 0.155672
R908 source.n47 source.n9 0.155672
R909 source.n39 source.n9 0.155672
R910 source.n39 source.n38 0.155672
R911 source.n38 source.n14 0.155672
R912 source.n31 source.n14 0.155672
R913 source.n31 source.n30 0.155672
R914 source.n30 source.n18 0.155672
R915 source.n23 source.n18 0.155672
R916 source.n137 source.n75 0.155672
R917 source.n130 source.n75 0.155672
R918 source.n130 source.n129 0.155672
R919 source.n129 source.n79 0.155672
R920 source.n122 source.n79 0.155672
R921 source.n122 source.n121 0.155672
R922 source.n121 source.n83 0.155672
R923 source.n113 source.n83 0.155672
R924 source.n113 source.n112 0.155672
R925 source.n112 source.n88 0.155672
R926 source.n105 source.n88 0.155672
R927 source.n105 source.n104 0.155672
R928 source.n104 source.n92 0.155672
R929 source.n97 source.n92 0.155672
R930 source.n203 source.n141 0.155672
R931 source.n196 source.n141 0.155672
R932 source.n196 source.n195 0.155672
R933 source.n195 source.n145 0.155672
R934 source.n188 source.n145 0.155672
R935 source.n188 source.n187 0.155672
R936 source.n187 source.n149 0.155672
R937 source.n179 source.n149 0.155672
R938 source.n179 source.n178 0.155672
R939 source.n178 source.n154 0.155672
R940 source.n171 source.n154 0.155672
R941 source.n171 source.n170 0.155672
R942 source.n170 source.n158 0.155672
R943 source.n163 source.n158 0.155672
R944 source.n277 source.n215 0.155672
R945 source.n270 source.n215 0.155672
R946 source.n270 source.n269 0.155672
R947 source.n269 source.n219 0.155672
R948 source.n262 source.n219 0.155672
R949 source.n262 source.n261 0.155672
R950 source.n261 source.n223 0.155672
R951 source.n253 source.n223 0.155672
R952 source.n253 source.n252 0.155672
R953 source.n252 source.n228 0.155672
R954 source.n245 source.n228 0.155672
R955 source.n245 source.n244 0.155672
R956 source.n244 source.n232 0.155672
R957 source.n237 source.n232 0.155672
R958 drain_left.n10 drain_left.n8 60.0527
R959 drain_left.n6 drain_left.n4 60.0525
R960 drain_left.n2 drain_left.n0 60.0525
R961 drain_left.n14 drain_left.n13 59.5527
R962 drain_left.n12 drain_left.n11 59.5527
R963 drain_left.n10 drain_left.n9 59.5527
R964 drain_left.n7 drain_left.n3 59.5525
R965 drain_left.n6 drain_left.n5 59.5525
R966 drain_left.n2 drain_left.n1 59.5525
R967 drain_left.n16 drain_left.n15 59.5525
R968 drain_left drain_left.n7 31.3671
R969 drain_left drain_left.n16 6.15322
R970 drain_left.n3 drain_left.t3 1.6505
R971 drain_left.n3 drain_left.t15 1.6505
R972 drain_left.n4 drain_left.t5 1.6505
R973 drain_left.n4 drain_left.t2 1.6505
R974 drain_left.n5 drain_left.t0 1.6505
R975 drain_left.n5 drain_left.t12 1.6505
R976 drain_left.n1 drain_left.t13 1.6505
R977 drain_left.n1 drain_left.t6 1.6505
R978 drain_left.n0 drain_left.t8 1.6505
R979 drain_left.n0 drain_left.t4 1.6505
R980 drain_left.n15 drain_left.t7 1.6505
R981 drain_left.n15 drain_left.t17 1.6505
R982 drain_left.n13 drain_left.t11 1.6505
R983 drain_left.n13 drain_left.t16 1.6505
R984 drain_left.n11 drain_left.t10 1.6505
R985 drain_left.n11 drain_left.t1 1.6505
R986 drain_left.n9 drain_left.t9 1.6505
R987 drain_left.n9 drain_left.t19 1.6505
R988 drain_left.n8 drain_left.t14 1.6505
R989 drain_left.n8 drain_left.t18 1.6505
R990 drain_left.n12 drain_left.n10 0.5005
R991 drain_left.n14 drain_left.n12 0.5005
R992 drain_left.n16 drain_left.n14 0.5005
R993 drain_left.n7 drain_left.n6 0.445154
R994 drain_left.n7 drain_left.n2 0.445154
R995 minus.n25 minus.t7 1334.7
R996 minus.n6 minus.t10 1334.7
R997 minus.n52 minus.t3 1334.7
R998 minus.n33 minus.t19 1334.7
R999 minus.n24 minus.t17 1282.12
R1000 minus.n22 minus.t5 1282.12
R1001 minus.n1 minus.t16 1282.12
R1002 minus.n17 minus.t6 1282.12
R1003 minus.n3 minus.t15 1282.12
R1004 minus.n11 minus.t0 1282.12
R1005 minus.n9 minus.t9 1282.12
R1006 minus.n5 minus.t1 1282.12
R1007 minus.n51 minus.t8 1282.12
R1008 minus.n49 minus.t12 1282.12
R1009 minus.n28 minus.t13 1282.12
R1010 minus.n44 minus.t18 1282.12
R1011 minus.n30 minus.t4 1282.12
R1012 minus.n38 minus.t11 1282.12
R1013 minus.n36 minus.t14 1282.12
R1014 minus.n32 minus.t2 1282.12
R1015 minus.n7 minus.n6 161.489
R1016 minus.n34 minus.n33 161.489
R1017 minus.n26 minus.n25 161.3
R1018 minus.n23 minus.n0 161.3
R1019 minus.n21 minus.n20 161.3
R1020 minus.n19 minus.n18 161.3
R1021 minus.n16 minus.n2 161.3
R1022 minus.n15 minus.n14 161.3
R1023 minus.n13 minus.n12 161.3
R1024 minus.n10 minus.n4 161.3
R1025 minus.n8 minus.n7 161.3
R1026 minus.n53 minus.n52 161.3
R1027 minus.n50 minus.n27 161.3
R1028 minus.n48 minus.n47 161.3
R1029 minus.n46 minus.n45 161.3
R1030 minus.n43 minus.n29 161.3
R1031 minus.n42 minus.n41 161.3
R1032 minus.n40 minus.n39 161.3
R1033 minus.n37 minus.n31 161.3
R1034 minus.n35 minus.n34 161.3
R1035 minus.n16 minus.n15 73.0308
R1036 minus.n43 minus.n42 73.0308
R1037 minus.n18 minus.n17 67.1884
R1038 minus.n12 minus.n3 67.1884
R1039 minus.n39 minus.n30 67.1884
R1040 minus.n45 minus.n44 67.1884
R1041 minus.n21 minus.n1 55.5035
R1042 minus.n11 minus.n10 55.5035
R1043 minus.n38 minus.n37 55.5035
R1044 minus.n48 minus.n28 55.5035
R1045 minus.n23 minus.n22 43.8187
R1046 minus.n9 minus.n8 43.8187
R1047 minus.n36 minus.n35 43.8187
R1048 minus.n50 minus.n49 43.8187
R1049 minus.n24 minus.n23 40.8975
R1050 minus.n8 minus.n5 40.8975
R1051 minus.n35 minus.n32 40.8975
R1052 minus.n51 minus.n50 40.8975
R1053 minus.n54 minus.n26 36.6634
R1054 minus.n25 minus.n24 32.1338
R1055 minus.n6 minus.n5 32.1338
R1056 minus.n33 minus.n32 32.1338
R1057 minus.n52 minus.n51 32.1338
R1058 minus.n22 minus.n21 29.2126
R1059 minus.n10 minus.n9 29.2126
R1060 minus.n37 minus.n36 29.2126
R1061 minus.n49 minus.n48 29.2126
R1062 minus.n18 minus.n1 17.5278
R1063 minus.n12 minus.n11 17.5278
R1064 minus.n39 minus.n38 17.5278
R1065 minus.n45 minus.n28 17.5278
R1066 minus.n54 minus.n53 6.49671
R1067 minus.n17 minus.n16 5.84292
R1068 minus.n15 minus.n3 5.84292
R1069 minus.n42 minus.n30 5.84292
R1070 minus.n44 minus.n43 5.84292
R1071 minus.n26 minus.n0 0.189894
R1072 minus.n20 minus.n0 0.189894
R1073 minus.n20 minus.n19 0.189894
R1074 minus.n19 minus.n2 0.189894
R1075 minus.n14 minus.n2 0.189894
R1076 minus.n14 minus.n13 0.189894
R1077 minus.n13 minus.n4 0.189894
R1078 minus.n7 minus.n4 0.189894
R1079 minus.n34 minus.n31 0.189894
R1080 minus.n40 minus.n31 0.189894
R1081 minus.n41 minus.n40 0.189894
R1082 minus.n41 minus.n29 0.189894
R1083 minus.n46 minus.n29 0.189894
R1084 minus.n47 minus.n46 0.189894
R1085 minus.n47 minus.n27 0.189894
R1086 minus.n53 minus.n27 0.189894
R1087 minus minus.n54 0.188
R1088 drain_right.n6 drain_right.n4 60.0525
R1089 drain_right.n2 drain_right.n0 60.0525
R1090 drain_right.n10 drain_right.n8 60.0525
R1091 drain_right.n10 drain_right.n9 59.5527
R1092 drain_right.n12 drain_right.n11 59.5527
R1093 drain_right.n14 drain_right.n13 59.5527
R1094 drain_right.n16 drain_right.n15 59.5527
R1095 drain_right.n7 drain_right.n3 59.5525
R1096 drain_right.n6 drain_right.n5 59.5525
R1097 drain_right.n2 drain_right.n1 59.5525
R1098 drain_right drain_right.n7 30.8138
R1099 drain_right drain_right.n16 6.15322
R1100 drain_right.n3 drain_right.t15 1.6505
R1101 drain_right.n3 drain_right.t1 1.6505
R1102 drain_right.n4 drain_right.t11 1.6505
R1103 drain_right.n4 drain_right.t16 1.6505
R1104 drain_right.n5 drain_right.t6 1.6505
R1105 drain_right.n5 drain_right.t7 1.6505
R1106 drain_right.n1 drain_right.t5 1.6505
R1107 drain_right.n1 drain_right.t8 1.6505
R1108 drain_right.n0 drain_right.t0 1.6505
R1109 drain_right.n0 drain_right.t17 1.6505
R1110 drain_right.n8 drain_right.t18 1.6505
R1111 drain_right.n8 drain_right.t9 1.6505
R1112 drain_right.n9 drain_right.t19 1.6505
R1113 drain_right.n9 drain_right.t10 1.6505
R1114 drain_right.n11 drain_right.t13 1.6505
R1115 drain_right.n11 drain_right.t4 1.6505
R1116 drain_right.n13 drain_right.t14 1.6505
R1117 drain_right.n13 drain_right.t3 1.6505
R1118 drain_right.n15 drain_right.t12 1.6505
R1119 drain_right.n15 drain_right.t2 1.6505
R1120 drain_right.n16 drain_right.n14 0.5005
R1121 drain_right.n14 drain_right.n12 0.5005
R1122 drain_right.n12 drain_right.n10 0.5005
R1123 drain_right.n7 drain_right.n6 0.445154
R1124 drain_right.n7 drain_right.n2 0.445154
C0 drain_right plus 0.349242f
C1 minus drain_left 0.171712f
C2 minus source 5.97207f
C3 source drain_left 40.8896f
C4 minus plus 5.63806f
C5 plus drain_left 6.46495f
C6 source plus 5.98611f
C7 drain_right minus 6.27045f
C8 drain_right drain_left 1.04652f
C9 drain_right source 40.8898f
C10 drain_right a_n1992_n3288# 7.0112f
C11 drain_left a_n1992_n3288# 7.32112f
C12 source a_n1992_n3288# 8.7117f
C13 minus a_n1992_n3288# 7.776731f
C14 plus a_n1992_n3288# 9.83018f
C15 drain_right.t0 a_n1992_n3288# 0.343273f
C16 drain_right.t17 a_n1992_n3288# 0.343273f
C17 drain_right.n0 a_n1992_n3288# 3.05822f
C18 drain_right.t5 a_n1992_n3288# 0.343273f
C19 drain_right.t8 a_n1992_n3288# 0.343273f
C20 drain_right.n1 a_n1992_n3288# 3.0546f
C21 drain_right.n2 a_n1992_n3288# 0.847292f
C22 drain_right.t15 a_n1992_n3288# 0.343273f
C23 drain_right.t1 a_n1992_n3288# 0.343273f
C24 drain_right.n3 a_n1992_n3288# 3.0546f
C25 drain_right.t11 a_n1992_n3288# 0.343273f
C26 drain_right.t16 a_n1992_n3288# 0.343273f
C27 drain_right.n4 a_n1992_n3288# 3.05822f
C28 drain_right.t6 a_n1992_n3288# 0.343273f
C29 drain_right.t7 a_n1992_n3288# 0.343273f
C30 drain_right.n5 a_n1992_n3288# 3.0546f
C31 drain_right.n6 a_n1992_n3288# 0.847292f
C32 drain_right.n7 a_n1992_n3288# 2.11523f
C33 drain_right.t18 a_n1992_n3288# 0.343273f
C34 drain_right.t9 a_n1992_n3288# 0.343273f
C35 drain_right.n8 a_n1992_n3288# 3.05822f
C36 drain_right.t19 a_n1992_n3288# 0.343273f
C37 drain_right.t10 a_n1992_n3288# 0.343273f
C38 drain_right.n9 a_n1992_n3288# 3.05461f
C39 drain_right.n10 a_n1992_n3288# 0.851848f
C40 drain_right.t13 a_n1992_n3288# 0.343273f
C41 drain_right.t4 a_n1992_n3288# 0.343273f
C42 drain_right.n11 a_n1992_n3288# 3.05461f
C43 drain_right.n12 a_n1992_n3288# 0.420439f
C44 drain_right.t14 a_n1992_n3288# 0.343273f
C45 drain_right.t3 a_n1992_n3288# 0.343273f
C46 drain_right.n13 a_n1992_n3288# 3.05461f
C47 drain_right.n14 a_n1992_n3288# 0.420439f
C48 drain_right.t12 a_n1992_n3288# 0.343273f
C49 drain_right.t2 a_n1992_n3288# 0.343273f
C50 drain_right.n15 a_n1992_n3288# 3.05461f
C51 drain_right.n16 a_n1992_n3288# 0.719242f
C52 minus.n0 a_n1992_n3288# 0.050969f
C53 minus.t7 a_n1992_n3288# 0.439082f
C54 minus.t17 a_n1992_n3288# 0.43209f
C55 minus.t5 a_n1992_n3288# 0.43209f
C56 minus.t16 a_n1992_n3288# 0.43209f
C57 minus.n1 a_n1992_n3288# 0.174026f
C58 minus.n2 a_n1992_n3288# 0.050969f
C59 minus.t6 a_n1992_n3288# 0.43209f
C60 minus.t15 a_n1992_n3288# 0.43209f
C61 minus.n3 a_n1992_n3288# 0.174026f
C62 minus.n4 a_n1992_n3288# 0.050969f
C63 minus.t0 a_n1992_n3288# 0.43209f
C64 minus.t9 a_n1992_n3288# 0.43209f
C65 minus.t1 a_n1992_n3288# 0.43209f
C66 minus.n5 a_n1992_n3288# 0.174026f
C67 minus.t10 a_n1992_n3288# 0.439082f
C68 minus.n6 a_n1992_n3288# 0.18999f
C69 minus.n7 a_n1992_n3288# 0.116631f
C70 minus.n8 a_n1992_n3288# 0.019422f
C71 minus.n9 a_n1992_n3288# 0.174026f
C72 minus.n10 a_n1992_n3288# 0.019422f
C73 minus.n11 a_n1992_n3288# 0.174026f
C74 minus.n12 a_n1992_n3288# 0.019422f
C75 minus.n13 a_n1992_n3288# 0.050969f
C76 minus.n14 a_n1992_n3288# 0.050969f
C77 minus.n15 a_n1992_n3288# 0.018165f
C78 minus.n16 a_n1992_n3288# 0.018165f
C79 minus.n17 a_n1992_n3288# 0.174026f
C80 minus.n18 a_n1992_n3288# 0.019422f
C81 minus.n19 a_n1992_n3288# 0.050969f
C82 minus.n20 a_n1992_n3288# 0.050969f
C83 minus.n21 a_n1992_n3288# 0.019422f
C84 minus.n22 a_n1992_n3288# 0.174026f
C85 minus.n23 a_n1992_n3288# 0.019422f
C86 minus.n24 a_n1992_n3288# 0.174026f
C87 minus.n25 a_n1992_n3288# 0.189913f
C88 minus.n26 a_n1992_n3288# 1.83775f
C89 minus.n27 a_n1992_n3288# 0.050969f
C90 minus.t8 a_n1992_n3288# 0.43209f
C91 minus.t12 a_n1992_n3288# 0.43209f
C92 minus.t13 a_n1992_n3288# 0.43209f
C93 minus.n28 a_n1992_n3288# 0.174026f
C94 minus.n29 a_n1992_n3288# 0.050969f
C95 minus.t18 a_n1992_n3288# 0.43209f
C96 minus.t4 a_n1992_n3288# 0.43209f
C97 minus.n30 a_n1992_n3288# 0.174026f
C98 minus.n31 a_n1992_n3288# 0.050969f
C99 minus.t11 a_n1992_n3288# 0.43209f
C100 minus.t14 a_n1992_n3288# 0.43209f
C101 minus.t2 a_n1992_n3288# 0.43209f
C102 minus.n32 a_n1992_n3288# 0.174026f
C103 minus.t19 a_n1992_n3288# 0.439082f
C104 minus.n33 a_n1992_n3288# 0.18999f
C105 minus.n34 a_n1992_n3288# 0.116631f
C106 minus.n35 a_n1992_n3288# 0.019422f
C107 minus.n36 a_n1992_n3288# 0.174026f
C108 minus.n37 a_n1992_n3288# 0.019422f
C109 minus.n38 a_n1992_n3288# 0.174026f
C110 minus.n39 a_n1992_n3288# 0.019422f
C111 minus.n40 a_n1992_n3288# 0.050969f
C112 minus.n41 a_n1992_n3288# 0.050969f
C113 minus.n42 a_n1992_n3288# 0.018165f
C114 minus.n43 a_n1992_n3288# 0.018165f
C115 minus.n44 a_n1992_n3288# 0.174026f
C116 minus.n45 a_n1992_n3288# 0.019422f
C117 minus.n46 a_n1992_n3288# 0.050969f
C118 minus.n47 a_n1992_n3288# 0.050969f
C119 minus.n48 a_n1992_n3288# 0.019422f
C120 minus.n49 a_n1992_n3288# 0.174026f
C121 minus.n50 a_n1992_n3288# 0.019422f
C122 minus.n51 a_n1992_n3288# 0.174026f
C123 minus.t3 a_n1992_n3288# 0.439082f
C124 minus.n52 a_n1992_n3288# 0.189913f
C125 minus.n53 a_n1992_n3288# 0.332829f
C126 minus.n54 a_n1992_n3288# 2.22939f
C127 drain_left.t8 a_n1992_n3288# 0.343696f
C128 drain_left.t4 a_n1992_n3288# 0.343696f
C129 drain_left.n0 a_n1992_n3288# 3.06199f
C130 drain_left.t13 a_n1992_n3288# 0.343696f
C131 drain_left.t6 a_n1992_n3288# 0.343696f
C132 drain_left.n1 a_n1992_n3288# 3.05837f
C133 drain_left.n2 a_n1992_n3288# 0.848338f
C134 drain_left.t3 a_n1992_n3288# 0.343696f
C135 drain_left.t15 a_n1992_n3288# 0.343696f
C136 drain_left.n3 a_n1992_n3288# 3.05837f
C137 drain_left.t5 a_n1992_n3288# 0.343696f
C138 drain_left.t2 a_n1992_n3288# 0.343696f
C139 drain_left.n4 a_n1992_n3288# 3.06199f
C140 drain_left.t0 a_n1992_n3288# 0.343696f
C141 drain_left.t12 a_n1992_n3288# 0.343696f
C142 drain_left.n5 a_n1992_n3288# 3.05837f
C143 drain_left.n6 a_n1992_n3288# 0.848338f
C144 drain_left.n7 a_n1992_n3288# 2.19281f
C145 drain_left.t14 a_n1992_n3288# 0.343696f
C146 drain_left.t18 a_n1992_n3288# 0.343696f
C147 drain_left.n8 a_n1992_n3288# 3.06201f
C148 drain_left.t9 a_n1992_n3288# 0.343696f
C149 drain_left.t19 a_n1992_n3288# 0.343696f
C150 drain_left.n9 a_n1992_n3288# 3.05838f
C151 drain_left.n10 a_n1992_n3288# 0.852886f
C152 drain_left.t10 a_n1992_n3288# 0.343696f
C153 drain_left.t1 a_n1992_n3288# 0.343696f
C154 drain_left.n11 a_n1992_n3288# 3.05838f
C155 drain_left.n12 a_n1992_n3288# 0.420957f
C156 drain_left.t11 a_n1992_n3288# 0.343696f
C157 drain_left.t16 a_n1992_n3288# 0.343696f
C158 drain_left.n13 a_n1992_n3288# 3.05838f
C159 drain_left.n14 a_n1992_n3288# 0.420957f
C160 drain_left.t7 a_n1992_n3288# 0.343696f
C161 drain_left.t17 a_n1992_n3288# 0.343696f
C162 drain_left.n15 a_n1992_n3288# 3.05837f
C163 drain_left.n16 a_n1992_n3288# 0.720142f
C164 source.n0 a_n1992_n3288# 0.041549f
C165 source.n1 a_n1992_n3288# 0.031366f
C166 source.n2 a_n1992_n3288# 0.016855f
C167 source.n3 a_n1992_n3288# 0.039839f
C168 source.n4 a_n1992_n3288# 0.017846f
C169 source.n5 a_n1992_n3288# 0.031366f
C170 source.n6 a_n1992_n3288# 0.016855f
C171 source.n7 a_n1992_n3288# 0.039839f
C172 source.n8 a_n1992_n3288# 0.017846f
C173 source.n9 a_n1992_n3288# 0.031366f
C174 source.n10 a_n1992_n3288# 0.017351f
C175 source.n11 a_n1992_n3288# 0.039839f
C176 source.n12 a_n1992_n3288# 0.016855f
C177 source.n13 a_n1992_n3288# 0.017846f
C178 source.n14 a_n1992_n3288# 0.031366f
C179 source.n15 a_n1992_n3288# 0.016855f
C180 source.n16 a_n1992_n3288# 0.039839f
C181 source.n17 a_n1992_n3288# 0.017846f
C182 source.n18 a_n1992_n3288# 0.031366f
C183 source.n19 a_n1992_n3288# 0.016855f
C184 source.n20 a_n1992_n3288# 0.029879f
C185 source.n21 a_n1992_n3288# 0.028163f
C186 source.t34 a_n1992_n3288# 0.067285f
C187 source.n22 a_n1992_n3288# 0.226147f
C188 source.n23 a_n1992_n3288# 1.58237f
C189 source.n24 a_n1992_n3288# 0.016855f
C190 source.n25 a_n1992_n3288# 0.017846f
C191 source.n26 a_n1992_n3288# 0.039839f
C192 source.n27 a_n1992_n3288# 0.039839f
C193 source.n28 a_n1992_n3288# 0.017846f
C194 source.n29 a_n1992_n3288# 0.016855f
C195 source.n30 a_n1992_n3288# 0.031366f
C196 source.n31 a_n1992_n3288# 0.031366f
C197 source.n32 a_n1992_n3288# 0.016855f
C198 source.n33 a_n1992_n3288# 0.017846f
C199 source.n34 a_n1992_n3288# 0.039839f
C200 source.n35 a_n1992_n3288# 0.039839f
C201 source.n36 a_n1992_n3288# 0.017846f
C202 source.n37 a_n1992_n3288# 0.016855f
C203 source.n38 a_n1992_n3288# 0.031366f
C204 source.n39 a_n1992_n3288# 0.031366f
C205 source.n40 a_n1992_n3288# 0.016855f
C206 source.n41 a_n1992_n3288# 0.017846f
C207 source.n42 a_n1992_n3288# 0.039839f
C208 source.n43 a_n1992_n3288# 0.039839f
C209 source.n44 a_n1992_n3288# 0.039839f
C210 source.n45 a_n1992_n3288# 0.017351f
C211 source.n46 a_n1992_n3288# 0.016855f
C212 source.n47 a_n1992_n3288# 0.031366f
C213 source.n48 a_n1992_n3288# 0.031366f
C214 source.n49 a_n1992_n3288# 0.016855f
C215 source.n50 a_n1992_n3288# 0.017846f
C216 source.n51 a_n1992_n3288# 0.039839f
C217 source.n52 a_n1992_n3288# 0.039839f
C218 source.n53 a_n1992_n3288# 0.017846f
C219 source.n54 a_n1992_n3288# 0.016855f
C220 source.n55 a_n1992_n3288# 0.031366f
C221 source.n56 a_n1992_n3288# 0.031366f
C222 source.n57 a_n1992_n3288# 0.016855f
C223 source.n58 a_n1992_n3288# 0.017846f
C224 source.n59 a_n1992_n3288# 0.039839f
C225 source.n60 a_n1992_n3288# 0.081753f
C226 source.n61 a_n1992_n3288# 0.017846f
C227 source.n62 a_n1992_n3288# 0.016855f
C228 source.n63 a_n1992_n3288# 0.06736f
C229 source.n64 a_n1992_n3288# 0.045119f
C230 source.n65 a_n1992_n3288# 1.25518f
C231 source.t22 a_n1992_n3288# 0.297438f
C232 source.t20 a_n1992_n3288# 0.297438f
C233 source.n66 a_n1992_n3288# 2.54667f
C234 source.n67 a_n1992_n3288# 0.421748f
C235 source.t33 a_n1992_n3288# 0.297438f
C236 source.t36 a_n1992_n3288# 0.297438f
C237 source.n68 a_n1992_n3288# 2.54667f
C238 source.n69 a_n1992_n3288# 0.421748f
C239 source.t24 a_n1992_n3288# 0.297438f
C240 source.t35 a_n1992_n3288# 0.297438f
C241 source.n70 a_n1992_n3288# 2.54667f
C242 source.n71 a_n1992_n3288# 0.421748f
C243 source.t28 a_n1992_n3288# 0.297438f
C244 source.t23 a_n1992_n3288# 0.297438f
C245 source.n72 a_n1992_n3288# 2.54667f
C246 source.n73 a_n1992_n3288# 0.421748f
C247 source.n74 a_n1992_n3288# 0.041549f
C248 source.n75 a_n1992_n3288# 0.031366f
C249 source.n76 a_n1992_n3288# 0.016855f
C250 source.n77 a_n1992_n3288# 0.039839f
C251 source.n78 a_n1992_n3288# 0.017846f
C252 source.n79 a_n1992_n3288# 0.031366f
C253 source.n80 a_n1992_n3288# 0.016855f
C254 source.n81 a_n1992_n3288# 0.039839f
C255 source.n82 a_n1992_n3288# 0.017846f
C256 source.n83 a_n1992_n3288# 0.031366f
C257 source.n84 a_n1992_n3288# 0.017351f
C258 source.n85 a_n1992_n3288# 0.039839f
C259 source.n86 a_n1992_n3288# 0.016855f
C260 source.n87 a_n1992_n3288# 0.017846f
C261 source.n88 a_n1992_n3288# 0.031366f
C262 source.n89 a_n1992_n3288# 0.016855f
C263 source.n90 a_n1992_n3288# 0.039839f
C264 source.n91 a_n1992_n3288# 0.017846f
C265 source.n92 a_n1992_n3288# 0.031366f
C266 source.n93 a_n1992_n3288# 0.016855f
C267 source.n94 a_n1992_n3288# 0.029879f
C268 source.n95 a_n1992_n3288# 0.028163f
C269 source.t18 a_n1992_n3288# 0.067285f
C270 source.n96 a_n1992_n3288# 0.226147f
C271 source.n97 a_n1992_n3288# 1.58237f
C272 source.n98 a_n1992_n3288# 0.016855f
C273 source.n99 a_n1992_n3288# 0.017846f
C274 source.n100 a_n1992_n3288# 0.039839f
C275 source.n101 a_n1992_n3288# 0.039839f
C276 source.n102 a_n1992_n3288# 0.017846f
C277 source.n103 a_n1992_n3288# 0.016855f
C278 source.n104 a_n1992_n3288# 0.031366f
C279 source.n105 a_n1992_n3288# 0.031366f
C280 source.n106 a_n1992_n3288# 0.016855f
C281 source.n107 a_n1992_n3288# 0.017846f
C282 source.n108 a_n1992_n3288# 0.039839f
C283 source.n109 a_n1992_n3288# 0.039839f
C284 source.n110 a_n1992_n3288# 0.017846f
C285 source.n111 a_n1992_n3288# 0.016855f
C286 source.n112 a_n1992_n3288# 0.031366f
C287 source.n113 a_n1992_n3288# 0.031366f
C288 source.n114 a_n1992_n3288# 0.016855f
C289 source.n115 a_n1992_n3288# 0.017846f
C290 source.n116 a_n1992_n3288# 0.039839f
C291 source.n117 a_n1992_n3288# 0.039839f
C292 source.n118 a_n1992_n3288# 0.039839f
C293 source.n119 a_n1992_n3288# 0.017351f
C294 source.n120 a_n1992_n3288# 0.016855f
C295 source.n121 a_n1992_n3288# 0.031366f
C296 source.n122 a_n1992_n3288# 0.031366f
C297 source.n123 a_n1992_n3288# 0.016855f
C298 source.n124 a_n1992_n3288# 0.017846f
C299 source.n125 a_n1992_n3288# 0.039839f
C300 source.n126 a_n1992_n3288# 0.039839f
C301 source.n127 a_n1992_n3288# 0.017846f
C302 source.n128 a_n1992_n3288# 0.016855f
C303 source.n129 a_n1992_n3288# 0.031366f
C304 source.n130 a_n1992_n3288# 0.031366f
C305 source.n131 a_n1992_n3288# 0.016855f
C306 source.n132 a_n1992_n3288# 0.017846f
C307 source.n133 a_n1992_n3288# 0.039839f
C308 source.n134 a_n1992_n3288# 0.081753f
C309 source.n135 a_n1992_n3288# 0.017846f
C310 source.n136 a_n1992_n3288# 0.016855f
C311 source.n137 a_n1992_n3288# 0.06736f
C312 source.n138 a_n1992_n3288# 0.045119f
C313 source.n139 a_n1992_n3288# 0.121912f
C314 source.n140 a_n1992_n3288# 0.041549f
C315 source.n141 a_n1992_n3288# 0.031366f
C316 source.n142 a_n1992_n3288# 0.016855f
C317 source.n143 a_n1992_n3288# 0.039839f
C318 source.n144 a_n1992_n3288# 0.017846f
C319 source.n145 a_n1992_n3288# 0.031366f
C320 source.n146 a_n1992_n3288# 0.016855f
C321 source.n147 a_n1992_n3288# 0.039839f
C322 source.n148 a_n1992_n3288# 0.017846f
C323 source.n149 a_n1992_n3288# 0.031366f
C324 source.n150 a_n1992_n3288# 0.017351f
C325 source.n151 a_n1992_n3288# 0.039839f
C326 source.n152 a_n1992_n3288# 0.016855f
C327 source.n153 a_n1992_n3288# 0.017846f
C328 source.n154 a_n1992_n3288# 0.031366f
C329 source.n155 a_n1992_n3288# 0.016855f
C330 source.n156 a_n1992_n3288# 0.039839f
C331 source.n157 a_n1992_n3288# 0.017846f
C332 source.n158 a_n1992_n3288# 0.031366f
C333 source.n159 a_n1992_n3288# 0.016855f
C334 source.n160 a_n1992_n3288# 0.029879f
C335 source.n161 a_n1992_n3288# 0.028163f
C336 source.t39 a_n1992_n3288# 0.067285f
C337 source.n162 a_n1992_n3288# 0.226147f
C338 source.n163 a_n1992_n3288# 1.58237f
C339 source.n164 a_n1992_n3288# 0.016855f
C340 source.n165 a_n1992_n3288# 0.017846f
C341 source.n166 a_n1992_n3288# 0.039839f
C342 source.n167 a_n1992_n3288# 0.039839f
C343 source.n168 a_n1992_n3288# 0.017846f
C344 source.n169 a_n1992_n3288# 0.016855f
C345 source.n170 a_n1992_n3288# 0.031366f
C346 source.n171 a_n1992_n3288# 0.031366f
C347 source.n172 a_n1992_n3288# 0.016855f
C348 source.n173 a_n1992_n3288# 0.017846f
C349 source.n174 a_n1992_n3288# 0.039839f
C350 source.n175 a_n1992_n3288# 0.039839f
C351 source.n176 a_n1992_n3288# 0.017846f
C352 source.n177 a_n1992_n3288# 0.016855f
C353 source.n178 a_n1992_n3288# 0.031366f
C354 source.n179 a_n1992_n3288# 0.031366f
C355 source.n180 a_n1992_n3288# 0.016855f
C356 source.n181 a_n1992_n3288# 0.017846f
C357 source.n182 a_n1992_n3288# 0.039839f
C358 source.n183 a_n1992_n3288# 0.039839f
C359 source.n184 a_n1992_n3288# 0.039839f
C360 source.n185 a_n1992_n3288# 0.017351f
C361 source.n186 a_n1992_n3288# 0.016855f
C362 source.n187 a_n1992_n3288# 0.031366f
C363 source.n188 a_n1992_n3288# 0.031366f
C364 source.n189 a_n1992_n3288# 0.016855f
C365 source.n190 a_n1992_n3288# 0.017846f
C366 source.n191 a_n1992_n3288# 0.039839f
C367 source.n192 a_n1992_n3288# 0.039839f
C368 source.n193 a_n1992_n3288# 0.017846f
C369 source.n194 a_n1992_n3288# 0.016855f
C370 source.n195 a_n1992_n3288# 0.031366f
C371 source.n196 a_n1992_n3288# 0.031366f
C372 source.n197 a_n1992_n3288# 0.016855f
C373 source.n198 a_n1992_n3288# 0.017846f
C374 source.n199 a_n1992_n3288# 0.039839f
C375 source.n200 a_n1992_n3288# 0.081753f
C376 source.n201 a_n1992_n3288# 0.017846f
C377 source.n202 a_n1992_n3288# 0.016855f
C378 source.n203 a_n1992_n3288# 0.06736f
C379 source.n204 a_n1992_n3288# 0.045119f
C380 source.n205 a_n1992_n3288# 0.121912f
C381 source.t3 a_n1992_n3288# 0.297438f
C382 source.t9 a_n1992_n3288# 0.297438f
C383 source.n206 a_n1992_n3288# 2.54667f
C384 source.n207 a_n1992_n3288# 0.421748f
C385 source.t12 a_n1992_n3288# 0.297438f
C386 source.t15 a_n1992_n3288# 0.297438f
C387 source.n208 a_n1992_n3288# 2.54667f
C388 source.n209 a_n1992_n3288# 0.421748f
C389 source.t17 a_n1992_n3288# 0.297438f
C390 source.t11 a_n1992_n3288# 0.297438f
C391 source.n210 a_n1992_n3288# 2.54667f
C392 source.n211 a_n1992_n3288# 0.421748f
C393 source.t38 a_n1992_n3288# 0.297438f
C394 source.t10 a_n1992_n3288# 0.297438f
C395 source.n212 a_n1992_n3288# 2.54667f
C396 source.n213 a_n1992_n3288# 0.421748f
C397 source.n214 a_n1992_n3288# 0.041549f
C398 source.n215 a_n1992_n3288# 0.031366f
C399 source.n216 a_n1992_n3288# 0.016855f
C400 source.n217 a_n1992_n3288# 0.039839f
C401 source.n218 a_n1992_n3288# 0.017846f
C402 source.n219 a_n1992_n3288# 0.031366f
C403 source.n220 a_n1992_n3288# 0.016855f
C404 source.n221 a_n1992_n3288# 0.039839f
C405 source.n222 a_n1992_n3288# 0.017846f
C406 source.n223 a_n1992_n3288# 0.031366f
C407 source.n224 a_n1992_n3288# 0.017351f
C408 source.n225 a_n1992_n3288# 0.039839f
C409 source.n226 a_n1992_n3288# 0.016855f
C410 source.n227 a_n1992_n3288# 0.017846f
C411 source.n228 a_n1992_n3288# 0.031366f
C412 source.n229 a_n1992_n3288# 0.016855f
C413 source.n230 a_n1992_n3288# 0.039839f
C414 source.n231 a_n1992_n3288# 0.017846f
C415 source.n232 a_n1992_n3288# 0.031366f
C416 source.n233 a_n1992_n3288# 0.016855f
C417 source.n234 a_n1992_n3288# 0.029879f
C418 source.n235 a_n1992_n3288# 0.028163f
C419 source.t16 a_n1992_n3288# 0.067285f
C420 source.n236 a_n1992_n3288# 0.226147f
C421 source.n237 a_n1992_n3288# 1.58237f
C422 source.n238 a_n1992_n3288# 0.016855f
C423 source.n239 a_n1992_n3288# 0.017846f
C424 source.n240 a_n1992_n3288# 0.039839f
C425 source.n241 a_n1992_n3288# 0.039839f
C426 source.n242 a_n1992_n3288# 0.017846f
C427 source.n243 a_n1992_n3288# 0.016855f
C428 source.n244 a_n1992_n3288# 0.031366f
C429 source.n245 a_n1992_n3288# 0.031366f
C430 source.n246 a_n1992_n3288# 0.016855f
C431 source.n247 a_n1992_n3288# 0.017846f
C432 source.n248 a_n1992_n3288# 0.039839f
C433 source.n249 a_n1992_n3288# 0.039839f
C434 source.n250 a_n1992_n3288# 0.017846f
C435 source.n251 a_n1992_n3288# 0.016855f
C436 source.n252 a_n1992_n3288# 0.031366f
C437 source.n253 a_n1992_n3288# 0.031366f
C438 source.n254 a_n1992_n3288# 0.016855f
C439 source.n255 a_n1992_n3288# 0.017846f
C440 source.n256 a_n1992_n3288# 0.039839f
C441 source.n257 a_n1992_n3288# 0.039839f
C442 source.n258 a_n1992_n3288# 0.039839f
C443 source.n259 a_n1992_n3288# 0.017351f
C444 source.n260 a_n1992_n3288# 0.016855f
C445 source.n261 a_n1992_n3288# 0.031366f
C446 source.n262 a_n1992_n3288# 0.031366f
C447 source.n263 a_n1992_n3288# 0.016855f
C448 source.n264 a_n1992_n3288# 0.017846f
C449 source.n265 a_n1992_n3288# 0.039839f
C450 source.n266 a_n1992_n3288# 0.039839f
C451 source.n267 a_n1992_n3288# 0.017846f
C452 source.n268 a_n1992_n3288# 0.016855f
C453 source.n269 a_n1992_n3288# 0.031366f
C454 source.n270 a_n1992_n3288# 0.031366f
C455 source.n271 a_n1992_n3288# 0.016855f
C456 source.n272 a_n1992_n3288# 0.017846f
C457 source.n273 a_n1992_n3288# 0.039839f
C458 source.n274 a_n1992_n3288# 0.081753f
C459 source.n275 a_n1992_n3288# 0.017846f
C460 source.n276 a_n1992_n3288# 0.016855f
C461 source.n277 a_n1992_n3288# 0.06736f
C462 source.n278 a_n1992_n3288# 0.045119f
C463 source.n279 a_n1992_n3288# 1.74683f
C464 source.n280 a_n1992_n3288# 0.041549f
C465 source.n281 a_n1992_n3288# 0.031366f
C466 source.n282 a_n1992_n3288# 0.016855f
C467 source.n283 a_n1992_n3288# 0.039839f
C468 source.n284 a_n1992_n3288# 0.017846f
C469 source.n285 a_n1992_n3288# 0.031366f
C470 source.n286 a_n1992_n3288# 0.016855f
C471 source.n287 a_n1992_n3288# 0.039839f
C472 source.n288 a_n1992_n3288# 0.017846f
C473 source.n289 a_n1992_n3288# 0.031366f
C474 source.n290 a_n1992_n3288# 0.017351f
C475 source.n291 a_n1992_n3288# 0.039839f
C476 source.n292 a_n1992_n3288# 0.017846f
C477 source.n293 a_n1992_n3288# 0.031366f
C478 source.n294 a_n1992_n3288# 0.016855f
C479 source.n295 a_n1992_n3288# 0.039839f
C480 source.n296 a_n1992_n3288# 0.017846f
C481 source.n297 a_n1992_n3288# 0.031366f
C482 source.n298 a_n1992_n3288# 0.016855f
C483 source.n299 a_n1992_n3288# 0.029879f
C484 source.n300 a_n1992_n3288# 0.028163f
C485 source.t26 a_n1992_n3288# 0.067285f
C486 source.n301 a_n1992_n3288# 0.226147f
C487 source.n302 a_n1992_n3288# 1.58237f
C488 source.n303 a_n1992_n3288# 0.016855f
C489 source.n304 a_n1992_n3288# 0.017846f
C490 source.n305 a_n1992_n3288# 0.039839f
C491 source.n306 a_n1992_n3288# 0.039839f
C492 source.n307 a_n1992_n3288# 0.017846f
C493 source.n308 a_n1992_n3288# 0.016855f
C494 source.n309 a_n1992_n3288# 0.031366f
C495 source.n310 a_n1992_n3288# 0.031366f
C496 source.n311 a_n1992_n3288# 0.016855f
C497 source.n312 a_n1992_n3288# 0.017846f
C498 source.n313 a_n1992_n3288# 0.039839f
C499 source.n314 a_n1992_n3288# 0.039839f
C500 source.n315 a_n1992_n3288# 0.017846f
C501 source.n316 a_n1992_n3288# 0.016855f
C502 source.n317 a_n1992_n3288# 0.031366f
C503 source.n318 a_n1992_n3288# 0.031366f
C504 source.n319 a_n1992_n3288# 0.016855f
C505 source.n320 a_n1992_n3288# 0.016855f
C506 source.n321 a_n1992_n3288# 0.017846f
C507 source.n322 a_n1992_n3288# 0.039839f
C508 source.n323 a_n1992_n3288# 0.039839f
C509 source.n324 a_n1992_n3288# 0.039839f
C510 source.n325 a_n1992_n3288# 0.017351f
C511 source.n326 a_n1992_n3288# 0.016855f
C512 source.n327 a_n1992_n3288# 0.031366f
C513 source.n328 a_n1992_n3288# 0.031366f
C514 source.n329 a_n1992_n3288# 0.016855f
C515 source.n330 a_n1992_n3288# 0.017846f
C516 source.n331 a_n1992_n3288# 0.039839f
C517 source.n332 a_n1992_n3288# 0.039839f
C518 source.n333 a_n1992_n3288# 0.017846f
C519 source.n334 a_n1992_n3288# 0.016855f
C520 source.n335 a_n1992_n3288# 0.031366f
C521 source.n336 a_n1992_n3288# 0.031366f
C522 source.n337 a_n1992_n3288# 0.016855f
C523 source.n338 a_n1992_n3288# 0.017846f
C524 source.n339 a_n1992_n3288# 0.039839f
C525 source.n340 a_n1992_n3288# 0.081753f
C526 source.n341 a_n1992_n3288# 0.017846f
C527 source.n342 a_n1992_n3288# 0.016855f
C528 source.n343 a_n1992_n3288# 0.06736f
C529 source.n344 a_n1992_n3288# 0.045119f
C530 source.n345 a_n1992_n3288# 1.74683f
C531 source.t30 a_n1992_n3288# 0.297438f
C532 source.t31 a_n1992_n3288# 0.297438f
C533 source.n346 a_n1992_n3288# 2.54666f
C534 source.n347 a_n1992_n3288# 0.421764f
C535 source.t19 a_n1992_n3288# 0.297438f
C536 source.t37 a_n1992_n3288# 0.297438f
C537 source.n348 a_n1992_n3288# 2.54666f
C538 source.n349 a_n1992_n3288# 0.421764f
C539 source.t25 a_n1992_n3288# 0.297438f
C540 source.t21 a_n1992_n3288# 0.297438f
C541 source.n350 a_n1992_n3288# 2.54666f
C542 source.n351 a_n1992_n3288# 0.421764f
C543 source.t29 a_n1992_n3288# 0.297438f
C544 source.t32 a_n1992_n3288# 0.297438f
C545 source.n352 a_n1992_n3288# 2.54666f
C546 source.n353 a_n1992_n3288# 0.421764f
C547 source.n354 a_n1992_n3288# 0.041549f
C548 source.n355 a_n1992_n3288# 0.031366f
C549 source.n356 a_n1992_n3288# 0.016855f
C550 source.n357 a_n1992_n3288# 0.039839f
C551 source.n358 a_n1992_n3288# 0.017846f
C552 source.n359 a_n1992_n3288# 0.031366f
C553 source.n360 a_n1992_n3288# 0.016855f
C554 source.n361 a_n1992_n3288# 0.039839f
C555 source.n362 a_n1992_n3288# 0.017846f
C556 source.n363 a_n1992_n3288# 0.031366f
C557 source.n364 a_n1992_n3288# 0.017351f
C558 source.n365 a_n1992_n3288# 0.039839f
C559 source.n366 a_n1992_n3288# 0.017846f
C560 source.n367 a_n1992_n3288# 0.031366f
C561 source.n368 a_n1992_n3288# 0.016855f
C562 source.n369 a_n1992_n3288# 0.039839f
C563 source.n370 a_n1992_n3288# 0.017846f
C564 source.n371 a_n1992_n3288# 0.031366f
C565 source.n372 a_n1992_n3288# 0.016855f
C566 source.n373 a_n1992_n3288# 0.029879f
C567 source.n374 a_n1992_n3288# 0.028163f
C568 source.t27 a_n1992_n3288# 0.067285f
C569 source.n375 a_n1992_n3288# 0.226147f
C570 source.n376 a_n1992_n3288# 1.58237f
C571 source.n377 a_n1992_n3288# 0.016855f
C572 source.n378 a_n1992_n3288# 0.017846f
C573 source.n379 a_n1992_n3288# 0.039839f
C574 source.n380 a_n1992_n3288# 0.039839f
C575 source.n381 a_n1992_n3288# 0.017846f
C576 source.n382 a_n1992_n3288# 0.016855f
C577 source.n383 a_n1992_n3288# 0.031366f
C578 source.n384 a_n1992_n3288# 0.031366f
C579 source.n385 a_n1992_n3288# 0.016855f
C580 source.n386 a_n1992_n3288# 0.017846f
C581 source.n387 a_n1992_n3288# 0.039839f
C582 source.n388 a_n1992_n3288# 0.039839f
C583 source.n389 a_n1992_n3288# 0.017846f
C584 source.n390 a_n1992_n3288# 0.016855f
C585 source.n391 a_n1992_n3288# 0.031366f
C586 source.n392 a_n1992_n3288# 0.031366f
C587 source.n393 a_n1992_n3288# 0.016855f
C588 source.n394 a_n1992_n3288# 0.016855f
C589 source.n395 a_n1992_n3288# 0.017846f
C590 source.n396 a_n1992_n3288# 0.039839f
C591 source.n397 a_n1992_n3288# 0.039839f
C592 source.n398 a_n1992_n3288# 0.039839f
C593 source.n399 a_n1992_n3288# 0.017351f
C594 source.n400 a_n1992_n3288# 0.016855f
C595 source.n401 a_n1992_n3288# 0.031366f
C596 source.n402 a_n1992_n3288# 0.031366f
C597 source.n403 a_n1992_n3288# 0.016855f
C598 source.n404 a_n1992_n3288# 0.017846f
C599 source.n405 a_n1992_n3288# 0.039839f
C600 source.n406 a_n1992_n3288# 0.039839f
C601 source.n407 a_n1992_n3288# 0.017846f
C602 source.n408 a_n1992_n3288# 0.016855f
C603 source.n409 a_n1992_n3288# 0.031366f
C604 source.n410 a_n1992_n3288# 0.031366f
C605 source.n411 a_n1992_n3288# 0.016855f
C606 source.n412 a_n1992_n3288# 0.017846f
C607 source.n413 a_n1992_n3288# 0.039839f
C608 source.n414 a_n1992_n3288# 0.081753f
C609 source.n415 a_n1992_n3288# 0.017846f
C610 source.n416 a_n1992_n3288# 0.016855f
C611 source.n417 a_n1992_n3288# 0.06736f
C612 source.n418 a_n1992_n3288# 0.045119f
C613 source.n419 a_n1992_n3288# 0.121912f
C614 source.n420 a_n1992_n3288# 0.041549f
C615 source.n421 a_n1992_n3288# 0.031366f
C616 source.n422 a_n1992_n3288# 0.016855f
C617 source.n423 a_n1992_n3288# 0.039839f
C618 source.n424 a_n1992_n3288# 0.017846f
C619 source.n425 a_n1992_n3288# 0.031366f
C620 source.n426 a_n1992_n3288# 0.016855f
C621 source.n427 a_n1992_n3288# 0.039839f
C622 source.n428 a_n1992_n3288# 0.017846f
C623 source.n429 a_n1992_n3288# 0.031366f
C624 source.n430 a_n1992_n3288# 0.017351f
C625 source.n431 a_n1992_n3288# 0.039839f
C626 source.n432 a_n1992_n3288# 0.017846f
C627 source.n433 a_n1992_n3288# 0.031366f
C628 source.n434 a_n1992_n3288# 0.016855f
C629 source.n435 a_n1992_n3288# 0.039839f
C630 source.n436 a_n1992_n3288# 0.017846f
C631 source.n437 a_n1992_n3288# 0.031366f
C632 source.n438 a_n1992_n3288# 0.016855f
C633 source.n439 a_n1992_n3288# 0.029879f
C634 source.n440 a_n1992_n3288# 0.028163f
C635 source.t7 a_n1992_n3288# 0.067285f
C636 source.n441 a_n1992_n3288# 0.226147f
C637 source.n442 a_n1992_n3288# 1.58237f
C638 source.n443 a_n1992_n3288# 0.016855f
C639 source.n444 a_n1992_n3288# 0.017846f
C640 source.n445 a_n1992_n3288# 0.039839f
C641 source.n446 a_n1992_n3288# 0.039839f
C642 source.n447 a_n1992_n3288# 0.017846f
C643 source.n448 a_n1992_n3288# 0.016855f
C644 source.n449 a_n1992_n3288# 0.031366f
C645 source.n450 a_n1992_n3288# 0.031366f
C646 source.n451 a_n1992_n3288# 0.016855f
C647 source.n452 a_n1992_n3288# 0.017846f
C648 source.n453 a_n1992_n3288# 0.039839f
C649 source.n454 a_n1992_n3288# 0.039839f
C650 source.n455 a_n1992_n3288# 0.017846f
C651 source.n456 a_n1992_n3288# 0.016855f
C652 source.n457 a_n1992_n3288# 0.031366f
C653 source.n458 a_n1992_n3288# 0.031366f
C654 source.n459 a_n1992_n3288# 0.016855f
C655 source.n460 a_n1992_n3288# 0.016855f
C656 source.n461 a_n1992_n3288# 0.017846f
C657 source.n462 a_n1992_n3288# 0.039839f
C658 source.n463 a_n1992_n3288# 0.039839f
C659 source.n464 a_n1992_n3288# 0.039839f
C660 source.n465 a_n1992_n3288# 0.017351f
C661 source.n466 a_n1992_n3288# 0.016855f
C662 source.n467 a_n1992_n3288# 0.031366f
C663 source.n468 a_n1992_n3288# 0.031366f
C664 source.n469 a_n1992_n3288# 0.016855f
C665 source.n470 a_n1992_n3288# 0.017846f
C666 source.n471 a_n1992_n3288# 0.039839f
C667 source.n472 a_n1992_n3288# 0.039839f
C668 source.n473 a_n1992_n3288# 0.017846f
C669 source.n474 a_n1992_n3288# 0.016855f
C670 source.n475 a_n1992_n3288# 0.031366f
C671 source.n476 a_n1992_n3288# 0.031366f
C672 source.n477 a_n1992_n3288# 0.016855f
C673 source.n478 a_n1992_n3288# 0.017846f
C674 source.n479 a_n1992_n3288# 0.039839f
C675 source.n480 a_n1992_n3288# 0.081753f
C676 source.n481 a_n1992_n3288# 0.017846f
C677 source.n482 a_n1992_n3288# 0.016855f
C678 source.n483 a_n1992_n3288# 0.06736f
C679 source.n484 a_n1992_n3288# 0.045119f
C680 source.n485 a_n1992_n3288# 0.121912f
C681 source.t8 a_n1992_n3288# 0.297438f
C682 source.t14 a_n1992_n3288# 0.297438f
C683 source.n486 a_n1992_n3288# 2.54666f
C684 source.n487 a_n1992_n3288# 0.421764f
C685 source.t5 a_n1992_n3288# 0.297438f
C686 source.t6 a_n1992_n3288# 0.297438f
C687 source.n488 a_n1992_n3288# 2.54666f
C688 source.n489 a_n1992_n3288# 0.421764f
C689 source.t13 a_n1992_n3288# 0.297438f
C690 source.t4 a_n1992_n3288# 0.297438f
C691 source.n490 a_n1992_n3288# 2.54666f
C692 source.n491 a_n1992_n3288# 0.421764f
C693 source.t0 a_n1992_n3288# 0.297438f
C694 source.t1 a_n1992_n3288# 0.297438f
C695 source.n492 a_n1992_n3288# 2.54666f
C696 source.n493 a_n1992_n3288# 0.421764f
C697 source.n494 a_n1992_n3288# 0.041549f
C698 source.n495 a_n1992_n3288# 0.031366f
C699 source.n496 a_n1992_n3288# 0.016855f
C700 source.n497 a_n1992_n3288# 0.039839f
C701 source.n498 a_n1992_n3288# 0.017846f
C702 source.n499 a_n1992_n3288# 0.031366f
C703 source.n500 a_n1992_n3288# 0.016855f
C704 source.n501 a_n1992_n3288# 0.039839f
C705 source.n502 a_n1992_n3288# 0.017846f
C706 source.n503 a_n1992_n3288# 0.031366f
C707 source.n504 a_n1992_n3288# 0.017351f
C708 source.n505 a_n1992_n3288# 0.039839f
C709 source.n506 a_n1992_n3288# 0.017846f
C710 source.n507 a_n1992_n3288# 0.031366f
C711 source.n508 a_n1992_n3288# 0.016855f
C712 source.n509 a_n1992_n3288# 0.039839f
C713 source.n510 a_n1992_n3288# 0.017846f
C714 source.n511 a_n1992_n3288# 0.031366f
C715 source.n512 a_n1992_n3288# 0.016855f
C716 source.n513 a_n1992_n3288# 0.029879f
C717 source.n514 a_n1992_n3288# 0.028163f
C718 source.t2 a_n1992_n3288# 0.067285f
C719 source.n515 a_n1992_n3288# 0.226147f
C720 source.n516 a_n1992_n3288# 1.58237f
C721 source.n517 a_n1992_n3288# 0.016855f
C722 source.n518 a_n1992_n3288# 0.017846f
C723 source.n519 a_n1992_n3288# 0.039839f
C724 source.n520 a_n1992_n3288# 0.039839f
C725 source.n521 a_n1992_n3288# 0.017846f
C726 source.n522 a_n1992_n3288# 0.016855f
C727 source.n523 a_n1992_n3288# 0.031366f
C728 source.n524 a_n1992_n3288# 0.031366f
C729 source.n525 a_n1992_n3288# 0.016855f
C730 source.n526 a_n1992_n3288# 0.017846f
C731 source.n527 a_n1992_n3288# 0.039839f
C732 source.n528 a_n1992_n3288# 0.039839f
C733 source.n529 a_n1992_n3288# 0.017846f
C734 source.n530 a_n1992_n3288# 0.016855f
C735 source.n531 a_n1992_n3288# 0.031366f
C736 source.n532 a_n1992_n3288# 0.031366f
C737 source.n533 a_n1992_n3288# 0.016855f
C738 source.n534 a_n1992_n3288# 0.016855f
C739 source.n535 a_n1992_n3288# 0.017846f
C740 source.n536 a_n1992_n3288# 0.039839f
C741 source.n537 a_n1992_n3288# 0.039839f
C742 source.n538 a_n1992_n3288# 0.039839f
C743 source.n539 a_n1992_n3288# 0.017351f
C744 source.n540 a_n1992_n3288# 0.016855f
C745 source.n541 a_n1992_n3288# 0.031366f
C746 source.n542 a_n1992_n3288# 0.031366f
C747 source.n543 a_n1992_n3288# 0.016855f
C748 source.n544 a_n1992_n3288# 0.017846f
C749 source.n545 a_n1992_n3288# 0.039839f
C750 source.n546 a_n1992_n3288# 0.039839f
C751 source.n547 a_n1992_n3288# 0.017846f
C752 source.n548 a_n1992_n3288# 0.016855f
C753 source.n549 a_n1992_n3288# 0.031366f
C754 source.n550 a_n1992_n3288# 0.031366f
C755 source.n551 a_n1992_n3288# 0.016855f
C756 source.n552 a_n1992_n3288# 0.017846f
C757 source.n553 a_n1992_n3288# 0.039839f
C758 source.n554 a_n1992_n3288# 0.081753f
C759 source.n555 a_n1992_n3288# 0.017846f
C760 source.n556 a_n1992_n3288# 0.016855f
C761 source.n557 a_n1992_n3288# 0.06736f
C762 source.n558 a_n1992_n3288# 0.045119f
C763 source.n559 a_n1992_n3288# 0.295487f
C764 source.n560 a_n1992_n3288# 1.96529f
C765 plus.n0 a_n1992_n3288# 0.051837f
C766 plus.t12 a_n1992_n3288# 0.439448f
C767 plus.t3 a_n1992_n3288# 0.439448f
C768 plus.t8 a_n1992_n3288# 0.439448f
C769 plus.n1 a_n1992_n3288# 0.17699f
C770 plus.n2 a_n1992_n3288# 0.051837f
C771 plus.t18 a_n1992_n3288# 0.439448f
C772 plus.t9 a_n1992_n3288# 0.439448f
C773 plus.n3 a_n1992_n3288# 0.17699f
C774 plus.n4 a_n1992_n3288# 0.051837f
C775 plus.t0 a_n1992_n3288# 0.439448f
C776 plus.t10 a_n1992_n3288# 0.439448f
C777 plus.t1 a_n1992_n3288# 0.439448f
C778 plus.n5 a_n1992_n3288# 0.17699f
C779 plus.t5 a_n1992_n3288# 0.446559f
C780 plus.n6 a_n1992_n3288# 0.193226f
C781 plus.n7 a_n1992_n3288# 0.118617f
C782 plus.n8 a_n1992_n3288# 0.019753f
C783 plus.n9 a_n1992_n3288# 0.17699f
C784 plus.n10 a_n1992_n3288# 0.019753f
C785 plus.n11 a_n1992_n3288# 0.17699f
C786 plus.n12 a_n1992_n3288# 0.019753f
C787 plus.n13 a_n1992_n3288# 0.051837f
C788 plus.n14 a_n1992_n3288# 0.051837f
C789 plus.n15 a_n1992_n3288# 0.018475f
C790 plus.n16 a_n1992_n3288# 0.018475f
C791 plus.n17 a_n1992_n3288# 0.17699f
C792 plus.n18 a_n1992_n3288# 0.019753f
C793 plus.n19 a_n1992_n3288# 0.051837f
C794 plus.n20 a_n1992_n3288# 0.051837f
C795 plus.n21 a_n1992_n3288# 0.019753f
C796 plus.n22 a_n1992_n3288# 0.17699f
C797 plus.n23 a_n1992_n3288# 0.019753f
C798 plus.n24 a_n1992_n3288# 0.17699f
C799 plus.t2 a_n1992_n3288# 0.446559f
C800 plus.n25 a_n1992_n3288# 0.193147f
C801 plus.n26 a_n1992_n3288# 0.579572f
C802 plus.n27 a_n1992_n3288# 0.051837f
C803 plus.t11 a_n1992_n3288# 0.446559f
C804 plus.t15 a_n1992_n3288# 0.439448f
C805 plus.t6 a_n1992_n3288# 0.439448f
C806 plus.t13 a_n1992_n3288# 0.439448f
C807 plus.n28 a_n1992_n3288# 0.17699f
C808 plus.n29 a_n1992_n3288# 0.051837f
C809 plus.t16 a_n1992_n3288# 0.439448f
C810 plus.t4 a_n1992_n3288# 0.439448f
C811 plus.n30 a_n1992_n3288# 0.17699f
C812 plus.n31 a_n1992_n3288# 0.051837f
C813 plus.t19 a_n1992_n3288# 0.439448f
C814 plus.t7 a_n1992_n3288# 0.439448f
C815 plus.t14 a_n1992_n3288# 0.439448f
C816 plus.n32 a_n1992_n3288# 0.17699f
C817 plus.t17 a_n1992_n3288# 0.446559f
C818 plus.n33 a_n1992_n3288# 0.193226f
C819 plus.n34 a_n1992_n3288# 0.118617f
C820 plus.n35 a_n1992_n3288# 0.019753f
C821 plus.n36 a_n1992_n3288# 0.17699f
C822 plus.n37 a_n1992_n3288# 0.019753f
C823 plus.n38 a_n1992_n3288# 0.17699f
C824 plus.n39 a_n1992_n3288# 0.019753f
C825 plus.n40 a_n1992_n3288# 0.051837f
C826 plus.n41 a_n1992_n3288# 0.051837f
C827 plus.n42 a_n1992_n3288# 0.018475f
C828 plus.n43 a_n1992_n3288# 0.018475f
C829 plus.n44 a_n1992_n3288# 0.17699f
C830 plus.n45 a_n1992_n3288# 0.019753f
C831 plus.n46 a_n1992_n3288# 0.051837f
C832 plus.n47 a_n1992_n3288# 0.051837f
C833 plus.n48 a_n1992_n3288# 0.019753f
C834 plus.n49 a_n1992_n3288# 0.17699f
C835 plus.n50 a_n1992_n3288# 0.019753f
C836 plus.n51 a_n1992_n3288# 0.17699f
C837 plus.n52 a_n1992_n3288# 0.193147f
C838 plus.n53 a_n1992_n3288# 1.58231f
.ends

