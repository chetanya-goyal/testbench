* NGSPICE file created from diffpair83.ext - technology: sky130A

.subckt diffpair83 minus drain_right drain_left source plus
X0 source.t10 minus.t0 drain_right.t0 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X1 a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X2 source.t11 plus.t0 drain_left.t7 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 drain_left.t6 plus.t1 source.t12 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 drain_right.t7 minus.t1 source.t9 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X5 a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X6 a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X7 a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X8 source.t8 minus.t2 drain_right.t5 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X9 source.t7 minus.t3 drain_right.t2 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 drain_right.t1 minus.t4 source.t6 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X11 source.t5 minus.t5 drain_right.t3 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X12 drain_right.t6 minus.t6 source.t4 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 source.t13 plus.t2 drain_left.t5 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t14 plus.t3 drain_left.t4 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X15 drain_right.t4 minus.t7 source.t3 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 drain_left.t3 plus.t4 source.t0 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X17 drain_left.t2 plus.t5 source.t15 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X18 source.t1 plus.t6 drain_left.t1 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 drain_left.t0 plus.t7 source.t2 a_n1366_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 minus.n5 minus.t5 599.58
R1 minus.n1 minus.t4 599.58
R2 minus.n12 minus.t1 599.58
R3 minus.n8 minus.t0 599.58
R4 minus.n4 minus.t7 530.201
R5 minus.n2 minus.t2 530.201
R6 minus.n11 minus.t3 530.201
R7 minus.n9 minus.t6 530.201
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 26.7997
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 drain_right.n5 drain_right.n3 101.356
R28 drain_right.n2 drain_right.n1 101.02
R29 drain_right.n2 drain_right.n0 101.02
R30 drain_right.n5 drain_right.n4 100.796
R31 drain_right drain_right.n2 21.1993
R32 drain_right.n1 drain_right.t2 15.0005
R33 drain_right.n1 drain_right.t7 15.0005
R34 drain_right.n0 drain_right.t0 15.0005
R35 drain_right.n0 drain_right.t6 15.0005
R36 drain_right.n3 drain_right.t5 15.0005
R37 drain_right.n3 drain_right.t1 15.0005
R38 drain_right.n4 drain_right.t3 15.0005
R39 drain_right.n4 drain_right.t4 15.0005
R40 drain_right drain_right.n5 6.21356
R41 source.n0 source.t0 99.1169
R42 source.n3 source.t14 99.1169
R43 source.n4 source.t6 99.1169
R44 source.n7 source.t5 99.1169
R45 source.n15 source.t9 99.1168
R46 source.n12 source.t10 99.1168
R47 source.n11 source.t15 99.1168
R48 source.n8 source.t11 99.1168
R49 source.n2 source.n1 84.1169
R50 source.n6 source.n5 84.1169
R51 source.n14 source.n13 84.1168
R52 source.n10 source.n9 84.1168
R53 source.n13 source.t4 15.0005
R54 source.n13 source.t7 15.0005
R55 source.n9 source.t12 15.0005
R56 source.n9 source.t13 15.0005
R57 source.n1 source.t2 15.0005
R58 source.n1 source.t1 15.0005
R59 source.n5 source.t3 15.0005
R60 source.n5 source.t8 15.0005
R61 source.n8 source.n7 14.2723
R62 source.n16 source.n0 8.72921
R63 source.n16 source.n15 5.5436
R64 source.n7 source.n6 0.560845
R65 source.n6 source.n4 0.560845
R66 source.n3 source.n2 0.560845
R67 source.n2 source.n0 0.560845
R68 source.n10 source.n8 0.560845
R69 source.n11 source.n10 0.560845
R70 source.n14 source.n12 0.560845
R71 source.n15 source.n14 0.560845
R72 source.n4 source.n3 0.470328
R73 source.n12 source.n11 0.470328
R74 source source.n16 0.188
R75 plus.n1 plus.t3 599.58
R76 plus.n5 plus.t4 599.58
R77 plus.n8 plus.t5 599.58
R78 plus.n12 plus.t0 599.58
R79 plus.n2 plus.t7 530.201
R80 plus.n4 plus.t6 530.201
R81 plus.n9 plus.t2 530.201
R82 plus.n11 plus.t1 530.201
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus.n2 plus.n1 25.5611
R94 plus.n5 plus.n4 25.5611
R95 plus.n12 plus.n11 25.5611
R96 plus.n9 plus.n8 25.5611
R97 plus plus.n13 24.4687
R98 plus plus.n6 8.43611
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 101.356
R102 drain_left.n2 drain_left.n1 101.02
R103 drain_left.n2 drain_left.n0 101.02
R104 drain_left.n5 drain_left.n4 100.796
R105 drain_left drain_left.n2 21.7525
R106 drain_left.n1 drain_left.t5 15.0005
R107 drain_left.n1 drain_left.t2 15.0005
R108 drain_left.n0 drain_left.t7 15.0005
R109 drain_left.n0 drain_left.t6 15.0005
R110 drain_left.n4 drain_left.t1 15.0005
R111 drain_left.n4 drain_left.t3 15.0005
R112 drain_left.n3 drain_left.t4 15.0005
R113 drain_left.n3 drain_left.t0 15.0005
R114 drain_left drain_left.n5 6.21356
C0 drain_right source 4.35965f
C1 drain_right plus 0.289056f
C2 drain_right minus 0.65096f
C3 source drain_left 4.36032f
C4 drain_left plus 0.780361f
C5 drain_left minus 0.176331f
C6 source plus 0.682733f
C7 source minus 0.66877f
C8 minus plus 2.99093f
C9 drain_right drain_left 0.640281f
C10 drain_right a_n1366_n1288# 3.09177f
C11 drain_left a_n1366_n1288# 3.2574f
C12 source a_n1366_n1288# 2.929171f
C13 minus a_n1366_n1288# 4.200463f
C14 plus a_n1366_n1288# 5.03788f
C15 drain_left.t7 a_n1366_n1288# 0.054748f
C16 drain_left.t6 a_n1366_n1288# 0.054748f
C17 drain_left.n0 a_n1366_n1288# 0.264776f
C18 drain_left.t5 a_n1366_n1288# 0.054748f
C19 drain_left.t2 a_n1366_n1288# 0.054748f
C20 drain_left.n1 a_n1366_n1288# 0.264776f
C21 drain_left.n2 a_n1366_n1288# 1.03377f
C22 drain_left.t4 a_n1366_n1288# 0.054748f
C23 drain_left.t0 a_n1366_n1288# 0.054748f
C24 drain_left.n3 a_n1366_n1288# 0.265708f
C25 drain_left.t1 a_n1366_n1288# 0.054748f
C26 drain_left.t3 a_n1366_n1288# 0.054748f
C27 drain_left.n4 a_n1366_n1288# 0.264233f
C28 drain_left.n5 a_n1366_n1288# 0.713761f
C29 plus.n0 a_n1366_n1288# 0.096087f
C30 plus.t6 a_n1366_n1288# 0.035816f
C31 plus.t7 a_n1366_n1288# 0.035816f
C32 plus.t3 a_n1366_n1288# 0.039796f
C33 plus.n1 a_n1366_n1288# 0.047691f
C34 plus.n2 a_n1366_n1288# 0.031268f
C35 plus.n3 a_n1366_n1288# 0.017211f
C36 plus.n4 a_n1366_n1288# 0.031268f
C37 plus.t4 a_n1366_n1288# 0.039796f
C38 plus.n5 a_n1366_n1288# 0.047626f
C39 plus.n6 a_n1366_n1288# 0.298079f
C40 plus.n7 a_n1366_n1288# 0.096087f
C41 plus.t0 a_n1366_n1288# 0.039796f
C42 plus.t1 a_n1366_n1288# 0.035816f
C43 plus.t2 a_n1366_n1288# 0.035816f
C44 plus.t5 a_n1366_n1288# 0.039796f
C45 plus.n8 a_n1366_n1288# 0.047691f
C46 plus.n9 a_n1366_n1288# 0.031268f
C47 plus.n10 a_n1366_n1288# 0.017211f
C48 plus.n11 a_n1366_n1288# 0.031268f
C49 plus.n12 a_n1366_n1288# 0.047626f
C50 plus.n13 a_n1366_n1288# 0.83433f
C51 source.t0 a_n1366_n1288# 0.281659f
C52 source.n0 a_n1366_n1288# 0.536834f
C53 source.t2 a_n1366_n1288# 0.053645f
C54 source.t1 a_n1366_n1288# 0.053645f
C55 source.n1 a_n1366_n1288# 0.225758f
C56 source.n2 a_n1366_n1288# 0.255064f
C57 source.t14 a_n1366_n1288# 0.281659f
C58 source.n3 a_n1366_n1288# 0.289191f
C59 source.t6 a_n1366_n1288# 0.281659f
C60 source.n4 a_n1366_n1288# 0.289191f
C61 source.t3 a_n1366_n1288# 0.053645f
C62 source.t8 a_n1366_n1288# 0.053645f
C63 source.n5 a_n1366_n1288# 0.225758f
C64 source.n6 a_n1366_n1288# 0.255064f
C65 source.t5 a_n1366_n1288# 0.281659f
C66 source.n7 a_n1366_n1288# 0.745969f
C67 source.t11 a_n1366_n1288# 0.281658f
C68 source.n8 a_n1366_n1288# 0.74597f
C69 source.t12 a_n1366_n1288# 0.053645f
C70 source.t13 a_n1366_n1288# 0.053645f
C71 source.n9 a_n1366_n1288# 0.225756f
C72 source.n10 a_n1366_n1288# 0.255065f
C73 source.t15 a_n1366_n1288# 0.281658f
C74 source.n11 a_n1366_n1288# 0.289192f
C75 source.t10 a_n1366_n1288# 0.281658f
C76 source.n12 a_n1366_n1288# 0.289192f
C77 source.t4 a_n1366_n1288# 0.053645f
C78 source.t7 a_n1366_n1288# 0.053645f
C79 source.n13 a_n1366_n1288# 0.225756f
C80 source.n14 a_n1366_n1288# 0.255065f
C81 source.t9 a_n1366_n1288# 0.281658f
C82 source.n15 a_n1366_n1288# 0.416646f
C83 source.n16 a_n1366_n1288# 0.554392f
C84 drain_right.t0 a_n1366_n1288# 0.055884f
C85 drain_right.t6 a_n1366_n1288# 0.055884f
C86 drain_right.n0 a_n1366_n1288# 0.27027f
C87 drain_right.t2 a_n1366_n1288# 0.055884f
C88 drain_right.t7 a_n1366_n1288# 0.055884f
C89 drain_right.n1 a_n1366_n1288# 0.27027f
C90 drain_right.n2 a_n1366_n1288# 1.00928f
C91 drain_right.t5 a_n1366_n1288# 0.055884f
C92 drain_right.t1 a_n1366_n1288# 0.055884f
C93 drain_right.n3 a_n1366_n1288# 0.271221f
C94 drain_right.t3 a_n1366_n1288# 0.055884f
C95 drain_right.t4 a_n1366_n1288# 0.055884f
C96 drain_right.n4 a_n1366_n1288# 0.269716f
C97 drain_right.n5 a_n1366_n1288# 0.728571f
C98 minus.n0 a_n1366_n1288# 0.093529f
C99 minus.t5 a_n1366_n1288# 0.038736f
C100 minus.t7 a_n1366_n1288# 0.034862f
C101 minus.t2 a_n1366_n1288# 0.034862f
C102 minus.t4 a_n1366_n1288# 0.038736f
C103 minus.n1 a_n1366_n1288# 0.046421f
C104 minus.n2 a_n1366_n1288# 0.030435f
C105 minus.n3 a_n1366_n1288# 0.016753f
C106 minus.n4 a_n1366_n1288# 0.030435f
C107 minus.n5 a_n1366_n1288# 0.046358f
C108 minus.n6 a_n1366_n1288# 0.845719f
C109 minus.n7 a_n1366_n1288# 0.093529f
C110 minus.t3 a_n1366_n1288# 0.034862f
C111 minus.t6 a_n1366_n1288# 0.034862f
C112 minus.t0 a_n1366_n1288# 0.038736f
C113 minus.n8 a_n1366_n1288# 0.046421f
C114 minus.n9 a_n1366_n1288# 0.030435f
C115 minus.n10 a_n1366_n1288# 0.016753f
C116 minus.n11 a_n1366_n1288# 0.030435f
C117 minus.t1 a_n1366_n1288# 0.038736f
C118 minus.n12 a_n1366_n1288# 0.046358f
C119 minus.n13 a_n1366_n1288# 0.265605f
C120 minus.n14 a_n1366_n1288# 1.04049f
.ends

