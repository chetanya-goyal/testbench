* NGSPICE file created from diffpair544.ext - technology: sky130A

.subckt diffpair544 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t16 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X1 drain_left.t9 plus.t0 source.t3 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X2 source.t6 plus.t1 drain_left.t8 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X3 drain_left.t7 plus.t2 source.t0 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X4 source.t11 minus.t1 drain_right.t8 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 source.t12 minus.t2 drain_right.t7 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X6 a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X7 a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X8 a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X9 drain_left.t6 plus.t3 source.t1 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X10 drain_left.t5 plus.t4 source.t5 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X11 drain_right.t6 minus.t3 source.t15 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X12 drain_right.t5 minus.t4 source.t14 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X13 source.t19 minus.t5 drain_right.t4 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X14 drain_right.t3 minus.t6 source.t17 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X15 a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X16 drain_right.t2 minus.t7 source.t13 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X17 source.t7 plus.t5 drain_left.t4 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X18 drain_right.t1 minus.t8 source.t18 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X19 source.t2 plus.t6 drain_left.t3 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X20 drain_left.t2 plus.t7 source.t4 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X21 source.t8 plus.t8 drain_left.t1 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X22 drain_left.t0 plus.t9 source.t9 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X23 source.t10 minus.t9 drain_right.t0 a_n1952_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
R0 minus.n3 minus.t8 595.295
R1 minus.n17 minus.t4 595.295
R2 minus.n4 minus.t1 572.548
R3 minus.n6 minus.t7 572.548
R4 minus.n10 minus.t9 572.548
R5 minus.n12 minus.t6 572.548
R6 minus.n18 minus.t5 572.548
R7 minus.n20 minus.t0 572.548
R8 minus.n24 minus.t2 572.548
R9 minus.n26 minus.t3 572.548
R10 minus.n13 minus.n12 161.3
R11 minus.n11 minus.n0 161.3
R12 minus.n10 minus.n9 161.3
R13 minus.n8 minus.n1 161.3
R14 minus.n7 minus.n6 161.3
R15 minus.n5 minus.n2 161.3
R16 minus.n27 minus.n26 161.3
R17 minus.n25 minus.n14 161.3
R18 minus.n24 minus.n23 161.3
R19 minus.n22 minus.n15 161.3
R20 minus.n21 minus.n20 161.3
R21 minus.n19 minus.n16 161.3
R22 minus.n3 minus.n2 44.8741
R23 minus.n17 minus.n16 44.8741
R24 minus.n28 minus.n13 38.9266
R25 minus.n12 minus.n11 30.6732
R26 minus.n26 minus.n25 30.6732
R27 minus.n5 minus.n4 26.2914
R28 minus.n10 minus.n1 26.2914
R29 minus.n19 minus.n18 26.2914
R30 minus.n24 minus.n15 26.2914
R31 minus.n6 minus.n5 21.9096
R32 minus.n6 minus.n1 21.9096
R33 minus.n20 minus.n19 21.9096
R34 minus.n20 minus.n15 21.9096
R35 minus.n4 minus.n3 19.0667
R36 minus.n18 minus.n17 19.0667
R37 minus.n11 minus.n10 17.5278
R38 minus.n25 minus.n24 17.5278
R39 minus.n28 minus.n27 6.63876
R40 minus.n13 minus.n0 0.189894
R41 minus.n9 minus.n0 0.189894
R42 minus.n9 minus.n8 0.189894
R43 minus.n8 minus.n7 0.189894
R44 minus.n7 minus.n2 0.189894
R45 minus.n21 minus.n16 0.189894
R46 minus.n22 minus.n21 0.189894
R47 minus.n23 minus.n22 0.189894
R48 minus.n23 minus.n14 0.189894
R49 minus.n27 minus.n14 0.189894
R50 minus minus.n28 0.188
R51 source.n5 source.t18 45.521
R52 source.n19 source.t15 45.5208
R53 source.n14 source.t3 45.5208
R54 source.n0 source.t1 45.5208
R55 source.n2 source.n1 44.201
R56 source.n4 source.n3 44.201
R57 source.n7 source.n6 44.201
R58 source.n9 source.n8 44.201
R59 source.n18 source.n17 44.2008
R60 source.n16 source.n15 44.2008
R61 source.n13 source.n12 44.2008
R62 source.n11 source.n10 44.2008
R63 source.n11 source.n9 25.3363
R64 source.n20 source.n0 18.7415
R65 source.n20 source.n19 5.7074
R66 source.n17 source.t16 1.3205
R67 source.n17 source.t12 1.3205
R68 source.n15 source.t14 1.3205
R69 source.n15 source.t19 1.3205
R70 source.n12 source.t9 1.3205
R71 source.n12 source.t6 1.3205
R72 source.n10 source.t4 1.3205
R73 source.n10 source.t2 1.3205
R74 source.n1 source.t0 1.3205
R75 source.n1 source.t7 1.3205
R76 source.n3 source.t5 1.3205
R77 source.n3 source.t8 1.3205
R78 source.n6 source.t13 1.3205
R79 source.n6 source.t11 1.3205
R80 source.n8 source.t17 1.3205
R81 source.n8 source.t10 1.3205
R82 source.n5 source.n4 0.914293
R83 source.n16 source.n14 0.914293
R84 source.n9 source.n7 0.888431
R85 source.n7 source.n5 0.888431
R86 source.n4 source.n2 0.888431
R87 source.n2 source.n0 0.888431
R88 source.n13 source.n11 0.888431
R89 source.n14 source.n13 0.888431
R90 source.n18 source.n16 0.888431
R91 source.n19 source.n18 0.888431
R92 source source.n20 0.188
R93 drain_right.n1 drain_right.t5 63.0875
R94 drain_right.n7 drain_right.t3 62.1998
R95 drain_right.n6 drain_right.n4 61.7676
R96 drain_right.n3 drain_right.n2 61.4902
R97 drain_right.n6 drain_right.n5 60.8798
R98 drain_right.n1 drain_right.n0 60.8796
R99 drain_right drain_right.n3 32.8603
R100 drain_right drain_right.n7 6.09718
R101 drain_right.n2 drain_right.t7 1.3205
R102 drain_right.n2 drain_right.t6 1.3205
R103 drain_right.n0 drain_right.t4 1.3205
R104 drain_right.n0 drain_right.t9 1.3205
R105 drain_right.n4 drain_right.t8 1.3205
R106 drain_right.n4 drain_right.t1 1.3205
R107 drain_right.n5 drain_right.t0 1.3205
R108 drain_right.n5 drain_right.t2 1.3205
R109 drain_right.n7 drain_right.n6 0.888431
R110 drain_right.n3 drain_right.n1 0.167137
R111 plus.n3 plus.t4 595.295
R112 plus.n17 plus.t0 595.295
R113 plus.n12 plus.t3 572.548
R114 plus.n10 plus.t5 572.548
R115 plus.n2 plus.t2 572.548
R116 plus.n4 plus.t8 572.548
R117 plus.n26 plus.t7 572.548
R118 plus.n24 plus.t6 572.548
R119 plus.n16 plus.t9 572.548
R120 plus.n18 plus.t1 572.548
R121 plus.n6 plus.n5 161.3
R122 plus.n7 plus.n2 161.3
R123 plus.n9 plus.n8 161.3
R124 plus.n10 plus.n1 161.3
R125 plus.n11 plus.n0 161.3
R126 plus.n13 plus.n12 161.3
R127 plus.n20 plus.n19 161.3
R128 plus.n21 plus.n16 161.3
R129 plus.n23 plus.n22 161.3
R130 plus.n24 plus.n15 161.3
R131 plus.n25 plus.n14 161.3
R132 plus.n27 plus.n26 161.3
R133 plus.n6 plus.n3 44.8741
R134 plus.n20 plus.n17 44.8741
R135 plus plus.n27 31.6714
R136 plus.n12 plus.n11 30.6732
R137 plus.n26 plus.n25 30.6732
R138 plus.n10 plus.n9 26.2914
R139 plus.n5 plus.n4 26.2914
R140 plus.n24 plus.n23 26.2914
R141 plus.n19 plus.n18 26.2914
R142 plus.n9 plus.n2 21.9096
R143 plus.n5 plus.n2 21.9096
R144 plus.n23 plus.n16 21.9096
R145 plus.n19 plus.n16 21.9096
R146 plus.n4 plus.n3 19.0667
R147 plus.n18 plus.n17 19.0667
R148 plus.n11 plus.n10 17.5278
R149 plus.n25 plus.n24 17.5278
R150 plus plus.n13 13.4191
R151 plus.n7 plus.n6 0.189894
R152 plus.n8 plus.n7 0.189894
R153 plus.n8 plus.n1 0.189894
R154 plus.n1 plus.n0 0.189894
R155 plus.n13 plus.n0 0.189894
R156 plus.n27 plus.n14 0.189894
R157 plus.n15 plus.n14 0.189894
R158 plus.n22 plus.n15 0.189894
R159 plus.n22 plus.n21 0.189894
R160 plus.n21 plus.n20 0.189894
R161 drain_left.n5 drain_left.t5 63.0877
R162 drain_left.n1 drain_left.t2 63.0875
R163 drain_left.n3 drain_left.n2 61.4902
R164 drain_left.n5 drain_left.n4 60.8798
R165 drain_left.n7 drain_left.n6 60.8796
R166 drain_left.n1 drain_left.n0 60.8796
R167 drain_left drain_left.n3 33.4135
R168 drain_left drain_left.n7 6.54115
R169 drain_left.n2 drain_left.t8 1.3205
R170 drain_left.n2 drain_left.t9 1.3205
R171 drain_left.n0 drain_left.t3 1.3205
R172 drain_left.n0 drain_left.t0 1.3205
R173 drain_left.n6 drain_left.t4 1.3205
R174 drain_left.n6 drain_left.t6 1.3205
R175 drain_left.n4 drain_left.t1 1.3205
R176 drain_left.n4 drain_left.t7 1.3205
R177 drain_left.n7 drain_left.n5 0.888431
R178 drain_left.n3 drain_left.n1 0.167137
C0 source minus 7.99491f
C1 minus plus 6.13266f
C2 drain_left minus 0.171897f
C3 source plus 8.00958f
C4 source drain_left 17.312302f
C5 drain_left plus 8.46795f
C6 drain_right minus 8.28059f
C7 source drain_right 17.3039f
C8 drain_right plus 0.347623f
C9 drain_right drain_left 0.970098f
C10 drain_right a_n1952_n3888# 7.78267f
C11 drain_left a_n1952_n3888# 8.080919f
C12 source a_n1952_n3888# 7.609848f
C13 minus a_n1952_n3888# 7.838418f
C14 plus a_n1952_n3888# 9.68802f
C15 drain_left.t2 a_n1952_n3888# 3.34298f
C16 drain_left.t3 a_n1952_n3888# 0.289324f
C17 drain_left.t0 a_n1952_n3888# 0.289324f
C18 drain_left.n0 a_n1952_n3888# 2.61515f
C19 drain_left.n1 a_n1952_n3888# 0.627083f
C20 drain_left.t8 a_n1952_n3888# 0.289324f
C21 drain_left.t9 a_n1952_n3888# 0.289324f
C22 drain_left.n2 a_n1952_n3888# 2.61842f
C23 drain_left.n3 a_n1952_n3888# 1.74283f
C24 drain_left.t5 a_n1952_n3888# 3.34298f
C25 drain_left.t1 a_n1952_n3888# 0.289324f
C26 drain_left.t7 a_n1952_n3888# 0.289324f
C27 drain_left.n4 a_n1952_n3888# 2.61515f
C28 drain_left.n5 a_n1952_n3888# 0.680412f
C29 drain_left.t4 a_n1952_n3888# 0.289324f
C30 drain_left.t6 a_n1952_n3888# 0.289324f
C31 drain_left.n6 a_n1952_n3888# 2.61515f
C32 drain_left.n7 a_n1952_n3888# 0.555492f
C33 plus.n0 a_n1952_n3888# 0.043105f
C34 plus.t3 a_n1952_n3888# 1.28616f
C35 plus.t5 a_n1952_n3888# 1.28616f
C36 plus.n1 a_n1952_n3888# 0.043105f
C37 plus.t2 a_n1952_n3888# 1.28616f
C38 plus.n2 a_n1952_n3888# 0.496332f
C39 plus.t4 a_n1952_n3888# 1.30512f
C40 plus.n3 a_n1952_n3888# 0.481301f
C41 plus.t8 a_n1952_n3888# 1.28616f
C42 plus.n4 a_n1952_n3888# 0.500675f
C43 plus.n5 a_n1952_n3888# 0.009781f
C44 plus.n6 a_n1952_n3888# 0.18004f
C45 plus.n7 a_n1952_n3888# 0.043105f
C46 plus.n8 a_n1952_n3888# 0.043105f
C47 plus.n9 a_n1952_n3888# 0.009781f
C48 plus.n10 a_n1952_n3888# 0.496332f
C49 plus.n11 a_n1952_n3888# 0.009781f
C50 plus.n12 a_n1952_n3888# 0.49394f
C51 plus.n13 a_n1952_n3888# 0.558755f
C52 plus.n14 a_n1952_n3888# 0.043105f
C53 plus.t7 a_n1952_n3888# 1.28616f
C54 plus.n15 a_n1952_n3888# 0.043105f
C55 plus.t6 a_n1952_n3888# 1.28616f
C56 plus.t9 a_n1952_n3888# 1.28616f
C57 plus.n16 a_n1952_n3888# 0.496332f
C58 plus.t0 a_n1952_n3888# 1.30512f
C59 plus.n17 a_n1952_n3888# 0.481301f
C60 plus.t1 a_n1952_n3888# 1.28616f
C61 plus.n18 a_n1952_n3888# 0.500675f
C62 plus.n19 a_n1952_n3888# 0.009781f
C63 plus.n20 a_n1952_n3888# 0.18004f
C64 plus.n21 a_n1952_n3888# 0.043105f
C65 plus.n22 a_n1952_n3888# 0.043105f
C66 plus.n23 a_n1952_n3888# 0.009781f
C67 plus.n24 a_n1952_n3888# 0.496332f
C68 plus.n25 a_n1952_n3888# 0.009781f
C69 plus.n26 a_n1952_n3888# 0.49394f
C70 plus.n27 a_n1952_n3888# 1.40949f
C71 drain_right.t5 a_n1952_n3888# 3.32939f
C72 drain_right.t4 a_n1952_n3888# 0.288148f
C73 drain_right.t9 a_n1952_n3888# 0.288148f
C74 drain_right.n0 a_n1952_n3888# 2.60452f
C75 drain_right.n1 a_n1952_n3888# 0.624533f
C76 drain_right.t7 a_n1952_n3888# 0.288148f
C77 drain_right.t6 a_n1952_n3888# 0.288148f
C78 drain_right.n2 a_n1952_n3888# 2.60777f
C79 drain_right.n3 a_n1952_n3888# 1.68522f
C80 drain_right.t8 a_n1952_n3888# 0.288148f
C81 drain_right.t1 a_n1952_n3888# 0.288148f
C82 drain_right.n4 a_n1952_n3888# 2.60952f
C83 drain_right.t0 a_n1952_n3888# 0.288148f
C84 drain_right.t2 a_n1952_n3888# 0.288148f
C85 drain_right.n5 a_n1952_n3888# 2.60452f
C86 drain_right.n6 a_n1952_n3888# 0.681213f
C87 drain_right.t3 a_n1952_n3888# 3.32454f
C88 drain_right.n7 a_n1952_n3888# 0.567698f
C89 source.t1 a_n1952_n3888# 3.34653f
C90 source.n0 a_n1952_n3888# 1.59517f
C91 source.t0 a_n1952_n3888# 0.298621f
C92 source.t7 a_n1952_n3888# 0.298621f
C93 source.n1 a_n1952_n3888# 2.62313f
C94 source.n2 a_n1952_n3888# 0.39231f
C95 source.t5 a_n1952_n3888# 0.298621f
C96 source.t8 a_n1952_n3888# 0.298621f
C97 source.n3 a_n1952_n3888# 2.62313f
C98 source.n4 a_n1952_n3888# 0.394409f
C99 source.t18 a_n1952_n3888# 3.34653f
C100 source.n5 a_n1952_n3888# 0.485432f
C101 source.t13 a_n1952_n3888# 0.298621f
C102 source.t11 a_n1952_n3888# 0.298621f
C103 source.n6 a_n1952_n3888# 2.62313f
C104 source.n7 a_n1952_n3888# 0.39231f
C105 source.t17 a_n1952_n3888# 0.298621f
C106 source.t10 a_n1952_n3888# 0.298621f
C107 source.n8 a_n1952_n3888# 2.62313f
C108 source.n9 a_n1952_n3888# 2.00594f
C109 source.t4 a_n1952_n3888# 0.298621f
C110 source.t2 a_n1952_n3888# 0.298621f
C111 source.n10 a_n1952_n3888# 2.62313f
C112 source.n11 a_n1952_n3888# 2.00594f
C113 source.t9 a_n1952_n3888# 0.298621f
C114 source.t6 a_n1952_n3888# 0.298621f
C115 source.n12 a_n1952_n3888# 2.62313f
C116 source.n13 a_n1952_n3888# 0.392313f
C117 source.t3 a_n1952_n3888# 3.34653f
C118 source.n14 a_n1952_n3888# 0.485436f
C119 source.t14 a_n1952_n3888# 0.298621f
C120 source.t19 a_n1952_n3888# 0.298621f
C121 source.n15 a_n1952_n3888# 2.62313f
C122 source.n16 a_n1952_n3888# 0.394413f
C123 source.t16 a_n1952_n3888# 0.298621f
C124 source.t12 a_n1952_n3888# 0.298621f
C125 source.n17 a_n1952_n3888# 2.62313f
C126 source.n18 a_n1952_n3888# 0.392313f
C127 source.t15 a_n1952_n3888# 3.34653f
C128 source.n19 a_n1952_n3888# 0.613729f
C129 source.n20 a_n1952_n3888# 1.85879f
C130 minus.n0 a_n1952_n3888# 0.042559f
C131 minus.n1 a_n1952_n3888# 0.009658f
C132 minus.t9 a_n1952_n3888# 1.26988f
C133 minus.n2 a_n1952_n3888# 0.177761f
C134 minus.t8 a_n1952_n3888# 1.2886f
C135 minus.n3 a_n1952_n3888# 0.475209f
C136 minus.t1 a_n1952_n3888# 1.26988f
C137 minus.n4 a_n1952_n3888# 0.494338f
C138 minus.n5 a_n1952_n3888# 0.009658f
C139 minus.t7 a_n1952_n3888# 1.26988f
C140 minus.n6 a_n1952_n3888# 0.490049f
C141 minus.n7 a_n1952_n3888# 0.042559f
C142 minus.n8 a_n1952_n3888# 0.042559f
C143 minus.n9 a_n1952_n3888# 0.042559f
C144 minus.n10 a_n1952_n3888# 0.490049f
C145 minus.n11 a_n1952_n3888# 0.009658f
C146 minus.t6 a_n1952_n3888# 1.26988f
C147 minus.n12 a_n1952_n3888# 0.487688f
C148 minus.n13 a_n1952_n3888# 1.68672f
C149 minus.n14 a_n1952_n3888# 0.042559f
C150 minus.n15 a_n1952_n3888# 0.009658f
C151 minus.n16 a_n1952_n3888# 0.177761f
C152 minus.t4 a_n1952_n3888# 1.2886f
C153 minus.n17 a_n1952_n3888# 0.475209f
C154 minus.t5 a_n1952_n3888# 1.26988f
C155 minus.n18 a_n1952_n3888# 0.494338f
C156 minus.n19 a_n1952_n3888# 0.009658f
C157 minus.t0 a_n1952_n3888# 1.26988f
C158 minus.n20 a_n1952_n3888# 0.490049f
C159 minus.n21 a_n1952_n3888# 0.042559f
C160 minus.n22 a_n1952_n3888# 0.042559f
C161 minus.n23 a_n1952_n3888# 0.042559f
C162 minus.t2 a_n1952_n3888# 1.26988f
C163 minus.n24 a_n1952_n3888# 0.490049f
C164 minus.n25 a_n1952_n3888# 0.009658f
C165 minus.t3 a_n1952_n3888# 1.26988f
C166 minus.n26 a_n1952_n3888# 0.487688f
C167 minus.n27 a_n1952_n3888# 0.292064f
C168 minus.n28 a_n1952_n3888# 2.02844f
.ends

