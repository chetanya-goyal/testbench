* NGSPICE file created from diffpair345.ext - technology: sky130A

.subckt diffpair345 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t20 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 drain_left.t10 plus.t1 source.t16 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 drain_right.t11 minus.t0 source.t4 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_left.t9 plus.t2 source.t19 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 source.t10 minus.t1 drain_right.t10 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 source.t9 minus.t2 drain_right.t9 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X6 source.t1 minus.t3 drain_right.t8 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X8 drain_left.t8 plus.t3 source.t12 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X9 source.t21 plus.t4 drain_left.t7 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X10 a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X11 source.t2 minus.t4 drain_right.t7 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X12 source.t22 plus.t5 drain_left.t6 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X13 source.t14 plus.t6 drain_left.t5 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X14 a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X15 drain_right.t6 minus.t5 source.t3 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X16 source.t13 plus.t7 drain_left.t4 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 drain_right.t5 minus.t6 source.t6 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X18 source.t8 minus.t7 drain_right.t4 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X19 drain_right.t3 minus.t8 source.t0 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X20 source.t23 plus.t8 drain_left.t3 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X21 drain_left.t2 plus.t9 source.t17 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X22 drain_right.t2 minus.t9 source.t7 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X23 source.t5 minus.t10 drain_right.t1 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X24 source.t15 plus.t10 drain_left.t1 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X25 drain_right.t0 minus.t11 source.t11 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X26 a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X27 drain_left.t0 plus.t11 source.t18 a_n1528_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
R0 plus.n2 plus.t4 1022.13
R1 plus.n13 plus.t11 1022.13
R2 plus.n17 plus.t9 1022.13
R3 plus.n28 plus.t8 1022.13
R4 plus.n3 plus.t1 992.92
R5 plus.n4 plus.t6 992.92
R6 plus.n10 plus.t0 992.92
R7 plus.n12 plus.t5 992.92
R8 plus.n19 plus.t7 992.92
R9 plus.n18 plus.t3 992.92
R10 plus.n25 plus.t10 992.92
R11 plus.n27 plus.t2 992.92
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 27.5899
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 10.9437
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n5 source.t21 51.0588
R53 source.n6 source.t0 51.0588
R54 source.n11 source.t2 51.0588
R55 source.n23 source.t7 51.0586
R56 source.n18 source.t5 51.0586
R57 source.n17 source.t17 51.0586
R58 source.n12 source.t23 51.0586
R59 source.n0 source.t18 51.0586
R60 source.n2 source.n1 48.8588
R61 source.n4 source.n3 48.8588
R62 source.n8 source.n7 48.8588
R63 source.n10 source.n9 48.8588
R64 source.n22 source.n21 48.8586
R65 source.n20 source.n19 48.8586
R66 source.n16 source.n15 48.8586
R67 source.n14 source.n13 48.8586
R68 source.n12 source.n11 19.515
R69 source.n24 source.n0 14.0021
R70 source.n24 source.n23 5.51343
R71 source.n21 source.t3 2.2005
R72 source.n21 source.t9 2.2005
R73 source.n19 source.t4 2.2005
R74 source.n19 source.t8 2.2005
R75 source.n15 source.t12 2.2005
R76 source.n15 source.t13 2.2005
R77 source.n13 source.t19 2.2005
R78 source.n13 source.t15 2.2005
R79 source.n1 source.t20 2.2005
R80 source.n1 source.t22 2.2005
R81 source.n3 source.t16 2.2005
R82 source.n3 source.t14 2.2005
R83 source.n7 source.t6 2.2005
R84 source.n7 source.t1 2.2005
R85 source.n9 source.t11 2.2005
R86 source.n9 source.t10 2.2005
R87 source.n11 source.n10 0.5005
R88 source.n10 source.n8 0.5005
R89 source.n8 source.n6 0.5005
R90 source.n5 source.n4 0.5005
R91 source.n4 source.n2 0.5005
R92 source.n2 source.n0 0.5005
R93 source.n14 source.n12 0.5005
R94 source.n16 source.n14 0.5005
R95 source.n17 source.n16 0.5005
R96 source.n20 source.n18 0.5005
R97 source.n22 source.n20 0.5005
R98 source.n23 source.n22 0.5005
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 66.0376
R103 drain_left.n3 drain_left.n2 65.982
R104 drain_left.n3 drain_left.n0 65.982
R105 drain_left.n6 drain_left.n5 65.5376
R106 drain_left.n8 drain_left.n7 65.5374
R107 drain_left.n3 drain_left.n1 65.5373
R108 drain_left drain_left.n3 27.5943
R109 drain_left drain_left.n8 6.15322
R110 drain_left.n1 drain_left.t1 2.2005
R111 drain_left.n1 drain_left.t8 2.2005
R112 drain_left.n2 drain_left.t4 2.2005
R113 drain_left.n2 drain_left.t2 2.2005
R114 drain_left.n0 drain_left.t3 2.2005
R115 drain_left.n0 drain_left.t9 2.2005
R116 drain_left.n7 drain_left.t6 2.2005
R117 drain_left.n7 drain_left.t0 2.2005
R118 drain_left.n5 drain_left.t5 2.2005
R119 drain_left.n5 drain_left.t11 2.2005
R120 drain_left.n4 drain_left.t7 2.2005
R121 drain_left.n4 drain_left.t10 2.2005
R122 drain_left.n8 drain_left.n6 0.5005
R123 minus.n13 minus.t4 1022.13
R124 minus.n2 minus.t8 1022.13
R125 minus.n28 minus.t9 1022.13
R126 minus.n17 minus.t10 1022.13
R127 minus.n12 minus.t11 992.92
R128 minus.n10 minus.t1 992.92
R129 minus.n3 minus.t6 992.92
R130 minus.n4 minus.t3 992.92
R131 minus.n27 minus.t2 992.92
R132 minus.n25 minus.t5 992.92
R133 minus.n19 minus.t7 992.92
R134 minus.n18 minus.t0 992.92
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 67.1884
R150 minus.n5 minus.n3 67.1884
R151 minus.n20 minus.n19 67.1884
R152 minus.n26 minus.n25 67.1884
R153 minus.n13 minus.n12 55.5035
R154 minus.n4 minus.n2 55.5035
R155 minus.n18 minus.n17 55.5035
R156 minus.n28 minus.n27 55.5035
R157 minus.n30 minus.n14 32.5725
R158 minus.n12 minus.n11 17.5278
R159 minus.n5 minus.n4 17.5278
R160 minus.n20 minus.n18 17.5278
R161 minus.n27 minus.n26 17.5278
R162 minus.n30 minus.n29 6.43611
R163 minus.n10 minus.n9 5.84292
R164 minus.n3 minus.n1 5.84292
R165 minus.n19 minus.n16 5.84292
R166 minus.n25 minus.n24 5.84292
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 66.0374
R177 drain_right.n3 drain_right.n2 65.982
R178 drain_right.n3 drain_right.n0 65.982
R179 drain_right.n6 drain_right.n5 65.5376
R180 drain_right.n8 drain_right.n7 65.5376
R181 drain_right.n3 drain_right.n1 65.5373
R182 drain_right drain_right.n3 27.0411
R183 drain_right drain_right.n8 6.15322
R184 drain_right.n1 drain_right.t4 2.2005
R185 drain_right.n1 drain_right.t6 2.2005
R186 drain_right.n2 drain_right.t9 2.2005
R187 drain_right.n2 drain_right.t2 2.2005
R188 drain_right.n0 drain_right.t1 2.2005
R189 drain_right.n0 drain_right.t11 2.2005
R190 drain_right.n4 drain_right.t8 2.2005
R191 drain_right.n4 drain_right.t3 2.2005
R192 drain_right.n5 drain_right.t10 2.2005
R193 drain_right.n5 drain_right.t5 2.2005
R194 drain_right.n7 drain_right.t7 2.2005
R195 drain_right.n7 drain_right.t0 2.2005
R196 drain_right.n8 drain_right.n6 0.5005
C0 minus plus 4.50667f
C1 source drain_right 19.752802f
C2 source minus 2.88691f
C3 source plus 2.90094f
C4 drain_right drain_left 0.751086f
C5 minus drain_left 0.171004f
C6 plus drain_left 3.31696f
C7 minus drain_right 3.17079f
C8 plus drain_right 0.300071f
C9 source drain_left 19.753399f
C10 drain_right a_n1528_n2688# 5.56649f
C11 drain_left a_n1528_n2688# 5.80769f
C12 source a_n1528_n2688# 6.9337f
C13 minus a_n1528_n2688# 5.72034f
C14 plus a_n1528_n2688# 7.51054f
C15 drain_right.t1 a_n1528_n2688# 0.251038f
C16 drain_right.t11 a_n1528_n2688# 0.251038f
C17 drain_right.n0 a_n1528_n2688# 2.19848f
C18 drain_right.t4 a_n1528_n2688# 0.251038f
C19 drain_right.t6 a_n1528_n2688# 0.251038f
C20 drain_right.n1 a_n1528_n2688# 2.19575f
C21 drain_right.t9 a_n1528_n2688# 0.251038f
C22 drain_right.t2 a_n1528_n2688# 0.251038f
C23 drain_right.n2 a_n1528_n2688# 2.19848f
C24 drain_right.n3 a_n1528_n2688# 2.44818f
C25 drain_right.t8 a_n1528_n2688# 0.251038f
C26 drain_right.t3 a_n1528_n2688# 0.251038f
C27 drain_right.n4 a_n1528_n2688# 2.19885f
C28 drain_right.t10 a_n1528_n2688# 0.251038f
C29 drain_right.t5 a_n1528_n2688# 0.251038f
C30 drain_right.n5 a_n1528_n2688# 2.19575f
C31 drain_right.n6 a_n1528_n2688# 0.804054f
C32 drain_right.t7 a_n1528_n2688# 0.251038f
C33 drain_right.t0 a_n1528_n2688# 0.251038f
C34 drain_right.n7 a_n1528_n2688# 2.19575f
C35 drain_right.n8 a_n1528_n2688# 0.687825f
C36 minus.n0 a_n1528_n2688# 0.053786f
C37 minus.t4 a_n1528_n2688# 0.347045f
C38 minus.t11 a_n1528_n2688# 0.342921f
C39 minus.t1 a_n1528_n2688# 0.342921f
C40 minus.n1 a_n1528_n2688# 0.019169f
C41 minus.t8 a_n1528_n2688# 0.347045f
C42 minus.n2 a_n1528_n2688# 0.160744f
C43 minus.t6 a_n1528_n2688# 0.342921f
C44 minus.n3 a_n1528_n2688# 0.145961f
C45 minus.t3 a_n1528_n2688# 0.342921f
C46 minus.n4 a_n1528_n2688# 0.145961f
C47 minus.n5 a_n1528_n2688# 0.020496f
C48 minus.n6 a_n1528_n2688# 0.112478f
C49 minus.n7 a_n1528_n2688# 0.053786f
C50 minus.n8 a_n1528_n2688# 0.053786f
C51 minus.n9 a_n1528_n2688# 0.019169f
C52 minus.n10 a_n1528_n2688# 0.145961f
C53 minus.n11 a_n1528_n2688# 0.020496f
C54 minus.n12 a_n1528_n2688# 0.145961f
C55 minus.n13 a_n1528_n2688# 0.160675f
C56 minus.n14 a_n1528_n2688# 1.60275f
C57 minus.n15 a_n1528_n2688# 0.053786f
C58 minus.t2 a_n1528_n2688# 0.342921f
C59 minus.t5 a_n1528_n2688# 0.342921f
C60 minus.n16 a_n1528_n2688# 0.019169f
C61 minus.t10 a_n1528_n2688# 0.347045f
C62 minus.n17 a_n1528_n2688# 0.160744f
C63 minus.t0 a_n1528_n2688# 0.342921f
C64 minus.n18 a_n1528_n2688# 0.145961f
C65 minus.t7 a_n1528_n2688# 0.342921f
C66 minus.n19 a_n1528_n2688# 0.145961f
C67 minus.n20 a_n1528_n2688# 0.020496f
C68 minus.n21 a_n1528_n2688# 0.112478f
C69 minus.n22 a_n1528_n2688# 0.053786f
C70 minus.n23 a_n1528_n2688# 0.053786f
C71 minus.n24 a_n1528_n2688# 0.019169f
C72 minus.n25 a_n1528_n2688# 0.145961f
C73 minus.n26 a_n1528_n2688# 0.020496f
C74 minus.n27 a_n1528_n2688# 0.145961f
C75 minus.t9 a_n1528_n2688# 0.347045f
C76 minus.n28 a_n1528_n2688# 0.160675f
C77 minus.n29 a_n1528_n2688# 0.34352f
C78 minus.n30 a_n1528_n2688# 1.97f
C79 drain_left.t3 a_n1528_n2688# 0.250625f
C80 drain_left.t9 a_n1528_n2688# 0.250625f
C81 drain_left.n0 a_n1528_n2688# 2.19486f
C82 drain_left.t1 a_n1528_n2688# 0.250625f
C83 drain_left.t8 a_n1528_n2688# 0.250625f
C84 drain_left.n1 a_n1528_n2688# 2.19213f
C85 drain_left.t4 a_n1528_n2688# 0.250625f
C86 drain_left.t2 a_n1528_n2688# 0.250625f
C87 drain_left.n2 a_n1528_n2688# 2.19486f
C88 drain_left.n3 a_n1528_n2688# 2.5171f
C89 drain_left.t7 a_n1528_n2688# 0.250625f
C90 drain_left.t10 a_n1528_n2688# 0.250625f
C91 drain_left.n4 a_n1528_n2688# 2.19524f
C92 drain_left.t5 a_n1528_n2688# 0.250625f
C93 drain_left.t11 a_n1528_n2688# 0.250625f
C94 drain_left.n5 a_n1528_n2688# 2.19214f
C95 drain_left.n6 a_n1528_n2688# 0.802722f
C96 drain_left.t6 a_n1528_n2688# 0.250625f
C97 drain_left.t0 a_n1528_n2688# 0.250625f
C98 drain_left.n7 a_n1528_n2688# 2.19213f
C99 drain_left.n8 a_n1528_n2688# 0.686703f
C100 source.t18 a_n1528_n2688# 2.16119f
C101 source.n0 a_n1528_n2688# 1.23612f
C102 source.t20 a_n1528_n2688# 0.202673f
C103 source.t22 a_n1528_n2688# 0.202673f
C104 source.n1 a_n1528_n2688# 1.69664f
C105 source.n2 a_n1528_n2688# 0.357421f
C106 source.t16 a_n1528_n2688# 0.202673f
C107 source.t14 a_n1528_n2688# 0.202673f
C108 source.n3 a_n1528_n2688# 1.69664f
C109 source.n4 a_n1528_n2688# 0.357421f
C110 source.t21 a_n1528_n2688# 2.1612f
C111 source.n5 a_n1528_n2688# 0.442839f
C112 source.t0 a_n1528_n2688# 2.1612f
C113 source.n6 a_n1528_n2688# 0.442839f
C114 source.t6 a_n1528_n2688# 0.202673f
C115 source.t1 a_n1528_n2688# 0.202673f
C116 source.n7 a_n1528_n2688# 1.69664f
C117 source.n8 a_n1528_n2688# 0.357421f
C118 source.t11 a_n1528_n2688# 0.202673f
C119 source.t10 a_n1528_n2688# 0.202673f
C120 source.n9 a_n1528_n2688# 1.69664f
C121 source.n10 a_n1528_n2688# 0.357421f
C122 source.t2 a_n1528_n2688# 2.1612f
C123 source.n11 a_n1528_n2688# 1.64888f
C124 source.t23 a_n1528_n2688# 2.16119f
C125 source.n12 a_n1528_n2688# 1.64889f
C126 source.t19 a_n1528_n2688# 0.202673f
C127 source.t15 a_n1528_n2688# 0.202673f
C128 source.n13 a_n1528_n2688# 1.69664f
C129 source.n14 a_n1528_n2688# 0.357426f
C130 source.t12 a_n1528_n2688# 0.202673f
C131 source.t13 a_n1528_n2688# 0.202673f
C132 source.n15 a_n1528_n2688# 1.69664f
C133 source.n16 a_n1528_n2688# 0.357426f
C134 source.t17 a_n1528_n2688# 2.16119f
C135 source.n17 a_n1528_n2688# 0.442844f
C136 source.t5 a_n1528_n2688# 2.16119f
C137 source.n18 a_n1528_n2688# 0.442844f
C138 source.t4 a_n1528_n2688# 0.202673f
C139 source.t8 a_n1528_n2688# 0.202673f
C140 source.n19 a_n1528_n2688# 1.69664f
C141 source.n20 a_n1528_n2688# 0.357426f
C142 source.t3 a_n1528_n2688# 0.202673f
C143 source.t9 a_n1528_n2688# 0.202673f
C144 source.n21 a_n1528_n2688# 1.69664f
C145 source.n22 a_n1528_n2688# 0.357426f
C146 source.t7 a_n1528_n2688# 2.16119f
C147 source.n23 a_n1528_n2688# 0.600541f
C148 source.n24 a_n1528_n2688# 1.48139f
C149 plus.n0 a_n1528_n2688# 0.054857f
C150 plus.t5 a_n1528_n2688# 0.349745f
C151 plus.t0 a_n1528_n2688# 0.349745f
C152 plus.n1 a_n1528_n2688# 0.019551f
C153 plus.t4 a_n1528_n2688# 0.353951f
C154 plus.n2 a_n1528_n2688# 0.163942f
C155 plus.t1 a_n1528_n2688# 0.349745f
C156 plus.n3 a_n1528_n2688# 0.148866f
C157 plus.t6 a_n1528_n2688# 0.349745f
C158 plus.n4 a_n1528_n2688# 0.148866f
C159 plus.n5 a_n1528_n2688# 0.020903f
C160 plus.n6 a_n1528_n2688# 0.114716f
C161 plus.n7 a_n1528_n2688# 0.054857f
C162 plus.n8 a_n1528_n2688# 0.054857f
C163 plus.n9 a_n1528_n2688# 0.019551f
C164 plus.n10 a_n1528_n2688# 0.148866f
C165 plus.n11 a_n1528_n2688# 0.020903f
C166 plus.n12 a_n1528_n2688# 0.148866f
C167 plus.t11 a_n1528_n2688# 0.353951f
C168 plus.n13 a_n1528_n2688# 0.163872f
C169 plus.n14 a_n1528_n2688# 0.530337f
C170 plus.n15 a_n1528_n2688# 0.054857f
C171 plus.t8 a_n1528_n2688# 0.353951f
C172 plus.t2 a_n1528_n2688# 0.349745f
C173 plus.t10 a_n1528_n2688# 0.349745f
C174 plus.n16 a_n1528_n2688# 0.019551f
C175 plus.t9 a_n1528_n2688# 0.353951f
C176 plus.n17 a_n1528_n2688# 0.163942f
C177 plus.t3 a_n1528_n2688# 0.349745f
C178 plus.n18 a_n1528_n2688# 0.148866f
C179 plus.t7 a_n1528_n2688# 0.349745f
C180 plus.n19 a_n1528_n2688# 0.148866f
C181 plus.n20 a_n1528_n2688# 0.020903f
C182 plus.n21 a_n1528_n2688# 0.114716f
C183 plus.n22 a_n1528_n2688# 0.054857f
C184 plus.n23 a_n1528_n2688# 0.054857f
C185 plus.n24 a_n1528_n2688# 0.019551f
C186 plus.n25 a_n1528_n2688# 0.148866f
C187 plus.n26 a_n1528_n2688# 0.020903f
C188 plus.n27 a_n1528_n2688# 0.148866f
C189 plus.n28 a_n1528_n2688# 0.163872f
C190 plus.n29 a_n1528_n2688# 1.42297f
.ends

