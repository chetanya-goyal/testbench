* NGSPICE file created from diffpair125.ext - technology: sky130A

.subckt diffpair125 minus drain_right drain_left source plus
X0 a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X1 drain_right.t11 minus.t0 source.t17 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X2 drain_right.t10 minus.t1 source.t10 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X3 source.t21 plus.t0 drain_left.t11 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X4 source.t22 plus.t1 drain_left.t10 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X5 source.t8 minus.t2 drain_right.t9 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X6 source.t2 plus.t2 drain_left.t9 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X7 source.t1 plus.t3 drain_left.t8 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X8 drain_right.t8 minus.t3 source.t9 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X9 drain_right.t7 minus.t4 source.t11 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X10 source.t16 minus.t5 drain_right.t6 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 drain_left.t7 plus.t4 source.t6 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X12 drain_left.t6 plus.t5 source.t3 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X13 source.t19 minus.t6 drain_right.t5 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X14 a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X15 drain_right.t4 minus.t7 source.t14 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X16 a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X17 a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X18 drain_left.t5 plus.t6 source.t5 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X19 source.t13 minus.t8 drain_right.t3 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X20 source.t12 minus.t9 drain_right.t2 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X21 drain_left.t4 plus.t7 source.t4 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X22 source.t15 minus.t10 drain_right.t1 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X23 source.t20 plus.t8 drain_left.t3 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X24 drain_right.t0 minus.t11 source.t18 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X25 source.t7 plus.t9 drain_left.t2 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X26 drain_left.t1 plus.t10 source.t0 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X27 drain_left.t0 plus.t11 source.t23 a_n1878_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
R0 minus.n3 minus.t7 201.636
R1 minus.n17 minus.t10 201.636
R2 minus.n4 minus.t2 174.966
R3 minus.n5 minus.t4 174.966
R4 minus.n1 minus.t9 174.966
R5 minus.n10 minus.t3 174.966
R6 minus.n12 minus.t6 174.966
R7 minus.n18 minus.t0 174.966
R8 minus.n19 minus.t8 174.966
R9 minus.n15 minus.t11 174.966
R10 minus.n24 minus.t5 174.966
R11 minus.n26 minus.t1 174.966
R12 minus.n13 minus.n12 161.3
R13 minus.n11 minus.n0 161.3
R14 minus.n10 minus.n9 161.3
R15 minus.n8 minus.n1 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n2 161.3
R18 minus.n27 minus.n26 161.3
R19 minus.n25 minus.n14 161.3
R20 minus.n24 minus.n23 161.3
R21 minus.n22 minus.n15 161.3
R22 minus.n21 minus.n20 161.3
R23 minus.n19 minus.n16 161.3
R24 minus.n5 minus.n4 48.2005
R25 minus.n10 minus.n1 48.2005
R26 minus.n19 minus.n18 48.2005
R27 minus.n24 minus.n15 48.2005
R28 minus.n12 minus.n11 47.4702
R29 minus.n26 minus.n25 47.4702
R30 minus.n3 minus.n2 45.1192
R31 minus.n17 minus.n16 45.1192
R32 minus.n28 minus.n13 28.6899
R33 minus.n6 minus.n1 24.1005
R34 minus.n6 minus.n5 24.1005
R35 minus.n20 minus.n19 24.1005
R36 minus.n20 minus.n15 24.1005
R37 minus.n4 minus.n3 13.6377
R38 minus.n18 minus.n17 13.6377
R39 minus.n28 minus.n27 6.5308
R40 minus.n11 minus.n10 0.730803
R41 minus.n25 minus.n24 0.730803
R42 minus.n13 minus.n0 0.189894
R43 minus.n9 minus.n0 0.189894
R44 minus.n9 minus.n8 0.189894
R45 minus.n8 minus.n7 0.189894
R46 minus.n7 minus.n2 0.189894
R47 minus.n21 minus.n16 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n14 0.189894
R51 minus.n27 minus.n14 0.189894
R52 minus minus.n28 0.188
R53 source.n74 source.n72 289.615
R54 source.n62 source.n60 289.615
R55 source.n54 source.n52 289.615
R56 source.n42 source.n40 289.615
R57 source.n2 source.n0 289.615
R58 source.n14 source.n12 289.615
R59 source.n22 source.n20 289.615
R60 source.n34 source.n32 289.615
R61 source.n75 source.n74 185
R62 source.n63 source.n62 185
R63 source.n55 source.n54 185
R64 source.n43 source.n42 185
R65 source.n3 source.n2 185
R66 source.n15 source.n14 185
R67 source.n23 source.n22 185
R68 source.n35 source.n34 185
R69 source.t10 source.n73 167.117
R70 source.t15 source.n61 167.117
R71 source.t0 source.n53 167.117
R72 source.t21 source.n41 167.117
R73 source.t23 source.n1 167.117
R74 source.t2 source.n13 167.117
R75 source.t14 source.n21 167.117
R76 source.t19 source.n33 167.117
R77 source.n9 source.n8 84.1169
R78 source.n11 source.n10 84.1169
R79 source.n29 source.n28 84.1169
R80 source.n31 source.n30 84.1169
R81 source.n71 source.n70 84.1168
R82 source.n69 source.n68 84.1168
R83 source.n51 source.n50 84.1168
R84 source.n49 source.n48 84.1168
R85 source.n74 source.t10 52.3082
R86 source.n62 source.t15 52.3082
R87 source.n54 source.t0 52.3082
R88 source.n42 source.t21 52.3082
R89 source.n2 source.t23 52.3082
R90 source.n14 source.t2 52.3082
R91 source.n22 source.t14 52.3082
R92 source.n34 source.t19 52.3082
R93 source.n79 source.n78 31.4096
R94 source.n67 source.n66 31.4096
R95 source.n59 source.n58 31.4096
R96 source.n47 source.n46 31.4096
R97 source.n7 source.n6 31.4096
R98 source.n19 source.n18 31.4096
R99 source.n27 source.n26 31.4096
R100 source.n39 source.n38 31.4096
R101 source.n47 source.n39 14.4275
R102 source.n70 source.t18 9.9005
R103 source.n70 source.t16 9.9005
R104 source.n68 source.t17 9.9005
R105 source.n68 source.t13 9.9005
R106 source.n50 source.t4 9.9005
R107 source.n50 source.t22 9.9005
R108 source.n48 source.t3 9.9005
R109 source.n48 source.t1 9.9005
R110 source.n8 source.t6 9.9005
R111 source.n8 source.t20 9.9005
R112 source.n10 source.t5 9.9005
R113 source.n10 source.t7 9.9005
R114 source.n28 source.t11 9.9005
R115 source.n28 source.t8 9.9005
R116 source.n30 source.t9 9.9005
R117 source.n30 source.t12 9.9005
R118 source.n75 source.n73 9.71174
R119 source.n63 source.n61 9.71174
R120 source.n55 source.n53 9.71174
R121 source.n43 source.n41 9.71174
R122 source.n3 source.n1 9.71174
R123 source.n15 source.n13 9.71174
R124 source.n23 source.n21 9.71174
R125 source.n35 source.n33 9.71174
R126 source.n78 source.n77 9.45567
R127 source.n66 source.n65 9.45567
R128 source.n58 source.n57 9.45567
R129 source.n46 source.n45 9.45567
R130 source.n6 source.n5 9.45567
R131 source.n18 source.n17 9.45567
R132 source.n26 source.n25 9.45567
R133 source.n38 source.n37 9.45567
R134 source.n77 source.n76 9.3005
R135 source.n65 source.n64 9.3005
R136 source.n57 source.n56 9.3005
R137 source.n45 source.n44 9.3005
R138 source.n5 source.n4 9.3005
R139 source.n17 source.n16 9.3005
R140 source.n25 source.n24 9.3005
R141 source.n37 source.n36 9.3005
R142 source.n80 source.n7 8.8068
R143 source.n78 source.n72 8.14595
R144 source.n66 source.n60 8.14595
R145 source.n58 source.n52 8.14595
R146 source.n46 source.n40 8.14595
R147 source.n6 source.n0 8.14595
R148 source.n18 source.n12 8.14595
R149 source.n26 source.n20 8.14595
R150 source.n38 source.n32 8.14595
R151 source.n76 source.n75 7.3702
R152 source.n64 source.n63 7.3702
R153 source.n56 source.n55 7.3702
R154 source.n44 source.n43 7.3702
R155 source.n4 source.n3 7.3702
R156 source.n16 source.n15 7.3702
R157 source.n24 source.n23 7.3702
R158 source.n36 source.n35 7.3702
R159 source.n76 source.n72 5.81868
R160 source.n64 source.n60 5.81868
R161 source.n56 source.n52 5.81868
R162 source.n44 source.n40 5.81868
R163 source.n4 source.n0 5.81868
R164 source.n16 source.n12 5.81868
R165 source.n24 source.n20 5.81868
R166 source.n36 source.n32 5.81868
R167 source.n80 source.n79 5.62119
R168 source.n77 source.n73 3.44771
R169 source.n65 source.n61 3.44771
R170 source.n57 source.n53 3.44771
R171 source.n45 source.n41 3.44771
R172 source.n5 source.n1 3.44771
R173 source.n17 source.n13 3.44771
R174 source.n25 source.n21 3.44771
R175 source.n37 source.n33 3.44771
R176 source.n39 source.n31 0.716017
R177 source.n31 source.n29 0.716017
R178 source.n29 source.n27 0.716017
R179 source.n19 source.n11 0.716017
R180 source.n11 source.n9 0.716017
R181 source.n9 source.n7 0.716017
R182 source.n49 source.n47 0.716017
R183 source.n51 source.n49 0.716017
R184 source.n59 source.n51 0.716017
R185 source.n69 source.n67 0.716017
R186 source.n71 source.n69 0.716017
R187 source.n79 source.n71 0.716017
R188 source.n27 source.n19 0.470328
R189 source.n67 source.n59 0.470328
R190 source source.n80 0.188
R191 drain_right.n6 drain_right.n4 101.511
R192 drain_right.n3 drain_right.n2 101.456
R193 drain_right.n3 drain_right.n0 101.456
R194 drain_right.n6 drain_right.n5 100.796
R195 drain_right.n8 drain_right.n7 100.796
R196 drain_right.n3 drain_right.n1 100.796
R197 drain_right drain_right.n3 22.8157
R198 drain_right.n1 drain_right.t3 9.9005
R199 drain_right.n1 drain_right.t0 9.9005
R200 drain_right.n2 drain_right.t6 9.9005
R201 drain_right.n2 drain_right.t10 9.9005
R202 drain_right.n0 drain_right.t1 9.9005
R203 drain_right.n0 drain_right.t11 9.9005
R204 drain_right.n4 drain_right.t9 9.9005
R205 drain_right.n4 drain_right.t4 9.9005
R206 drain_right.n5 drain_right.t2 9.9005
R207 drain_right.n5 drain_right.t7 9.9005
R208 drain_right.n7 drain_right.t5 9.9005
R209 drain_right.n7 drain_right.t8 9.9005
R210 drain_right drain_right.n8 6.36873
R211 drain_right.n8 drain_right.n6 0.716017
R212 plus.n5 plus.t2 201.636
R213 plus.n19 plus.t10 201.636
R214 plus.n12 plus.t11 174.966
R215 plus.n10 plus.t8 174.966
R216 plus.n9 plus.t4 174.966
R217 plus.n3 plus.t9 174.966
R218 plus.n4 plus.t6 174.966
R219 plus.n26 plus.t0 174.966
R220 plus.n24 plus.t5 174.966
R221 plus.n23 plus.t3 174.966
R222 plus.n17 plus.t7 174.966
R223 plus.n18 plus.t1 174.966
R224 plus.n6 plus.n3 161.3
R225 plus.n8 plus.n7 161.3
R226 plus.n9 plus.n2 161.3
R227 plus.n10 plus.n1 161.3
R228 plus.n11 plus.n0 161.3
R229 plus.n13 plus.n12 161.3
R230 plus.n20 plus.n17 161.3
R231 plus.n22 plus.n21 161.3
R232 plus.n23 plus.n16 161.3
R233 plus.n24 plus.n15 161.3
R234 plus.n25 plus.n14 161.3
R235 plus.n27 plus.n26 161.3
R236 plus.n10 plus.n9 48.2005
R237 plus.n4 plus.n3 48.2005
R238 plus.n24 plus.n23 48.2005
R239 plus.n18 plus.n17 48.2005
R240 plus.n12 plus.n11 47.4702
R241 plus.n26 plus.n25 47.4702
R242 plus.n6 plus.n5 45.1192
R243 plus.n20 plus.n19 45.1192
R244 plus plus.n27 26.3589
R245 plus.n8 plus.n3 24.1005
R246 plus.n9 plus.n8 24.1005
R247 plus.n23 plus.n22 24.1005
R248 plus.n22 plus.n17 24.1005
R249 plus.n5 plus.n4 13.6377
R250 plus.n19 plus.n18 13.6377
R251 plus plus.n13 8.38686
R252 plus.n11 plus.n10 0.730803
R253 plus.n25 plus.n24 0.730803
R254 plus.n7 plus.n6 0.189894
R255 plus.n7 plus.n2 0.189894
R256 plus.n2 plus.n1 0.189894
R257 plus.n1 plus.n0 0.189894
R258 plus.n13 plus.n0 0.189894
R259 plus.n27 plus.n14 0.189894
R260 plus.n15 plus.n14 0.189894
R261 plus.n16 plus.n15 0.189894
R262 plus.n21 plus.n16 0.189894
R263 plus.n21 plus.n20 0.189894
R264 drain_left.n6 drain_left.n4 101.511
R265 drain_left.n3 drain_left.n2 101.456
R266 drain_left.n3 drain_left.n0 101.456
R267 drain_left.n8 drain_left.n7 100.796
R268 drain_left.n6 drain_left.n5 100.796
R269 drain_left.n3 drain_left.n1 100.796
R270 drain_left drain_left.n3 23.3689
R271 drain_left.n1 drain_left.t8 9.9005
R272 drain_left.n1 drain_left.t4 9.9005
R273 drain_left.n2 drain_left.t10 9.9005
R274 drain_left.n2 drain_left.t1 9.9005
R275 drain_left.n0 drain_left.t11 9.9005
R276 drain_left.n0 drain_left.t6 9.9005
R277 drain_left.n7 drain_left.t3 9.9005
R278 drain_left.n7 drain_left.t0 9.9005
R279 drain_left.n5 drain_left.t2 9.9005
R280 drain_left.n5 drain_left.t7 9.9005
R281 drain_left.n4 drain_left.t9 9.9005
R282 drain_left.n4 drain_left.t5 9.9005
R283 drain_left drain_left.n8 6.36873
R284 drain_left.n8 drain_left.n6 0.716017
C0 plus drain_right 0.343944f
C1 drain_left drain_right 0.936595f
C2 plus drain_left 1.65097f
C3 minus drain_right 1.46842f
C4 plus minus 3.64913f
C5 drain_left minus 0.177489f
C6 drain_right source 5.17326f
C7 plus source 1.76591f
C8 drain_left source 5.17229f
C9 minus source 1.75195f
C10 drain_right a_n1878_n1288# 3.63748f
C11 drain_left a_n1878_n1288# 3.87974f
C12 source a_n1878_n1288# 3.110602f
C13 minus a_n1878_n1288# 6.548949f
C14 plus a_n1878_n1288# 7.093791f
C15 drain_left.t11 a_n1878_n1288# 0.033537f
C16 drain_left.t6 a_n1878_n1288# 0.033537f
C17 drain_left.n0 a_n1878_n1288# 0.212422f
C18 drain_left.t8 a_n1878_n1288# 0.033537f
C19 drain_left.t4 a_n1878_n1288# 0.033537f
C20 drain_left.n1 a_n1878_n1288# 0.210692f
C21 drain_left.t10 a_n1878_n1288# 0.033537f
C22 drain_left.t1 a_n1878_n1288# 0.033537f
C23 drain_left.n2 a_n1878_n1288# 0.212422f
C24 drain_left.n3 a_n1878_n1288# 1.36361f
C25 drain_left.t9 a_n1878_n1288# 0.033537f
C26 drain_left.t5 a_n1878_n1288# 0.033537f
C27 drain_left.n4 a_n1878_n1288# 0.212588f
C28 drain_left.t2 a_n1878_n1288# 0.033537f
C29 drain_left.t7 a_n1878_n1288# 0.033537f
C30 drain_left.n5 a_n1878_n1288# 0.210693f
C31 drain_left.n6 a_n1878_n1288# 0.527178f
C32 drain_left.t3 a_n1878_n1288# 0.033537f
C33 drain_left.t0 a_n1878_n1288# 0.033537f
C34 drain_left.n7 a_n1878_n1288# 0.210693f
C35 drain_left.n8 a_n1878_n1288# 0.442572f
C36 plus.n0 a_n1878_n1288# 0.025532f
C37 plus.t11 a_n1878_n1288# 0.079067f
C38 plus.t8 a_n1878_n1288# 0.079067f
C39 plus.n1 a_n1878_n1288# 0.025532f
C40 plus.t4 a_n1878_n1288# 0.079067f
C41 plus.n2 a_n1878_n1288# 0.025532f
C42 plus.t9 a_n1878_n1288# 0.079067f
C43 plus.n3 a_n1878_n1288# 0.059552f
C44 plus.t6 a_n1878_n1288# 0.079067f
C45 plus.n4 a_n1878_n1288# 0.06263f
C46 plus.t2 a_n1878_n1288# 0.086604f
C47 plus.n5 a_n1878_n1288# 0.050043f
C48 plus.n6 a_n1878_n1288# 0.103984f
C49 plus.n7 a_n1878_n1288# 0.025532f
C50 plus.n8 a_n1878_n1288# 0.005794f
C51 plus.n9 a_n1878_n1288# 0.059552f
C52 plus.n10 a_n1878_n1288# 0.057033f
C53 plus.n11 a_n1878_n1288# 0.005794f
C54 plus.n12 a_n1878_n1288# 0.056876f
C55 plus.n13 a_n1878_n1288# 0.184479f
C56 plus.n14 a_n1878_n1288# 0.025532f
C57 plus.t0 a_n1878_n1288# 0.079067f
C58 plus.n15 a_n1878_n1288# 0.025532f
C59 plus.t5 a_n1878_n1288# 0.079067f
C60 plus.n16 a_n1878_n1288# 0.025532f
C61 plus.t3 a_n1878_n1288# 0.079067f
C62 plus.t7 a_n1878_n1288# 0.079067f
C63 plus.n17 a_n1878_n1288# 0.059552f
C64 plus.t10 a_n1878_n1288# 0.086604f
C65 plus.t1 a_n1878_n1288# 0.079067f
C66 plus.n18 a_n1878_n1288# 0.06263f
C67 plus.n19 a_n1878_n1288# 0.050043f
C68 plus.n20 a_n1878_n1288# 0.103984f
C69 plus.n21 a_n1878_n1288# 0.025532f
C70 plus.n22 a_n1878_n1288# 0.005794f
C71 plus.n23 a_n1878_n1288# 0.059552f
C72 plus.n24 a_n1878_n1288# 0.057033f
C73 plus.n25 a_n1878_n1288# 0.005794f
C74 plus.n26 a_n1878_n1288# 0.056876f
C75 plus.n27 a_n1878_n1288# 0.587699f
C76 drain_right.t1 a_n1878_n1288# 0.034081f
C77 drain_right.t11 a_n1878_n1288# 0.034081f
C78 drain_right.n0 a_n1878_n1288# 0.215868f
C79 drain_right.t3 a_n1878_n1288# 0.034081f
C80 drain_right.t0 a_n1878_n1288# 0.034081f
C81 drain_right.n1 a_n1878_n1288# 0.21411f
C82 drain_right.t6 a_n1878_n1288# 0.034081f
C83 drain_right.t10 a_n1878_n1288# 0.034081f
C84 drain_right.n2 a_n1878_n1288# 0.215868f
C85 drain_right.n3 a_n1878_n1288# 1.3435f
C86 drain_right.t9 a_n1878_n1288# 0.034081f
C87 drain_right.t4 a_n1878_n1288# 0.034081f
C88 drain_right.n4 a_n1878_n1288# 0.216037f
C89 drain_right.t2 a_n1878_n1288# 0.034081f
C90 drain_right.t7 a_n1878_n1288# 0.034081f
C91 drain_right.n5 a_n1878_n1288# 0.214111f
C92 drain_right.n6 a_n1878_n1288# 0.53573f
C93 drain_right.t5 a_n1878_n1288# 0.034081f
C94 drain_right.t8 a_n1878_n1288# 0.034081f
C95 drain_right.n7 a_n1878_n1288# 0.214111f
C96 drain_right.n8 a_n1878_n1288# 0.449752f
C97 source.n0 a_n1878_n1288# 0.032109f
C98 source.n1 a_n1878_n1288# 0.071045f
C99 source.t23 a_n1878_n1288# 0.053316f
C100 source.n2 a_n1878_n1288# 0.055603f
C101 source.n3 a_n1878_n1288# 0.017924f
C102 source.n4 a_n1878_n1288# 0.011821f
C103 source.n5 a_n1878_n1288# 0.156601f
C104 source.n6 a_n1878_n1288# 0.035199f
C105 source.n7 a_n1878_n1288# 0.353837f
C106 source.t6 a_n1878_n1288# 0.034769f
C107 source.t20 a_n1878_n1288# 0.034769f
C108 source.n8 a_n1878_n1288# 0.185873f
C109 source.n9 a_n1878_n1288# 0.272473f
C110 source.t5 a_n1878_n1288# 0.034769f
C111 source.t7 a_n1878_n1288# 0.034769f
C112 source.n10 a_n1878_n1288# 0.185873f
C113 source.n11 a_n1878_n1288# 0.272473f
C114 source.n12 a_n1878_n1288# 0.032109f
C115 source.n13 a_n1878_n1288# 0.071045f
C116 source.t2 a_n1878_n1288# 0.053316f
C117 source.n14 a_n1878_n1288# 0.055603f
C118 source.n15 a_n1878_n1288# 0.017924f
C119 source.n16 a_n1878_n1288# 0.011821f
C120 source.n17 a_n1878_n1288# 0.156601f
C121 source.n18 a_n1878_n1288# 0.035199f
C122 source.n19 a_n1878_n1288# 0.102135f
C123 source.n20 a_n1878_n1288# 0.032109f
C124 source.n21 a_n1878_n1288# 0.071045f
C125 source.t14 a_n1878_n1288# 0.053316f
C126 source.n22 a_n1878_n1288# 0.055603f
C127 source.n23 a_n1878_n1288# 0.017924f
C128 source.n24 a_n1878_n1288# 0.011821f
C129 source.n25 a_n1878_n1288# 0.156601f
C130 source.n26 a_n1878_n1288# 0.035199f
C131 source.n27 a_n1878_n1288# 0.102135f
C132 source.t11 a_n1878_n1288# 0.034769f
C133 source.t8 a_n1878_n1288# 0.034769f
C134 source.n28 a_n1878_n1288# 0.185873f
C135 source.n29 a_n1878_n1288# 0.272473f
C136 source.t9 a_n1878_n1288# 0.034769f
C137 source.t12 a_n1878_n1288# 0.034769f
C138 source.n30 a_n1878_n1288# 0.185873f
C139 source.n31 a_n1878_n1288# 0.272473f
C140 source.n32 a_n1878_n1288# 0.032109f
C141 source.n33 a_n1878_n1288# 0.071045f
C142 source.t19 a_n1878_n1288# 0.053316f
C143 source.n34 a_n1878_n1288# 0.055603f
C144 source.n35 a_n1878_n1288# 0.017924f
C145 source.n36 a_n1878_n1288# 0.011821f
C146 source.n37 a_n1878_n1288# 0.156601f
C147 source.n38 a_n1878_n1288# 0.035199f
C148 source.n39 a_n1878_n1288# 0.561692f
C149 source.n40 a_n1878_n1288# 0.032109f
C150 source.n41 a_n1878_n1288# 0.071045f
C151 source.t21 a_n1878_n1288# 0.053316f
C152 source.n42 a_n1878_n1288# 0.055603f
C153 source.n43 a_n1878_n1288# 0.017924f
C154 source.n44 a_n1878_n1288# 0.011821f
C155 source.n45 a_n1878_n1288# 0.156601f
C156 source.n46 a_n1878_n1288# 0.035199f
C157 source.n47 a_n1878_n1288# 0.561692f
C158 source.t3 a_n1878_n1288# 0.034769f
C159 source.t1 a_n1878_n1288# 0.034769f
C160 source.n48 a_n1878_n1288# 0.185871f
C161 source.n49 a_n1878_n1288# 0.272474f
C162 source.t4 a_n1878_n1288# 0.034769f
C163 source.t22 a_n1878_n1288# 0.034769f
C164 source.n50 a_n1878_n1288# 0.185871f
C165 source.n51 a_n1878_n1288# 0.272474f
C166 source.n52 a_n1878_n1288# 0.032109f
C167 source.n53 a_n1878_n1288# 0.071045f
C168 source.t0 a_n1878_n1288# 0.053316f
C169 source.n54 a_n1878_n1288# 0.055603f
C170 source.n55 a_n1878_n1288# 0.017924f
C171 source.n56 a_n1878_n1288# 0.011821f
C172 source.n57 a_n1878_n1288# 0.156601f
C173 source.n58 a_n1878_n1288# 0.035199f
C174 source.n59 a_n1878_n1288# 0.102135f
C175 source.n60 a_n1878_n1288# 0.032109f
C176 source.n61 a_n1878_n1288# 0.071045f
C177 source.t15 a_n1878_n1288# 0.053316f
C178 source.n62 a_n1878_n1288# 0.055603f
C179 source.n63 a_n1878_n1288# 0.017924f
C180 source.n64 a_n1878_n1288# 0.011821f
C181 source.n65 a_n1878_n1288# 0.156601f
C182 source.n66 a_n1878_n1288# 0.035199f
C183 source.n67 a_n1878_n1288# 0.102135f
C184 source.t17 a_n1878_n1288# 0.034769f
C185 source.t13 a_n1878_n1288# 0.034769f
C186 source.n68 a_n1878_n1288# 0.185871f
C187 source.n69 a_n1878_n1288# 0.272474f
C188 source.t18 a_n1878_n1288# 0.034769f
C189 source.t16 a_n1878_n1288# 0.034769f
C190 source.n70 a_n1878_n1288# 0.185871f
C191 source.n71 a_n1878_n1288# 0.272474f
C192 source.n72 a_n1878_n1288# 0.032109f
C193 source.n73 a_n1878_n1288# 0.071045f
C194 source.t10 a_n1878_n1288# 0.053316f
C195 source.n74 a_n1878_n1288# 0.055603f
C196 source.n75 a_n1878_n1288# 0.017924f
C197 source.n76 a_n1878_n1288# 0.011821f
C198 source.n77 a_n1878_n1288# 0.156601f
C199 source.n78 a_n1878_n1288# 0.035199f
C200 source.n79 a_n1878_n1288# 0.236032f
C201 source.n80 a_n1878_n1288# 0.549163f
C202 minus.n0 a_n1878_n1288# 0.025171f
C203 minus.t9 a_n1878_n1288# 0.077949f
C204 minus.n1 a_n1878_n1288# 0.05871f
C205 minus.t3 a_n1878_n1288# 0.077949f
C206 minus.n2 a_n1878_n1288# 0.102514f
C207 minus.t7 a_n1878_n1288# 0.085379f
C208 minus.n3 a_n1878_n1288# 0.049336f
C209 minus.t2 a_n1878_n1288# 0.077949f
C210 minus.n4 a_n1878_n1288# 0.061744f
C211 minus.t4 a_n1878_n1288# 0.077949f
C212 minus.n5 a_n1878_n1288# 0.05871f
C213 minus.n6 a_n1878_n1288# 0.005712f
C214 minus.n7 a_n1878_n1288# 0.025171f
C215 minus.n8 a_n1878_n1288# 0.025171f
C216 minus.n9 a_n1878_n1288# 0.025171f
C217 minus.n10 a_n1878_n1288# 0.056227f
C218 minus.n11 a_n1878_n1288# 0.005712f
C219 minus.t6 a_n1878_n1288# 0.077949f
C220 minus.n12 a_n1878_n1288# 0.056072f
C221 minus.n13 a_n1878_n1288# 0.60696f
C222 minus.n14 a_n1878_n1288# 0.025171f
C223 minus.t11 a_n1878_n1288# 0.077949f
C224 minus.n15 a_n1878_n1288# 0.05871f
C225 minus.n16 a_n1878_n1288# 0.102514f
C226 minus.t10 a_n1878_n1288# 0.085379f
C227 minus.n17 a_n1878_n1288# 0.049336f
C228 minus.t0 a_n1878_n1288# 0.077949f
C229 minus.n18 a_n1878_n1288# 0.061744f
C230 minus.t8 a_n1878_n1288# 0.077949f
C231 minus.n19 a_n1878_n1288# 0.05871f
C232 minus.n20 a_n1878_n1288# 0.005712f
C233 minus.n21 a_n1878_n1288# 0.025171f
C234 minus.n22 a_n1878_n1288# 0.025171f
C235 minus.n23 a_n1878_n1288# 0.025171f
C236 minus.t5 a_n1878_n1288# 0.077949f
C237 minus.n24 a_n1878_n1288# 0.056227f
C238 minus.n25 a_n1878_n1288# 0.005712f
C239 minus.t1 a_n1878_n1288# 0.077949f
C240 minus.n26 a_n1878_n1288# 0.056072f
C241 minus.n27 a_n1878_n1288# 0.166388f
C242 minus.n28 a_n1878_n1288# 0.749032f
.ends

