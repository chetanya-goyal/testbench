* NGSPICE file created from diffpair465.ext - technology: sky130A

.subckt diffpair465 minus drain_right drain_left source plus
X0 source.t20 plus.t0 drain_left.t6 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X1 source.t23 minus.t0 drain_right.t11 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X2 source.t19 plus.t1 drain_left.t5 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X3 source.t3 minus.t1 drain_right.t10 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X4 drain_right.t9 minus.t2 source.t2 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X5 source.t18 plus.t2 drain_left.t8 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X6 source.t17 plus.t3 drain_left.t11 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X7 source.t16 plus.t4 drain_left.t9 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X8 drain_right.t8 minus.t3 source.t21 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X9 drain_left.t10 plus.t5 source.t15 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X10 drain_right.t7 minus.t4 source.t22 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X11 drain_left.t7 plus.t6 source.t14 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X12 drain_left.t0 plus.t7 source.t13 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X13 a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X14 drain_right.t6 minus.t5 source.t7 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X15 drain_left.t2 plus.t8 source.t12 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X16 drain_left.t4 plus.t9 source.t11 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X17 a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X18 drain_right.t5 minus.t6 source.t0 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X19 drain_left.t1 plus.t10 source.t10 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X20 source.t1 minus.t7 drain_right.t4 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X21 source.t9 plus.t11 drain_left.t3 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X22 drain_right.t3 minus.t8 source.t6 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X23 source.t4 minus.t9 drain_right.t2 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X24 source.t8 minus.t10 drain_right.t1 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X25 a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X26 source.t5 minus.t11 drain_right.t0 a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X27 a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# a_n2158_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
R0 plus.n5 plus.t3 492.565
R1 plus.n23 plus.t10 492.565
R2 plus.n16 plus.t7 469.262
R3 plus.n14 plus.t2 469.262
R4 plus.n2 plus.t6 469.262
R5 plus.n8 plus.t1 469.262
R6 plus.n4 plus.t8 469.262
R7 plus.n34 plus.t0 469.262
R8 plus.n32 plus.t5 469.262
R9 plus.n20 plus.t4 469.262
R10 plus.n26 plus.t9 469.262
R11 plus.n22 plus.t11 469.262
R12 plus.n7 plus.n6 161.3
R13 plus.n8 plus.n3 161.3
R14 plus.n10 plus.n9 161.3
R15 plus.n11 plus.n2 161.3
R16 plus.n13 plus.n12 161.3
R17 plus.n14 plus.n1 161.3
R18 plus.n15 plus.n0 161.3
R19 plus.n17 plus.n16 161.3
R20 plus.n25 plus.n24 161.3
R21 plus.n26 plus.n21 161.3
R22 plus.n28 plus.n27 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus.n16 plus.n15 32.8641
R31 plus.n34 plus.n33 32.8641
R32 plus plus.n35 31.321
R33 plus.n14 plus.n13 28.4823
R34 plus.n7 plus.n4 28.4823
R35 plus.n32 plus.n31 28.4823
R36 plus.n25 plus.n22 28.4823
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 12.2884
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 drain_left.n6 drain_left.n4 60.4406
R65 drain_left.n3 drain_left.n2 60.3851
R66 drain_left.n3 drain_left.n0 60.3851
R67 drain_left.n6 drain_left.n5 59.5527
R68 drain_left.n3 drain_left.n1 59.5525
R69 drain_left.n8 drain_left.n7 59.5525
R70 drain_left drain_left.n3 31.8067
R71 drain_left drain_left.n8 6.54115
R72 drain_left.n1 drain_left.t9 1.6505
R73 drain_left.n1 drain_left.t4 1.6505
R74 drain_left.n2 drain_left.t3 1.6505
R75 drain_left.n2 drain_left.t1 1.6505
R76 drain_left.n0 drain_left.t6 1.6505
R77 drain_left.n0 drain_left.t10 1.6505
R78 drain_left.n7 drain_left.t8 1.6505
R79 drain_left.n7 drain_left.t0 1.6505
R80 drain_left.n5 drain_left.t5 1.6505
R81 drain_left.n5 drain_left.t7 1.6505
R82 drain_left.n4 drain_left.t11 1.6505
R83 drain_left.n4 drain_left.t2 1.6505
R84 drain_left.n8 drain_left.n6 0.888431
R85 source.n538 source.n478 289.615
R86 source.n468 source.n408 289.615
R87 source.n402 source.n342 289.615
R88 source.n332 source.n272 289.615
R89 source.n60 source.n0 289.615
R90 source.n130 source.n70 289.615
R91 source.n196 source.n136 289.615
R92 source.n266 source.n206 289.615
R93 source.n498 source.n497 185
R94 source.n503 source.n502 185
R95 source.n505 source.n504 185
R96 source.n494 source.n493 185
R97 source.n511 source.n510 185
R98 source.n513 source.n512 185
R99 source.n490 source.n489 185
R100 source.n520 source.n519 185
R101 source.n521 source.n488 185
R102 source.n523 source.n522 185
R103 source.n486 source.n485 185
R104 source.n529 source.n528 185
R105 source.n531 source.n530 185
R106 source.n482 source.n481 185
R107 source.n537 source.n536 185
R108 source.n539 source.n538 185
R109 source.n428 source.n427 185
R110 source.n433 source.n432 185
R111 source.n435 source.n434 185
R112 source.n424 source.n423 185
R113 source.n441 source.n440 185
R114 source.n443 source.n442 185
R115 source.n420 source.n419 185
R116 source.n450 source.n449 185
R117 source.n451 source.n418 185
R118 source.n453 source.n452 185
R119 source.n416 source.n415 185
R120 source.n459 source.n458 185
R121 source.n461 source.n460 185
R122 source.n412 source.n411 185
R123 source.n467 source.n466 185
R124 source.n469 source.n468 185
R125 source.n362 source.n361 185
R126 source.n367 source.n366 185
R127 source.n369 source.n368 185
R128 source.n358 source.n357 185
R129 source.n375 source.n374 185
R130 source.n377 source.n376 185
R131 source.n354 source.n353 185
R132 source.n384 source.n383 185
R133 source.n385 source.n352 185
R134 source.n387 source.n386 185
R135 source.n350 source.n349 185
R136 source.n393 source.n392 185
R137 source.n395 source.n394 185
R138 source.n346 source.n345 185
R139 source.n401 source.n400 185
R140 source.n403 source.n402 185
R141 source.n292 source.n291 185
R142 source.n297 source.n296 185
R143 source.n299 source.n298 185
R144 source.n288 source.n287 185
R145 source.n305 source.n304 185
R146 source.n307 source.n306 185
R147 source.n284 source.n283 185
R148 source.n314 source.n313 185
R149 source.n315 source.n282 185
R150 source.n317 source.n316 185
R151 source.n280 source.n279 185
R152 source.n323 source.n322 185
R153 source.n325 source.n324 185
R154 source.n276 source.n275 185
R155 source.n331 source.n330 185
R156 source.n333 source.n332 185
R157 source.n61 source.n60 185
R158 source.n59 source.n58 185
R159 source.n4 source.n3 185
R160 source.n53 source.n52 185
R161 source.n51 source.n50 185
R162 source.n8 source.n7 185
R163 source.n45 source.n44 185
R164 source.n43 source.n10 185
R165 source.n42 source.n41 185
R166 source.n13 source.n11 185
R167 source.n36 source.n35 185
R168 source.n34 source.n33 185
R169 source.n17 source.n16 185
R170 source.n28 source.n27 185
R171 source.n26 source.n25 185
R172 source.n21 source.n20 185
R173 source.n131 source.n130 185
R174 source.n129 source.n128 185
R175 source.n74 source.n73 185
R176 source.n123 source.n122 185
R177 source.n121 source.n120 185
R178 source.n78 source.n77 185
R179 source.n115 source.n114 185
R180 source.n113 source.n80 185
R181 source.n112 source.n111 185
R182 source.n83 source.n81 185
R183 source.n106 source.n105 185
R184 source.n104 source.n103 185
R185 source.n87 source.n86 185
R186 source.n98 source.n97 185
R187 source.n96 source.n95 185
R188 source.n91 source.n90 185
R189 source.n197 source.n196 185
R190 source.n195 source.n194 185
R191 source.n140 source.n139 185
R192 source.n189 source.n188 185
R193 source.n187 source.n186 185
R194 source.n144 source.n143 185
R195 source.n181 source.n180 185
R196 source.n179 source.n146 185
R197 source.n178 source.n177 185
R198 source.n149 source.n147 185
R199 source.n172 source.n171 185
R200 source.n170 source.n169 185
R201 source.n153 source.n152 185
R202 source.n164 source.n163 185
R203 source.n162 source.n161 185
R204 source.n157 source.n156 185
R205 source.n267 source.n266 185
R206 source.n265 source.n264 185
R207 source.n210 source.n209 185
R208 source.n259 source.n258 185
R209 source.n257 source.n256 185
R210 source.n214 source.n213 185
R211 source.n251 source.n250 185
R212 source.n249 source.n216 185
R213 source.n248 source.n247 185
R214 source.n219 source.n217 185
R215 source.n242 source.n241 185
R216 source.n240 source.n239 185
R217 source.n223 source.n222 185
R218 source.n234 source.n233 185
R219 source.n232 source.n231 185
R220 source.n227 source.n226 185
R221 source.n499 source.t0 149.524
R222 source.n429 source.t23 149.524
R223 source.n363 source.t10 149.524
R224 source.n293 source.t20 149.524
R225 source.n22 source.t13 149.524
R226 source.n92 source.t17 149.524
R227 source.n158 source.t7 149.524
R228 source.n228 source.t8 149.524
R229 source.n503 source.n497 104.615
R230 source.n504 source.n503 104.615
R231 source.n504 source.n493 104.615
R232 source.n511 source.n493 104.615
R233 source.n512 source.n511 104.615
R234 source.n512 source.n489 104.615
R235 source.n520 source.n489 104.615
R236 source.n521 source.n520 104.615
R237 source.n522 source.n521 104.615
R238 source.n522 source.n485 104.615
R239 source.n529 source.n485 104.615
R240 source.n530 source.n529 104.615
R241 source.n530 source.n481 104.615
R242 source.n537 source.n481 104.615
R243 source.n538 source.n537 104.615
R244 source.n433 source.n427 104.615
R245 source.n434 source.n433 104.615
R246 source.n434 source.n423 104.615
R247 source.n441 source.n423 104.615
R248 source.n442 source.n441 104.615
R249 source.n442 source.n419 104.615
R250 source.n450 source.n419 104.615
R251 source.n451 source.n450 104.615
R252 source.n452 source.n451 104.615
R253 source.n452 source.n415 104.615
R254 source.n459 source.n415 104.615
R255 source.n460 source.n459 104.615
R256 source.n460 source.n411 104.615
R257 source.n467 source.n411 104.615
R258 source.n468 source.n467 104.615
R259 source.n367 source.n361 104.615
R260 source.n368 source.n367 104.615
R261 source.n368 source.n357 104.615
R262 source.n375 source.n357 104.615
R263 source.n376 source.n375 104.615
R264 source.n376 source.n353 104.615
R265 source.n384 source.n353 104.615
R266 source.n385 source.n384 104.615
R267 source.n386 source.n385 104.615
R268 source.n386 source.n349 104.615
R269 source.n393 source.n349 104.615
R270 source.n394 source.n393 104.615
R271 source.n394 source.n345 104.615
R272 source.n401 source.n345 104.615
R273 source.n402 source.n401 104.615
R274 source.n297 source.n291 104.615
R275 source.n298 source.n297 104.615
R276 source.n298 source.n287 104.615
R277 source.n305 source.n287 104.615
R278 source.n306 source.n305 104.615
R279 source.n306 source.n283 104.615
R280 source.n314 source.n283 104.615
R281 source.n315 source.n314 104.615
R282 source.n316 source.n315 104.615
R283 source.n316 source.n279 104.615
R284 source.n323 source.n279 104.615
R285 source.n324 source.n323 104.615
R286 source.n324 source.n275 104.615
R287 source.n331 source.n275 104.615
R288 source.n332 source.n331 104.615
R289 source.n60 source.n59 104.615
R290 source.n59 source.n3 104.615
R291 source.n52 source.n3 104.615
R292 source.n52 source.n51 104.615
R293 source.n51 source.n7 104.615
R294 source.n44 source.n7 104.615
R295 source.n44 source.n43 104.615
R296 source.n43 source.n42 104.615
R297 source.n42 source.n11 104.615
R298 source.n35 source.n11 104.615
R299 source.n35 source.n34 104.615
R300 source.n34 source.n16 104.615
R301 source.n27 source.n16 104.615
R302 source.n27 source.n26 104.615
R303 source.n26 source.n20 104.615
R304 source.n130 source.n129 104.615
R305 source.n129 source.n73 104.615
R306 source.n122 source.n73 104.615
R307 source.n122 source.n121 104.615
R308 source.n121 source.n77 104.615
R309 source.n114 source.n77 104.615
R310 source.n114 source.n113 104.615
R311 source.n113 source.n112 104.615
R312 source.n112 source.n81 104.615
R313 source.n105 source.n81 104.615
R314 source.n105 source.n104 104.615
R315 source.n104 source.n86 104.615
R316 source.n97 source.n86 104.615
R317 source.n97 source.n96 104.615
R318 source.n96 source.n90 104.615
R319 source.n196 source.n195 104.615
R320 source.n195 source.n139 104.615
R321 source.n188 source.n139 104.615
R322 source.n188 source.n187 104.615
R323 source.n187 source.n143 104.615
R324 source.n180 source.n143 104.615
R325 source.n180 source.n179 104.615
R326 source.n179 source.n178 104.615
R327 source.n178 source.n147 104.615
R328 source.n171 source.n147 104.615
R329 source.n171 source.n170 104.615
R330 source.n170 source.n152 104.615
R331 source.n163 source.n152 104.615
R332 source.n163 source.n162 104.615
R333 source.n162 source.n156 104.615
R334 source.n266 source.n265 104.615
R335 source.n265 source.n209 104.615
R336 source.n258 source.n209 104.615
R337 source.n258 source.n257 104.615
R338 source.n257 source.n213 104.615
R339 source.n250 source.n213 104.615
R340 source.n250 source.n249 104.615
R341 source.n249 source.n248 104.615
R342 source.n248 source.n217 104.615
R343 source.n241 source.n217 104.615
R344 source.n241 source.n240 104.615
R345 source.n240 source.n222 104.615
R346 source.n233 source.n222 104.615
R347 source.n233 source.n232 104.615
R348 source.n232 source.n226 104.615
R349 source.t0 source.n497 52.3082
R350 source.t23 source.n427 52.3082
R351 source.t10 source.n361 52.3082
R352 source.t20 source.n291 52.3082
R353 source.t13 source.n20 52.3082
R354 source.t17 source.n90 52.3082
R355 source.t7 source.n156 52.3082
R356 source.t8 source.n226 52.3082
R357 source.n67 source.n66 42.8739
R358 source.n69 source.n68 42.8739
R359 source.n203 source.n202 42.8739
R360 source.n205 source.n204 42.8739
R361 source.n477 source.n476 42.8737
R362 source.n475 source.n474 42.8737
R363 source.n341 source.n340 42.8737
R364 source.n339 source.n338 42.8737
R365 source.n543 source.n542 29.8581
R366 source.n473 source.n472 29.8581
R367 source.n407 source.n406 29.8581
R368 source.n337 source.n336 29.8581
R369 source.n65 source.n64 29.8581
R370 source.n135 source.n134 29.8581
R371 source.n201 source.n200 29.8581
R372 source.n271 source.n270 29.8581
R373 source.n337 source.n271 22.1757
R374 source.n544 source.n65 16.4688
R375 source.n523 source.n488 13.1884
R376 source.n453 source.n418 13.1884
R377 source.n387 source.n352 13.1884
R378 source.n317 source.n282 13.1884
R379 source.n45 source.n10 13.1884
R380 source.n115 source.n80 13.1884
R381 source.n181 source.n146 13.1884
R382 source.n251 source.n216 13.1884
R383 source.n519 source.n518 12.8005
R384 source.n524 source.n486 12.8005
R385 source.n449 source.n448 12.8005
R386 source.n454 source.n416 12.8005
R387 source.n383 source.n382 12.8005
R388 source.n388 source.n350 12.8005
R389 source.n313 source.n312 12.8005
R390 source.n318 source.n280 12.8005
R391 source.n46 source.n8 12.8005
R392 source.n41 source.n12 12.8005
R393 source.n116 source.n78 12.8005
R394 source.n111 source.n82 12.8005
R395 source.n182 source.n144 12.8005
R396 source.n177 source.n148 12.8005
R397 source.n252 source.n214 12.8005
R398 source.n247 source.n218 12.8005
R399 source.n517 source.n490 12.0247
R400 source.n528 source.n527 12.0247
R401 source.n447 source.n420 12.0247
R402 source.n458 source.n457 12.0247
R403 source.n381 source.n354 12.0247
R404 source.n392 source.n391 12.0247
R405 source.n311 source.n284 12.0247
R406 source.n322 source.n321 12.0247
R407 source.n50 source.n49 12.0247
R408 source.n40 source.n13 12.0247
R409 source.n120 source.n119 12.0247
R410 source.n110 source.n83 12.0247
R411 source.n186 source.n185 12.0247
R412 source.n176 source.n149 12.0247
R413 source.n256 source.n255 12.0247
R414 source.n246 source.n219 12.0247
R415 source.n514 source.n513 11.249
R416 source.n531 source.n484 11.249
R417 source.n444 source.n443 11.249
R418 source.n461 source.n414 11.249
R419 source.n378 source.n377 11.249
R420 source.n395 source.n348 11.249
R421 source.n308 source.n307 11.249
R422 source.n325 source.n278 11.249
R423 source.n53 source.n6 11.249
R424 source.n37 source.n36 11.249
R425 source.n123 source.n76 11.249
R426 source.n107 source.n106 11.249
R427 source.n189 source.n142 11.249
R428 source.n173 source.n172 11.249
R429 source.n259 source.n212 11.249
R430 source.n243 source.n242 11.249
R431 source.n510 source.n492 10.4732
R432 source.n532 source.n482 10.4732
R433 source.n440 source.n422 10.4732
R434 source.n462 source.n412 10.4732
R435 source.n374 source.n356 10.4732
R436 source.n396 source.n346 10.4732
R437 source.n304 source.n286 10.4732
R438 source.n326 source.n276 10.4732
R439 source.n54 source.n4 10.4732
R440 source.n33 source.n15 10.4732
R441 source.n124 source.n74 10.4732
R442 source.n103 source.n85 10.4732
R443 source.n190 source.n140 10.4732
R444 source.n169 source.n151 10.4732
R445 source.n260 source.n210 10.4732
R446 source.n239 source.n221 10.4732
R447 source.n499 source.n498 10.2747
R448 source.n429 source.n428 10.2747
R449 source.n363 source.n362 10.2747
R450 source.n293 source.n292 10.2747
R451 source.n22 source.n21 10.2747
R452 source.n92 source.n91 10.2747
R453 source.n158 source.n157 10.2747
R454 source.n228 source.n227 10.2747
R455 source.n509 source.n494 9.69747
R456 source.n536 source.n535 9.69747
R457 source.n439 source.n424 9.69747
R458 source.n466 source.n465 9.69747
R459 source.n373 source.n358 9.69747
R460 source.n400 source.n399 9.69747
R461 source.n303 source.n288 9.69747
R462 source.n330 source.n329 9.69747
R463 source.n58 source.n57 9.69747
R464 source.n32 source.n17 9.69747
R465 source.n128 source.n127 9.69747
R466 source.n102 source.n87 9.69747
R467 source.n194 source.n193 9.69747
R468 source.n168 source.n153 9.69747
R469 source.n264 source.n263 9.69747
R470 source.n238 source.n223 9.69747
R471 source.n542 source.n541 9.45567
R472 source.n472 source.n471 9.45567
R473 source.n406 source.n405 9.45567
R474 source.n336 source.n335 9.45567
R475 source.n64 source.n63 9.45567
R476 source.n134 source.n133 9.45567
R477 source.n200 source.n199 9.45567
R478 source.n270 source.n269 9.45567
R479 source.n541 source.n540 9.3005
R480 source.n480 source.n479 9.3005
R481 source.n535 source.n534 9.3005
R482 source.n533 source.n532 9.3005
R483 source.n484 source.n483 9.3005
R484 source.n527 source.n526 9.3005
R485 source.n525 source.n524 9.3005
R486 source.n501 source.n500 9.3005
R487 source.n496 source.n495 9.3005
R488 source.n507 source.n506 9.3005
R489 source.n509 source.n508 9.3005
R490 source.n492 source.n491 9.3005
R491 source.n515 source.n514 9.3005
R492 source.n517 source.n516 9.3005
R493 source.n518 source.n487 9.3005
R494 source.n471 source.n470 9.3005
R495 source.n410 source.n409 9.3005
R496 source.n465 source.n464 9.3005
R497 source.n463 source.n462 9.3005
R498 source.n414 source.n413 9.3005
R499 source.n457 source.n456 9.3005
R500 source.n455 source.n454 9.3005
R501 source.n431 source.n430 9.3005
R502 source.n426 source.n425 9.3005
R503 source.n437 source.n436 9.3005
R504 source.n439 source.n438 9.3005
R505 source.n422 source.n421 9.3005
R506 source.n445 source.n444 9.3005
R507 source.n447 source.n446 9.3005
R508 source.n448 source.n417 9.3005
R509 source.n405 source.n404 9.3005
R510 source.n344 source.n343 9.3005
R511 source.n399 source.n398 9.3005
R512 source.n397 source.n396 9.3005
R513 source.n348 source.n347 9.3005
R514 source.n391 source.n390 9.3005
R515 source.n389 source.n388 9.3005
R516 source.n365 source.n364 9.3005
R517 source.n360 source.n359 9.3005
R518 source.n371 source.n370 9.3005
R519 source.n373 source.n372 9.3005
R520 source.n356 source.n355 9.3005
R521 source.n379 source.n378 9.3005
R522 source.n381 source.n380 9.3005
R523 source.n382 source.n351 9.3005
R524 source.n335 source.n334 9.3005
R525 source.n274 source.n273 9.3005
R526 source.n329 source.n328 9.3005
R527 source.n327 source.n326 9.3005
R528 source.n278 source.n277 9.3005
R529 source.n321 source.n320 9.3005
R530 source.n319 source.n318 9.3005
R531 source.n295 source.n294 9.3005
R532 source.n290 source.n289 9.3005
R533 source.n301 source.n300 9.3005
R534 source.n303 source.n302 9.3005
R535 source.n286 source.n285 9.3005
R536 source.n309 source.n308 9.3005
R537 source.n311 source.n310 9.3005
R538 source.n312 source.n281 9.3005
R539 source.n24 source.n23 9.3005
R540 source.n19 source.n18 9.3005
R541 source.n30 source.n29 9.3005
R542 source.n32 source.n31 9.3005
R543 source.n15 source.n14 9.3005
R544 source.n38 source.n37 9.3005
R545 source.n40 source.n39 9.3005
R546 source.n12 source.n9 9.3005
R547 source.n63 source.n62 9.3005
R548 source.n2 source.n1 9.3005
R549 source.n57 source.n56 9.3005
R550 source.n55 source.n54 9.3005
R551 source.n6 source.n5 9.3005
R552 source.n49 source.n48 9.3005
R553 source.n47 source.n46 9.3005
R554 source.n94 source.n93 9.3005
R555 source.n89 source.n88 9.3005
R556 source.n100 source.n99 9.3005
R557 source.n102 source.n101 9.3005
R558 source.n85 source.n84 9.3005
R559 source.n108 source.n107 9.3005
R560 source.n110 source.n109 9.3005
R561 source.n82 source.n79 9.3005
R562 source.n133 source.n132 9.3005
R563 source.n72 source.n71 9.3005
R564 source.n127 source.n126 9.3005
R565 source.n125 source.n124 9.3005
R566 source.n76 source.n75 9.3005
R567 source.n119 source.n118 9.3005
R568 source.n117 source.n116 9.3005
R569 source.n160 source.n159 9.3005
R570 source.n155 source.n154 9.3005
R571 source.n166 source.n165 9.3005
R572 source.n168 source.n167 9.3005
R573 source.n151 source.n150 9.3005
R574 source.n174 source.n173 9.3005
R575 source.n176 source.n175 9.3005
R576 source.n148 source.n145 9.3005
R577 source.n199 source.n198 9.3005
R578 source.n138 source.n137 9.3005
R579 source.n193 source.n192 9.3005
R580 source.n191 source.n190 9.3005
R581 source.n142 source.n141 9.3005
R582 source.n185 source.n184 9.3005
R583 source.n183 source.n182 9.3005
R584 source.n230 source.n229 9.3005
R585 source.n225 source.n224 9.3005
R586 source.n236 source.n235 9.3005
R587 source.n238 source.n237 9.3005
R588 source.n221 source.n220 9.3005
R589 source.n244 source.n243 9.3005
R590 source.n246 source.n245 9.3005
R591 source.n218 source.n215 9.3005
R592 source.n269 source.n268 9.3005
R593 source.n208 source.n207 9.3005
R594 source.n263 source.n262 9.3005
R595 source.n261 source.n260 9.3005
R596 source.n212 source.n211 9.3005
R597 source.n255 source.n254 9.3005
R598 source.n253 source.n252 9.3005
R599 source.n506 source.n505 8.92171
R600 source.n539 source.n480 8.92171
R601 source.n436 source.n435 8.92171
R602 source.n469 source.n410 8.92171
R603 source.n370 source.n369 8.92171
R604 source.n403 source.n344 8.92171
R605 source.n300 source.n299 8.92171
R606 source.n333 source.n274 8.92171
R607 source.n61 source.n2 8.92171
R608 source.n29 source.n28 8.92171
R609 source.n131 source.n72 8.92171
R610 source.n99 source.n98 8.92171
R611 source.n197 source.n138 8.92171
R612 source.n165 source.n164 8.92171
R613 source.n267 source.n208 8.92171
R614 source.n235 source.n234 8.92171
R615 source.n502 source.n496 8.14595
R616 source.n540 source.n478 8.14595
R617 source.n432 source.n426 8.14595
R618 source.n470 source.n408 8.14595
R619 source.n366 source.n360 8.14595
R620 source.n404 source.n342 8.14595
R621 source.n296 source.n290 8.14595
R622 source.n334 source.n272 8.14595
R623 source.n62 source.n0 8.14595
R624 source.n25 source.n19 8.14595
R625 source.n132 source.n70 8.14595
R626 source.n95 source.n89 8.14595
R627 source.n198 source.n136 8.14595
R628 source.n161 source.n155 8.14595
R629 source.n268 source.n206 8.14595
R630 source.n231 source.n225 8.14595
R631 source.n501 source.n498 7.3702
R632 source.n431 source.n428 7.3702
R633 source.n365 source.n362 7.3702
R634 source.n295 source.n292 7.3702
R635 source.n24 source.n21 7.3702
R636 source.n94 source.n91 7.3702
R637 source.n160 source.n157 7.3702
R638 source.n230 source.n227 7.3702
R639 source.n502 source.n501 5.81868
R640 source.n542 source.n478 5.81868
R641 source.n432 source.n431 5.81868
R642 source.n472 source.n408 5.81868
R643 source.n366 source.n365 5.81868
R644 source.n406 source.n342 5.81868
R645 source.n296 source.n295 5.81868
R646 source.n336 source.n272 5.81868
R647 source.n64 source.n0 5.81868
R648 source.n25 source.n24 5.81868
R649 source.n134 source.n70 5.81868
R650 source.n95 source.n94 5.81868
R651 source.n200 source.n136 5.81868
R652 source.n161 source.n160 5.81868
R653 source.n270 source.n206 5.81868
R654 source.n231 source.n230 5.81868
R655 source.n544 source.n543 5.7074
R656 source.n505 source.n496 5.04292
R657 source.n540 source.n539 5.04292
R658 source.n435 source.n426 5.04292
R659 source.n470 source.n469 5.04292
R660 source.n369 source.n360 5.04292
R661 source.n404 source.n403 5.04292
R662 source.n299 source.n290 5.04292
R663 source.n334 source.n333 5.04292
R664 source.n62 source.n61 5.04292
R665 source.n28 source.n19 5.04292
R666 source.n132 source.n131 5.04292
R667 source.n98 source.n89 5.04292
R668 source.n198 source.n197 5.04292
R669 source.n164 source.n155 5.04292
R670 source.n268 source.n267 5.04292
R671 source.n234 source.n225 5.04292
R672 source.n506 source.n494 4.26717
R673 source.n536 source.n480 4.26717
R674 source.n436 source.n424 4.26717
R675 source.n466 source.n410 4.26717
R676 source.n370 source.n358 4.26717
R677 source.n400 source.n344 4.26717
R678 source.n300 source.n288 4.26717
R679 source.n330 source.n274 4.26717
R680 source.n58 source.n2 4.26717
R681 source.n29 source.n17 4.26717
R682 source.n128 source.n72 4.26717
R683 source.n99 source.n87 4.26717
R684 source.n194 source.n138 4.26717
R685 source.n165 source.n153 4.26717
R686 source.n264 source.n208 4.26717
R687 source.n235 source.n223 4.26717
R688 source.n510 source.n509 3.49141
R689 source.n535 source.n482 3.49141
R690 source.n440 source.n439 3.49141
R691 source.n465 source.n412 3.49141
R692 source.n374 source.n373 3.49141
R693 source.n399 source.n346 3.49141
R694 source.n304 source.n303 3.49141
R695 source.n329 source.n276 3.49141
R696 source.n57 source.n4 3.49141
R697 source.n33 source.n32 3.49141
R698 source.n127 source.n74 3.49141
R699 source.n103 source.n102 3.49141
R700 source.n193 source.n140 3.49141
R701 source.n169 source.n168 3.49141
R702 source.n263 source.n210 3.49141
R703 source.n239 source.n238 3.49141
R704 source.n500 source.n499 2.84303
R705 source.n430 source.n429 2.84303
R706 source.n364 source.n363 2.84303
R707 source.n294 source.n293 2.84303
R708 source.n23 source.n22 2.84303
R709 source.n93 source.n92 2.84303
R710 source.n159 source.n158 2.84303
R711 source.n229 source.n228 2.84303
R712 source.n513 source.n492 2.71565
R713 source.n532 source.n531 2.71565
R714 source.n443 source.n422 2.71565
R715 source.n462 source.n461 2.71565
R716 source.n377 source.n356 2.71565
R717 source.n396 source.n395 2.71565
R718 source.n307 source.n286 2.71565
R719 source.n326 source.n325 2.71565
R720 source.n54 source.n53 2.71565
R721 source.n36 source.n15 2.71565
R722 source.n124 source.n123 2.71565
R723 source.n106 source.n85 2.71565
R724 source.n190 source.n189 2.71565
R725 source.n172 source.n151 2.71565
R726 source.n260 source.n259 2.71565
R727 source.n242 source.n221 2.71565
R728 source.n514 source.n490 1.93989
R729 source.n528 source.n484 1.93989
R730 source.n444 source.n420 1.93989
R731 source.n458 source.n414 1.93989
R732 source.n378 source.n354 1.93989
R733 source.n392 source.n348 1.93989
R734 source.n308 source.n284 1.93989
R735 source.n322 source.n278 1.93989
R736 source.n50 source.n6 1.93989
R737 source.n37 source.n13 1.93989
R738 source.n120 source.n76 1.93989
R739 source.n107 source.n83 1.93989
R740 source.n186 source.n142 1.93989
R741 source.n173 source.n149 1.93989
R742 source.n256 source.n212 1.93989
R743 source.n243 source.n219 1.93989
R744 source.n476 source.t6 1.6505
R745 source.n476 source.t5 1.6505
R746 source.n474 source.t2 1.6505
R747 source.n474 source.t1 1.6505
R748 source.n340 source.t11 1.6505
R749 source.n340 source.t9 1.6505
R750 source.n338 source.t15 1.6505
R751 source.n338 source.t16 1.6505
R752 source.n66 source.t14 1.6505
R753 source.n66 source.t18 1.6505
R754 source.n68 source.t12 1.6505
R755 source.n68 source.t19 1.6505
R756 source.n202 source.t22 1.6505
R757 source.n202 source.t3 1.6505
R758 source.n204 source.t21 1.6505
R759 source.n204 source.t4 1.6505
R760 source.n519 source.n517 1.16414
R761 source.n527 source.n486 1.16414
R762 source.n449 source.n447 1.16414
R763 source.n457 source.n416 1.16414
R764 source.n383 source.n381 1.16414
R765 source.n391 source.n350 1.16414
R766 source.n313 source.n311 1.16414
R767 source.n321 source.n280 1.16414
R768 source.n49 source.n8 1.16414
R769 source.n41 source.n40 1.16414
R770 source.n119 source.n78 1.16414
R771 source.n111 source.n110 1.16414
R772 source.n185 source.n144 1.16414
R773 source.n177 source.n176 1.16414
R774 source.n255 source.n214 1.16414
R775 source.n247 source.n246 1.16414
R776 source.n271 source.n205 0.888431
R777 source.n205 source.n203 0.888431
R778 source.n203 source.n201 0.888431
R779 source.n135 source.n69 0.888431
R780 source.n69 source.n67 0.888431
R781 source.n67 source.n65 0.888431
R782 source.n339 source.n337 0.888431
R783 source.n341 source.n339 0.888431
R784 source.n407 source.n341 0.888431
R785 source.n475 source.n473 0.888431
R786 source.n477 source.n475 0.888431
R787 source.n543 source.n477 0.888431
R788 source.n201 source.n135 0.470328
R789 source.n473 source.n407 0.470328
R790 source.n518 source.n488 0.388379
R791 source.n524 source.n523 0.388379
R792 source.n448 source.n418 0.388379
R793 source.n454 source.n453 0.388379
R794 source.n382 source.n352 0.388379
R795 source.n388 source.n387 0.388379
R796 source.n312 source.n282 0.388379
R797 source.n318 source.n317 0.388379
R798 source.n46 source.n45 0.388379
R799 source.n12 source.n10 0.388379
R800 source.n116 source.n115 0.388379
R801 source.n82 source.n80 0.388379
R802 source.n182 source.n181 0.388379
R803 source.n148 source.n146 0.388379
R804 source.n252 source.n251 0.388379
R805 source.n218 source.n216 0.388379
R806 source source.n544 0.188
R807 source.n500 source.n495 0.155672
R808 source.n507 source.n495 0.155672
R809 source.n508 source.n507 0.155672
R810 source.n508 source.n491 0.155672
R811 source.n515 source.n491 0.155672
R812 source.n516 source.n515 0.155672
R813 source.n516 source.n487 0.155672
R814 source.n525 source.n487 0.155672
R815 source.n526 source.n525 0.155672
R816 source.n526 source.n483 0.155672
R817 source.n533 source.n483 0.155672
R818 source.n534 source.n533 0.155672
R819 source.n534 source.n479 0.155672
R820 source.n541 source.n479 0.155672
R821 source.n430 source.n425 0.155672
R822 source.n437 source.n425 0.155672
R823 source.n438 source.n437 0.155672
R824 source.n438 source.n421 0.155672
R825 source.n445 source.n421 0.155672
R826 source.n446 source.n445 0.155672
R827 source.n446 source.n417 0.155672
R828 source.n455 source.n417 0.155672
R829 source.n456 source.n455 0.155672
R830 source.n456 source.n413 0.155672
R831 source.n463 source.n413 0.155672
R832 source.n464 source.n463 0.155672
R833 source.n464 source.n409 0.155672
R834 source.n471 source.n409 0.155672
R835 source.n364 source.n359 0.155672
R836 source.n371 source.n359 0.155672
R837 source.n372 source.n371 0.155672
R838 source.n372 source.n355 0.155672
R839 source.n379 source.n355 0.155672
R840 source.n380 source.n379 0.155672
R841 source.n380 source.n351 0.155672
R842 source.n389 source.n351 0.155672
R843 source.n390 source.n389 0.155672
R844 source.n390 source.n347 0.155672
R845 source.n397 source.n347 0.155672
R846 source.n398 source.n397 0.155672
R847 source.n398 source.n343 0.155672
R848 source.n405 source.n343 0.155672
R849 source.n294 source.n289 0.155672
R850 source.n301 source.n289 0.155672
R851 source.n302 source.n301 0.155672
R852 source.n302 source.n285 0.155672
R853 source.n309 source.n285 0.155672
R854 source.n310 source.n309 0.155672
R855 source.n310 source.n281 0.155672
R856 source.n319 source.n281 0.155672
R857 source.n320 source.n319 0.155672
R858 source.n320 source.n277 0.155672
R859 source.n327 source.n277 0.155672
R860 source.n328 source.n327 0.155672
R861 source.n328 source.n273 0.155672
R862 source.n335 source.n273 0.155672
R863 source.n63 source.n1 0.155672
R864 source.n56 source.n1 0.155672
R865 source.n56 source.n55 0.155672
R866 source.n55 source.n5 0.155672
R867 source.n48 source.n5 0.155672
R868 source.n48 source.n47 0.155672
R869 source.n47 source.n9 0.155672
R870 source.n39 source.n9 0.155672
R871 source.n39 source.n38 0.155672
R872 source.n38 source.n14 0.155672
R873 source.n31 source.n14 0.155672
R874 source.n31 source.n30 0.155672
R875 source.n30 source.n18 0.155672
R876 source.n23 source.n18 0.155672
R877 source.n133 source.n71 0.155672
R878 source.n126 source.n71 0.155672
R879 source.n126 source.n125 0.155672
R880 source.n125 source.n75 0.155672
R881 source.n118 source.n75 0.155672
R882 source.n118 source.n117 0.155672
R883 source.n117 source.n79 0.155672
R884 source.n109 source.n79 0.155672
R885 source.n109 source.n108 0.155672
R886 source.n108 source.n84 0.155672
R887 source.n101 source.n84 0.155672
R888 source.n101 source.n100 0.155672
R889 source.n100 source.n88 0.155672
R890 source.n93 source.n88 0.155672
R891 source.n199 source.n137 0.155672
R892 source.n192 source.n137 0.155672
R893 source.n192 source.n191 0.155672
R894 source.n191 source.n141 0.155672
R895 source.n184 source.n141 0.155672
R896 source.n184 source.n183 0.155672
R897 source.n183 source.n145 0.155672
R898 source.n175 source.n145 0.155672
R899 source.n175 source.n174 0.155672
R900 source.n174 source.n150 0.155672
R901 source.n167 source.n150 0.155672
R902 source.n167 source.n166 0.155672
R903 source.n166 source.n154 0.155672
R904 source.n159 source.n154 0.155672
R905 source.n269 source.n207 0.155672
R906 source.n262 source.n207 0.155672
R907 source.n262 source.n261 0.155672
R908 source.n261 source.n211 0.155672
R909 source.n254 source.n211 0.155672
R910 source.n254 source.n253 0.155672
R911 source.n253 source.n215 0.155672
R912 source.n245 source.n215 0.155672
R913 source.n245 source.n244 0.155672
R914 source.n244 source.n220 0.155672
R915 source.n237 source.n220 0.155672
R916 source.n237 source.n236 0.155672
R917 source.n236 source.n224 0.155672
R918 source.n229 source.n224 0.155672
R919 minus.n5 minus.t5 492.565
R920 minus.n23 minus.t0 492.565
R921 minus.n4 minus.t1 469.262
R922 minus.n8 minus.t4 469.262
R923 minus.n10 minus.t9 469.262
R924 minus.n14 minus.t3 469.262
R925 minus.n16 minus.t10 469.262
R926 minus.n22 minus.t2 469.262
R927 minus.n26 minus.t7 469.262
R928 minus.n28 minus.t8 469.262
R929 minus.n32 minus.t11 469.262
R930 minus.n34 minus.t6 469.262
R931 minus.n17 minus.n16 161.3
R932 minus.n15 minus.n0 161.3
R933 minus.n14 minus.n13 161.3
R934 minus.n12 minus.n1 161.3
R935 minus.n11 minus.n10 161.3
R936 minus.n9 minus.n2 161.3
R937 minus.n8 minus.n7 161.3
R938 minus.n6 minus.n3 161.3
R939 minus.n35 minus.n34 161.3
R940 minus.n33 minus.n18 161.3
R941 minus.n32 minus.n31 161.3
R942 minus.n30 minus.n19 161.3
R943 minus.n29 minus.n28 161.3
R944 minus.n27 minus.n20 161.3
R945 minus.n26 minus.n25 161.3
R946 minus.n24 minus.n21 161.3
R947 minus.n6 minus.n5 44.8907
R948 minus.n24 minus.n23 44.8907
R949 minus.n36 minus.n17 37.4399
R950 minus.n16 minus.n15 32.8641
R951 minus.n34 minus.n33 32.8641
R952 minus.n4 minus.n3 28.4823
R953 minus.n14 minus.n1 28.4823
R954 minus.n22 minus.n21 28.4823
R955 minus.n32 minus.n19 28.4823
R956 minus.n10 minus.n9 24.1005
R957 minus.n9 minus.n8 24.1005
R958 minus.n27 minus.n26 24.1005
R959 minus.n28 minus.n27 24.1005
R960 minus.n8 minus.n3 19.7187
R961 minus.n10 minus.n1 19.7187
R962 minus.n26 minus.n21 19.7187
R963 minus.n28 minus.n19 19.7187
R964 minus.n5 minus.n4 18.4104
R965 minus.n23 minus.n22 18.4104
R966 minus.n15 minus.n14 15.3369
R967 minus.n33 minus.n32 15.3369
R968 minus.n36 minus.n35 6.64444
R969 minus.n17 minus.n0 0.189894
R970 minus.n13 minus.n0 0.189894
R971 minus.n13 minus.n12 0.189894
R972 minus.n12 minus.n11 0.189894
R973 minus.n11 minus.n2 0.189894
R974 minus.n7 minus.n2 0.189894
R975 minus.n7 minus.n6 0.189894
R976 minus.n25 minus.n24 0.189894
R977 minus.n25 minus.n20 0.189894
R978 minus.n29 minus.n20 0.189894
R979 minus.n30 minus.n29 0.189894
R980 minus.n31 minus.n30 0.189894
R981 minus.n31 minus.n18 0.189894
R982 minus.n35 minus.n18 0.189894
R983 minus minus.n36 0.188
R984 drain_right.n6 drain_right.n4 60.4404
R985 drain_right.n3 drain_right.n2 60.3851
R986 drain_right.n3 drain_right.n0 60.3851
R987 drain_right.n6 drain_right.n5 59.5527
R988 drain_right.n8 drain_right.n7 59.5527
R989 drain_right.n3 drain_right.n1 59.5525
R990 drain_right drain_right.n3 31.2535
R991 drain_right drain_right.n8 6.54115
R992 drain_right.n1 drain_right.t4 1.6505
R993 drain_right.n1 drain_right.t3 1.6505
R994 drain_right.n2 drain_right.t0 1.6505
R995 drain_right.n2 drain_right.t5 1.6505
R996 drain_right.n0 drain_right.t11 1.6505
R997 drain_right.n0 drain_right.t9 1.6505
R998 drain_right.n4 drain_right.t10 1.6505
R999 drain_right.n4 drain_right.t6 1.6505
R1000 drain_right.n5 drain_right.t2 1.6505
R1001 drain_right.n5 drain_right.t7 1.6505
R1002 drain_right.n7 drain_right.t1 1.6505
R1003 drain_right.n7 drain_right.t8 1.6505
R1004 drain_right.n8 drain_right.n6 0.888431
C0 plus drain_left 8.09882f
C1 drain_left drain_right 1.08491f
C2 drain_left minus 0.17184f
C3 plus drain_right 0.366822f
C4 plus minus 5.83479f
C5 drain_left source 15.505099f
C6 minus drain_right 7.88707f
C7 plus source 7.79416f
C8 drain_right source 15.5071f
C9 minus source 7.78012f
C10 drain_right a_n2158_n3288# 6.2102f
C11 drain_left a_n2158_n3288# 6.52051f
C12 source a_n2158_n3288# 9.101151f
C13 minus a_n2158_n3288# 8.509627f
C14 plus a_n2158_n3288# 10.214849f
C15 drain_right.t11 a_n2158_n3288# 0.257089f
C16 drain_right.t9 a_n2158_n3288# 0.257089f
C17 drain_right.n0 a_n2158_n3288# 2.29306f
C18 drain_right.t4 a_n2158_n3288# 0.257089f
C19 drain_right.t3 a_n2158_n3288# 0.257089f
C20 drain_right.n1 a_n2158_n3288# 2.28769f
C21 drain_right.t0 a_n2158_n3288# 0.257089f
C22 drain_right.t5 a_n2158_n3288# 0.257089f
C23 drain_right.n2 a_n2158_n3288# 2.29306f
C24 drain_right.n3 a_n2158_n3288# 2.45998f
C25 drain_right.t10 a_n2158_n3288# 0.257089f
C26 drain_right.t6 a_n2158_n3288# 0.257089f
C27 drain_right.n4 a_n2158_n3288# 2.29347f
C28 drain_right.t2 a_n2158_n3288# 0.257089f
C29 drain_right.t7 a_n2158_n3288# 0.257089f
C30 drain_right.n5 a_n2158_n3288# 2.2877f
C31 drain_right.n6 a_n2158_n3288# 0.770464f
C32 drain_right.t1 a_n2158_n3288# 0.257089f
C33 drain_right.t8 a_n2158_n3288# 0.257089f
C34 drain_right.n7 a_n2158_n3288# 2.2877f
C35 drain_right.n8 a_n2158_n3288# 0.622458f
C36 minus.n0 a_n2158_n3288# 0.041782f
C37 minus.n1 a_n2158_n3288# 0.009481f
C38 minus.t3 a_n2158_n3288# 1.0008f
C39 minus.n2 a_n2158_n3288# 0.041782f
C40 minus.n3 a_n2158_n3288# 0.009481f
C41 minus.t4 a_n2158_n3288# 1.0008f
C42 minus.t5 a_n2158_n3288# 1.01968f
C43 minus.t1 a_n2158_n3288# 1.0008f
C44 minus.n4 a_n2158_n3288# 0.40381f
C45 minus.n5 a_n2158_n3288# 0.383996f
C46 minus.n6 a_n2158_n3288# 0.175281f
C47 minus.n7 a_n2158_n3288# 0.041782f
C48 minus.n8 a_n2158_n3288# 0.399137f
C49 minus.n9 a_n2158_n3288# 0.009481f
C50 minus.t9 a_n2158_n3288# 1.0008f
C51 minus.n10 a_n2158_n3288# 0.399137f
C52 minus.n11 a_n2158_n3288# 0.041782f
C53 minus.n12 a_n2158_n3288# 0.041782f
C54 minus.n13 a_n2158_n3288# 0.041782f
C55 minus.n14 a_n2158_n3288# 0.399137f
C56 minus.n15 a_n2158_n3288# 0.009481f
C57 minus.t10 a_n2158_n3288# 1.0008f
C58 minus.n16 a_n2158_n3288# 0.397204f
C59 minus.n17 a_n2158_n3288# 1.56079f
C60 minus.n18 a_n2158_n3288# 0.041782f
C61 minus.n19 a_n2158_n3288# 0.009481f
C62 minus.n20 a_n2158_n3288# 0.041782f
C63 minus.n21 a_n2158_n3288# 0.009481f
C64 minus.t0 a_n2158_n3288# 1.01968f
C65 minus.t2 a_n2158_n3288# 1.0008f
C66 minus.n22 a_n2158_n3288# 0.40381f
C67 minus.n23 a_n2158_n3288# 0.383996f
C68 minus.n24 a_n2158_n3288# 0.175281f
C69 minus.n25 a_n2158_n3288# 0.041782f
C70 minus.t7 a_n2158_n3288# 1.0008f
C71 minus.n26 a_n2158_n3288# 0.399137f
C72 minus.n27 a_n2158_n3288# 0.009481f
C73 minus.t8 a_n2158_n3288# 1.0008f
C74 minus.n28 a_n2158_n3288# 0.399137f
C75 minus.n29 a_n2158_n3288# 0.041782f
C76 minus.n30 a_n2158_n3288# 0.041782f
C77 minus.n31 a_n2158_n3288# 0.041782f
C78 minus.t11 a_n2158_n3288# 1.0008f
C79 minus.n32 a_n2158_n3288# 0.399137f
C80 minus.n33 a_n2158_n3288# 0.009481f
C81 minus.t6 a_n2158_n3288# 1.0008f
C82 minus.n34 a_n2158_n3288# 0.397204f
C83 minus.n35 a_n2158_n3288# 0.287284f
C84 minus.n36 a_n2158_n3288# 1.88453f
C85 source.n0 a_n2158_n3288# 0.029163f
C86 source.n1 a_n2158_n3288# 0.022016f
C87 source.n2 a_n2158_n3288# 0.01183f
C88 source.n3 a_n2158_n3288# 0.027963f
C89 source.n4 a_n2158_n3288# 0.012526f
C90 source.n5 a_n2158_n3288# 0.022016f
C91 source.n6 a_n2158_n3288# 0.01183f
C92 source.n7 a_n2158_n3288# 0.027963f
C93 source.n8 a_n2158_n3288# 0.012526f
C94 source.n9 a_n2158_n3288# 0.022016f
C95 source.n10 a_n2158_n3288# 0.012178f
C96 source.n11 a_n2158_n3288# 0.027963f
C97 source.n12 a_n2158_n3288# 0.01183f
C98 source.n13 a_n2158_n3288# 0.012526f
C99 source.n14 a_n2158_n3288# 0.022016f
C100 source.n15 a_n2158_n3288# 0.01183f
C101 source.n16 a_n2158_n3288# 0.027963f
C102 source.n17 a_n2158_n3288# 0.012526f
C103 source.n18 a_n2158_n3288# 0.022016f
C104 source.n19 a_n2158_n3288# 0.01183f
C105 source.n20 a_n2158_n3288# 0.020972f
C106 source.n21 a_n2158_n3288# 0.019768f
C107 source.t13 a_n2158_n3288# 0.047227f
C108 source.n22 a_n2158_n3288# 0.158732f
C109 source.n23 a_n2158_n3288# 1.11066f
C110 source.n24 a_n2158_n3288# 0.01183f
C111 source.n25 a_n2158_n3288# 0.012526f
C112 source.n26 a_n2158_n3288# 0.027963f
C113 source.n27 a_n2158_n3288# 0.027963f
C114 source.n28 a_n2158_n3288# 0.012526f
C115 source.n29 a_n2158_n3288# 0.01183f
C116 source.n30 a_n2158_n3288# 0.022016f
C117 source.n31 a_n2158_n3288# 0.022016f
C118 source.n32 a_n2158_n3288# 0.01183f
C119 source.n33 a_n2158_n3288# 0.012526f
C120 source.n34 a_n2158_n3288# 0.027963f
C121 source.n35 a_n2158_n3288# 0.027963f
C122 source.n36 a_n2158_n3288# 0.012526f
C123 source.n37 a_n2158_n3288# 0.01183f
C124 source.n38 a_n2158_n3288# 0.022016f
C125 source.n39 a_n2158_n3288# 0.022016f
C126 source.n40 a_n2158_n3288# 0.01183f
C127 source.n41 a_n2158_n3288# 0.012526f
C128 source.n42 a_n2158_n3288# 0.027963f
C129 source.n43 a_n2158_n3288# 0.027963f
C130 source.n44 a_n2158_n3288# 0.027963f
C131 source.n45 a_n2158_n3288# 0.012178f
C132 source.n46 a_n2158_n3288# 0.01183f
C133 source.n47 a_n2158_n3288# 0.022016f
C134 source.n48 a_n2158_n3288# 0.022016f
C135 source.n49 a_n2158_n3288# 0.01183f
C136 source.n50 a_n2158_n3288# 0.012526f
C137 source.n51 a_n2158_n3288# 0.027963f
C138 source.n52 a_n2158_n3288# 0.027963f
C139 source.n53 a_n2158_n3288# 0.012526f
C140 source.n54 a_n2158_n3288# 0.01183f
C141 source.n55 a_n2158_n3288# 0.022016f
C142 source.n56 a_n2158_n3288# 0.022016f
C143 source.n57 a_n2158_n3288# 0.01183f
C144 source.n58 a_n2158_n3288# 0.012526f
C145 source.n59 a_n2158_n3288# 0.027963f
C146 source.n60 a_n2158_n3288# 0.057382f
C147 source.n61 a_n2158_n3288# 0.012526f
C148 source.n62 a_n2158_n3288# 0.01183f
C149 source.n63 a_n2158_n3288# 0.047279f
C150 source.n64 a_n2158_n3288# 0.031669f
C151 source.n65 a_n2158_n3288# 0.926127f
C152 source.t14 a_n2158_n3288# 0.208771f
C153 source.t18 a_n2158_n3288# 0.208771f
C154 source.n66 a_n2158_n3288# 1.7875f
C155 source.n67 a_n2158_n3288# 0.351064f
C156 source.t12 a_n2158_n3288# 0.208771f
C157 source.t19 a_n2158_n3288# 0.208771f
C158 source.n68 a_n2158_n3288# 1.7875f
C159 source.n69 a_n2158_n3288# 0.351064f
C160 source.n70 a_n2158_n3288# 0.029163f
C161 source.n71 a_n2158_n3288# 0.022016f
C162 source.n72 a_n2158_n3288# 0.01183f
C163 source.n73 a_n2158_n3288# 0.027963f
C164 source.n74 a_n2158_n3288# 0.012526f
C165 source.n75 a_n2158_n3288# 0.022016f
C166 source.n76 a_n2158_n3288# 0.01183f
C167 source.n77 a_n2158_n3288# 0.027963f
C168 source.n78 a_n2158_n3288# 0.012526f
C169 source.n79 a_n2158_n3288# 0.022016f
C170 source.n80 a_n2158_n3288# 0.012178f
C171 source.n81 a_n2158_n3288# 0.027963f
C172 source.n82 a_n2158_n3288# 0.01183f
C173 source.n83 a_n2158_n3288# 0.012526f
C174 source.n84 a_n2158_n3288# 0.022016f
C175 source.n85 a_n2158_n3288# 0.01183f
C176 source.n86 a_n2158_n3288# 0.027963f
C177 source.n87 a_n2158_n3288# 0.012526f
C178 source.n88 a_n2158_n3288# 0.022016f
C179 source.n89 a_n2158_n3288# 0.01183f
C180 source.n90 a_n2158_n3288# 0.020972f
C181 source.n91 a_n2158_n3288# 0.019768f
C182 source.t17 a_n2158_n3288# 0.047227f
C183 source.n92 a_n2158_n3288# 0.158732f
C184 source.n93 a_n2158_n3288# 1.11066f
C185 source.n94 a_n2158_n3288# 0.01183f
C186 source.n95 a_n2158_n3288# 0.012526f
C187 source.n96 a_n2158_n3288# 0.027963f
C188 source.n97 a_n2158_n3288# 0.027963f
C189 source.n98 a_n2158_n3288# 0.012526f
C190 source.n99 a_n2158_n3288# 0.01183f
C191 source.n100 a_n2158_n3288# 0.022016f
C192 source.n101 a_n2158_n3288# 0.022016f
C193 source.n102 a_n2158_n3288# 0.01183f
C194 source.n103 a_n2158_n3288# 0.012526f
C195 source.n104 a_n2158_n3288# 0.027963f
C196 source.n105 a_n2158_n3288# 0.027963f
C197 source.n106 a_n2158_n3288# 0.012526f
C198 source.n107 a_n2158_n3288# 0.01183f
C199 source.n108 a_n2158_n3288# 0.022016f
C200 source.n109 a_n2158_n3288# 0.022016f
C201 source.n110 a_n2158_n3288# 0.01183f
C202 source.n111 a_n2158_n3288# 0.012526f
C203 source.n112 a_n2158_n3288# 0.027963f
C204 source.n113 a_n2158_n3288# 0.027963f
C205 source.n114 a_n2158_n3288# 0.027963f
C206 source.n115 a_n2158_n3288# 0.012178f
C207 source.n116 a_n2158_n3288# 0.01183f
C208 source.n117 a_n2158_n3288# 0.022016f
C209 source.n118 a_n2158_n3288# 0.022016f
C210 source.n119 a_n2158_n3288# 0.01183f
C211 source.n120 a_n2158_n3288# 0.012526f
C212 source.n121 a_n2158_n3288# 0.027963f
C213 source.n122 a_n2158_n3288# 0.027963f
C214 source.n123 a_n2158_n3288# 0.012526f
C215 source.n124 a_n2158_n3288# 0.01183f
C216 source.n125 a_n2158_n3288# 0.022016f
C217 source.n126 a_n2158_n3288# 0.022016f
C218 source.n127 a_n2158_n3288# 0.01183f
C219 source.n128 a_n2158_n3288# 0.012526f
C220 source.n129 a_n2158_n3288# 0.027963f
C221 source.n130 a_n2158_n3288# 0.057382f
C222 source.n131 a_n2158_n3288# 0.012526f
C223 source.n132 a_n2158_n3288# 0.01183f
C224 source.n133 a_n2158_n3288# 0.047279f
C225 source.n134 a_n2158_n3288# 0.031669f
C226 source.n135 a_n2158_n3288# 0.11309f
C227 source.n136 a_n2158_n3288# 0.029163f
C228 source.n137 a_n2158_n3288# 0.022016f
C229 source.n138 a_n2158_n3288# 0.01183f
C230 source.n139 a_n2158_n3288# 0.027963f
C231 source.n140 a_n2158_n3288# 0.012526f
C232 source.n141 a_n2158_n3288# 0.022016f
C233 source.n142 a_n2158_n3288# 0.01183f
C234 source.n143 a_n2158_n3288# 0.027963f
C235 source.n144 a_n2158_n3288# 0.012526f
C236 source.n145 a_n2158_n3288# 0.022016f
C237 source.n146 a_n2158_n3288# 0.012178f
C238 source.n147 a_n2158_n3288# 0.027963f
C239 source.n148 a_n2158_n3288# 0.01183f
C240 source.n149 a_n2158_n3288# 0.012526f
C241 source.n150 a_n2158_n3288# 0.022016f
C242 source.n151 a_n2158_n3288# 0.01183f
C243 source.n152 a_n2158_n3288# 0.027963f
C244 source.n153 a_n2158_n3288# 0.012526f
C245 source.n154 a_n2158_n3288# 0.022016f
C246 source.n155 a_n2158_n3288# 0.01183f
C247 source.n156 a_n2158_n3288# 0.020972f
C248 source.n157 a_n2158_n3288# 0.019768f
C249 source.t7 a_n2158_n3288# 0.047227f
C250 source.n158 a_n2158_n3288# 0.158732f
C251 source.n159 a_n2158_n3288# 1.11066f
C252 source.n160 a_n2158_n3288# 0.01183f
C253 source.n161 a_n2158_n3288# 0.012526f
C254 source.n162 a_n2158_n3288# 0.027963f
C255 source.n163 a_n2158_n3288# 0.027963f
C256 source.n164 a_n2158_n3288# 0.012526f
C257 source.n165 a_n2158_n3288# 0.01183f
C258 source.n166 a_n2158_n3288# 0.022016f
C259 source.n167 a_n2158_n3288# 0.022016f
C260 source.n168 a_n2158_n3288# 0.01183f
C261 source.n169 a_n2158_n3288# 0.012526f
C262 source.n170 a_n2158_n3288# 0.027963f
C263 source.n171 a_n2158_n3288# 0.027963f
C264 source.n172 a_n2158_n3288# 0.012526f
C265 source.n173 a_n2158_n3288# 0.01183f
C266 source.n174 a_n2158_n3288# 0.022016f
C267 source.n175 a_n2158_n3288# 0.022016f
C268 source.n176 a_n2158_n3288# 0.01183f
C269 source.n177 a_n2158_n3288# 0.012526f
C270 source.n178 a_n2158_n3288# 0.027963f
C271 source.n179 a_n2158_n3288# 0.027963f
C272 source.n180 a_n2158_n3288# 0.027963f
C273 source.n181 a_n2158_n3288# 0.012178f
C274 source.n182 a_n2158_n3288# 0.01183f
C275 source.n183 a_n2158_n3288# 0.022016f
C276 source.n184 a_n2158_n3288# 0.022016f
C277 source.n185 a_n2158_n3288# 0.01183f
C278 source.n186 a_n2158_n3288# 0.012526f
C279 source.n187 a_n2158_n3288# 0.027963f
C280 source.n188 a_n2158_n3288# 0.027963f
C281 source.n189 a_n2158_n3288# 0.012526f
C282 source.n190 a_n2158_n3288# 0.01183f
C283 source.n191 a_n2158_n3288# 0.022016f
C284 source.n192 a_n2158_n3288# 0.022016f
C285 source.n193 a_n2158_n3288# 0.01183f
C286 source.n194 a_n2158_n3288# 0.012526f
C287 source.n195 a_n2158_n3288# 0.027963f
C288 source.n196 a_n2158_n3288# 0.057382f
C289 source.n197 a_n2158_n3288# 0.012526f
C290 source.n198 a_n2158_n3288# 0.01183f
C291 source.n199 a_n2158_n3288# 0.047279f
C292 source.n200 a_n2158_n3288# 0.031669f
C293 source.n201 a_n2158_n3288# 0.11309f
C294 source.t22 a_n2158_n3288# 0.208771f
C295 source.t3 a_n2158_n3288# 0.208771f
C296 source.n202 a_n2158_n3288# 1.7875f
C297 source.n203 a_n2158_n3288# 0.351064f
C298 source.t21 a_n2158_n3288# 0.208771f
C299 source.t4 a_n2158_n3288# 0.208771f
C300 source.n204 a_n2158_n3288# 1.7875f
C301 source.n205 a_n2158_n3288# 0.351064f
C302 source.n206 a_n2158_n3288# 0.029163f
C303 source.n207 a_n2158_n3288# 0.022016f
C304 source.n208 a_n2158_n3288# 0.01183f
C305 source.n209 a_n2158_n3288# 0.027963f
C306 source.n210 a_n2158_n3288# 0.012526f
C307 source.n211 a_n2158_n3288# 0.022016f
C308 source.n212 a_n2158_n3288# 0.01183f
C309 source.n213 a_n2158_n3288# 0.027963f
C310 source.n214 a_n2158_n3288# 0.012526f
C311 source.n215 a_n2158_n3288# 0.022016f
C312 source.n216 a_n2158_n3288# 0.012178f
C313 source.n217 a_n2158_n3288# 0.027963f
C314 source.n218 a_n2158_n3288# 0.01183f
C315 source.n219 a_n2158_n3288# 0.012526f
C316 source.n220 a_n2158_n3288# 0.022016f
C317 source.n221 a_n2158_n3288# 0.01183f
C318 source.n222 a_n2158_n3288# 0.027963f
C319 source.n223 a_n2158_n3288# 0.012526f
C320 source.n224 a_n2158_n3288# 0.022016f
C321 source.n225 a_n2158_n3288# 0.01183f
C322 source.n226 a_n2158_n3288# 0.020972f
C323 source.n227 a_n2158_n3288# 0.019768f
C324 source.t8 a_n2158_n3288# 0.047227f
C325 source.n228 a_n2158_n3288# 0.158732f
C326 source.n229 a_n2158_n3288# 1.11066f
C327 source.n230 a_n2158_n3288# 0.01183f
C328 source.n231 a_n2158_n3288# 0.012526f
C329 source.n232 a_n2158_n3288# 0.027963f
C330 source.n233 a_n2158_n3288# 0.027963f
C331 source.n234 a_n2158_n3288# 0.012526f
C332 source.n235 a_n2158_n3288# 0.01183f
C333 source.n236 a_n2158_n3288# 0.022016f
C334 source.n237 a_n2158_n3288# 0.022016f
C335 source.n238 a_n2158_n3288# 0.01183f
C336 source.n239 a_n2158_n3288# 0.012526f
C337 source.n240 a_n2158_n3288# 0.027963f
C338 source.n241 a_n2158_n3288# 0.027963f
C339 source.n242 a_n2158_n3288# 0.012526f
C340 source.n243 a_n2158_n3288# 0.01183f
C341 source.n244 a_n2158_n3288# 0.022016f
C342 source.n245 a_n2158_n3288# 0.022016f
C343 source.n246 a_n2158_n3288# 0.01183f
C344 source.n247 a_n2158_n3288# 0.012526f
C345 source.n248 a_n2158_n3288# 0.027963f
C346 source.n249 a_n2158_n3288# 0.027963f
C347 source.n250 a_n2158_n3288# 0.027963f
C348 source.n251 a_n2158_n3288# 0.012178f
C349 source.n252 a_n2158_n3288# 0.01183f
C350 source.n253 a_n2158_n3288# 0.022016f
C351 source.n254 a_n2158_n3288# 0.022016f
C352 source.n255 a_n2158_n3288# 0.01183f
C353 source.n256 a_n2158_n3288# 0.012526f
C354 source.n257 a_n2158_n3288# 0.027963f
C355 source.n258 a_n2158_n3288# 0.027963f
C356 source.n259 a_n2158_n3288# 0.012526f
C357 source.n260 a_n2158_n3288# 0.01183f
C358 source.n261 a_n2158_n3288# 0.022016f
C359 source.n262 a_n2158_n3288# 0.022016f
C360 source.n263 a_n2158_n3288# 0.01183f
C361 source.n264 a_n2158_n3288# 0.012526f
C362 source.n265 a_n2158_n3288# 0.027963f
C363 source.n266 a_n2158_n3288# 0.057382f
C364 source.n267 a_n2158_n3288# 0.012526f
C365 source.n268 a_n2158_n3288# 0.01183f
C366 source.n269 a_n2158_n3288# 0.047279f
C367 source.n270 a_n2158_n3288# 0.031669f
C368 source.n271 a_n2158_n3288# 1.28113f
C369 source.n272 a_n2158_n3288# 0.029163f
C370 source.n273 a_n2158_n3288# 0.022016f
C371 source.n274 a_n2158_n3288# 0.01183f
C372 source.n275 a_n2158_n3288# 0.027963f
C373 source.n276 a_n2158_n3288# 0.012526f
C374 source.n277 a_n2158_n3288# 0.022016f
C375 source.n278 a_n2158_n3288# 0.01183f
C376 source.n279 a_n2158_n3288# 0.027963f
C377 source.n280 a_n2158_n3288# 0.012526f
C378 source.n281 a_n2158_n3288# 0.022016f
C379 source.n282 a_n2158_n3288# 0.012178f
C380 source.n283 a_n2158_n3288# 0.027963f
C381 source.n284 a_n2158_n3288# 0.012526f
C382 source.n285 a_n2158_n3288# 0.022016f
C383 source.n286 a_n2158_n3288# 0.01183f
C384 source.n287 a_n2158_n3288# 0.027963f
C385 source.n288 a_n2158_n3288# 0.012526f
C386 source.n289 a_n2158_n3288# 0.022016f
C387 source.n290 a_n2158_n3288# 0.01183f
C388 source.n291 a_n2158_n3288# 0.020972f
C389 source.n292 a_n2158_n3288# 0.019768f
C390 source.t20 a_n2158_n3288# 0.047227f
C391 source.n293 a_n2158_n3288# 0.158732f
C392 source.n294 a_n2158_n3288# 1.11066f
C393 source.n295 a_n2158_n3288# 0.01183f
C394 source.n296 a_n2158_n3288# 0.012526f
C395 source.n297 a_n2158_n3288# 0.027963f
C396 source.n298 a_n2158_n3288# 0.027963f
C397 source.n299 a_n2158_n3288# 0.012526f
C398 source.n300 a_n2158_n3288# 0.01183f
C399 source.n301 a_n2158_n3288# 0.022016f
C400 source.n302 a_n2158_n3288# 0.022016f
C401 source.n303 a_n2158_n3288# 0.01183f
C402 source.n304 a_n2158_n3288# 0.012526f
C403 source.n305 a_n2158_n3288# 0.027963f
C404 source.n306 a_n2158_n3288# 0.027963f
C405 source.n307 a_n2158_n3288# 0.012526f
C406 source.n308 a_n2158_n3288# 0.01183f
C407 source.n309 a_n2158_n3288# 0.022016f
C408 source.n310 a_n2158_n3288# 0.022016f
C409 source.n311 a_n2158_n3288# 0.01183f
C410 source.n312 a_n2158_n3288# 0.01183f
C411 source.n313 a_n2158_n3288# 0.012526f
C412 source.n314 a_n2158_n3288# 0.027963f
C413 source.n315 a_n2158_n3288# 0.027963f
C414 source.n316 a_n2158_n3288# 0.027963f
C415 source.n317 a_n2158_n3288# 0.012178f
C416 source.n318 a_n2158_n3288# 0.01183f
C417 source.n319 a_n2158_n3288# 0.022016f
C418 source.n320 a_n2158_n3288# 0.022016f
C419 source.n321 a_n2158_n3288# 0.01183f
C420 source.n322 a_n2158_n3288# 0.012526f
C421 source.n323 a_n2158_n3288# 0.027963f
C422 source.n324 a_n2158_n3288# 0.027963f
C423 source.n325 a_n2158_n3288# 0.012526f
C424 source.n326 a_n2158_n3288# 0.01183f
C425 source.n327 a_n2158_n3288# 0.022016f
C426 source.n328 a_n2158_n3288# 0.022016f
C427 source.n329 a_n2158_n3288# 0.01183f
C428 source.n330 a_n2158_n3288# 0.012526f
C429 source.n331 a_n2158_n3288# 0.027963f
C430 source.n332 a_n2158_n3288# 0.057382f
C431 source.n333 a_n2158_n3288# 0.012526f
C432 source.n334 a_n2158_n3288# 0.01183f
C433 source.n335 a_n2158_n3288# 0.047279f
C434 source.n336 a_n2158_n3288# 0.031669f
C435 source.n337 a_n2158_n3288# 1.28113f
C436 source.t15 a_n2158_n3288# 0.208771f
C437 source.t16 a_n2158_n3288# 0.208771f
C438 source.n338 a_n2158_n3288# 1.78749f
C439 source.n339 a_n2158_n3288# 0.351075f
C440 source.t11 a_n2158_n3288# 0.208771f
C441 source.t9 a_n2158_n3288# 0.208771f
C442 source.n340 a_n2158_n3288# 1.78749f
C443 source.n341 a_n2158_n3288# 0.351075f
C444 source.n342 a_n2158_n3288# 0.029163f
C445 source.n343 a_n2158_n3288# 0.022016f
C446 source.n344 a_n2158_n3288# 0.01183f
C447 source.n345 a_n2158_n3288# 0.027963f
C448 source.n346 a_n2158_n3288# 0.012526f
C449 source.n347 a_n2158_n3288# 0.022016f
C450 source.n348 a_n2158_n3288# 0.01183f
C451 source.n349 a_n2158_n3288# 0.027963f
C452 source.n350 a_n2158_n3288# 0.012526f
C453 source.n351 a_n2158_n3288# 0.022016f
C454 source.n352 a_n2158_n3288# 0.012178f
C455 source.n353 a_n2158_n3288# 0.027963f
C456 source.n354 a_n2158_n3288# 0.012526f
C457 source.n355 a_n2158_n3288# 0.022016f
C458 source.n356 a_n2158_n3288# 0.01183f
C459 source.n357 a_n2158_n3288# 0.027963f
C460 source.n358 a_n2158_n3288# 0.012526f
C461 source.n359 a_n2158_n3288# 0.022016f
C462 source.n360 a_n2158_n3288# 0.01183f
C463 source.n361 a_n2158_n3288# 0.020972f
C464 source.n362 a_n2158_n3288# 0.019768f
C465 source.t10 a_n2158_n3288# 0.047227f
C466 source.n363 a_n2158_n3288# 0.158732f
C467 source.n364 a_n2158_n3288# 1.11066f
C468 source.n365 a_n2158_n3288# 0.01183f
C469 source.n366 a_n2158_n3288# 0.012526f
C470 source.n367 a_n2158_n3288# 0.027963f
C471 source.n368 a_n2158_n3288# 0.027963f
C472 source.n369 a_n2158_n3288# 0.012526f
C473 source.n370 a_n2158_n3288# 0.01183f
C474 source.n371 a_n2158_n3288# 0.022016f
C475 source.n372 a_n2158_n3288# 0.022016f
C476 source.n373 a_n2158_n3288# 0.01183f
C477 source.n374 a_n2158_n3288# 0.012526f
C478 source.n375 a_n2158_n3288# 0.027963f
C479 source.n376 a_n2158_n3288# 0.027963f
C480 source.n377 a_n2158_n3288# 0.012526f
C481 source.n378 a_n2158_n3288# 0.01183f
C482 source.n379 a_n2158_n3288# 0.022016f
C483 source.n380 a_n2158_n3288# 0.022016f
C484 source.n381 a_n2158_n3288# 0.01183f
C485 source.n382 a_n2158_n3288# 0.01183f
C486 source.n383 a_n2158_n3288# 0.012526f
C487 source.n384 a_n2158_n3288# 0.027963f
C488 source.n385 a_n2158_n3288# 0.027963f
C489 source.n386 a_n2158_n3288# 0.027963f
C490 source.n387 a_n2158_n3288# 0.012178f
C491 source.n388 a_n2158_n3288# 0.01183f
C492 source.n389 a_n2158_n3288# 0.022016f
C493 source.n390 a_n2158_n3288# 0.022016f
C494 source.n391 a_n2158_n3288# 0.01183f
C495 source.n392 a_n2158_n3288# 0.012526f
C496 source.n393 a_n2158_n3288# 0.027963f
C497 source.n394 a_n2158_n3288# 0.027963f
C498 source.n395 a_n2158_n3288# 0.012526f
C499 source.n396 a_n2158_n3288# 0.01183f
C500 source.n397 a_n2158_n3288# 0.022016f
C501 source.n398 a_n2158_n3288# 0.022016f
C502 source.n399 a_n2158_n3288# 0.01183f
C503 source.n400 a_n2158_n3288# 0.012526f
C504 source.n401 a_n2158_n3288# 0.027963f
C505 source.n402 a_n2158_n3288# 0.057382f
C506 source.n403 a_n2158_n3288# 0.012526f
C507 source.n404 a_n2158_n3288# 0.01183f
C508 source.n405 a_n2158_n3288# 0.047279f
C509 source.n406 a_n2158_n3288# 0.031669f
C510 source.n407 a_n2158_n3288# 0.11309f
C511 source.n408 a_n2158_n3288# 0.029163f
C512 source.n409 a_n2158_n3288# 0.022016f
C513 source.n410 a_n2158_n3288# 0.01183f
C514 source.n411 a_n2158_n3288# 0.027963f
C515 source.n412 a_n2158_n3288# 0.012526f
C516 source.n413 a_n2158_n3288# 0.022016f
C517 source.n414 a_n2158_n3288# 0.01183f
C518 source.n415 a_n2158_n3288# 0.027963f
C519 source.n416 a_n2158_n3288# 0.012526f
C520 source.n417 a_n2158_n3288# 0.022016f
C521 source.n418 a_n2158_n3288# 0.012178f
C522 source.n419 a_n2158_n3288# 0.027963f
C523 source.n420 a_n2158_n3288# 0.012526f
C524 source.n421 a_n2158_n3288# 0.022016f
C525 source.n422 a_n2158_n3288# 0.01183f
C526 source.n423 a_n2158_n3288# 0.027963f
C527 source.n424 a_n2158_n3288# 0.012526f
C528 source.n425 a_n2158_n3288# 0.022016f
C529 source.n426 a_n2158_n3288# 0.01183f
C530 source.n427 a_n2158_n3288# 0.020972f
C531 source.n428 a_n2158_n3288# 0.019768f
C532 source.t23 a_n2158_n3288# 0.047227f
C533 source.n429 a_n2158_n3288# 0.158732f
C534 source.n430 a_n2158_n3288# 1.11066f
C535 source.n431 a_n2158_n3288# 0.01183f
C536 source.n432 a_n2158_n3288# 0.012526f
C537 source.n433 a_n2158_n3288# 0.027963f
C538 source.n434 a_n2158_n3288# 0.027963f
C539 source.n435 a_n2158_n3288# 0.012526f
C540 source.n436 a_n2158_n3288# 0.01183f
C541 source.n437 a_n2158_n3288# 0.022016f
C542 source.n438 a_n2158_n3288# 0.022016f
C543 source.n439 a_n2158_n3288# 0.01183f
C544 source.n440 a_n2158_n3288# 0.012526f
C545 source.n441 a_n2158_n3288# 0.027963f
C546 source.n442 a_n2158_n3288# 0.027963f
C547 source.n443 a_n2158_n3288# 0.012526f
C548 source.n444 a_n2158_n3288# 0.01183f
C549 source.n445 a_n2158_n3288# 0.022016f
C550 source.n446 a_n2158_n3288# 0.022016f
C551 source.n447 a_n2158_n3288# 0.01183f
C552 source.n448 a_n2158_n3288# 0.01183f
C553 source.n449 a_n2158_n3288# 0.012526f
C554 source.n450 a_n2158_n3288# 0.027963f
C555 source.n451 a_n2158_n3288# 0.027963f
C556 source.n452 a_n2158_n3288# 0.027963f
C557 source.n453 a_n2158_n3288# 0.012178f
C558 source.n454 a_n2158_n3288# 0.01183f
C559 source.n455 a_n2158_n3288# 0.022016f
C560 source.n456 a_n2158_n3288# 0.022016f
C561 source.n457 a_n2158_n3288# 0.01183f
C562 source.n458 a_n2158_n3288# 0.012526f
C563 source.n459 a_n2158_n3288# 0.027963f
C564 source.n460 a_n2158_n3288# 0.027963f
C565 source.n461 a_n2158_n3288# 0.012526f
C566 source.n462 a_n2158_n3288# 0.01183f
C567 source.n463 a_n2158_n3288# 0.022016f
C568 source.n464 a_n2158_n3288# 0.022016f
C569 source.n465 a_n2158_n3288# 0.01183f
C570 source.n466 a_n2158_n3288# 0.012526f
C571 source.n467 a_n2158_n3288# 0.027963f
C572 source.n468 a_n2158_n3288# 0.057382f
C573 source.n469 a_n2158_n3288# 0.012526f
C574 source.n470 a_n2158_n3288# 0.01183f
C575 source.n471 a_n2158_n3288# 0.047279f
C576 source.n472 a_n2158_n3288# 0.031669f
C577 source.n473 a_n2158_n3288# 0.11309f
C578 source.t2 a_n2158_n3288# 0.208771f
C579 source.t1 a_n2158_n3288# 0.208771f
C580 source.n474 a_n2158_n3288# 1.78749f
C581 source.n475 a_n2158_n3288# 0.351075f
C582 source.t6 a_n2158_n3288# 0.208771f
C583 source.t5 a_n2158_n3288# 0.208771f
C584 source.n476 a_n2158_n3288# 1.78749f
C585 source.n477 a_n2158_n3288# 0.351075f
C586 source.n478 a_n2158_n3288# 0.029163f
C587 source.n479 a_n2158_n3288# 0.022016f
C588 source.n480 a_n2158_n3288# 0.01183f
C589 source.n481 a_n2158_n3288# 0.027963f
C590 source.n482 a_n2158_n3288# 0.012526f
C591 source.n483 a_n2158_n3288# 0.022016f
C592 source.n484 a_n2158_n3288# 0.01183f
C593 source.n485 a_n2158_n3288# 0.027963f
C594 source.n486 a_n2158_n3288# 0.012526f
C595 source.n487 a_n2158_n3288# 0.022016f
C596 source.n488 a_n2158_n3288# 0.012178f
C597 source.n489 a_n2158_n3288# 0.027963f
C598 source.n490 a_n2158_n3288# 0.012526f
C599 source.n491 a_n2158_n3288# 0.022016f
C600 source.n492 a_n2158_n3288# 0.01183f
C601 source.n493 a_n2158_n3288# 0.027963f
C602 source.n494 a_n2158_n3288# 0.012526f
C603 source.n495 a_n2158_n3288# 0.022016f
C604 source.n496 a_n2158_n3288# 0.01183f
C605 source.n497 a_n2158_n3288# 0.020972f
C606 source.n498 a_n2158_n3288# 0.019768f
C607 source.t0 a_n2158_n3288# 0.047227f
C608 source.n499 a_n2158_n3288# 0.158732f
C609 source.n500 a_n2158_n3288# 1.11066f
C610 source.n501 a_n2158_n3288# 0.01183f
C611 source.n502 a_n2158_n3288# 0.012526f
C612 source.n503 a_n2158_n3288# 0.027963f
C613 source.n504 a_n2158_n3288# 0.027963f
C614 source.n505 a_n2158_n3288# 0.012526f
C615 source.n506 a_n2158_n3288# 0.01183f
C616 source.n507 a_n2158_n3288# 0.022016f
C617 source.n508 a_n2158_n3288# 0.022016f
C618 source.n509 a_n2158_n3288# 0.01183f
C619 source.n510 a_n2158_n3288# 0.012526f
C620 source.n511 a_n2158_n3288# 0.027963f
C621 source.n512 a_n2158_n3288# 0.027963f
C622 source.n513 a_n2158_n3288# 0.012526f
C623 source.n514 a_n2158_n3288# 0.01183f
C624 source.n515 a_n2158_n3288# 0.022016f
C625 source.n516 a_n2158_n3288# 0.022016f
C626 source.n517 a_n2158_n3288# 0.01183f
C627 source.n518 a_n2158_n3288# 0.01183f
C628 source.n519 a_n2158_n3288# 0.012526f
C629 source.n520 a_n2158_n3288# 0.027963f
C630 source.n521 a_n2158_n3288# 0.027963f
C631 source.n522 a_n2158_n3288# 0.027963f
C632 source.n523 a_n2158_n3288# 0.012178f
C633 source.n524 a_n2158_n3288# 0.01183f
C634 source.n525 a_n2158_n3288# 0.022016f
C635 source.n526 a_n2158_n3288# 0.022016f
C636 source.n527 a_n2158_n3288# 0.01183f
C637 source.n528 a_n2158_n3288# 0.012526f
C638 source.n529 a_n2158_n3288# 0.027963f
C639 source.n530 a_n2158_n3288# 0.027963f
C640 source.n531 a_n2158_n3288# 0.012526f
C641 source.n532 a_n2158_n3288# 0.01183f
C642 source.n533 a_n2158_n3288# 0.022016f
C643 source.n534 a_n2158_n3288# 0.022016f
C644 source.n535 a_n2158_n3288# 0.01183f
C645 source.n536 a_n2158_n3288# 0.012526f
C646 source.n537 a_n2158_n3288# 0.027963f
C647 source.n538 a_n2158_n3288# 0.057382f
C648 source.n539 a_n2158_n3288# 0.012526f
C649 source.n540 a_n2158_n3288# 0.01183f
C650 source.n541 a_n2158_n3288# 0.047279f
C651 source.n542 a_n2158_n3288# 0.031669f
C652 source.n543 a_n2158_n3288# 0.2567f
C653 source.n544 a_n2158_n3288# 1.3951f
C654 drain_left.t6 a_n2158_n3288# 0.258116f
C655 drain_left.t10 a_n2158_n3288# 0.258116f
C656 drain_left.n0 a_n2158_n3288# 2.30223f
C657 drain_left.t9 a_n2158_n3288# 0.258116f
C658 drain_left.t4 a_n2158_n3288# 0.258116f
C659 drain_left.n1 a_n2158_n3288# 2.29683f
C660 drain_left.t3 a_n2158_n3288# 0.258116f
C661 drain_left.t1 a_n2158_n3288# 0.258116f
C662 drain_left.n2 a_n2158_n3288# 2.30223f
C663 drain_left.n3 a_n2158_n3288# 2.52598f
C664 drain_left.t11 a_n2158_n3288# 0.258116f
C665 drain_left.t2 a_n2158_n3288# 0.258116f
C666 drain_left.n4 a_n2158_n3288# 2.30265f
C667 drain_left.t5 a_n2158_n3288# 0.258116f
C668 drain_left.t7 a_n2158_n3288# 0.258116f
C669 drain_left.n5 a_n2158_n3288# 2.29684f
C670 drain_left.n6 a_n2158_n3288# 0.773534f
C671 drain_left.t8 a_n2158_n3288# 0.258116f
C672 drain_left.t0 a_n2158_n3288# 0.258116f
C673 drain_left.n7 a_n2158_n3288# 2.29683f
C674 drain_left.n8 a_n2158_n3288# 0.624955f
C675 plus.n0 a_n2158_n3288# 0.042337f
C676 plus.t7 a_n2158_n3288# 1.01409f
C677 plus.t2 a_n2158_n3288# 1.01409f
C678 plus.n1 a_n2158_n3288# 0.042337f
C679 plus.t6 a_n2158_n3288# 1.01409f
C680 plus.n2 a_n2158_n3288# 0.404439f
C681 plus.n3 a_n2158_n3288# 0.042337f
C682 plus.t1 a_n2158_n3288# 1.01409f
C683 plus.t8 a_n2158_n3288# 1.01409f
C684 plus.n4 a_n2158_n3288# 0.409174f
C685 plus.t3 a_n2158_n3288# 1.03322f
C686 plus.n5 a_n2158_n3288# 0.389097f
C687 plus.n6 a_n2158_n3288# 0.17761f
C688 plus.n7 a_n2158_n3288# 0.009607f
C689 plus.n8 a_n2158_n3288# 0.404439f
C690 plus.n9 a_n2158_n3288# 0.009607f
C691 plus.n10 a_n2158_n3288# 0.042337f
C692 plus.n11 a_n2158_n3288# 0.042337f
C693 plus.n12 a_n2158_n3288# 0.042337f
C694 plus.n13 a_n2158_n3288# 0.009607f
C695 plus.n14 a_n2158_n3288# 0.404439f
C696 plus.n15 a_n2158_n3288# 0.009607f
C697 plus.n16 a_n2158_n3288# 0.402481f
C698 plus.n17 a_n2158_n3288# 0.488256f
C699 plus.n18 a_n2158_n3288# 0.042337f
C700 plus.t0 a_n2158_n3288# 1.01409f
C701 plus.n19 a_n2158_n3288# 0.042337f
C702 plus.t5 a_n2158_n3288# 1.01409f
C703 plus.t4 a_n2158_n3288# 1.01409f
C704 plus.n20 a_n2158_n3288# 0.404439f
C705 plus.n21 a_n2158_n3288# 0.042337f
C706 plus.t9 a_n2158_n3288# 1.01409f
C707 plus.t11 a_n2158_n3288# 1.01409f
C708 plus.n22 a_n2158_n3288# 0.409174f
C709 plus.t10 a_n2158_n3288# 1.03322f
C710 plus.n23 a_n2158_n3288# 0.389097f
C711 plus.n24 a_n2158_n3288# 0.17761f
C712 plus.n25 a_n2158_n3288# 0.009607f
C713 plus.n26 a_n2158_n3288# 0.404439f
C714 plus.n27 a_n2158_n3288# 0.009607f
C715 plus.n28 a_n2158_n3288# 0.042337f
C716 plus.n29 a_n2158_n3288# 0.042337f
C717 plus.n30 a_n2158_n3288# 0.042337f
C718 plus.n31 a_n2158_n3288# 0.009607f
C719 plus.n32 a_n2158_n3288# 0.404439f
C720 plus.n33 a_n2158_n3288# 0.009607f
C721 plus.n34 a_n2158_n3288# 0.402481f
C722 plus.n35 a_n2158_n3288# 1.34298f
.ends

