* NGSPICE file created from diffpair511.ext - technology: sky130A

.subckt diffpair511 minus drain_right drain_left source plus
X0 drain_right minus source a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X1 source plus drain_left a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X2 drain_right minus source a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X3 source minus drain_right a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X4 a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X5 drain_left plus source a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X6 a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X7 source minus drain_right a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X8 a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X9 source plus drain_left a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X10 a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X11 drain_left plus source a_n1094_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
.ends

