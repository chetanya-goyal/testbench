* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t4 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 source.t26 plus.t1 drain_left.t5 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t2 plus.t2 source.t25 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t24 plus.t3 drain_left.t0 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X5 source.t0 minus.t0 drain_right.t13 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 source.t12 minus.t1 drain_right.t12 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X7 source.t23 plus.t4 drain_left.t6 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X8 drain_left.t3 plus.t5 source.t22 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X9 source.t2 minus.t2 drain_right.t11 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X10 source.t8 minus.t3 drain_right.t10 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X11 source.t10 minus.t4 drain_right.t9 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 drain_right.t8 minus.t5 source.t6 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X13 drain_left.t1 plus.t6 source.t21 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X14 drain_left.t7 plus.t7 source.t20 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X15 drain_left.t9 plus.t8 source.t19 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X16 drain_right.t7 minus.t6 source.t13 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X17 drain_right.t6 minus.t7 source.t7 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X18 a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X19 drain_right.t5 minus.t8 source.t9 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X20 drain_right.t4 minus.t9 source.t11 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X21 drain_right.t3 minus.t10 source.t4 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X22 a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X23 source.t1 minus.t11 drain_right.t2 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X24 source.t18 plus.t9 drain_left.t10 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X25 drain_right.t1 minus.t12 source.t3 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X26 drain_right.t0 minus.t13 source.t5 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X27 drain_left.t8 plus.t10 source.t17 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X28 drain_left.t13 plus.t11 source.t16 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X29 source.t15 plus.t12 drain_left.t11 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X30 a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X31 drain_left.t12 plus.t13 source.t14 a_n1644_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
R0 plus.n3 plus.t5 353.175
R1 plus.n15 plus.t6 353.175
R2 plus.n20 plus.t11 353.175
R3 plus.n32 plus.t13 353.175
R4 plus.n1 plus.t0 318.12
R5 plus.n4 plus.t1 318.12
R6 plus.n6 plus.t8 318.12
R7 plus.n12 plus.t7 318.12
R8 plus.n14 plus.t12 318.12
R9 plus.n18 plus.t4 318.12
R10 plus.n21 plus.t9 318.12
R11 plus.n23 plus.t2 318.12
R12 plus.n29 plus.t10 318.12
R13 plus.n31 plus.t3 318.12
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 25.393
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus.n7 plus.n6 11.6853
R46 plus.n12 plus.n11 11.6853
R47 plus.n29 plus.n28 11.6853
R48 plus.n24 plus.n23 11.6853
R49 plus plus.n16 8.30732
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n2 drain_left.n0 289.615
R61 drain_left.n15 drain_left.n13 289.615
R62 drain_left.n3 drain_left.n2 185
R63 drain_left.n16 drain_left.n15 185
R64 drain_left.t12 drain_left.n1 167.117
R65 drain_left.t3 drain_left.n14 167.117
R66 drain_left.n11 drain_left.n9 101.296
R67 drain_left.n25 drain_left.n24 100.796
R68 drain_left.n23 drain_left.n22 100.796
R69 drain_left.n21 drain_left.n20 100.796
R70 drain_left.n11 drain_left.n10 100.796
R71 drain_left.n8 drain_left.n7 100.796
R72 drain_left.n2 drain_left.t12 52.3082
R73 drain_left.n15 drain_left.t3 52.3082
R74 drain_left.n8 drain_left.n6 48.5884
R75 drain_left.n21 drain_left.n19 48.5884
R76 drain_left drain_left.n12 22.6663
R77 drain_left.n9 drain_left.t10 9.9005
R78 drain_left.n9 drain_left.t13 9.9005
R79 drain_left.n10 drain_left.t6 9.9005
R80 drain_left.n10 drain_left.t2 9.9005
R81 drain_left.n7 drain_left.t0 9.9005
R82 drain_left.n7 drain_left.t8 9.9005
R83 drain_left.n24 drain_left.t11 9.9005
R84 drain_left.n24 drain_left.t1 9.9005
R85 drain_left.n22 drain_left.t4 9.9005
R86 drain_left.n22 drain_left.t7 9.9005
R87 drain_left.n20 drain_left.t5 9.9005
R88 drain_left.n20 drain_left.t9 9.9005
R89 drain_left.n3 drain_left.n1 9.71174
R90 drain_left.n16 drain_left.n14 9.71174
R91 drain_left.n6 drain_left.n5 9.45567
R92 drain_left.n19 drain_left.n18 9.45567
R93 drain_left.n5 drain_left.n4 9.3005
R94 drain_left.n18 drain_left.n17 9.3005
R95 drain_left.n6 drain_left.n0 8.14595
R96 drain_left.n19 drain_left.n13 8.14595
R97 drain_left.n4 drain_left.n3 7.3702
R98 drain_left.n17 drain_left.n16 7.3702
R99 drain_left drain_left.n25 6.15322
R100 drain_left.n4 drain_left.n0 5.81868
R101 drain_left.n17 drain_left.n13 5.81868
R102 drain_left.n5 drain_left.n1 3.44771
R103 drain_left.n18 drain_left.n14 3.44771
R104 drain_left.n23 drain_left.n21 0.5005
R105 drain_left.n25 drain_left.n23 0.5005
R106 drain_left.n12 drain_left.n8 0.320154
R107 drain_left.n12 drain_left.n11 0.070154
R108 source.n50 source.n48 289.615
R109 source.n36 source.n34 289.615
R110 source.n2 source.n0 289.615
R111 source.n16 source.n14 289.615
R112 source.n51 source.n50 185
R113 source.n37 source.n36 185
R114 source.n3 source.n2 185
R115 source.n17 source.n16 185
R116 source.t4 source.n49 167.117
R117 source.t16 source.n35 167.117
R118 source.t21 source.n1 167.117
R119 source.t11 source.n15 167.117
R120 source.n9 source.n8 84.1169
R121 source.n11 source.n10 84.1169
R122 source.n13 source.n12 84.1169
R123 source.n23 source.n22 84.1169
R124 source.n25 source.n24 84.1169
R125 source.n27 source.n26 84.1169
R126 source.n47 source.n46 84.1168
R127 source.n45 source.n44 84.1168
R128 source.n43 source.n42 84.1168
R129 source.n33 source.n32 84.1168
R130 source.n31 source.n30 84.1168
R131 source.n29 source.n28 84.1168
R132 source.n50 source.t4 52.3082
R133 source.n36 source.t16 52.3082
R134 source.n2 source.t21 52.3082
R135 source.n16 source.t11 52.3082
R136 source.n55 source.n54 31.4096
R137 source.n41 source.n40 31.4096
R138 source.n7 source.n6 31.4096
R139 source.n21 source.n20 31.4096
R140 source.n29 source.n27 14.712
R141 source.n46 source.t13 9.9005
R142 source.n46 source.t1 9.9005
R143 source.n44 source.t6 9.9005
R144 source.n44 source.t10 9.9005
R145 source.n42 source.t7 9.9005
R146 source.n42 source.t2 9.9005
R147 source.n32 source.t25 9.9005
R148 source.n32 source.t18 9.9005
R149 source.n30 source.t17 9.9005
R150 source.n30 source.t23 9.9005
R151 source.n28 source.t14 9.9005
R152 source.n28 source.t24 9.9005
R153 source.n8 source.t20 9.9005
R154 source.n8 source.t15 9.9005
R155 source.n10 source.t19 9.9005
R156 source.n10 source.t27 9.9005
R157 source.n12 source.t22 9.9005
R158 source.n12 source.t26 9.9005
R159 source.n22 source.t9 9.9005
R160 source.n22 source.t12 9.9005
R161 source.n24 source.t3 9.9005
R162 source.n24 source.t0 9.9005
R163 source.n26 source.t5 9.9005
R164 source.n26 source.t8 9.9005
R165 source.n51 source.n49 9.71174
R166 source.n37 source.n35 9.71174
R167 source.n3 source.n1 9.71174
R168 source.n17 source.n15 9.71174
R169 source.n54 source.n53 9.45567
R170 source.n40 source.n39 9.45567
R171 source.n6 source.n5 9.45567
R172 source.n20 source.n19 9.45567
R173 source.n53 source.n52 9.3005
R174 source.n39 source.n38 9.3005
R175 source.n5 source.n4 9.3005
R176 source.n19 source.n18 9.3005
R177 source.n56 source.n7 8.69904
R178 source.n54 source.n48 8.14595
R179 source.n40 source.n34 8.14595
R180 source.n6 source.n0 8.14595
R181 source.n20 source.n14 8.14595
R182 source.n52 source.n51 7.3702
R183 source.n38 source.n37 7.3702
R184 source.n4 source.n3 7.3702
R185 source.n18 source.n17 7.3702
R186 source.n52 source.n48 5.81868
R187 source.n38 source.n34 5.81868
R188 source.n4 source.n0 5.81868
R189 source.n18 source.n14 5.81868
R190 source.n56 source.n55 5.51343
R191 source.n53 source.n49 3.44771
R192 source.n39 source.n35 3.44771
R193 source.n5 source.n1 3.44771
R194 source.n19 source.n15 3.44771
R195 source.n21 source.n13 0.720328
R196 source.n43 source.n41 0.720328
R197 source.n27 source.n25 0.5005
R198 source.n25 source.n23 0.5005
R199 source.n23 source.n21 0.5005
R200 source.n13 source.n11 0.5005
R201 source.n11 source.n9 0.5005
R202 source.n9 source.n7 0.5005
R203 source.n31 source.n29 0.5005
R204 source.n33 source.n31 0.5005
R205 source.n41 source.n33 0.5005
R206 source.n45 source.n43 0.5005
R207 source.n47 source.n45 0.5005
R208 source.n55 source.n47 0.5005
R209 source source.n56 0.188
R210 minus.n15 minus.t13 353.175
R211 minus.n3 minus.t9 353.175
R212 minus.n32 minus.t10 353.175
R213 minus.n20 minus.t7 353.175
R214 minus.n1 minus.t0 318.12
R215 minus.n14 minus.t3 318.12
R216 minus.n12 minus.t12 318.12
R217 minus.n6 minus.t8 318.12
R218 minus.n4 minus.t1 318.12
R219 minus.n18 minus.t4 318.12
R220 minus.n31 minus.t11 318.12
R221 minus.n29 minus.t6 318.12
R222 minus.n23 minus.t5 318.12
R223 minus.n21 minus.t2 318.12
R224 minus.n3 minus.n2 161.489
R225 minus.n20 minus.n19 161.489
R226 minus.n16 minus.n15 161.3
R227 minus.n13 minus.n0 161.3
R228 minus.n11 minus.n10 161.3
R229 minus.n9 minus.n1 161.3
R230 minus.n8 minus.n7 161.3
R231 minus.n5 minus.n2 161.3
R232 minus.n33 minus.n32 161.3
R233 minus.n30 minus.n17 161.3
R234 minus.n28 minus.n27 161.3
R235 minus.n26 minus.n18 161.3
R236 minus.n25 minus.n24 161.3
R237 minus.n22 minus.n19 161.3
R238 minus.n11 minus.n1 73.0308
R239 minus.n7 minus.n1 73.0308
R240 minus.n24 minus.n18 73.0308
R241 minus.n28 minus.n18 73.0308
R242 minus.n13 minus.n12 61.346
R243 minus.n6 minus.n5 61.346
R244 minus.n23 minus.n22 61.346
R245 minus.n30 minus.n29 61.346
R246 minus.n15 minus.n14 49.6611
R247 minus.n4 minus.n3 49.6611
R248 minus.n21 minus.n20 49.6611
R249 minus.n32 minus.n31 49.6611
R250 minus.n34 minus.n16 27.724
R251 minus.n14 minus.n13 23.3702
R252 minus.n5 minus.n4 23.3702
R253 minus.n22 minus.n21 23.3702
R254 minus.n31 minus.n30 23.3702
R255 minus.n12 minus.n11 11.6853
R256 minus.n7 minus.n6 11.6853
R257 minus.n24 minus.n23 11.6853
R258 minus.n29 minus.n28 11.6853
R259 minus.n34 minus.n33 6.45126
R260 minus.n16 minus.n0 0.189894
R261 minus.n10 minus.n0 0.189894
R262 minus.n10 minus.n9 0.189894
R263 minus.n9 minus.n8 0.189894
R264 minus.n8 minus.n2 0.189894
R265 minus.n25 minus.n19 0.189894
R266 minus.n26 minus.n25 0.189894
R267 minus.n27 minus.n26 0.189894
R268 minus.n27 minus.n17 0.189894
R269 minus.n33 minus.n17 0.189894
R270 minus minus.n34 0.188
R271 drain_right.n2 drain_right.n0 289.615
R272 drain_right.n20 drain_right.n18 289.615
R273 drain_right.n3 drain_right.n2 185
R274 drain_right.n21 drain_right.n20 185
R275 drain_right.t6 drain_right.n1 167.117
R276 drain_right.t0 drain_right.n19 167.117
R277 drain_right.n15 drain_right.n13 101.296
R278 drain_right.n11 drain_right.n9 101.296
R279 drain_right.n15 drain_right.n14 100.796
R280 drain_right.n17 drain_right.n16 100.796
R281 drain_right.n11 drain_right.n10 100.796
R282 drain_right.n8 drain_right.n7 100.796
R283 drain_right.n2 drain_right.t6 52.3082
R284 drain_right.n20 drain_right.t0 52.3082
R285 drain_right.n8 drain_right.n6 48.5884
R286 drain_right.n25 drain_right.n24 48.0884
R287 drain_right drain_right.n12 22.1131
R288 drain_right.n9 drain_right.t2 9.9005
R289 drain_right.n9 drain_right.t3 9.9005
R290 drain_right.n10 drain_right.t9 9.9005
R291 drain_right.n10 drain_right.t7 9.9005
R292 drain_right.n7 drain_right.t11 9.9005
R293 drain_right.n7 drain_right.t8 9.9005
R294 drain_right.n13 drain_right.t12 9.9005
R295 drain_right.n13 drain_right.t4 9.9005
R296 drain_right.n14 drain_right.t13 9.9005
R297 drain_right.n14 drain_right.t5 9.9005
R298 drain_right.n16 drain_right.t10 9.9005
R299 drain_right.n16 drain_right.t1 9.9005
R300 drain_right.n3 drain_right.n1 9.71174
R301 drain_right.n21 drain_right.n19 9.71174
R302 drain_right.n6 drain_right.n5 9.45567
R303 drain_right.n24 drain_right.n23 9.45567
R304 drain_right.n5 drain_right.n4 9.3005
R305 drain_right.n23 drain_right.n22 9.3005
R306 drain_right.n6 drain_right.n0 8.14595
R307 drain_right.n24 drain_right.n18 8.14595
R308 drain_right.n4 drain_right.n3 7.3702
R309 drain_right.n22 drain_right.n21 7.3702
R310 drain_right drain_right.n25 5.90322
R311 drain_right.n4 drain_right.n0 5.81868
R312 drain_right.n22 drain_right.n18 5.81868
R313 drain_right.n5 drain_right.n1 3.44771
R314 drain_right.n23 drain_right.n19 3.44771
R315 drain_right.n25 drain_right.n17 0.5005
R316 drain_right.n17 drain_right.n15 0.5005
R317 drain_right.n12 drain_right.n8 0.320154
R318 drain_right.n12 drain_right.n11 0.070154
C0 source drain_right 7.22696f
C1 source drain_left 7.22975f
C2 drain_left drain_right 0.83691f
C3 plus minus 3.36217f
C4 minus source 1.30613f
C5 minus drain_right 1.15667f
C6 minus drain_left 0.177925f
C7 plus source 1.32021f
C8 plus drain_right 0.32016f
C9 plus drain_left 1.31449f
C10 drain_right a_n1644_n1288# 3.90951f
C11 drain_left a_n1644_n1288# 4.14758f
C12 source a_n1644_n1288# 2.519798f
C13 minus a_n1644_n1288# 5.588917f
C14 plus a_n1644_n1288# 6.244725f
C15 drain_right.n0 a_n1644_n1288# 0.038271f
C16 drain_right.n1 a_n1644_n1288# 0.084679f
C17 drain_right.t6 a_n1644_n1288# 0.063547f
C18 drain_right.n2 a_n1644_n1288# 0.066273f
C19 drain_right.n3 a_n1644_n1288# 0.021364f
C20 drain_right.n4 a_n1644_n1288# 0.01409f
C21 drain_right.n5 a_n1644_n1288# 0.186652f
C22 drain_right.n6 a_n1644_n1288# 0.061016f
C23 drain_right.t11 a_n1644_n1288# 0.041441f
C24 drain_right.t8 a_n1644_n1288# 0.041441f
C25 drain_right.n7 a_n1644_n1288# 0.260343f
C26 drain_right.n8 a_n1644_n1288# 0.362812f
C27 drain_right.t2 a_n1644_n1288# 0.041441f
C28 drain_right.t3 a_n1644_n1288# 0.041441f
C29 drain_right.n9 a_n1644_n1288# 0.261803f
C30 drain_right.t9 a_n1644_n1288# 0.041441f
C31 drain_right.t7 a_n1644_n1288# 0.041441f
C32 drain_right.n10 a_n1644_n1288# 0.260343f
C33 drain_right.n11 a_n1644_n1288# 0.551828f
C34 drain_right.n12 a_n1644_n1288# 0.636882f
C35 drain_right.t12 a_n1644_n1288# 0.041441f
C36 drain_right.t4 a_n1644_n1288# 0.041441f
C37 drain_right.n13 a_n1644_n1288# 0.261804f
C38 drain_right.t13 a_n1644_n1288# 0.041441f
C39 drain_right.t5 a_n1644_n1288# 0.041441f
C40 drain_right.n14 a_n1644_n1288# 0.260344f
C41 drain_right.n15 a_n1644_n1288# 0.579458f
C42 drain_right.t10 a_n1644_n1288# 0.041441f
C43 drain_right.t1 a_n1644_n1288# 0.041441f
C44 drain_right.n16 a_n1644_n1288# 0.260344f
C45 drain_right.n17 a_n1644_n1288# 0.285178f
C46 drain_right.n18 a_n1644_n1288# 0.038271f
C47 drain_right.n19 a_n1644_n1288# 0.084679f
C48 drain_right.t0 a_n1644_n1288# 0.063547f
C49 drain_right.n20 a_n1644_n1288# 0.066273f
C50 drain_right.n21 a_n1644_n1288# 0.021364f
C51 drain_right.n22 a_n1644_n1288# 0.01409f
C52 drain_right.n23 a_n1644_n1288# 0.186652f
C53 drain_right.n24 a_n1644_n1288# 0.06007f
C54 drain_right.n25 a_n1644_n1288# 0.307848f
C55 minus.n0 a_n1644_n1288# 0.030649f
C56 minus.t13 a_n1644_n1288# 0.048358f
C57 minus.t3 a_n1644_n1288# 0.045094f
C58 minus.t12 a_n1644_n1288# 0.045094f
C59 minus.t0 a_n1644_n1288# 0.045094f
C60 minus.n1 a_n1644_n1288# 0.043236f
C61 minus.n2 a_n1644_n1288# 0.065604f
C62 minus.t8 a_n1644_n1288# 0.045094f
C63 minus.t1 a_n1644_n1288# 0.045094f
C64 minus.t9 a_n1644_n1288# 0.048358f
C65 minus.n3 a_n1644_n1288# 0.041337f
C66 minus.n4 a_n1644_n1288# 0.033069f
C67 minus.n5 a_n1644_n1288# 0.011679f
C68 minus.n6 a_n1644_n1288# 0.033069f
C69 minus.n7 a_n1644_n1288# 0.011679f
C70 minus.n8 a_n1644_n1288# 0.030649f
C71 minus.n9 a_n1644_n1288# 0.030649f
C72 minus.n10 a_n1644_n1288# 0.030649f
C73 minus.n11 a_n1644_n1288# 0.011679f
C74 minus.n12 a_n1644_n1288# 0.033069f
C75 minus.n13 a_n1644_n1288# 0.011679f
C76 minus.n14 a_n1644_n1288# 0.033069f
C77 minus.n15 a_n1644_n1288# 0.041296f
C78 minus.n16 a_n1644_n1288# 0.693364f
C79 minus.n17 a_n1644_n1288# 0.030649f
C80 minus.t11 a_n1644_n1288# 0.045094f
C81 minus.t6 a_n1644_n1288# 0.045094f
C82 minus.t4 a_n1644_n1288# 0.045094f
C83 minus.n18 a_n1644_n1288# 0.043236f
C84 minus.n19 a_n1644_n1288# 0.065604f
C85 minus.t5 a_n1644_n1288# 0.045094f
C86 minus.t2 a_n1644_n1288# 0.045094f
C87 minus.t7 a_n1644_n1288# 0.048358f
C88 minus.n20 a_n1644_n1288# 0.041337f
C89 minus.n21 a_n1644_n1288# 0.033069f
C90 minus.n22 a_n1644_n1288# 0.011679f
C91 minus.n23 a_n1644_n1288# 0.033069f
C92 minus.n24 a_n1644_n1288# 0.011679f
C93 minus.n25 a_n1644_n1288# 0.030649f
C94 minus.n26 a_n1644_n1288# 0.030649f
C95 minus.n27 a_n1644_n1288# 0.030649f
C96 minus.n28 a_n1644_n1288# 0.011679f
C97 minus.n29 a_n1644_n1288# 0.033069f
C98 minus.n30 a_n1644_n1288# 0.011679f
C99 minus.n31 a_n1644_n1288# 0.033069f
C100 minus.t10 a_n1644_n1288# 0.048358f
C101 minus.n32 a_n1644_n1288# 0.041296f
C102 minus.n33 a_n1644_n1288# 0.196849f
C103 minus.n34 a_n1644_n1288# 0.859164f
C104 source.n0 a_n1644_n1288# 0.046178f
C105 source.n1 a_n1644_n1288# 0.102174f
C106 source.t21 a_n1644_n1288# 0.076676f
C107 source.n2 a_n1644_n1288# 0.079965f
C108 source.n3 a_n1644_n1288# 0.025778f
C109 source.n4 a_n1644_n1288# 0.017001f
C110 source.n5 a_n1644_n1288# 0.225216f
C111 source.n6 a_n1644_n1288# 0.050621f
C112 source.n7 a_n1644_n1288# 0.46987f
C113 source.t20 a_n1644_n1288# 0.050003f
C114 source.t15 a_n1644_n1288# 0.050003f
C115 source.n8 a_n1644_n1288# 0.267312f
C116 source.n9 a_n1644_n1288# 0.347915f
C117 source.t19 a_n1644_n1288# 0.050003f
C118 source.t27 a_n1644_n1288# 0.050003f
C119 source.n10 a_n1644_n1288# 0.267312f
C120 source.n11 a_n1644_n1288# 0.347915f
C121 source.t22 a_n1644_n1288# 0.050003f
C122 source.t26 a_n1644_n1288# 0.050003f
C123 source.n12 a_n1644_n1288# 0.267312f
C124 source.n13 a_n1644_n1288# 0.370326f
C125 source.n14 a_n1644_n1288# 0.046178f
C126 source.n15 a_n1644_n1288# 0.102174f
C127 source.t11 a_n1644_n1288# 0.076676f
C128 source.n16 a_n1644_n1288# 0.079965f
C129 source.n17 a_n1644_n1288# 0.025778f
C130 source.n18 a_n1644_n1288# 0.017001f
C131 source.n19 a_n1644_n1288# 0.225216f
C132 source.n20 a_n1644_n1288# 0.050621f
C133 source.n21 a_n1644_n1288# 0.150401f
C134 source.t9 a_n1644_n1288# 0.050003f
C135 source.t12 a_n1644_n1288# 0.050003f
C136 source.n22 a_n1644_n1288# 0.267312f
C137 source.n23 a_n1644_n1288# 0.347915f
C138 source.t3 a_n1644_n1288# 0.050003f
C139 source.t0 a_n1644_n1288# 0.050003f
C140 source.n24 a_n1644_n1288# 0.267312f
C141 source.n25 a_n1644_n1288# 0.347915f
C142 source.t5 a_n1644_n1288# 0.050003f
C143 source.t8 a_n1644_n1288# 0.050003f
C144 source.n26 a_n1644_n1288# 0.267312f
C145 source.n27 a_n1644_n1288# 1.03475f
C146 source.t14 a_n1644_n1288# 0.050003f
C147 source.t24 a_n1644_n1288# 0.050003f
C148 source.n28 a_n1644_n1288# 0.267311f
C149 source.n29 a_n1644_n1288# 1.03476f
C150 source.t17 a_n1644_n1288# 0.050003f
C151 source.t23 a_n1644_n1288# 0.050003f
C152 source.n30 a_n1644_n1288# 0.267311f
C153 source.n31 a_n1644_n1288# 0.347917f
C154 source.t25 a_n1644_n1288# 0.050003f
C155 source.t18 a_n1644_n1288# 0.050003f
C156 source.n32 a_n1644_n1288# 0.267311f
C157 source.n33 a_n1644_n1288# 0.347917f
C158 source.n34 a_n1644_n1288# 0.046178f
C159 source.n35 a_n1644_n1288# 0.102174f
C160 source.t16 a_n1644_n1288# 0.076676f
C161 source.n36 a_n1644_n1288# 0.079965f
C162 source.n37 a_n1644_n1288# 0.025778f
C163 source.n38 a_n1644_n1288# 0.017001f
C164 source.n39 a_n1644_n1288# 0.225216f
C165 source.n40 a_n1644_n1288# 0.050621f
C166 source.n41 a_n1644_n1288# 0.150401f
C167 source.t7 a_n1644_n1288# 0.050003f
C168 source.t2 a_n1644_n1288# 0.050003f
C169 source.n42 a_n1644_n1288# 0.267311f
C170 source.n43 a_n1644_n1288# 0.370327f
C171 source.t6 a_n1644_n1288# 0.050003f
C172 source.t10 a_n1644_n1288# 0.050003f
C173 source.n44 a_n1644_n1288# 0.267311f
C174 source.n45 a_n1644_n1288# 0.347917f
C175 source.t13 a_n1644_n1288# 0.050003f
C176 source.t1 a_n1644_n1288# 0.050003f
C177 source.n46 a_n1644_n1288# 0.267311f
C178 source.n47 a_n1644_n1288# 0.347917f
C179 source.n48 a_n1644_n1288# 0.046178f
C180 source.n49 a_n1644_n1288# 0.102174f
C181 source.t4 a_n1644_n1288# 0.076676f
C182 source.n50 a_n1644_n1288# 0.079965f
C183 source.n51 a_n1644_n1288# 0.025778f
C184 source.n52 a_n1644_n1288# 0.017001f
C185 source.n53 a_n1644_n1288# 0.225216f
C186 source.n54 a_n1644_n1288# 0.050621f
C187 source.n55 a_n1644_n1288# 0.299993f
C188 source.n56 a_n1644_n1288# 0.780352f
C189 drain_left.n0 a_n1644_n1288# 0.037733f
C190 drain_left.n1 a_n1644_n1288# 0.083489f
C191 drain_left.t12 a_n1644_n1288# 0.062654f
C192 drain_left.n2 a_n1644_n1288# 0.065342f
C193 drain_left.n3 a_n1644_n1288# 0.021064f
C194 drain_left.n4 a_n1644_n1288# 0.013892f
C195 drain_left.n5 a_n1644_n1288# 0.184031f
C196 drain_left.n6 a_n1644_n1288# 0.060159f
C197 drain_left.t0 a_n1644_n1288# 0.040859f
C198 drain_left.t8 a_n1644_n1288# 0.040859f
C199 drain_left.n7 a_n1644_n1288# 0.256686f
C200 drain_left.n8 a_n1644_n1288# 0.357716f
C201 drain_left.t10 a_n1644_n1288# 0.040859f
C202 drain_left.t13 a_n1644_n1288# 0.040859f
C203 drain_left.n9 a_n1644_n1288# 0.258126f
C204 drain_left.t6 a_n1644_n1288# 0.040859f
C205 drain_left.t2 a_n1644_n1288# 0.040859f
C206 drain_left.n10 a_n1644_n1288# 0.256686f
C207 drain_left.n11 a_n1644_n1288# 0.544077f
C208 drain_left.n12 a_n1644_n1288# 0.678682f
C209 drain_left.n13 a_n1644_n1288# 0.037733f
C210 drain_left.n14 a_n1644_n1288# 0.083489f
C211 drain_left.t3 a_n1644_n1288# 0.062654f
C212 drain_left.n15 a_n1644_n1288# 0.065342f
C213 drain_left.n16 a_n1644_n1288# 0.021064f
C214 drain_left.n17 a_n1644_n1288# 0.013892f
C215 drain_left.n18 a_n1644_n1288# 0.184031f
C216 drain_left.n19 a_n1644_n1288# 0.060159f
C217 drain_left.t5 a_n1644_n1288# 0.040859f
C218 drain_left.t9 a_n1644_n1288# 0.040859f
C219 drain_left.n20 a_n1644_n1288# 0.256687f
C220 drain_left.n21 a_n1644_n1288# 0.370863f
C221 drain_left.t4 a_n1644_n1288# 0.040859f
C222 drain_left.t7 a_n1644_n1288# 0.040859f
C223 drain_left.n22 a_n1644_n1288# 0.256687f
C224 drain_left.n23 a_n1644_n1288# 0.281172f
C225 drain_left.t11 a_n1644_n1288# 0.040859f
C226 drain_left.t1 a_n1644_n1288# 0.040859f
C227 drain_left.n24 a_n1644_n1288# 0.256687f
C228 drain_left.n25 a_n1644_n1288# 0.494566f
C229 plus.n0 a_n1644_n1288# 0.031218f
C230 plus.t12 a_n1644_n1288# 0.045931f
C231 plus.t7 a_n1644_n1288# 0.045931f
C232 plus.t0 a_n1644_n1288# 0.045931f
C233 plus.n1 a_n1644_n1288# 0.044039f
C234 plus.n2 a_n1644_n1288# 0.066822f
C235 plus.t8 a_n1644_n1288# 0.045931f
C236 plus.t1 a_n1644_n1288# 0.045931f
C237 plus.t5 a_n1644_n1288# 0.049256f
C238 plus.n3 a_n1644_n1288# 0.042104f
C239 plus.n4 a_n1644_n1288# 0.033683f
C240 plus.n5 a_n1644_n1288# 0.011896f
C241 plus.n6 a_n1644_n1288# 0.033683f
C242 plus.n7 a_n1644_n1288# 0.011896f
C243 plus.n8 a_n1644_n1288# 0.031218f
C244 plus.n9 a_n1644_n1288# 0.031218f
C245 plus.n10 a_n1644_n1288# 0.031218f
C246 plus.n11 a_n1644_n1288# 0.011896f
C247 plus.n12 a_n1644_n1288# 0.033683f
C248 plus.n13 a_n1644_n1288# 0.011896f
C249 plus.n14 a_n1644_n1288# 0.033683f
C250 plus.t6 a_n1644_n1288# 0.049256f
C251 plus.n15 a_n1644_n1288# 0.042062f
C252 plus.n16 a_n1644_n1288# 0.219392f
C253 plus.n17 a_n1644_n1288# 0.031218f
C254 plus.t13 a_n1644_n1288# 0.049256f
C255 plus.t3 a_n1644_n1288# 0.045931f
C256 plus.t10 a_n1644_n1288# 0.045931f
C257 plus.t4 a_n1644_n1288# 0.045931f
C258 plus.n18 a_n1644_n1288# 0.044039f
C259 plus.n19 a_n1644_n1288# 0.066822f
C260 plus.t2 a_n1644_n1288# 0.045931f
C261 plus.t9 a_n1644_n1288# 0.045931f
C262 plus.t11 a_n1644_n1288# 0.049256f
C263 plus.n20 a_n1644_n1288# 0.042104f
C264 plus.n21 a_n1644_n1288# 0.033683f
C265 plus.n22 a_n1644_n1288# 0.011896f
C266 plus.n23 a_n1644_n1288# 0.033683f
C267 plus.n24 a_n1644_n1288# 0.011896f
C268 plus.n25 a_n1644_n1288# 0.031218f
C269 plus.n26 a_n1644_n1288# 0.031218f
C270 plus.n27 a_n1644_n1288# 0.031218f
C271 plus.n28 a_n1644_n1288# 0.011896f
C272 plus.n29 a_n1644_n1288# 0.033683f
C273 plus.n30 a_n1644_n1288# 0.011896f
C274 plus.n31 a_n1644_n1288# 0.033683f
C275 plus.n32 a_n1644_n1288# 0.042062f
C276 plus.n33 a_n1644_n1288# 0.675482f
.ends

