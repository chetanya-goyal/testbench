* NGSPICE file created from diffpair363.ext - technology: sky130A

.subckt diffpair363 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t7 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 source.t1 minus.t0 drain_right.t7 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 source.t8 plus.t1 drain_left.t6 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X3 drain_right.t6 minus.t1 source.t2 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X4 a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X5 drain_right.t5 minus.t2 source.t3 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 source.t0 minus.t3 drain_right.t4 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X7 drain_left.t5 plus.t2 source.t9 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X8 a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X9 drain_right.t3 minus.t4 source.t15 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X10 drain_left.t4 plus.t3 source.t10 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 drain_left.t3 plus.t4 source.t13 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X12 source.t11 plus.t5 drain_left.t2 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 source.t4 minus.t5 drain_right.t2 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X14 source.t14 plus.t6 drain_left.t1 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X15 a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X16 source.t12 plus.t7 drain_left.t0 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 drain_right.t1 minus.t6 source.t6 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 source.t5 minus.t7 drain_right.t0 a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X19 a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# a_n1546_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 plus.n2 plus.t1 533.348
R1 plus.n10 plus.t4 533.348
R2 plus.n6 plus.t2 512.366
R3 plus.n5 plus.t7 512.366
R4 plus.n1 plus.t3 512.366
R5 plus.n14 plus.t6 512.366
R6 plus.n13 plus.t0 512.366
R7 plus.n9 plus.t5 512.366
R8 plus.n4 plus.n3 161.3
R9 plus.n5 plus.n0 161.3
R10 plus.n7 plus.n6 161.3
R11 plus.n12 plus.n11 161.3
R12 plus.n13 plus.n8 161.3
R13 plus.n15 plus.n14 161.3
R14 plus.n3 plus.n2 70.4033
R15 plus.n11 plus.n10 70.4033
R16 plus.n6 plus.n5 48.2005
R17 plus.n14 plus.n13 48.2005
R18 plus plus.n15 27.8172
R19 plus.n4 plus.n1 24.1005
R20 plus.n5 plus.n4 24.1005
R21 plus.n13 plus.n12 24.1005
R22 plus.n12 plus.n9 24.1005
R23 plus.n2 plus.n1 20.9576
R24 plus.n10 plus.n9 20.9576
R25 plus plus.n7 11.1028
R26 plus.n3 plus.n0 0.189894
R27 plus.n7 plus.n0 0.189894
R28 plus.n15 plus.n8 0.189894
R29 plus.n11 plus.n8 0.189894
R30 source.n3 source.t8 51.0588
R31 source.n4 source.t15 51.0588
R32 source.n7 source.t4 51.0588
R33 source.n15 source.t2 51.0586
R34 source.n12 source.t5 51.0586
R35 source.n11 source.t13 51.0586
R36 source.n8 source.t14 51.0586
R37 source.n0 source.t9 51.0586
R38 source.n2 source.n1 48.8588
R39 source.n6 source.n5 48.8588
R40 source.n14 source.n13 48.8586
R41 source.n10 source.n9 48.8586
R42 source.n8 source.n7 19.7305
R43 source.n16 source.n0 14.1098
R44 source.n16 source.n15 5.62119
R45 source.n13 source.t6 2.2005
R46 source.n13 source.t0 2.2005
R47 source.n9 source.t7 2.2005
R48 source.n9 source.t11 2.2005
R49 source.n1 source.t10 2.2005
R50 source.n1 source.t12 2.2005
R51 source.n5 source.t3 2.2005
R52 source.n5 source.t1 2.2005
R53 source.n7 source.n6 0.716017
R54 source.n6 source.n4 0.716017
R55 source.n3 source.n2 0.716017
R56 source.n2 source.n0 0.716017
R57 source.n10 source.n8 0.716017
R58 source.n11 source.n10 0.716017
R59 source.n14 source.n12 0.716017
R60 source.n15 source.n14 0.716017
R61 source.n4 source.n3 0.470328
R62 source.n12 source.n11 0.470328
R63 source source.n16 0.188
R64 drain_left.n5 drain_left.n3 66.2531
R65 drain_left.n2 drain_left.n1 65.8397
R66 drain_left.n2 drain_left.n0 65.8397
R67 drain_left.n5 drain_left.n4 65.5374
R68 drain_left drain_left.n2 27.5987
R69 drain_left drain_left.n5 6.36873
R70 drain_left.n1 drain_left.t2 2.2005
R71 drain_left.n1 drain_left.t3 2.2005
R72 drain_left.n0 drain_left.t1 2.2005
R73 drain_left.n0 drain_left.t7 2.2005
R74 drain_left.n4 drain_left.t0 2.2005
R75 drain_left.n4 drain_left.t5 2.2005
R76 drain_left.n3 drain_left.t6 2.2005
R77 drain_left.n3 drain_left.t4 2.2005
R78 minus.n2 minus.t4 533.348
R79 minus.n10 minus.t7 533.348
R80 minus.n1 minus.t0 512.366
R81 minus.n5 minus.t2 512.366
R82 minus.n6 minus.t5 512.366
R83 minus.n9 minus.t6 512.366
R84 minus.n13 minus.t3 512.366
R85 minus.n14 minus.t1 512.366
R86 minus.n7 minus.n6 161.3
R87 minus.n5 minus.n0 161.3
R88 minus.n4 minus.n3 161.3
R89 minus.n15 minus.n14 161.3
R90 minus.n13 minus.n8 161.3
R91 minus.n12 minus.n11 161.3
R92 minus.n3 minus.n2 70.4033
R93 minus.n11 minus.n10 70.4033
R94 minus.n6 minus.n5 48.2005
R95 minus.n14 minus.n13 48.2005
R96 minus.n16 minus.n7 32.7997
R97 minus.n5 minus.n4 24.1005
R98 minus.n4 minus.n1 24.1005
R99 minus.n12 minus.n9 24.1005
R100 minus.n13 minus.n12 24.1005
R101 minus.n2 minus.n1 20.9576
R102 minus.n10 minus.n9 20.9576
R103 minus.n16 minus.n15 6.5952
R104 minus.n7 minus.n0 0.189894
R105 minus.n3 minus.n0 0.189894
R106 minus.n11 minus.n8 0.189894
R107 minus.n15 minus.n8 0.189894
R108 minus minus.n16 0.188
R109 drain_right.n5 drain_right.n3 66.2529
R110 drain_right.n2 drain_right.n1 65.8397
R111 drain_right.n2 drain_right.n0 65.8397
R112 drain_right.n5 drain_right.n4 65.5376
R113 drain_right drain_right.n2 27.0454
R114 drain_right drain_right.n5 6.36873
R115 drain_right.n1 drain_right.t4 2.2005
R116 drain_right.n1 drain_right.t6 2.2005
R117 drain_right.n0 drain_right.t0 2.2005
R118 drain_right.n0 drain_right.t1 2.2005
R119 drain_right.n3 drain_right.t7 2.2005
R120 drain_right.n3 drain_right.t3 2.2005
R121 drain_right.n4 drain_right.t2 2.2005
R122 drain_right.n4 drain_right.t5 2.2005
C0 drain_right plus 0.302201f
C1 source drain_right 10.3145f
C2 source plus 3.3423f
C3 minus drain_left 0.171215f
C4 drain_right drain_left 0.727126f
C5 drain_left plus 3.67827f
C6 source drain_left 10.314f
C7 minus drain_right 3.53025f
C8 minus plus 4.51612f
C9 source minus 3.32826f
C10 drain_right a_n1546_n2688# 5.00728f
C11 drain_left a_n1546_n2688# 5.252691f
C12 source a_n1546_n2688# 7.082566f
C13 minus a_n1546_n2688# 5.758883f
C14 plus a_n1546_n2688# 7.40293f
C15 drain_right.t0 a_n1546_n2688# 0.203389f
C16 drain_right.t1 a_n1546_n2688# 0.203389f
C17 drain_right.n0 a_n1546_n2688# 1.78052f
C18 drain_right.t4 a_n1546_n2688# 0.203389f
C19 drain_right.t6 a_n1546_n2688# 0.203389f
C20 drain_right.n1 a_n1546_n2688# 1.78052f
C21 drain_right.n2 a_n1546_n2688# 1.74345f
C22 drain_right.t7 a_n1546_n2688# 0.203389f
C23 drain_right.t3 a_n1546_n2688# 0.203389f
C24 drain_right.n3 a_n1546_n2688# 1.78299f
C25 drain_right.t2 a_n1546_n2688# 0.203389f
C26 drain_right.t5 a_n1546_n2688# 0.203389f
C27 drain_right.n4 a_n1546_n2688# 1.77898f
C28 drain_right.n5 a_n1546_n2688# 0.975067f
C29 minus.n0 a_n1546_n2688# 0.048826f
C30 minus.t0 a_n1546_n2688# 0.630113f
C31 minus.n1 a_n1546_n2688# 0.27352f
C32 minus.t4 a_n1546_n2688# 0.640681f
C33 minus.n2 a_n1546_n2688# 0.258362f
C34 minus.n3 a_n1546_n2688# 0.160851f
C35 minus.n4 a_n1546_n2688# 0.01108f
C36 minus.t2 a_n1546_n2688# 0.630113f
C37 minus.n5 a_n1546_n2688# 0.27352f
C38 minus.t5 a_n1546_n2688# 0.630113f
C39 minus.n6 a_n1546_n2688# 0.268552f
C40 minus.n7 a_n1546_n2688# 1.47824f
C41 minus.n8 a_n1546_n2688# 0.048826f
C42 minus.t6 a_n1546_n2688# 0.630113f
C43 minus.n9 a_n1546_n2688# 0.27352f
C44 minus.t7 a_n1546_n2688# 0.640681f
C45 minus.n10 a_n1546_n2688# 0.258362f
C46 minus.n11 a_n1546_n2688# 0.160851f
C47 minus.n12 a_n1546_n2688# 0.01108f
C48 minus.t3 a_n1546_n2688# 0.630113f
C49 minus.n13 a_n1546_n2688# 0.27352f
C50 minus.t1 a_n1546_n2688# 0.630113f
C51 minus.n14 a_n1546_n2688# 0.268552f
C52 minus.n15 a_n1546_n2688# 0.330111f
C53 minus.n16 a_n1546_n2688# 1.80813f
C54 drain_left.t1 a_n1546_n2688# 0.204678f
C55 drain_left.t7 a_n1546_n2688# 0.204678f
C56 drain_left.n0 a_n1546_n2688# 1.7918f
C57 drain_left.t2 a_n1546_n2688# 0.204678f
C58 drain_left.t3 a_n1546_n2688# 0.204678f
C59 drain_left.n1 a_n1546_n2688# 1.7918f
C60 drain_left.n2 a_n1546_n2688# 1.81407f
C61 drain_left.t6 a_n1546_n2688# 0.204678f
C62 drain_left.t4 a_n1546_n2688# 0.204678f
C63 drain_left.n3 a_n1546_n2688# 1.7943f
C64 drain_left.t0 a_n1546_n2688# 0.204678f
C65 drain_left.t5 a_n1546_n2688# 0.204678f
C66 drain_left.n4 a_n1546_n2688# 1.79024f
C67 drain_left.n5 a_n1546_n2688# 0.981244f
C68 source.t9 a_n1546_n2688# 1.6348f
C69 source.n0 a_n1546_n2688# 0.960092f
C70 source.t10 a_n1546_n2688# 0.153309f
C71 source.t12 a_n1546_n2688# 0.153309f
C72 source.n1 a_n1546_n2688# 1.2834f
C73 source.n2 a_n1546_n2688# 0.300304f
C74 source.t8 a_n1546_n2688# 1.63481f
C75 source.n3 a_n1546_n2688# 0.349948f
C76 source.t15 a_n1546_n2688# 1.63481f
C77 source.n4 a_n1546_n2688# 0.349948f
C78 source.t3 a_n1546_n2688# 0.153309f
C79 source.t1 a_n1546_n2688# 0.153309f
C80 source.n5 a_n1546_n2688# 1.2834f
C81 source.n6 a_n1546_n2688# 0.300304f
C82 source.t4 a_n1546_n2688# 1.63481f
C83 source.n7 a_n1546_n2688# 1.27721f
C84 source.t14 a_n1546_n2688# 1.6348f
C85 source.n8 a_n1546_n2688# 1.27722f
C86 source.t7 a_n1546_n2688# 0.153309f
C87 source.t11 a_n1546_n2688# 0.153309f
C88 source.n9 a_n1546_n2688# 1.2834f
C89 source.n10 a_n1546_n2688# 0.300308f
C90 source.t13 a_n1546_n2688# 1.6348f
C91 source.n11 a_n1546_n2688# 0.349952f
C92 source.t5 a_n1546_n2688# 1.6348f
C93 source.n12 a_n1546_n2688# 0.349952f
C94 source.t6 a_n1546_n2688# 0.153309f
C95 source.t0 a_n1546_n2688# 0.153309f
C96 source.n13 a_n1546_n2688# 1.2834f
C97 source.n14 a_n1546_n2688# 0.300308f
C98 source.t2 a_n1546_n2688# 1.6348f
C99 source.n15 a_n1546_n2688# 0.481153f
C100 source.n16 a_n1546_n2688# 1.12852f
C101 plus.n0 a_n1546_n2688# 0.050128f
C102 plus.t2 a_n1546_n2688# 0.646918f
C103 plus.t7 a_n1546_n2688# 0.646918f
C104 plus.t3 a_n1546_n2688# 0.646918f
C105 plus.n1 a_n1546_n2688# 0.280814f
C106 plus.t1 a_n1546_n2688# 0.657768f
C107 plus.n2 a_n1546_n2688# 0.265252f
C108 plus.n3 a_n1546_n2688# 0.165141f
C109 plus.n4 a_n1546_n2688# 0.011375f
C110 plus.n5 a_n1546_n2688# 0.280814f
C111 plus.n6 a_n1546_n2688# 0.275715f
C112 plus.n7 a_n1546_n2688# 0.503948f
C113 plus.n8 a_n1546_n2688# 0.050128f
C114 plus.t6 a_n1546_n2688# 0.646918f
C115 plus.t0 a_n1546_n2688# 0.646918f
C116 plus.t5 a_n1546_n2688# 0.646918f
C117 plus.n9 a_n1546_n2688# 0.280814f
C118 plus.t4 a_n1546_n2688# 0.657768f
C119 plus.n10 a_n1546_n2688# 0.265252f
C120 plus.n11 a_n1546_n2688# 0.165141f
C121 plus.n12 a_n1546_n2688# 0.011375f
C122 plus.n13 a_n1546_n2688# 0.280814f
C123 plus.n14 a_n1546_n2688# 0.275715f
C124 plus.n15 a_n1546_n2688# 1.32347f
.ends

