* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t11 plus.t0 drain_left.t4 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 drain_right.t5 minus.t0 source.t3 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X2 source.t2 minus.t1 drain_right.t4 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 drain_right.t3 minus.t2 source.t0 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X4 drain_left.t1 plus.t1 source.t10 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X5 a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X6 source.t9 plus.t2 drain_left.t0 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X7 drain_left.t5 plus.t3 source.t8 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X8 a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X9 drain_left.t3 plus.t4 source.t7 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X10 drain_right.t2 minus.t3 source.t5 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X11 drain_right.t1 minus.t4 source.t1 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X12 drain_left.t2 plus.t5 source.t6 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X13 a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X14 source.t4 minus.t5 drain_right.t0 a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X15 a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# a_n1180_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
R0 plus.n0 plus.t1 269.921
R1 plus.n2 plus.t3 269.921
R2 plus.n4 plus.t4 269.921
R3 plus.n6 plus.t5 269.921
R4 plus.n1 plus.t0 221.72
R5 plus.n5 plus.t2 221.72
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 23.2907
R15 plus plus.n3 7.96262
R16 drain_left.n3 drain_left.t1 260.433
R17 drain_left.n1 drain_left.t2 260.252
R18 drain_left.n1 drain_left.n0 240.202
R19 drain_left.n3 drain_left.n2 240.132
R20 drain_left drain_left.n1 20.4087
R21 drain_left.n0 drain_left.t0 19.8005
R22 drain_left.n0 drain_left.t3 19.8005
R23 drain_left.n2 drain_left.t4 19.8005
R24 drain_left.n2 drain_left.t5 19.8005
R25 drain_left drain_left.n3 6.15322
R26 source.n0 source.t8 243.255
R27 source.n3 source.t1 243.255
R28 source.n11 source.t3 243.254
R29 source.n8 source.t7 243.254
R30 source.n2 source.n1 223.454
R31 source.n5 source.n4 223.454
R32 source.n10 source.n9 223.453
R33 source.n7 source.n6 223.453
R34 source.n9 source.t0 19.8005
R35 source.n9 source.t4 19.8005
R36 source.n6 source.t6 19.8005
R37 source.n6 source.t9 19.8005
R38 source.n1 source.t10 19.8005
R39 source.n1 source.t11 19.8005
R40 source.n4 source.t5 19.8005
R41 source.n4 source.t2 19.8005
R42 source.n7 source.n5 13.9544
R43 source.n12 source.n0 7.94146
R44 source.n12 source.n11 5.51343
R45 source.n3 source.n2 0.720328
R46 source.n10 source.n8 0.720328
R47 source.n5 source.n3 0.5005
R48 source.n2 source.n0 0.5005
R49 source.n8 source.n7 0.5005
R50 source.n11 source.n10 0.5005
R51 source source.n12 0.188
R52 minus.n2 minus.t3 269.921
R53 minus.n0 minus.t4 269.921
R54 minus.n6 minus.t0 269.921
R55 minus.n4 minus.t2 269.921
R56 minus.n1 minus.t1 221.72
R57 minus.n5 minus.t5 221.72
R58 minus.n3 minus.n0 161.489
R59 minus.n7 minus.n4 161.489
R60 minus.n3 minus.n2 161.3
R61 minus.n7 minus.n6 161.3
R62 minus.n2 minus.n1 36.5157
R63 minus.n1 minus.n0 36.5157
R64 minus.n5 minus.n4 36.5157
R65 minus.n6 minus.n5 36.5157
R66 minus.n8 minus.n3 25.2429
R67 minus.n8 minus.n7 6.48535
R68 minus minus.n8 0.188
R69 drain_right.n1 drain_right.t3 260.252
R70 drain_right.n3 drain_right.t2 259.933
R71 drain_right.n3 drain_right.n2 240.632
R72 drain_right.n1 drain_right.n0 240.202
R73 drain_right drain_right.n1 19.8555
R74 drain_right.n0 drain_right.t0 19.8005
R75 drain_right.n0 drain_right.t5 19.8005
R76 drain_right.n2 drain_right.t4 19.8005
R77 drain_right.n2 drain_right.t1 19.8005
R78 drain_right drain_right.n3 5.90322
C0 source drain_right 2.74272f
C1 minus drain_right 0.489067f
C2 minus source 0.60138f
C3 drain_left plus 0.598799f
C4 drain_left drain_right 0.547385f
C5 drain_left source 2.74581f
C6 drain_right plus 0.272027f
C7 minus drain_left 0.178167f
C8 source plus 0.6153f
C9 minus plus 2.59426f
C10 drain_right a_n1180_n1088# 2.718115f
C11 drain_left a_n1180_n1088# 2.862884f
C12 source a_n1180_n1088# 1.897006f
C13 minus a_n1180_n1088# 3.624647f
C14 plus a_n1180_n1088# 4.384402f
C15 drain_right.t3 a_n1180_n1088# 0.10565f
C16 drain_right.t0 a_n1180_n1088# 0.017043f
C17 drain_right.t5 a_n1180_n1088# 0.017043f
C18 drain_right.n0 a_n1180_n1088# 0.066283f
C19 drain_right.n1 a_n1180_n1088# 0.790257f
C20 drain_right.t4 a_n1180_n1088# 0.017043f
C21 drain_right.t1 a_n1180_n1088# 0.017043f
C22 drain_right.n2 a_n1180_n1088# 0.066699f
C23 drain_right.t2 a_n1180_n1088# 0.105416f
C24 drain_right.n3 a_n1180_n1088# 0.607669f
C25 minus.t4 a_n1180_n1088# 0.037982f
C26 minus.n0 a_n1180_n1088# 0.045617f
C27 minus.t3 a_n1180_n1088# 0.037982f
C28 minus.t1 a_n1180_n1088# 0.03146f
C29 minus.n1 a_n1180_n1088# 0.034511f
C30 minus.n2 a_n1180_n1088# 0.045557f
C31 minus.n3 a_n1180_n1088# 0.830201f
C32 minus.t2 a_n1180_n1088# 0.037982f
C33 minus.n4 a_n1180_n1088# 0.045617f
C34 minus.t5 a_n1180_n1088# 0.03146f
C35 minus.n5 a_n1180_n1088# 0.034511f
C36 minus.t0 a_n1180_n1088# 0.037982f
C37 minus.n6 a_n1180_n1088# 0.045557f
C38 minus.n7 a_n1180_n1088# 0.316551f
C39 minus.n8 a_n1180_n1088# 0.960218f
C40 source.t8 a_n1180_n1088# 0.127312f
C41 source.n0 a_n1180_n1088# 0.539452f
C42 source.t10 a_n1180_n1088# 0.022874f
C43 source.t11 a_n1180_n1088# 0.022874f
C44 source.n1 a_n1180_n1088# 0.074184f
C45 source.n2 a_n1180_n1088# 0.291548f
C46 source.t1 a_n1180_n1088# 0.127312f
C47 source.n3 a_n1180_n1088# 0.300803f
C48 source.t5 a_n1180_n1088# 0.022874f
C49 source.t2 a_n1180_n1088# 0.022874f
C50 source.n4 a_n1180_n1088# 0.074184f
C51 source.n5 a_n1180_n1088# 0.807943f
C52 source.t6 a_n1180_n1088# 0.022874f
C53 source.t9 a_n1180_n1088# 0.022874f
C54 source.n6 a_n1180_n1088# 0.074183f
C55 source.n7 a_n1180_n1088# 0.807943f
C56 source.t7 a_n1180_n1088# 0.127312f
C57 source.n8 a_n1180_n1088# 0.300803f
C58 source.t0 a_n1180_n1088# 0.022874f
C59 source.t4 a_n1180_n1088# 0.022874f
C60 source.n9 a_n1180_n1088# 0.074183f
C61 source.n10 a_n1180_n1088# 0.291548f
C62 source.t3 a_n1180_n1088# 0.127312f
C63 source.n11 a_n1180_n1088# 0.437666f
C64 source.n12 a_n1180_n1088# 0.584594f
C65 drain_left.t2 a_n1180_n1088# 0.102449f
C66 drain_left.t0 a_n1180_n1088# 0.016526f
C67 drain_left.t3 a_n1180_n1088# 0.016526f
C68 drain_left.n0 a_n1180_n1088# 0.064274f
C69 drain_left.n1 a_n1180_n1088# 0.806906f
C70 drain_left.t1 a_n1180_n1088# 0.102597f
C71 drain_left.t4 a_n1180_n1088# 0.016526f
C72 drain_left.t5 a_n1180_n1088# 0.016526f
C73 drain_left.n2 a_n1180_n1088# 0.064216f
C74 drain_left.n3 a_n1180_n1088# 0.581318f
C75 plus.t1 a_n1180_n1088# 0.039228f
C76 plus.n0 a_n1180_n1088# 0.047113f
C77 plus.t0 a_n1180_n1088# 0.032492f
C78 plus.n1 a_n1180_n1088# 0.035643f
C79 plus.t3 a_n1180_n1088# 0.039228f
C80 plus.n2 a_n1180_n1088# 0.047051f
C81 plus.n3 a_n1180_n1088# 0.340271f
C82 plus.t4 a_n1180_n1088# 0.039228f
C83 plus.n4 a_n1180_n1088# 0.047113f
C84 plus.t5 a_n1180_n1088# 0.039228f
C85 plus.t2 a_n1180_n1088# 0.032492f
C86 plus.n5 a_n1180_n1088# 0.035643f
C87 plus.n6 a_n1180_n1088# 0.047051f
C88 plus.n7 a_n1180_n1088# 0.841537f
.ends

