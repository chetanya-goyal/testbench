* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 drain_right.t9 minus.t0 source.t14 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X3 drain_left.t9 plus.t0 source.t7 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X4 a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X5 a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X6 drain_right.t8 minus.t1 source.t12 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X7 drain_right.t7 minus.t2 source.t19 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_right.t6 minus.t3 source.t18 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X9 drain_left.t8 plus.t1 source.t1 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X10 drain_left.t7 plus.t2 source.t5 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X11 source.t17 minus.t4 drain_right.t5 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X12 drain_right.t4 minus.t5 source.t16 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X13 source.t13 minus.t6 drain_right.t3 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X14 drain_right.t2 minus.t7 source.t15 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X15 source.t6 plus.t3 drain_left.t6 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X16 source.t11 minus.t8 drain_right.t1 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X17 source.t10 minus.t9 drain_right.t0 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_left.t5 plus.t4 source.t0 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X19 drain_left.t4 plus.t5 source.t2 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X20 source.t9 plus.t6 drain_left.t3 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 source.t8 plus.t7 drain_left.t2 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 drain_left.t1 plus.t8 source.t4 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X23 source.t3 plus.t9 drain_left.t0 a_n2072_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n9 minus.n8 161.3
R1 minus.n7 minus.n0 161.3
R2 minus.n19 minus.n18 161.3
R3 minus.n17 minus.n10 161.3
R4 minus.n3 minus.t5 102.425
R5 minus.n13 minus.t2 102.425
R6 minus.n6 minus.n5 80.6037
R7 minus.n4 minus.n1 80.6037
R8 minus.n16 minus.n15 80.6037
R9 minus.n14 minus.n11 80.6037
R10 minus.n2 minus.t4 79.2293
R11 minus.n1 minus.t3 79.2293
R12 minus.n6 minus.t6 79.2293
R13 minus.n8 minus.t7 79.2293
R14 minus.n12 minus.t9 79.2293
R15 minus.n11 minus.t1 79.2293
R16 minus.n16 minus.t8 79.2293
R17 minus.n18 minus.t0 79.2293
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n7 minus.n6 32.1338
R23 minus.n17 minus.n16 32.1338
R24 minus.n4 minus.n3 31.8629
R25 minus.n14 minus.n13 31.8629
R26 minus.n20 minus.n9 28.813
R27 minus.n3 minus.n2 16.2333
R28 minus.n13 minus.n12 16.2333
R29 minus.n8 minus.n7 16.0672
R30 minus.n18 minus.n17 16.0672
R31 minus.n20 minus.n19 6.67664
R32 minus.n5 minus.n4 0.380177
R33 minus.n15 minus.n14 0.380177
R34 minus.n5 minus.n0 0.285035
R35 minus.n15 minus.n10 0.285035
R36 minus.n9 minus.n0 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 source.n0 source.t2 243.255
R40 source.n5 source.t16 243.255
R41 source.n19 source.t14 243.254
R42 source.n14 source.t1 243.254
R43 source.n2 source.n1 223.454
R44 source.n4 source.n3 223.454
R45 source.n7 source.n6 223.454
R46 source.n9 source.n8 223.454
R47 source.n18 source.n17 223.453
R48 source.n16 source.n15 223.453
R49 source.n13 source.n12 223.453
R50 source.n11 source.n10 223.453
R51 source.n17 source.t12 19.8005
R52 source.n17 source.t11 19.8005
R53 source.n15 source.t19 19.8005
R54 source.n15 source.t10 19.8005
R55 source.n12 source.t5 19.8005
R56 source.n12 source.t8 19.8005
R57 source.n10 source.t7 19.8005
R58 source.n10 source.t3 19.8005
R59 source.n1 source.t0 19.8005
R60 source.n1 source.t6 19.8005
R61 source.n3 source.t4 19.8005
R62 source.n3 source.t9 19.8005
R63 source.n6 source.t18 19.8005
R64 source.n6 source.t17 19.8005
R65 source.n8 source.t15 19.8005
R66 source.n8 source.t13 19.8005
R67 source.n11 source.n9 14.9027
R68 source.n20 source.n0 8.17853
R69 source.n20 source.n19 5.7505
R70 source.n9 source.n7 0.974638
R71 source.n7 source.n5 0.974638
R72 source.n4 source.n2 0.974638
R73 source.n2 source.n0 0.974638
R74 source.n13 source.n11 0.974638
R75 source.n14 source.n13 0.974638
R76 source.n18 source.n16 0.974638
R77 source.n19 source.n18 0.974638
R78 source.n5 source.n4 0.957397
R79 source.n16 source.n14 0.957397
R80 source source.n20 0.188
R81 drain_right.n1 drain_right.t7 260.906
R82 drain_right.n7 drain_right.t2 259.933
R83 drain_right.n6 drain_right.n4 241.107
R84 drain_right.n3 drain_right.n2 240.808
R85 drain_right.n6 drain_right.n5 240.132
R86 drain_right.n1 drain_right.n0 240.131
R87 drain_right drain_right.n3 22.6206
R88 drain_right.n2 drain_right.t1 19.8005
R89 drain_right.n2 drain_right.t9 19.8005
R90 drain_right.n0 drain_right.t0 19.8005
R91 drain_right.n0 drain_right.t8 19.8005
R92 drain_right.n4 drain_right.t5 19.8005
R93 drain_right.n4 drain_right.t4 19.8005
R94 drain_right.n5 drain_right.t3 19.8005
R95 drain_right.n5 drain_right.t6 19.8005
R96 drain_right drain_right.n7 6.14028
R97 drain_right.n7 drain_right.n6 0.974638
R98 drain_right.n3 drain_right.n1 0.188688
R99 plus.n7 plus.n0 161.3
R100 plus.n9 plus.n8 161.3
R101 plus.n17 plus.n10 161.3
R102 plus.n19 plus.n18 161.3
R103 plus.n3 plus.t8 102.425
R104 plus.n13 plus.t1 102.425
R105 plus.n5 plus.n2 80.6037
R106 plus.n6 plus.n1 80.6037
R107 plus.n15 plus.n12 80.6037
R108 plus.n16 plus.n11 80.6037
R109 plus.n8 plus.t5 79.2293
R110 plus.n6 plus.t3 79.2293
R111 plus.n5 plus.t4 79.2293
R112 plus.n4 plus.t6 79.2293
R113 plus.n18 plus.t0 79.2293
R114 plus.n16 plus.t9 79.2293
R115 plus.n15 plus.t2 79.2293
R116 plus.n14 plus.t7 79.2293
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n7 plus.n6 32.1338
R122 plus.n17 plus.n16 32.1338
R123 plus.n3 plus.n2 31.8629
R124 plus.n13 plus.n12 31.8629
R125 plus plus.n19 26.8608
R126 plus.n4 plus.n3 16.2333
R127 plus.n14 plus.n13 16.2333
R128 plus.n8 plus.n7 16.0672
R129 plus.n18 plus.n17 16.0672
R130 plus plus.n9 8.15391
R131 plus.n2 plus.n1 0.380177
R132 plus.n12 plus.n11 0.380177
R133 plus.n1 plus.n0 0.285035
R134 plus.n11 plus.n10 0.285035
R135 plus.n9 plus.n0 0.189894
R136 plus.n19 plus.n10 0.189894
R137 drain_left.n5 drain_left.t1 260.906
R138 drain_left.n1 drain_left.t9 260.906
R139 drain_left.n3 drain_left.n2 240.808
R140 drain_left.n7 drain_left.n6 240.132
R141 drain_left.n5 drain_left.n4 240.132
R142 drain_left.n1 drain_left.n0 240.131
R143 drain_left drain_left.n3 23.1738
R144 drain_left.n2 drain_left.t2 19.8005
R145 drain_left.n2 drain_left.t8 19.8005
R146 drain_left.n0 drain_left.t0 19.8005
R147 drain_left.n0 drain_left.t7 19.8005
R148 drain_left.n6 drain_left.t6 19.8005
R149 drain_left.n6 drain_left.t4 19.8005
R150 drain_left.n4 drain_left.t3 19.8005
R151 drain_left.n4 drain_left.t5 19.8005
R152 drain_left drain_left.n7 6.62735
R153 drain_left.n7 drain_left.n5 0.974638
R154 drain_left.n3 drain_left.n1 0.188688
C0 drain_left minus 0.180282f
C1 drain_right minus 1.00766f
C2 drain_left source 3.5924f
C3 drain_right source 3.5934f
C4 drain_left plus 1.21005f
C5 drain_right plus 0.367711f
C6 drain_left drain_right 1.03066f
C7 minus source 1.51963f
C8 plus minus 3.69666f
C9 plus source 1.53353f
C10 drain_right a_n2072_n1088# 3.673105f
C11 drain_left a_n2072_n1088# 3.94356f
C12 source a_n2072_n1088# 2.242486f
C13 minus a_n2072_n1088# 7.196236f
C14 plus a_n2072_n1088# 7.802946f
C15 drain_left.t9 a_n2072_n1088# 0.091711f
C16 drain_left.t0 a_n2072_n1088# 0.014705f
C17 drain_left.t7 a_n2072_n1088# 0.014705f
C18 drain_left.n0 a_n2072_n1088# 0.057139f
C19 drain_left.n1 a_n2072_n1088# 0.403681f
C20 drain_left.t2 a_n2072_n1088# 0.014705f
C21 drain_left.t8 a_n2072_n1088# 0.014705f
C22 drain_left.n2 a_n2072_n1088# 0.057804f
C23 drain_left.n3 a_n2072_n1088# 0.798789f
C24 drain_left.t1 a_n2072_n1088# 0.091711f
C25 drain_left.t3 a_n2072_n1088# 0.014705f
C26 drain_left.t5 a_n2072_n1088# 0.014705f
C27 drain_left.n4 a_n2072_n1088# 0.057139f
C28 drain_left.n5 a_n2072_n1088# 0.448514f
C29 drain_left.t6 a_n2072_n1088# 0.014705f
C30 drain_left.t4 a_n2072_n1088# 0.014705f
C31 drain_left.n6 a_n2072_n1088# 0.057139f
C32 drain_left.n7 a_n2072_n1088# 0.413808f
C33 plus.n0 a_n2072_n1088# 0.036893f
C34 plus.t5 a_n2072_n1088# 0.075004f
C35 plus.t3 a_n2072_n1088# 0.075004f
C36 plus.n1 a_n2072_n1088# 0.046051f
C37 plus.t4 a_n2072_n1088# 0.075004f
C38 plus.n2 a_n2072_n1088# 0.169667f
C39 plus.t6 a_n2072_n1088# 0.075004f
C40 plus.t8 a_n2072_n1088# 0.091787f
C41 plus.n3 a_n2072_n1088# 0.060463f
C42 plus.n4 a_n2072_n1088# 0.079857f
C43 plus.n5 a_n2072_n1088# 0.080526f
C44 plus.n6 a_n2072_n1088# 0.078651f
C45 plus.n7 a_n2072_n1088# 0.006274f
C46 plus.n8 a_n2072_n1088# 0.070502f
C47 plus.n9 a_n2072_n1088# 0.201589f
C48 plus.n10 a_n2072_n1088# 0.036893f
C49 plus.t0 a_n2072_n1088# 0.075004f
C50 plus.n11 a_n2072_n1088# 0.046051f
C51 plus.t9 a_n2072_n1088# 0.075004f
C52 plus.n12 a_n2072_n1088# 0.169667f
C53 plus.t2 a_n2072_n1088# 0.075004f
C54 plus.t1 a_n2072_n1088# 0.091787f
C55 plus.n13 a_n2072_n1088# 0.060463f
C56 plus.t7 a_n2072_n1088# 0.075004f
C57 plus.n14 a_n2072_n1088# 0.079857f
C58 plus.n15 a_n2072_n1088# 0.080526f
C59 plus.n16 a_n2072_n1088# 0.078651f
C60 plus.n17 a_n2072_n1088# 0.006274f
C61 plus.n18 a_n2072_n1088# 0.070502f
C62 plus.n19 a_n2072_n1088# 0.653941f
C63 drain_right.t7 a_n2072_n1088# 0.093604f
C64 drain_right.t0 a_n2072_n1088# 0.015008f
C65 drain_right.t8 a_n2072_n1088# 0.015008f
C66 drain_right.n0 a_n2072_n1088# 0.058318f
C67 drain_right.n1 a_n2072_n1088# 0.412012f
C68 drain_right.t1 a_n2072_n1088# 0.015008f
C69 drain_right.t9 a_n2072_n1088# 0.015008f
C70 drain_right.n2 a_n2072_n1088# 0.058997f
C71 drain_right.n3 a_n2072_n1088# 0.778616f
C72 drain_right.t5 a_n2072_n1088# 0.015008f
C73 drain_right.t4 a_n2072_n1088# 0.015008f
C74 drain_right.n4 a_n2072_n1088# 0.059367f
C75 drain_right.t3 a_n2072_n1088# 0.015008f
C76 drain_right.t6 a_n2072_n1088# 0.015008f
C77 drain_right.n5 a_n2072_n1088# 0.058318f
C78 drain_right.n6 a_n2072_n1088# 0.51069f
C79 drain_right.t2 a_n2072_n1088# 0.092833f
C80 drain_right.n7 a_n2072_n1088# 0.385024f
C81 source.t2 a_n2072_n1088# 0.114221f
C82 source.n0 a_n2072_n1088# 0.554802f
C83 source.t0 a_n2072_n1088# 0.020522f
C84 source.t6 a_n2072_n1088# 0.020522f
C85 source.n1 a_n2072_n1088# 0.066555f
C86 source.n2 a_n2072_n1088# 0.322523f
C87 source.t4 a_n2072_n1088# 0.020522f
C88 source.t9 a_n2072_n1088# 0.020522f
C89 source.n3 a_n2072_n1088# 0.066555f
C90 source.n4 a_n2072_n1088# 0.321081f
C91 source.t16 a_n2072_n1088# 0.114221f
C92 source.n5 a_n2072_n1088# 0.329383f
C93 source.t18 a_n2072_n1088# 0.020522f
C94 source.t17 a_n2072_n1088# 0.020522f
C95 source.n6 a_n2072_n1088# 0.066555f
C96 source.n7 a_n2072_n1088# 0.322523f
C97 source.t15 a_n2072_n1088# 0.020522f
C98 source.t13 a_n2072_n1088# 0.020522f
C99 source.n8 a_n2072_n1088# 0.066555f
C100 source.n9 a_n2072_n1088# 0.843886f
C101 source.t7 a_n2072_n1088# 0.020522f
C102 source.t3 a_n2072_n1088# 0.020522f
C103 source.n10 a_n2072_n1088# 0.066555f
C104 source.n11 a_n2072_n1088# 0.843886f
C105 source.t5 a_n2072_n1088# 0.020522f
C106 source.t8 a_n2072_n1088# 0.020522f
C107 source.n12 a_n2072_n1088# 0.066555f
C108 source.n13 a_n2072_n1088# 0.322524f
C109 source.t1 a_n2072_n1088# 0.114221f
C110 source.n14 a_n2072_n1088# 0.329383f
C111 source.t19 a_n2072_n1088# 0.020522f
C112 source.t10 a_n2072_n1088# 0.020522f
C113 source.n15 a_n2072_n1088# 0.066555f
C114 source.n16 a_n2072_n1088# 0.321081f
C115 source.t12 a_n2072_n1088# 0.020522f
C116 source.t11 a_n2072_n1088# 0.020522f
C117 source.n17 a_n2072_n1088# 0.066555f
C118 source.n18 a_n2072_n1088# 0.322524f
C119 source.t14 a_n2072_n1088# 0.114221f
C120 source.n19 a_n2072_n1088# 0.463647f
C121 source.n20 a_n2072_n1088# 0.541371f
C122 minus.n0 a_n2072_n1088# 0.036344f
C123 minus.t3 a_n2072_n1088# 0.073887f
C124 minus.n1 a_n2072_n1088# 0.079328f
C125 minus.t6 a_n2072_n1088# 0.073887f
C126 minus.t5 a_n2072_n1088# 0.09042f
C127 minus.t4 a_n2072_n1088# 0.073887f
C128 minus.n2 a_n2072_n1088# 0.078669f
C129 minus.n3 a_n2072_n1088# 0.059563f
C130 minus.n4 a_n2072_n1088# 0.167142f
C131 minus.n5 a_n2072_n1088# 0.045366f
C132 minus.n6 a_n2072_n1088# 0.07748f
C133 minus.n7 a_n2072_n1088# 0.006181f
C134 minus.t7 a_n2072_n1088# 0.073887f
C135 minus.n8 a_n2072_n1088# 0.069453f
C136 minus.n9 a_n2072_n1088# 0.665524f
C137 minus.n10 a_n2072_n1088# 0.036344f
C138 minus.t1 a_n2072_n1088# 0.073887f
C139 minus.n11 a_n2072_n1088# 0.079328f
C140 minus.t2 a_n2072_n1088# 0.09042f
C141 minus.t9 a_n2072_n1088# 0.073887f
C142 minus.n12 a_n2072_n1088# 0.078669f
C143 minus.n13 a_n2072_n1088# 0.059563f
C144 minus.n14 a_n2072_n1088# 0.167142f
C145 minus.n15 a_n2072_n1088# 0.045366f
C146 minus.t8 a_n2072_n1088# 0.073887f
C147 minus.n16 a_n2072_n1088# 0.07748f
C148 minus.n17 a_n2072_n1088# 0.006181f
C149 minus.t0 a_n2072_n1088# 0.073887f
C150 minus.n18 a_n2072_n1088# 0.069453f
C151 minus.n19 a_n2072_n1088# 0.189307f
C152 minus.n20 a_n2072_n1088# 0.816298f
.ends

