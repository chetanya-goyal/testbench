* NGSPICE file created from diffpair645.ext - technology: sky130A

.subckt diffpair645 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t17 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X2 source.t20 minus.t1 drain_right.t10 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X3 source.t3 plus.t0 drain_left.t11 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X4 a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X5 a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X6 drain_left.t10 plus.t1 source.t7 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X7 source.t12 minus.t2 drain_right.t9 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X8 source.t4 plus.t2 drain_left.t9 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X9 drain_right.t8 minus.t3 source.t23 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X10 drain_right.t7 minus.t4 source.t19 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X11 source.t15 minus.t5 drain_right.t6 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X12 drain_left.t8 plus.t3 source.t6 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X13 source.t18 minus.t6 drain_right.t5 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X14 drain_left.t7 plus.t4 source.t8 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X15 source.t0 plus.t5 drain_left.t6 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X16 drain_right.t4 minus.t7 source.t22 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 drain_right.t3 minus.t8 source.t13 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X18 drain_left.t5 plus.t6 source.t10 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 source.t21 minus.t9 drain_right.t2 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X20 drain_right.t1 minus.t10 source.t14 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X21 source.t1 plus.t7 drain_left.t4 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 source.t5 plus.t8 drain_left.t3 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X23 a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X24 drain_left.t2 plus.t9 source.t2 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X25 drain_left.t1 plus.t10 source.t9 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X26 source.t16 minus.t11 drain_right.t0 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X27 source.t11 plus.t11 drain_left.t0 a_n1626_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
R0 minus.n13 minus.t9 4280.31
R1 minus.n2 minus.t3 4280.31
R2 minus.n28 minus.t10 4280.31
R3 minus.n17 minus.t1 4280.31
R4 minus.n12 minus.t4 4225.53
R5 minus.n10 minus.t6 4225.53
R6 minus.n3 minus.t7 4225.53
R7 minus.n4 minus.t2 4225.53
R8 minus.n27 minus.t5 4225.53
R9 minus.n25 minus.t0 4225.53
R10 minus.n19 minus.t11 4225.53
R11 minus.n18 minus.t8 4225.53
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 62.0763
R27 minus.n5 minus.n3 62.0763
R28 minus.n20 minus.n19 62.0763
R29 minus.n26 minus.n25 62.0763
R30 minus.n30 minus.n14 45.171
R31 minus.n13 minus.n12 40.1672
R32 minus.n4 minus.n2 40.1672
R33 minus.n18 minus.n17 40.1672
R34 minus.n28 minus.n27 40.1672
R35 minus.n12 minus.n11 32.8641
R36 minus.n5 minus.n4 32.8641
R37 minus.n20 minus.n18 32.8641
R38 minus.n27 minus.n26 32.8641
R39 minus.n10 minus.n9 10.955
R40 minus.n3 minus.n1 10.955
R41 minus.n19 minus.n16 10.955
R42 minus.n25 minus.n24 10.955
R43 minus.n30 minus.n29 6.54217
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 source.n5 source.t0 43.2366
R54 source.n6 source.t23 43.2366
R55 source.n11 source.t21 43.2366
R56 source.n23 source.t14 43.2365
R57 source.n18 source.t20 43.2365
R58 source.n17 source.t6 43.2365
R59 source.n12 source.t3 43.2365
R60 source.n0 source.t2 43.2365
R61 source.n22 source.n21 42.0366
R62 source.n20 source.n19 42.0366
R63 source.n16 source.n15 42.0366
R64 source.n14 source.n13 42.0366
R65 source.n2 source.n1 42.0366
R66 source.n4 source.n3 42.0366
R67 source.n8 source.n7 42.0366
R68 source.n10 source.n9 42.0366
R69 source.n12 source.n11 31.6966
R70 source.n24 source.n0 26.1535
R71 source.n24 source.n23 5.5436
R72 source.n21 source.t17 1.2005
R73 source.n21 source.t15 1.2005
R74 source.n19 source.t13 1.2005
R75 source.n19 source.t16 1.2005
R76 source.n15 source.t7 1.2005
R77 source.n15 source.t1 1.2005
R78 source.n13 source.t8 1.2005
R79 source.n13 source.t4 1.2005
R80 source.n1 source.t10 1.2005
R81 source.n1 source.t11 1.2005
R82 source.n3 source.t9 1.2005
R83 source.n3 source.t5 1.2005
R84 source.n7 source.t22 1.2005
R85 source.n7 source.t12 1.2005
R86 source.n9 source.t19 1.2005
R87 source.n9 source.t18 1.2005
R88 source.n11 source.n10 0.560845
R89 source.n10 source.n8 0.560845
R90 source.n8 source.n6 0.560845
R91 source.n5 source.n4 0.560845
R92 source.n4 source.n2 0.560845
R93 source.n2 source.n0 0.560845
R94 source.n14 source.n12 0.560845
R95 source.n16 source.n14 0.560845
R96 source.n17 source.n16 0.560845
R97 source.n20 source.n18 0.560845
R98 source.n22 source.n20 0.560845
R99 source.n23 source.n22 0.560845
R100 source.n6 source.n5 0.470328
R101 source.n18 source.n17 0.470328
R102 source source.n24 0.188
R103 drain_right.n6 drain_right.n4 59.2756
R104 drain_right.n3 drain_right.n2 59.2204
R105 drain_right.n3 drain_right.n0 59.2204
R106 drain_right.n3 drain_right.n1 58.7154
R107 drain_right.n6 drain_right.n5 58.7154
R108 drain_right.n8 drain_right.n7 58.7154
R109 drain_right drain_right.n3 39.4641
R110 drain_right drain_right.n8 6.21356
R111 drain_right.n1 drain_right.t0 1.2005
R112 drain_right.n1 drain_right.t11 1.2005
R113 drain_right.n2 drain_right.t6 1.2005
R114 drain_right.n2 drain_right.t1 1.2005
R115 drain_right.n0 drain_right.t10 1.2005
R116 drain_right.n0 drain_right.t3 1.2005
R117 drain_right.n4 drain_right.t9 1.2005
R118 drain_right.n4 drain_right.t8 1.2005
R119 drain_right.n5 drain_right.t5 1.2005
R120 drain_right.n5 drain_right.t4 1.2005
R121 drain_right.n7 drain_right.t2 1.2005
R122 drain_right.n7 drain_right.t7 1.2005
R123 drain_right.n8 drain_right.n6 0.560845
R124 plus.n2 plus.t5 4280.31
R125 plus.n13 plus.t9 4280.31
R126 plus.n17 plus.t3 4280.31
R127 plus.n28 plus.t0 4280.31
R128 plus.n3 plus.t10 4225.53
R129 plus.n4 plus.t8 4225.53
R130 plus.n10 plus.t6 4225.53
R131 plus.n12 plus.t11 4225.53
R132 plus.n19 plus.t7 4225.53
R133 plus.n18 plus.t1 4225.53
R134 plus.n25 plus.t2 4225.53
R135 plus.n27 plus.t4 4225.53
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 62.0763
R151 plus.n11 plus.n10 62.0763
R152 plus.n26 plus.n25 62.0763
R153 plus.n20 plus.n18 62.0763
R154 plus.n3 plus.n2 40.1672
R155 plus.n13 plus.n12 40.1672
R156 plus.n28 plus.n27 40.1672
R157 plus.n19 plus.n17 40.1672
R158 plus plus.n29 34.1278
R159 plus.n5 plus.n3 32.8641
R160 plus.n12 plus.n11 32.8641
R161 plus.n27 plus.n26 32.8641
R162 plus.n20 plus.n19 32.8641
R163 plus plus.n14 17.1103
R164 plus.n4 plus.n1 10.955
R165 plus.n10 plus.n9 10.955
R166 plus.n25 plus.n24 10.955
R167 plus.n18 plus.n16 10.955
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 59.2758
R177 drain_left.n3 drain_left.n2 59.2204
R178 drain_left.n3 drain_left.n0 59.2204
R179 drain_left.n3 drain_left.n1 58.7154
R180 drain_left.n6 drain_left.n5 58.7154
R181 drain_left.n8 drain_left.n7 58.7153
R182 drain_left drain_left.n3 40.0173
R183 drain_left drain_left.n8 6.21356
R184 drain_left.n1 drain_left.t9 1.2005
R185 drain_left.n1 drain_left.t10 1.2005
R186 drain_left.n2 drain_left.t4 1.2005
R187 drain_left.n2 drain_left.t8 1.2005
R188 drain_left.n0 drain_left.t11 1.2005
R189 drain_left.n0 drain_left.t7 1.2005
R190 drain_left.n7 drain_left.t0 1.2005
R191 drain_left.n7 drain_left.t2 1.2005
R192 drain_left.n5 drain_left.t3 1.2005
R193 drain_left.n5 drain_left.t5 1.2005
R194 drain_left.n4 drain_left.t6 1.2005
R195 drain_left.n4 drain_left.t1 1.2005
R196 drain_left.n8 drain_left.n6 0.560845
C0 drain_left drain_right 0.801529f
C1 plus source 4.35321f
C2 plus minus 7.57115f
C3 drain_right source 47.465f
C4 drain_right minus 5.48942f
C5 drain_left source 47.4651f
C6 drain_left minus 0.170585f
C7 drain_right plus 0.309819f
C8 drain_left plus 5.64591f
C9 minus source 4.33917f
C10 drain_right a_n1626_n5888# 8.11366f
C11 drain_left a_n1626_n5888# 8.35622f
C12 source a_n1626_n5888# 15.746701f
C13 minus a_n1626_n5888# 6.857574f
C14 plus a_n1626_n5888# 10.00658f
C15 drain_left.t11 a_n1626_n5888# 0.845917f
C16 drain_left.t7 a_n1626_n5888# 0.845917f
C17 drain_left.n0 a_n1626_n5888# 5.72358f
C18 drain_left.t9 a_n1626_n5888# 0.845917f
C19 drain_left.t10 a_n1626_n5888# 0.845917f
C20 drain_left.n1 a_n1626_n5888# 5.72061f
C21 drain_left.t4 a_n1626_n5888# 0.845917f
C22 drain_left.t8 a_n1626_n5888# 0.845917f
C23 drain_left.n2 a_n1626_n5888# 5.72358f
C24 drain_left.n3 a_n1626_n5888# 3.23221f
C25 drain_left.t6 a_n1626_n5888# 0.845917f
C26 drain_left.t1 a_n1626_n5888# 0.845917f
C27 drain_left.n4 a_n1626_n5888# 5.72394f
C28 drain_left.t3 a_n1626_n5888# 0.845917f
C29 drain_left.t5 a_n1626_n5888# 0.845917f
C30 drain_left.n5 a_n1626_n5888# 5.72061f
C31 drain_left.n6 a_n1626_n5888# 0.689917f
C32 drain_left.t0 a_n1626_n5888# 0.845917f
C33 drain_left.t2 a_n1626_n5888# 0.845917f
C34 drain_left.n7 a_n1626_n5888# 5.7206f
C35 drain_left.n8 a_n1626_n5888# 0.576949f
C36 plus.n0 a_n1626_n5888# 0.058124f
C37 plus.t11 a_n1626_n5888# 0.613281f
C38 plus.t6 a_n1626_n5888# 0.613281f
C39 plus.n1 a_n1626_n5888# 0.021969f
C40 plus.t5 a_n1626_n5888# 0.616263f
C41 plus.n2 a_n1626_n5888# 0.254775f
C42 plus.t10 a_n1626_n5888# 0.613281f
C43 plus.n3 a_n1626_n5888# 0.232118f
C44 plus.t8 a_n1626_n5888# 0.613281f
C45 plus.n4 a_n1626_n5888# 0.232118f
C46 plus.n5 a_n1626_n5888# 0.024657f
C47 plus.n6 a_n1626_n5888# 0.130497f
C48 plus.n7 a_n1626_n5888# 0.058124f
C49 plus.n8 a_n1626_n5888# 0.058124f
C50 plus.n9 a_n1626_n5888# 0.021969f
C51 plus.n10 a_n1626_n5888# 0.232118f
C52 plus.n11 a_n1626_n5888# 0.024657f
C53 plus.n12 a_n1626_n5888# 0.232118f
C54 plus.t9 a_n1626_n5888# 0.616263f
C55 plus.n13 a_n1626_n5888# 0.25469f
C56 plus.n14 a_n1626_n5888# 1.04306f
C57 plus.n15 a_n1626_n5888# 0.058124f
C58 plus.t0 a_n1626_n5888# 0.616263f
C59 plus.t4 a_n1626_n5888# 0.613281f
C60 plus.t2 a_n1626_n5888# 0.613281f
C61 plus.n16 a_n1626_n5888# 0.021969f
C62 plus.t3 a_n1626_n5888# 0.616263f
C63 plus.n17 a_n1626_n5888# 0.254775f
C64 plus.t1 a_n1626_n5888# 0.613281f
C65 plus.n18 a_n1626_n5888# 0.232118f
C66 plus.t7 a_n1626_n5888# 0.613281f
C67 plus.n19 a_n1626_n5888# 0.232118f
C68 plus.n20 a_n1626_n5888# 0.024657f
C69 plus.n21 a_n1626_n5888# 0.130497f
C70 plus.n22 a_n1626_n5888# 0.058124f
C71 plus.n23 a_n1626_n5888# 0.058124f
C72 plus.n24 a_n1626_n5888# 0.021969f
C73 plus.n25 a_n1626_n5888# 0.232118f
C74 plus.n26 a_n1626_n5888# 0.024657f
C75 plus.n27 a_n1626_n5888# 0.232118f
C76 plus.n28 a_n1626_n5888# 0.25469f
C77 plus.n29 a_n1626_n5888# 2.18341f
C78 drain_right.t10 a_n1626_n5888# 0.846086f
C79 drain_right.t3 a_n1626_n5888# 0.846086f
C80 drain_right.n0 a_n1626_n5888# 5.72472f
C81 drain_right.t0 a_n1626_n5888# 0.846086f
C82 drain_right.t11 a_n1626_n5888# 0.846086f
C83 drain_right.n1 a_n1626_n5888# 5.72175f
C84 drain_right.t6 a_n1626_n5888# 0.846086f
C85 drain_right.t1 a_n1626_n5888# 0.846086f
C86 drain_right.n2 a_n1626_n5888# 5.72472f
C87 drain_right.n3 a_n1626_n5888# 3.17409f
C88 drain_right.t9 a_n1626_n5888# 0.846086f
C89 drain_right.t8 a_n1626_n5888# 0.846086f
C90 drain_right.n4 a_n1626_n5888# 5.72507f
C91 drain_right.t5 a_n1626_n5888# 0.846086f
C92 drain_right.t4 a_n1626_n5888# 0.846086f
C93 drain_right.n5 a_n1626_n5888# 5.72175f
C94 drain_right.n6 a_n1626_n5888# 0.690067f
C95 drain_right.t2 a_n1626_n5888# 0.846086f
C96 drain_right.t7 a_n1626_n5888# 0.846086f
C97 drain_right.n7 a_n1626_n5888# 5.72175f
C98 drain_right.n8 a_n1626_n5888# 0.577052f
C99 source.t2 a_n1626_n5888# 5.45484f
C100 source.n0 a_n1626_n5888# 2.08728f
C101 source.t10 a_n1626_n5888# 0.661496f
C102 source.t11 a_n1626_n5888# 0.661496f
C103 source.n1 a_n1626_n5888# 4.401f
C104 source.n2 a_n1626_n5888# 0.309016f
C105 source.t9 a_n1626_n5888# 0.661496f
C106 source.t5 a_n1626_n5888# 0.661496f
C107 source.n3 a_n1626_n5888# 4.401f
C108 source.n4 a_n1626_n5888# 0.309016f
C109 source.t0 a_n1626_n5888# 5.45485f
C110 source.n5 a_n1626_n5888# 0.439406f
C111 source.t23 a_n1626_n5888# 5.45485f
C112 source.n6 a_n1626_n5888# 0.439406f
C113 source.t22 a_n1626_n5888# 0.661496f
C114 source.t12 a_n1626_n5888# 0.661496f
C115 source.n7 a_n1626_n5888# 4.401f
C116 source.n8 a_n1626_n5888# 0.309016f
C117 source.t19 a_n1626_n5888# 0.661496f
C118 source.t18 a_n1626_n5888# 0.661496f
C119 source.n9 a_n1626_n5888# 4.401f
C120 source.n10 a_n1626_n5888# 0.309016f
C121 source.t21 a_n1626_n5888# 5.45485f
C122 source.n11 a_n1626_n5888# 2.49665f
C123 source.t3 a_n1626_n5888# 5.45484f
C124 source.n12 a_n1626_n5888# 2.49666f
C125 source.t8 a_n1626_n5888# 0.661496f
C126 source.t4 a_n1626_n5888# 0.661496f
C127 source.n13 a_n1626_n5888# 4.401f
C128 source.n14 a_n1626_n5888# 0.309018f
C129 source.t7 a_n1626_n5888# 0.661496f
C130 source.t1 a_n1626_n5888# 0.661496f
C131 source.n15 a_n1626_n5888# 4.401f
C132 source.n16 a_n1626_n5888# 0.309018f
C133 source.t6 a_n1626_n5888# 5.45484f
C134 source.n17 a_n1626_n5888# 0.43942f
C135 source.t20 a_n1626_n5888# 5.45484f
C136 source.n18 a_n1626_n5888# 0.43942f
C137 source.t13 a_n1626_n5888# 0.661496f
C138 source.t16 a_n1626_n5888# 0.661496f
C139 source.n19 a_n1626_n5888# 4.401f
C140 source.n20 a_n1626_n5888# 0.309018f
C141 source.t17 a_n1626_n5888# 0.661496f
C142 source.t15 a_n1626_n5888# 0.661496f
C143 source.n21 a_n1626_n5888# 4.401f
C144 source.n22 a_n1626_n5888# 0.309018f
C145 source.t14 a_n1626_n5888# 5.45484f
C146 source.n23 a_n1626_n5888# 0.565151f
C147 source.n24 a_n1626_n5888# 2.35661f
C148 minus.n0 a_n1626_n5888# 0.057082f
C149 minus.t9 a_n1626_n5888# 0.605218f
C150 minus.t4 a_n1626_n5888# 0.60229f
C151 minus.t6 a_n1626_n5888# 0.60229f
C152 minus.n1 a_n1626_n5888# 0.021576f
C153 minus.t3 a_n1626_n5888# 0.605218f
C154 minus.n2 a_n1626_n5888# 0.250208f
C155 minus.t7 a_n1626_n5888# 0.60229f
C156 minus.n3 a_n1626_n5888# 0.227958f
C157 minus.t2 a_n1626_n5888# 0.60229f
C158 minus.n4 a_n1626_n5888# 0.227958f
C159 minus.n5 a_n1626_n5888# 0.024215f
C160 minus.n6 a_n1626_n5888# 0.128158f
C161 minus.n7 a_n1626_n5888# 0.057082f
C162 minus.n8 a_n1626_n5888# 0.057082f
C163 minus.n9 a_n1626_n5888# 0.021576f
C164 minus.n10 a_n1626_n5888# 0.227958f
C165 minus.n11 a_n1626_n5888# 0.024215f
C166 minus.n12 a_n1626_n5888# 0.227958f
C167 minus.n13 a_n1626_n5888# 0.250125f
C168 minus.n14 a_n1626_n5888# 2.81145f
C169 minus.n15 a_n1626_n5888# 0.057082f
C170 minus.t5 a_n1626_n5888# 0.60229f
C171 minus.t0 a_n1626_n5888# 0.60229f
C172 minus.n16 a_n1626_n5888# 0.021576f
C173 minus.t1 a_n1626_n5888# 0.605218f
C174 minus.n17 a_n1626_n5888# 0.250208f
C175 minus.t8 a_n1626_n5888# 0.60229f
C176 minus.n18 a_n1626_n5888# 0.227958f
C177 minus.t11 a_n1626_n5888# 0.60229f
C178 minus.n19 a_n1626_n5888# 0.227958f
C179 minus.n20 a_n1626_n5888# 0.024215f
C180 minus.n21 a_n1626_n5888# 0.128158f
C181 minus.n22 a_n1626_n5888# 0.057082f
C182 minus.n23 a_n1626_n5888# 0.057082f
C183 minus.n24 a_n1626_n5888# 0.021576f
C184 minus.n25 a_n1626_n5888# 0.227958f
C185 minus.n26 a_n1626_n5888# 0.024215f
C186 minus.n27 a_n1626_n5888# 0.227958f
C187 minus.t10 a_n1626_n5888# 0.605218f
C188 minus.n28 a_n1626_n5888# 0.250125f
C189 minus.n29 a_n1626_n5888# 0.378847f
C190 minus.n30 a_n1626_n5888# 3.32672f
.ends

