* NGSPICE file created from diffpair318.ext - technology: sky130A

.subckt diffpair318 minus drain_right drain_left source plus
X0 a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X1 source.t37 plus.t0 drain_left.t2 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 drain_left.t11 plus.t1 source.t36 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X3 a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X4 a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X5 drain_right.t19 minus.t0 source.t8 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X6 drain_left.t9 plus.t2 source.t35 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X7 a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X8 drain_left.t12 plus.t3 source.t34 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X9 drain_left.t7 plus.t4 source.t33 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X10 source.t7 minus.t1 drain_right.t18 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X11 source.t13 minus.t2 drain_right.t17 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X12 source.t3 minus.t3 drain_right.t16 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X13 source.t14 minus.t4 drain_right.t15 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X14 source.t32 plus.t5 drain_left.t8 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X15 drain_right.t14 minus.t5 source.t5 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X16 drain_left.t3 plus.t6 source.t31 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X17 source.t1 minus.t6 drain_right.t13 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X18 drain_left.t1 plus.t7 source.t30 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X19 source.t9 minus.t7 drain_right.t12 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X20 drain_right.t11 minus.t8 source.t0 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X21 source.t15 minus.t9 drain_right.t10 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X22 source.t29 plus.t8 drain_left.t0 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X23 drain_right.t9 minus.t10 source.t2 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X24 source.t28 plus.t9 drain_left.t14 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X25 source.t38 minus.t11 drain_right.t8 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X26 drain_right.t7 minus.t12 source.t16 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X27 drain_left.t15 plus.t10 source.t27 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X28 source.t12 minus.t13 drain_right.t6 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X29 drain_right.t5 minus.t14 source.t6 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X30 drain_right.t4 minus.t15 source.t4 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X31 drain_right.t3 minus.t16 source.t10 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X32 source.t26 plus.t11 drain_left.t5 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X33 source.t25 plus.t12 drain_left.t4 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X34 drain_left.t18 plus.t13 source.t24 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X35 drain_left.t17 plus.t14 source.t23 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X36 source.t17 minus.t17 drain_right.t2 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X37 source.t22 plus.t15 drain_left.t16 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X38 drain_right.t1 minus.t18 source.t39 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X39 source.t21 plus.t16 drain_left.t6 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X40 drain_left.t19 plus.t17 source.t20 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X41 source.t19 plus.t18 drain_left.t10 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X42 drain_right.t0 minus.t19 source.t11 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X43 source.t18 plus.t19 drain_left.t13 a_n3202_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
R0 plus.n9 plus.t18 251.644
R1 plus.n39 plus.t6 251.644
R2 plus.n28 plus.t7 229.855
R3 plus.n26 plus.t9 229.855
R4 plus.n2 plus.t10 229.855
R5 plus.n21 plus.t11 229.855
R6 plus.n19 plus.t13 229.855
R7 plus.n5 plus.t16 229.855
R8 plus.n13 plus.t14 229.855
R9 plus.n12 plus.t15 229.855
R10 plus.n8 plus.t17 229.855
R11 plus.n58 plus.t5 229.855
R12 plus.n56 plus.t1 229.855
R13 plus.n32 plus.t12 229.855
R14 plus.n51 plus.t2 229.855
R15 plus.n49 plus.t8 229.855
R16 plus.n35 plus.t4 229.855
R17 plus.n43 plus.t19 229.855
R18 plus.n42 plus.t3 229.855
R19 plus.n38 plus.t0 229.855
R20 plus.n11 plus.n10 161.3
R21 plus.n15 plus.n14 161.3
R22 plus.n16 plus.n5 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n4 161.3
R25 plus.n20 plus.n3 161.3
R26 plus.n25 plus.n24 161.3
R27 plus.n26 plus.n1 161.3
R28 plus.n27 plus.n0 161.3
R29 plus.n29 plus.n28 161.3
R30 plus.n41 plus.n40 161.3
R31 plus.n45 plus.n44 161.3
R32 plus.n46 plus.n35 161.3
R33 plus.n48 plus.n47 161.3
R34 plus.n49 plus.n34 161.3
R35 plus.n50 plus.n33 161.3
R36 plus.n55 plus.n54 161.3
R37 plus.n56 plus.n31 161.3
R38 plus.n57 plus.n30 161.3
R39 plus.n59 plus.n58 161.3
R40 plus.n12 plus.n7 80.6037
R41 plus.n13 plus.n6 80.6037
R42 plus.n22 plus.n21 80.6037
R43 plus.n23 plus.n2 80.6037
R44 plus.n42 plus.n37 80.6037
R45 plus.n43 plus.n36 80.6037
R46 plus.n52 plus.n51 80.6037
R47 plus.n53 plus.n32 80.6037
R48 plus.n21 plus.n2 48.2005
R49 plus.n13 plus.n12 48.2005
R50 plus.n51 plus.n32 48.2005
R51 plus.n43 plus.n42 48.2005
R52 plus.n40 plus.n39 44.8565
R53 plus.n10 plus.n9 44.8565
R54 plus.n21 plus.n20 43.0884
R55 plus.n14 plus.n13 43.0884
R56 plus.n51 plus.n50 43.0884
R57 plus.n44 plus.n43 43.0884
R58 plus.n25 plus.n2 40.1672
R59 plus.n12 plus.n11 40.1672
R60 plus.n55 plus.n32 40.1672
R61 plus.n42 plus.n41 40.1672
R62 plus plus.n59 33.0634
R63 plus.n28 plus.n27 27.0217
R64 plus.n58 plus.n57 27.0217
R65 plus.n18 plus.n5 24.1005
R66 plus.n19 plus.n18 24.1005
R67 plus.n49 plus.n48 24.1005
R68 plus.n48 plus.n35 24.1005
R69 plus.n27 plus.n26 21.1793
R70 plus.n57 plus.n56 21.1793
R71 plus.n39 plus.n38 20.1275
R72 plus.n9 plus.n8 20.1275
R73 plus plus.n29 10.0763
R74 plus.n26 plus.n25 8.03383
R75 plus.n11 plus.n8 8.03383
R76 plus.n56 plus.n55 8.03383
R77 plus.n41 plus.n38 8.03383
R78 plus.n20 plus.n19 5.11262
R79 plus.n14 plus.n5 5.11262
R80 plus.n50 plus.n49 5.11262
R81 plus.n44 plus.n35 5.11262
R82 plus.n7 plus.n6 0.380177
R83 plus.n23 plus.n22 0.380177
R84 plus.n53 plus.n52 0.380177
R85 plus.n37 plus.n36 0.380177
R86 plus.n10 plus.n7 0.285035
R87 plus.n15 plus.n6 0.285035
R88 plus.n22 plus.n3 0.285035
R89 plus.n24 plus.n23 0.285035
R90 plus.n54 plus.n53 0.285035
R91 plus.n52 plus.n33 0.285035
R92 plus.n45 plus.n36 0.285035
R93 plus.n40 plus.n37 0.285035
R94 plus.n16 plus.n15 0.189894
R95 plus.n17 plus.n16 0.189894
R96 plus.n17 plus.n4 0.189894
R97 plus.n4 plus.n3 0.189894
R98 plus.n24 plus.n1 0.189894
R99 plus.n1 plus.n0 0.189894
R100 plus.n29 plus.n0 0.189894
R101 plus.n59 plus.n30 0.189894
R102 plus.n31 plus.n30 0.189894
R103 plus.n54 plus.n31 0.189894
R104 plus.n34 plus.n33 0.189894
R105 plus.n47 plus.n34 0.189894
R106 plus.n47 plus.n46 0.189894
R107 plus.n46 plus.n45 0.189894
R108 drain_left.n10 drain_left.n8 68.165
R109 drain_left.n6 drain_left.n4 68.1648
R110 drain_left.n2 drain_left.n0 68.1648
R111 drain_left.n14 drain_left.n13 67.1908
R112 drain_left.n12 drain_left.n11 67.1908
R113 drain_left.n10 drain_left.n9 67.1908
R114 drain_left.n16 drain_left.n15 67.1907
R115 drain_left.n7 drain_left.n3 67.1907
R116 drain_left.n6 drain_left.n5 67.1907
R117 drain_left.n2 drain_left.n1 67.1907
R118 drain_left drain_left.n7 30.6147
R119 drain_left drain_left.n16 6.62735
R120 drain_left.n3 drain_left.t0 3.3005
R121 drain_left.n3 drain_left.t7 3.3005
R122 drain_left.n4 drain_left.t2 3.3005
R123 drain_left.n4 drain_left.t3 3.3005
R124 drain_left.n5 drain_left.t13 3.3005
R125 drain_left.n5 drain_left.t12 3.3005
R126 drain_left.n1 drain_left.t4 3.3005
R127 drain_left.n1 drain_left.t9 3.3005
R128 drain_left.n0 drain_left.t8 3.3005
R129 drain_left.n0 drain_left.t11 3.3005
R130 drain_left.n15 drain_left.t14 3.3005
R131 drain_left.n15 drain_left.t1 3.3005
R132 drain_left.n13 drain_left.t5 3.3005
R133 drain_left.n13 drain_left.t15 3.3005
R134 drain_left.n11 drain_left.t6 3.3005
R135 drain_left.n11 drain_left.t18 3.3005
R136 drain_left.n9 drain_left.t16 3.3005
R137 drain_left.n9 drain_left.t17 3.3005
R138 drain_left.n8 drain_left.t10 3.3005
R139 drain_left.n8 drain_left.t19 3.3005
R140 drain_left.n12 drain_left.n10 0.974638
R141 drain_left.n14 drain_left.n12 0.974638
R142 drain_left.n16 drain_left.n14 0.974638
R143 drain_left.n7 drain_left.n6 0.919292
R144 drain_left.n7 drain_left.n2 0.919292
R145 source.n282 source.n256 289.615
R146 source.n242 source.n216 289.615
R147 source.n210 source.n184 289.615
R148 source.n170 source.n144 289.615
R149 source.n26 source.n0 289.615
R150 source.n66 source.n40 289.615
R151 source.n98 source.n72 289.615
R152 source.n138 source.n112 289.615
R153 source.n267 source.n266 185
R154 source.n264 source.n263 185
R155 source.n273 source.n272 185
R156 source.n275 source.n274 185
R157 source.n260 source.n259 185
R158 source.n281 source.n280 185
R159 source.n283 source.n282 185
R160 source.n227 source.n226 185
R161 source.n224 source.n223 185
R162 source.n233 source.n232 185
R163 source.n235 source.n234 185
R164 source.n220 source.n219 185
R165 source.n241 source.n240 185
R166 source.n243 source.n242 185
R167 source.n195 source.n194 185
R168 source.n192 source.n191 185
R169 source.n201 source.n200 185
R170 source.n203 source.n202 185
R171 source.n188 source.n187 185
R172 source.n209 source.n208 185
R173 source.n211 source.n210 185
R174 source.n155 source.n154 185
R175 source.n152 source.n151 185
R176 source.n161 source.n160 185
R177 source.n163 source.n162 185
R178 source.n148 source.n147 185
R179 source.n169 source.n168 185
R180 source.n171 source.n170 185
R181 source.n27 source.n26 185
R182 source.n25 source.n24 185
R183 source.n4 source.n3 185
R184 source.n19 source.n18 185
R185 source.n17 source.n16 185
R186 source.n8 source.n7 185
R187 source.n11 source.n10 185
R188 source.n67 source.n66 185
R189 source.n65 source.n64 185
R190 source.n44 source.n43 185
R191 source.n59 source.n58 185
R192 source.n57 source.n56 185
R193 source.n48 source.n47 185
R194 source.n51 source.n50 185
R195 source.n99 source.n98 185
R196 source.n97 source.n96 185
R197 source.n76 source.n75 185
R198 source.n91 source.n90 185
R199 source.n89 source.n88 185
R200 source.n80 source.n79 185
R201 source.n83 source.n82 185
R202 source.n139 source.n138 185
R203 source.n137 source.n136 185
R204 source.n116 source.n115 185
R205 source.n131 source.n130 185
R206 source.n129 source.n128 185
R207 source.n120 source.n119 185
R208 source.n123 source.n122 185
R209 source.t10 source.n265 147.661
R210 source.t15 source.n225 147.661
R211 source.t31 source.n193 147.661
R212 source.t32 source.n153 147.661
R213 source.t30 source.n9 147.661
R214 source.t19 source.n49 147.661
R215 source.t2 source.n81 147.661
R216 source.t13 source.n121 147.661
R217 source.n266 source.n263 104.615
R218 source.n273 source.n263 104.615
R219 source.n274 source.n273 104.615
R220 source.n274 source.n259 104.615
R221 source.n281 source.n259 104.615
R222 source.n282 source.n281 104.615
R223 source.n226 source.n223 104.615
R224 source.n233 source.n223 104.615
R225 source.n234 source.n233 104.615
R226 source.n234 source.n219 104.615
R227 source.n241 source.n219 104.615
R228 source.n242 source.n241 104.615
R229 source.n194 source.n191 104.615
R230 source.n201 source.n191 104.615
R231 source.n202 source.n201 104.615
R232 source.n202 source.n187 104.615
R233 source.n209 source.n187 104.615
R234 source.n210 source.n209 104.615
R235 source.n154 source.n151 104.615
R236 source.n161 source.n151 104.615
R237 source.n162 source.n161 104.615
R238 source.n162 source.n147 104.615
R239 source.n169 source.n147 104.615
R240 source.n170 source.n169 104.615
R241 source.n26 source.n25 104.615
R242 source.n25 source.n3 104.615
R243 source.n18 source.n3 104.615
R244 source.n18 source.n17 104.615
R245 source.n17 source.n7 104.615
R246 source.n10 source.n7 104.615
R247 source.n66 source.n65 104.615
R248 source.n65 source.n43 104.615
R249 source.n58 source.n43 104.615
R250 source.n58 source.n57 104.615
R251 source.n57 source.n47 104.615
R252 source.n50 source.n47 104.615
R253 source.n98 source.n97 104.615
R254 source.n97 source.n75 104.615
R255 source.n90 source.n75 104.615
R256 source.n90 source.n89 104.615
R257 source.n89 source.n79 104.615
R258 source.n82 source.n79 104.615
R259 source.n138 source.n137 104.615
R260 source.n137 source.n115 104.615
R261 source.n130 source.n115 104.615
R262 source.n130 source.n129 104.615
R263 source.n129 source.n119 104.615
R264 source.n122 source.n119 104.615
R265 source.n266 source.t10 52.3082
R266 source.n226 source.t15 52.3082
R267 source.n194 source.t31 52.3082
R268 source.n154 source.t32 52.3082
R269 source.n10 source.t30 52.3082
R270 source.n50 source.t19 52.3082
R271 source.n82 source.t2 52.3082
R272 source.n122 source.t13 52.3082
R273 source.n33 source.n32 50.512
R274 source.n35 source.n34 50.512
R275 source.n37 source.n36 50.512
R276 source.n39 source.n38 50.512
R277 source.n105 source.n104 50.512
R278 source.n107 source.n106 50.512
R279 source.n109 source.n108 50.512
R280 source.n111 source.n110 50.512
R281 source.n255 source.n254 50.5119
R282 source.n253 source.n252 50.5119
R283 source.n251 source.n250 50.5119
R284 source.n249 source.n248 50.5119
R285 source.n183 source.n182 50.5119
R286 source.n181 source.n180 50.5119
R287 source.n179 source.n178 50.5119
R288 source.n177 source.n176 50.5119
R289 source.n287 source.n286 32.1853
R290 source.n247 source.n246 32.1853
R291 source.n215 source.n214 32.1853
R292 source.n175 source.n174 32.1853
R293 source.n31 source.n30 32.1853
R294 source.n71 source.n70 32.1853
R295 source.n103 source.n102 32.1853
R296 source.n143 source.n142 32.1853
R297 source.n175 source.n143 17.7164
R298 source.n267 source.n265 15.6674
R299 source.n227 source.n225 15.6674
R300 source.n195 source.n193 15.6674
R301 source.n155 source.n153 15.6674
R302 source.n11 source.n9 15.6674
R303 source.n51 source.n49 15.6674
R304 source.n83 source.n81 15.6674
R305 source.n123 source.n121 15.6674
R306 source.n268 source.n264 12.8005
R307 source.n228 source.n224 12.8005
R308 source.n196 source.n192 12.8005
R309 source.n156 source.n152 12.8005
R310 source.n12 source.n8 12.8005
R311 source.n52 source.n48 12.8005
R312 source.n84 source.n80 12.8005
R313 source.n124 source.n120 12.8005
R314 source.n272 source.n271 12.0247
R315 source.n232 source.n231 12.0247
R316 source.n200 source.n199 12.0247
R317 source.n160 source.n159 12.0247
R318 source.n16 source.n15 12.0247
R319 source.n56 source.n55 12.0247
R320 source.n88 source.n87 12.0247
R321 source.n128 source.n127 12.0247
R322 source.n288 source.n31 11.9664
R323 source.n275 source.n262 11.249
R324 source.n235 source.n222 11.249
R325 source.n203 source.n190 11.249
R326 source.n163 source.n150 11.249
R327 source.n19 source.n6 11.249
R328 source.n59 source.n46 11.249
R329 source.n91 source.n78 11.249
R330 source.n131 source.n118 11.249
R331 source.n276 source.n260 10.4732
R332 source.n236 source.n220 10.4732
R333 source.n204 source.n188 10.4732
R334 source.n164 source.n148 10.4732
R335 source.n20 source.n4 10.4732
R336 source.n60 source.n44 10.4732
R337 source.n92 source.n76 10.4732
R338 source.n132 source.n116 10.4732
R339 source.n280 source.n279 9.69747
R340 source.n240 source.n239 9.69747
R341 source.n208 source.n207 9.69747
R342 source.n168 source.n167 9.69747
R343 source.n24 source.n23 9.69747
R344 source.n64 source.n63 9.69747
R345 source.n96 source.n95 9.69747
R346 source.n136 source.n135 9.69747
R347 source.n286 source.n285 9.45567
R348 source.n246 source.n245 9.45567
R349 source.n214 source.n213 9.45567
R350 source.n174 source.n173 9.45567
R351 source.n30 source.n29 9.45567
R352 source.n70 source.n69 9.45567
R353 source.n102 source.n101 9.45567
R354 source.n142 source.n141 9.45567
R355 source.n285 source.n284 9.3005
R356 source.n258 source.n257 9.3005
R357 source.n279 source.n278 9.3005
R358 source.n277 source.n276 9.3005
R359 source.n262 source.n261 9.3005
R360 source.n271 source.n270 9.3005
R361 source.n269 source.n268 9.3005
R362 source.n245 source.n244 9.3005
R363 source.n218 source.n217 9.3005
R364 source.n239 source.n238 9.3005
R365 source.n237 source.n236 9.3005
R366 source.n222 source.n221 9.3005
R367 source.n231 source.n230 9.3005
R368 source.n229 source.n228 9.3005
R369 source.n213 source.n212 9.3005
R370 source.n186 source.n185 9.3005
R371 source.n207 source.n206 9.3005
R372 source.n205 source.n204 9.3005
R373 source.n190 source.n189 9.3005
R374 source.n199 source.n198 9.3005
R375 source.n197 source.n196 9.3005
R376 source.n173 source.n172 9.3005
R377 source.n146 source.n145 9.3005
R378 source.n167 source.n166 9.3005
R379 source.n165 source.n164 9.3005
R380 source.n150 source.n149 9.3005
R381 source.n159 source.n158 9.3005
R382 source.n157 source.n156 9.3005
R383 source.n29 source.n28 9.3005
R384 source.n2 source.n1 9.3005
R385 source.n23 source.n22 9.3005
R386 source.n21 source.n20 9.3005
R387 source.n6 source.n5 9.3005
R388 source.n15 source.n14 9.3005
R389 source.n13 source.n12 9.3005
R390 source.n69 source.n68 9.3005
R391 source.n42 source.n41 9.3005
R392 source.n63 source.n62 9.3005
R393 source.n61 source.n60 9.3005
R394 source.n46 source.n45 9.3005
R395 source.n55 source.n54 9.3005
R396 source.n53 source.n52 9.3005
R397 source.n101 source.n100 9.3005
R398 source.n74 source.n73 9.3005
R399 source.n95 source.n94 9.3005
R400 source.n93 source.n92 9.3005
R401 source.n78 source.n77 9.3005
R402 source.n87 source.n86 9.3005
R403 source.n85 source.n84 9.3005
R404 source.n141 source.n140 9.3005
R405 source.n114 source.n113 9.3005
R406 source.n135 source.n134 9.3005
R407 source.n133 source.n132 9.3005
R408 source.n118 source.n117 9.3005
R409 source.n127 source.n126 9.3005
R410 source.n125 source.n124 9.3005
R411 source.n283 source.n258 8.92171
R412 source.n243 source.n218 8.92171
R413 source.n211 source.n186 8.92171
R414 source.n171 source.n146 8.92171
R415 source.n27 source.n2 8.92171
R416 source.n67 source.n42 8.92171
R417 source.n99 source.n74 8.92171
R418 source.n139 source.n114 8.92171
R419 source.n284 source.n256 8.14595
R420 source.n244 source.n216 8.14595
R421 source.n212 source.n184 8.14595
R422 source.n172 source.n144 8.14595
R423 source.n28 source.n0 8.14595
R424 source.n68 source.n40 8.14595
R425 source.n100 source.n72 8.14595
R426 source.n140 source.n112 8.14595
R427 source.n286 source.n256 5.81868
R428 source.n246 source.n216 5.81868
R429 source.n214 source.n184 5.81868
R430 source.n174 source.n144 5.81868
R431 source.n30 source.n0 5.81868
R432 source.n70 source.n40 5.81868
R433 source.n102 source.n72 5.81868
R434 source.n142 source.n112 5.81868
R435 source.n288 source.n287 5.7505
R436 source.n284 source.n283 5.04292
R437 source.n244 source.n243 5.04292
R438 source.n212 source.n211 5.04292
R439 source.n172 source.n171 5.04292
R440 source.n28 source.n27 5.04292
R441 source.n68 source.n67 5.04292
R442 source.n100 source.n99 5.04292
R443 source.n140 source.n139 5.04292
R444 source.n269 source.n265 4.38594
R445 source.n229 source.n225 4.38594
R446 source.n197 source.n193 4.38594
R447 source.n157 source.n153 4.38594
R448 source.n13 source.n9 4.38594
R449 source.n53 source.n49 4.38594
R450 source.n85 source.n81 4.38594
R451 source.n125 source.n121 4.38594
R452 source.n280 source.n258 4.26717
R453 source.n240 source.n218 4.26717
R454 source.n208 source.n186 4.26717
R455 source.n168 source.n146 4.26717
R456 source.n24 source.n2 4.26717
R457 source.n64 source.n42 4.26717
R458 source.n96 source.n74 4.26717
R459 source.n136 source.n114 4.26717
R460 source.n279 source.n260 3.49141
R461 source.n239 source.n220 3.49141
R462 source.n207 source.n188 3.49141
R463 source.n167 source.n148 3.49141
R464 source.n23 source.n4 3.49141
R465 source.n63 source.n44 3.49141
R466 source.n95 source.n76 3.49141
R467 source.n135 source.n116 3.49141
R468 source.n254 source.t16 3.3005
R469 source.n254 source.t3 3.3005
R470 source.n252 source.t39 3.3005
R471 source.n252 source.t7 3.3005
R472 source.n250 source.t11 3.3005
R473 source.n250 source.t1 3.3005
R474 source.n248 source.t8 3.3005
R475 source.n248 source.t14 3.3005
R476 source.n182 source.t34 3.3005
R477 source.n182 source.t37 3.3005
R478 source.n180 source.t33 3.3005
R479 source.n180 source.t18 3.3005
R480 source.n178 source.t35 3.3005
R481 source.n178 source.t29 3.3005
R482 source.n176 source.t36 3.3005
R483 source.n176 source.t25 3.3005
R484 source.n32 source.t27 3.3005
R485 source.n32 source.t28 3.3005
R486 source.n34 source.t24 3.3005
R487 source.n34 source.t26 3.3005
R488 source.n36 source.t23 3.3005
R489 source.n36 source.t21 3.3005
R490 source.n38 source.t20 3.3005
R491 source.n38 source.t22 3.3005
R492 source.n104 source.t5 3.3005
R493 source.n104 source.t9 3.3005
R494 source.n106 source.t4 3.3005
R495 source.n106 source.t12 3.3005
R496 source.n108 source.t0 3.3005
R497 source.n108 source.t38 3.3005
R498 source.n110 source.t6 3.3005
R499 source.n110 source.t17 3.3005
R500 source.n276 source.n275 2.71565
R501 source.n236 source.n235 2.71565
R502 source.n204 source.n203 2.71565
R503 source.n164 source.n163 2.71565
R504 source.n20 source.n19 2.71565
R505 source.n60 source.n59 2.71565
R506 source.n92 source.n91 2.71565
R507 source.n132 source.n131 2.71565
R508 source.n272 source.n262 1.93989
R509 source.n232 source.n222 1.93989
R510 source.n200 source.n190 1.93989
R511 source.n160 source.n150 1.93989
R512 source.n16 source.n6 1.93989
R513 source.n56 source.n46 1.93989
R514 source.n88 source.n78 1.93989
R515 source.n128 source.n118 1.93989
R516 source.n271 source.n264 1.16414
R517 source.n231 source.n224 1.16414
R518 source.n199 source.n192 1.16414
R519 source.n159 source.n152 1.16414
R520 source.n15 source.n8 1.16414
R521 source.n55 source.n48 1.16414
R522 source.n87 source.n80 1.16414
R523 source.n127 source.n120 1.16414
R524 source.n143 source.n111 0.974638
R525 source.n111 source.n109 0.974638
R526 source.n109 source.n107 0.974638
R527 source.n107 source.n105 0.974638
R528 source.n105 source.n103 0.974638
R529 source.n71 source.n39 0.974638
R530 source.n39 source.n37 0.974638
R531 source.n37 source.n35 0.974638
R532 source.n35 source.n33 0.974638
R533 source.n33 source.n31 0.974638
R534 source.n177 source.n175 0.974638
R535 source.n179 source.n177 0.974638
R536 source.n181 source.n179 0.974638
R537 source.n183 source.n181 0.974638
R538 source.n215 source.n183 0.974638
R539 source.n249 source.n247 0.974638
R540 source.n251 source.n249 0.974638
R541 source.n253 source.n251 0.974638
R542 source.n255 source.n253 0.974638
R543 source.n287 source.n255 0.974638
R544 source.n103 source.n71 0.470328
R545 source.n247 source.n215 0.470328
R546 source.n268 source.n267 0.388379
R547 source.n228 source.n227 0.388379
R548 source.n196 source.n195 0.388379
R549 source.n156 source.n155 0.388379
R550 source.n12 source.n11 0.388379
R551 source.n52 source.n51 0.388379
R552 source.n84 source.n83 0.388379
R553 source.n124 source.n123 0.388379
R554 source source.n288 0.188
R555 source.n270 source.n269 0.155672
R556 source.n270 source.n261 0.155672
R557 source.n277 source.n261 0.155672
R558 source.n278 source.n277 0.155672
R559 source.n278 source.n257 0.155672
R560 source.n285 source.n257 0.155672
R561 source.n230 source.n229 0.155672
R562 source.n230 source.n221 0.155672
R563 source.n237 source.n221 0.155672
R564 source.n238 source.n237 0.155672
R565 source.n238 source.n217 0.155672
R566 source.n245 source.n217 0.155672
R567 source.n198 source.n197 0.155672
R568 source.n198 source.n189 0.155672
R569 source.n205 source.n189 0.155672
R570 source.n206 source.n205 0.155672
R571 source.n206 source.n185 0.155672
R572 source.n213 source.n185 0.155672
R573 source.n158 source.n157 0.155672
R574 source.n158 source.n149 0.155672
R575 source.n165 source.n149 0.155672
R576 source.n166 source.n165 0.155672
R577 source.n166 source.n145 0.155672
R578 source.n173 source.n145 0.155672
R579 source.n29 source.n1 0.155672
R580 source.n22 source.n1 0.155672
R581 source.n22 source.n21 0.155672
R582 source.n21 source.n5 0.155672
R583 source.n14 source.n5 0.155672
R584 source.n14 source.n13 0.155672
R585 source.n69 source.n41 0.155672
R586 source.n62 source.n41 0.155672
R587 source.n62 source.n61 0.155672
R588 source.n61 source.n45 0.155672
R589 source.n54 source.n45 0.155672
R590 source.n54 source.n53 0.155672
R591 source.n101 source.n73 0.155672
R592 source.n94 source.n73 0.155672
R593 source.n94 source.n93 0.155672
R594 source.n93 source.n77 0.155672
R595 source.n86 source.n77 0.155672
R596 source.n86 source.n85 0.155672
R597 source.n141 source.n113 0.155672
R598 source.n134 source.n113 0.155672
R599 source.n134 source.n133 0.155672
R600 source.n133 source.n117 0.155672
R601 source.n126 source.n117 0.155672
R602 source.n126 source.n125 0.155672
R603 minus.n7 minus.t10 251.644
R604 minus.n37 minus.t9 251.644
R605 minus.n8 minus.t7 229.855
R606 minus.n10 minus.t5 229.855
R607 minus.n5 minus.t13 229.855
R608 minus.n15 minus.t15 229.855
R609 minus.n3 minus.t11 229.855
R610 minus.n21 minus.t8 229.855
R611 minus.n22 minus.t17 229.855
R612 minus.n26 minus.t14 229.855
R613 minus.n28 minus.t2 229.855
R614 minus.n38 minus.t0 229.855
R615 minus.n40 minus.t4 229.855
R616 minus.n35 minus.t19 229.855
R617 minus.n45 minus.t6 229.855
R618 minus.n33 minus.t18 229.855
R619 minus.n51 minus.t1 229.855
R620 minus.n52 minus.t12 229.855
R621 minus.n56 minus.t3 229.855
R622 minus.n58 minus.t16 229.855
R623 minus.n29 minus.n28 161.3
R624 minus.n27 minus.n0 161.3
R625 minus.n26 minus.n25 161.3
R626 minus.n24 minus.n1 161.3
R627 minus.n20 minus.n19 161.3
R628 minus.n18 minus.n3 161.3
R629 minus.n17 minus.n16 161.3
R630 minus.n15 minus.n4 161.3
R631 minus.n14 minus.n13 161.3
R632 minus.n9 minus.n6 161.3
R633 minus.n59 minus.n58 161.3
R634 minus.n57 minus.n30 161.3
R635 minus.n56 minus.n55 161.3
R636 minus.n54 minus.n31 161.3
R637 minus.n50 minus.n49 161.3
R638 minus.n48 minus.n33 161.3
R639 minus.n47 minus.n46 161.3
R640 minus.n45 minus.n34 161.3
R641 minus.n44 minus.n43 161.3
R642 minus.n39 minus.n36 161.3
R643 minus.n23 minus.n22 80.6037
R644 minus.n21 minus.n2 80.6037
R645 minus.n12 minus.n5 80.6037
R646 minus.n11 minus.n10 80.6037
R647 minus.n53 minus.n52 80.6037
R648 minus.n51 minus.n32 80.6037
R649 minus.n42 minus.n35 80.6037
R650 minus.n41 minus.n40 80.6037
R651 minus.n10 minus.n5 48.2005
R652 minus.n22 minus.n21 48.2005
R653 minus.n40 minus.n35 48.2005
R654 minus.n52 minus.n51 48.2005
R655 minus.n7 minus.n6 44.8565
R656 minus.n37 minus.n36 44.8565
R657 minus.n14 minus.n5 43.0884
R658 minus.n21 minus.n20 43.0884
R659 minus.n44 minus.n35 43.0884
R660 minus.n51 minus.n50 43.0884
R661 minus.n10 minus.n9 40.1672
R662 minus.n22 minus.n1 40.1672
R663 minus.n40 minus.n39 40.1672
R664 minus.n52 minus.n31 40.1672
R665 minus.n60 minus.n29 36.9096
R666 minus.n28 minus.n27 27.0217
R667 minus.n58 minus.n57 27.0217
R668 minus.n16 minus.n3 24.1005
R669 minus.n16 minus.n15 24.1005
R670 minus.n46 minus.n45 24.1005
R671 minus.n46 minus.n33 24.1005
R672 minus.n27 minus.n26 21.1793
R673 minus.n57 minus.n56 21.1793
R674 minus.n8 minus.n7 20.1275
R675 minus.n38 minus.n37 20.1275
R676 minus.n9 minus.n8 8.03383
R677 minus.n26 minus.n1 8.03383
R678 minus.n39 minus.n38 8.03383
R679 minus.n56 minus.n31 8.03383
R680 minus.n60 minus.n59 6.70505
R681 minus.n15 minus.n14 5.11262
R682 minus.n20 minus.n3 5.11262
R683 minus.n45 minus.n44 5.11262
R684 minus.n50 minus.n33 5.11262
R685 minus.n23 minus.n2 0.380177
R686 minus.n12 minus.n11 0.380177
R687 minus.n42 minus.n41 0.380177
R688 minus.n53 minus.n32 0.380177
R689 minus.n24 minus.n23 0.285035
R690 minus.n19 minus.n2 0.285035
R691 minus.n13 minus.n12 0.285035
R692 minus.n11 minus.n6 0.285035
R693 minus.n41 minus.n36 0.285035
R694 minus.n43 minus.n42 0.285035
R695 minus.n49 minus.n32 0.285035
R696 minus.n54 minus.n53 0.285035
R697 minus.n29 minus.n0 0.189894
R698 minus.n25 minus.n0 0.189894
R699 minus.n25 minus.n24 0.189894
R700 minus.n19 minus.n18 0.189894
R701 minus.n18 minus.n17 0.189894
R702 minus.n17 minus.n4 0.189894
R703 minus.n13 minus.n4 0.189894
R704 minus.n43 minus.n34 0.189894
R705 minus.n47 minus.n34 0.189894
R706 minus.n48 minus.n47 0.189894
R707 minus.n49 minus.n48 0.189894
R708 minus.n55 minus.n54 0.189894
R709 minus.n55 minus.n30 0.189894
R710 minus.n59 minus.n30 0.189894
R711 minus minus.n60 0.188
R712 drain_right.n6 drain_right.n4 68.1648
R713 drain_right.n2 drain_right.n0 68.1648
R714 drain_right.n10 drain_right.n8 68.1648
R715 drain_right.n10 drain_right.n9 67.1908
R716 drain_right.n12 drain_right.n11 67.1908
R717 drain_right.n14 drain_right.n13 67.1908
R718 drain_right.n16 drain_right.n15 67.1908
R719 drain_right.n7 drain_right.n3 67.1907
R720 drain_right.n6 drain_right.n5 67.1907
R721 drain_right.n2 drain_right.n1 67.1907
R722 drain_right drain_right.n7 30.0615
R723 drain_right drain_right.n16 6.62735
R724 drain_right.n3 drain_right.t13 3.3005
R725 drain_right.n3 drain_right.t1 3.3005
R726 drain_right.n4 drain_right.t16 3.3005
R727 drain_right.n4 drain_right.t3 3.3005
R728 drain_right.n5 drain_right.t18 3.3005
R729 drain_right.n5 drain_right.t7 3.3005
R730 drain_right.n1 drain_right.t15 3.3005
R731 drain_right.n1 drain_right.t0 3.3005
R732 drain_right.n0 drain_right.t10 3.3005
R733 drain_right.n0 drain_right.t19 3.3005
R734 drain_right.n8 drain_right.t12 3.3005
R735 drain_right.n8 drain_right.t9 3.3005
R736 drain_right.n9 drain_right.t6 3.3005
R737 drain_right.n9 drain_right.t14 3.3005
R738 drain_right.n11 drain_right.t8 3.3005
R739 drain_right.n11 drain_right.t4 3.3005
R740 drain_right.n13 drain_right.t2 3.3005
R741 drain_right.n13 drain_right.t11 3.3005
R742 drain_right.n15 drain_right.t17 3.3005
R743 drain_right.n15 drain_right.t5 3.3005
R744 drain_right.n16 drain_right.n14 0.974638
R745 drain_right.n14 drain_right.n12 0.974638
R746 drain_right.n12 drain_right.n10 0.974638
R747 drain_right.n7 drain_right.n6 0.919292
R748 drain_right.n7 drain_right.n2 0.919292
C0 source drain_left 13.4091f
C1 plus drain_right 0.478206f
C2 drain_right minus 7.12407f
C3 drain_right drain_left 1.72917f
C4 plus minus 6.02719f
C5 plus drain_left 7.44451f
C6 minus drain_left 0.17405f
C7 drain_right source 13.412f
C8 plus source 7.73958f
C9 minus source 7.72556f
C10 drain_right a_n3202_n2088# 6.39501f
C11 drain_left a_n3202_n2088# 6.84478f
C12 source a_n3202_n2088# 5.908512f
C13 minus a_n3202_n2088# 12.388208f
C14 plus a_n3202_n2088# 13.90121f
C15 drain_right.t10 a_n3202_n2088# 0.125175f
C16 drain_right.t19 a_n3202_n2088# 0.125175f
C17 drain_right.n0 a_n3202_n2088# 1.04954f
C18 drain_right.t15 a_n3202_n2088# 0.125175f
C19 drain_right.t0 a_n3202_n2088# 0.125175f
C20 drain_right.n1 a_n3202_n2088# 1.04396f
C21 drain_right.n2 a_n3202_n2088# 0.761035f
C22 drain_right.t13 a_n3202_n2088# 0.125175f
C23 drain_right.t1 a_n3202_n2088# 0.125175f
C24 drain_right.n3 a_n3202_n2088# 1.04396f
C25 drain_right.t16 a_n3202_n2088# 0.125175f
C26 drain_right.t3 a_n3202_n2088# 0.125175f
C27 drain_right.n4 a_n3202_n2088# 1.04954f
C28 drain_right.t18 a_n3202_n2088# 0.125175f
C29 drain_right.t7 a_n3202_n2088# 0.125175f
C30 drain_right.n5 a_n3202_n2088# 1.04396f
C31 drain_right.n6 a_n3202_n2088# 0.761035f
C32 drain_right.n7 a_n3202_n2088# 1.59122f
C33 drain_right.t12 a_n3202_n2088# 0.125175f
C34 drain_right.t9 a_n3202_n2088# 0.125175f
C35 drain_right.n8 a_n3202_n2088# 1.04954f
C36 drain_right.t6 a_n3202_n2088# 0.125175f
C37 drain_right.t14 a_n3202_n2088# 0.125175f
C38 drain_right.n9 a_n3202_n2088# 1.04397f
C39 drain_right.n10 a_n3202_n2088# 0.765072f
C40 drain_right.t8 a_n3202_n2088# 0.125175f
C41 drain_right.t4 a_n3202_n2088# 0.125175f
C42 drain_right.n11 a_n3202_n2088# 1.04397f
C43 drain_right.n12 a_n3202_n2088# 0.380008f
C44 drain_right.t2 a_n3202_n2088# 0.125175f
C45 drain_right.t11 a_n3202_n2088# 0.125175f
C46 drain_right.n13 a_n3202_n2088# 1.04397f
C47 drain_right.n14 a_n3202_n2088# 0.380008f
C48 drain_right.t17 a_n3202_n2088# 0.125175f
C49 drain_right.t5 a_n3202_n2088# 0.125175f
C50 drain_right.n15 a_n3202_n2088# 1.04397f
C51 drain_right.n16 a_n3202_n2088# 0.61674f
C52 minus.n0 a_n3202_n2088# 0.038539f
C53 minus.n1 a_n3202_n2088# 0.008745f
C54 minus.t14 a_n3202_n2088# 0.536567f
C55 minus.n2 a_n3202_n2088# 0.064192f
C56 minus.t11 a_n3202_n2088# 0.536567f
C57 minus.n3 a_n3202_n2088# 0.244418f
C58 minus.n4 a_n3202_n2088# 0.038539f
C59 minus.t13 a_n3202_n2088# 0.536567f
C60 minus.n5 a_n3202_n2088# 0.255421f
C61 minus.n6 a_n3202_n2088# 0.177394f
C62 minus.t10 a_n3202_n2088# 0.557918f
C63 minus.n7 a_n3202_n2088# 0.229033f
C64 minus.t7 a_n3202_n2088# 0.536567f
C65 minus.n8 a_n3202_n2088# 0.247658f
C66 minus.n9 a_n3202_n2088# 0.008745f
C67 minus.t5 a_n3202_n2088# 0.536567f
C68 minus.n10 a_n3202_n2088# 0.254946f
C69 minus.n11 a_n3202_n2088# 0.064192f
C70 minus.n12 a_n3202_n2088# 0.064192f
C71 minus.n13 a_n3202_n2088# 0.051426f
C72 minus.n14 a_n3202_n2088# 0.008745f
C73 minus.t15 a_n3202_n2088# 0.536567f
C74 minus.n15 a_n3202_n2088# 0.244418f
C75 minus.n16 a_n3202_n2088# 0.008745f
C76 minus.n17 a_n3202_n2088# 0.038539f
C77 minus.n18 a_n3202_n2088# 0.038539f
C78 minus.n19 a_n3202_n2088# 0.051426f
C79 minus.n20 a_n3202_n2088# 0.008745f
C80 minus.t8 a_n3202_n2088# 0.536567f
C81 minus.n21 a_n3202_n2088# 0.255421f
C82 minus.t17 a_n3202_n2088# 0.536567f
C83 minus.n22 a_n3202_n2088# 0.254946f
C84 minus.n23 a_n3202_n2088# 0.064192f
C85 minus.n24 a_n3202_n2088# 0.051426f
C86 minus.n25 a_n3202_n2088# 0.038539f
C87 minus.n26 a_n3202_n2088# 0.244418f
C88 minus.n27 a_n3202_n2088# 0.008745f
C89 minus.t2 a_n3202_n2088# 0.536567f
C90 minus.n28 a_n3202_n2088# 0.244062f
C91 minus.n29 a_n3202_n2088# 1.41016f
C92 minus.n30 a_n3202_n2088# 0.038539f
C93 minus.n31 a_n3202_n2088# 0.008745f
C94 minus.n32 a_n3202_n2088# 0.064192f
C95 minus.t18 a_n3202_n2088# 0.536567f
C96 minus.n33 a_n3202_n2088# 0.244418f
C97 minus.n34 a_n3202_n2088# 0.038539f
C98 minus.t19 a_n3202_n2088# 0.536567f
C99 minus.n35 a_n3202_n2088# 0.255421f
C100 minus.n36 a_n3202_n2088# 0.177394f
C101 minus.t9 a_n3202_n2088# 0.557918f
C102 minus.n37 a_n3202_n2088# 0.229033f
C103 minus.t0 a_n3202_n2088# 0.536567f
C104 minus.n38 a_n3202_n2088# 0.247658f
C105 minus.n39 a_n3202_n2088# 0.008745f
C106 minus.t4 a_n3202_n2088# 0.536567f
C107 minus.n40 a_n3202_n2088# 0.254946f
C108 minus.n41 a_n3202_n2088# 0.064192f
C109 minus.n42 a_n3202_n2088# 0.064192f
C110 minus.n43 a_n3202_n2088# 0.051426f
C111 minus.n44 a_n3202_n2088# 0.008745f
C112 minus.t6 a_n3202_n2088# 0.536567f
C113 minus.n45 a_n3202_n2088# 0.244418f
C114 minus.n46 a_n3202_n2088# 0.008745f
C115 minus.n47 a_n3202_n2088# 0.038539f
C116 minus.n48 a_n3202_n2088# 0.038539f
C117 minus.n49 a_n3202_n2088# 0.051426f
C118 minus.n50 a_n3202_n2088# 0.008745f
C119 minus.t1 a_n3202_n2088# 0.536567f
C120 minus.n51 a_n3202_n2088# 0.255421f
C121 minus.t12 a_n3202_n2088# 0.536567f
C122 minus.n52 a_n3202_n2088# 0.254946f
C123 minus.n53 a_n3202_n2088# 0.064192f
C124 minus.n54 a_n3202_n2088# 0.051426f
C125 minus.n55 a_n3202_n2088# 0.038539f
C126 minus.t3 a_n3202_n2088# 0.536567f
C127 minus.n56 a_n3202_n2088# 0.244418f
C128 minus.n57 a_n3202_n2088# 0.008745f
C129 minus.t16 a_n3202_n2088# 0.536567f
C130 minus.n58 a_n3202_n2088# 0.244062f
C131 minus.n59 a_n3202_n2088# 0.2704f
C132 minus.n60 a_n3202_n2088# 1.7034f
C133 source.n0 a_n3202_n2088# 0.036082f
C134 source.n1 a_n3202_n2088# 0.025671f
C135 source.n2 a_n3202_n2088# 0.013794f
C136 source.n3 a_n3202_n2088# 0.032604f
C137 source.n4 a_n3202_n2088# 0.014606f
C138 source.n5 a_n3202_n2088# 0.025671f
C139 source.n6 a_n3202_n2088# 0.013794f
C140 source.n7 a_n3202_n2088# 0.032604f
C141 source.n8 a_n3202_n2088# 0.014606f
C142 source.n9 a_n3202_n2088# 0.109852f
C143 source.t30 a_n3202_n2088# 0.053141f
C144 source.n10 a_n3202_n2088# 0.024453f
C145 source.n11 a_n3202_n2088# 0.019259f
C146 source.n12 a_n3202_n2088# 0.013794f
C147 source.n13 a_n3202_n2088# 0.610805f
C148 source.n14 a_n3202_n2088# 0.025671f
C149 source.n15 a_n3202_n2088# 0.013794f
C150 source.n16 a_n3202_n2088# 0.014606f
C151 source.n17 a_n3202_n2088# 0.032604f
C152 source.n18 a_n3202_n2088# 0.032604f
C153 source.n19 a_n3202_n2088# 0.014606f
C154 source.n20 a_n3202_n2088# 0.013794f
C155 source.n21 a_n3202_n2088# 0.025671f
C156 source.n22 a_n3202_n2088# 0.025671f
C157 source.n23 a_n3202_n2088# 0.013794f
C158 source.n24 a_n3202_n2088# 0.014606f
C159 source.n25 a_n3202_n2088# 0.032604f
C160 source.n26 a_n3202_n2088# 0.070583f
C161 source.n27 a_n3202_n2088# 0.014606f
C162 source.n28 a_n3202_n2088# 0.013794f
C163 source.n29 a_n3202_n2088# 0.059336f
C164 source.n30 a_n3202_n2088# 0.039494f
C165 source.n31 a_n3202_n2088# 0.682782f
C166 source.t27 a_n3202_n2088# 0.121714f
C167 source.t28 a_n3202_n2088# 0.121714f
C168 source.n32 a_n3202_n2088# 0.947916f
C169 source.n33 a_n3202_n2088# 0.40179f
C170 source.t24 a_n3202_n2088# 0.121714f
C171 source.t26 a_n3202_n2088# 0.121714f
C172 source.n34 a_n3202_n2088# 0.947916f
C173 source.n35 a_n3202_n2088# 0.40179f
C174 source.t23 a_n3202_n2088# 0.121714f
C175 source.t21 a_n3202_n2088# 0.121714f
C176 source.n36 a_n3202_n2088# 0.947916f
C177 source.n37 a_n3202_n2088# 0.40179f
C178 source.t20 a_n3202_n2088# 0.121714f
C179 source.t22 a_n3202_n2088# 0.121714f
C180 source.n38 a_n3202_n2088# 0.947916f
C181 source.n39 a_n3202_n2088# 0.40179f
C182 source.n40 a_n3202_n2088# 0.036082f
C183 source.n41 a_n3202_n2088# 0.025671f
C184 source.n42 a_n3202_n2088# 0.013794f
C185 source.n43 a_n3202_n2088# 0.032604f
C186 source.n44 a_n3202_n2088# 0.014606f
C187 source.n45 a_n3202_n2088# 0.025671f
C188 source.n46 a_n3202_n2088# 0.013794f
C189 source.n47 a_n3202_n2088# 0.032604f
C190 source.n48 a_n3202_n2088# 0.014606f
C191 source.n49 a_n3202_n2088# 0.109852f
C192 source.t19 a_n3202_n2088# 0.053141f
C193 source.n50 a_n3202_n2088# 0.024453f
C194 source.n51 a_n3202_n2088# 0.019259f
C195 source.n52 a_n3202_n2088# 0.013794f
C196 source.n53 a_n3202_n2088# 0.610805f
C197 source.n54 a_n3202_n2088# 0.025671f
C198 source.n55 a_n3202_n2088# 0.013794f
C199 source.n56 a_n3202_n2088# 0.014606f
C200 source.n57 a_n3202_n2088# 0.032604f
C201 source.n58 a_n3202_n2088# 0.032604f
C202 source.n59 a_n3202_n2088# 0.014606f
C203 source.n60 a_n3202_n2088# 0.013794f
C204 source.n61 a_n3202_n2088# 0.025671f
C205 source.n62 a_n3202_n2088# 0.025671f
C206 source.n63 a_n3202_n2088# 0.013794f
C207 source.n64 a_n3202_n2088# 0.014606f
C208 source.n65 a_n3202_n2088# 0.032604f
C209 source.n66 a_n3202_n2088# 0.070583f
C210 source.n67 a_n3202_n2088# 0.014606f
C211 source.n68 a_n3202_n2088# 0.013794f
C212 source.n69 a_n3202_n2088# 0.059336f
C213 source.n70 a_n3202_n2088# 0.039494f
C214 source.n71 a_n3202_n2088# 0.141364f
C215 source.n72 a_n3202_n2088# 0.036082f
C216 source.n73 a_n3202_n2088# 0.025671f
C217 source.n74 a_n3202_n2088# 0.013794f
C218 source.n75 a_n3202_n2088# 0.032604f
C219 source.n76 a_n3202_n2088# 0.014606f
C220 source.n77 a_n3202_n2088# 0.025671f
C221 source.n78 a_n3202_n2088# 0.013794f
C222 source.n79 a_n3202_n2088# 0.032604f
C223 source.n80 a_n3202_n2088# 0.014606f
C224 source.n81 a_n3202_n2088# 0.109852f
C225 source.t2 a_n3202_n2088# 0.053141f
C226 source.n82 a_n3202_n2088# 0.024453f
C227 source.n83 a_n3202_n2088# 0.019259f
C228 source.n84 a_n3202_n2088# 0.013794f
C229 source.n85 a_n3202_n2088# 0.610805f
C230 source.n86 a_n3202_n2088# 0.025671f
C231 source.n87 a_n3202_n2088# 0.013794f
C232 source.n88 a_n3202_n2088# 0.014606f
C233 source.n89 a_n3202_n2088# 0.032604f
C234 source.n90 a_n3202_n2088# 0.032604f
C235 source.n91 a_n3202_n2088# 0.014606f
C236 source.n92 a_n3202_n2088# 0.013794f
C237 source.n93 a_n3202_n2088# 0.025671f
C238 source.n94 a_n3202_n2088# 0.025671f
C239 source.n95 a_n3202_n2088# 0.013794f
C240 source.n96 a_n3202_n2088# 0.014606f
C241 source.n97 a_n3202_n2088# 0.032604f
C242 source.n98 a_n3202_n2088# 0.070583f
C243 source.n99 a_n3202_n2088# 0.014606f
C244 source.n100 a_n3202_n2088# 0.013794f
C245 source.n101 a_n3202_n2088# 0.059336f
C246 source.n102 a_n3202_n2088# 0.039494f
C247 source.n103 a_n3202_n2088# 0.141364f
C248 source.t5 a_n3202_n2088# 0.121714f
C249 source.t9 a_n3202_n2088# 0.121714f
C250 source.n104 a_n3202_n2088# 0.947916f
C251 source.n105 a_n3202_n2088# 0.40179f
C252 source.t4 a_n3202_n2088# 0.121714f
C253 source.t12 a_n3202_n2088# 0.121714f
C254 source.n106 a_n3202_n2088# 0.947916f
C255 source.n107 a_n3202_n2088# 0.40179f
C256 source.t0 a_n3202_n2088# 0.121714f
C257 source.t38 a_n3202_n2088# 0.121714f
C258 source.n108 a_n3202_n2088# 0.947916f
C259 source.n109 a_n3202_n2088# 0.40179f
C260 source.t6 a_n3202_n2088# 0.121714f
C261 source.t17 a_n3202_n2088# 0.121714f
C262 source.n110 a_n3202_n2088# 0.947916f
C263 source.n111 a_n3202_n2088# 0.40179f
C264 source.n112 a_n3202_n2088# 0.036082f
C265 source.n113 a_n3202_n2088# 0.025671f
C266 source.n114 a_n3202_n2088# 0.013794f
C267 source.n115 a_n3202_n2088# 0.032604f
C268 source.n116 a_n3202_n2088# 0.014606f
C269 source.n117 a_n3202_n2088# 0.025671f
C270 source.n118 a_n3202_n2088# 0.013794f
C271 source.n119 a_n3202_n2088# 0.032604f
C272 source.n120 a_n3202_n2088# 0.014606f
C273 source.n121 a_n3202_n2088# 0.109852f
C274 source.t13 a_n3202_n2088# 0.053141f
C275 source.n122 a_n3202_n2088# 0.024453f
C276 source.n123 a_n3202_n2088# 0.019259f
C277 source.n124 a_n3202_n2088# 0.013794f
C278 source.n125 a_n3202_n2088# 0.610805f
C279 source.n126 a_n3202_n2088# 0.025671f
C280 source.n127 a_n3202_n2088# 0.013794f
C281 source.n128 a_n3202_n2088# 0.014606f
C282 source.n129 a_n3202_n2088# 0.032604f
C283 source.n130 a_n3202_n2088# 0.032604f
C284 source.n131 a_n3202_n2088# 0.014606f
C285 source.n132 a_n3202_n2088# 0.013794f
C286 source.n133 a_n3202_n2088# 0.025671f
C287 source.n134 a_n3202_n2088# 0.025671f
C288 source.n135 a_n3202_n2088# 0.013794f
C289 source.n136 a_n3202_n2088# 0.014606f
C290 source.n137 a_n3202_n2088# 0.032604f
C291 source.n138 a_n3202_n2088# 0.070583f
C292 source.n139 a_n3202_n2088# 0.014606f
C293 source.n140 a_n3202_n2088# 0.013794f
C294 source.n141 a_n3202_n2088# 0.059336f
C295 source.n142 a_n3202_n2088# 0.039494f
C296 source.n143 a_n3202_n2088# 1.02358f
C297 source.n144 a_n3202_n2088# 0.036082f
C298 source.n145 a_n3202_n2088# 0.025671f
C299 source.n146 a_n3202_n2088# 0.013794f
C300 source.n147 a_n3202_n2088# 0.032604f
C301 source.n148 a_n3202_n2088# 0.014606f
C302 source.n149 a_n3202_n2088# 0.025671f
C303 source.n150 a_n3202_n2088# 0.013794f
C304 source.n151 a_n3202_n2088# 0.032604f
C305 source.n152 a_n3202_n2088# 0.014606f
C306 source.n153 a_n3202_n2088# 0.109852f
C307 source.t32 a_n3202_n2088# 0.053141f
C308 source.n154 a_n3202_n2088# 0.024453f
C309 source.n155 a_n3202_n2088# 0.019259f
C310 source.n156 a_n3202_n2088# 0.013794f
C311 source.n157 a_n3202_n2088# 0.610805f
C312 source.n158 a_n3202_n2088# 0.025671f
C313 source.n159 a_n3202_n2088# 0.013794f
C314 source.n160 a_n3202_n2088# 0.014606f
C315 source.n161 a_n3202_n2088# 0.032604f
C316 source.n162 a_n3202_n2088# 0.032604f
C317 source.n163 a_n3202_n2088# 0.014606f
C318 source.n164 a_n3202_n2088# 0.013794f
C319 source.n165 a_n3202_n2088# 0.025671f
C320 source.n166 a_n3202_n2088# 0.025671f
C321 source.n167 a_n3202_n2088# 0.013794f
C322 source.n168 a_n3202_n2088# 0.014606f
C323 source.n169 a_n3202_n2088# 0.032604f
C324 source.n170 a_n3202_n2088# 0.070583f
C325 source.n171 a_n3202_n2088# 0.014606f
C326 source.n172 a_n3202_n2088# 0.013794f
C327 source.n173 a_n3202_n2088# 0.059336f
C328 source.n174 a_n3202_n2088# 0.039494f
C329 source.n175 a_n3202_n2088# 1.02358f
C330 source.t36 a_n3202_n2088# 0.121714f
C331 source.t25 a_n3202_n2088# 0.121714f
C332 source.n176 a_n3202_n2088# 0.94791f
C333 source.n177 a_n3202_n2088# 0.401797f
C334 source.t35 a_n3202_n2088# 0.121714f
C335 source.t29 a_n3202_n2088# 0.121714f
C336 source.n178 a_n3202_n2088# 0.94791f
C337 source.n179 a_n3202_n2088# 0.401797f
C338 source.t33 a_n3202_n2088# 0.121714f
C339 source.t18 a_n3202_n2088# 0.121714f
C340 source.n180 a_n3202_n2088# 0.94791f
C341 source.n181 a_n3202_n2088# 0.401797f
C342 source.t34 a_n3202_n2088# 0.121714f
C343 source.t37 a_n3202_n2088# 0.121714f
C344 source.n182 a_n3202_n2088# 0.94791f
C345 source.n183 a_n3202_n2088# 0.401797f
C346 source.n184 a_n3202_n2088# 0.036082f
C347 source.n185 a_n3202_n2088# 0.025671f
C348 source.n186 a_n3202_n2088# 0.013794f
C349 source.n187 a_n3202_n2088# 0.032604f
C350 source.n188 a_n3202_n2088# 0.014606f
C351 source.n189 a_n3202_n2088# 0.025671f
C352 source.n190 a_n3202_n2088# 0.013794f
C353 source.n191 a_n3202_n2088# 0.032604f
C354 source.n192 a_n3202_n2088# 0.014606f
C355 source.n193 a_n3202_n2088# 0.109852f
C356 source.t31 a_n3202_n2088# 0.053141f
C357 source.n194 a_n3202_n2088# 0.024453f
C358 source.n195 a_n3202_n2088# 0.019259f
C359 source.n196 a_n3202_n2088# 0.013794f
C360 source.n197 a_n3202_n2088# 0.610805f
C361 source.n198 a_n3202_n2088# 0.025671f
C362 source.n199 a_n3202_n2088# 0.013794f
C363 source.n200 a_n3202_n2088# 0.014606f
C364 source.n201 a_n3202_n2088# 0.032604f
C365 source.n202 a_n3202_n2088# 0.032604f
C366 source.n203 a_n3202_n2088# 0.014606f
C367 source.n204 a_n3202_n2088# 0.013794f
C368 source.n205 a_n3202_n2088# 0.025671f
C369 source.n206 a_n3202_n2088# 0.025671f
C370 source.n207 a_n3202_n2088# 0.013794f
C371 source.n208 a_n3202_n2088# 0.014606f
C372 source.n209 a_n3202_n2088# 0.032604f
C373 source.n210 a_n3202_n2088# 0.070583f
C374 source.n211 a_n3202_n2088# 0.014606f
C375 source.n212 a_n3202_n2088# 0.013794f
C376 source.n213 a_n3202_n2088# 0.059336f
C377 source.n214 a_n3202_n2088# 0.039494f
C378 source.n215 a_n3202_n2088# 0.141364f
C379 source.n216 a_n3202_n2088# 0.036082f
C380 source.n217 a_n3202_n2088# 0.025671f
C381 source.n218 a_n3202_n2088# 0.013794f
C382 source.n219 a_n3202_n2088# 0.032604f
C383 source.n220 a_n3202_n2088# 0.014606f
C384 source.n221 a_n3202_n2088# 0.025671f
C385 source.n222 a_n3202_n2088# 0.013794f
C386 source.n223 a_n3202_n2088# 0.032604f
C387 source.n224 a_n3202_n2088# 0.014606f
C388 source.n225 a_n3202_n2088# 0.109852f
C389 source.t15 a_n3202_n2088# 0.053141f
C390 source.n226 a_n3202_n2088# 0.024453f
C391 source.n227 a_n3202_n2088# 0.019259f
C392 source.n228 a_n3202_n2088# 0.013794f
C393 source.n229 a_n3202_n2088# 0.610805f
C394 source.n230 a_n3202_n2088# 0.025671f
C395 source.n231 a_n3202_n2088# 0.013794f
C396 source.n232 a_n3202_n2088# 0.014606f
C397 source.n233 a_n3202_n2088# 0.032604f
C398 source.n234 a_n3202_n2088# 0.032604f
C399 source.n235 a_n3202_n2088# 0.014606f
C400 source.n236 a_n3202_n2088# 0.013794f
C401 source.n237 a_n3202_n2088# 0.025671f
C402 source.n238 a_n3202_n2088# 0.025671f
C403 source.n239 a_n3202_n2088# 0.013794f
C404 source.n240 a_n3202_n2088# 0.014606f
C405 source.n241 a_n3202_n2088# 0.032604f
C406 source.n242 a_n3202_n2088# 0.070583f
C407 source.n243 a_n3202_n2088# 0.014606f
C408 source.n244 a_n3202_n2088# 0.013794f
C409 source.n245 a_n3202_n2088# 0.059336f
C410 source.n246 a_n3202_n2088# 0.039494f
C411 source.n247 a_n3202_n2088# 0.141364f
C412 source.t8 a_n3202_n2088# 0.121714f
C413 source.t14 a_n3202_n2088# 0.121714f
C414 source.n248 a_n3202_n2088# 0.94791f
C415 source.n249 a_n3202_n2088# 0.401797f
C416 source.t11 a_n3202_n2088# 0.121714f
C417 source.t1 a_n3202_n2088# 0.121714f
C418 source.n250 a_n3202_n2088# 0.94791f
C419 source.n251 a_n3202_n2088# 0.401797f
C420 source.t39 a_n3202_n2088# 0.121714f
C421 source.t7 a_n3202_n2088# 0.121714f
C422 source.n252 a_n3202_n2088# 0.94791f
C423 source.n253 a_n3202_n2088# 0.401797f
C424 source.t16 a_n3202_n2088# 0.121714f
C425 source.t3 a_n3202_n2088# 0.121714f
C426 source.n254 a_n3202_n2088# 0.94791f
C427 source.n255 a_n3202_n2088# 0.401797f
C428 source.n256 a_n3202_n2088# 0.036082f
C429 source.n257 a_n3202_n2088# 0.025671f
C430 source.n258 a_n3202_n2088# 0.013794f
C431 source.n259 a_n3202_n2088# 0.032604f
C432 source.n260 a_n3202_n2088# 0.014606f
C433 source.n261 a_n3202_n2088# 0.025671f
C434 source.n262 a_n3202_n2088# 0.013794f
C435 source.n263 a_n3202_n2088# 0.032604f
C436 source.n264 a_n3202_n2088# 0.014606f
C437 source.n265 a_n3202_n2088# 0.109852f
C438 source.t10 a_n3202_n2088# 0.053141f
C439 source.n266 a_n3202_n2088# 0.024453f
C440 source.n267 a_n3202_n2088# 0.019259f
C441 source.n268 a_n3202_n2088# 0.013794f
C442 source.n269 a_n3202_n2088# 0.610805f
C443 source.n270 a_n3202_n2088# 0.025671f
C444 source.n271 a_n3202_n2088# 0.013794f
C445 source.n272 a_n3202_n2088# 0.014606f
C446 source.n273 a_n3202_n2088# 0.032604f
C447 source.n274 a_n3202_n2088# 0.032604f
C448 source.n275 a_n3202_n2088# 0.014606f
C449 source.n276 a_n3202_n2088# 0.013794f
C450 source.n277 a_n3202_n2088# 0.025671f
C451 source.n278 a_n3202_n2088# 0.025671f
C452 source.n279 a_n3202_n2088# 0.013794f
C453 source.n280 a_n3202_n2088# 0.014606f
C454 source.n281 a_n3202_n2088# 0.032604f
C455 source.n282 a_n3202_n2088# 0.070583f
C456 source.n283 a_n3202_n2088# 0.014606f
C457 source.n284 a_n3202_n2088# 0.013794f
C458 source.n285 a_n3202_n2088# 0.059336f
C459 source.n286 a_n3202_n2088# 0.039494f
C460 source.n287 a_n3202_n2088# 0.314371f
C461 source.n288 a_n3202_n2088# 1.06826f
C462 drain_left.t8 a_n3202_n2088# 0.12637f
C463 drain_left.t11 a_n3202_n2088# 0.12637f
C464 drain_left.n0 a_n3202_n2088# 1.05957f
C465 drain_left.t4 a_n3202_n2088# 0.12637f
C466 drain_left.t9 a_n3202_n2088# 0.12637f
C467 drain_left.n1 a_n3202_n2088# 1.05393f
C468 drain_left.n2 a_n3202_n2088# 0.768302f
C469 drain_left.t0 a_n3202_n2088# 0.12637f
C470 drain_left.t7 a_n3202_n2088# 0.12637f
C471 drain_left.n3 a_n3202_n2088# 1.05393f
C472 drain_left.t2 a_n3202_n2088# 0.12637f
C473 drain_left.t3 a_n3202_n2088# 0.12637f
C474 drain_left.n4 a_n3202_n2088# 1.05957f
C475 drain_left.t13 a_n3202_n2088# 0.12637f
C476 drain_left.t12 a_n3202_n2088# 0.12637f
C477 drain_left.n5 a_n3202_n2088# 1.05393f
C478 drain_left.n6 a_n3202_n2088# 0.768302f
C479 drain_left.n7 a_n3202_n2088# 1.65945f
C480 drain_left.t10 a_n3202_n2088# 0.12637f
C481 drain_left.t19 a_n3202_n2088# 0.12637f
C482 drain_left.n8 a_n3202_n2088# 1.05957f
C483 drain_left.t16 a_n3202_n2088# 0.12637f
C484 drain_left.t17 a_n3202_n2088# 0.12637f
C485 drain_left.n9 a_n3202_n2088# 1.05393f
C486 drain_left.n10 a_n3202_n2088# 0.772373f
C487 drain_left.t6 a_n3202_n2088# 0.12637f
C488 drain_left.t18 a_n3202_n2088# 0.12637f
C489 drain_left.n11 a_n3202_n2088# 1.05393f
C490 drain_left.n12 a_n3202_n2088# 0.383637f
C491 drain_left.t5 a_n3202_n2088# 0.12637f
C492 drain_left.t15 a_n3202_n2088# 0.12637f
C493 drain_left.n13 a_n3202_n2088# 1.05393f
C494 drain_left.n14 a_n3202_n2088# 0.383637f
C495 drain_left.t14 a_n3202_n2088# 0.12637f
C496 drain_left.t1 a_n3202_n2088# 0.12637f
C497 drain_left.n15 a_n3202_n2088# 1.05393f
C498 drain_left.n16 a_n3202_n2088# 0.622634f
C499 plus.n0 a_n3202_n2088# 0.039242f
C500 plus.t7 a_n3202_n2088# 0.546353f
C501 plus.t9 a_n3202_n2088# 0.546353f
C502 plus.n1 a_n3202_n2088# 0.039242f
C503 plus.t10 a_n3202_n2088# 0.546353f
C504 plus.n2 a_n3202_n2088# 0.259596f
C505 plus.n3 a_n3202_n2088# 0.052363f
C506 plus.t11 a_n3202_n2088# 0.546353f
C507 plus.t13 a_n3202_n2088# 0.546353f
C508 plus.n4 a_n3202_n2088# 0.039242f
C509 plus.t16 a_n3202_n2088# 0.546353f
C510 plus.n5 a_n3202_n2088# 0.248876f
C511 plus.n6 a_n3202_n2088# 0.065362f
C512 plus.t14 a_n3202_n2088# 0.546353f
C513 plus.t15 a_n3202_n2088# 0.546353f
C514 plus.n7 a_n3202_n2088# 0.065362f
C515 plus.t17 a_n3202_n2088# 0.546353f
C516 plus.n8 a_n3202_n2088# 0.252175f
C517 plus.t18 a_n3202_n2088# 0.568093f
C518 plus.n9 a_n3202_n2088# 0.23321f
C519 plus.n10 a_n3202_n2088# 0.18063f
C520 plus.n11 a_n3202_n2088# 0.008905f
C521 plus.n12 a_n3202_n2088# 0.259596f
C522 plus.n13 a_n3202_n2088# 0.26008f
C523 plus.n14 a_n3202_n2088# 0.008905f
C524 plus.n15 a_n3202_n2088# 0.052363f
C525 plus.n16 a_n3202_n2088# 0.039242f
C526 plus.n17 a_n3202_n2088# 0.039242f
C527 plus.n18 a_n3202_n2088# 0.008905f
C528 plus.n19 a_n3202_n2088# 0.248876f
C529 plus.n20 a_n3202_n2088# 0.008905f
C530 plus.n21 a_n3202_n2088# 0.26008f
C531 plus.n22 a_n3202_n2088# 0.065362f
C532 plus.n23 a_n3202_n2088# 0.065362f
C533 plus.n24 a_n3202_n2088# 0.052363f
C534 plus.n25 a_n3202_n2088# 0.008905f
C535 plus.n26 a_n3202_n2088# 0.248876f
C536 plus.n27 a_n3202_n2088# 0.008905f
C537 plus.n28 a_n3202_n2088# 0.248513f
C538 plus.n29 a_n3202_n2088# 0.355899f
C539 plus.n30 a_n3202_n2088# 0.039242f
C540 plus.t5 a_n3202_n2088# 0.546353f
C541 plus.n31 a_n3202_n2088# 0.039242f
C542 plus.t1 a_n3202_n2088# 0.546353f
C543 plus.t12 a_n3202_n2088# 0.546353f
C544 plus.n32 a_n3202_n2088# 0.259596f
C545 plus.n33 a_n3202_n2088# 0.052363f
C546 plus.t2 a_n3202_n2088# 0.546353f
C547 plus.n34 a_n3202_n2088# 0.039242f
C548 plus.t8 a_n3202_n2088# 0.546353f
C549 plus.t4 a_n3202_n2088# 0.546353f
C550 plus.n35 a_n3202_n2088# 0.248876f
C551 plus.n36 a_n3202_n2088# 0.065362f
C552 plus.t19 a_n3202_n2088# 0.546353f
C553 plus.n37 a_n3202_n2088# 0.065362f
C554 plus.t3 a_n3202_n2088# 0.546353f
C555 plus.t0 a_n3202_n2088# 0.546353f
C556 plus.n38 a_n3202_n2088# 0.252175f
C557 plus.t6 a_n3202_n2088# 0.568093f
C558 plus.n39 a_n3202_n2088# 0.23321f
C559 plus.n40 a_n3202_n2088# 0.18063f
C560 plus.n41 a_n3202_n2088# 0.008905f
C561 plus.n42 a_n3202_n2088# 0.259596f
C562 plus.n43 a_n3202_n2088# 0.26008f
C563 plus.n44 a_n3202_n2088# 0.008905f
C564 plus.n45 a_n3202_n2088# 0.052363f
C565 plus.n46 a_n3202_n2088# 0.039242f
C566 plus.n47 a_n3202_n2088# 0.039242f
C567 plus.n48 a_n3202_n2088# 0.008905f
C568 plus.n49 a_n3202_n2088# 0.248876f
C569 plus.n50 a_n3202_n2088# 0.008905f
C570 plus.n51 a_n3202_n2088# 0.26008f
C571 plus.n52 a_n3202_n2088# 0.065362f
C572 plus.n53 a_n3202_n2088# 0.065362f
C573 plus.n54 a_n3202_n2088# 0.052363f
C574 plus.n55 a_n3202_n2088# 0.008905f
C575 plus.n56 a_n3202_n2088# 0.248876f
C576 plus.n57 a_n3202_n2088# 0.008905f
C577 plus.n58 a_n3202_n2088# 0.248513f
C578 plus.n59 a_n3202_n2088# 1.30397f
.ends

