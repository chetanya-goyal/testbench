* NGSPICE file created from diffpair537.ext - technology: sky130A

.subckt diffpair537 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t31 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X1 drain_left.t15 plus.t0 source.t3 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X2 source.t9 plus.t1 drain_left.t14 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X3 drain_left.t13 plus.t2 source.t14 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X4 source.t2 plus.t3 drain_left.t12 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X5 source.t13 plus.t4 drain_left.t11 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X6 drain_left.t10 plus.t5 source.t4 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X7 source.t22 minus.t1 drain_right.t14 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X8 drain_right.t13 minus.t2 source.t16 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X9 drain_right.t12 minus.t3 source.t17 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X10 drain_right.t11 minus.t4 source.t24 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X11 source.t28 minus.t5 drain_right.t10 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X12 drain_left.t9 plus.t6 source.t15 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X13 source.t21 minus.t6 drain_right.t9 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X14 drain_right.t8 minus.t7 source.t27 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X15 source.t1 plus.t7 drain_left.t8 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X16 a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.6
X17 source.t7 plus.t8 drain_left.t7 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X18 source.t26 minus.t8 drain_right.t7 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X19 drain_right.t6 minus.t9 source.t30 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X20 source.t23 minus.t10 drain_right.t5 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X21 a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X22 source.t11 plus.t9 drain_left.t6 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X23 a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X24 drain_left.t5 plus.t10 source.t5 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X25 source.t25 minus.t11 drain_right.t4 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X26 source.t6 plus.t11 drain_left.t4 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X27 drain_right.t3 minus.t12 source.t18 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X28 drain_left.t3 plus.t12 source.t10 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X29 source.t0 plus.t13 drain_left.t2 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X30 a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X31 source.t29 minus.t13 drain_right.t2 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X32 source.t19 minus.t14 drain_right.t1 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X33 drain_left.t1 plus.t14 source.t8 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X34 drain_left.t0 plus.t15 source.t12 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X35 drain_right.t0 minus.t15 source.t20 a_n2390_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
R0 minus.n6 minus.t12 688.953
R1 minus.n30 minus.t14 688.953
R2 minus.n5 minus.t11 667.972
R3 minus.n9 minus.t9 667.972
R4 minus.n3 minus.t8 667.972
R5 minus.n15 minus.t3 667.972
R6 minus.n1 minus.t5 667.972
R7 minus.n21 minus.t4 667.972
R8 minus.n22 minus.t1 667.972
R9 minus.n29 minus.t7 667.972
R10 minus.n33 minus.t10 667.972
R11 minus.n27 minus.t0 667.972
R12 minus.n39 minus.t6 667.972
R13 minus.n25 minus.t2 667.972
R14 minus.n45 minus.t13 667.972
R15 minus.n46 minus.t15 667.972
R16 minus.n23 minus.n22 161.3
R17 minus.n21 minus.n0 161.3
R18 minus.n20 minus.n19 161.3
R19 minus.n18 minus.n1 161.3
R20 minus.n17 minus.n16 161.3
R21 minus.n15 minus.n2 161.3
R22 minus.n14 minus.n13 161.3
R23 minus.n12 minus.n3 161.3
R24 minus.n11 minus.n10 161.3
R25 minus.n9 minus.n4 161.3
R26 minus.n8 minus.n7 161.3
R27 minus.n47 minus.n46 161.3
R28 minus.n45 minus.n24 161.3
R29 minus.n44 minus.n43 161.3
R30 minus.n42 minus.n25 161.3
R31 minus.n41 minus.n40 161.3
R32 minus.n39 minus.n26 161.3
R33 minus.n38 minus.n37 161.3
R34 minus.n36 minus.n27 161.3
R35 minus.n35 minus.n34 161.3
R36 minus.n33 minus.n28 161.3
R37 minus.n32 minus.n31 161.3
R38 minus.n7 minus.n6 70.4033
R39 minus.n31 minus.n30 70.4033
R40 minus.n22 minus.n21 48.2005
R41 minus.n46 minus.n45 48.2005
R42 minus.n9 minus.n8 44.549
R43 minus.n20 minus.n1 44.549
R44 minus.n33 minus.n32 44.549
R45 minus.n44 minus.n25 44.549
R46 minus.n48 minus.n23 40.6028
R47 minus.n10 minus.n3 34.3247
R48 minus.n16 minus.n15 34.3247
R49 minus.n34 minus.n27 34.3247
R50 minus.n40 minus.n39 34.3247
R51 minus.n15 minus.n14 24.1005
R52 minus.n14 minus.n3 24.1005
R53 minus.n38 minus.n27 24.1005
R54 minus.n39 minus.n38 24.1005
R55 minus.n6 minus.n5 20.9576
R56 minus.n30 minus.n29 20.9576
R57 minus.n10 minus.n9 13.8763
R58 minus.n16 minus.n1 13.8763
R59 minus.n34 minus.n33 13.8763
R60 minus.n40 minus.n25 13.8763
R61 minus.n48 minus.n47 6.6558
R62 minus.n8 minus.n5 3.65202
R63 minus.n21 minus.n20 3.65202
R64 minus.n32 minus.n29 3.65202
R65 minus.n45 minus.n44 3.65202
R66 minus.n23 minus.n0 0.189894
R67 minus.n19 minus.n0 0.189894
R68 minus.n19 minus.n18 0.189894
R69 minus.n18 minus.n17 0.189894
R70 minus.n17 minus.n2 0.189894
R71 minus.n13 minus.n2 0.189894
R72 minus.n13 minus.n12 0.189894
R73 minus.n12 minus.n11 0.189894
R74 minus.n11 minus.n4 0.189894
R75 minus.n7 minus.n4 0.189894
R76 minus.n31 minus.n28 0.189894
R77 minus.n35 minus.n28 0.189894
R78 minus.n36 minus.n35 0.189894
R79 minus.n37 minus.n36 0.189894
R80 minus.n37 minus.n26 0.189894
R81 minus.n41 minus.n26 0.189894
R82 minus.n42 minus.n41 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n24 0.189894
R85 minus.n47 minus.n24 0.189894
R86 minus minus.n48 0.188
R87 source.n7 source.t0 45.521
R88 source.n8 source.t18 45.521
R89 source.n15 source.t22 45.521
R90 source.n31 source.t20 45.5208
R91 source.n24 source.t19 45.5208
R92 source.n23 source.t3 45.5208
R93 source.n16 source.t2 45.5208
R94 source.n0 source.t14 45.5208
R95 source.n2 source.n1 44.201
R96 source.n4 source.n3 44.201
R97 source.n6 source.n5 44.201
R98 source.n10 source.n9 44.201
R99 source.n12 source.n11 44.201
R100 source.n14 source.n13 44.201
R101 source.n30 source.n29 44.2008
R102 source.n28 source.n27 44.2008
R103 source.n26 source.n25 44.2008
R104 source.n22 source.n21 44.2008
R105 source.n20 source.n19 44.2008
R106 source.n18 source.n17 44.2008
R107 source.n16 source.n15 24.3622
R108 source.n32 source.n0 18.6984
R109 source.n32 source.n31 5.66429
R110 source.n29 source.t16 1.3205
R111 source.n29 source.t29 1.3205
R112 source.n27 source.t31 1.3205
R113 source.n27 source.t21 1.3205
R114 source.n25 source.t27 1.3205
R115 source.n25 source.t23 1.3205
R116 source.n21 source.t8 1.3205
R117 source.n21 source.t11 1.3205
R118 source.n19 source.t15 1.3205
R119 source.n19 source.t9 1.3205
R120 source.n17 source.t12 1.3205
R121 source.n17 source.t1 1.3205
R122 source.n1 source.t4 1.3205
R123 source.n1 source.t13 1.3205
R124 source.n3 source.t5 1.3205
R125 source.n3 source.t7 1.3205
R126 source.n5 source.t10 1.3205
R127 source.n5 source.t6 1.3205
R128 source.n9 source.t30 1.3205
R129 source.n9 source.t25 1.3205
R130 source.n11 source.t17 1.3205
R131 source.n11 source.t26 1.3205
R132 source.n13 source.t24 1.3205
R133 source.n13 source.t28 1.3205
R134 source.n15 source.n14 0.802224
R135 source.n14 source.n12 0.802224
R136 source.n12 source.n10 0.802224
R137 source.n10 source.n8 0.802224
R138 source.n7 source.n6 0.802224
R139 source.n6 source.n4 0.802224
R140 source.n4 source.n2 0.802224
R141 source.n2 source.n0 0.802224
R142 source.n18 source.n16 0.802224
R143 source.n20 source.n18 0.802224
R144 source.n22 source.n20 0.802224
R145 source.n23 source.n22 0.802224
R146 source.n26 source.n24 0.802224
R147 source.n28 source.n26 0.802224
R148 source.n30 source.n28 0.802224
R149 source.n31 source.n30 0.802224
R150 source.n8 source.n7 0.470328
R151 source.n24 source.n23 0.470328
R152 source source.n32 0.188
R153 drain_right.n9 drain_right.n7 61.6814
R154 drain_right.n5 drain_right.n3 61.6813
R155 drain_right.n2 drain_right.n0 61.6813
R156 drain_right.n9 drain_right.n8 60.8798
R157 drain_right.n11 drain_right.n10 60.8798
R158 drain_right.n13 drain_right.n12 60.8798
R159 drain_right.n5 drain_right.n4 60.8796
R160 drain_right.n2 drain_right.n1 60.8796
R161 drain_right drain_right.n6 34.2978
R162 drain_right drain_right.n13 6.45494
R163 drain_right.n3 drain_right.t2 1.3205
R164 drain_right.n3 drain_right.t0 1.3205
R165 drain_right.n4 drain_right.t9 1.3205
R166 drain_right.n4 drain_right.t13 1.3205
R167 drain_right.n1 drain_right.t5 1.3205
R168 drain_right.n1 drain_right.t15 1.3205
R169 drain_right.n0 drain_right.t1 1.3205
R170 drain_right.n0 drain_right.t8 1.3205
R171 drain_right.n7 drain_right.t4 1.3205
R172 drain_right.n7 drain_right.t3 1.3205
R173 drain_right.n8 drain_right.t7 1.3205
R174 drain_right.n8 drain_right.t6 1.3205
R175 drain_right.n10 drain_right.t10 1.3205
R176 drain_right.n10 drain_right.t12 1.3205
R177 drain_right.n12 drain_right.t14 1.3205
R178 drain_right.n12 drain_right.t11 1.3205
R179 drain_right.n13 drain_right.n11 0.802224
R180 drain_right.n11 drain_right.n9 0.802224
R181 drain_right.n6 drain_right.n5 0.346016
R182 drain_right.n6 drain_right.n2 0.346016
R183 plus.n6 plus.t13 688.953
R184 plus.n30 plus.t0 688.953
R185 plus.n22 plus.t2 667.972
R186 plus.n21 plus.t4 667.972
R187 plus.n1 plus.t5 667.972
R188 plus.n15 plus.t8 667.972
R189 plus.n3 plus.t10 667.972
R190 plus.n9 plus.t11 667.972
R191 plus.n5 plus.t12 667.972
R192 plus.n46 plus.t3 667.972
R193 plus.n45 plus.t15 667.972
R194 plus.n25 plus.t7 667.972
R195 plus.n39 plus.t6 667.972
R196 plus.n27 plus.t1 667.972
R197 plus.n33 plus.t14 667.972
R198 plus.n29 plus.t9 667.972
R199 plus.n8 plus.n7 161.3
R200 plus.n9 plus.n4 161.3
R201 plus.n11 plus.n10 161.3
R202 plus.n12 plus.n3 161.3
R203 plus.n14 plus.n13 161.3
R204 plus.n15 plus.n2 161.3
R205 plus.n17 plus.n16 161.3
R206 plus.n18 plus.n1 161.3
R207 plus.n20 plus.n19 161.3
R208 plus.n21 plus.n0 161.3
R209 plus.n23 plus.n22 161.3
R210 plus.n32 plus.n31 161.3
R211 plus.n33 plus.n28 161.3
R212 plus.n35 plus.n34 161.3
R213 plus.n36 plus.n27 161.3
R214 plus.n38 plus.n37 161.3
R215 plus.n39 plus.n26 161.3
R216 plus.n41 plus.n40 161.3
R217 plus.n42 plus.n25 161.3
R218 plus.n44 plus.n43 161.3
R219 plus.n45 plus.n24 161.3
R220 plus.n47 plus.n46 161.3
R221 plus.n7 plus.n6 70.4033
R222 plus.n31 plus.n30 70.4033
R223 plus.n22 plus.n21 48.2005
R224 plus.n46 plus.n45 48.2005
R225 plus.n20 plus.n1 44.549
R226 plus.n9 plus.n8 44.549
R227 plus.n44 plus.n25 44.549
R228 plus.n33 plus.n32 44.549
R229 plus.n16 plus.n15 34.3247
R230 plus.n10 plus.n3 34.3247
R231 plus.n40 plus.n39 34.3247
R232 plus.n34 plus.n27 34.3247
R233 plus plus.n47 33.3475
R234 plus.n14 plus.n3 24.1005
R235 plus.n15 plus.n14 24.1005
R236 plus.n39 plus.n38 24.1005
R237 plus.n38 plus.n27 24.1005
R238 plus.n6 plus.n5 20.9576
R239 plus.n30 plus.n29 20.9576
R240 plus.n16 plus.n1 13.8763
R241 plus.n10 plus.n9 13.8763
R242 plus.n40 plus.n25 13.8763
R243 plus.n34 plus.n33 13.8763
R244 plus plus.n23 13.4361
R245 plus.n21 plus.n20 3.65202
R246 plus.n8 plus.n5 3.65202
R247 plus.n45 plus.n44 3.65202
R248 plus.n32 plus.n29 3.65202
R249 plus.n7 plus.n4 0.189894
R250 plus.n11 plus.n4 0.189894
R251 plus.n12 plus.n11 0.189894
R252 plus.n13 plus.n12 0.189894
R253 plus.n13 plus.n2 0.189894
R254 plus.n17 plus.n2 0.189894
R255 plus.n18 plus.n17 0.189894
R256 plus.n19 plus.n18 0.189894
R257 plus.n19 plus.n0 0.189894
R258 plus.n23 plus.n0 0.189894
R259 plus.n47 plus.n24 0.189894
R260 plus.n43 plus.n24 0.189894
R261 plus.n43 plus.n42 0.189894
R262 plus.n42 plus.n41 0.189894
R263 plus.n41 plus.n26 0.189894
R264 plus.n37 plus.n26 0.189894
R265 plus.n37 plus.n36 0.189894
R266 plus.n36 plus.n35 0.189894
R267 plus.n35 plus.n28 0.189894
R268 plus.n31 plus.n28 0.189894
R269 drain_left.n9 drain_left.n7 61.6815
R270 drain_left.n5 drain_left.n3 61.6813
R271 drain_left.n2 drain_left.n0 61.6813
R272 drain_left.n11 drain_left.n10 60.8798
R273 drain_left.n9 drain_left.n8 60.8798
R274 drain_left.n13 drain_left.n12 60.8796
R275 drain_left.n5 drain_left.n4 60.8796
R276 drain_left.n2 drain_left.n1 60.8796
R277 drain_left drain_left.n6 34.851
R278 drain_left drain_left.n13 6.45494
R279 drain_left.n3 drain_left.t6 1.3205
R280 drain_left.n3 drain_left.t15 1.3205
R281 drain_left.n4 drain_left.t14 1.3205
R282 drain_left.n4 drain_left.t1 1.3205
R283 drain_left.n1 drain_left.t8 1.3205
R284 drain_left.n1 drain_left.t9 1.3205
R285 drain_left.n0 drain_left.t12 1.3205
R286 drain_left.n0 drain_left.t0 1.3205
R287 drain_left.n12 drain_left.t11 1.3205
R288 drain_left.n12 drain_left.t13 1.3205
R289 drain_left.n10 drain_left.t7 1.3205
R290 drain_left.n10 drain_left.t10 1.3205
R291 drain_left.n8 drain_left.t4 1.3205
R292 drain_left.n8 drain_left.t5 1.3205
R293 drain_left.n7 drain_left.t2 1.3205
R294 drain_left.n7 drain_left.t3 1.3205
R295 drain_left.n11 drain_left.n9 0.802224
R296 drain_left.n13 drain_left.n11 0.802224
R297 drain_left.n6 drain_left.n5 0.346016
R298 drain_left.n6 drain_left.n2 0.346016
C0 drain_left source 25.9375f
C1 drain_left drain_right 1.24373f
C2 plus minus 6.6798f
C3 source drain_right 25.9392f
C4 drain_left minus 0.172752f
C5 drain_left plus 11.7944f
C6 source minus 11.4009f
C7 drain_right minus 11.558499f
C8 source plus 11.414901f
C9 drain_right plus 0.391974f
C10 drain_right a_n2390_n3888# 7.23827f
C11 drain_left a_n2390_n3888# 7.578239f
C12 source a_n2390_n3888# 10.82193f
C13 minus a_n2390_n3888# 9.685987f
C14 plus a_n2390_n3888# 11.65742f
C15 drain_left.t12 a_n2390_n3888# 0.333599f
C16 drain_left.t0 a_n2390_n3888# 0.333599f
C17 drain_left.n0 a_n2390_n3888# 3.02038f
C18 drain_left.t8 a_n2390_n3888# 0.333599f
C19 drain_left.t9 a_n2390_n3888# 0.333599f
C20 drain_left.n1 a_n2390_n3888# 3.01535f
C21 drain_left.n2 a_n2390_n3888# 0.718664f
C22 drain_left.t6 a_n2390_n3888# 0.333599f
C23 drain_left.t15 a_n2390_n3888# 0.333599f
C24 drain_left.n3 a_n2390_n3888# 3.02038f
C25 drain_left.t14 a_n2390_n3888# 0.333599f
C26 drain_left.t1 a_n2390_n3888# 0.333599f
C27 drain_left.n4 a_n2390_n3888# 3.01535f
C28 drain_left.n5 a_n2390_n3888# 0.718664f
C29 drain_left.n6 a_n2390_n3888# 1.75816f
C30 drain_left.t2 a_n2390_n3888# 0.333599f
C31 drain_left.t3 a_n2390_n3888# 0.333599f
C32 drain_left.n7 a_n2390_n3888# 3.02038f
C33 drain_left.t4 a_n2390_n3888# 0.333599f
C34 drain_left.t5 a_n2390_n3888# 0.333599f
C35 drain_left.n8 a_n2390_n3888# 3.01535f
C36 drain_left.n9 a_n2390_n3888# 0.758142f
C37 drain_left.t7 a_n2390_n3888# 0.333599f
C38 drain_left.t10 a_n2390_n3888# 0.333599f
C39 drain_left.n10 a_n2390_n3888# 3.01535f
C40 drain_left.n11 a_n2390_n3888# 0.37592f
C41 drain_left.t11 a_n2390_n3888# 0.333599f
C42 drain_left.t13 a_n2390_n3888# 0.333599f
C43 drain_left.n12 a_n2390_n3888# 3.01534f
C44 drain_left.n13 a_n2390_n3888# 0.621341f
C45 plus.n0 a_n2390_n3888# 0.043107f
C46 plus.t2 a_n2390_n3888# 1.10248f
C47 plus.t4 a_n2390_n3888# 1.10248f
C48 plus.t5 a_n2390_n3888# 1.10248f
C49 plus.n1 a_n2390_n3888# 0.42939f
C50 plus.n2 a_n2390_n3888# 0.043107f
C51 plus.t8 a_n2390_n3888# 1.10248f
C52 plus.t10 a_n2390_n3888# 1.10248f
C53 plus.n3 a_n2390_n3888# 0.42939f
C54 plus.n4 a_n2390_n3888# 0.043107f
C55 plus.t11 a_n2390_n3888# 1.10248f
C56 plus.t12 a_n2390_n3888# 1.10248f
C57 plus.n5 a_n2390_n3888# 0.428194f
C58 plus.t13 a_n2390_n3888# 1.1155f
C59 plus.n6 a_n2390_n3888# 0.414852f
C60 plus.n7 a_n2390_n3888# 0.145188f
C61 plus.n8 a_n2390_n3888# 0.009782f
C62 plus.n9 a_n2390_n3888# 0.42939f
C63 plus.n10 a_n2390_n3888# 0.009782f
C64 plus.n11 a_n2390_n3888# 0.043107f
C65 plus.n12 a_n2390_n3888# 0.043107f
C66 plus.n13 a_n2390_n3888# 0.043107f
C67 plus.n14 a_n2390_n3888# 0.009782f
C68 plus.n15 a_n2390_n3888# 0.42939f
C69 plus.n16 a_n2390_n3888# 0.009782f
C70 plus.n17 a_n2390_n3888# 0.043107f
C71 plus.n18 a_n2390_n3888# 0.043107f
C72 plus.n19 a_n2390_n3888# 0.043107f
C73 plus.n20 a_n2390_n3888# 0.009782f
C74 plus.n21 a_n2390_n3888# 0.428194f
C75 plus.n22 a_n2390_n3888# 0.42753f
C76 plus.n23 a_n2390_n3888# 0.560503f
C77 plus.n24 a_n2390_n3888# 0.043107f
C78 plus.t3 a_n2390_n3888# 1.10248f
C79 plus.t15 a_n2390_n3888# 1.10248f
C80 plus.t7 a_n2390_n3888# 1.10248f
C81 plus.n25 a_n2390_n3888# 0.42939f
C82 plus.n26 a_n2390_n3888# 0.043107f
C83 plus.t6 a_n2390_n3888# 1.10248f
C84 plus.t1 a_n2390_n3888# 1.10248f
C85 plus.n27 a_n2390_n3888# 0.42939f
C86 plus.n28 a_n2390_n3888# 0.043107f
C87 plus.t14 a_n2390_n3888# 1.10248f
C88 plus.t9 a_n2390_n3888# 1.10248f
C89 plus.n29 a_n2390_n3888# 0.428194f
C90 plus.t0 a_n2390_n3888# 1.1155f
C91 plus.n30 a_n2390_n3888# 0.414852f
C92 plus.n31 a_n2390_n3888# 0.145188f
C93 plus.n32 a_n2390_n3888# 0.009782f
C94 plus.n33 a_n2390_n3888# 0.42939f
C95 plus.n34 a_n2390_n3888# 0.009782f
C96 plus.n35 a_n2390_n3888# 0.043107f
C97 plus.n36 a_n2390_n3888# 0.043107f
C98 plus.n37 a_n2390_n3888# 0.043107f
C99 plus.n38 a_n2390_n3888# 0.009782f
C100 plus.n39 a_n2390_n3888# 0.42939f
C101 plus.n40 a_n2390_n3888# 0.009782f
C102 plus.n41 a_n2390_n3888# 0.043107f
C103 plus.n42 a_n2390_n3888# 0.043107f
C104 plus.n43 a_n2390_n3888# 0.043107f
C105 plus.n44 a_n2390_n3888# 0.009782f
C106 plus.n45 a_n2390_n3888# 0.428194f
C107 plus.n46 a_n2390_n3888# 0.42753f
C108 plus.n47 a_n2390_n3888# 1.50964f
C109 drain_right.t1 a_n2390_n3888# 0.332802f
C110 drain_right.t8 a_n2390_n3888# 0.332802f
C111 drain_right.n0 a_n2390_n3888# 3.01316f
C112 drain_right.t5 a_n2390_n3888# 0.332802f
C113 drain_right.t15 a_n2390_n3888# 0.332802f
C114 drain_right.n1 a_n2390_n3888# 3.00814f
C115 drain_right.n2 a_n2390_n3888# 0.716945f
C116 drain_right.t2 a_n2390_n3888# 0.332802f
C117 drain_right.t0 a_n2390_n3888# 0.332802f
C118 drain_right.n3 a_n2390_n3888# 3.01316f
C119 drain_right.t9 a_n2390_n3888# 0.332802f
C120 drain_right.t13 a_n2390_n3888# 0.332802f
C121 drain_right.n4 a_n2390_n3888# 3.00814f
C122 drain_right.n5 a_n2390_n3888# 0.716945f
C123 drain_right.n6 a_n2390_n3888# 1.69602f
C124 drain_right.t4 a_n2390_n3888# 0.332802f
C125 drain_right.t3 a_n2390_n3888# 0.332802f
C126 drain_right.n7 a_n2390_n3888# 3.01315f
C127 drain_right.t7 a_n2390_n3888# 0.332802f
C128 drain_right.t6 a_n2390_n3888# 0.332802f
C129 drain_right.n8 a_n2390_n3888# 3.00814f
C130 drain_right.n9 a_n2390_n3888# 0.756339f
C131 drain_right.t10 a_n2390_n3888# 0.332802f
C132 drain_right.t12 a_n2390_n3888# 0.332802f
C133 drain_right.n10 a_n2390_n3888# 3.00814f
C134 drain_right.n11 a_n2390_n3888# 0.375021f
C135 drain_right.t14 a_n2390_n3888# 0.332802f
C136 drain_right.t11 a_n2390_n3888# 0.332802f
C137 drain_right.n12 a_n2390_n3888# 3.00814f
C138 drain_right.n13 a_n2390_n3888# 0.619844f
C139 source.t14 a_n2390_n3888# 3.12728f
C140 source.n0 a_n2390_n3888# 1.48013f
C141 source.t4 a_n2390_n3888# 0.279057f
C142 source.t13 a_n2390_n3888# 0.279057f
C143 source.n1 a_n2390_n3888# 2.45128f
C144 source.n2 a_n2390_n3888# 0.353529f
C145 source.t5 a_n2390_n3888# 0.279057f
C146 source.t7 a_n2390_n3888# 0.279057f
C147 source.n3 a_n2390_n3888# 2.45128f
C148 source.n4 a_n2390_n3888# 0.353529f
C149 source.t10 a_n2390_n3888# 0.279057f
C150 source.t6 a_n2390_n3888# 0.279057f
C151 source.n5 a_n2390_n3888# 2.45128f
C152 source.n6 a_n2390_n3888# 0.353529f
C153 source.t0 a_n2390_n3888# 3.12729f
C154 source.n7 a_n2390_n3888# 0.413411f
C155 source.t18 a_n2390_n3888# 3.12729f
C156 source.n8 a_n2390_n3888# 0.413411f
C157 source.t30 a_n2390_n3888# 0.279057f
C158 source.t25 a_n2390_n3888# 0.279057f
C159 source.n9 a_n2390_n3888# 2.45128f
C160 source.n10 a_n2390_n3888# 0.353529f
C161 source.t17 a_n2390_n3888# 0.279057f
C162 source.t26 a_n2390_n3888# 0.279057f
C163 source.n11 a_n2390_n3888# 2.45128f
C164 source.n12 a_n2390_n3888# 0.353529f
C165 source.t24 a_n2390_n3888# 0.279057f
C166 source.t28 a_n2390_n3888# 0.279057f
C167 source.n13 a_n2390_n3888# 2.45128f
C168 source.n14 a_n2390_n3888# 0.353529f
C169 source.t22 a_n2390_n3888# 3.12729f
C170 source.n15 a_n2390_n3888# 1.87914f
C171 source.t2 a_n2390_n3888# 3.12728f
C172 source.n16 a_n2390_n3888# 1.87915f
C173 source.t12 a_n2390_n3888# 0.279057f
C174 source.t1 a_n2390_n3888# 0.279057f
C175 source.n17 a_n2390_n3888# 2.45128f
C176 source.n18 a_n2390_n3888# 0.353532f
C177 source.t15 a_n2390_n3888# 0.279057f
C178 source.t9 a_n2390_n3888# 0.279057f
C179 source.n19 a_n2390_n3888# 2.45128f
C180 source.n20 a_n2390_n3888# 0.353532f
C181 source.t8 a_n2390_n3888# 0.279057f
C182 source.t11 a_n2390_n3888# 0.279057f
C183 source.n21 a_n2390_n3888# 2.45128f
C184 source.n22 a_n2390_n3888# 0.353532f
C185 source.t3 a_n2390_n3888# 3.12728f
C186 source.n23 a_n2390_n3888# 0.413415f
C187 source.t19 a_n2390_n3888# 3.12728f
C188 source.n24 a_n2390_n3888# 0.413415f
C189 source.t27 a_n2390_n3888# 0.279057f
C190 source.t23 a_n2390_n3888# 0.279057f
C191 source.n25 a_n2390_n3888# 2.45128f
C192 source.n26 a_n2390_n3888# 0.353532f
C193 source.t31 a_n2390_n3888# 0.279057f
C194 source.t21 a_n2390_n3888# 0.279057f
C195 source.n27 a_n2390_n3888# 2.45128f
C196 source.n28 a_n2390_n3888# 0.353532f
C197 source.t16 a_n2390_n3888# 0.279057f
C198 source.t29 a_n2390_n3888# 0.279057f
C199 source.n29 a_n2390_n3888# 2.45128f
C200 source.n30 a_n2390_n3888# 0.353532f
C201 source.t20 a_n2390_n3888# 3.12728f
C202 source.n31 a_n2390_n3888# 0.561858f
C203 source.n32 a_n2390_n3888# 1.73306f
C204 minus.n0 a_n2390_n3888# 0.042694f
C205 minus.t5 a_n2390_n3888# 1.09192f
C206 minus.n1 a_n2390_n3888# 0.425278f
C207 minus.n2 a_n2390_n3888# 0.042694f
C208 minus.t8 a_n2390_n3888# 1.09192f
C209 minus.n3 a_n2390_n3888# 0.425278f
C210 minus.n4 a_n2390_n3888# 0.042694f
C211 minus.t11 a_n2390_n3888# 1.09192f
C212 minus.n5 a_n2390_n3888# 0.424094f
C213 minus.t12 a_n2390_n3888# 1.10482f
C214 minus.n6 a_n2390_n3888# 0.410879f
C215 minus.n7 a_n2390_n3888# 0.143798f
C216 minus.n8 a_n2390_n3888# 0.009688f
C217 minus.t9 a_n2390_n3888# 1.09192f
C218 minus.n9 a_n2390_n3888# 0.425278f
C219 minus.n10 a_n2390_n3888# 0.009688f
C220 minus.n11 a_n2390_n3888# 0.042694f
C221 minus.n12 a_n2390_n3888# 0.042694f
C222 minus.n13 a_n2390_n3888# 0.042694f
C223 minus.n14 a_n2390_n3888# 0.009688f
C224 minus.t3 a_n2390_n3888# 1.09192f
C225 minus.n15 a_n2390_n3888# 0.425278f
C226 minus.n16 a_n2390_n3888# 0.009688f
C227 minus.n17 a_n2390_n3888# 0.042694f
C228 minus.n18 a_n2390_n3888# 0.042694f
C229 minus.n19 a_n2390_n3888# 0.042694f
C230 minus.n20 a_n2390_n3888# 0.009688f
C231 minus.t4 a_n2390_n3888# 1.09192f
C232 minus.n21 a_n2390_n3888# 0.424094f
C233 minus.t1 a_n2390_n3888# 1.09192f
C234 minus.n22 a_n2390_n3888# 0.423435f
C235 minus.n23 a_n2390_n3888# 1.80288f
C236 minus.n24 a_n2390_n3888# 0.042694f
C237 minus.t2 a_n2390_n3888# 1.09192f
C238 minus.n25 a_n2390_n3888# 0.425278f
C239 minus.n26 a_n2390_n3888# 0.042694f
C240 minus.t0 a_n2390_n3888# 1.09192f
C241 minus.n27 a_n2390_n3888# 0.425278f
C242 minus.n28 a_n2390_n3888# 0.042694f
C243 minus.t7 a_n2390_n3888# 1.09192f
C244 minus.n29 a_n2390_n3888# 0.424094f
C245 minus.t14 a_n2390_n3888# 1.10482f
C246 minus.n30 a_n2390_n3888# 0.410879f
C247 minus.n31 a_n2390_n3888# 0.143798f
C248 minus.n32 a_n2390_n3888# 0.009688f
C249 minus.t10 a_n2390_n3888# 1.09192f
C250 minus.n33 a_n2390_n3888# 0.425278f
C251 minus.n34 a_n2390_n3888# 0.009688f
C252 minus.n35 a_n2390_n3888# 0.042694f
C253 minus.n36 a_n2390_n3888# 0.042694f
C254 minus.n37 a_n2390_n3888# 0.042694f
C255 minus.n38 a_n2390_n3888# 0.009688f
C256 minus.t6 a_n2390_n3888# 1.09192f
C257 minus.n39 a_n2390_n3888# 0.425278f
C258 minus.n40 a_n2390_n3888# 0.009688f
C259 minus.n41 a_n2390_n3888# 0.042694f
C260 minus.n42 a_n2390_n3888# 0.042694f
C261 minus.n43 a_n2390_n3888# 0.042694f
C262 minus.n44 a_n2390_n3888# 0.009688f
C263 minus.t13 a_n2390_n3888# 1.09192f
C264 minus.n45 a_n2390_n3888# 0.424094f
C265 minus.t15 a_n2390_n3888# 1.09192f
C266 minus.n46 a_n2390_n3888# 0.423435f
C267 minus.n47 a_n2390_n3888# 0.294682f
C268 minus.n48 a_n2390_n3888# 2.15769f
.ends

