* NGSPICE file created from diffpair356.ext - technology: sky130A

.subckt diffpair356 minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t5 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X1 drain_left.t13 plus.t0 source.t7 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 drain_left.t12 plus.t1 source.t11 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X3 drain_right.t11 minus.t1 source.t26 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 drain_left.t11 plus.t2 source.t1 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X5 drain_right.t12 minus.t2 source.t25 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X6 drain_right.t8 minus.t3 source.t24 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X7 drain_right.t7 minus.t4 source.t23 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X8 source.t10 plus.t3 drain_left.t10 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X10 drain_left.t9 plus.t4 source.t2 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 source.t13 plus.t5 drain_left.t8 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X12 source.t0 plus.t6 drain_left.t7 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X13 source.t6 plus.t7 drain_left.t6 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X14 source.t22 minus.t5 drain_right.t13 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 source.t21 minus.t6 drain_right.t2 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X16 a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X17 source.t20 minus.t7 drain_right.t0 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X18 source.t19 minus.t8 drain_right.t9 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X19 drain_right.t3 minus.t9 source.t18 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X20 source.t9 plus.t8 drain_left.t5 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X21 drain_left.t4 plus.t9 source.t4 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X22 drain_left.t3 plus.t10 source.t5 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X23 drain_left.t2 plus.t11 source.t8 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X24 drain_right.t6 minus.t10 source.t17 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X25 a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X26 a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X27 source.t16 minus.t11 drain_right.t1 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X28 drain_right.t10 minus.t12 source.t15 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X29 drain_right.t4 minus.t13 source.t14 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X30 drain_left.t1 plus.t12 source.t3 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X31 source.t12 plus.t13 drain_left.t0 a_n1724_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 minus.n15 minus.t4 884.398
R1 minus.n3 minus.t9 884.398
R2 minus.n32 minus.t2 884.398
R3 minus.n20 minus.t13 884.398
R4 minus.n1 minus.t7 827.433
R5 minus.n14 minus.t0 827.433
R6 minus.n12 minus.t10 827.433
R7 minus.n6 minus.t1 827.433
R8 minus.n4 minus.t11 827.433
R9 minus.n18 minus.t5 827.433
R10 minus.n31 minus.t8 827.433
R11 minus.n29 minus.t3 827.433
R12 minus.n23 minus.t12 827.433
R13 minus.n21 minus.t6 827.433
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n15 minus.n14 35.055
R41 minus.n4 minus.n3 35.055
R42 minus.n21 minus.n20 35.055
R43 minus.n32 minus.n31 35.055
R44 minus.n34 minus.n16 33.4153
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n1 drain_right.t4 68.2804
R62 drain_right.n11 drain_right.t7 67.7376
R63 drain_right.n8 drain_right.n6 66.0805
R64 drain_right.n4 drain_right.n2 66.0804
R65 drain_right.n8 drain_right.n7 65.5376
R66 drain_right.n10 drain_right.n9 65.5376
R67 drain_right.n4 drain_right.n3 65.5373
R68 drain_right.n1 drain_right.n0 65.5373
R69 drain_right drain_right.n5 27.664
R70 drain_right drain_right.n11 5.92477
R71 drain_right.n2 drain_right.t9 2.2005
R72 drain_right.n2 drain_right.t12 2.2005
R73 drain_right.n3 drain_right.t13 2.2005
R74 drain_right.n3 drain_right.t8 2.2005
R75 drain_right.n0 drain_right.t2 2.2005
R76 drain_right.n0 drain_right.t10 2.2005
R77 drain_right.n6 drain_right.t1 2.2005
R78 drain_right.n6 drain_right.t3 2.2005
R79 drain_right.n7 drain_right.t0 2.2005
R80 drain_right.n7 drain_right.t11 2.2005
R81 drain_right.n9 drain_right.t5 2.2005
R82 drain_right.n9 drain_right.t6 2.2005
R83 drain_right.n11 drain_right.n10 0.543603
R84 drain_right.n10 drain_right.n8 0.543603
R85 drain_right.n5 drain_right.n1 0.352482
R86 drain_right.n5 drain_right.n4 0.0809298
R87 source.n7 source.t18 51.0588
R88 source.n27 source.t25 51.0586
R89 source.n20 source.t4 51.0586
R90 source.n0 source.t3 51.0586
R91 source.n2 source.n1 48.8588
R92 source.n4 source.n3 48.8588
R93 source.n6 source.n5 48.8588
R94 source.n9 source.n8 48.8588
R95 source.n11 source.n10 48.8588
R96 source.n13 source.n12 48.8588
R97 source.n26 source.n25 48.8586
R98 source.n24 source.n23 48.8586
R99 source.n22 source.n21 48.8586
R100 source.n19 source.n18 48.8586
R101 source.n17 source.n16 48.8586
R102 source.n15 source.n14 48.8586
R103 source.n15 source.n13 20.1012
R104 source.n28 source.n0 14.0236
R105 source.n28 source.n27 5.53498
R106 source.n25 source.t24 2.2005
R107 source.n25 source.t19 2.2005
R108 source.n23 source.t15 2.2005
R109 source.n23 source.t22 2.2005
R110 source.n21 source.t14 2.2005
R111 source.n21 source.t21 2.2005
R112 source.n18 source.t8 2.2005
R113 source.n18 source.t10 2.2005
R114 source.n16 source.t7 2.2005
R115 source.n16 source.t13 2.2005
R116 source.n14 source.t11 2.2005
R117 source.n14 source.t0 2.2005
R118 source.n1 source.t2 2.2005
R119 source.n1 source.t9 2.2005
R120 source.n3 source.t5 2.2005
R121 source.n3 source.t12 2.2005
R122 source.n5 source.t1 2.2005
R123 source.n5 source.t6 2.2005
R124 source.n8 source.t26 2.2005
R125 source.n8 source.t16 2.2005
R126 source.n10 source.t17 2.2005
R127 source.n10 source.t20 2.2005
R128 source.n12 source.t23 2.2005
R129 source.n12 source.t27 2.2005
R130 source.n7 source.n6 0.741879
R131 source.n22 source.n20 0.741879
R132 source.n13 source.n11 0.543603
R133 source.n11 source.n9 0.543603
R134 source.n9 source.n7 0.543603
R135 source.n6 source.n4 0.543603
R136 source.n4 source.n2 0.543603
R137 source.n2 source.n0 0.543603
R138 source.n17 source.n15 0.543603
R139 source.n19 source.n17 0.543603
R140 source.n20 source.n19 0.543603
R141 source.n24 source.n22 0.543603
R142 source.n26 source.n24 0.543603
R143 source.n27 source.n26 0.543603
R144 source source.n28 0.188
R145 plus.n3 plus.t2 884.398
R146 plus.n15 plus.t12 884.398
R147 plus.n20 plus.t9 884.398
R148 plus.n32 plus.t1 884.398
R149 plus.n1 plus.t13 827.433
R150 plus.n4 plus.t7 827.433
R151 plus.n6 plus.t10 827.433
R152 plus.n12 plus.t4 827.433
R153 plus.n14 plus.t8 827.433
R154 plus.n18 plus.t5 827.433
R155 plus.n21 plus.t3 827.433
R156 plus.n23 plus.t11 827.433
R157 plus.n29 plus.t0 827.433
R158 plus.n31 plus.t6 827.433
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 54.0429
R178 plus.n13 plus.n12 54.0429
R179 plus.n30 plus.n29 54.0429
R180 plus.n23 plus.n22 54.0429
R181 plus.n5 plus.n4 37.9763
R182 plus.n14 plus.n13 37.9763
R183 plus.n31 plus.n30 37.9763
R184 plus.n22 plus.n21 37.9763
R185 plus.n4 plus.n3 35.055
R186 plus.n15 plus.n14 35.055
R187 plus.n32 plus.n31 35.055
R188 plus.n21 plus.n20 35.055
R189 plus plus.n33 28.4327
R190 plus.n7 plus.n6 18.9884
R191 plus.n12 plus.n11 18.9884
R192 plus.n29 plus.n28 18.9884
R193 plus.n24 plus.n23 18.9884
R194 plus plus.n16 11.0441
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t11 68.2807
R206 drain_left.n1 drain_left.t12 68.2804
R207 drain_left.n4 drain_left.n2 66.0804
R208 drain_left.n9 drain_left.n8 65.5376
R209 drain_left.n7 drain_left.n6 65.5376
R210 drain_left.n11 drain_left.n10 65.5374
R211 drain_left.n4 drain_left.n3 65.5373
R212 drain_left.n1 drain_left.n0 65.5373
R213 drain_left drain_left.n5 28.2172
R214 drain_left drain_left.n11 6.19632
R215 drain_left.n2 drain_left.t10 2.2005
R216 drain_left.n2 drain_left.t4 2.2005
R217 drain_left.n3 drain_left.t8 2.2005
R218 drain_left.n3 drain_left.t2 2.2005
R219 drain_left.n0 drain_left.t7 2.2005
R220 drain_left.n0 drain_left.t13 2.2005
R221 drain_left.n10 drain_left.t5 2.2005
R222 drain_left.n10 drain_left.t1 2.2005
R223 drain_left.n8 drain_left.t0 2.2005
R224 drain_left.n8 drain_left.t9 2.2005
R225 drain_left.n6 drain_left.t6 2.2005
R226 drain_left.n6 drain_left.t3 2.2005
R227 drain_left.n9 drain_left.n7 0.543603
R228 drain_left.n11 drain_left.n9 0.543603
R229 drain_left.n5 drain_left.n1 0.352482
R230 drain_left.n5 drain_left.n4 0.0809298
C0 drain_right drain_left 0.882512f
C1 drain_right source 21.6653f
C2 minus drain_left 0.171678f
C3 plus drain_left 4.233971f
C4 minus source 3.85929f
C5 plus source 3.87382f
C6 source drain_left 21.673302f
C7 drain_right minus 4.06944f
C8 drain_right plus 0.322849f
C9 plus minus 4.74362f
C10 drain_right a_n1724_n2688# 6.44917f
C11 drain_left a_n1724_n2688# 6.72177f
C12 source a_n1724_n2688# 5.156964f
C13 minus a_n1724_n2688# 6.501832f
C14 plus a_n1724_n2688# 8.27621f
C15 drain_left.t12 a_n1724_n2688# 2.43283f
C16 drain_left.t7 a_n1724_n2688# 0.218233f
C17 drain_left.t13 a_n1724_n2688# 0.218233f
C18 drain_left.n0 a_n1724_n2688# 1.90881f
C19 drain_left.n1 a_n1724_n2688# 0.719326f
C20 drain_left.t10 a_n1724_n2688# 0.218233f
C21 drain_left.t4 a_n1724_n2688# 0.218233f
C22 drain_left.n2 a_n1724_n2688# 1.91182f
C23 drain_left.t8 a_n1724_n2688# 0.218233f
C24 drain_left.t2 a_n1724_n2688# 0.218233f
C25 drain_left.n3 a_n1724_n2688# 1.90881f
C26 drain_left.n4 a_n1724_n2688# 0.678827f
C27 drain_left.n5 a_n1724_n2688# 1.25261f
C28 drain_left.t11 a_n1724_n2688# 2.43283f
C29 drain_left.t6 a_n1724_n2688# 0.218233f
C30 drain_left.t3 a_n1724_n2688# 0.218233f
C31 drain_left.n6 a_n1724_n2688# 1.90882f
C32 drain_left.n7 a_n1724_n2688# 0.736194f
C33 drain_left.t0 a_n1724_n2688# 0.218233f
C34 drain_left.t9 a_n1724_n2688# 0.218233f
C35 drain_left.n8 a_n1724_n2688# 1.90882f
C36 drain_left.n9 a_n1724_n2688# 0.353183f
C37 drain_left.t5 a_n1724_n2688# 0.218233f
C38 drain_left.t1 a_n1724_n2688# 0.218233f
C39 drain_left.n10 a_n1724_n2688# 1.90881f
C40 drain_left.n11 a_n1724_n2688# 0.6086f
C41 plus.n0 a_n1724_n2688# 0.052214f
C42 plus.t8 a_n1724_n2688# 0.399477f
C43 plus.t4 a_n1724_n2688# 0.399477f
C44 plus.t13 a_n1724_n2688# 0.399477f
C45 plus.n1 a_n1724_n2688# 0.184136f
C46 plus.n2 a_n1724_n2688# 0.123017f
C47 plus.t10 a_n1724_n2688# 0.399477f
C48 plus.t7 a_n1724_n2688# 0.399477f
C49 plus.t2 a_n1724_n2688# 0.410616f
C50 plus.n3 a_n1724_n2688# 0.183382f
C51 plus.n4 a_n1724_n2688# 0.166815f
C52 plus.n5 a_n1724_n2688# 0.021506f
C53 plus.n6 a_n1724_n2688# 0.166815f
C54 plus.n7 a_n1724_n2688# 0.021506f
C55 plus.n8 a_n1724_n2688# 0.052214f
C56 plus.n9 a_n1724_n2688# 0.052214f
C57 plus.n10 a_n1724_n2688# 0.052214f
C58 plus.n11 a_n1724_n2688# 0.021506f
C59 plus.n12 a_n1724_n2688# 0.166815f
C60 plus.n13 a_n1724_n2688# 0.021506f
C61 plus.n14 a_n1724_n2688# 0.166815f
C62 plus.t12 a_n1724_n2688# 0.410616f
C63 plus.n15 a_n1724_n2688# 0.183299f
C64 plus.n16 a_n1724_n2688# 0.517515f
C65 plus.n17 a_n1724_n2688# 0.052214f
C66 plus.t1 a_n1724_n2688# 0.410616f
C67 plus.t6 a_n1724_n2688# 0.399477f
C68 plus.t0 a_n1724_n2688# 0.399477f
C69 plus.t5 a_n1724_n2688# 0.399477f
C70 plus.n18 a_n1724_n2688# 0.184136f
C71 plus.n19 a_n1724_n2688# 0.123017f
C72 plus.t11 a_n1724_n2688# 0.399477f
C73 plus.t3 a_n1724_n2688# 0.399477f
C74 plus.t9 a_n1724_n2688# 0.410616f
C75 plus.n20 a_n1724_n2688# 0.183382f
C76 plus.n21 a_n1724_n2688# 0.166815f
C77 plus.n22 a_n1724_n2688# 0.021506f
C78 plus.n23 a_n1724_n2688# 0.166815f
C79 plus.n24 a_n1724_n2688# 0.021506f
C80 plus.n25 a_n1724_n2688# 0.052214f
C81 plus.n26 a_n1724_n2688# 0.052214f
C82 plus.n27 a_n1724_n2688# 0.052214f
C83 plus.n28 a_n1724_n2688# 0.021506f
C84 plus.n29 a_n1724_n2688# 0.166815f
C85 plus.n30 a_n1724_n2688# 0.021506f
C86 plus.n31 a_n1724_n2688# 0.166815f
C87 plus.n32 a_n1724_n2688# 0.183299f
C88 plus.n33 a_n1724_n2688# 1.41841f
C89 source.t3 a_n1724_n2688# 2.45238f
C90 source.n0 a_n1724_n2688# 1.41018f
C91 source.t2 a_n1724_n2688# 0.22998f
C92 source.t9 a_n1724_n2688# 0.22998f
C93 source.n1 a_n1724_n2688# 1.92524f
C94 source.n2 a_n1724_n2688# 0.41456f
C95 source.t5 a_n1724_n2688# 0.22998f
C96 source.t12 a_n1724_n2688# 0.22998f
C97 source.n3 a_n1724_n2688# 1.92524f
C98 source.n4 a_n1724_n2688# 0.41456f
C99 source.t1 a_n1724_n2688# 0.22998f
C100 source.t6 a_n1724_n2688# 0.22998f
C101 source.n5 a_n1724_n2688# 1.92524f
C102 source.n6 a_n1724_n2688# 0.435219f
C103 source.t18 a_n1724_n2688# 2.45239f
C104 source.n7 a_n1724_n2688# 0.53529f
C105 source.t26 a_n1724_n2688# 0.22998f
C106 source.t16 a_n1724_n2688# 0.22998f
C107 source.n8 a_n1724_n2688# 1.92524f
C108 source.n9 a_n1724_n2688# 0.41456f
C109 source.t17 a_n1724_n2688# 0.22998f
C110 source.t20 a_n1724_n2688# 0.22998f
C111 source.n10 a_n1724_n2688# 1.92524f
C112 source.n11 a_n1724_n2688# 0.41456f
C113 source.t23 a_n1724_n2688# 0.22998f
C114 source.t27 a_n1724_n2688# 0.22998f
C115 source.n12 a_n1724_n2688# 1.92524f
C116 source.n13 a_n1724_n2688# 1.83655f
C117 source.t11 a_n1724_n2688# 0.22998f
C118 source.t0 a_n1724_n2688# 0.22998f
C119 source.n14 a_n1724_n2688# 1.92523f
C120 source.n15 a_n1724_n2688# 1.83655f
C121 source.t7 a_n1724_n2688# 0.22998f
C122 source.t13 a_n1724_n2688# 0.22998f
C123 source.n16 a_n1724_n2688# 1.92523f
C124 source.n17 a_n1724_n2688# 0.414565f
C125 source.t8 a_n1724_n2688# 0.22998f
C126 source.t10 a_n1724_n2688# 0.22998f
C127 source.n18 a_n1724_n2688# 1.92523f
C128 source.n19 a_n1724_n2688# 0.414565f
C129 source.t4 a_n1724_n2688# 2.45238f
C130 source.n20 a_n1724_n2688# 0.535296f
C131 source.t14 a_n1724_n2688# 0.22998f
C132 source.t21 a_n1724_n2688# 0.22998f
C133 source.n21 a_n1724_n2688# 1.92523f
C134 source.n22 a_n1724_n2688# 0.435225f
C135 source.t15 a_n1724_n2688# 0.22998f
C136 source.t22 a_n1724_n2688# 0.22998f
C137 source.n23 a_n1724_n2688# 1.92523f
C138 source.n24 a_n1724_n2688# 0.414565f
C139 source.t24 a_n1724_n2688# 0.22998f
C140 source.t19 a_n1724_n2688# 0.22998f
C141 source.n25 a_n1724_n2688# 1.92523f
C142 source.n26 a_n1724_n2688# 0.414565f
C143 source.t25 a_n1724_n2688# 2.45238f
C144 source.n27 a_n1724_n2688# 0.689541f
C145 source.n28 a_n1724_n2688# 1.68334f
C146 drain_right.t4 a_n1724_n2688# 2.43472f
C147 drain_right.t2 a_n1724_n2688# 0.218403f
C148 drain_right.t10 a_n1724_n2688# 0.218403f
C149 drain_right.n0 a_n1724_n2688# 1.9103f
C150 drain_right.n1 a_n1724_n2688# 0.719885f
C151 drain_right.t9 a_n1724_n2688# 0.218403f
C152 drain_right.t12 a_n1724_n2688# 0.218403f
C153 drain_right.n2 a_n1724_n2688# 1.9133f
C154 drain_right.t13 a_n1724_n2688# 0.218403f
C155 drain_right.t8 a_n1724_n2688# 0.218403f
C156 drain_right.n3 a_n1724_n2688# 1.9103f
C157 drain_right.n4 a_n1724_n2688# 0.679354f
C158 drain_right.n5 a_n1724_n2688# 1.19024f
C159 drain_right.t1 a_n1724_n2688# 0.218403f
C160 drain_right.t3 a_n1724_n2688# 0.218403f
C161 drain_right.n6 a_n1724_n2688# 1.9133f
C162 drain_right.t0 a_n1724_n2688# 0.218403f
C163 drain_right.t11 a_n1724_n2688# 0.218403f
C164 drain_right.n7 a_n1724_n2688# 1.9103f
C165 drain_right.n8 a_n1724_n2688# 0.716285f
C166 drain_right.t5 a_n1724_n2688# 0.218403f
C167 drain_right.t6 a_n1724_n2688# 0.218403f
C168 drain_right.n9 a_n1724_n2688# 1.9103f
C169 drain_right.n10 a_n1724_n2688# 0.353458f
C170 drain_right.t7 a_n1724_n2688# 2.43165f
C171 drain_right.n11 a_n1724_n2688# 0.642569f
C172 minus.n0 a_n1724_n2688# 0.051382f
C173 minus.t4 a_n1724_n2688# 0.404075f
C174 minus.t0 a_n1724_n2688# 0.393114f
C175 minus.t10 a_n1724_n2688# 0.393114f
C176 minus.t7 a_n1724_n2688# 0.393114f
C177 minus.n1 a_n1724_n2688# 0.181203f
C178 minus.n2 a_n1724_n2688# 0.121057f
C179 minus.t1 a_n1724_n2688# 0.393114f
C180 minus.t11 a_n1724_n2688# 0.393114f
C181 minus.t9 a_n1724_n2688# 0.404075f
C182 minus.n3 a_n1724_n2688# 0.180461f
C183 minus.n4 a_n1724_n2688# 0.164157f
C184 minus.n5 a_n1724_n2688# 0.021164f
C185 minus.n6 a_n1724_n2688# 0.164157f
C186 minus.n7 a_n1724_n2688# 0.021164f
C187 minus.n8 a_n1724_n2688# 0.051382f
C188 minus.n9 a_n1724_n2688# 0.051382f
C189 minus.n10 a_n1724_n2688# 0.051382f
C190 minus.n11 a_n1724_n2688# 0.021164f
C191 minus.n12 a_n1724_n2688# 0.164157f
C192 minus.n13 a_n1724_n2688# 0.021164f
C193 minus.n14 a_n1724_n2688# 0.164157f
C194 minus.n15 a_n1724_n2688# 0.180379f
C195 minus.n16 a_n1724_n2688# 1.60072f
C196 minus.n17 a_n1724_n2688# 0.051382f
C197 minus.t8 a_n1724_n2688# 0.393114f
C198 minus.t3 a_n1724_n2688# 0.393114f
C199 minus.t5 a_n1724_n2688# 0.393114f
C200 minus.n18 a_n1724_n2688# 0.181203f
C201 minus.n19 a_n1724_n2688# 0.121057f
C202 minus.t12 a_n1724_n2688# 0.393114f
C203 minus.t6 a_n1724_n2688# 0.393114f
C204 minus.t13 a_n1724_n2688# 0.404075f
C205 minus.n20 a_n1724_n2688# 0.180461f
C206 minus.n21 a_n1724_n2688# 0.164157f
C207 minus.n22 a_n1724_n2688# 0.021164f
C208 minus.n23 a_n1724_n2688# 0.164157f
C209 minus.n24 a_n1724_n2688# 0.021164f
C210 minus.n25 a_n1724_n2688# 0.051382f
C211 minus.n26 a_n1724_n2688# 0.051382f
C212 minus.n27 a_n1724_n2688# 0.051382f
C213 minus.n28 a_n1724_n2688# 0.021164f
C214 minus.n29 a_n1724_n2688# 0.164157f
C215 minus.n30 a_n1724_n2688# 0.021164f
C216 minus.n31 a_n1724_n2688# 0.164157f
C217 minus.t2 a_n1724_n2688# 0.404075f
C218 minus.n32 a_n1724_n2688# 0.180379f
C219 minus.n33 a_n1724_n2688# 0.340334f
C220 minus.n34 a_n1724_n2688# 1.95795f
.ends

