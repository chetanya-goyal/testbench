* NGSPICE file created from diffpair195.ext - technology: sky130A

.subckt diffpair195 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t22 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 source.t19 minus.t1 drain_right.t10 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X2 drain_right.t9 minus.t2 source.t14 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X3 drain_left.t11 plus.t0 source.t5 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X4 drain_right.t8 minus.t3 source.t16 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X5 a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X6 source.t23 minus.t4 drain_right.t7 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X7 a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X8 source.t2 plus.t1 drain_left.t10 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X9 drain_left.t9 plus.t2 source.t9 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X10 a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X11 source.t15 minus.t5 drain_right.t6 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X12 source.t8 plus.t3 drain_left.t8 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X13 source.t3 plus.t4 drain_left.t7 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X14 drain_left.t6 plus.t5 source.t4 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X15 drain_right.t5 minus.t6 source.t20 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X16 source.t17 minus.t7 drain_right.t4 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X17 drain_right.t3 minus.t8 source.t13 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X18 drain_left.t5 plus.t6 source.t6 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X19 source.t0 plus.t7 drain_left.t4 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X20 a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X21 drain_left.t3 plus.t8 source.t1 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X22 drain_right.t2 minus.t9 source.t12 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X23 source.t18 minus.t10 drain_right.t1 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X24 source.t21 minus.t11 drain_right.t0 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X25 source.t7 plus.t9 drain_left.t2 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X26 source.t10 plus.t10 drain_left.t1 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X27 drain_left.t0 plus.t11 source.t11 a_n1598_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n13 minus.t1 392.904
R1 minus.n2 minus.t8 392.904
R2 minus.n28 minus.t2 392.904
R3 minus.n17 minus.t5 392.904
R4 minus.n12 minus.t9 345.433
R5 minus.n10 minus.t7 345.433
R6 minus.n3 minus.t3 345.433
R7 minus.n4 minus.t10 345.433
R8 minus.n27 minus.t4 345.433
R9 minus.n25 minus.t6 345.433
R10 minus.n19 minus.t11 345.433
R11 minus.n18 minus.t0 345.433
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n13 minus.n12 44.549
R31 minus.n4 minus.n2 44.549
R32 minus.n18 minus.n17 44.549
R33 minus.n28 minus.n27 44.549
R34 minus.n12 minus.n11 28.4823
R35 minus.n5 minus.n4 28.4823
R36 minus.n20 minus.n18 28.4823
R37 minus.n27 minus.n26 28.4823
R38 minus.n30 minus.n14 28.3679
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 source.n0 source.t6 69.6943
R54 source.n5 source.t2 69.6943
R55 source.n6 source.t13 69.6943
R56 source.n11 source.t19 69.6943
R57 source.n23 source.t14 69.6942
R58 source.n18 source.t15 69.6942
R59 source.n17 source.t9 69.6942
R60 source.n12 source.t10 69.6942
R61 source.n2 source.n1 63.0943
R62 source.n4 source.n3 63.0943
R63 source.n8 source.n7 63.0943
R64 source.n10 source.n9 63.0943
R65 source.n22 source.n21 63.0942
R66 source.n20 source.n19 63.0942
R67 source.n16 source.n15 63.0942
R68 source.n14 source.n13 63.0942
R69 source.n12 source.n11 15.0126
R70 source.n24 source.n0 9.47816
R71 source.n21 source.t20 6.6005
R72 source.n21 source.t23 6.6005
R73 source.n19 source.t22 6.6005
R74 source.n19 source.t21 6.6005
R75 source.n15 source.t1 6.6005
R76 source.n15 source.t7 6.6005
R77 source.n13 source.t5 6.6005
R78 source.n13 source.t3 6.6005
R79 source.n1 source.t11 6.6005
R80 source.n1 source.t8 6.6005
R81 source.n3 source.t4 6.6005
R82 source.n3 source.t0 6.6005
R83 source.n7 source.t16 6.6005
R84 source.n7 source.t18 6.6005
R85 source.n9 source.t12 6.6005
R86 source.n9 source.t17 6.6005
R87 source.n24 source.n23 5.53498
R88 source.n11 source.n10 0.543603
R89 source.n10 source.n8 0.543603
R90 source.n8 source.n6 0.543603
R91 source.n5 source.n4 0.543603
R92 source.n4 source.n2 0.543603
R93 source.n2 source.n0 0.543603
R94 source.n14 source.n12 0.543603
R95 source.n16 source.n14 0.543603
R96 source.n17 source.n16 0.543603
R97 source.n20 source.n18 0.543603
R98 source.n22 source.n20 0.543603
R99 source.n23 source.n22 0.543603
R100 source.n6 source.n5 0.470328
R101 source.n18 source.n17 0.470328
R102 source source.n24 0.188
R103 drain_right.n6 drain_right.n4 80.3162
R104 drain_right.n3 drain_right.n2 80.2608
R105 drain_right.n3 drain_right.n0 80.2608
R106 drain_right.n6 drain_right.n5 79.7731
R107 drain_right.n8 drain_right.n7 79.7731
R108 drain_right.n3 drain_right.n1 79.773
R109 drain_right drain_right.n3 22.7112
R110 drain_right.n1 drain_right.t0 6.6005
R111 drain_right.n1 drain_right.t5 6.6005
R112 drain_right.n2 drain_right.t7 6.6005
R113 drain_right.n2 drain_right.t9 6.6005
R114 drain_right.n0 drain_right.t6 6.6005
R115 drain_right.n0 drain_right.t11 6.6005
R116 drain_right.n4 drain_right.t1 6.6005
R117 drain_right.n4 drain_right.t3 6.6005
R118 drain_right.n5 drain_right.t4 6.6005
R119 drain_right.n5 drain_right.t8 6.6005
R120 drain_right.n7 drain_right.t10 6.6005
R121 drain_right.n7 drain_right.t2 6.6005
R122 drain_right drain_right.n8 6.19632
R123 drain_right.n8 drain_right.n6 0.543603
R124 plus.n2 plus.t1 392.904
R125 plus.n13 plus.t6 392.904
R126 plus.n17 plus.t2 392.904
R127 plus.n28 plus.t10 392.904
R128 plus.n3 plus.t5 345.433
R129 plus.n4 plus.t7 345.433
R130 plus.n10 plus.t11 345.433
R131 plus.n12 plus.t3 345.433
R132 plus.n19 plus.t9 345.433
R133 plus.n18 plus.t8 345.433
R134 plus.n25 plus.t4 345.433
R135 plus.n27 plus.t0 345.433
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 63.5369
R151 plus.n11 plus.n10 63.5369
R152 plus.n26 plus.n25 63.5369
R153 plus.n20 plus.n18 63.5369
R154 plus.n3 plus.n2 44.549
R155 plus.n13 plus.n12 44.549
R156 plus.n28 plus.n27 44.549
R157 plus.n19 plus.n17 44.549
R158 plus.n5 plus.n3 28.4823
R159 plus.n12 plus.n11 28.4823
R160 plus.n27 plus.n26 28.4823
R161 plus.n20 plus.n19 28.4823
R162 plus plus.n29 25.6581
R163 plus.n4 plus.n1 9.49444
R164 plus.n10 plus.n9 9.49444
R165 plus.n25 plus.n24 9.49444
R166 plus.n18 plus.n16 9.49444
R167 plus plus.n14 8.74671
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 80.3162
R177 drain_left.n3 drain_left.n2 80.2608
R178 drain_left.n3 drain_left.n0 80.2608
R179 drain_left.n8 drain_left.n7 79.7731
R180 drain_left.n6 drain_left.n5 79.7731
R181 drain_left.n3 drain_left.n1 79.773
R182 drain_left drain_left.n3 23.2644
R183 drain_left.n1 drain_left.t7 6.6005
R184 drain_left.n1 drain_left.t3 6.6005
R185 drain_left.n2 drain_left.t2 6.6005
R186 drain_left.n2 drain_left.t9 6.6005
R187 drain_left.n0 drain_left.t1 6.6005
R188 drain_left.n0 drain_left.t11 6.6005
R189 drain_left.n7 drain_left.t8 6.6005
R190 drain_left.n7 drain_left.t5 6.6005
R191 drain_left.n5 drain_left.t4 6.6005
R192 drain_left.n5 drain_left.t0 6.6005
R193 drain_left.n4 drain_left.t10 6.6005
R194 drain_left.n4 drain_left.t6 6.6005
R195 drain_left drain_left.n8 6.19632
R196 drain_left.n8 drain_left.n6 0.543603
C0 drain_right drain_left 0.78581f
C1 minus drain_left 0.175831f
C2 plus drain_left 1.64365f
C3 minus drain_right 1.49021f
C4 plus drain_right 0.312678f
C5 source drain_left 7.61714f
C6 minus plus 3.48345f
C7 source drain_right 7.6169f
C8 source minus 1.56747f
C9 source plus 1.58147f
C10 drain_right a_n1598_n1488# 3.75296f
C11 drain_left a_n1598_n1488# 3.97225f
C12 source a_n1598_n1488# 3.568497f
C13 minus a_n1598_n1488# 5.479291f
C14 plus a_n1598_n1488# 6.106687f
C15 drain_left.t1 a_n1598_n1488# 0.061452f
C16 drain_left.t11 a_n1598_n1488# 0.061452f
C17 drain_left.n0 a_n1598_n1488# 0.445039f
C18 drain_left.t7 a_n1598_n1488# 0.061452f
C19 drain_left.t3 a_n1598_n1488# 0.061452f
C20 drain_left.n1 a_n1598_n1488# 0.443183f
C21 drain_left.t2 a_n1598_n1488# 0.061452f
C22 drain_left.t9 a_n1598_n1488# 0.061452f
C23 drain_left.n2 a_n1598_n1488# 0.445039f
C24 drain_left.n3 a_n1598_n1488# 1.58334f
C25 drain_left.t10 a_n1598_n1488# 0.061452f
C26 drain_left.t6 a_n1598_n1488# 0.061452f
C27 drain_left.n4 a_n1598_n1488# 0.445273f
C28 drain_left.t4 a_n1598_n1488# 0.061452f
C29 drain_left.t0 a_n1598_n1488# 0.061452f
C30 drain_left.n5 a_n1598_n1488# 0.443186f
C31 drain_left.n6 a_n1598_n1488# 0.604793f
C32 drain_left.t8 a_n1598_n1488# 0.061452f
C33 drain_left.t5 a_n1598_n1488# 0.061452f
C34 drain_left.n7 a_n1598_n1488# 0.443186f
C35 drain_left.n8 a_n1598_n1488# 0.51398f
C36 plus.n0 a_n1598_n1488# 0.028435f
C37 plus.t3 a_n1598_n1488# 0.074111f
C38 plus.t11 a_n1598_n1488# 0.074111f
C39 plus.n1 a_n1598_n1488# 0.010573f
C40 plus.t1 a_n1598_n1488# 0.079575f
C41 plus.n2 a_n1598_n1488# 0.051514f
C42 plus.t5 a_n1598_n1488# 0.074111f
C43 plus.n3 a_n1598_n1488# 0.043032f
C44 plus.t7 a_n1598_n1488# 0.074111f
C45 plus.n4 a_n1598_n1488# 0.043032f
C46 plus.n5 a_n1598_n1488# 0.011712f
C47 plus.n6 a_n1598_n1488# 0.064717f
C48 plus.n7 a_n1598_n1488# 0.028435f
C49 plus.n8 a_n1598_n1488# 0.028435f
C50 plus.n9 a_n1598_n1488# 0.010573f
C51 plus.n10 a_n1598_n1488# 0.043032f
C52 plus.n11 a_n1598_n1488# 0.011712f
C53 plus.n12 a_n1598_n1488# 0.043032f
C54 plus.t6 a_n1598_n1488# 0.079575f
C55 plus.n13 a_n1598_n1488# 0.051472f
C56 plus.n14 a_n1598_n1488# 0.213245f
C57 plus.n15 a_n1598_n1488# 0.028435f
C58 plus.t10 a_n1598_n1488# 0.079575f
C59 plus.t0 a_n1598_n1488# 0.074111f
C60 plus.t4 a_n1598_n1488# 0.074111f
C61 plus.n16 a_n1598_n1488# 0.010573f
C62 plus.t2 a_n1598_n1488# 0.079575f
C63 plus.n17 a_n1598_n1488# 0.051514f
C64 plus.t8 a_n1598_n1488# 0.074111f
C65 plus.n18 a_n1598_n1488# 0.043032f
C66 plus.t9 a_n1598_n1488# 0.074111f
C67 plus.n19 a_n1598_n1488# 0.043032f
C68 plus.n20 a_n1598_n1488# 0.011712f
C69 plus.n21 a_n1598_n1488# 0.064717f
C70 plus.n22 a_n1598_n1488# 0.028435f
C71 plus.n23 a_n1598_n1488# 0.028435f
C72 plus.n24 a_n1598_n1488# 0.010573f
C73 plus.n25 a_n1598_n1488# 0.043032f
C74 plus.n26 a_n1598_n1488# 0.011712f
C75 plus.n27 a_n1598_n1488# 0.043032f
C76 plus.n28 a_n1598_n1488# 0.051472f
C77 plus.n29 a_n1598_n1488# 0.633058f
C78 drain_right.t6 a_n1598_n1488# 0.062283f
C79 drain_right.t11 a_n1598_n1488# 0.062283f
C80 drain_right.n0 a_n1598_n1488# 0.451057f
C81 drain_right.t0 a_n1598_n1488# 0.062283f
C82 drain_right.t5 a_n1598_n1488# 0.062283f
C83 drain_right.n1 a_n1598_n1488# 0.449176f
C84 drain_right.t7 a_n1598_n1488# 0.062283f
C85 drain_right.t9 a_n1598_n1488# 0.062283f
C86 drain_right.n2 a_n1598_n1488# 0.451057f
C87 drain_right.n3 a_n1598_n1488# 1.55253f
C88 drain_right.t1 a_n1598_n1488# 0.062283f
C89 drain_right.t3 a_n1598_n1488# 0.062283f
C90 drain_right.n4 a_n1598_n1488# 0.451294f
C91 drain_right.t4 a_n1598_n1488# 0.062283f
C92 drain_right.t8 a_n1598_n1488# 0.062283f
C93 drain_right.n5 a_n1598_n1488# 0.449179f
C94 drain_right.n6 a_n1598_n1488# 0.612972f
C95 drain_right.t10 a_n1598_n1488# 0.062283f
C96 drain_right.t2 a_n1598_n1488# 0.062283f
C97 drain_right.n7 a_n1598_n1488# 0.449179f
C98 drain_right.n8 a_n1598_n1488# 0.52093f
C99 source.t6 a_n1598_n1488# 0.482598f
C100 source.n0 a_n1598_n1488# 0.658426f
C101 source.t11 a_n1598_n1488# 0.058118f
C102 source.t8 a_n1598_n1488# 0.058118f
C103 source.n1 a_n1598_n1488# 0.368499f
C104 source.n2 a_n1598_n1488# 0.29936f
C105 source.t4 a_n1598_n1488# 0.058118f
C106 source.t0 a_n1598_n1488# 0.058118f
C107 source.n3 a_n1598_n1488# 0.368499f
C108 source.n4 a_n1598_n1488# 0.29936f
C109 source.t2 a_n1598_n1488# 0.482598f
C110 source.n5 a_n1598_n1488# 0.337975f
C111 source.t13 a_n1598_n1488# 0.482598f
C112 source.n6 a_n1598_n1488# 0.337975f
C113 source.t16 a_n1598_n1488# 0.058118f
C114 source.t18 a_n1598_n1488# 0.058118f
C115 source.n7 a_n1598_n1488# 0.368499f
C116 source.n8 a_n1598_n1488# 0.29936f
C117 source.t12 a_n1598_n1488# 0.058118f
C118 source.t17 a_n1598_n1488# 0.058118f
C119 source.n9 a_n1598_n1488# 0.368499f
C120 source.n10 a_n1598_n1488# 0.29936f
C121 source.t19 a_n1598_n1488# 0.482598f
C122 source.n11 a_n1598_n1488# 0.913962f
C123 source.t10 a_n1598_n1488# 0.482596f
C124 source.n12 a_n1598_n1488# 0.913965f
C125 source.t5 a_n1598_n1488# 0.058118f
C126 source.t3 a_n1598_n1488# 0.058118f
C127 source.n13 a_n1598_n1488# 0.368496f
C128 source.n14 a_n1598_n1488# 0.299363f
C129 source.t1 a_n1598_n1488# 0.058118f
C130 source.t7 a_n1598_n1488# 0.058118f
C131 source.n15 a_n1598_n1488# 0.368496f
C132 source.n16 a_n1598_n1488# 0.299363f
C133 source.t9 a_n1598_n1488# 0.482596f
C134 source.n17 a_n1598_n1488# 0.337978f
C135 source.t15 a_n1598_n1488# 0.482596f
C136 source.n18 a_n1598_n1488# 0.337978f
C137 source.t22 a_n1598_n1488# 0.058118f
C138 source.t21 a_n1598_n1488# 0.058118f
C139 source.n19 a_n1598_n1488# 0.368496f
C140 source.n20 a_n1598_n1488# 0.299363f
C141 source.t20 a_n1598_n1488# 0.058118f
C142 source.t23 a_n1598_n1488# 0.058118f
C143 source.n21 a_n1598_n1488# 0.368496f
C144 source.n22 a_n1598_n1488# 0.299363f
C145 source.t14 a_n1598_n1488# 0.482596f
C146 source.n23 a_n1598_n1488# 0.476365f
C147 source.n24 a_n1598_n1488# 0.710573f
C148 minus.n0 a_n1598_n1488# 0.027976f
C149 minus.t1 a_n1598_n1488# 0.078288f
C150 minus.t9 a_n1598_n1488# 0.072913f
C151 minus.t7 a_n1598_n1488# 0.072913f
C152 minus.n1 a_n1598_n1488# 0.010402f
C153 minus.t8 a_n1598_n1488# 0.078288f
C154 minus.n2 a_n1598_n1488# 0.050682f
C155 minus.t3 a_n1598_n1488# 0.072913f
C156 minus.n3 a_n1598_n1488# 0.042337f
C157 minus.t10 a_n1598_n1488# 0.072913f
C158 minus.n4 a_n1598_n1488# 0.042337f
C159 minus.n5 a_n1598_n1488# 0.011523f
C160 minus.n6 a_n1598_n1488# 0.063671f
C161 minus.n7 a_n1598_n1488# 0.027976f
C162 minus.n8 a_n1598_n1488# 0.027976f
C163 minus.n9 a_n1598_n1488# 0.010402f
C164 minus.n10 a_n1598_n1488# 0.042337f
C165 minus.n11 a_n1598_n1488# 0.011523f
C166 minus.n12 a_n1598_n1488# 0.042337f
C167 minus.n13 a_n1598_n1488# 0.05064f
C168 minus.n14 a_n1598_n1488# 0.660873f
C169 minus.n15 a_n1598_n1488# 0.027976f
C170 minus.t4 a_n1598_n1488# 0.072913f
C171 minus.t6 a_n1598_n1488# 0.072913f
C172 minus.n16 a_n1598_n1488# 0.010402f
C173 minus.t5 a_n1598_n1488# 0.078288f
C174 minus.n17 a_n1598_n1488# 0.050682f
C175 minus.t0 a_n1598_n1488# 0.072913f
C176 minus.n18 a_n1598_n1488# 0.042337f
C177 minus.t11 a_n1598_n1488# 0.072913f
C178 minus.n19 a_n1598_n1488# 0.042337f
C179 minus.n20 a_n1598_n1488# 0.011523f
C180 minus.n21 a_n1598_n1488# 0.063671f
C181 minus.n22 a_n1598_n1488# 0.027976f
C182 minus.n23 a_n1598_n1488# 0.027976f
C183 minus.n24 a_n1598_n1488# 0.010402f
C184 minus.n25 a_n1598_n1488# 0.042337f
C185 minus.n26 a_n1598_n1488# 0.011523f
C186 minus.n27 a_n1598_n1488# 0.042337f
C187 minus.t2 a_n1598_n1488# 0.078288f
C188 minus.n28 a_n1598_n1488# 0.05064f
C189 minus.n29 a_n1598_n1488# 0.183679f
C190 minus.n30 a_n1598_n1488# 0.81639f
.ends

