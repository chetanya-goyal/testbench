* NGSPICE file created from diffpair614.ext - technology: sky130A

.subckt diffpair614 minus drain_right drain_left source plus
X0 a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X1 source.t17 minus.t0 drain_right.t3 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X2 drain_left.t9 plus.t0 source.t1 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X3 source.t19 plus.t1 drain_left.t8 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X4 drain_right.t9 minus.t1 source.t16 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X5 drain_left.t7 plus.t2 source.t3 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X6 a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X7 drain_right.t5 minus.t2 source.t15 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X8 source.t14 minus.t3 drain_right.t4 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X9 drain_left.t6 plus.t3 source.t4 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X10 source.t13 minus.t4 drain_right.t1 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X11 drain_right.t2 minus.t5 source.t12 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X12 drain_right.t0 minus.t6 source.t11 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X13 source.t6 plus.t4 drain_left.t5 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X14 source.t2 plus.t5 drain_left.t4 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X15 source.t10 minus.t7 drain_right.t8 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X16 drain_left.t3 plus.t6 source.t18 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X17 drain_right.t7 minus.t8 source.t9 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X18 source.t5 plus.t7 drain_left.t2 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X19 drain_left.t1 plus.t8 source.t0 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X20 a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X21 drain_right.t6 minus.t9 source.t8 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X22 a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X23 drain_left.t0 plus.t9 source.t7 a_n1832_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
R0 minus.n3 minus.t8 895.006
R1 minus.n13 minus.t9 895.006
R2 minus.n2 minus.t7 868.806
R3 minus.n1 minus.t6 868.806
R4 minus.n6 minus.t4 868.806
R5 minus.n8 minus.t1 868.806
R6 minus.n12 minus.t3 868.806
R7 minus.n11 minus.t5 868.806
R8 minus.n16 minus.t0 868.806
R9 minus.n18 minus.t2 868.806
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n6 minus.n5 161.3
R13 minus.n19 minus.n18 161.3
R14 minus.n17 minus.n10 161.3
R15 minus.n16 minus.n15 161.3
R16 minus.n4 minus.n1 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n8 minus.n7 45.2793
R23 minus.n18 minus.n17 45.2793
R24 minus.n4 minus.n3 45.1669
R25 minus.n14 minus.n13 45.1669
R26 minus.n20 minus.n9 42.2221
R27 minus.n3 minus.n2 14.3992
R28 minus.n13 minus.n12 14.3992
R29 minus.n20 minus.n19 6.60088
R30 minus.n7 minus.n6 2.92171
R31 minus.n17 minus.n16 2.92171
R32 minus.n5 minus.n4 0.285035
R33 minus.n15 minus.n14 0.285035
R34 minus.n9 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n15 minus.n10 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 drain_right.n1 drain_right.t6 61.61
R40 drain_right.n7 drain_right.t9 60.8084
R41 drain_right.n6 drain_right.n4 60.6202
R42 drain_right.n3 drain_right.n2 60.3644
R43 drain_right.n6 drain_right.n5 59.8185
R44 drain_right.n1 drain_right.n0 59.8184
R45 drain_right drain_right.n3 36.2818
R46 drain_right drain_right.n7 6.05408
R47 drain_right.n2 drain_right.t3 0.9905
R48 drain_right.n2 drain_right.t5 0.9905
R49 drain_right.n0 drain_right.t4 0.9905
R50 drain_right.n0 drain_right.t2 0.9905
R51 drain_right.n4 drain_right.t8 0.9905
R52 drain_right.n4 drain_right.t7 0.9905
R53 drain_right.n5 drain_right.t1 0.9905
R54 drain_right.n5 drain_right.t0 0.9905
R55 drain_right.n7 drain_right.n6 0.802224
R56 drain_right.n3 drain_right.n1 0.145585
R57 source.n0 source.t4 44.1297
R58 source.n5 source.t9 44.1296
R59 source.n19 source.t15 44.1295
R60 source.n14 source.t1 44.1295
R61 source.n2 source.n1 43.1397
R62 source.n4 source.n3 43.1397
R63 source.n7 source.n6 43.1397
R64 source.n9 source.n8 43.1397
R65 source.n18 source.n17 43.1396
R66 source.n16 source.n15 43.1396
R67 source.n13 source.n12 43.1396
R68 source.n11 source.n10 43.1396
R69 source.n11 source.n9 28.9518
R70 source.n20 source.n0 22.4863
R71 source.n20 source.n19 5.66429
R72 source.n17 source.t12 0.9905
R73 source.n17 source.t17 0.9905
R74 source.n15 source.t8 0.9905
R75 source.n15 source.t14 0.9905
R76 source.n12 source.t7 0.9905
R77 source.n12 source.t6 0.9905
R78 source.n10 source.t3 0.9905
R79 source.n10 source.t19 0.9905
R80 source.n1 source.t18 0.9905
R81 source.n1 source.t2 0.9905
R82 source.n3 source.t0 0.9905
R83 source.n3 source.t5 0.9905
R84 source.n6 source.t11 0.9905
R85 source.n6 source.t10 0.9905
R86 source.n8 source.t16 0.9905
R87 source.n8 source.t13 0.9905
R88 source.n5 source.n4 0.87119
R89 source.n16 source.n14 0.87119
R90 source.n9 source.n7 0.802224
R91 source.n7 source.n5 0.802224
R92 source.n4 source.n2 0.802224
R93 source.n2 source.n0 0.802224
R94 source.n13 source.n11 0.802224
R95 source.n14 source.n13 0.802224
R96 source.n18 source.n16 0.802224
R97 source.n19 source.n18 0.802224
R98 source source.n20 0.188
R99 plus.n3 plus.t8 895.006
R100 plus.n13 plus.t0 895.006
R101 plus.n8 plus.t3 868.806
R102 plus.n6 plus.t5 868.806
R103 plus.n5 plus.t6 868.806
R104 plus.n4 plus.t7 868.806
R105 plus.n18 plus.t2 868.806
R106 plus.n16 plus.t1 868.806
R107 plus.n15 plus.t9 868.806
R108 plus.n14 plus.t4 868.806
R109 plus.n6 plus.n1 161.3
R110 plus.n7 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n16 plus.n11 161.3
R113 plus.n17 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n5 plus.n2 80.6037
R116 plus.n15 plus.n12 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n8 plus.n7 45.2793
R122 plus.n18 plus.n17 45.2793
R123 plus.n3 plus.n2 45.1669
R124 plus.n13 plus.n12 45.1669
R125 plus plus.n19 33.0729
R126 plus plus.n9 15.2751
R127 plus.n4 plus.n3 14.3992
R128 plus.n14 plus.n13 14.3992
R129 plus.n7 plus.n6 2.92171
R130 plus.n17 plus.n16 2.92171
R131 plus.n2 plus.n1 0.285035
R132 plus.n12 plus.n11 0.285035
R133 plus.n1 plus.n0 0.189894
R134 plus.n9 plus.n0 0.189894
R135 plus.n19 plus.n10 0.189894
R136 plus.n11 plus.n10 0.189894
R137 drain_left.n5 drain_left.t1 61.6101
R138 drain_left.n1 drain_left.t7 61.61
R139 drain_left.n3 drain_left.n2 60.3644
R140 drain_left.n7 drain_left.n6 59.8185
R141 drain_left.n5 drain_left.n4 59.8185
R142 drain_left.n1 drain_left.n0 59.8184
R143 drain_left drain_left.n3 36.835
R144 drain_left drain_left.n7 6.45494
R145 drain_left.n2 drain_left.t5 0.9905
R146 drain_left.n2 drain_left.t9 0.9905
R147 drain_left.n0 drain_left.t8 0.9905
R148 drain_left.n0 drain_left.t0 0.9905
R149 drain_left.n6 drain_left.t4 0.9905
R150 drain_left.n6 drain_left.t6 0.9905
R151 drain_left.n4 drain_left.t2 0.9905
R152 drain_left.n4 drain_left.t3 0.9905
R153 drain_left.n7 drain_left.n5 0.802224
R154 drain_left.n3 drain_left.n1 0.145585
C0 drain_right minus 9.98426f
C1 drain_left source 23.979801f
C2 drain_right source 23.9669f
C3 drain_left plus 10.158f
C4 drain_right plus 0.336175f
C5 drain_left drain_right 0.912619f
C6 minus source 9.43982f
C7 plus minus 6.91127f
C8 plus source 9.45475f
C9 drain_left minus 0.172117f
C10 drain_right a_n1832_n4888# 9.1077f
C11 drain_left a_n1832_n4888# 9.391471f
C12 source a_n1832_n4888# 9.365002f
C13 minus a_n1832_n4888# 7.683152f
C14 plus a_n1832_n4888# 9.88996f
C15 drain_left.t7 a_n1832_n4888# 4.64508f
C16 drain_left.t8 a_n1832_n4888# 0.396873f
C17 drain_left.t0 a_n1832_n4888# 0.396873f
C18 drain_left.n0 a_n1832_n4888# 3.6283f
C19 drain_left.n1 a_n1832_n4888# 0.645014f
C20 drain_left.t5 a_n1832_n4888# 0.396873f
C21 drain_left.t9 a_n1832_n4888# 0.396873f
C22 drain_left.n2 a_n1832_n4888# 3.63131f
C23 drain_left.n3 a_n1832_n4888# 2.06477f
C24 drain_left.t1 a_n1832_n4888# 4.6451f
C25 drain_left.t2 a_n1832_n4888# 0.396873f
C26 drain_left.t3 a_n1832_n4888# 0.396873f
C27 drain_left.n4 a_n1832_n4888# 3.6283f
C28 drain_left.n5 a_n1832_n4888# 0.69412f
C29 drain_left.t4 a_n1832_n4888# 0.396873f
C30 drain_left.t6 a_n1832_n4888# 0.396873f
C31 drain_left.n6 a_n1832_n4888# 3.6283f
C32 drain_left.n7 a_n1832_n4888# 0.560617f
C33 plus.n0 a_n1832_n4888# 0.045378f
C34 plus.t3 a_n1832_n4888# 1.54208f
C35 plus.t5 a_n1832_n4888# 1.54208f
C36 plus.n1 a_n1832_n4888# 0.060552f
C37 plus.t6 a_n1832_n4888# 1.54208f
C38 plus.n2 a_n1832_n4888# 0.219334f
C39 plus.t7 a_n1832_n4888# 1.54208f
C40 plus.t8 a_n1832_n4888# 1.55898f
C41 plus.n3 a_n1832_n4888# 0.562432f
C42 plus.n4 a_n1832_n4888# 0.586764f
C43 plus.n5 a_n1832_n4888# 0.587525f
C44 plus.n6 a_n1832_n4888# 0.577788f
C45 plus.n7 a_n1832_n4888# 0.010297f
C46 plus.n8 a_n1832_n4888# 0.576669f
C47 plus.n9 a_n1832_n4888# 0.69955f
C48 plus.n10 a_n1832_n4888# 0.045378f
C49 plus.t2 a_n1832_n4888# 1.54208f
C50 plus.n11 a_n1832_n4888# 0.060552f
C51 plus.t1 a_n1832_n4888# 1.54208f
C52 plus.n12 a_n1832_n4888# 0.219334f
C53 plus.t9 a_n1832_n4888# 1.54208f
C54 plus.t0 a_n1832_n4888# 1.55898f
C55 plus.n13 a_n1832_n4888# 0.562432f
C56 plus.t4 a_n1832_n4888# 1.54208f
C57 plus.n14 a_n1832_n4888# 0.586764f
C58 plus.n15 a_n1832_n4888# 0.587525f
C59 plus.n16 a_n1832_n4888# 0.577788f
C60 plus.n17 a_n1832_n4888# 0.010297f
C61 plus.n18 a_n1832_n4888# 0.576669f
C62 plus.n19 a_n1832_n4888# 1.60607f
C63 source.t4 a_n1832_n4888# 4.60758f
C64 source.n0 a_n1832_n4888# 1.99326f
C65 source.t18 a_n1832_n4888# 0.40317f
C66 source.t2 a_n1832_n4888# 0.40317f
C67 source.n1 a_n1832_n4888# 3.60451f
C68 source.n2 a_n1832_n4888# 0.393749f
C69 source.t0 a_n1832_n4888# 0.40317f
C70 source.t5 a_n1832_n4888# 0.40317f
C71 source.n3 a_n1832_n4888# 3.60451f
C72 source.n4 a_n1832_n4888# 0.399417f
C73 source.t9 a_n1832_n4888# 4.60759f
C74 source.n5 a_n1832_n4888# 0.495894f
C75 source.t11 a_n1832_n4888# 0.40317f
C76 source.t10 a_n1832_n4888# 0.40317f
C77 source.n6 a_n1832_n4888# 3.60451f
C78 source.n7 a_n1832_n4888# 0.393749f
C79 source.t16 a_n1832_n4888# 0.40317f
C80 source.t13 a_n1832_n4888# 0.40317f
C81 source.n8 a_n1832_n4888# 3.60451f
C82 source.n9 a_n1832_n4888# 2.42376f
C83 source.t3 a_n1832_n4888# 0.40317f
C84 source.t19 a_n1832_n4888# 0.40317f
C85 source.n10 a_n1832_n4888# 3.60452f
C86 source.n11 a_n1832_n4888# 2.42375f
C87 source.t7 a_n1832_n4888# 0.40317f
C88 source.t6 a_n1832_n4888# 0.40317f
C89 source.n12 a_n1832_n4888# 3.60452f
C90 source.n13 a_n1832_n4888# 0.393741f
C91 source.t1 a_n1832_n4888# 4.60756f
C92 source.n14 a_n1832_n4888# 0.49592f
C93 source.t8 a_n1832_n4888# 0.40317f
C94 source.t14 a_n1832_n4888# 0.40317f
C95 source.n15 a_n1832_n4888# 3.60452f
C96 source.n16 a_n1832_n4888# 0.39941f
C97 source.t12 a_n1832_n4888# 0.40317f
C98 source.t17 a_n1832_n4888# 0.40317f
C99 source.n17 a_n1832_n4888# 3.60452f
C100 source.n18 a_n1832_n4888# 0.393741f
C101 source.t15 a_n1832_n4888# 4.60756f
C102 source.n19 a_n1832_n4888# 0.623817f
C103 source.n20 a_n1832_n4888# 2.30977f
C104 drain_right.t6 a_n1832_n4888# 4.63122f
C105 drain_right.t4 a_n1832_n4888# 0.395689f
C106 drain_right.t2 a_n1832_n4888# 0.395689f
C107 drain_right.n0 a_n1832_n4888# 3.61747f
C108 drain_right.n1 a_n1832_n4888# 0.643089f
C109 drain_right.t3 a_n1832_n4888# 0.395689f
C110 drain_right.t5 a_n1832_n4888# 0.395689f
C111 drain_right.n2 a_n1832_n4888# 3.62047f
C112 drain_right.n3 a_n1832_n4888# 2.00647f
C113 drain_right.t8 a_n1832_n4888# 0.395689f
C114 drain_right.t7 a_n1832_n4888# 0.395689f
C115 drain_right.n4 a_n1832_n4888# 3.62211f
C116 drain_right.t1 a_n1832_n4888# 0.395689f
C117 drain_right.t0 a_n1832_n4888# 0.395689f
C118 drain_right.n5 a_n1832_n4888# 3.61747f
C119 drain_right.n6 a_n1832_n4888# 0.686706f
C120 drain_right.t9 a_n1832_n4888# 4.62661f
C121 drain_right.n7 a_n1832_n4888# 0.580881f
C122 minus.n0 a_n1832_n4888# 0.044712f
C123 minus.t6 a_n1832_n4888# 1.51945f
C124 minus.n1 a_n1832_n4888# 0.578902f
C125 minus.t4 a_n1832_n4888# 1.51945f
C126 minus.t8 a_n1832_n4888# 1.5361f
C127 minus.t7 a_n1832_n4888# 1.51945f
C128 minus.n2 a_n1832_n4888# 0.578151f
C129 minus.n3 a_n1832_n4888# 0.554177f
C130 minus.n4 a_n1832_n4888# 0.216115f
C131 minus.n5 a_n1832_n4888# 0.059663f
C132 minus.n6 a_n1832_n4888# 0.569307f
C133 minus.n7 a_n1832_n4888# 0.010146f
C134 minus.t1 a_n1832_n4888# 1.51945f
C135 minus.n8 a_n1832_n4888# 0.568205f
C136 minus.n9 a_n1832_n4888# 1.99856f
C137 minus.n10 a_n1832_n4888# 0.044712f
C138 minus.t5 a_n1832_n4888# 1.51945f
C139 minus.n11 a_n1832_n4888# 0.578902f
C140 minus.t9 a_n1832_n4888# 1.5361f
C141 minus.t3 a_n1832_n4888# 1.51945f
C142 minus.n12 a_n1832_n4888# 0.578151f
C143 minus.n13 a_n1832_n4888# 0.554177f
C144 minus.n14 a_n1832_n4888# 0.216115f
C145 minus.n15 a_n1832_n4888# 0.059663f
C146 minus.t0 a_n1832_n4888# 1.51945f
C147 minus.n16 a_n1832_n4888# 0.569307f
C148 minus.n17 a_n1832_n4888# 0.010146f
C149 minus.t2 a_n1832_n4888# 1.51945f
C150 minus.n18 a_n1832_n4888# 0.568205f
C151 minus.n19 a_n1832_n4888# 0.302894f
C152 minus.n20 a_n1832_n4888# 2.38265f
.ends

