* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t24 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X1 source.t20 plus.t1 drain_left.t12 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X2 drain_left.t11 plus.t2 source.t26 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X3 source.t25 plus.t3 drain_left.t10 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X4 drain_right.t13 minus.t0 source.t12 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 drain_right.t12 minus.t1 source.t13 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X6 source.t10 minus.t2 drain_right.t11 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X7 drain_right.t10 minus.t3 source.t2 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X9 drain_right.t9 minus.t4 source.t3 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X10 source.t5 minus.t5 drain_right.t8 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 source.t27 plus.t4 drain_left.t9 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X12 drain_left.t8 plus.t5 source.t16 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 source.t7 minus.t6 drain_right.t7 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 drain_right.t6 minus.t7 source.t9 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 drain_left.t7 plus.t6 source.t19 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X16 source.t17 plus.t7 drain_left.t6 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X17 source.t0 minus.t8 drain_right.t5 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X18 drain_left.t5 plus.t8 source.t21 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X19 a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X20 drain_left.t4 plus.t9 source.t22 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 drain_right.t4 minus.t9 source.t1 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X22 a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X23 source.t15 plus.t10 drain_left.t3 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X24 drain_left.t2 plus.t11 source.t23 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X25 a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X26 drain_right.t3 minus.t10 source.t4 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X27 source.t14 plus.t12 drain_left.t1 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X28 source.t6 minus.t11 drain_right.t2 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X29 source.t8 minus.t12 drain_right.t1 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X30 drain_right.t0 minus.t13 source.t11 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X31 drain_left.t0 plus.t13 source.t18 a_n2204_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n7 plus.n6 161.3
R1 plus.n8 plus.n3 161.3
R2 plus.n11 plus.n2 161.3
R3 plus.n13 plus.n12 161.3
R4 plus.n14 plus.n1 161.3
R5 plus.n15 plus.n0 161.3
R6 plus.n17 plus.n16 161.3
R7 plus.n25 plus.n24 161.3
R8 plus.n26 plus.n21 161.3
R9 plus.n29 plus.n20 161.3
R10 plus.n31 plus.n30 161.3
R11 plus.n32 plus.n19 161.3
R12 plus.n33 plus.n18 161.3
R13 plus.n35 plus.n34 161.3
R14 plus.n5 plus.t11 129.486
R15 plus.n23 plus.t6 129.486
R16 plus.n16 plus.t2 105.638
R17 plus.n14 plus.t3 105.638
R18 plus.n2 plus.t5 105.638
R19 plus.n9 plus.t7 105.638
R20 plus.n8 plus.t9 105.638
R21 plus.n4 plus.t10 105.638
R22 plus.n34 plus.t0 105.638
R23 plus.n32 plus.t4 105.638
R24 plus.n20 plus.t8 105.638
R25 plus.n27 plus.t12 105.638
R26 plus.n26 plus.t13 105.638
R27 plus.n22 plus.t1 105.638
R28 plus.n10 plus.n9 80.6037
R29 plus.n28 plus.n27 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n14 plus.n13 45.2793
R35 plus.n7 plus.n4 45.2793
R36 plus.n32 plus.n31 45.2793
R37 plus.n25 plus.n22 45.2793
R38 plus.n24 plus.n23 44.9119
R39 plus.n6 plus.n5 44.9119
R40 plus.n16 plus.n15 35.055
R41 plus.n34 plus.n33 35.055
R42 plus plus.n35 27.2585
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n15 plus.n14 13.146
R46 plus.n33 plus.n32 13.146
R47 plus plus.n17 8.05164
R48 plus.n13 plus.n2 2.92171
R49 plus.n8 plus.n7 2.92171
R50 plus.n31 plus.n20 2.92171
R51 plus.n26 plus.n25 2.92171
R52 plus.n10 plus.n3 0.285035
R53 plus.n11 plus.n10 0.285035
R54 plus.n29 plus.n28 0.285035
R55 plus.n28 plus.n21 0.285035
R56 plus.n6 plus.n3 0.189894
R57 plus.n12 plus.n11 0.189894
R58 plus.n12 plus.n1 0.189894
R59 plus.n1 plus.n0 0.189894
R60 plus.n17 plus.n0 0.189894
R61 plus.n35 plus.n18 0.189894
R62 plus.n19 plus.n18 0.189894
R63 plus.n30 plus.n19 0.189894
R64 plus.n30 plus.n29 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n0 source.t26 243.255
R67 source.n7 source.t1 243.255
R68 source.n27 source.t3 243.254
R69 source.n20 source.t19 243.254
R70 source.n2 source.n1 223.454
R71 source.n4 source.n3 223.454
R72 source.n6 source.n5 223.454
R73 source.n9 source.n8 223.454
R74 source.n11 source.n10 223.454
R75 source.n13 source.n12 223.454
R76 source.n26 source.n25 223.453
R77 source.n24 source.n23 223.453
R78 source.n22 source.n21 223.453
R79 source.n19 source.n18 223.453
R80 source.n17 source.n16 223.453
R81 source.n15 source.n14 223.453
R82 source.n25 source.t4 19.8005
R83 source.n25 source.t6 19.8005
R84 source.n23 source.t2 19.8005
R85 source.n23 source.t8 19.8005
R86 source.n21 source.t11 19.8005
R87 source.n21 source.t5 19.8005
R88 source.n18 source.t18 19.8005
R89 source.n18 source.t20 19.8005
R90 source.n16 source.t21 19.8005
R91 source.n16 source.t14 19.8005
R92 source.n14 source.t24 19.8005
R93 source.n14 source.t27 19.8005
R94 source.n1 source.t16 19.8005
R95 source.n1 source.t25 19.8005
R96 source.n3 source.t22 19.8005
R97 source.n3 source.t17 19.8005
R98 source.n5 source.t23 19.8005
R99 source.n5 source.t15 19.8005
R100 source.n8 source.t9 19.8005
R101 source.n8 source.t0 19.8005
R102 source.n10 source.t12 19.8005
R103 source.n10 source.t7 19.8005
R104 source.n12 source.t13 19.8005
R105 source.n12 source.t10 19.8005
R106 source.n15 source.n13 14.5578
R107 source.n28 source.n0 8.09232
R108 source.n28 source.n27 5.66429
R109 source.n7 source.n6 0.87119
R110 source.n22 source.n20 0.87119
R111 source.n13 source.n11 0.802224
R112 source.n11 source.n9 0.802224
R113 source.n9 source.n7 0.802224
R114 source.n6 source.n4 0.802224
R115 source.n4 source.n2 0.802224
R116 source.n2 source.n0 0.802224
R117 source.n17 source.n15 0.802224
R118 source.n19 source.n17 0.802224
R119 source.n20 source.n19 0.802224
R120 source.n24 source.n22 0.802224
R121 source.n26 source.n24 0.802224
R122 source.n27 source.n26 0.802224
R123 source source.n28 0.188
R124 drain_left.n7 drain_left.t2 260.735
R125 drain_left.n1 drain_left.t13 260.733
R126 drain_left.n4 drain_left.n2 240.934
R127 drain_left.n11 drain_left.n10 240.132
R128 drain_left.n9 drain_left.n8 240.132
R129 drain_left.n7 drain_left.n6 240.132
R130 drain_left.n4 drain_left.n3 240.131
R131 drain_left.n1 drain_left.n0 240.131
R132 drain_left drain_left.n5 23.6437
R133 drain_left.n2 drain_left.t12 19.8005
R134 drain_left.n2 drain_left.t7 19.8005
R135 drain_left.n3 drain_left.t1 19.8005
R136 drain_left.n3 drain_left.t0 19.8005
R137 drain_left.n0 drain_left.t9 19.8005
R138 drain_left.n0 drain_left.t5 19.8005
R139 drain_left.n10 drain_left.t10 19.8005
R140 drain_left.n10 drain_left.t11 19.8005
R141 drain_left.n8 drain_left.t6 19.8005
R142 drain_left.n8 drain_left.t8 19.8005
R143 drain_left.n6 drain_left.t3 19.8005
R144 drain_left.n6 drain_left.t4 19.8005
R145 drain_left drain_left.n11 6.45494
R146 drain_left.n9 drain_left.n7 0.802224
R147 drain_left.n11 drain_left.n9 0.802224
R148 drain_left.n5 drain_left.n1 0.546447
R149 drain_left.n5 drain_left.n4 0.145585
R150 minus.n17 minus.n16 161.3
R151 minus.n15 minus.n0 161.3
R152 minus.n14 minus.n13 161.3
R153 minus.n12 minus.n1 161.3
R154 minus.n11 minus.n10 161.3
R155 minus.n8 minus.n7 161.3
R156 minus.n6 minus.n3 161.3
R157 minus.n35 minus.n34 161.3
R158 minus.n33 minus.n18 161.3
R159 minus.n32 minus.n31 161.3
R160 minus.n30 minus.n19 161.3
R161 minus.n29 minus.n28 161.3
R162 minus.n26 minus.n25 161.3
R163 minus.n24 minus.n21 161.3
R164 minus.n5 minus.t9 129.486
R165 minus.n23 minus.t13 129.486
R166 minus.n4 minus.t8 105.638
R167 minus.n8 minus.t7 105.638
R168 minus.n9 minus.t6 105.638
R169 minus.n10 minus.t0 105.638
R170 minus.n14 minus.t2 105.638
R171 minus.n16 minus.t1 105.638
R172 minus.n22 minus.t5 105.638
R173 minus.n26 minus.t3 105.638
R174 minus.n27 minus.t12 105.638
R175 minus.n28 minus.t10 105.638
R176 minus.n32 minus.t11 105.638
R177 minus.n34 minus.t4 105.638
R178 minus.n9 minus.n2 80.6037
R179 minus.n27 minus.n20 80.6037
R180 minus.n9 minus.n8 48.2005
R181 minus.n10 minus.n9 48.2005
R182 minus.n27 minus.n26 48.2005
R183 minus.n28 minus.n27 48.2005
R184 minus.n4 minus.n3 45.2793
R185 minus.n14 minus.n1 45.2793
R186 minus.n22 minus.n21 45.2793
R187 minus.n32 minus.n19 45.2793
R188 minus.n6 minus.n5 44.9119
R189 minus.n24 minus.n23 44.9119
R190 minus.n16 minus.n15 35.055
R191 minus.n34 minus.n33 35.055
R192 minus.n36 minus.n17 29.2107
R193 minus.n5 minus.n4 17.739
R194 minus.n23 minus.n22 17.739
R195 minus.n15 minus.n14 13.146
R196 minus.n33 minus.n32 13.146
R197 minus.n36 minus.n35 6.57436
R198 minus.n8 minus.n3 2.92171
R199 minus.n10 minus.n1 2.92171
R200 minus.n26 minus.n21 2.92171
R201 minus.n28 minus.n19 2.92171
R202 minus.n11 minus.n2 0.285035
R203 minus.n7 minus.n2 0.285035
R204 minus.n25 minus.n20 0.285035
R205 minus.n29 minus.n20 0.285035
R206 minus.n17 minus.n0 0.189894
R207 minus.n13 minus.n0 0.189894
R208 minus.n13 minus.n12 0.189894
R209 minus.n12 minus.n11 0.189894
R210 minus.n7 minus.n6 0.189894
R211 minus.n25 minus.n24 0.189894
R212 minus.n30 minus.n29 0.189894
R213 minus.n31 minus.n30 0.189894
R214 minus.n31 minus.n18 0.189894
R215 minus.n35 minus.n18 0.189894
R216 minus minus.n36 0.188
R217 drain_right.n1 drain_right.t0 260.733
R218 drain_right.n11 drain_right.t12 259.933
R219 drain_right.n8 drain_right.n6 240.935
R220 drain_right.n4 drain_right.n2 240.934
R221 drain_right.n8 drain_right.n7 240.132
R222 drain_right.n10 drain_right.n9 240.132
R223 drain_right.n4 drain_right.n3 240.131
R224 drain_right.n1 drain_right.n0 240.131
R225 drain_right drain_right.n5 23.0904
R226 drain_right.n2 drain_right.t2 19.8005
R227 drain_right.n2 drain_right.t9 19.8005
R228 drain_right.n3 drain_right.t1 19.8005
R229 drain_right.n3 drain_right.t3 19.8005
R230 drain_right.n0 drain_right.t8 19.8005
R231 drain_right.n0 drain_right.t10 19.8005
R232 drain_right.n6 drain_right.t5 19.8005
R233 drain_right.n6 drain_right.t4 19.8005
R234 drain_right.n7 drain_right.t7 19.8005
R235 drain_right.n7 drain_right.t6 19.8005
R236 drain_right.n9 drain_right.t11 19.8005
R237 drain_right.n9 drain_right.t13 19.8005
R238 drain_right drain_right.n11 6.05408
R239 drain_right.n11 drain_right.n10 0.802224
R240 drain_right.n10 drain_right.n8 0.802224
R241 drain_right.n5 drain_right.n1 0.546447
R242 drain_right.n5 drain_right.n4 0.145585
C0 plus minus 3.87071f
C1 source plus 1.71257f
C2 drain_left plus 1.38593f
C3 drain_right minus 1.16983f
C4 source drain_right 4.47439f
C5 drain_left drain_right 1.14465f
C6 source minus 1.69866f
C7 drain_left minus 0.180773f
C8 source drain_left 4.47432f
C9 drain_right plus 0.382038f
C10 drain_right a_n2204_n1088# 3.97432f
C11 drain_left a_n2204_n1088# 4.26719f
C12 source a_n2204_n1088# 2.303602f
C13 minus a_n2204_n1088# 7.805969f
C14 plus a_n2204_n1088# 8.419283f
C15 drain_right.t0 a_n2204_n1088# 0.100588f
C16 drain_right.t8 a_n2204_n1088# 0.016157f
C17 drain_right.t10 a_n2204_n1088# 0.016157f
C18 drain_right.n0 a_n2204_n1088# 0.062782f
C19 drain_right.n1 a_n2204_n1088# 0.442937f
C20 drain_right.t2 a_n2204_n1088# 0.016157f
C21 drain_right.t9 a_n2204_n1088# 0.016157f
C22 drain_right.n2 a_n2204_n1088# 0.063637f
C23 drain_right.t1 a_n2204_n1088# 0.016157f
C24 drain_right.t3 a_n2204_n1088# 0.016157f
C25 drain_right.n3 a_n2204_n1088# 0.062782f
C26 drain_right.n4 a_n2204_n1088# 0.464631f
C27 drain_right.n5 a_n2204_n1088# 0.595096f
C28 drain_right.t5 a_n2204_n1088# 0.016157f
C29 drain_right.t4 a_n2204_n1088# 0.016157f
C30 drain_right.n6 a_n2204_n1088# 0.063637f
C31 drain_right.t7 a_n2204_n1088# 0.016157f
C32 drain_right.t6 a_n2204_n1088# 0.016157f
C33 drain_right.n7 a_n2204_n1088# 0.062782f
C34 drain_right.n8 a_n2204_n1088# 0.504625f
C35 drain_right.t11 a_n2204_n1088# 0.016157f
C36 drain_right.t13 a_n2204_n1088# 0.016157f
C37 drain_right.n9 a_n2204_n1088# 0.062782f
C38 drain_right.n10 a_n2204_n1088# 0.248622f
C39 drain_right.t12 a_n2204_n1088# 0.09994f
C40 drain_right.n11 a_n2204_n1088# 0.394556f
C41 minus.n0 a_n2204_n1088# 0.026907f
C42 minus.n1 a_n2204_n1088# 0.006106f
C43 minus.t2 a_n2204_n1088# 0.054745f
C44 minus.n2 a_n2204_n1088# 0.03582f
C45 minus.n3 a_n2204_n1088# 0.006106f
C46 minus.t7 a_n2204_n1088# 0.054745f
C47 minus.t9 a_n2204_n1088# 0.06492f
C48 minus.t8 a_n2204_n1088# 0.054745f
C49 minus.n4 a_n2204_n1088# 0.060217f
C50 minus.n5 a_n2204_n1088# 0.047363f
C51 minus.n6 a_n2204_n1088# 0.11008f
C52 minus.n7 a_n2204_n1088# 0.035904f
C53 minus.n8 a_n2204_n1088# 0.056055f
C54 minus.t6 a_n2204_n1088# 0.054745f
C55 minus.n9 a_n2204_n1088# 0.061829f
C56 minus.t0 a_n2204_n1088# 0.054745f
C57 minus.n10 a_n2204_n1088# 0.056055f
C58 minus.n11 a_n2204_n1088# 0.035904f
C59 minus.n12 a_n2204_n1088# 0.026907f
C60 minus.n13 a_n2204_n1088# 0.026907f
C61 minus.n14 a_n2204_n1088# 0.056884f
C62 minus.n15 a_n2204_n1088# 0.006106f
C63 minus.t1 a_n2204_n1088# 0.054745f
C64 minus.n16 a_n2204_n1088# 0.05423f
C65 minus.n17 a_n2204_n1088# 0.670518f
C66 minus.n18 a_n2204_n1088# 0.026907f
C67 minus.n19 a_n2204_n1088# 0.006106f
C68 minus.n20 a_n2204_n1088# 0.03582f
C69 minus.n21 a_n2204_n1088# 0.006106f
C70 minus.t13 a_n2204_n1088# 0.06492f
C71 minus.t5 a_n2204_n1088# 0.054745f
C72 minus.n22 a_n2204_n1088# 0.060217f
C73 minus.n23 a_n2204_n1088# 0.047363f
C74 minus.n24 a_n2204_n1088# 0.11008f
C75 minus.n25 a_n2204_n1088# 0.035904f
C76 minus.t3 a_n2204_n1088# 0.054745f
C77 minus.n26 a_n2204_n1088# 0.056055f
C78 minus.t12 a_n2204_n1088# 0.054745f
C79 minus.n27 a_n2204_n1088# 0.061829f
C80 minus.t10 a_n2204_n1088# 0.054745f
C81 minus.n28 a_n2204_n1088# 0.056055f
C82 minus.n29 a_n2204_n1088# 0.035904f
C83 minus.n30 a_n2204_n1088# 0.026907f
C84 minus.n31 a_n2204_n1088# 0.026907f
C85 minus.t11 a_n2204_n1088# 0.054745f
C86 minus.n32 a_n2204_n1088# 0.056884f
C87 minus.n33 a_n2204_n1088# 0.006106f
C88 minus.t4 a_n2204_n1088# 0.054745f
C89 minus.n34 a_n2204_n1088# 0.05423f
C90 minus.n35 a_n2204_n1088# 0.180609f
C91 minus.n36 a_n2204_n1088# 0.825667f
C92 drain_left.t13 a_n2204_n1088# 0.098831f
C93 drain_left.t9 a_n2204_n1088# 0.015875f
C94 drain_left.t5 a_n2204_n1088# 0.015875f
C95 drain_left.n0 a_n2204_n1088# 0.061686f
C96 drain_left.n1 a_n2204_n1088# 0.435202f
C97 drain_left.t12 a_n2204_n1088# 0.015875f
C98 drain_left.t7 a_n2204_n1088# 0.015875f
C99 drain_left.n2 a_n2204_n1088# 0.062526f
C100 drain_left.t1 a_n2204_n1088# 0.015875f
C101 drain_left.t0 a_n2204_n1088# 0.015875f
C102 drain_left.n3 a_n2204_n1088# 0.061686f
C103 drain_left.n4 a_n2204_n1088# 0.456517f
C104 drain_left.n5 a_n2204_n1088# 0.623439f
C105 drain_left.t2 a_n2204_n1088# 0.098832f
C106 drain_left.t3 a_n2204_n1088# 0.015875f
C107 drain_left.t4 a_n2204_n1088# 0.015875f
C108 drain_left.n6 a_n2204_n1088# 0.061686f
C109 drain_left.n7 a_n2204_n1088# 0.450905f
C110 drain_left.t6 a_n2204_n1088# 0.015875f
C111 drain_left.t8 a_n2204_n1088# 0.015875f
C112 drain_left.n8 a_n2204_n1088# 0.061686f
C113 drain_left.n9 a_n2204_n1088# 0.24428f
C114 drain_left.t10 a_n2204_n1088# 0.015875f
C115 drain_left.t11 a_n2204_n1088# 0.015875f
C116 drain_left.n10 a_n2204_n1088# 0.061686f
C117 drain_left.n11 a_n2204_n1088# 0.419457f
C118 source.t26 a_n2204_n1088# 0.121528f
C119 source.n0 a_n2204_n1088# 0.562978f
C120 source.t16 a_n2204_n1088# 0.021835f
C121 source.t25 a_n2204_n1088# 0.021835f
C122 source.n1 a_n2204_n1088# 0.070813f
C123 source.n2 a_n2204_n1088# 0.312457f
C124 source.t22 a_n2204_n1088# 0.021835f
C125 source.t17 a_n2204_n1088# 0.021835f
C126 source.n3 a_n2204_n1088# 0.070813f
C127 source.n4 a_n2204_n1088# 0.312457f
C128 source.t23 a_n2204_n1088# 0.021835f
C129 source.t15 a_n2204_n1088# 0.021835f
C130 source.n5 a_n2204_n1088# 0.070813f
C131 source.n6 a_n2204_n1088# 0.318598f
C132 source.t1 a_n2204_n1088# 0.121528f
C133 source.n7 a_n2204_n1088# 0.327431f
C134 source.t9 a_n2204_n1088# 0.021835f
C135 source.t0 a_n2204_n1088# 0.021835f
C136 source.n8 a_n2204_n1088# 0.070813f
C137 source.n9 a_n2204_n1088# 0.312457f
C138 source.t12 a_n2204_n1088# 0.021835f
C139 source.t7 a_n2204_n1088# 0.021835f
C140 source.n10 a_n2204_n1088# 0.070813f
C141 source.n11 a_n2204_n1088# 0.312457f
C142 source.t13 a_n2204_n1088# 0.021835f
C143 source.t10 a_n2204_n1088# 0.021835f
C144 source.n12 a_n2204_n1088# 0.070813f
C145 source.n13 a_n2204_n1088# 0.851826f
C146 source.t24 a_n2204_n1088# 0.021835f
C147 source.t27 a_n2204_n1088# 0.021835f
C148 source.n14 a_n2204_n1088# 0.070813f
C149 source.n15 a_n2204_n1088# 0.851826f
C150 source.t21 a_n2204_n1088# 0.021835f
C151 source.t14 a_n2204_n1088# 0.021835f
C152 source.n16 a_n2204_n1088# 0.070813f
C153 source.n17 a_n2204_n1088# 0.312458f
C154 source.t18 a_n2204_n1088# 0.021835f
C155 source.t20 a_n2204_n1088# 0.021835f
C156 source.n18 a_n2204_n1088# 0.070813f
C157 source.n19 a_n2204_n1088# 0.312458f
C158 source.t19 a_n2204_n1088# 0.121528f
C159 source.n20 a_n2204_n1088# 0.327432f
C160 source.t11 a_n2204_n1088# 0.021835f
C161 source.t5 a_n2204_n1088# 0.021835f
C162 source.n21 a_n2204_n1088# 0.070813f
C163 source.n22 a_n2204_n1088# 0.318598f
C164 source.t2 a_n2204_n1088# 0.021835f
C165 source.t8 a_n2204_n1088# 0.021835f
C166 source.n23 a_n2204_n1088# 0.070813f
C167 source.n24 a_n2204_n1088# 0.312458f
C168 source.t4 a_n2204_n1088# 0.021835f
C169 source.t6 a_n2204_n1088# 0.021835f
C170 source.n25 a_n2204_n1088# 0.070813f
C171 source.n26 a_n2204_n1088# 0.312458f
C172 source.t3 a_n2204_n1088# 0.121528f
C173 source.n27 a_n2204_n1088# 0.465964f
C174 source.n28 a_n2204_n1088# 0.569272f
C175 plus.n0 a_n2204_n1088# 0.027288f
C176 plus.t2 a_n2204_n1088# 0.05552f
C177 plus.t3 a_n2204_n1088# 0.05552f
C178 plus.n1 a_n2204_n1088# 0.027288f
C179 plus.t5 a_n2204_n1088# 0.05552f
C180 plus.n2 a_n2204_n1088# 0.056848f
C181 plus.n3 a_n2204_n1088# 0.036412f
C182 plus.t7 a_n2204_n1088# 0.05552f
C183 plus.t9 a_n2204_n1088# 0.05552f
C184 plus.t10 a_n2204_n1088# 0.05552f
C185 plus.n4 a_n2204_n1088# 0.061069f
C186 plus.t11 a_n2204_n1088# 0.065838f
C187 plus.n5 a_n2204_n1088# 0.048033f
C188 plus.n6 a_n2204_n1088# 0.111637f
C189 plus.n7 a_n2204_n1088# 0.006192f
C190 plus.n8 a_n2204_n1088# 0.056848f
C191 plus.n9 a_n2204_n1088# 0.062704f
C192 plus.n10 a_n2204_n1088# 0.036327f
C193 plus.n11 a_n2204_n1088# 0.036412f
C194 plus.n12 a_n2204_n1088# 0.027288f
C195 plus.n13 a_n2204_n1088# 0.006192f
C196 plus.n14 a_n2204_n1088# 0.057689f
C197 plus.n15 a_n2204_n1088# 0.006192f
C198 plus.n16 a_n2204_n1088# 0.054997f
C199 plus.n17 a_n2204_n1088# 0.192107f
C200 plus.n18 a_n2204_n1088# 0.027288f
C201 plus.t0 a_n2204_n1088# 0.05552f
C202 plus.n19 a_n2204_n1088# 0.027288f
C203 plus.t4 a_n2204_n1088# 0.05552f
C204 plus.t8 a_n2204_n1088# 0.05552f
C205 plus.n20 a_n2204_n1088# 0.056848f
C206 plus.n21 a_n2204_n1088# 0.036412f
C207 plus.t12 a_n2204_n1088# 0.05552f
C208 plus.t13 a_n2204_n1088# 0.05552f
C209 plus.t1 a_n2204_n1088# 0.05552f
C210 plus.n22 a_n2204_n1088# 0.061069f
C211 plus.t6 a_n2204_n1088# 0.065838f
C212 plus.n23 a_n2204_n1088# 0.048033f
C213 plus.n24 a_n2204_n1088# 0.111637f
C214 plus.n25 a_n2204_n1088# 0.006192f
C215 plus.n26 a_n2204_n1088# 0.056848f
C216 plus.n27 a_n2204_n1088# 0.062704f
C217 plus.n28 a_n2204_n1088# 0.036327f
C218 plus.n29 a_n2204_n1088# 0.036412f
C219 plus.n30 a_n2204_n1088# 0.027288f
C220 plus.n31 a_n2204_n1088# 0.006192f
C221 plus.n32 a_n2204_n1088# 0.057689f
C222 plus.n33 a_n2204_n1088# 0.006192f
C223 plus.n34 a_n2204_n1088# 0.054997f
C224 plus.n35 a_n2204_n1088# 0.657376f
.ends

