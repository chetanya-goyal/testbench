* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t29 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X1 drain_right.t19 minus.t0 source.t9 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X2 drain_left.t18 plus.t1 source.t26 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X3 source.t28 plus.t2 drain_left.t17 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X4 drain_left.t16 plus.t3 source.t27 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t13 minus.t1 drain_right.t18 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X6 source.t39 plus.t4 drain_left.t15 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 drain_right.t17 minus.t2 source.t7 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X8 source.t8 minus.t3 drain_right.t16 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_left.t14 plus.t5 source.t30 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X10 source.t19 minus.t4 drain_right.t15 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X11 source.t25 plus.t6 drain_left.t13 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X12 source.t10 minus.t5 drain_right.t14 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X13 drain_right.t13 minus.t6 source.t3 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 drain_right.t12 minus.t7 source.t5 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 drain_right.t11 minus.t8 source.t11 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 drain_right.t10 minus.t9 source.t14 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 source.t0 minus.t10 drain_right.t9 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X18 source.t22 plus.t7 drain_left.t12 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X20 source.t16 minus.t11 drain_right.t8 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X21 a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X22 a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X23 drain_left.t11 plus.t8 source.t32 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X24 a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X25 drain_left.t10 plus.t9 source.t33 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X26 source.t21 plus.t10 drain_left.t9 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X27 source.t34 plus.t11 drain_left.t8 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X28 source.t2 minus.t12 drain_right.t7 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X29 drain_right.t6 minus.t13 source.t1 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X30 drain_left.t7 plus.t12 source.t35 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X31 source.t18 minus.t14 drain_right.t5 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X32 source.t36 plus.t13 drain_left.t6 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X33 drain_right.t4 minus.t15 source.t4 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X34 drain_right.t3 minus.t16 source.t17 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X35 source.t6 minus.t17 drain_right.t2 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X36 source.t24 plus.t14 drain_left.t5 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X37 drain_left.t4 plus.t15 source.t38 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X38 source.t37 plus.t16 drain_left.t3 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X39 source.t12 minus.t18 drain_right.t1 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X40 source.t31 plus.t17 drain_left.t2 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X41 drain_right.t0 minus.t19 source.t15 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X42 drain_left.t1 plus.t18 source.t23 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X43 drain_left.t0 plus.t19 source.t20 a_n2762_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
R0 plus.n8 plus.t16 172.626
R1 plus.n36 plus.t18 172.626
R2 plus.n9 plus.n6 161.3
R3 plus.n11 plus.n10 161.3
R4 plus.n12 plus.n5 161.3
R5 plus.n14 plus.n13 161.3
R6 plus.n15 plus.n4 161.3
R7 plus.n17 plus.n16 161.3
R8 plus.n18 plus.n3 161.3
R9 plus.n20 plus.n19 161.3
R10 plus.n21 plus.n2 161.3
R11 plus.n23 plus.n22 161.3
R12 plus.n24 plus.n1 161.3
R13 plus.n27 plus.n26 161.3
R14 plus.n37 plus.n34 161.3
R15 plus.n39 plus.n38 161.3
R16 plus.n40 plus.n33 161.3
R17 plus.n42 plus.n41 161.3
R18 plus.n43 plus.n32 161.3
R19 plus.n45 plus.n44 161.3
R20 plus.n46 plus.n31 161.3
R21 plus.n48 plus.n47 161.3
R22 plus.n49 plus.n30 161.3
R23 plus.n51 plus.n50 161.3
R24 plus.n52 plus.n29 161.3
R25 plus.n55 plus.n54 161.3
R26 plus.n26 plus.t0 145.805
R27 plus.n25 plus.t2 145.805
R28 plus.n24 plus.t3 145.805
R29 plus.n2 plus.t4 145.805
R30 plus.n18 plus.t5 145.805
R31 plus.n4 plus.t10 145.805
R32 plus.n12 plus.t12 145.805
R33 plus.n6 plus.t13 145.805
R34 plus.n7 plus.t15 145.805
R35 plus.n54 plus.t14 145.805
R36 plus.n53 plus.t1 145.805
R37 plus.n52 plus.t7 145.805
R38 plus.n30 plus.t9 145.805
R39 plus.n46 plus.t17 145.805
R40 plus.n32 plus.t19 145.805
R41 plus.n40 plus.t6 145.805
R42 plus.n34 plus.t8 145.805
R43 plus.n35 plus.t11 145.805
R44 plus.n25 plus.n0 80.6037
R45 plus.n53 plus.n28 80.6037
R46 plus.n26 plus.n25 48.2005
R47 plus.n25 plus.n24 48.2005
R48 plus.n7 plus.n6 48.2005
R49 plus.n54 plus.n53 48.2005
R50 plus.n53 plus.n52 48.2005
R51 plus.n35 plus.n34 48.2005
R52 plus.n9 plus.n8 45.1367
R53 plus.n37 plus.n36 45.1367
R54 plus.n23 plus.n2 44.549
R55 plus.n12 plus.n11 44.549
R56 plus.n51 plus.n30 44.549
R57 plus.n40 plus.n39 44.549
R58 plus.n19 plus.n18 34.3247
R59 plus.n13 plus.n4 34.3247
R60 plus.n47 plus.n46 34.3247
R61 plus.n41 plus.n32 34.3247
R62 plus plus.n55 29.8058
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n19 plus.n2 13.8763
R68 plus.n13 plus.n12 13.8763
R69 plus.n47 plus.n30 13.8763
R70 plus.n41 plus.n40 13.8763
R71 plus.n8 plus.n7 13.3799
R72 plus.n36 plus.n35 13.3799
R73 plus plus.n27 8.48535
R74 plus.n24 plus.n23 3.65202
R75 plus.n11 plus.n6 3.65202
R76 plus.n52 plus.n51 3.65202
R77 plus.n39 plus.n34 3.65202
R78 plus.n1 plus.n0 0.285035
R79 plus.n27 plus.n0 0.285035
R80 plus.n55 plus.n28 0.285035
R81 plus.n29 plus.n28 0.285035
R82 plus.n10 plus.n9 0.189894
R83 plus.n10 plus.n5 0.189894
R84 plus.n14 plus.n5 0.189894
R85 plus.n15 plus.n14 0.189894
R86 plus.n16 plus.n15 0.189894
R87 plus.n16 plus.n3 0.189894
R88 plus.n20 plus.n3 0.189894
R89 plus.n21 plus.n20 0.189894
R90 plus.n22 plus.n21 0.189894
R91 plus.n22 plus.n1 0.189894
R92 plus.n50 plus.n29 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n48 0.189894
R95 plus.n48 plus.n31 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n38 plus.n33 0.189894
R101 plus.n38 plus.n37 0.189894
R102 source.n90 source.n88 289.615
R103 source.n74 source.n72 289.615
R104 source.n66 source.n64 289.615
R105 source.n50 source.n48 289.615
R106 source.n2 source.n0 289.615
R107 source.n18 source.n16 289.615
R108 source.n26 source.n24 289.615
R109 source.n42 source.n40 289.615
R110 source.n91 source.n90 185
R111 source.n75 source.n74 185
R112 source.n67 source.n66 185
R113 source.n51 source.n50 185
R114 source.n3 source.n2 185
R115 source.n19 source.n18 185
R116 source.n27 source.n26 185
R117 source.n43 source.n42 185
R118 source.t9 source.n89 167.117
R119 source.t0 source.n73 167.117
R120 source.t23 source.n65 167.117
R121 source.t24 source.n49 167.117
R122 source.t29 source.n1 167.117
R123 source.t37 source.n17 167.117
R124 source.t4 source.n25 167.117
R125 source.t13 source.n41 167.117
R126 source.n9 source.n8 84.1169
R127 source.n11 source.n10 84.1169
R128 source.n13 source.n12 84.1169
R129 source.n15 source.n14 84.1169
R130 source.n33 source.n32 84.1169
R131 source.n35 source.n34 84.1169
R132 source.n37 source.n36 84.1169
R133 source.n39 source.n38 84.1169
R134 source.n87 source.n86 84.1168
R135 source.n85 source.n84 84.1168
R136 source.n83 source.n82 84.1168
R137 source.n81 source.n80 84.1168
R138 source.n63 source.n62 84.1168
R139 source.n61 source.n60 84.1168
R140 source.n59 source.n58 84.1168
R141 source.n57 source.n56 84.1168
R142 source.n90 source.t9 52.3082
R143 source.n74 source.t0 52.3082
R144 source.n66 source.t23 52.3082
R145 source.n50 source.t24 52.3082
R146 source.n2 source.t29 52.3082
R147 source.n18 source.t37 52.3082
R148 source.n26 source.t4 52.3082
R149 source.n42 source.t13 52.3082
R150 source.n95 source.n94 31.4096
R151 source.n79 source.n78 31.4096
R152 source.n71 source.n70 31.4096
R153 source.n55 source.n54 31.4096
R154 source.n7 source.n6 31.4096
R155 source.n23 source.n22 31.4096
R156 source.n31 source.n30 31.4096
R157 source.n47 source.n46 31.4096
R158 source.n55 source.n47 14.5137
R159 source.n86 source.t17 9.9005
R160 source.n86 source.t10 9.9005
R161 source.n84 source.t3 9.9005
R162 source.n84 source.t12 9.9005
R163 source.n82 source.t14 9.9005
R164 source.n82 source.t8 9.9005
R165 source.n80 source.t15 9.9005
R166 source.n80 source.t6 9.9005
R167 source.n62 source.t32 9.9005
R168 source.n62 source.t34 9.9005
R169 source.n60 source.t20 9.9005
R170 source.n60 source.t25 9.9005
R171 source.n58 source.t33 9.9005
R172 source.n58 source.t31 9.9005
R173 source.n56 source.t26 9.9005
R174 source.n56 source.t22 9.9005
R175 source.n8 source.t27 9.9005
R176 source.n8 source.t28 9.9005
R177 source.n10 source.t30 9.9005
R178 source.n10 source.t39 9.9005
R179 source.n12 source.t35 9.9005
R180 source.n12 source.t21 9.9005
R181 source.n14 source.t38 9.9005
R182 source.n14 source.t36 9.9005
R183 source.n32 source.t1 9.9005
R184 source.n32 source.t18 9.9005
R185 source.n34 source.t5 9.9005
R186 source.n34 source.t2 9.9005
R187 source.n36 source.t11 9.9005
R188 source.n36 source.t16 9.9005
R189 source.n38 source.t7 9.9005
R190 source.n38 source.t19 9.9005
R191 source.n91 source.n89 9.71174
R192 source.n75 source.n73 9.71174
R193 source.n67 source.n65 9.71174
R194 source.n51 source.n49 9.71174
R195 source.n3 source.n1 9.71174
R196 source.n19 source.n17 9.71174
R197 source.n27 source.n25 9.71174
R198 source.n43 source.n41 9.71174
R199 source.n94 source.n93 9.45567
R200 source.n78 source.n77 9.45567
R201 source.n70 source.n69 9.45567
R202 source.n54 source.n53 9.45567
R203 source.n6 source.n5 9.45567
R204 source.n22 source.n21 9.45567
R205 source.n30 source.n29 9.45567
R206 source.n46 source.n45 9.45567
R207 source.n93 source.n92 9.3005
R208 source.n77 source.n76 9.3005
R209 source.n69 source.n68 9.3005
R210 source.n53 source.n52 9.3005
R211 source.n5 source.n4 9.3005
R212 source.n21 source.n20 9.3005
R213 source.n29 source.n28 9.3005
R214 source.n45 source.n44 9.3005
R215 source.n96 source.n7 8.8499
R216 source.n94 source.n88 8.14595
R217 source.n78 source.n72 8.14595
R218 source.n70 source.n64 8.14595
R219 source.n54 source.n48 8.14595
R220 source.n6 source.n0 8.14595
R221 source.n22 source.n16 8.14595
R222 source.n30 source.n24 8.14595
R223 source.n46 source.n40 8.14595
R224 source.n92 source.n91 7.3702
R225 source.n76 source.n75 7.3702
R226 source.n68 source.n67 7.3702
R227 source.n52 source.n51 7.3702
R228 source.n4 source.n3 7.3702
R229 source.n20 source.n19 7.3702
R230 source.n28 source.n27 7.3702
R231 source.n44 source.n43 7.3702
R232 source.n92 source.n88 5.81868
R233 source.n76 source.n72 5.81868
R234 source.n68 source.n64 5.81868
R235 source.n52 source.n48 5.81868
R236 source.n4 source.n0 5.81868
R237 source.n20 source.n16 5.81868
R238 source.n28 source.n24 5.81868
R239 source.n44 source.n40 5.81868
R240 source.n96 source.n95 5.66429
R241 source.n93 source.n89 3.44771
R242 source.n77 source.n73 3.44771
R243 source.n69 source.n65 3.44771
R244 source.n53 source.n49 3.44771
R245 source.n5 source.n1 3.44771
R246 source.n21 source.n17 3.44771
R247 source.n29 source.n25 3.44771
R248 source.n45 source.n41 3.44771
R249 source.n47 source.n39 0.802224
R250 source.n39 source.n37 0.802224
R251 source.n37 source.n35 0.802224
R252 source.n35 source.n33 0.802224
R253 source.n33 source.n31 0.802224
R254 source.n23 source.n15 0.802224
R255 source.n15 source.n13 0.802224
R256 source.n13 source.n11 0.802224
R257 source.n11 source.n9 0.802224
R258 source.n9 source.n7 0.802224
R259 source.n57 source.n55 0.802224
R260 source.n59 source.n57 0.802224
R261 source.n61 source.n59 0.802224
R262 source.n63 source.n61 0.802224
R263 source.n71 source.n63 0.802224
R264 source.n81 source.n79 0.802224
R265 source.n83 source.n81 0.802224
R266 source.n85 source.n83 0.802224
R267 source.n87 source.n85 0.802224
R268 source.n95 source.n87 0.802224
R269 source.n31 source.n23 0.470328
R270 source.n79 source.n71 0.470328
R271 source source.n96 0.188
R272 drain_left.n10 drain_left.n8 101.597
R273 drain_left.n6 drain_left.n4 101.597
R274 drain_left.n2 drain_left.n0 101.597
R275 drain_left.n16 drain_left.n15 100.796
R276 drain_left.n14 drain_left.n13 100.796
R277 drain_left.n12 drain_left.n11 100.796
R278 drain_left.n10 drain_left.n9 100.796
R279 drain_left.n7 drain_left.n3 100.796
R280 drain_left.n6 drain_left.n5 100.796
R281 drain_left.n2 drain_left.n1 100.796
R282 drain_left drain_left.n7 26.2051
R283 drain_left.n3 drain_left.t2 9.9005
R284 drain_left.n3 drain_left.t0 9.9005
R285 drain_left.n4 drain_left.t8 9.9005
R286 drain_left.n4 drain_left.t1 9.9005
R287 drain_left.n5 drain_left.t13 9.9005
R288 drain_left.n5 drain_left.t11 9.9005
R289 drain_left.n1 drain_left.t12 9.9005
R290 drain_left.n1 drain_left.t10 9.9005
R291 drain_left.n0 drain_left.t5 9.9005
R292 drain_left.n0 drain_left.t18 9.9005
R293 drain_left.n15 drain_left.t17 9.9005
R294 drain_left.n15 drain_left.t19 9.9005
R295 drain_left.n13 drain_left.t15 9.9005
R296 drain_left.n13 drain_left.t16 9.9005
R297 drain_left.n11 drain_left.t9 9.9005
R298 drain_left.n11 drain_left.t14 9.9005
R299 drain_left.n9 drain_left.t6 9.9005
R300 drain_left.n9 drain_left.t7 9.9005
R301 drain_left.n8 drain_left.t3 9.9005
R302 drain_left.n8 drain_left.t4 9.9005
R303 drain_left drain_left.n16 6.45494
R304 drain_left.n12 drain_left.n10 0.802224
R305 drain_left.n14 drain_left.n12 0.802224
R306 drain_left.n16 drain_left.n14 0.802224
R307 drain_left.n7 drain_left.n6 0.746878
R308 drain_left.n7 drain_left.n2 0.746878
R309 minus.n6 minus.t15 172.626
R310 minus.n34 minus.t10 172.626
R311 minus.n27 minus.n26 161.3
R312 minus.n24 minus.n23 161.3
R313 minus.n22 minus.n1 161.3
R314 minus.n21 minus.n20 161.3
R315 minus.n19 minus.n2 161.3
R316 minus.n18 minus.n17 161.3
R317 minus.n16 minus.n3 161.3
R318 minus.n15 minus.n14 161.3
R319 minus.n13 minus.n4 161.3
R320 minus.n12 minus.n11 161.3
R321 minus.n10 minus.n5 161.3
R322 minus.n9 minus.n8 161.3
R323 minus.n55 minus.n54 161.3
R324 minus.n52 minus.n51 161.3
R325 minus.n50 minus.n29 161.3
R326 minus.n49 minus.n48 161.3
R327 minus.n47 minus.n30 161.3
R328 minus.n46 minus.n45 161.3
R329 minus.n44 minus.n31 161.3
R330 minus.n43 minus.n42 161.3
R331 minus.n41 minus.n32 161.3
R332 minus.n40 minus.n39 161.3
R333 minus.n38 minus.n33 161.3
R334 minus.n37 minus.n36 161.3
R335 minus.n7 minus.t14 145.805
R336 minus.n8 minus.t13 145.805
R337 minus.n12 minus.t12 145.805
R338 minus.n14 minus.t7 145.805
R339 minus.n18 minus.t11 145.805
R340 minus.n20 minus.t8 145.805
R341 minus.n24 minus.t4 145.805
R342 minus.n25 minus.t2 145.805
R343 minus.n26 minus.t1 145.805
R344 minus.n35 minus.t19 145.805
R345 minus.n36 minus.t17 145.805
R346 minus.n40 minus.t9 145.805
R347 minus.n42 minus.t3 145.805
R348 minus.n46 minus.t6 145.805
R349 minus.n48 minus.t18 145.805
R350 minus.n52 minus.t16 145.805
R351 minus.n53 minus.t5 145.805
R352 minus.n54 minus.t0 145.805
R353 minus.n25 minus.n0 80.6037
R354 minus.n53 minus.n28 80.6037
R355 minus.n8 minus.n7 48.2005
R356 minus.n25 minus.n24 48.2005
R357 minus.n26 minus.n25 48.2005
R358 minus.n36 minus.n35 48.2005
R359 minus.n53 minus.n52 48.2005
R360 minus.n54 minus.n53 48.2005
R361 minus.n9 minus.n6 45.1367
R362 minus.n37 minus.n34 45.1367
R363 minus.n12 minus.n5 44.549
R364 minus.n20 minus.n1 44.549
R365 minus.n40 minus.n33 44.549
R366 minus.n48 minus.n29 44.549
R367 minus.n14 minus.n13 34.3247
R368 minus.n19 minus.n18 34.3247
R369 minus.n42 minus.n41 34.3247
R370 minus.n47 minus.n46 34.3247
R371 minus.n56 minus.n27 32.1369
R372 minus.n18 minus.n3 24.1005
R373 minus.n14 minus.n3 24.1005
R374 minus.n42 minus.n31 24.1005
R375 minus.n46 minus.n31 24.1005
R376 minus.n13 minus.n12 13.8763
R377 minus.n20 minus.n19 13.8763
R378 minus.n41 minus.n40 13.8763
R379 minus.n48 minus.n47 13.8763
R380 minus.n7 minus.n6 13.3799
R381 minus.n35 minus.n34 13.3799
R382 minus.n56 minus.n55 6.62929
R383 minus.n8 minus.n5 3.65202
R384 minus.n24 minus.n1 3.65202
R385 minus.n36 minus.n33 3.65202
R386 minus.n52 minus.n29 3.65202
R387 minus.n27 minus.n0 0.285035
R388 minus.n23 minus.n0 0.285035
R389 minus.n51 minus.n28 0.285035
R390 minus.n55 minus.n28 0.285035
R391 minus.n23 minus.n22 0.189894
R392 minus.n22 minus.n21 0.189894
R393 minus.n21 minus.n2 0.189894
R394 minus.n17 minus.n2 0.189894
R395 minus.n17 minus.n16 0.189894
R396 minus.n16 minus.n15 0.189894
R397 minus.n15 minus.n4 0.189894
R398 minus.n11 minus.n4 0.189894
R399 minus.n11 minus.n10 0.189894
R400 minus.n10 minus.n9 0.189894
R401 minus.n38 minus.n37 0.189894
R402 minus.n39 minus.n38 0.189894
R403 minus.n39 minus.n32 0.189894
R404 minus.n43 minus.n32 0.189894
R405 minus.n44 minus.n43 0.189894
R406 minus.n45 minus.n44 0.189894
R407 minus.n45 minus.n30 0.189894
R408 minus.n49 minus.n30 0.189894
R409 minus.n50 minus.n49 0.189894
R410 minus.n51 minus.n50 0.189894
R411 minus minus.n56 0.188
R412 drain_right.n10 drain_right.n8 101.597
R413 drain_right.n6 drain_right.n4 101.597
R414 drain_right.n2 drain_right.n0 101.597
R415 drain_right.n10 drain_right.n9 100.796
R416 drain_right.n12 drain_right.n11 100.796
R417 drain_right.n14 drain_right.n13 100.796
R418 drain_right.n16 drain_right.n15 100.796
R419 drain_right.n7 drain_right.n3 100.796
R420 drain_right.n6 drain_right.n5 100.796
R421 drain_right.n2 drain_right.n1 100.796
R422 drain_right drain_right.n7 25.6519
R423 drain_right.n3 drain_right.t16 9.9005
R424 drain_right.n3 drain_right.t13 9.9005
R425 drain_right.n4 drain_right.t14 9.9005
R426 drain_right.n4 drain_right.t19 9.9005
R427 drain_right.n5 drain_right.t1 9.9005
R428 drain_right.n5 drain_right.t3 9.9005
R429 drain_right.n1 drain_right.t2 9.9005
R430 drain_right.n1 drain_right.t10 9.9005
R431 drain_right.n0 drain_right.t9 9.9005
R432 drain_right.n0 drain_right.t0 9.9005
R433 drain_right.n8 drain_right.t5 9.9005
R434 drain_right.n8 drain_right.t4 9.9005
R435 drain_right.n9 drain_right.t7 9.9005
R436 drain_right.n9 drain_right.t6 9.9005
R437 drain_right.n11 drain_right.t8 9.9005
R438 drain_right.n11 drain_right.t12 9.9005
R439 drain_right.n13 drain_right.t15 9.9005
R440 drain_right.n13 drain_right.t11 9.9005
R441 drain_right.n15 drain_right.t18 9.9005
R442 drain_right.n15 drain_right.t17 9.9005
R443 drain_right drain_right.n16 6.45494
R444 drain_right.n16 drain_right.n14 0.802224
R445 drain_right.n14 drain_right.n12 0.802224
R446 drain_right.n12 drain_right.n10 0.802224
R447 drain_right.n7 drain_right.n6 0.746878
R448 drain_right.n7 drain_right.n2 0.746878
C0 source drain_right 7.5894f
C1 source plus 3.10756f
C2 drain_right plus 0.438563f
C3 minus drain_left 0.179543f
C4 source minus 3.09359f
C5 minus drain_right 2.46985f
C6 minus plus 4.74895f
C7 source drain_left 7.58756f
C8 drain_right drain_left 1.48701f
C9 drain_left plus 2.74437f
C10 drain_right a_n2762_n1288# 5.1715f
C11 drain_left a_n2762_n1288# 5.56926f
C12 source a_n2762_n1288# 3.459466f
C13 minus a_n2762_n1288# 10.227885f
C14 plus a_n2762_n1288# 11.58139f
C15 drain_right.t9 a_n2762_n1288# 0.043534f
C16 drain_right.t0 a_n2762_n1288# 0.043534f
C17 drain_right.n0 a_n2762_n1288# 0.276369f
C18 drain_right.t2 a_n2762_n1288# 0.043534f
C19 drain_right.t10 a_n2762_n1288# 0.043534f
C20 drain_right.n1 a_n2762_n1288# 0.273494f
C21 drain_right.n2 a_n2762_n1288# 0.710454f
C22 drain_right.t16 a_n2762_n1288# 0.043534f
C23 drain_right.t13 a_n2762_n1288# 0.043534f
C24 drain_right.n3 a_n2762_n1288# 0.273494f
C25 drain_right.t14 a_n2762_n1288# 0.043534f
C26 drain_right.t19 a_n2762_n1288# 0.043534f
C27 drain_right.n4 a_n2762_n1288# 0.276369f
C28 drain_right.t1 a_n2762_n1288# 0.043534f
C29 drain_right.t3 a_n2762_n1288# 0.043534f
C30 drain_right.n5 a_n2762_n1288# 0.273494f
C31 drain_right.n6 a_n2762_n1288# 0.710454f
C32 drain_right.n7 a_n2762_n1288# 1.28576f
C33 drain_right.t5 a_n2762_n1288# 0.043534f
C34 drain_right.t4 a_n2762_n1288# 0.043534f
C35 drain_right.n8 a_n2762_n1288# 0.27637f
C36 drain_right.t7 a_n2762_n1288# 0.043534f
C37 drain_right.t6 a_n2762_n1288# 0.043534f
C38 drain_right.n9 a_n2762_n1288# 0.273495f
C39 drain_right.n10 a_n2762_n1288# 0.714508f
C40 drain_right.t8 a_n2762_n1288# 0.043534f
C41 drain_right.t12 a_n2762_n1288# 0.043534f
C42 drain_right.n11 a_n2762_n1288# 0.273495f
C43 drain_right.n12 a_n2762_n1288# 0.353144f
C44 drain_right.t15 a_n2762_n1288# 0.043534f
C45 drain_right.t11 a_n2762_n1288# 0.043534f
C46 drain_right.n13 a_n2762_n1288# 0.273495f
C47 drain_right.n14 a_n2762_n1288# 0.353144f
C48 drain_right.t18 a_n2762_n1288# 0.043534f
C49 drain_right.t17 a_n2762_n1288# 0.043534f
C50 drain_right.n15 a_n2762_n1288# 0.273495f
C51 drain_right.n16 a_n2762_n1288# 0.593335f
C52 minus.n0 a_n2762_n1288# 0.058152f
C53 minus.n1 a_n2762_n1288# 0.009912f
C54 minus.t4 a_n2762_n1288# 0.162327f
C55 minus.n2 a_n2762_n1288# 0.043682f
C56 minus.n3 a_n2762_n1288# 0.009912f
C57 minus.t11 a_n2762_n1288# 0.162327f
C58 minus.n4 a_n2762_n1288# 0.043682f
C59 minus.n5 a_n2762_n1288# 0.009912f
C60 minus.t12 a_n2762_n1288# 0.162327f
C61 minus.t15 a_n2762_n1288# 0.180206f
C62 minus.n6 a_n2762_n1288# 0.098007f
C63 minus.t14 a_n2762_n1288# 0.162327f
C64 minus.n7 a_n2762_n1288# 0.12486f
C65 minus.t13 a_n2762_n1288# 0.162327f
C66 minus.n8 a_n2762_n1288# 0.115621f
C67 minus.n9 a_n2762_n1288# 0.18645f
C68 minus.n10 a_n2762_n1288# 0.043682f
C69 minus.n11 a_n2762_n1288# 0.043682f
C70 minus.n12 a_n2762_n1288# 0.116833f
C71 minus.n13 a_n2762_n1288# 0.009912f
C72 minus.t7 a_n2762_n1288# 0.162327f
C73 minus.n14 a_n2762_n1288# 0.116833f
C74 minus.n15 a_n2762_n1288# 0.043682f
C75 minus.n16 a_n2762_n1288# 0.043682f
C76 minus.n17 a_n2762_n1288# 0.043682f
C77 minus.n18 a_n2762_n1288# 0.116833f
C78 minus.n19 a_n2762_n1288# 0.009912f
C79 minus.t8 a_n2762_n1288# 0.162327f
C80 minus.n20 a_n2762_n1288# 0.116833f
C81 minus.n21 a_n2762_n1288# 0.043682f
C82 minus.n22 a_n2762_n1288# 0.043682f
C83 minus.n23 a_n2762_n1288# 0.058289f
C84 minus.n24 a_n2762_n1288# 0.115621f
C85 minus.t2 a_n2762_n1288# 0.162327f
C86 minus.n25 a_n2762_n1288# 0.12486f
C87 minus.t1 a_n2762_n1288# 0.162327f
C88 minus.n26 a_n2762_n1288# 0.114948f
C89 minus.n27 a_n2762_n1288# 1.295f
C90 minus.n28 a_n2762_n1288# 0.058152f
C91 minus.n29 a_n2762_n1288# 0.009912f
C92 minus.n30 a_n2762_n1288# 0.043682f
C93 minus.n31 a_n2762_n1288# 0.009912f
C94 minus.n32 a_n2762_n1288# 0.043682f
C95 minus.n33 a_n2762_n1288# 0.009912f
C96 minus.t10 a_n2762_n1288# 0.180206f
C97 minus.n34 a_n2762_n1288# 0.098007f
C98 minus.t19 a_n2762_n1288# 0.162327f
C99 minus.n35 a_n2762_n1288# 0.12486f
C100 minus.t17 a_n2762_n1288# 0.162327f
C101 minus.n36 a_n2762_n1288# 0.115621f
C102 minus.n37 a_n2762_n1288# 0.18645f
C103 minus.n38 a_n2762_n1288# 0.043682f
C104 minus.n39 a_n2762_n1288# 0.043682f
C105 minus.t9 a_n2762_n1288# 0.162327f
C106 minus.n40 a_n2762_n1288# 0.116833f
C107 minus.n41 a_n2762_n1288# 0.009912f
C108 minus.t3 a_n2762_n1288# 0.162327f
C109 minus.n42 a_n2762_n1288# 0.116833f
C110 minus.n43 a_n2762_n1288# 0.043682f
C111 minus.n44 a_n2762_n1288# 0.043682f
C112 minus.n45 a_n2762_n1288# 0.043682f
C113 minus.t6 a_n2762_n1288# 0.162327f
C114 minus.n46 a_n2762_n1288# 0.116833f
C115 minus.n47 a_n2762_n1288# 0.009912f
C116 minus.t18 a_n2762_n1288# 0.162327f
C117 minus.n48 a_n2762_n1288# 0.116833f
C118 minus.n49 a_n2762_n1288# 0.043682f
C119 minus.n50 a_n2762_n1288# 0.043682f
C120 minus.n51 a_n2762_n1288# 0.058289f
C121 minus.t16 a_n2762_n1288# 0.162327f
C122 minus.n52 a_n2762_n1288# 0.115621f
C123 minus.t5 a_n2762_n1288# 0.162327f
C124 minus.n53 a_n2762_n1288# 0.12486f
C125 minus.t0 a_n2762_n1288# 0.162327f
C126 minus.n54 a_n2762_n1288# 0.114948f
C127 minus.n55 a_n2762_n1288# 0.313416f
C128 minus.n56 a_n2762_n1288# 1.56691f
C129 drain_left.t5 a_n2762_n1288# 0.043927f
C130 drain_left.t18 a_n2762_n1288# 0.043927f
C131 drain_left.n0 a_n2762_n1288# 0.278866f
C132 drain_left.t12 a_n2762_n1288# 0.043927f
C133 drain_left.t10 a_n2762_n1288# 0.043927f
C134 drain_left.n1 a_n2762_n1288# 0.275966f
C135 drain_left.n2 a_n2762_n1288# 0.716874f
C136 drain_left.t2 a_n2762_n1288# 0.043927f
C137 drain_left.t0 a_n2762_n1288# 0.043927f
C138 drain_left.n3 a_n2762_n1288# 0.275966f
C139 drain_left.t8 a_n2762_n1288# 0.043927f
C140 drain_left.t1 a_n2762_n1288# 0.043927f
C141 drain_left.n4 a_n2762_n1288# 0.278866f
C142 drain_left.t13 a_n2762_n1288# 0.043927f
C143 drain_left.t11 a_n2762_n1288# 0.043927f
C144 drain_left.n5 a_n2762_n1288# 0.275966f
C145 drain_left.n6 a_n2762_n1288# 0.716874f
C146 drain_left.n7 a_n2762_n1288# 1.35136f
C147 drain_left.t3 a_n2762_n1288# 0.043927f
C148 drain_left.t4 a_n2762_n1288# 0.043927f
C149 drain_left.n8 a_n2762_n1288# 0.278867f
C150 drain_left.t6 a_n2762_n1288# 0.043927f
C151 drain_left.t7 a_n2762_n1288# 0.043927f
C152 drain_left.n9 a_n2762_n1288# 0.275967f
C153 drain_left.n10 a_n2762_n1288# 0.720965f
C154 drain_left.t9 a_n2762_n1288# 0.043927f
C155 drain_left.t14 a_n2762_n1288# 0.043927f
C156 drain_left.n11 a_n2762_n1288# 0.275967f
C157 drain_left.n12 a_n2762_n1288# 0.356335f
C158 drain_left.t15 a_n2762_n1288# 0.043927f
C159 drain_left.t16 a_n2762_n1288# 0.043927f
C160 drain_left.n13 a_n2762_n1288# 0.275967f
C161 drain_left.n14 a_n2762_n1288# 0.356335f
C162 drain_left.t17 a_n2762_n1288# 0.043927f
C163 drain_left.t19 a_n2762_n1288# 0.043927f
C164 drain_left.n15 a_n2762_n1288# 0.275967f
C165 drain_left.n16 a_n2762_n1288# 0.598697f
C166 source.n0 a_n2762_n1288# 0.046141f
C167 source.n1 a_n2762_n1288# 0.102093f
C168 source.t29 a_n2762_n1288# 0.076616f
C169 source.n2 a_n2762_n1288# 0.079902f
C170 source.n3 a_n2762_n1288# 0.025757f
C171 source.n4 a_n2762_n1288# 0.016987f
C172 source.n5 a_n2762_n1288# 0.225039f
C173 source.n6 a_n2762_n1288# 0.050582f
C174 source.n7 a_n2762_n1288# 0.524017f
C175 source.t27 a_n2762_n1288# 0.049963f
C176 source.t28 a_n2762_n1288# 0.049963f
C177 source.n8 a_n2762_n1288# 0.267102f
C178 source.n9 a_n2762_n1288# 0.409112f
C179 source.t30 a_n2762_n1288# 0.049963f
C180 source.t39 a_n2762_n1288# 0.049963f
C181 source.n10 a_n2762_n1288# 0.267102f
C182 source.n11 a_n2762_n1288# 0.409112f
C183 source.t35 a_n2762_n1288# 0.049963f
C184 source.t21 a_n2762_n1288# 0.049963f
C185 source.n12 a_n2762_n1288# 0.267102f
C186 source.n13 a_n2762_n1288# 0.409112f
C187 source.t38 a_n2762_n1288# 0.049963f
C188 source.t36 a_n2762_n1288# 0.049963f
C189 source.n14 a_n2762_n1288# 0.267102f
C190 source.n15 a_n2762_n1288# 0.409112f
C191 source.n16 a_n2762_n1288# 0.046141f
C192 source.n17 a_n2762_n1288# 0.102093f
C193 source.t37 a_n2762_n1288# 0.076616f
C194 source.n18 a_n2762_n1288# 0.079902f
C195 source.n19 a_n2762_n1288# 0.025757f
C196 source.n20 a_n2762_n1288# 0.016987f
C197 source.n21 a_n2762_n1288# 0.225039f
C198 source.n22 a_n2762_n1288# 0.050582f
C199 source.n23 a_n2762_n1288# 0.155551f
C200 source.n24 a_n2762_n1288# 0.046141f
C201 source.n25 a_n2762_n1288# 0.102093f
C202 source.t4 a_n2762_n1288# 0.076616f
C203 source.n26 a_n2762_n1288# 0.079902f
C204 source.n27 a_n2762_n1288# 0.025757f
C205 source.n28 a_n2762_n1288# 0.016987f
C206 source.n29 a_n2762_n1288# 0.225039f
C207 source.n30 a_n2762_n1288# 0.050582f
C208 source.n31 a_n2762_n1288# 0.155551f
C209 source.t1 a_n2762_n1288# 0.049963f
C210 source.t18 a_n2762_n1288# 0.049963f
C211 source.n32 a_n2762_n1288# 0.267102f
C212 source.n33 a_n2762_n1288# 0.409112f
C213 source.t5 a_n2762_n1288# 0.049963f
C214 source.t2 a_n2762_n1288# 0.049963f
C215 source.n34 a_n2762_n1288# 0.267102f
C216 source.n35 a_n2762_n1288# 0.409112f
C217 source.t11 a_n2762_n1288# 0.049963f
C218 source.t16 a_n2762_n1288# 0.049963f
C219 source.n36 a_n2762_n1288# 0.267102f
C220 source.n37 a_n2762_n1288# 0.409112f
C221 source.t7 a_n2762_n1288# 0.049963f
C222 source.t19 a_n2762_n1288# 0.049963f
C223 source.n38 a_n2762_n1288# 0.267102f
C224 source.n39 a_n2762_n1288# 0.409112f
C225 source.n40 a_n2762_n1288# 0.046141f
C226 source.n41 a_n2762_n1288# 0.102093f
C227 source.t13 a_n2762_n1288# 0.076616f
C228 source.n42 a_n2762_n1288# 0.079902f
C229 source.n43 a_n2762_n1288# 0.025757f
C230 source.n44 a_n2762_n1288# 0.016987f
C231 source.n45 a_n2762_n1288# 0.225039f
C232 source.n46 a_n2762_n1288# 0.050582f
C233 source.n47 a_n2762_n1288# 0.824725f
C234 source.n48 a_n2762_n1288# 0.046141f
C235 source.n49 a_n2762_n1288# 0.102093f
C236 source.t24 a_n2762_n1288# 0.076616f
C237 source.n50 a_n2762_n1288# 0.079902f
C238 source.n51 a_n2762_n1288# 0.025757f
C239 source.n52 a_n2762_n1288# 0.016987f
C240 source.n53 a_n2762_n1288# 0.225039f
C241 source.n54 a_n2762_n1288# 0.050582f
C242 source.n55 a_n2762_n1288# 0.824725f
C243 source.t26 a_n2762_n1288# 0.049963f
C244 source.t22 a_n2762_n1288# 0.049963f
C245 source.n56 a_n2762_n1288# 0.267101f
C246 source.n57 a_n2762_n1288# 0.409113f
C247 source.t33 a_n2762_n1288# 0.049963f
C248 source.t31 a_n2762_n1288# 0.049963f
C249 source.n58 a_n2762_n1288# 0.267101f
C250 source.n59 a_n2762_n1288# 0.409113f
C251 source.t20 a_n2762_n1288# 0.049963f
C252 source.t25 a_n2762_n1288# 0.049963f
C253 source.n60 a_n2762_n1288# 0.267101f
C254 source.n61 a_n2762_n1288# 0.409113f
C255 source.t32 a_n2762_n1288# 0.049963f
C256 source.t34 a_n2762_n1288# 0.049963f
C257 source.n62 a_n2762_n1288# 0.267101f
C258 source.n63 a_n2762_n1288# 0.409113f
C259 source.n64 a_n2762_n1288# 0.046141f
C260 source.n65 a_n2762_n1288# 0.102093f
C261 source.t23 a_n2762_n1288# 0.076616f
C262 source.n66 a_n2762_n1288# 0.079902f
C263 source.n67 a_n2762_n1288# 0.025757f
C264 source.n68 a_n2762_n1288# 0.016987f
C265 source.n69 a_n2762_n1288# 0.225039f
C266 source.n70 a_n2762_n1288# 0.050582f
C267 source.n71 a_n2762_n1288# 0.155551f
C268 source.n72 a_n2762_n1288# 0.046141f
C269 source.n73 a_n2762_n1288# 0.102093f
C270 source.t0 a_n2762_n1288# 0.076616f
C271 source.n74 a_n2762_n1288# 0.079902f
C272 source.n75 a_n2762_n1288# 0.025757f
C273 source.n76 a_n2762_n1288# 0.016987f
C274 source.n77 a_n2762_n1288# 0.225039f
C275 source.n78 a_n2762_n1288# 0.050582f
C276 source.n79 a_n2762_n1288# 0.155551f
C277 source.t15 a_n2762_n1288# 0.049963f
C278 source.t6 a_n2762_n1288# 0.049963f
C279 source.n80 a_n2762_n1288# 0.267101f
C280 source.n81 a_n2762_n1288# 0.409113f
C281 source.t14 a_n2762_n1288# 0.049963f
C282 source.t8 a_n2762_n1288# 0.049963f
C283 source.n82 a_n2762_n1288# 0.267101f
C284 source.n83 a_n2762_n1288# 0.409113f
C285 source.t3 a_n2762_n1288# 0.049963f
C286 source.t12 a_n2762_n1288# 0.049963f
C287 source.n84 a_n2762_n1288# 0.267101f
C288 source.n85 a_n2762_n1288# 0.409113f
C289 source.t17 a_n2762_n1288# 0.049963f
C290 source.t10 a_n2762_n1288# 0.049963f
C291 source.n86 a_n2762_n1288# 0.267101f
C292 source.n87 a_n2762_n1288# 0.409113f
C293 source.n88 a_n2762_n1288# 0.046141f
C294 source.n89 a_n2762_n1288# 0.102093f
C295 source.t9 a_n2762_n1288# 0.076616f
C296 source.n90 a_n2762_n1288# 0.079902f
C297 source.n91 a_n2762_n1288# 0.025757f
C298 source.n92 a_n2762_n1288# 0.016987f
C299 source.n93 a_n2762_n1288# 0.225039f
C300 source.n94 a_n2762_n1288# 0.050582f
C301 source.n95 a_n2762_n1288# 0.354883f
C302 source.n96 a_n2762_n1288# 0.793036f
C303 plus.n0 a_n2762_n1288# 0.059794f
C304 plus.t0 a_n2762_n1288# 0.166911f
C305 plus.t2 a_n2762_n1288# 0.166911f
C306 plus.t3 a_n2762_n1288# 0.166911f
C307 plus.n1 a_n2762_n1288# 0.059935f
C308 plus.t4 a_n2762_n1288# 0.166911f
C309 plus.n2 a_n2762_n1288# 0.120132f
C310 plus.n3 a_n2762_n1288# 0.044916f
C311 plus.t5 a_n2762_n1288# 0.166911f
C312 plus.t10 a_n2762_n1288# 0.166911f
C313 plus.n4 a_n2762_n1288# 0.120132f
C314 plus.n5 a_n2762_n1288# 0.044916f
C315 plus.t12 a_n2762_n1288# 0.166911f
C316 plus.t13 a_n2762_n1288# 0.166911f
C317 plus.n6 a_n2762_n1288# 0.118886f
C318 plus.t15 a_n2762_n1288# 0.166911f
C319 plus.n7 a_n2762_n1288# 0.128386f
C320 plus.t16 a_n2762_n1288# 0.185294f
C321 plus.n8 a_n2762_n1288# 0.100774f
C322 plus.n9 a_n2762_n1288# 0.191715f
C323 plus.n10 a_n2762_n1288# 0.044916f
C324 plus.n11 a_n2762_n1288# 0.010192f
C325 plus.n12 a_n2762_n1288# 0.120132f
C326 plus.n13 a_n2762_n1288# 0.010192f
C327 plus.n14 a_n2762_n1288# 0.044916f
C328 plus.n15 a_n2762_n1288# 0.044916f
C329 plus.n16 a_n2762_n1288# 0.044916f
C330 plus.n17 a_n2762_n1288# 0.010192f
C331 plus.n18 a_n2762_n1288# 0.120132f
C332 plus.n19 a_n2762_n1288# 0.010192f
C333 plus.n20 a_n2762_n1288# 0.044916f
C334 plus.n21 a_n2762_n1288# 0.044916f
C335 plus.n22 a_n2762_n1288# 0.044916f
C336 plus.n23 a_n2762_n1288# 0.010192f
C337 plus.n24 a_n2762_n1288# 0.118886f
C338 plus.n25 a_n2762_n1288# 0.128386f
C339 plus.n26 a_n2762_n1288# 0.118193f
C340 plus.n27 a_n2762_n1288# 0.350459f
C341 plus.n28 a_n2762_n1288# 0.059794f
C342 plus.t14 a_n2762_n1288# 0.166911f
C343 plus.t1 a_n2762_n1288# 0.166911f
C344 plus.n29 a_n2762_n1288# 0.059935f
C345 plus.t7 a_n2762_n1288# 0.166911f
C346 plus.t9 a_n2762_n1288# 0.166911f
C347 plus.n30 a_n2762_n1288# 0.120132f
C348 plus.n31 a_n2762_n1288# 0.044916f
C349 plus.t17 a_n2762_n1288# 0.166911f
C350 plus.t19 a_n2762_n1288# 0.166911f
C351 plus.n32 a_n2762_n1288# 0.120132f
C352 plus.n33 a_n2762_n1288# 0.044916f
C353 plus.t6 a_n2762_n1288# 0.166911f
C354 plus.t8 a_n2762_n1288# 0.166911f
C355 plus.n34 a_n2762_n1288# 0.118886f
C356 plus.t11 a_n2762_n1288# 0.166911f
C357 plus.n35 a_n2762_n1288# 0.128386f
C358 plus.t18 a_n2762_n1288# 0.185294f
C359 plus.n36 a_n2762_n1288# 0.100774f
C360 plus.n37 a_n2762_n1288# 0.191715f
C361 plus.n38 a_n2762_n1288# 0.044916f
C362 plus.n39 a_n2762_n1288# 0.010192f
C363 plus.n40 a_n2762_n1288# 0.120132f
C364 plus.n41 a_n2762_n1288# 0.010192f
C365 plus.n42 a_n2762_n1288# 0.044916f
C366 plus.n43 a_n2762_n1288# 0.044916f
C367 plus.n44 a_n2762_n1288# 0.044916f
C368 plus.n45 a_n2762_n1288# 0.010192f
C369 plus.n46 a_n2762_n1288# 0.120132f
C370 plus.n47 a_n2762_n1288# 0.010192f
C371 plus.n48 a_n2762_n1288# 0.044916f
C372 plus.n49 a_n2762_n1288# 0.044916f
C373 plus.n50 a_n2762_n1288# 0.044916f
C374 plus.n51 a_n2762_n1288# 0.010192f
C375 plus.n52 a_n2762_n1288# 0.118886f
C376 plus.n53 a_n2762_n1288# 0.128386f
C377 plus.n54 a_n2762_n1288# 0.118193f
C378 plus.n55 a_n2762_n1288# 1.2669f
.ends

