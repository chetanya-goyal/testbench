* NGSPICE file created from diffpair479.ext - technology: sky130A

.subckt diffpair479 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t22 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X1 drain_right.t22 minus.t1 source.t26 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X2 a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X3 source.t5 plus.t0 drain_left.t23 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X4 drain_right.t21 minus.t2 source.t31 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X5 drain_right.t20 minus.t3 source.t38 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X6 a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X7 source.t10 plus.t1 drain_left.t22 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X8 source.t28 minus.t4 drain_right.t19 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X9 source.t7 plus.t2 drain_left.t21 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X10 drain_left.t20 plus.t3 source.t44 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X11 source.t35 minus.t5 drain_right.t18 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X12 drain_left.t19 plus.t4 source.t15 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X13 drain_left.t18 plus.t5 source.t16 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X14 drain_right.t17 minus.t6 source.t20 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X15 drain_left.t17 plus.t6 source.t47 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X16 source.t2 plus.t7 drain_left.t16 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X17 drain_right.t16 minus.t7 source.t43 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X18 drain_left.t15 plus.t8 source.t17 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X19 source.t32 minus.t8 drain_right.t15 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X20 source.t42 minus.t9 drain_right.t14 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X21 drain_right.t13 minus.t10 source.t41 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X22 drain_right.t12 minus.t11 source.t30 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X23 drain_right.t11 minus.t12 source.t29 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X24 source.t14 plus.t9 drain_left.t14 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X25 source.t36 minus.t13 drain_right.t10 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X26 drain_left.t13 plus.t10 source.t12 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X27 drain_left.t12 plus.t11 source.t4 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X28 source.t23 minus.t14 drain_right.t9 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X29 drain_right.t8 minus.t15 source.t25 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X30 drain_left.t11 plus.t12 source.t18 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X31 drain_right.t7 minus.t16 source.t39 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X32 source.t37 minus.t17 drain_right.t6 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X33 source.t0 plus.t13 drain_left.t10 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X34 a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X35 source.t40 minus.t18 drain_right.t5 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X36 source.t21 minus.t19 drain_right.t4 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X37 drain_left.t9 plus.t14 source.t46 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X38 drain_left.t8 plus.t15 source.t45 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X39 source.t33 minus.t20 drain_right.t3 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X40 source.t8 plus.t16 drain_left.t7 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X41 source.t13 plus.t17 drain_left.t6 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X42 drain_left.t5 plus.t18 source.t6 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X43 source.t1 plus.t19 drain_left.t4 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X44 drain_left.t3 plus.t20 source.t3 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X45 drain_right.t2 minus.t21 source.t34 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X46 a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X47 source.t27 minus.t22 drain_right.t1 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X48 source.t9 plus.t21 drain_left.t2 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X49 source.t24 minus.t23 drain_right.t0 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X50 source.t19 plus.t22 drain_left.t1 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X51 source.t11 plus.t23 drain_left.t0 a_n3654_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
R0 minus.n8 minus.t12 432.041
R1 minus.n44 minus.t23 432.041
R2 minus.n9 minus.t8 410.604
R3 minus.n10 minus.t7 410.604
R4 minus.n14 minus.t14 410.604
R5 minus.n16 minus.t16 410.604
R6 minus.n20 minus.t13 410.604
R7 minus.n21 minus.t10 410.604
R8 minus.n3 minus.t20 410.604
R9 minus.n27 minus.t15 410.604
R10 minus.n1 minus.t5 410.604
R11 minus.n32 minus.t11 410.604
R12 minus.n34 minus.t9 410.604
R13 minus.n45 minus.t6 410.604
R14 minus.n46 minus.t19 410.604
R15 minus.n50 minus.t3 410.604
R16 minus.n52 minus.t22 410.604
R17 minus.n56 minus.t2 410.604
R18 minus.n57 minus.t17 410.604
R19 minus.n39 minus.t0 410.604
R20 minus.n63 minus.t18 410.604
R21 minus.n37 minus.t1 410.604
R22 minus.n68 minus.t4 410.604
R23 minus.n70 minus.t21 410.604
R24 minus.n35 minus.n34 161.3
R25 minus.n33 minus.n0 161.3
R26 minus.n29 minus.n28 161.3
R27 minus.n27 minus.n2 161.3
R28 minus.n26 minus.n25 161.3
R29 minus.n24 minus.n3 161.3
R30 minus.n23 minus.n22 161.3
R31 minus.n18 minus.n5 161.3
R32 minus.n17 minus.n16 161.3
R33 minus.n15 minus.n6 161.3
R34 minus.n14 minus.n13 161.3
R35 minus.n12 minus.n7 161.3
R36 minus.n71 minus.n70 161.3
R37 minus.n69 minus.n36 161.3
R38 minus.n65 minus.n64 161.3
R39 minus.n63 minus.n38 161.3
R40 minus.n62 minus.n61 161.3
R41 minus.n60 minus.n39 161.3
R42 minus.n59 minus.n58 161.3
R43 minus.n54 minus.n41 161.3
R44 minus.n53 minus.n52 161.3
R45 minus.n51 minus.n42 161.3
R46 minus.n50 minus.n49 161.3
R47 minus.n48 minus.n43 161.3
R48 minus.n32 minus.n31 80.6037
R49 minus.n30 minus.n1 80.6037
R50 minus.n21 minus.n4 80.6037
R51 minus.n20 minus.n19 80.6037
R52 minus.n11 minus.n10 80.6037
R53 minus.n68 minus.n67 80.6037
R54 minus.n66 minus.n37 80.6037
R55 minus.n57 minus.n40 80.6037
R56 minus.n56 minus.n55 80.6037
R57 minus.n47 minus.n46 80.6037
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n72 minus.n35 43.1217
R69 minus.n20 minus.n5 41.6278
R70 minus.n22 minus.n21 41.6278
R71 minus.n56 minus.n41 41.6278
R72 minus.n58 minus.n57 41.6278
R73 minus.n33 minus.n32 38.7066
R74 minus.n69 minus.n68 38.7066
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 source.n562 source.n502 289.615
R132 source.n486 source.n426 289.615
R133 source.n420 source.n360 289.615
R134 source.n344 source.n284 289.615
R135 source.n60 source.n0 289.615
R136 source.n136 source.n76 289.615
R137 source.n202 source.n142 289.615
R138 source.n278 source.n218 289.615
R139 source.n522 source.n521 185
R140 source.n527 source.n526 185
R141 source.n529 source.n528 185
R142 source.n518 source.n517 185
R143 source.n535 source.n534 185
R144 source.n537 source.n536 185
R145 source.n514 source.n513 185
R146 source.n544 source.n543 185
R147 source.n545 source.n512 185
R148 source.n547 source.n546 185
R149 source.n510 source.n509 185
R150 source.n553 source.n552 185
R151 source.n555 source.n554 185
R152 source.n506 source.n505 185
R153 source.n561 source.n560 185
R154 source.n563 source.n562 185
R155 source.n446 source.n445 185
R156 source.n451 source.n450 185
R157 source.n453 source.n452 185
R158 source.n442 source.n441 185
R159 source.n459 source.n458 185
R160 source.n461 source.n460 185
R161 source.n438 source.n437 185
R162 source.n468 source.n467 185
R163 source.n469 source.n436 185
R164 source.n471 source.n470 185
R165 source.n434 source.n433 185
R166 source.n477 source.n476 185
R167 source.n479 source.n478 185
R168 source.n430 source.n429 185
R169 source.n485 source.n484 185
R170 source.n487 source.n486 185
R171 source.n380 source.n379 185
R172 source.n385 source.n384 185
R173 source.n387 source.n386 185
R174 source.n376 source.n375 185
R175 source.n393 source.n392 185
R176 source.n395 source.n394 185
R177 source.n372 source.n371 185
R178 source.n402 source.n401 185
R179 source.n403 source.n370 185
R180 source.n405 source.n404 185
R181 source.n368 source.n367 185
R182 source.n411 source.n410 185
R183 source.n413 source.n412 185
R184 source.n364 source.n363 185
R185 source.n419 source.n418 185
R186 source.n421 source.n420 185
R187 source.n304 source.n303 185
R188 source.n309 source.n308 185
R189 source.n311 source.n310 185
R190 source.n300 source.n299 185
R191 source.n317 source.n316 185
R192 source.n319 source.n318 185
R193 source.n296 source.n295 185
R194 source.n326 source.n325 185
R195 source.n327 source.n294 185
R196 source.n329 source.n328 185
R197 source.n292 source.n291 185
R198 source.n335 source.n334 185
R199 source.n337 source.n336 185
R200 source.n288 source.n287 185
R201 source.n343 source.n342 185
R202 source.n345 source.n344 185
R203 source.n61 source.n60 185
R204 source.n59 source.n58 185
R205 source.n4 source.n3 185
R206 source.n53 source.n52 185
R207 source.n51 source.n50 185
R208 source.n8 source.n7 185
R209 source.n45 source.n44 185
R210 source.n43 source.n10 185
R211 source.n42 source.n41 185
R212 source.n13 source.n11 185
R213 source.n36 source.n35 185
R214 source.n34 source.n33 185
R215 source.n17 source.n16 185
R216 source.n28 source.n27 185
R217 source.n26 source.n25 185
R218 source.n21 source.n20 185
R219 source.n137 source.n136 185
R220 source.n135 source.n134 185
R221 source.n80 source.n79 185
R222 source.n129 source.n128 185
R223 source.n127 source.n126 185
R224 source.n84 source.n83 185
R225 source.n121 source.n120 185
R226 source.n119 source.n86 185
R227 source.n118 source.n117 185
R228 source.n89 source.n87 185
R229 source.n112 source.n111 185
R230 source.n110 source.n109 185
R231 source.n93 source.n92 185
R232 source.n104 source.n103 185
R233 source.n102 source.n101 185
R234 source.n97 source.n96 185
R235 source.n203 source.n202 185
R236 source.n201 source.n200 185
R237 source.n146 source.n145 185
R238 source.n195 source.n194 185
R239 source.n193 source.n192 185
R240 source.n150 source.n149 185
R241 source.n187 source.n186 185
R242 source.n185 source.n152 185
R243 source.n184 source.n183 185
R244 source.n155 source.n153 185
R245 source.n178 source.n177 185
R246 source.n176 source.n175 185
R247 source.n159 source.n158 185
R248 source.n170 source.n169 185
R249 source.n168 source.n167 185
R250 source.n163 source.n162 185
R251 source.n279 source.n278 185
R252 source.n277 source.n276 185
R253 source.n222 source.n221 185
R254 source.n271 source.n270 185
R255 source.n269 source.n268 185
R256 source.n226 source.n225 185
R257 source.n263 source.n262 185
R258 source.n261 source.n228 185
R259 source.n260 source.n259 185
R260 source.n231 source.n229 185
R261 source.n254 source.n253 185
R262 source.n252 source.n251 185
R263 source.n235 source.n234 185
R264 source.n246 source.n245 185
R265 source.n244 source.n243 185
R266 source.n239 source.n238 185
R267 source.n523 source.t34 149.524
R268 source.n447 source.t24 149.524
R269 source.n381 source.t6 149.524
R270 source.n305 source.t11 149.524
R271 source.n22 source.t15 149.524
R272 source.n98 source.t9 149.524
R273 source.n164 source.t29 149.524
R274 source.n240 source.t42 149.524
R275 source.n527 source.n521 104.615
R276 source.n528 source.n527 104.615
R277 source.n528 source.n517 104.615
R278 source.n535 source.n517 104.615
R279 source.n536 source.n535 104.615
R280 source.n536 source.n513 104.615
R281 source.n544 source.n513 104.615
R282 source.n545 source.n544 104.615
R283 source.n546 source.n545 104.615
R284 source.n546 source.n509 104.615
R285 source.n553 source.n509 104.615
R286 source.n554 source.n553 104.615
R287 source.n554 source.n505 104.615
R288 source.n561 source.n505 104.615
R289 source.n562 source.n561 104.615
R290 source.n451 source.n445 104.615
R291 source.n452 source.n451 104.615
R292 source.n452 source.n441 104.615
R293 source.n459 source.n441 104.615
R294 source.n460 source.n459 104.615
R295 source.n460 source.n437 104.615
R296 source.n468 source.n437 104.615
R297 source.n469 source.n468 104.615
R298 source.n470 source.n469 104.615
R299 source.n470 source.n433 104.615
R300 source.n477 source.n433 104.615
R301 source.n478 source.n477 104.615
R302 source.n478 source.n429 104.615
R303 source.n485 source.n429 104.615
R304 source.n486 source.n485 104.615
R305 source.n385 source.n379 104.615
R306 source.n386 source.n385 104.615
R307 source.n386 source.n375 104.615
R308 source.n393 source.n375 104.615
R309 source.n394 source.n393 104.615
R310 source.n394 source.n371 104.615
R311 source.n402 source.n371 104.615
R312 source.n403 source.n402 104.615
R313 source.n404 source.n403 104.615
R314 source.n404 source.n367 104.615
R315 source.n411 source.n367 104.615
R316 source.n412 source.n411 104.615
R317 source.n412 source.n363 104.615
R318 source.n419 source.n363 104.615
R319 source.n420 source.n419 104.615
R320 source.n309 source.n303 104.615
R321 source.n310 source.n309 104.615
R322 source.n310 source.n299 104.615
R323 source.n317 source.n299 104.615
R324 source.n318 source.n317 104.615
R325 source.n318 source.n295 104.615
R326 source.n326 source.n295 104.615
R327 source.n327 source.n326 104.615
R328 source.n328 source.n327 104.615
R329 source.n328 source.n291 104.615
R330 source.n335 source.n291 104.615
R331 source.n336 source.n335 104.615
R332 source.n336 source.n287 104.615
R333 source.n343 source.n287 104.615
R334 source.n344 source.n343 104.615
R335 source.n60 source.n59 104.615
R336 source.n59 source.n3 104.615
R337 source.n52 source.n3 104.615
R338 source.n52 source.n51 104.615
R339 source.n51 source.n7 104.615
R340 source.n44 source.n7 104.615
R341 source.n44 source.n43 104.615
R342 source.n43 source.n42 104.615
R343 source.n42 source.n11 104.615
R344 source.n35 source.n11 104.615
R345 source.n35 source.n34 104.615
R346 source.n34 source.n16 104.615
R347 source.n27 source.n16 104.615
R348 source.n27 source.n26 104.615
R349 source.n26 source.n20 104.615
R350 source.n136 source.n135 104.615
R351 source.n135 source.n79 104.615
R352 source.n128 source.n79 104.615
R353 source.n128 source.n127 104.615
R354 source.n127 source.n83 104.615
R355 source.n120 source.n83 104.615
R356 source.n120 source.n119 104.615
R357 source.n119 source.n118 104.615
R358 source.n118 source.n87 104.615
R359 source.n111 source.n87 104.615
R360 source.n111 source.n110 104.615
R361 source.n110 source.n92 104.615
R362 source.n103 source.n92 104.615
R363 source.n103 source.n102 104.615
R364 source.n102 source.n96 104.615
R365 source.n202 source.n201 104.615
R366 source.n201 source.n145 104.615
R367 source.n194 source.n145 104.615
R368 source.n194 source.n193 104.615
R369 source.n193 source.n149 104.615
R370 source.n186 source.n149 104.615
R371 source.n186 source.n185 104.615
R372 source.n185 source.n184 104.615
R373 source.n184 source.n153 104.615
R374 source.n177 source.n153 104.615
R375 source.n177 source.n176 104.615
R376 source.n176 source.n158 104.615
R377 source.n169 source.n158 104.615
R378 source.n169 source.n168 104.615
R379 source.n168 source.n162 104.615
R380 source.n278 source.n277 104.615
R381 source.n277 source.n221 104.615
R382 source.n270 source.n221 104.615
R383 source.n270 source.n269 104.615
R384 source.n269 source.n225 104.615
R385 source.n262 source.n225 104.615
R386 source.n262 source.n261 104.615
R387 source.n261 source.n260 104.615
R388 source.n260 source.n229 104.615
R389 source.n253 source.n229 104.615
R390 source.n253 source.n252 104.615
R391 source.n252 source.n234 104.615
R392 source.n245 source.n234 104.615
R393 source.n245 source.n244 104.615
R394 source.n244 source.n238 104.615
R395 source.t34 source.n521 52.3082
R396 source.t24 source.n445 52.3082
R397 source.t6 source.n379 52.3082
R398 source.t11 source.n303 52.3082
R399 source.t15 source.n20 52.3082
R400 source.t9 source.n96 52.3082
R401 source.t29 source.n162 52.3082
R402 source.t42 source.n238 52.3082
R403 source.n67 source.n66 42.8739
R404 source.n69 source.n68 42.8739
R405 source.n71 source.n70 42.8739
R406 source.n73 source.n72 42.8739
R407 source.n75 source.n74 42.8739
R408 source.n209 source.n208 42.8739
R409 source.n211 source.n210 42.8739
R410 source.n213 source.n212 42.8739
R411 source.n215 source.n214 42.8739
R412 source.n217 source.n216 42.8739
R413 source.n501 source.n500 42.8737
R414 source.n499 source.n498 42.8737
R415 source.n497 source.n496 42.8737
R416 source.n495 source.n494 42.8737
R417 source.n493 source.n492 42.8737
R418 source.n359 source.n358 42.8737
R419 source.n357 source.n356 42.8737
R420 source.n355 source.n354 42.8737
R421 source.n353 source.n352 42.8737
R422 source.n351 source.n350 42.8737
R423 source.n567 source.n566 29.8581
R424 source.n491 source.n490 29.8581
R425 source.n425 source.n424 29.8581
R426 source.n349 source.n348 29.8581
R427 source.n65 source.n64 29.8581
R428 source.n141 source.n140 29.8581
R429 source.n207 source.n206 29.8581
R430 source.n283 source.n282 29.8581
R431 source.n349 source.n283 22.2619
R432 source.n568 source.n65 16.5119
R433 source.n547 source.n512 13.1884
R434 source.n471 source.n436 13.1884
R435 source.n405 source.n370 13.1884
R436 source.n329 source.n294 13.1884
R437 source.n45 source.n10 13.1884
R438 source.n121 source.n86 13.1884
R439 source.n187 source.n152 13.1884
R440 source.n263 source.n228 13.1884
R441 source.n543 source.n542 12.8005
R442 source.n548 source.n510 12.8005
R443 source.n467 source.n466 12.8005
R444 source.n472 source.n434 12.8005
R445 source.n401 source.n400 12.8005
R446 source.n406 source.n368 12.8005
R447 source.n325 source.n324 12.8005
R448 source.n330 source.n292 12.8005
R449 source.n46 source.n8 12.8005
R450 source.n41 source.n12 12.8005
R451 source.n122 source.n84 12.8005
R452 source.n117 source.n88 12.8005
R453 source.n188 source.n150 12.8005
R454 source.n183 source.n154 12.8005
R455 source.n264 source.n226 12.8005
R456 source.n259 source.n230 12.8005
R457 source.n541 source.n514 12.0247
R458 source.n552 source.n551 12.0247
R459 source.n465 source.n438 12.0247
R460 source.n476 source.n475 12.0247
R461 source.n399 source.n372 12.0247
R462 source.n410 source.n409 12.0247
R463 source.n323 source.n296 12.0247
R464 source.n334 source.n333 12.0247
R465 source.n50 source.n49 12.0247
R466 source.n40 source.n13 12.0247
R467 source.n126 source.n125 12.0247
R468 source.n116 source.n89 12.0247
R469 source.n192 source.n191 12.0247
R470 source.n182 source.n155 12.0247
R471 source.n268 source.n267 12.0247
R472 source.n258 source.n231 12.0247
R473 source.n538 source.n537 11.249
R474 source.n555 source.n508 11.249
R475 source.n462 source.n461 11.249
R476 source.n479 source.n432 11.249
R477 source.n396 source.n395 11.249
R478 source.n413 source.n366 11.249
R479 source.n320 source.n319 11.249
R480 source.n337 source.n290 11.249
R481 source.n53 source.n6 11.249
R482 source.n37 source.n36 11.249
R483 source.n129 source.n82 11.249
R484 source.n113 source.n112 11.249
R485 source.n195 source.n148 11.249
R486 source.n179 source.n178 11.249
R487 source.n271 source.n224 11.249
R488 source.n255 source.n254 11.249
R489 source.n534 source.n516 10.4732
R490 source.n556 source.n506 10.4732
R491 source.n458 source.n440 10.4732
R492 source.n480 source.n430 10.4732
R493 source.n392 source.n374 10.4732
R494 source.n414 source.n364 10.4732
R495 source.n316 source.n298 10.4732
R496 source.n338 source.n288 10.4732
R497 source.n54 source.n4 10.4732
R498 source.n33 source.n15 10.4732
R499 source.n130 source.n80 10.4732
R500 source.n109 source.n91 10.4732
R501 source.n196 source.n146 10.4732
R502 source.n175 source.n157 10.4732
R503 source.n272 source.n222 10.4732
R504 source.n251 source.n233 10.4732
R505 source.n523 source.n522 10.2747
R506 source.n447 source.n446 10.2747
R507 source.n381 source.n380 10.2747
R508 source.n305 source.n304 10.2747
R509 source.n22 source.n21 10.2747
R510 source.n98 source.n97 10.2747
R511 source.n164 source.n163 10.2747
R512 source.n240 source.n239 10.2747
R513 source.n533 source.n518 9.69747
R514 source.n560 source.n559 9.69747
R515 source.n457 source.n442 9.69747
R516 source.n484 source.n483 9.69747
R517 source.n391 source.n376 9.69747
R518 source.n418 source.n417 9.69747
R519 source.n315 source.n300 9.69747
R520 source.n342 source.n341 9.69747
R521 source.n58 source.n57 9.69747
R522 source.n32 source.n17 9.69747
R523 source.n134 source.n133 9.69747
R524 source.n108 source.n93 9.69747
R525 source.n200 source.n199 9.69747
R526 source.n174 source.n159 9.69747
R527 source.n276 source.n275 9.69747
R528 source.n250 source.n235 9.69747
R529 source.n566 source.n565 9.45567
R530 source.n490 source.n489 9.45567
R531 source.n424 source.n423 9.45567
R532 source.n348 source.n347 9.45567
R533 source.n64 source.n63 9.45567
R534 source.n140 source.n139 9.45567
R535 source.n206 source.n205 9.45567
R536 source.n282 source.n281 9.45567
R537 source.n565 source.n564 9.3005
R538 source.n504 source.n503 9.3005
R539 source.n559 source.n558 9.3005
R540 source.n557 source.n556 9.3005
R541 source.n508 source.n507 9.3005
R542 source.n551 source.n550 9.3005
R543 source.n549 source.n548 9.3005
R544 source.n525 source.n524 9.3005
R545 source.n520 source.n519 9.3005
R546 source.n531 source.n530 9.3005
R547 source.n533 source.n532 9.3005
R548 source.n516 source.n515 9.3005
R549 source.n539 source.n538 9.3005
R550 source.n541 source.n540 9.3005
R551 source.n542 source.n511 9.3005
R552 source.n489 source.n488 9.3005
R553 source.n428 source.n427 9.3005
R554 source.n483 source.n482 9.3005
R555 source.n481 source.n480 9.3005
R556 source.n432 source.n431 9.3005
R557 source.n475 source.n474 9.3005
R558 source.n473 source.n472 9.3005
R559 source.n449 source.n448 9.3005
R560 source.n444 source.n443 9.3005
R561 source.n455 source.n454 9.3005
R562 source.n457 source.n456 9.3005
R563 source.n440 source.n439 9.3005
R564 source.n463 source.n462 9.3005
R565 source.n465 source.n464 9.3005
R566 source.n466 source.n435 9.3005
R567 source.n423 source.n422 9.3005
R568 source.n362 source.n361 9.3005
R569 source.n417 source.n416 9.3005
R570 source.n415 source.n414 9.3005
R571 source.n366 source.n365 9.3005
R572 source.n409 source.n408 9.3005
R573 source.n407 source.n406 9.3005
R574 source.n383 source.n382 9.3005
R575 source.n378 source.n377 9.3005
R576 source.n389 source.n388 9.3005
R577 source.n391 source.n390 9.3005
R578 source.n374 source.n373 9.3005
R579 source.n397 source.n396 9.3005
R580 source.n399 source.n398 9.3005
R581 source.n400 source.n369 9.3005
R582 source.n347 source.n346 9.3005
R583 source.n286 source.n285 9.3005
R584 source.n341 source.n340 9.3005
R585 source.n339 source.n338 9.3005
R586 source.n290 source.n289 9.3005
R587 source.n333 source.n332 9.3005
R588 source.n331 source.n330 9.3005
R589 source.n307 source.n306 9.3005
R590 source.n302 source.n301 9.3005
R591 source.n313 source.n312 9.3005
R592 source.n315 source.n314 9.3005
R593 source.n298 source.n297 9.3005
R594 source.n321 source.n320 9.3005
R595 source.n323 source.n322 9.3005
R596 source.n324 source.n293 9.3005
R597 source.n24 source.n23 9.3005
R598 source.n19 source.n18 9.3005
R599 source.n30 source.n29 9.3005
R600 source.n32 source.n31 9.3005
R601 source.n15 source.n14 9.3005
R602 source.n38 source.n37 9.3005
R603 source.n40 source.n39 9.3005
R604 source.n12 source.n9 9.3005
R605 source.n63 source.n62 9.3005
R606 source.n2 source.n1 9.3005
R607 source.n57 source.n56 9.3005
R608 source.n55 source.n54 9.3005
R609 source.n6 source.n5 9.3005
R610 source.n49 source.n48 9.3005
R611 source.n47 source.n46 9.3005
R612 source.n100 source.n99 9.3005
R613 source.n95 source.n94 9.3005
R614 source.n106 source.n105 9.3005
R615 source.n108 source.n107 9.3005
R616 source.n91 source.n90 9.3005
R617 source.n114 source.n113 9.3005
R618 source.n116 source.n115 9.3005
R619 source.n88 source.n85 9.3005
R620 source.n139 source.n138 9.3005
R621 source.n78 source.n77 9.3005
R622 source.n133 source.n132 9.3005
R623 source.n131 source.n130 9.3005
R624 source.n82 source.n81 9.3005
R625 source.n125 source.n124 9.3005
R626 source.n123 source.n122 9.3005
R627 source.n166 source.n165 9.3005
R628 source.n161 source.n160 9.3005
R629 source.n172 source.n171 9.3005
R630 source.n174 source.n173 9.3005
R631 source.n157 source.n156 9.3005
R632 source.n180 source.n179 9.3005
R633 source.n182 source.n181 9.3005
R634 source.n154 source.n151 9.3005
R635 source.n205 source.n204 9.3005
R636 source.n144 source.n143 9.3005
R637 source.n199 source.n198 9.3005
R638 source.n197 source.n196 9.3005
R639 source.n148 source.n147 9.3005
R640 source.n191 source.n190 9.3005
R641 source.n189 source.n188 9.3005
R642 source.n242 source.n241 9.3005
R643 source.n237 source.n236 9.3005
R644 source.n248 source.n247 9.3005
R645 source.n250 source.n249 9.3005
R646 source.n233 source.n232 9.3005
R647 source.n256 source.n255 9.3005
R648 source.n258 source.n257 9.3005
R649 source.n230 source.n227 9.3005
R650 source.n281 source.n280 9.3005
R651 source.n220 source.n219 9.3005
R652 source.n275 source.n274 9.3005
R653 source.n273 source.n272 9.3005
R654 source.n224 source.n223 9.3005
R655 source.n267 source.n266 9.3005
R656 source.n265 source.n264 9.3005
R657 source.n530 source.n529 8.92171
R658 source.n563 source.n504 8.92171
R659 source.n454 source.n453 8.92171
R660 source.n487 source.n428 8.92171
R661 source.n388 source.n387 8.92171
R662 source.n421 source.n362 8.92171
R663 source.n312 source.n311 8.92171
R664 source.n345 source.n286 8.92171
R665 source.n61 source.n2 8.92171
R666 source.n29 source.n28 8.92171
R667 source.n137 source.n78 8.92171
R668 source.n105 source.n104 8.92171
R669 source.n203 source.n144 8.92171
R670 source.n171 source.n170 8.92171
R671 source.n279 source.n220 8.92171
R672 source.n247 source.n246 8.92171
R673 source.n526 source.n520 8.14595
R674 source.n564 source.n502 8.14595
R675 source.n450 source.n444 8.14595
R676 source.n488 source.n426 8.14595
R677 source.n384 source.n378 8.14595
R678 source.n422 source.n360 8.14595
R679 source.n308 source.n302 8.14595
R680 source.n346 source.n284 8.14595
R681 source.n62 source.n0 8.14595
R682 source.n25 source.n19 8.14595
R683 source.n138 source.n76 8.14595
R684 source.n101 source.n95 8.14595
R685 source.n204 source.n142 8.14595
R686 source.n167 source.n161 8.14595
R687 source.n280 source.n218 8.14595
R688 source.n243 source.n237 8.14595
R689 source.n525 source.n522 7.3702
R690 source.n449 source.n446 7.3702
R691 source.n383 source.n380 7.3702
R692 source.n307 source.n304 7.3702
R693 source.n24 source.n21 7.3702
R694 source.n100 source.n97 7.3702
R695 source.n166 source.n163 7.3702
R696 source.n242 source.n239 7.3702
R697 source.n526 source.n525 5.81868
R698 source.n566 source.n502 5.81868
R699 source.n450 source.n449 5.81868
R700 source.n490 source.n426 5.81868
R701 source.n384 source.n383 5.81868
R702 source.n424 source.n360 5.81868
R703 source.n308 source.n307 5.81868
R704 source.n348 source.n284 5.81868
R705 source.n64 source.n0 5.81868
R706 source.n25 source.n24 5.81868
R707 source.n140 source.n76 5.81868
R708 source.n101 source.n100 5.81868
R709 source.n206 source.n142 5.81868
R710 source.n167 source.n166 5.81868
R711 source.n282 source.n218 5.81868
R712 source.n243 source.n242 5.81868
R713 source.n568 source.n567 5.7505
R714 source.n529 source.n520 5.04292
R715 source.n564 source.n563 5.04292
R716 source.n453 source.n444 5.04292
R717 source.n488 source.n487 5.04292
R718 source.n387 source.n378 5.04292
R719 source.n422 source.n421 5.04292
R720 source.n311 source.n302 5.04292
R721 source.n346 source.n345 5.04292
R722 source.n62 source.n61 5.04292
R723 source.n28 source.n19 5.04292
R724 source.n138 source.n137 5.04292
R725 source.n104 source.n95 5.04292
R726 source.n204 source.n203 5.04292
R727 source.n170 source.n161 5.04292
R728 source.n280 source.n279 5.04292
R729 source.n246 source.n237 5.04292
R730 source.n530 source.n518 4.26717
R731 source.n560 source.n504 4.26717
R732 source.n454 source.n442 4.26717
R733 source.n484 source.n428 4.26717
R734 source.n388 source.n376 4.26717
R735 source.n418 source.n362 4.26717
R736 source.n312 source.n300 4.26717
R737 source.n342 source.n286 4.26717
R738 source.n58 source.n2 4.26717
R739 source.n29 source.n17 4.26717
R740 source.n134 source.n78 4.26717
R741 source.n105 source.n93 4.26717
R742 source.n200 source.n144 4.26717
R743 source.n171 source.n159 4.26717
R744 source.n276 source.n220 4.26717
R745 source.n247 source.n235 4.26717
R746 source.n534 source.n533 3.49141
R747 source.n559 source.n506 3.49141
R748 source.n458 source.n457 3.49141
R749 source.n483 source.n430 3.49141
R750 source.n392 source.n391 3.49141
R751 source.n417 source.n364 3.49141
R752 source.n316 source.n315 3.49141
R753 source.n341 source.n288 3.49141
R754 source.n57 source.n4 3.49141
R755 source.n33 source.n32 3.49141
R756 source.n133 source.n80 3.49141
R757 source.n109 source.n108 3.49141
R758 source.n199 source.n146 3.49141
R759 source.n175 source.n174 3.49141
R760 source.n275 source.n222 3.49141
R761 source.n251 source.n250 3.49141
R762 source.n524 source.n523 2.84303
R763 source.n448 source.n447 2.84303
R764 source.n382 source.n381 2.84303
R765 source.n306 source.n305 2.84303
R766 source.n23 source.n22 2.84303
R767 source.n99 source.n98 2.84303
R768 source.n165 source.n164 2.84303
R769 source.n241 source.n240 2.84303
R770 source.n537 source.n516 2.71565
R771 source.n556 source.n555 2.71565
R772 source.n461 source.n440 2.71565
R773 source.n480 source.n479 2.71565
R774 source.n395 source.n374 2.71565
R775 source.n414 source.n413 2.71565
R776 source.n319 source.n298 2.71565
R777 source.n338 source.n337 2.71565
R778 source.n54 source.n53 2.71565
R779 source.n36 source.n15 2.71565
R780 source.n130 source.n129 2.71565
R781 source.n112 source.n91 2.71565
R782 source.n196 source.n195 2.71565
R783 source.n178 source.n157 2.71565
R784 source.n272 source.n271 2.71565
R785 source.n254 source.n233 2.71565
R786 source.n538 source.n514 1.93989
R787 source.n552 source.n508 1.93989
R788 source.n462 source.n438 1.93989
R789 source.n476 source.n432 1.93989
R790 source.n396 source.n372 1.93989
R791 source.n410 source.n366 1.93989
R792 source.n320 source.n296 1.93989
R793 source.n334 source.n290 1.93989
R794 source.n50 source.n6 1.93989
R795 source.n37 source.n13 1.93989
R796 source.n126 source.n82 1.93989
R797 source.n113 source.n89 1.93989
R798 source.n192 source.n148 1.93989
R799 source.n179 source.n155 1.93989
R800 source.n268 source.n224 1.93989
R801 source.n255 source.n231 1.93989
R802 source.n500 source.t26 1.6505
R803 source.n500 source.t28 1.6505
R804 source.n498 source.t22 1.6505
R805 source.n498 source.t40 1.6505
R806 source.n496 source.t31 1.6505
R807 source.n496 source.t37 1.6505
R808 source.n494 source.t38 1.6505
R809 source.n494 source.t27 1.6505
R810 source.n492 source.t20 1.6505
R811 source.n492 source.t21 1.6505
R812 source.n358 source.t18 1.6505
R813 source.n358 source.t7 1.6505
R814 source.n356 source.t12 1.6505
R815 source.n356 source.t10 1.6505
R816 source.n354 source.t47 1.6505
R817 source.n354 source.t19 1.6505
R818 source.n352 source.t44 1.6505
R819 source.n352 source.t5 1.6505
R820 source.n350 source.t16 1.6505
R821 source.n350 source.t13 1.6505
R822 source.n66 source.t17 1.6505
R823 source.n66 source.t2 1.6505
R824 source.n68 source.t4 1.6505
R825 source.n68 source.t14 1.6505
R826 source.n70 source.t46 1.6505
R827 source.n70 source.t0 1.6505
R828 source.n72 source.t45 1.6505
R829 source.n72 source.t1 1.6505
R830 source.n74 source.t3 1.6505
R831 source.n74 source.t8 1.6505
R832 source.n208 source.t43 1.6505
R833 source.n208 source.t32 1.6505
R834 source.n210 source.t39 1.6505
R835 source.n210 source.t23 1.6505
R836 source.n212 source.t41 1.6505
R837 source.n212 source.t36 1.6505
R838 source.n214 source.t25 1.6505
R839 source.n214 source.t33 1.6505
R840 source.n216 source.t30 1.6505
R841 source.n216 source.t35 1.6505
R842 source.n543 source.n541 1.16414
R843 source.n551 source.n510 1.16414
R844 source.n467 source.n465 1.16414
R845 source.n475 source.n434 1.16414
R846 source.n401 source.n399 1.16414
R847 source.n409 source.n368 1.16414
R848 source.n325 source.n323 1.16414
R849 source.n333 source.n292 1.16414
R850 source.n49 source.n8 1.16414
R851 source.n41 source.n40 1.16414
R852 source.n125 source.n84 1.16414
R853 source.n117 source.n116 1.16414
R854 source.n191 source.n150 1.16414
R855 source.n183 source.n182 1.16414
R856 source.n267 source.n226 1.16414
R857 source.n259 source.n258 1.16414
R858 source.n283 source.n217 0.974638
R859 source.n217 source.n215 0.974638
R860 source.n215 source.n213 0.974638
R861 source.n213 source.n211 0.974638
R862 source.n211 source.n209 0.974638
R863 source.n209 source.n207 0.974638
R864 source.n141 source.n75 0.974638
R865 source.n75 source.n73 0.974638
R866 source.n73 source.n71 0.974638
R867 source.n71 source.n69 0.974638
R868 source.n69 source.n67 0.974638
R869 source.n67 source.n65 0.974638
R870 source.n351 source.n349 0.974638
R871 source.n353 source.n351 0.974638
R872 source.n355 source.n353 0.974638
R873 source.n357 source.n355 0.974638
R874 source.n359 source.n357 0.974638
R875 source.n425 source.n359 0.974638
R876 source.n493 source.n491 0.974638
R877 source.n495 source.n493 0.974638
R878 source.n497 source.n495 0.974638
R879 source.n499 source.n497 0.974638
R880 source.n501 source.n499 0.974638
R881 source.n567 source.n501 0.974638
R882 source.n207 source.n141 0.470328
R883 source.n491 source.n425 0.470328
R884 source.n542 source.n512 0.388379
R885 source.n548 source.n547 0.388379
R886 source.n466 source.n436 0.388379
R887 source.n472 source.n471 0.388379
R888 source.n400 source.n370 0.388379
R889 source.n406 source.n405 0.388379
R890 source.n324 source.n294 0.388379
R891 source.n330 source.n329 0.388379
R892 source.n46 source.n45 0.388379
R893 source.n12 source.n10 0.388379
R894 source.n122 source.n121 0.388379
R895 source.n88 source.n86 0.388379
R896 source.n188 source.n187 0.388379
R897 source.n154 source.n152 0.388379
R898 source.n264 source.n263 0.388379
R899 source.n230 source.n228 0.388379
R900 source source.n568 0.188
R901 source.n524 source.n519 0.155672
R902 source.n531 source.n519 0.155672
R903 source.n532 source.n531 0.155672
R904 source.n532 source.n515 0.155672
R905 source.n539 source.n515 0.155672
R906 source.n540 source.n539 0.155672
R907 source.n540 source.n511 0.155672
R908 source.n549 source.n511 0.155672
R909 source.n550 source.n549 0.155672
R910 source.n550 source.n507 0.155672
R911 source.n557 source.n507 0.155672
R912 source.n558 source.n557 0.155672
R913 source.n558 source.n503 0.155672
R914 source.n565 source.n503 0.155672
R915 source.n448 source.n443 0.155672
R916 source.n455 source.n443 0.155672
R917 source.n456 source.n455 0.155672
R918 source.n456 source.n439 0.155672
R919 source.n463 source.n439 0.155672
R920 source.n464 source.n463 0.155672
R921 source.n464 source.n435 0.155672
R922 source.n473 source.n435 0.155672
R923 source.n474 source.n473 0.155672
R924 source.n474 source.n431 0.155672
R925 source.n481 source.n431 0.155672
R926 source.n482 source.n481 0.155672
R927 source.n482 source.n427 0.155672
R928 source.n489 source.n427 0.155672
R929 source.n382 source.n377 0.155672
R930 source.n389 source.n377 0.155672
R931 source.n390 source.n389 0.155672
R932 source.n390 source.n373 0.155672
R933 source.n397 source.n373 0.155672
R934 source.n398 source.n397 0.155672
R935 source.n398 source.n369 0.155672
R936 source.n407 source.n369 0.155672
R937 source.n408 source.n407 0.155672
R938 source.n408 source.n365 0.155672
R939 source.n415 source.n365 0.155672
R940 source.n416 source.n415 0.155672
R941 source.n416 source.n361 0.155672
R942 source.n423 source.n361 0.155672
R943 source.n306 source.n301 0.155672
R944 source.n313 source.n301 0.155672
R945 source.n314 source.n313 0.155672
R946 source.n314 source.n297 0.155672
R947 source.n321 source.n297 0.155672
R948 source.n322 source.n321 0.155672
R949 source.n322 source.n293 0.155672
R950 source.n331 source.n293 0.155672
R951 source.n332 source.n331 0.155672
R952 source.n332 source.n289 0.155672
R953 source.n339 source.n289 0.155672
R954 source.n340 source.n339 0.155672
R955 source.n340 source.n285 0.155672
R956 source.n347 source.n285 0.155672
R957 source.n63 source.n1 0.155672
R958 source.n56 source.n1 0.155672
R959 source.n56 source.n55 0.155672
R960 source.n55 source.n5 0.155672
R961 source.n48 source.n5 0.155672
R962 source.n48 source.n47 0.155672
R963 source.n47 source.n9 0.155672
R964 source.n39 source.n9 0.155672
R965 source.n39 source.n38 0.155672
R966 source.n38 source.n14 0.155672
R967 source.n31 source.n14 0.155672
R968 source.n31 source.n30 0.155672
R969 source.n30 source.n18 0.155672
R970 source.n23 source.n18 0.155672
R971 source.n139 source.n77 0.155672
R972 source.n132 source.n77 0.155672
R973 source.n132 source.n131 0.155672
R974 source.n131 source.n81 0.155672
R975 source.n124 source.n81 0.155672
R976 source.n124 source.n123 0.155672
R977 source.n123 source.n85 0.155672
R978 source.n115 source.n85 0.155672
R979 source.n115 source.n114 0.155672
R980 source.n114 source.n90 0.155672
R981 source.n107 source.n90 0.155672
R982 source.n107 source.n106 0.155672
R983 source.n106 source.n94 0.155672
R984 source.n99 source.n94 0.155672
R985 source.n205 source.n143 0.155672
R986 source.n198 source.n143 0.155672
R987 source.n198 source.n197 0.155672
R988 source.n197 source.n147 0.155672
R989 source.n190 source.n147 0.155672
R990 source.n190 source.n189 0.155672
R991 source.n189 source.n151 0.155672
R992 source.n181 source.n151 0.155672
R993 source.n181 source.n180 0.155672
R994 source.n180 source.n156 0.155672
R995 source.n173 source.n156 0.155672
R996 source.n173 source.n172 0.155672
R997 source.n172 source.n160 0.155672
R998 source.n165 source.n160 0.155672
R999 source.n281 source.n219 0.155672
R1000 source.n274 source.n219 0.155672
R1001 source.n274 source.n273 0.155672
R1002 source.n273 source.n223 0.155672
R1003 source.n266 source.n223 0.155672
R1004 source.n266 source.n265 0.155672
R1005 source.n265 source.n227 0.155672
R1006 source.n257 source.n227 0.155672
R1007 source.n257 source.n256 0.155672
R1008 source.n256 source.n232 0.155672
R1009 source.n249 source.n232 0.155672
R1010 source.n249 source.n248 0.155672
R1011 source.n248 source.n236 0.155672
R1012 source.n241 source.n236 0.155672
R1013 drain_right.n7 drain_right.n5 60.5266
R1014 drain_right.n2 drain_right.n0 60.5266
R1015 drain_right.n13 drain_right.n11 60.5266
R1016 drain_right.n13 drain_right.n12 59.5527
R1017 drain_right.n15 drain_right.n14 59.5527
R1018 drain_right.n17 drain_right.n16 59.5527
R1019 drain_right.n19 drain_right.n18 59.5527
R1020 drain_right.n21 drain_right.n20 59.5527
R1021 drain_right.n7 drain_right.n6 59.5525
R1022 drain_right.n9 drain_right.n8 59.5525
R1023 drain_right.n4 drain_right.n3 59.5525
R1024 drain_right.n2 drain_right.n1 59.5525
R1025 drain_right drain_right.n10 36.0682
R1026 drain_right drain_right.n21 6.62735
R1027 drain_right.n5 drain_right.t19 1.6505
R1028 drain_right.n5 drain_right.t2 1.6505
R1029 drain_right.n6 drain_right.t5 1.6505
R1030 drain_right.n6 drain_right.t22 1.6505
R1031 drain_right.n8 drain_right.t6 1.6505
R1032 drain_right.n8 drain_right.t23 1.6505
R1033 drain_right.n3 drain_right.t1 1.6505
R1034 drain_right.n3 drain_right.t21 1.6505
R1035 drain_right.n1 drain_right.t4 1.6505
R1036 drain_right.n1 drain_right.t20 1.6505
R1037 drain_right.n0 drain_right.t0 1.6505
R1038 drain_right.n0 drain_right.t17 1.6505
R1039 drain_right.n11 drain_right.t15 1.6505
R1040 drain_right.n11 drain_right.t11 1.6505
R1041 drain_right.n12 drain_right.t9 1.6505
R1042 drain_right.n12 drain_right.t16 1.6505
R1043 drain_right.n14 drain_right.t10 1.6505
R1044 drain_right.n14 drain_right.t7 1.6505
R1045 drain_right.n16 drain_right.t3 1.6505
R1046 drain_right.n16 drain_right.t13 1.6505
R1047 drain_right.n18 drain_right.t18 1.6505
R1048 drain_right.n18 drain_right.t8 1.6505
R1049 drain_right.n20 drain_right.t14 1.6505
R1050 drain_right.n20 drain_right.t12 1.6505
R1051 drain_right.n9 drain_right.n7 0.974638
R1052 drain_right.n4 drain_right.n2 0.974638
R1053 drain_right.n21 drain_right.n19 0.974638
R1054 drain_right.n19 drain_right.n17 0.974638
R1055 drain_right.n17 drain_right.n15 0.974638
R1056 drain_right.n15 drain_right.n13 0.974638
R1057 drain_right.n10 drain_right.n9 0.432223
R1058 drain_right.n10 drain_right.n4 0.432223
R1059 plus.n10 plus.t21 432.041
R1060 plus.n46 plus.t18 432.041
R1061 plus.n34 plus.t4 410.604
R1062 plus.n32 plus.t7 410.604
R1063 plus.n31 plus.t8 410.604
R1064 plus.n3 plus.t9 410.604
R1065 plus.n25 plus.t11 410.604
R1066 plus.n5 plus.t13 410.604
R1067 plus.n20 plus.t14 410.604
R1068 plus.n18 plus.t19 410.604
R1069 plus.n8 plus.t15 410.604
R1070 plus.n12 plus.t16 410.604
R1071 plus.n11 plus.t20 410.604
R1072 plus.n70 plus.t23 410.604
R1073 plus.n68 plus.t5 410.604
R1074 plus.n67 plus.t17 410.604
R1075 plus.n39 plus.t3 410.604
R1076 plus.n61 plus.t0 410.604
R1077 plus.n41 plus.t6 410.604
R1078 plus.n56 plus.t22 410.604
R1079 plus.n54 plus.t10 410.604
R1080 plus.n44 plus.t1 410.604
R1081 plus.n48 plus.t12 410.604
R1082 plus.n47 plus.t2 410.604
R1083 plus.n14 plus.n13 161.3
R1084 plus.n15 plus.n8 161.3
R1085 plus.n17 plus.n16 161.3
R1086 plus.n18 plus.n7 161.3
R1087 plus.n19 plus.n6 161.3
R1088 plus.n24 plus.n23 161.3
R1089 plus.n25 plus.n4 161.3
R1090 plus.n27 plus.n26 161.3
R1091 plus.n28 plus.n3 161.3
R1092 plus.n30 plus.n29 161.3
R1093 plus.n33 plus.n0 161.3
R1094 plus.n35 plus.n34 161.3
R1095 plus.n50 plus.n49 161.3
R1096 plus.n51 plus.n44 161.3
R1097 plus.n53 plus.n52 161.3
R1098 plus.n54 plus.n43 161.3
R1099 plus.n55 plus.n42 161.3
R1100 plus.n60 plus.n59 161.3
R1101 plus.n61 plus.n40 161.3
R1102 plus.n63 plus.n62 161.3
R1103 plus.n64 plus.n39 161.3
R1104 plus.n66 plus.n65 161.3
R1105 plus.n69 plus.n36 161.3
R1106 plus.n71 plus.n70 161.3
R1107 plus.n12 plus.n9 80.6037
R1108 plus.n21 plus.n20 80.6037
R1109 plus.n22 plus.n5 80.6037
R1110 plus.n31 plus.n2 80.6037
R1111 plus.n32 plus.n1 80.6037
R1112 plus.n48 plus.n45 80.6037
R1113 plus.n57 plus.n56 80.6037
R1114 plus.n58 plus.n41 80.6037
R1115 plus.n67 plus.n38 80.6037
R1116 plus.n68 plus.n37 80.6037
R1117 plus.n32 plus.n31 48.2005
R1118 plus.n20 plus.n5 48.2005
R1119 plus.n12 plus.n11 48.2005
R1120 plus.n68 plus.n67 48.2005
R1121 plus.n56 plus.n41 48.2005
R1122 plus.n48 plus.n47 48.2005
R1123 plus.n31 plus.n30 44.549
R1124 plus.n13 plus.n12 44.549
R1125 plus.n67 plus.n66 44.549
R1126 plus.n49 plus.n48 44.549
R1127 plus.n24 plus.n5 41.6278
R1128 plus.n20 plus.n19 41.6278
R1129 plus.n60 plus.n41 41.6278
R1130 plus.n56 plus.n55 41.6278
R1131 plus.n33 plus.n32 38.7066
R1132 plus.n69 plus.n68 38.7066
R1133 plus plus.n71 37.0028
R1134 plus.n10 plus.n9 31.6825
R1135 plus.n46 plus.n45 31.6825
R1136 plus.n26 plus.n3 25.5611
R1137 plus.n17 plus.n8 25.5611
R1138 plus.n62 plus.n39 25.5611
R1139 plus.n53 plus.n44 25.5611
R1140 plus.n26 plus.n25 22.6399
R1141 plus.n18 plus.n17 22.6399
R1142 plus.n62 plus.n61 22.6399
R1143 plus.n54 plus.n53 22.6399
R1144 plus.n11 plus.n10 17.2341
R1145 plus.n47 plus.n46 17.2341
R1146 plus plus.n35 12.3035
R1147 plus.n34 plus.n33 9.49444
R1148 plus.n70 plus.n69 9.49444
R1149 plus.n25 plus.n24 6.57323
R1150 plus.n19 plus.n18 6.57323
R1151 plus.n61 plus.n60 6.57323
R1152 plus.n55 plus.n54 6.57323
R1153 plus.n30 plus.n3 3.65202
R1154 plus.n13 plus.n8 3.65202
R1155 plus.n66 plus.n39 3.65202
R1156 plus.n49 plus.n44 3.65202
R1157 plus.n22 plus.n21 0.380177
R1158 plus.n2 plus.n1 0.380177
R1159 plus.n38 plus.n37 0.380177
R1160 plus.n58 plus.n57 0.380177
R1161 plus.n14 plus.n9 0.285035
R1162 plus.n21 plus.n6 0.285035
R1163 plus.n23 plus.n22 0.285035
R1164 plus.n29 plus.n2 0.285035
R1165 plus.n1 plus.n0 0.285035
R1166 plus.n37 plus.n36 0.285035
R1167 plus.n65 plus.n38 0.285035
R1168 plus.n59 plus.n58 0.285035
R1169 plus.n57 plus.n42 0.285035
R1170 plus.n50 plus.n45 0.285035
R1171 plus.n15 plus.n14 0.189894
R1172 plus.n16 plus.n15 0.189894
R1173 plus.n16 plus.n7 0.189894
R1174 plus.n7 plus.n6 0.189894
R1175 plus.n23 plus.n4 0.189894
R1176 plus.n27 plus.n4 0.189894
R1177 plus.n28 plus.n27 0.189894
R1178 plus.n29 plus.n28 0.189894
R1179 plus.n35 plus.n0 0.189894
R1180 plus.n71 plus.n36 0.189894
R1181 plus.n65 plus.n64 0.189894
R1182 plus.n64 plus.n63 0.189894
R1183 plus.n63 plus.n40 0.189894
R1184 plus.n59 plus.n40 0.189894
R1185 plus.n43 plus.n42 0.189894
R1186 plus.n52 plus.n43 0.189894
R1187 plus.n52 plus.n51 0.189894
R1188 plus.n51 plus.n50 0.189894
R1189 drain_left.n13 drain_left.n11 60.5268
R1190 drain_left.n7 drain_left.n5 60.5266
R1191 drain_left.n2 drain_left.n0 60.5266
R1192 drain_left.n19 drain_left.n18 59.5527
R1193 drain_left.n17 drain_left.n16 59.5527
R1194 drain_left.n15 drain_left.n14 59.5527
R1195 drain_left.n13 drain_left.n12 59.5527
R1196 drain_left.n7 drain_left.n6 59.5525
R1197 drain_left.n9 drain_left.n8 59.5525
R1198 drain_left.n4 drain_left.n3 59.5525
R1199 drain_left.n2 drain_left.n1 59.5525
R1200 drain_left.n21 drain_left.n20 59.5525
R1201 drain_left drain_left.n10 36.6214
R1202 drain_left drain_left.n21 6.62735
R1203 drain_left.n5 drain_left.t21 1.6505
R1204 drain_left.n5 drain_left.t5 1.6505
R1205 drain_left.n6 drain_left.t22 1.6505
R1206 drain_left.n6 drain_left.t11 1.6505
R1207 drain_left.n8 drain_left.t1 1.6505
R1208 drain_left.n8 drain_left.t13 1.6505
R1209 drain_left.n3 drain_left.t23 1.6505
R1210 drain_left.n3 drain_left.t17 1.6505
R1211 drain_left.n1 drain_left.t6 1.6505
R1212 drain_left.n1 drain_left.t20 1.6505
R1213 drain_left.n0 drain_left.t0 1.6505
R1214 drain_left.n0 drain_left.t18 1.6505
R1215 drain_left.n20 drain_left.t16 1.6505
R1216 drain_left.n20 drain_left.t19 1.6505
R1217 drain_left.n18 drain_left.t14 1.6505
R1218 drain_left.n18 drain_left.t15 1.6505
R1219 drain_left.n16 drain_left.t10 1.6505
R1220 drain_left.n16 drain_left.t12 1.6505
R1221 drain_left.n14 drain_left.t4 1.6505
R1222 drain_left.n14 drain_left.t9 1.6505
R1223 drain_left.n12 drain_left.t7 1.6505
R1224 drain_left.n12 drain_left.t8 1.6505
R1225 drain_left.n11 drain_left.t2 1.6505
R1226 drain_left.n11 drain_left.t3 1.6505
R1227 drain_left.n9 drain_left.n7 0.974638
R1228 drain_left.n4 drain_left.n2 0.974638
R1229 drain_left.n15 drain_left.n13 0.974638
R1230 drain_left.n17 drain_left.n15 0.974638
R1231 drain_left.n19 drain_left.n17 0.974638
R1232 drain_left.n21 drain_left.n19 0.974638
R1233 drain_left.n10 drain_left.n9 0.432223
R1234 drain_left.n10 drain_left.n4 0.432223
C0 drain_right minus 16.068901f
C1 plus drain_left 16.4364f
C2 plus source 16.4871f
C3 plus drain_right 0.526806f
C4 drain_left source 26.4633f
C5 plus minus 7.70879f
C6 drain_right drain_left 2.02887f
C7 drain_left minus 0.175388f
C8 drain_right source 26.4664f
C9 source minus 16.4731f
C10 drain_right a_n3654_n3288# 8.26849f
C11 drain_left a_n3654_n3288# 8.767981f
C12 source a_n3654_n3288# 9.738027f
C13 minus a_n3654_n3288# 14.874453f
C14 plus a_n3654_n3288# 16.7159f
C15 drain_left.t0 a_n3654_n3288# 0.264495f
C16 drain_left.t18 a_n3654_n3288# 0.264495f
C17 drain_left.n0 a_n3654_n3288# 2.36036f
C18 drain_left.t6 a_n3654_n3288# 0.264495f
C19 drain_left.t20 a_n3654_n3288# 0.264495f
C20 drain_left.n1 a_n3654_n3288# 2.3536f
C21 drain_left.n2 a_n3654_n3288# 0.822843f
C22 drain_left.t23 a_n3654_n3288# 0.264495f
C23 drain_left.t17 a_n3654_n3288# 0.264495f
C24 drain_left.n3 a_n3654_n3288# 2.3536f
C25 drain_left.n4 a_n3654_n3288# 0.361936f
C26 drain_left.t21 a_n3654_n3288# 0.264495f
C27 drain_left.t5 a_n3654_n3288# 0.264495f
C28 drain_left.n5 a_n3654_n3288# 2.36036f
C29 drain_left.t22 a_n3654_n3288# 0.264495f
C30 drain_left.t11 a_n3654_n3288# 0.264495f
C31 drain_left.n6 a_n3654_n3288# 2.3536f
C32 drain_left.n7 a_n3654_n3288# 0.822843f
C33 drain_left.t1 a_n3654_n3288# 0.264495f
C34 drain_left.t13 a_n3654_n3288# 0.264495f
C35 drain_left.n8 a_n3654_n3288# 2.3536f
C36 drain_left.n9 a_n3654_n3288# 0.361936f
C37 drain_left.n10 a_n3654_n3288# 1.9222f
C38 drain_left.t2 a_n3654_n3288# 0.264495f
C39 drain_left.t3 a_n3654_n3288# 0.264495f
C40 drain_left.n11 a_n3654_n3288# 2.36037f
C41 drain_left.t7 a_n3654_n3288# 0.264495f
C42 drain_left.t8 a_n3654_n3288# 0.264495f
C43 drain_left.n12 a_n3654_n3288# 2.3536f
C44 drain_left.n13 a_n3654_n3288# 0.822824f
C45 drain_left.t4 a_n3654_n3288# 0.264495f
C46 drain_left.t9 a_n3654_n3288# 0.264495f
C47 drain_left.n14 a_n3654_n3288# 2.3536f
C48 drain_left.n15 a_n3654_n3288# 0.409178f
C49 drain_left.t10 a_n3654_n3288# 0.264495f
C50 drain_left.t12 a_n3654_n3288# 0.264495f
C51 drain_left.n16 a_n3654_n3288# 2.3536f
C52 drain_left.n17 a_n3654_n3288# 0.409178f
C53 drain_left.t14 a_n3654_n3288# 0.264495f
C54 drain_left.t15 a_n3654_n3288# 0.264495f
C55 drain_left.n18 a_n3654_n3288# 2.3536f
C56 drain_left.n19 a_n3654_n3288# 0.409178f
C57 drain_left.t16 a_n3654_n3288# 0.264495f
C58 drain_left.t19 a_n3654_n3288# 0.264495f
C59 drain_left.n20 a_n3654_n3288# 2.3536f
C60 drain_left.n21 a_n3654_n3288# 0.659295f
C61 plus.n0 a_n3654_n3288# 0.050151f
C62 plus.t4 a_n3654_n3288# 1.02883f
C63 plus.t7 a_n3654_n3288# 1.02883f
C64 plus.n1 a_n3654_n3288# 0.0626f
C65 plus.t8 a_n3654_n3288# 1.02883f
C66 plus.n2 a_n3654_n3288# 0.0626f
C67 plus.t9 a_n3654_n3288# 1.02883f
C68 plus.n3 a_n3654_n3288# 0.406881f
C69 plus.n4 a_n3654_n3288# 0.037584f
C70 plus.t11 a_n3654_n3288# 1.02883f
C71 plus.t13 a_n3654_n3288# 1.02883f
C72 plus.n5 a_n3654_n3288# 0.417379f
C73 plus.n6 a_n3654_n3288# 0.050151f
C74 plus.t14 a_n3654_n3288# 1.02883f
C75 plus.t19 a_n3654_n3288# 1.02883f
C76 plus.n7 a_n3654_n3288# 0.037584f
C77 plus.t15 a_n3654_n3288# 1.02883f
C78 plus.n8 a_n3654_n3288# 0.406881f
C79 plus.n9 a_n3654_n3288# 0.216016f
C80 plus.t16 a_n3654_n3288# 1.02883f
C81 plus.t20 a_n3654_n3288# 1.02883f
C82 plus.t21 a_n3654_n3288# 1.04917f
C83 plus.n10 a_n3654_n3288# 0.393276f
C84 plus.n11 a_n3654_n3288# 0.417823f
C85 plus.n12 a_n3654_n3288# 0.417842f
C86 plus.n13 a_n3654_n3288# 0.008528f
C87 plus.n14 a_n3654_n3288# 0.050151f
C88 plus.n15 a_n3654_n3288# 0.037584f
C89 plus.n16 a_n3654_n3288# 0.037584f
C90 plus.n17 a_n3654_n3288# 0.008528f
C91 plus.n18 a_n3654_n3288# 0.406881f
C92 plus.n19 a_n3654_n3288# 0.008528f
C93 plus.n20 a_n3654_n3288# 0.417379f
C94 plus.n21 a_n3654_n3288# 0.0626f
C95 plus.n22 a_n3654_n3288# 0.0626f
C96 plus.n23 a_n3654_n3288# 0.050151f
C97 plus.n24 a_n3654_n3288# 0.008528f
C98 plus.n25 a_n3654_n3288# 0.406881f
C99 plus.n26 a_n3654_n3288# 0.008528f
C100 plus.n27 a_n3654_n3288# 0.037584f
C101 plus.n28 a_n3654_n3288# 0.037584f
C102 plus.n29 a_n3654_n3288# 0.050151f
C103 plus.n30 a_n3654_n3288# 0.008528f
C104 plus.n31 a_n3654_n3288# 0.417842f
C105 plus.n32 a_n3654_n3288# 0.416915f
C106 plus.n33 a_n3654_n3288# 0.008528f
C107 plus.n34 a_n3654_n3288# 0.403752f
C108 plus.n35 a_n3654_n3288# 0.434784f
C109 plus.n36 a_n3654_n3288# 0.050151f
C110 plus.t23 a_n3654_n3288# 1.02883f
C111 plus.n37 a_n3654_n3288# 0.0626f
C112 plus.t5 a_n3654_n3288# 1.02883f
C113 plus.n38 a_n3654_n3288# 0.0626f
C114 plus.t17 a_n3654_n3288# 1.02883f
C115 plus.t3 a_n3654_n3288# 1.02883f
C116 plus.n39 a_n3654_n3288# 0.406881f
C117 plus.n40 a_n3654_n3288# 0.037584f
C118 plus.t0 a_n3654_n3288# 1.02883f
C119 plus.t6 a_n3654_n3288# 1.02883f
C120 plus.n41 a_n3654_n3288# 0.417379f
C121 plus.n42 a_n3654_n3288# 0.050151f
C122 plus.t22 a_n3654_n3288# 1.02883f
C123 plus.n43 a_n3654_n3288# 0.037584f
C124 plus.t10 a_n3654_n3288# 1.02883f
C125 plus.t1 a_n3654_n3288# 1.02883f
C126 plus.n44 a_n3654_n3288# 0.406881f
C127 plus.n45 a_n3654_n3288# 0.216016f
C128 plus.t12 a_n3654_n3288# 1.02883f
C129 plus.t18 a_n3654_n3288# 1.04917f
C130 plus.n46 a_n3654_n3288# 0.393276f
C131 plus.t2 a_n3654_n3288# 1.02883f
C132 plus.n47 a_n3654_n3288# 0.417823f
C133 plus.n48 a_n3654_n3288# 0.417842f
C134 plus.n49 a_n3654_n3288# 0.008528f
C135 plus.n50 a_n3654_n3288# 0.050151f
C136 plus.n51 a_n3654_n3288# 0.037584f
C137 plus.n52 a_n3654_n3288# 0.037584f
C138 plus.n53 a_n3654_n3288# 0.008528f
C139 plus.n54 a_n3654_n3288# 0.406881f
C140 plus.n55 a_n3654_n3288# 0.008528f
C141 plus.n56 a_n3654_n3288# 0.417379f
C142 plus.n57 a_n3654_n3288# 0.0626f
C143 plus.n58 a_n3654_n3288# 0.0626f
C144 plus.n59 a_n3654_n3288# 0.050151f
C145 plus.n60 a_n3654_n3288# 0.008528f
C146 plus.n61 a_n3654_n3288# 0.406881f
C147 plus.n62 a_n3654_n3288# 0.008528f
C148 plus.n63 a_n3654_n3288# 0.037584f
C149 plus.n64 a_n3654_n3288# 0.037584f
C150 plus.n65 a_n3654_n3288# 0.050151f
C151 plus.n66 a_n3654_n3288# 0.008528f
C152 plus.n67 a_n3654_n3288# 0.417842f
C153 plus.n68 a_n3654_n3288# 0.416915f
C154 plus.n69 a_n3654_n3288# 0.008528f
C155 plus.n70 a_n3654_n3288# 0.403752f
C156 plus.n71 a_n3654_n3288# 1.49422f
C157 drain_right.t0 a_n3654_n3288# 0.263368f
C158 drain_right.t17 a_n3654_n3288# 0.263368f
C159 drain_right.n0 a_n3654_n3288# 2.3503f
C160 drain_right.t4 a_n3654_n3288# 0.263368f
C161 drain_right.t20 a_n3654_n3288# 0.263368f
C162 drain_right.n1 a_n3654_n3288# 2.34356f
C163 drain_right.n2 a_n3654_n3288# 0.819336f
C164 drain_right.t1 a_n3654_n3288# 0.263368f
C165 drain_right.t21 a_n3654_n3288# 0.263368f
C166 drain_right.n3 a_n3654_n3288# 2.34356f
C167 drain_right.n4 a_n3654_n3288# 0.360393f
C168 drain_right.t19 a_n3654_n3288# 0.263368f
C169 drain_right.t2 a_n3654_n3288# 0.263368f
C170 drain_right.n5 a_n3654_n3288# 2.3503f
C171 drain_right.t5 a_n3654_n3288# 0.263368f
C172 drain_right.t22 a_n3654_n3288# 0.263368f
C173 drain_right.n6 a_n3654_n3288# 2.34356f
C174 drain_right.n7 a_n3654_n3288# 0.819336f
C175 drain_right.t6 a_n3654_n3288# 0.263368f
C176 drain_right.t23 a_n3654_n3288# 0.263368f
C177 drain_right.n8 a_n3654_n3288# 2.34356f
C178 drain_right.n9 a_n3654_n3288# 0.360393f
C179 drain_right.n10 a_n3654_n3288# 1.85796f
C180 drain_right.t15 a_n3654_n3288# 0.263368f
C181 drain_right.t11 a_n3654_n3288# 0.263368f
C182 drain_right.n11 a_n3654_n3288# 2.3503f
C183 drain_right.t9 a_n3654_n3288# 0.263368f
C184 drain_right.t16 a_n3654_n3288# 0.263368f
C185 drain_right.n12 a_n3654_n3288# 2.34357f
C186 drain_right.n13 a_n3654_n3288# 0.819326f
C187 drain_right.t10 a_n3654_n3288# 0.263368f
C188 drain_right.t7 a_n3654_n3288# 0.263368f
C189 drain_right.n14 a_n3654_n3288# 2.34357f
C190 drain_right.n15 a_n3654_n3288# 0.407434f
C191 drain_right.t3 a_n3654_n3288# 0.263368f
C192 drain_right.t13 a_n3654_n3288# 0.263368f
C193 drain_right.n16 a_n3654_n3288# 2.34357f
C194 drain_right.n17 a_n3654_n3288# 0.407434f
C195 drain_right.t18 a_n3654_n3288# 0.263368f
C196 drain_right.t8 a_n3654_n3288# 0.263368f
C197 drain_right.n18 a_n3654_n3288# 2.34357f
C198 drain_right.n19 a_n3654_n3288# 0.407434f
C199 drain_right.t14 a_n3654_n3288# 0.263368f
C200 drain_right.t12 a_n3654_n3288# 0.263368f
C201 drain_right.n20 a_n3654_n3288# 2.34357f
C202 drain_right.n21 a_n3654_n3288# 0.656475f
C203 source.n0 a_n3654_n3288# 0.032323f
C204 source.n1 a_n3654_n3288# 0.024402f
C205 source.n2 a_n3654_n3288# 0.013112f
C206 source.n3 a_n3654_n3288# 0.030993f
C207 source.n4 a_n3654_n3288# 0.013884f
C208 source.n5 a_n3654_n3288# 0.024402f
C209 source.n6 a_n3654_n3288# 0.013112f
C210 source.n7 a_n3654_n3288# 0.030993f
C211 source.n8 a_n3654_n3288# 0.013884f
C212 source.n9 a_n3654_n3288# 0.024402f
C213 source.n10 a_n3654_n3288# 0.013498f
C214 source.n11 a_n3654_n3288# 0.030993f
C215 source.n12 a_n3654_n3288# 0.013112f
C216 source.n13 a_n3654_n3288# 0.013884f
C217 source.n14 a_n3654_n3288# 0.024402f
C218 source.n15 a_n3654_n3288# 0.013112f
C219 source.n16 a_n3654_n3288# 0.030993f
C220 source.n17 a_n3654_n3288# 0.013884f
C221 source.n18 a_n3654_n3288# 0.024402f
C222 source.n19 a_n3654_n3288# 0.013112f
C223 source.n20 a_n3654_n3288# 0.023245f
C224 source.n21 a_n3654_n3288# 0.02191f
C225 source.t15 a_n3654_n3288# 0.052345f
C226 source.n22 a_n3654_n3288# 0.175934f
C227 source.n23 a_n3654_n3288# 1.23103f
C228 source.n24 a_n3654_n3288# 0.013112f
C229 source.n25 a_n3654_n3288# 0.013884f
C230 source.n26 a_n3654_n3288# 0.030993f
C231 source.n27 a_n3654_n3288# 0.030993f
C232 source.n28 a_n3654_n3288# 0.013884f
C233 source.n29 a_n3654_n3288# 0.013112f
C234 source.n30 a_n3654_n3288# 0.024402f
C235 source.n31 a_n3654_n3288# 0.024402f
C236 source.n32 a_n3654_n3288# 0.013112f
C237 source.n33 a_n3654_n3288# 0.013884f
C238 source.n34 a_n3654_n3288# 0.030993f
C239 source.n35 a_n3654_n3288# 0.030993f
C240 source.n36 a_n3654_n3288# 0.013884f
C241 source.n37 a_n3654_n3288# 0.013112f
C242 source.n38 a_n3654_n3288# 0.024402f
C243 source.n39 a_n3654_n3288# 0.024402f
C244 source.n40 a_n3654_n3288# 0.013112f
C245 source.n41 a_n3654_n3288# 0.013884f
C246 source.n42 a_n3654_n3288# 0.030993f
C247 source.n43 a_n3654_n3288# 0.030993f
C248 source.n44 a_n3654_n3288# 0.030993f
C249 source.n45 a_n3654_n3288# 0.013498f
C250 source.n46 a_n3654_n3288# 0.013112f
C251 source.n47 a_n3654_n3288# 0.024402f
C252 source.n48 a_n3654_n3288# 0.024402f
C253 source.n49 a_n3654_n3288# 0.013112f
C254 source.n50 a_n3654_n3288# 0.013884f
C255 source.n51 a_n3654_n3288# 0.030993f
C256 source.n52 a_n3654_n3288# 0.030993f
C257 source.n53 a_n3654_n3288# 0.013884f
C258 source.n54 a_n3654_n3288# 0.013112f
C259 source.n55 a_n3654_n3288# 0.024402f
C260 source.n56 a_n3654_n3288# 0.024402f
C261 source.n57 a_n3654_n3288# 0.013112f
C262 source.n58 a_n3654_n3288# 0.013884f
C263 source.n59 a_n3654_n3288# 0.030993f
C264 source.n60 a_n3654_n3288# 0.063601f
C265 source.n61 a_n3654_n3288# 0.013884f
C266 source.n62 a_n3654_n3288# 0.013112f
C267 source.n63 a_n3654_n3288# 0.052403f
C268 source.n64 a_n3654_n3288# 0.035101f
C269 source.n65 a_n3654_n3288# 1.03759f
C270 source.t17 a_n3654_n3288# 0.231396f
C271 source.t2 a_n3654_n3288# 0.231396f
C272 source.n66 a_n3654_n3288# 1.98122f
C273 source.n67 a_n3654_n3288# 0.402665f
C274 source.t4 a_n3654_n3288# 0.231396f
C275 source.t14 a_n3654_n3288# 0.231396f
C276 source.n68 a_n3654_n3288# 1.98122f
C277 source.n69 a_n3654_n3288# 0.402665f
C278 source.t46 a_n3654_n3288# 0.231396f
C279 source.t0 a_n3654_n3288# 0.231396f
C280 source.n70 a_n3654_n3288# 1.98122f
C281 source.n71 a_n3654_n3288# 0.402665f
C282 source.t45 a_n3654_n3288# 0.231396f
C283 source.t1 a_n3654_n3288# 0.231396f
C284 source.n72 a_n3654_n3288# 1.98122f
C285 source.n73 a_n3654_n3288# 0.402665f
C286 source.t3 a_n3654_n3288# 0.231396f
C287 source.t8 a_n3654_n3288# 0.231396f
C288 source.n74 a_n3654_n3288# 1.98122f
C289 source.n75 a_n3654_n3288# 0.402665f
C290 source.n76 a_n3654_n3288# 0.032323f
C291 source.n77 a_n3654_n3288# 0.024402f
C292 source.n78 a_n3654_n3288# 0.013112f
C293 source.n79 a_n3654_n3288# 0.030993f
C294 source.n80 a_n3654_n3288# 0.013884f
C295 source.n81 a_n3654_n3288# 0.024402f
C296 source.n82 a_n3654_n3288# 0.013112f
C297 source.n83 a_n3654_n3288# 0.030993f
C298 source.n84 a_n3654_n3288# 0.013884f
C299 source.n85 a_n3654_n3288# 0.024402f
C300 source.n86 a_n3654_n3288# 0.013498f
C301 source.n87 a_n3654_n3288# 0.030993f
C302 source.n88 a_n3654_n3288# 0.013112f
C303 source.n89 a_n3654_n3288# 0.013884f
C304 source.n90 a_n3654_n3288# 0.024402f
C305 source.n91 a_n3654_n3288# 0.013112f
C306 source.n92 a_n3654_n3288# 0.030993f
C307 source.n93 a_n3654_n3288# 0.013884f
C308 source.n94 a_n3654_n3288# 0.024402f
C309 source.n95 a_n3654_n3288# 0.013112f
C310 source.n96 a_n3654_n3288# 0.023245f
C311 source.n97 a_n3654_n3288# 0.02191f
C312 source.t9 a_n3654_n3288# 0.052345f
C313 source.n98 a_n3654_n3288# 0.175934f
C314 source.n99 a_n3654_n3288# 1.23103f
C315 source.n100 a_n3654_n3288# 0.013112f
C316 source.n101 a_n3654_n3288# 0.013884f
C317 source.n102 a_n3654_n3288# 0.030993f
C318 source.n103 a_n3654_n3288# 0.030993f
C319 source.n104 a_n3654_n3288# 0.013884f
C320 source.n105 a_n3654_n3288# 0.013112f
C321 source.n106 a_n3654_n3288# 0.024402f
C322 source.n107 a_n3654_n3288# 0.024402f
C323 source.n108 a_n3654_n3288# 0.013112f
C324 source.n109 a_n3654_n3288# 0.013884f
C325 source.n110 a_n3654_n3288# 0.030993f
C326 source.n111 a_n3654_n3288# 0.030993f
C327 source.n112 a_n3654_n3288# 0.013884f
C328 source.n113 a_n3654_n3288# 0.013112f
C329 source.n114 a_n3654_n3288# 0.024402f
C330 source.n115 a_n3654_n3288# 0.024402f
C331 source.n116 a_n3654_n3288# 0.013112f
C332 source.n117 a_n3654_n3288# 0.013884f
C333 source.n118 a_n3654_n3288# 0.030993f
C334 source.n119 a_n3654_n3288# 0.030993f
C335 source.n120 a_n3654_n3288# 0.030993f
C336 source.n121 a_n3654_n3288# 0.013498f
C337 source.n122 a_n3654_n3288# 0.013112f
C338 source.n123 a_n3654_n3288# 0.024402f
C339 source.n124 a_n3654_n3288# 0.024402f
C340 source.n125 a_n3654_n3288# 0.013112f
C341 source.n126 a_n3654_n3288# 0.013884f
C342 source.n127 a_n3654_n3288# 0.030993f
C343 source.n128 a_n3654_n3288# 0.030993f
C344 source.n129 a_n3654_n3288# 0.013884f
C345 source.n130 a_n3654_n3288# 0.013112f
C346 source.n131 a_n3654_n3288# 0.024402f
C347 source.n132 a_n3654_n3288# 0.024402f
C348 source.n133 a_n3654_n3288# 0.013112f
C349 source.n134 a_n3654_n3288# 0.013884f
C350 source.n135 a_n3654_n3288# 0.030993f
C351 source.n136 a_n3654_n3288# 0.063601f
C352 source.n137 a_n3654_n3288# 0.013884f
C353 source.n138 a_n3654_n3288# 0.013112f
C354 source.n139 a_n3654_n3288# 0.052403f
C355 source.n140 a_n3654_n3288# 0.035101f
C356 source.n141 a_n3654_n3288# 0.132123f
C357 source.n142 a_n3654_n3288# 0.032323f
C358 source.n143 a_n3654_n3288# 0.024402f
C359 source.n144 a_n3654_n3288# 0.013112f
C360 source.n145 a_n3654_n3288# 0.030993f
C361 source.n146 a_n3654_n3288# 0.013884f
C362 source.n147 a_n3654_n3288# 0.024402f
C363 source.n148 a_n3654_n3288# 0.013112f
C364 source.n149 a_n3654_n3288# 0.030993f
C365 source.n150 a_n3654_n3288# 0.013884f
C366 source.n151 a_n3654_n3288# 0.024402f
C367 source.n152 a_n3654_n3288# 0.013498f
C368 source.n153 a_n3654_n3288# 0.030993f
C369 source.n154 a_n3654_n3288# 0.013112f
C370 source.n155 a_n3654_n3288# 0.013884f
C371 source.n156 a_n3654_n3288# 0.024402f
C372 source.n157 a_n3654_n3288# 0.013112f
C373 source.n158 a_n3654_n3288# 0.030993f
C374 source.n159 a_n3654_n3288# 0.013884f
C375 source.n160 a_n3654_n3288# 0.024402f
C376 source.n161 a_n3654_n3288# 0.013112f
C377 source.n162 a_n3654_n3288# 0.023245f
C378 source.n163 a_n3654_n3288# 0.02191f
C379 source.t29 a_n3654_n3288# 0.052345f
C380 source.n164 a_n3654_n3288# 0.175934f
C381 source.n165 a_n3654_n3288# 1.23103f
C382 source.n166 a_n3654_n3288# 0.013112f
C383 source.n167 a_n3654_n3288# 0.013884f
C384 source.n168 a_n3654_n3288# 0.030993f
C385 source.n169 a_n3654_n3288# 0.030993f
C386 source.n170 a_n3654_n3288# 0.013884f
C387 source.n171 a_n3654_n3288# 0.013112f
C388 source.n172 a_n3654_n3288# 0.024402f
C389 source.n173 a_n3654_n3288# 0.024402f
C390 source.n174 a_n3654_n3288# 0.013112f
C391 source.n175 a_n3654_n3288# 0.013884f
C392 source.n176 a_n3654_n3288# 0.030993f
C393 source.n177 a_n3654_n3288# 0.030993f
C394 source.n178 a_n3654_n3288# 0.013884f
C395 source.n179 a_n3654_n3288# 0.013112f
C396 source.n180 a_n3654_n3288# 0.024402f
C397 source.n181 a_n3654_n3288# 0.024402f
C398 source.n182 a_n3654_n3288# 0.013112f
C399 source.n183 a_n3654_n3288# 0.013884f
C400 source.n184 a_n3654_n3288# 0.030993f
C401 source.n185 a_n3654_n3288# 0.030993f
C402 source.n186 a_n3654_n3288# 0.030993f
C403 source.n187 a_n3654_n3288# 0.013498f
C404 source.n188 a_n3654_n3288# 0.013112f
C405 source.n189 a_n3654_n3288# 0.024402f
C406 source.n190 a_n3654_n3288# 0.024402f
C407 source.n191 a_n3654_n3288# 0.013112f
C408 source.n192 a_n3654_n3288# 0.013884f
C409 source.n193 a_n3654_n3288# 0.030993f
C410 source.n194 a_n3654_n3288# 0.030993f
C411 source.n195 a_n3654_n3288# 0.013884f
C412 source.n196 a_n3654_n3288# 0.013112f
C413 source.n197 a_n3654_n3288# 0.024402f
C414 source.n198 a_n3654_n3288# 0.024402f
C415 source.n199 a_n3654_n3288# 0.013112f
C416 source.n200 a_n3654_n3288# 0.013884f
C417 source.n201 a_n3654_n3288# 0.030993f
C418 source.n202 a_n3654_n3288# 0.063601f
C419 source.n203 a_n3654_n3288# 0.013884f
C420 source.n204 a_n3654_n3288# 0.013112f
C421 source.n205 a_n3654_n3288# 0.052403f
C422 source.n206 a_n3654_n3288# 0.035101f
C423 source.n207 a_n3654_n3288# 0.132123f
C424 source.t43 a_n3654_n3288# 0.231396f
C425 source.t32 a_n3654_n3288# 0.231396f
C426 source.n208 a_n3654_n3288# 1.98122f
C427 source.n209 a_n3654_n3288# 0.402665f
C428 source.t39 a_n3654_n3288# 0.231396f
C429 source.t23 a_n3654_n3288# 0.231396f
C430 source.n210 a_n3654_n3288# 1.98122f
C431 source.n211 a_n3654_n3288# 0.402665f
C432 source.t41 a_n3654_n3288# 0.231396f
C433 source.t36 a_n3654_n3288# 0.231396f
C434 source.n212 a_n3654_n3288# 1.98122f
C435 source.n213 a_n3654_n3288# 0.402665f
C436 source.t25 a_n3654_n3288# 0.231396f
C437 source.t33 a_n3654_n3288# 0.231396f
C438 source.n214 a_n3654_n3288# 1.98122f
C439 source.n215 a_n3654_n3288# 0.402665f
C440 source.t30 a_n3654_n3288# 0.231396f
C441 source.t35 a_n3654_n3288# 0.231396f
C442 source.n216 a_n3654_n3288# 1.98122f
C443 source.n217 a_n3654_n3288# 0.402665f
C444 source.n218 a_n3654_n3288# 0.032323f
C445 source.n219 a_n3654_n3288# 0.024402f
C446 source.n220 a_n3654_n3288# 0.013112f
C447 source.n221 a_n3654_n3288# 0.030993f
C448 source.n222 a_n3654_n3288# 0.013884f
C449 source.n223 a_n3654_n3288# 0.024402f
C450 source.n224 a_n3654_n3288# 0.013112f
C451 source.n225 a_n3654_n3288# 0.030993f
C452 source.n226 a_n3654_n3288# 0.013884f
C453 source.n227 a_n3654_n3288# 0.024402f
C454 source.n228 a_n3654_n3288# 0.013498f
C455 source.n229 a_n3654_n3288# 0.030993f
C456 source.n230 a_n3654_n3288# 0.013112f
C457 source.n231 a_n3654_n3288# 0.013884f
C458 source.n232 a_n3654_n3288# 0.024402f
C459 source.n233 a_n3654_n3288# 0.013112f
C460 source.n234 a_n3654_n3288# 0.030993f
C461 source.n235 a_n3654_n3288# 0.013884f
C462 source.n236 a_n3654_n3288# 0.024402f
C463 source.n237 a_n3654_n3288# 0.013112f
C464 source.n238 a_n3654_n3288# 0.023245f
C465 source.n239 a_n3654_n3288# 0.02191f
C466 source.t42 a_n3654_n3288# 0.052345f
C467 source.n240 a_n3654_n3288# 0.175934f
C468 source.n241 a_n3654_n3288# 1.23103f
C469 source.n242 a_n3654_n3288# 0.013112f
C470 source.n243 a_n3654_n3288# 0.013884f
C471 source.n244 a_n3654_n3288# 0.030993f
C472 source.n245 a_n3654_n3288# 0.030993f
C473 source.n246 a_n3654_n3288# 0.013884f
C474 source.n247 a_n3654_n3288# 0.013112f
C475 source.n248 a_n3654_n3288# 0.024402f
C476 source.n249 a_n3654_n3288# 0.024402f
C477 source.n250 a_n3654_n3288# 0.013112f
C478 source.n251 a_n3654_n3288# 0.013884f
C479 source.n252 a_n3654_n3288# 0.030993f
C480 source.n253 a_n3654_n3288# 0.030993f
C481 source.n254 a_n3654_n3288# 0.013884f
C482 source.n255 a_n3654_n3288# 0.013112f
C483 source.n256 a_n3654_n3288# 0.024402f
C484 source.n257 a_n3654_n3288# 0.024402f
C485 source.n258 a_n3654_n3288# 0.013112f
C486 source.n259 a_n3654_n3288# 0.013884f
C487 source.n260 a_n3654_n3288# 0.030993f
C488 source.n261 a_n3654_n3288# 0.030993f
C489 source.n262 a_n3654_n3288# 0.030993f
C490 source.n263 a_n3654_n3288# 0.013498f
C491 source.n264 a_n3654_n3288# 0.013112f
C492 source.n265 a_n3654_n3288# 0.024402f
C493 source.n266 a_n3654_n3288# 0.024402f
C494 source.n267 a_n3654_n3288# 0.013112f
C495 source.n268 a_n3654_n3288# 0.013884f
C496 source.n269 a_n3654_n3288# 0.030993f
C497 source.n270 a_n3654_n3288# 0.030993f
C498 source.n271 a_n3654_n3288# 0.013884f
C499 source.n272 a_n3654_n3288# 0.013112f
C500 source.n273 a_n3654_n3288# 0.024402f
C501 source.n274 a_n3654_n3288# 0.024402f
C502 source.n275 a_n3654_n3288# 0.013112f
C503 source.n276 a_n3654_n3288# 0.013884f
C504 source.n277 a_n3654_n3288# 0.030993f
C505 source.n278 a_n3654_n3288# 0.063601f
C506 source.n279 a_n3654_n3288# 0.013884f
C507 source.n280 a_n3654_n3288# 0.013112f
C508 source.n281 a_n3654_n3288# 0.052403f
C509 source.n282 a_n3654_n3288# 0.035101f
C510 source.n283 a_n3654_n3288# 1.43353f
C511 source.n284 a_n3654_n3288# 0.032323f
C512 source.n285 a_n3654_n3288# 0.024402f
C513 source.n286 a_n3654_n3288# 0.013112f
C514 source.n287 a_n3654_n3288# 0.030993f
C515 source.n288 a_n3654_n3288# 0.013884f
C516 source.n289 a_n3654_n3288# 0.024402f
C517 source.n290 a_n3654_n3288# 0.013112f
C518 source.n291 a_n3654_n3288# 0.030993f
C519 source.n292 a_n3654_n3288# 0.013884f
C520 source.n293 a_n3654_n3288# 0.024402f
C521 source.n294 a_n3654_n3288# 0.013498f
C522 source.n295 a_n3654_n3288# 0.030993f
C523 source.n296 a_n3654_n3288# 0.013884f
C524 source.n297 a_n3654_n3288# 0.024402f
C525 source.n298 a_n3654_n3288# 0.013112f
C526 source.n299 a_n3654_n3288# 0.030993f
C527 source.n300 a_n3654_n3288# 0.013884f
C528 source.n301 a_n3654_n3288# 0.024402f
C529 source.n302 a_n3654_n3288# 0.013112f
C530 source.n303 a_n3654_n3288# 0.023245f
C531 source.n304 a_n3654_n3288# 0.02191f
C532 source.t11 a_n3654_n3288# 0.052345f
C533 source.n305 a_n3654_n3288# 0.175934f
C534 source.n306 a_n3654_n3288# 1.23103f
C535 source.n307 a_n3654_n3288# 0.013112f
C536 source.n308 a_n3654_n3288# 0.013884f
C537 source.n309 a_n3654_n3288# 0.030993f
C538 source.n310 a_n3654_n3288# 0.030993f
C539 source.n311 a_n3654_n3288# 0.013884f
C540 source.n312 a_n3654_n3288# 0.013112f
C541 source.n313 a_n3654_n3288# 0.024402f
C542 source.n314 a_n3654_n3288# 0.024402f
C543 source.n315 a_n3654_n3288# 0.013112f
C544 source.n316 a_n3654_n3288# 0.013884f
C545 source.n317 a_n3654_n3288# 0.030993f
C546 source.n318 a_n3654_n3288# 0.030993f
C547 source.n319 a_n3654_n3288# 0.013884f
C548 source.n320 a_n3654_n3288# 0.013112f
C549 source.n321 a_n3654_n3288# 0.024402f
C550 source.n322 a_n3654_n3288# 0.024402f
C551 source.n323 a_n3654_n3288# 0.013112f
C552 source.n324 a_n3654_n3288# 0.013112f
C553 source.n325 a_n3654_n3288# 0.013884f
C554 source.n326 a_n3654_n3288# 0.030993f
C555 source.n327 a_n3654_n3288# 0.030993f
C556 source.n328 a_n3654_n3288# 0.030993f
C557 source.n329 a_n3654_n3288# 0.013498f
C558 source.n330 a_n3654_n3288# 0.013112f
C559 source.n331 a_n3654_n3288# 0.024402f
C560 source.n332 a_n3654_n3288# 0.024402f
C561 source.n333 a_n3654_n3288# 0.013112f
C562 source.n334 a_n3654_n3288# 0.013884f
C563 source.n335 a_n3654_n3288# 0.030993f
C564 source.n336 a_n3654_n3288# 0.030993f
C565 source.n337 a_n3654_n3288# 0.013884f
C566 source.n338 a_n3654_n3288# 0.013112f
C567 source.n339 a_n3654_n3288# 0.024402f
C568 source.n340 a_n3654_n3288# 0.024402f
C569 source.n341 a_n3654_n3288# 0.013112f
C570 source.n342 a_n3654_n3288# 0.013884f
C571 source.n343 a_n3654_n3288# 0.030993f
C572 source.n344 a_n3654_n3288# 0.063601f
C573 source.n345 a_n3654_n3288# 0.013884f
C574 source.n346 a_n3654_n3288# 0.013112f
C575 source.n347 a_n3654_n3288# 0.052403f
C576 source.n348 a_n3654_n3288# 0.035101f
C577 source.n349 a_n3654_n3288# 1.43353f
C578 source.t16 a_n3654_n3288# 0.231396f
C579 source.t13 a_n3654_n3288# 0.231396f
C580 source.n350 a_n3654_n3288# 1.9812f
C581 source.n351 a_n3654_n3288# 0.402677f
C582 source.t44 a_n3654_n3288# 0.231396f
C583 source.t5 a_n3654_n3288# 0.231396f
C584 source.n352 a_n3654_n3288# 1.9812f
C585 source.n353 a_n3654_n3288# 0.402677f
C586 source.t47 a_n3654_n3288# 0.231396f
C587 source.t19 a_n3654_n3288# 0.231396f
C588 source.n354 a_n3654_n3288# 1.9812f
C589 source.n355 a_n3654_n3288# 0.402677f
C590 source.t12 a_n3654_n3288# 0.231396f
C591 source.t10 a_n3654_n3288# 0.231396f
C592 source.n356 a_n3654_n3288# 1.9812f
C593 source.n357 a_n3654_n3288# 0.402677f
C594 source.t18 a_n3654_n3288# 0.231396f
C595 source.t7 a_n3654_n3288# 0.231396f
C596 source.n358 a_n3654_n3288# 1.9812f
C597 source.n359 a_n3654_n3288# 0.402677f
C598 source.n360 a_n3654_n3288# 0.032323f
C599 source.n361 a_n3654_n3288# 0.024402f
C600 source.n362 a_n3654_n3288# 0.013112f
C601 source.n363 a_n3654_n3288# 0.030993f
C602 source.n364 a_n3654_n3288# 0.013884f
C603 source.n365 a_n3654_n3288# 0.024402f
C604 source.n366 a_n3654_n3288# 0.013112f
C605 source.n367 a_n3654_n3288# 0.030993f
C606 source.n368 a_n3654_n3288# 0.013884f
C607 source.n369 a_n3654_n3288# 0.024402f
C608 source.n370 a_n3654_n3288# 0.013498f
C609 source.n371 a_n3654_n3288# 0.030993f
C610 source.n372 a_n3654_n3288# 0.013884f
C611 source.n373 a_n3654_n3288# 0.024402f
C612 source.n374 a_n3654_n3288# 0.013112f
C613 source.n375 a_n3654_n3288# 0.030993f
C614 source.n376 a_n3654_n3288# 0.013884f
C615 source.n377 a_n3654_n3288# 0.024402f
C616 source.n378 a_n3654_n3288# 0.013112f
C617 source.n379 a_n3654_n3288# 0.023245f
C618 source.n380 a_n3654_n3288# 0.02191f
C619 source.t6 a_n3654_n3288# 0.052345f
C620 source.n381 a_n3654_n3288# 0.175934f
C621 source.n382 a_n3654_n3288# 1.23103f
C622 source.n383 a_n3654_n3288# 0.013112f
C623 source.n384 a_n3654_n3288# 0.013884f
C624 source.n385 a_n3654_n3288# 0.030993f
C625 source.n386 a_n3654_n3288# 0.030993f
C626 source.n387 a_n3654_n3288# 0.013884f
C627 source.n388 a_n3654_n3288# 0.013112f
C628 source.n389 a_n3654_n3288# 0.024402f
C629 source.n390 a_n3654_n3288# 0.024402f
C630 source.n391 a_n3654_n3288# 0.013112f
C631 source.n392 a_n3654_n3288# 0.013884f
C632 source.n393 a_n3654_n3288# 0.030993f
C633 source.n394 a_n3654_n3288# 0.030993f
C634 source.n395 a_n3654_n3288# 0.013884f
C635 source.n396 a_n3654_n3288# 0.013112f
C636 source.n397 a_n3654_n3288# 0.024402f
C637 source.n398 a_n3654_n3288# 0.024402f
C638 source.n399 a_n3654_n3288# 0.013112f
C639 source.n400 a_n3654_n3288# 0.013112f
C640 source.n401 a_n3654_n3288# 0.013884f
C641 source.n402 a_n3654_n3288# 0.030993f
C642 source.n403 a_n3654_n3288# 0.030993f
C643 source.n404 a_n3654_n3288# 0.030993f
C644 source.n405 a_n3654_n3288# 0.013498f
C645 source.n406 a_n3654_n3288# 0.013112f
C646 source.n407 a_n3654_n3288# 0.024402f
C647 source.n408 a_n3654_n3288# 0.024402f
C648 source.n409 a_n3654_n3288# 0.013112f
C649 source.n410 a_n3654_n3288# 0.013884f
C650 source.n411 a_n3654_n3288# 0.030993f
C651 source.n412 a_n3654_n3288# 0.030993f
C652 source.n413 a_n3654_n3288# 0.013884f
C653 source.n414 a_n3654_n3288# 0.013112f
C654 source.n415 a_n3654_n3288# 0.024402f
C655 source.n416 a_n3654_n3288# 0.024402f
C656 source.n417 a_n3654_n3288# 0.013112f
C657 source.n418 a_n3654_n3288# 0.013884f
C658 source.n419 a_n3654_n3288# 0.030993f
C659 source.n420 a_n3654_n3288# 0.063601f
C660 source.n421 a_n3654_n3288# 0.013884f
C661 source.n422 a_n3654_n3288# 0.013112f
C662 source.n423 a_n3654_n3288# 0.052403f
C663 source.n424 a_n3654_n3288# 0.035101f
C664 source.n425 a_n3654_n3288# 0.132123f
C665 source.n426 a_n3654_n3288# 0.032323f
C666 source.n427 a_n3654_n3288# 0.024402f
C667 source.n428 a_n3654_n3288# 0.013112f
C668 source.n429 a_n3654_n3288# 0.030993f
C669 source.n430 a_n3654_n3288# 0.013884f
C670 source.n431 a_n3654_n3288# 0.024402f
C671 source.n432 a_n3654_n3288# 0.013112f
C672 source.n433 a_n3654_n3288# 0.030993f
C673 source.n434 a_n3654_n3288# 0.013884f
C674 source.n435 a_n3654_n3288# 0.024402f
C675 source.n436 a_n3654_n3288# 0.013498f
C676 source.n437 a_n3654_n3288# 0.030993f
C677 source.n438 a_n3654_n3288# 0.013884f
C678 source.n439 a_n3654_n3288# 0.024402f
C679 source.n440 a_n3654_n3288# 0.013112f
C680 source.n441 a_n3654_n3288# 0.030993f
C681 source.n442 a_n3654_n3288# 0.013884f
C682 source.n443 a_n3654_n3288# 0.024402f
C683 source.n444 a_n3654_n3288# 0.013112f
C684 source.n445 a_n3654_n3288# 0.023245f
C685 source.n446 a_n3654_n3288# 0.02191f
C686 source.t24 a_n3654_n3288# 0.052345f
C687 source.n447 a_n3654_n3288# 0.175934f
C688 source.n448 a_n3654_n3288# 1.23103f
C689 source.n449 a_n3654_n3288# 0.013112f
C690 source.n450 a_n3654_n3288# 0.013884f
C691 source.n451 a_n3654_n3288# 0.030993f
C692 source.n452 a_n3654_n3288# 0.030993f
C693 source.n453 a_n3654_n3288# 0.013884f
C694 source.n454 a_n3654_n3288# 0.013112f
C695 source.n455 a_n3654_n3288# 0.024402f
C696 source.n456 a_n3654_n3288# 0.024402f
C697 source.n457 a_n3654_n3288# 0.013112f
C698 source.n458 a_n3654_n3288# 0.013884f
C699 source.n459 a_n3654_n3288# 0.030993f
C700 source.n460 a_n3654_n3288# 0.030993f
C701 source.n461 a_n3654_n3288# 0.013884f
C702 source.n462 a_n3654_n3288# 0.013112f
C703 source.n463 a_n3654_n3288# 0.024402f
C704 source.n464 a_n3654_n3288# 0.024402f
C705 source.n465 a_n3654_n3288# 0.013112f
C706 source.n466 a_n3654_n3288# 0.013112f
C707 source.n467 a_n3654_n3288# 0.013884f
C708 source.n468 a_n3654_n3288# 0.030993f
C709 source.n469 a_n3654_n3288# 0.030993f
C710 source.n470 a_n3654_n3288# 0.030993f
C711 source.n471 a_n3654_n3288# 0.013498f
C712 source.n472 a_n3654_n3288# 0.013112f
C713 source.n473 a_n3654_n3288# 0.024402f
C714 source.n474 a_n3654_n3288# 0.024402f
C715 source.n475 a_n3654_n3288# 0.013112f
C716 source.n476 a_n3654_n3288# 0.013884f
C717 source.n477 a_n3654_n3288# 0.030993f
C718 source.n478 a_n3654_n3288# 0.030993f
C719 source.n479 a_n3654_n3288# 0.013884f
C720 source.n480 a_n3654_n3288# 0.013112f
C721 source.n481 a_n3654_n3288# 0.024402f
C722 source.n482 a_n3654_n3288# 0.024402f
C723 source.n483 a_n3654_n3288# 0.013112f
C724 source.n484 a_n3654_n3288# 0.013884f
C725 source.n485 a_n3654_n3288# 0.030993f
C726 source.n486 a_n3654_n3288# 0.063601f
C727 source.n487 a_n3654_n3288# 0.013884f
C728 source.n488 a_n3654_n3288# 0.013112f
C729 source.n489 a_n3654_n3288# 0.052403f
C730 source.n490 a_n3654_n3288# 0.035101f
C731 source.n491 a_n3654_n3288# 0.132123f
C732 source.t20 a_n3654_n3288# 0.231396f
C733 source.t21 a_n3654_n3288# 0.231396f
C734 source.n492 a_n3654_n3288# 1.9812f
C735 source.n493 a_n3654_n3288# 0.402677f
C736 source.t38 a_n3654_n3288# 0.231396f
C737 source.t27 a_n3654_n3288# 0.231396f
C738 source.n494 a_n3654_n3288# 1.9812f
C739 source.n495 a_n3654_n3288# 0.402677f
C740 source.t31 a_n3654_n3288# 0.231396f
C741 source.t37 a_n3654_n3288# 0.231396f
C742 source.n496 a_n3654_n3288# 1.9812f
C743 source.n497 a_n3654_n3288# 0.402677f
C744 source.t22 a_n3654_n3288# 0.231396f
C745 source.t40 a_n3654_n3288# 0.231396f
C746 source.n498 a_n3654_n3288# 1.9812f
C747 source.n499 a_n3654_n3288# 0.402677f
C748 source.t26 a_n3654_n3288# 0.231396f
C749 source.t28 a_n3654_n3288# 0.231396f
C750 source.n500 a_n3654_n3288# 1.9812f
C751 source.n501 a_n3654_n3288# 0.402677f
C752 source.n502 a_n3654_n3288# 0.032323f
C753 source.n503 a_n3654_n3288# 0.024402f
C754 source.n504 a_n3654_n3288# 0.013112f
C755 source.n505 a_n3654_n3288# 0.030993f
C756 source.n506 a_n3654_n3288# 0.013884f
C757 source.n507 a_n3654_n3288# 0.024402f
C758 source.n508 a_n3654_n3288# 0.013112f
C759 source.n509 a_n3654_n3288# 0.030993f
C760 source.n510 a_n3654_n3288# 0.013884f
C761 source.n511 a_n3654_n3288# 0.024402f
C762 source.n512 a_n3654_n3288# 0.013498f
C763 source.n513 a_n3654_n3288# 0.030993f
C764 source.n514 a_n3654_n3288# 0.013884f
C765 source.n515 a_n3654_n3288# 0.024402f
C766 source.n516 a_n3654_n3288# 0.013112f
C767 source.n517 a_n3654_n3288# 0.030993f
C768 source.n518 a_n3654_n3288# 0.013884f
C769 source.n519 a_n3654_n3288# 0.024402f
C770 source.n520 a_n3654_n3288# 0.013112f
C771 source.n521 a_n3654_n3288# 0.023245f
C772 source.n522 a_n3654_n3288# 0.02191f
C773 source.t34 a_n3654_n3288# 0.052345f
C774 source.n523 a_n3654_n3288# 0.175934f
C775 source.n524 a_n3654_n3288# 1.23103f
C776 source.n525 a_n3654_n3288# 0.013112f
C777 source.n526 a_n3654_n3288# 0.013884f
C778 source.n527 a_n3654_n3288# 0.030993f
C779 source.n528 a_n3654_n3288# 0.030993f
C780 source.n529 a_n3654_n3288# 0.013884f
C781 source.n530 a_n3654_n3288# 0.013112f
C782 source.n531 a_n3654_n3288# 0.024402f
C783 source.n532 a_n3654_n3288# 0.024402f
C784 source.n533 a_n3654_n3288# 0.013112f
C785 source.n534 a_n3654_n3288# 0.013884f
C786 source.n535 a_n3654_n3288# 0.030993f
C787 source.n536 a_n3654_n3288# 0.030993f
C788 source.n537 a_n3654_n3288# 0.013884f
C789 source.n538 a_n3654_n3288# 0.013112f
C790 source.n539 a_n3654_n3288# 0.024402f
C791 source.n540 a_n3654_n3288# 0.024402f
C792 source.n541 a_n3654_n3288# 0.013112f
C793 source.n542 a_n3654_n3288# 0.013112f
C794 source.n543 a_n3654_n3288# 0.013884f
C795 source.n544 a_n3654_n3288# 0.030993f
C796 source.n545 a_n3654_n3288# 0.030993f
C797 source.n546 a_n3654_n3288# 0.030993f
C798 source.n547 a_n3654_n3288# 0.013498f
C799 source.n548 a_n3654_n3288# 0.013112f
C800 source.n549 a_n3654_n3288# 0.024402f
C801 source.n550 a_n3654_n3288# 0.024402f
C802 source.n551 a_n3654_n3288# 0.013112f
C803 source.n552 a_n3654_n3288# 0.013884f
C804 source.n553 a_n3654_n3288# 0.030993f
C805 source.n554 a_n3654_n3288# 0.030993f
C806 source.n555 a_n3654_n3288# 0.013884f
C807 source.n556 a_n3654_n3288# 0.013112f
C808 source.n557 a_n3654_n3288# 0.024402f
C809 source.n558 a_n3654_n3288# 0.024402f
C810 source.n559 a_n3654_n3288# 0.013112f
C811 source.n560 a_n3654_n3288# 0.013884f
C812 source.n561 a_n3654_n3288# 0.030993f
C813 source.n562 a_n3654_n3288# 0.063601f
C814 source.n563 a_n3654_n3288# 0.013884f
C815 source.n564 a_n3654_n3288# 0.013112f
C816 source.n565 a_n3654_n3288# 0.052403f
C817 source.n566 a_n3654_n3288# 0.035101f
C818 source.n567 a_n3654_n3288# 0.29658f
C819 source.n568 a_n3654_n3288# 1.55024f
C820 minus.n0 a_n3654_n3288# 0.049687f
C821 minus.t5 a_n3654_n3288# 1.01932f
C822 minus.n1 a_n3654_n3288# 0.41398f
C823 minus.t11 a_n3654_n3288# 1.01932f
C824 minus.n2 a_n3654_n3288# 0.037236f
C825 minus.t20 a_n3654_n3288# 1.01932f
C826 minus.n3 a_n3654_n3288# 0.403119f
C827 minus.n4 a_n3654_n3288# 0.062021f
C828 minus.n5 a_n3654_n3288# 0.00845f
C829 minus.t13 a_n3654_n3288# 1.01932f
C830 minus.n6 a_n3654_n3288# 0.037236f
C831 minus.n7 a_n3654_n3288# 0.00845f
C832 minus.t14 a_n3654_n3288# 1.01932f
C833 minus.t12 a_n3654_n3288# 1.03948f
C834 minus.n8 a_n3654_n3288# 0.38964f
C835 minus.t8 a_n3654_n3288# 1.01932f
C836 minus.n9 a_n3654_n3288# 0.41396f
C837 minus.t7 a_n3654_n3288# 1.01932f
C838 minus.n10 a_n3654_n3288# 0.41398f
C839 minus.n11 a_n3654_n3288# 0.214019f
C840 minus.n12 a_n3654_n3288# 0.049687f
C841 minus.n13 a_n3654_n3288# 0.037236f
C842 minus.n14 a_n3654_n3288# 0.403119f
C843 minus.n15 a_n3654_n3288# 0.00845f
C844 minus.t16 a_n3654_n3288# 1.01932f
C845 minus.n16 a_n3654_n3288# 0.403119f
C846 minus.n17 a_n3654_n3288# 0.037236f
C847 minus.n18 a_n3654_n3288# 0.049687f
C848 minus.n19 a_n3654_n3288# 0.062021f
C849 minus.n20 a_n3654_n3288# 0.41352f
C850 minus.t10 a_n3654_n3288# 1.01932f
C851 minus.n21 a_n3654_n3288# 0.41352f
C852 minus.n22 a_n3654_n3288# 0.00845f
C853 minus.n23 a_n3654_n3288# 0.049687f
C854 minus.n24 a_n3654_n3288# 0.037236f
C855 minus.n25 a_n3654_n3288# 0.037236f
C856 minus.n26 a_n3654_n3288# 0.00845f
C857 minus.t15 a_n3654_n3288# 1.01932f
C858 minus.n27 a_n3654_n3288# 0.403119f
C859 minus.n28 a_n3654_n3288# 0.00845f
C860 minus.n29 a_n3654_n3288# 0.049687f
C861 minus.n30 a_n3654_n3288# 0.062021f
C862 minus.n31 a_n3654_n3288# 0.062021f
C863 minus.n32 a_n3654_n3288# 0.413061f
C864 minus.n33 a_n3654_n3288# 0.00845f
C865 minus.t9 a_n3654_n3288# 1.01932f
C866 minus.n34 a_n3654_n3288# 0.40002f
C867 minus.n35 a_n3654_n3288# 1.71784f
C868 minus.n36 a_n3654_n3288# 0.049687f
C869 minus.t1 a_n3654_n3288# 1.01932f
C870 minus.n37 a_n3654_n3288# 0.41398f
C871 minus.n38 a_n3654_n3288# 0.037236f
C872 minus.t0 a_n3654_n3288# 1.01932f
C873 minus.n39 a_n3654_n3288# 0.403119f
C874 minus.n40 a_n3654_n3288# 0.062021f
C875 minus.n41 a_n3654_n3288# 0.00845f
C876 minus.n42 a_n3654_n3288# 0.037236f
C877 minus.n43 a_n3654_n3288# 0.00845f
C878 minus.t23 a_n3654_n3288# 1.03948f
C879 minus.n44 a_n3654_n3288# 0.38964f
C880 minus.t6 a_n3654_n3288# 1.01932f
C881 minus.n45 a_n3654_n3288# 0.41396f
C882 minus.t19 a_n3654_n3288# 1.01932f
C883 minus.n46 a_n3654_n3288# 0.41398f
C884 minus.n47 a_n3654_n3288# 0.214019f
C885 minus.n48 a_n3654_n3288# 0.049687f
C886 minus.n49 a_n3654_n3288# 0.037236f
C887 minus.t3 a_n3654_n3288# 1.01932f
C888 minus.n50 a_n3654_n3288# 0.403119f
C889 minus.n51 a_n3654_n3288# 0.00845f
C890 minus.t22 a_n3654_n3288# 1.01932f
C891 minus.n52 a_n3654_n3288# 0.403119f
C892 minus.n53 a_n3654_n3288# 0.037236f
C893 minus.n54 a_n3654_n3288# 0.049687f
C894 minus.n55 a_n3654_n3288# 0.062021f
C895 minus.t2 a_n3654_n3288# 1.01932f
C896 minus.n56 a_n3654_n3288# 0.41352f
C897 minus.t17 a_n3654_n3288# 1.01932f
C898 minus.n57 a_n3654_n3288# 0.41352f
C899 minus.n58 a_n3654_n3288# 0.00845f
C900 minus.n59 a_n3654_n3288# 0.049687f
C901 minus.n60 a_n3654_n3288# 0.037236f
C902 minus.n61 a_n3654_n3288# 0.037236f
C903 minus.n62 a_n3654_n3288# 0.00845f
C904 minus.t18 a_n3654_n3288# 1.01932f
C905 minus.n63 a_n3654_n3288# 0.403119f
C906 minus.n64 a_n3654_n3288# 0.00845f
C907 minus.n65 a_n3654_n3288# 0.049687f
C908 minus.n66 a_n3654_n3288# 0.062021f
C909 minus.n67 a_n3654_n3288# 0.062021f
C910 minus.t4 a_n3654_n3288# 1.01932f
C911 minus.n68 a_n3654_n3288# 0.413061f
C912 minus.n69 a_n3654_n3288# 0.00845f
C913 minus.t21 a_n3654_n3288# 1.01932f
C914 minus.n70 a_n3654_n3288# 0.40002f
C915 minus.n71 a_n3654_n3288# 0.257336f
C916 minus.n72 a_n3654_n3288# 2.04187f
.ends

