* NGSPICE file created from diffpair648.ext - technology: sky130A

.subckt diffpair648 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t27 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 source.t12 plus.t0 drain_left.t19 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X2 drain_right.t18 minus.t1 source.t19 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X3 source.t37 minus.t2 drain_right.t17 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X4 a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X5 source.t15 plus.t1 drain_left.t18 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X6 a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X7 a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X8 drain_left.t17 plus.t2 source.t3 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X9 source.t7 plus.t3 drain_left.t16 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X10 drain_left.t15 plus.t4 source.t2 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X11 source.t25 minus.t3 drain_right.t16 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X12 source.t0 plus.t5 drain_left.t14 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X13 a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X14 drain_left.t13 plus.t6 source.t17 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X15 drain_right.t15 minus.t4 source.t23 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X16 drain_right.t14 minus.t5 source.t30 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 source.t32 minus.t6 drain_right.t13 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X18 source.t34 minus.t7 drain_right.t12 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 drain_left.t12 plus.t7 source.t16 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X20 source.t36 minus.t8 drain_right.t11 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X21 drain_right.t10 minus.t9 source.t21 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 drain_left.t11 plus.t8 source.t9 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X23 drain_left.t10 plus.t9 source.t8 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X24 source.t38 plus.t10 drain_left.t9 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X25 drain_right.t9 minus.t10 source.t28 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X26 drain_right.t8 minus.t11 source.t20 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X27 drain_right.t7 minus.t12 source.t26 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X28 source.t18 minus.t13 drain_right.t6 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X29 drain_left.t8 plus.t11 source.t39 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X30 source.t35 minus.t14 drain_right.t5 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X31 drain_right.t4 minus.t15 source.t24 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X32 drain_right.t3 minus.t16 source.t22 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X33 source.t4 plus.t12 drain_left.t7 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X34 drain_left.t6 plus.t13 source.t6 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X35 source.t1 plus.t14 drain_left.t5 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X36 source.t11 plus.t15 drain_left.t4 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X37 source.t29 minus.t17 drain_right.t2 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X38 source.t14 plus.t16 drain_left.t3 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X39 drain_left.t2 plus.t17 source.t5 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X40 drain_left.t1 plus.t18 source.t10 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X41 source.t31 minus.t18 drain_right.t1 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X42 source.t13 plus.t19 drain_left.t0 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X43 source.t33 minus.t19 drain_right.t0 a_n2146_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
R0 minus.n27 minus.t17 4287.61
R1 minus.n7 minus.t4 4287.61
R2 minus.n56 minus.t16 4287.61
R3 minus.n35 minus.t2 4287.61
R4 minus.n26 minus.t9 4225.53
R5 minus.n24 minus.t13 4225.53
R6 minus.n3 minus.t11 4225.53
R7 minus.n18 minus.t14 4225.53
R8 minus.n16 minus.t5 4225.53
R9 minus.n4 minus.t8 4225.53
R10 minus.n10 minus.t10 4225.53
R11 minus.n6 minus.t3 4225.53
R12 minus.n55 minus.t7 4225.53
R13 minus.n53 minus.t1 4225.53
R14 minus.n47 minus.t19 4225.53
R15 minus.n46 minus.t15 4225.53
R16 minus.n44 minus.t6 4225.53
R17 minus.n32 minus.t0 4225.53
R18 minus.n38 minus.t18 4225.53
R19 minus.n34 minus.t12 4225.53
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 69.3793
R47 minus.n15 minus.n4 69.3793
R48 minus.n43 minus.n32 69.3793
R49 minus.n48 minus.n47 69.3793
R50 minus.n25 minus.n24 54.7732
R51 minus.n10 minus.n9 54.7732
R52 minus.n38 minus.n37 54.7732
R53 minus.n54 minus.n53 54.7732
R54 minus.n18 minus.n17 47.4702
R55 minus.n17 minus.n16 47.4702
R56 minus.n45 minus.n44 47.4702
R57 minus.n46 minus.n45 47.4702
R58 minus.n58 minus.n28 47.1596
R59 minus.n26 minus.n25 40.1672
R60 minus.n9 minus.n6 40.1672
R61 minus.n37 minus.n34 40.1672
R62 minus.n55 minus.n54 40.1672
R63 minus.n27 minus.n26 32.8641
R64 minus.n7 minus.n6 32.8641
R65 minus.n35 minus.n34 32.8641
R66 minus.n56 minus.n55 32.8641
R67 minus.n19 minus.n18 25.5611
R68 minus.n16 minus.n15 25.5611
R69 minus.n44 minus.n43 25.5611
R70 minus.n48 minus.n46 25.5611
R71 minus.n24 minus.n23 18.2581
R72 minus.n11 minus.n10 18.2581
R73 minus.n39 minus.n38 18.2581
R74 minus.n53 minus.n52 18.2581
R75 minus.n58 minus.n57 6.56111
R76 minus.n3 minus.n1 3.65202
R77 minus.n12 minus.n4 3.65202
R78 minus.n40 minus.n32 3.65202
R79 minus.n47 minus.n30 3.65202
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 source.n9 source.t38 43.2366
R100 source.n10 source.t23 43.2366
R101 source.n19 source.t29 43.2366
R102 source.n39 source.t22 43.2365
R103 source.n30 source.t37 43.2365
R104 source.n29 source.t16 43.2365
R105 source.n20 source.t12 43.2365
R106 source.n0 source.t6 43.2365
R107 source.n38 source.n37 42.0366
R108 source.n36 source.n35 42.0366
R109 source.n34 source.n33 42.0366
R110 source.n32 source.n31 42.0366
R111 source.n28 source.n27 42.0366
R112 source.n26 source.n25 42.0366
R113 source.n24 source.n23 42.0366
R114 source.n22 source.n21 42.0366
R115 source.n2 source.n1 42.0366
R116 source.n4 source.n3 42.0366
R117 source.n6 source.n5 42.0366
R118 source.n8 source.n7 42.0366
R119 source.n12 source.n11 42.0366
R120 source.n14 source.n13 42.0366
R121 source.n16 source.n15 42.0366
R122 source.n18 source.n17 42.0366
R123 source.n20 source.n19 31.6966
R124 source.n40 source.n0 26.1535
R125 source.n40 source.n39 5.5436
R126 source.n37 source.t19 1.2005
R127 source.n37 source.t34 1.2005
R128 source.n35 source.t24 1.2005
R129 source.n35 source.t33 1.2005
R130 source.n33 source.t27 1.2005
R131 source.n33 source.t32 1.2005
R132 source.n31 source.t26 1.2005
R133 source.n31 source.t31 1.2005
R134 source.n27 source.t3 1.2005
R135 source.n27 source.t4 1.2005
R136 source.n25 source.t9 1.2005
R137 source.n25 source.t0 1.2005
R138 source.n23 source.t2 1.2005
R139 source.n23 source.t15 1.2005
R140 source.n21 source.t17 1.2005
R141 source.n21 source.t7 1.2005
R142 source.n1 source.t8 1.2005
R143 source.n1 source.t14 1.2005
R144 source.n3 source.t5 1.2005
R145 source.n3 source.t1 1.2005
R146 source.n5 source.t39 1.2005
R147 source.n5 source.t13 1.2005
R148 source.n7 source.t10 1.2005
R149 source.n7 source.t11 1.2005
R150 source.n11 source.t28 1.2005
R151 source.n11 source.t25 1.2005
R152 source.n13 source.t30 1.2005
R153 source.n13 source.t36 1.2005
R154 source.n15 source.t20 1.2005
R155 source.n15 source.t35 1.2005
R156 source.n17 source.t21 1.2005
R157 source.n17 source.t18 1.2005
R158 source.n19 source.n18 0.560845
R159 source.n18 source.n16 0.560845
R160 source.n16 source.n14 0.560845
R161 source.n14 source.n12 0.560845
R162 source.n12 source.n10 0.560845
R163 source.n9 source.n8 0.560845
R164 source.n8 source.n6 0.560845
R165 source.n6 source.n4 0.560845
R166 source.n4 source.n2 0.560845
R167 source.n2 source.n0 0.560845
R168 source.n22 source.n20 0.560845
R169 source.n24 source.n22 0.560845
R170 source.n26 source.n24 0.560845
R171 source.n28 source.n26 0.560845
R172 source.n29 source.n28 0.560845
R173 source.n32 source.n30 0.560845
R174 source.n34 source.n32 0.560845
R175 source.n36 source.n34 0.560845
R176 source.n38 source.n36 0.560845
R177 source.n39 source.n38 0.560845
R178 source.n10 source.n9 0.470328
R179 source.n30 source.n29 0.470328
R180 source source.n40 0.188
R181 drain_right.n6 drain_right.n4 59.2758
R182 drain_right.n2 drain_right.n0 59.2758
R183 drain_right.n10 drain_right.n8 59.2756
R184 drain_right.n7 drain_right.n3 58.7154
R185 drain_right.n6 drain_right.n5 58.7154
R186 drain_right.n2 drain_right.n1 58.7154
R187 drain_right.n10 drain_right.n9 58.7154
R188 drain_right.n12 drain_right.n11 58.7154
R189 drain_right.n14 drain_right.n13 58.7154
R190 drain_right.n16 drain_right.n15 58.7154
R191 drain_right drain_right.n7 41.1451
R192 drain_right drain_right.n16 6.21356
R193 drain_right.n3 drain_right.t13 1.2005
R194 drain_right.n3 drain_right.t4 1.2005
R195 drain_right.n4 drain_right.t12 1.2005
R196 drain_right.n4 drain_right.t3 1.2005
R197 drain_right.n5 drain_right.t0 1.2005
R198 drain_right.n5 drain_right.t18 1.2005
R199 drain_right.n1 drain_right.t1 1.2005
R200 drain_right.n1 drain_right.t19 1.2005
R201 drain_right.n0 drain_right.t17 1.2005
R202 drain_right.n0 drain_right.t7 1.2005
R203 drain_right.n8 drain_right.t16 1.2005
R204 drain_right.n8 drain_right.t15 1.2005
R205 drain_right.n9 drain_right.t11 1.2005
R206 drain_right.n9 drain_right.t9 1.2005
R207 drain_right.n11 drain_right.t5 1.2005
R208 drain_right.n11 drain_right.t14 1.2005
R209 drain_right.n13 drain_right.t6 1.2005
R210 drain_right.n13 drain_right.t8 1.2005
R211 drain_right.n15 drain_right.t2 1.2005
R212 drain_right.n15 drain_right.t10 1.2005
R213 drain_right.n16 drain_right.n14 0.560845
R214 drain_right.n14 drain_right.n12 0.560845
R215 drain_right.n12 drain_right.n10 0.560845
R216 drain_right.n7 drain_right.n6 0.505499
R217 drain_right.n7 drain_right.n2 0.505499
R218 plus.n6 plus.t10 4287.61
R219 plus.n27 plus.t13 4287.61
R220 plus.n36 plus.t7 4287.61
R221 plus.n56 plus.t0 4287.61
R222 plus.n5 plus.t18 4225.53
R223 plus.n9 plus.t15 4225.53
R224 plus.n3 plus.t11 4225.53
R225 plus.n15 plus.t19 4225.53
R226 plus.n17 plus.t17 4225.53
R227 plus.n18 plus.t14 4225.53
R228 plus.n24 plus.t9 4225.53
R229 plus.n26 plus.t16 4225.53
R230 plus.n35 plus.t12 4225.53
R231 plus.n39 plus.t2 4225.53
R232 plus.n33 plus.t5 4225.53
R233 plus.n45 plus.t8 4225.53
R234 plus.n47 plus.t1 4225.53
R235 plus.n32 plus.t4 4225.53
R236 plus.n53 plus.t3 4225.53
R237 plus.n55 plus.t6 4225.53
R238 plus.n7 plus.n6 161.489
R239 plus.n37 plus.n36 161.489
R240 plus.n8 plus.n7 161.3
R241 plus.n10 plus.n4 161.3
R242 plus.n12 plus.n11 161.3
R243 plus.n14 plus.n13 161.3
R244 plus.n16 plus.n2 161.3
R245 plus.n20 plus.n19 161.3
R246 plus.n21 plus.n1 161.3
R247 plus.n23 plus.n22 161.3
R248 plus.n25 plus.n0 161.3
R249 plus.n28 plus.n27 161.3
R250 plus.n38 plus.n37 161.3
R251 plus.n40 plus.n34 161.3
R252 plus.n42 plus.n41 161.3
R253 plus.n44 plus.n43 161.3
R254 plus.n46 plus.n31 161.3
R255 plus.n49 plus.n48 161.3
R256 plus.n50 plus.n30 161.3
R257 plus.n52 plus.n51 161.3
R258 plus.n54 plus.n29 161.3
R259 plus.n57 plus.n56 161.3
R260 plus.n11 plus.n10 73.0308
R261 plus.n23 plus.n1 73.0308
R262 plus.n52 plus.n30 73.0308
R263 plus.n41 plus.n40 73.0308
R264 plus.n14 plus.n3 69.3793
R265 plus.n19 plus.n18 69.3793
R266 plus.n48 plus.n32 69.3793
R267 plus.n44 plus.n33 69.3793
R268 plus.n9 plus.n8 54.7732
R269 plus.n25 plus.n24 54.7732
R270 plus.n54 plus.n53 54.7732
R271 plus.n39 plus.n38 54.7732
R272 plus.n16 plus.n15 47.4702
R273 plus.n17 plus.n16 47.4702
R274 plus.n47 plus.n46 47.4702
R275 plus.n46 plus.n45 47.4702
R276 plus.n8 plus.n5 40.1672
R277 plus.n26 plus.n25 40.1672
R278 plus.n55 plus.n54 40.1672
R279 plus.n38 plus.n35 40.1672
R280 plus plus.n57 36.1164
R281 plus.n6 plus.n5 32.8641
R282 plus.n27 plus.n26 32.8641
R283 plus.n56 plus.n55 32.8641
R284 plus.n36 plus.n35 32.8641
R285 plus.n15 plus.n14 25.5611
R286 plus.n19 plus.n17 25.5611
R287 plus.n48 plus.n47 25.5611
R288 plus.n45 plus.n44 25.5611
R289 plus.n10 plus.n9 18.2581
R290 plus.n24 plus.n23 18.2581
R291 plus.n53 plus.n52 18.2581
R292 plus.n40 plus.n39 18.2581
R293 plus plus.n28 17.1293
R294 plus.n11 plus.n3 3.65202
R295 plus.n18 plus.n1 3.65202
R296 plus.n32 plus.n30 3.65202
R297 plus.n41 plus.n33 3.65202
R298 plus.n7 plus.n4 0.189894
R299 plus.n12 plus.n4 0.189894
R300 plus.n13 plus.n12 0.189894
R301 plus.n13 plus.n2 0.189894
R302 plus.n20 plus.n2 0.189894
R303 plus.n21 plus.n20 0.189894
R304 plus.n22 plus.n21 0.189894
R305 plus.n22 plus.n0 0.189894
R306 plus.n28 plus.n0 0.189894
R307 plus.n57 plus.n29 0.189894
R308 plus.n51 plus.n29 0.189894
R309 plus.n51 plus.n50 0.189894
R310 plus.n50 plus.n49 0.189894
R311 plus.n49 plus.n31 0.189894
R312 plus.n43 plus.n31 0.189894
R313 plus.n43 plus.n42 0.189894
R314 plus.n42 plus.n34 0.189894
R315 plus.n37 plus.n34 0.189894
R316 drain_left.n6 drain_left.n4 59.2758
R317 drain_left.n2 drain_left.n0 59.2758
R318 drain_left.n10 drain_left.n8 59.2758
R319 drain_left.n7 drain_left.n3 58.7154
R320 drain_left.n6 drain_left.n5 58.7154
R321 drain_left.n2 drain_left.n1 58.7154
R322 drain_left.n14 drain_left.n13 58.7154
R323 drain_left.n12 drain_left.n11 58.7154
R324 drain_left.n10 drain_left.n9 58.7154
R325 drain_left.n16 drain_left.n15 58.7153
R326 drain_left drain_left.n7 41.6983
R327 drain_left drain_left.n16 6.21356
R328 drain_left.n3 drain_left.t18 1.2005
R329 drain_left.n3 drain_left.t11 1.2005
R330 drain_left.n4 drain_left.t7 1.2005
R331 drain_left.n4 drain_left.t12 1.2005
R332 drain_left.n5 drain_left.t14 1.2005
R333 drain_left.n5 drain_left.t17 1.2005
R334 drain_left.n1 drain_left.t16 1.2005
R335 drain_left.n1 drain_left.t15 1.2005
R336 drain_left.n0 drain_left.t19 1.2005
R337 drain_left.n0 drain_left.t13 1.2005
R338 drain_left.n15 drain_left.t3 1.2005
R339 drain_left.n15 drain_left.t6 1.2005
R340 drain_left.n13 drain_left.t5 1.2005
R341 drain_left.n13 drain_left.t10 1.2005
R342 drain_left.n11 drain_left.t0 1.2005
R343 drain_left.n11 drain_left.t2 1.2005
R344 drain_left.n9 drain_left.t4 1.2005
R345 drain_left.n9 drain_left.t8 1.2005
R346 drain_left.n8 drain_left.t9 1.2005
R347 drain_left.n8 drain_left.t1 1.2005
R348 drain_left.n12 drain_left.n10 0.560845
R349 drain_left.n14 drain_left.n12 0.560845
R350 drain_left.n16 drain_left.n14 0.560845
R351 drain_left.n7 drain_left.n6 0.505499
R352 drain_left.n7 drain_left.n2 0.505499
C0 plus minus 8.220281f
C1 drain_right minus 8.13969f
C2 plus drain_left 8.35037f
C3 drain_left drain_right 1.13563f
C4 plus source 7.07977f
C5 drain_right source 76.01679f
C6 plus drain_right 0.364841f
C7 drain_left minus 0.171338f
C8 source minus 7.06573f
C9 drain_left source 76.0163f
C10 drain_right a_n2146_n5888# 8.81905f
C11 drain_left a_n2146_n5888# 9.13696f
C12 source a_n2146_n5888# 15.873385f
C13 minus a_n2146_n5888# 8.804264f
C14 plus a_n2146_n5888# 11.89727f
C15 drain_left.t19 a_n2146_n5888# 0.84572f
C16 drain_left.t13 a_n2146_n5888# 0.84572f
C17 drain_left.n0 a_n2146_n5888# 5.72261f
C18 drain_left.t16 a_n2146_n5888# 0.84572f
C19 drain_left.t15 a_n2146_n5888# 0.84572f
C20 drain_left.n1 a_n2146_n5888# 5.71928f
C21 drain_left.n2 a_n2146_n5888# 0.686018f
C22 drain_left.t18 a_n2146_n5888# 0.84572f
C23 drain_left.t11 a_n2146_n5888# 0.84572f
C24 drain_left.n3 a_n2146_n5888# 5.71928f
C25 drain_left.t7 a_n2146_n5888# 0.84572f
C26 drain_left.t12 a_n2146_n5888# 0.84572f
C27 drain_left.n4 a_n2146_n5888# 5.72261f
C28 drain_left.t14 a_n2146_n5888# 0.84572f
C29 drain_left.t17 a_n2146_n5888# 0.84572f
C30 drain_left.n5 a_n2146_n5888# 5.71928f
C31 drain_left.n6 a_n2146_n5888# 0.686018f
C32 drain_left.n7 a_n2146_n5888# 2.69193f
C33 drain_left.t9 a_n2146_n5888# 0.84572f
C34 drain_left.t1 a_n2146_n5888# 0.84572f
C35 drain_left.n8 a_n2146_n5888# 5.72261f
C36 drain_left.t4 a_n2146_n5888# 0.84572f
C37 drain_left.t8 a_n2146_n5888# 0.84572f
C38 drain_left.n9 a_n2146_n5888# 5.71928f
C39 drain_left.n10 a_n2146_n5888# 0.689756f
C40 drain_left.t0 a_n2146_n5888# 0.84572f
C41 drain_left.t2 a_n2146_n5888# 0.84572f
C42 drain_left.n11 a_n2146_n5888# 5.71928f
C43 drain_left.n12 a_n2146_n5888# 0.340853f
C44 drain_left.t5 a_n2146_n5888# 0.84572f
C45 drain_left.t10 a_n2146_n5888# 0.84572f
C46 drain_left.n13 a_n2146_n5888# 5.71928f
C47 drain_left.n14 a_n2146_n5888# 0.340853f
C48 drain_left.t3 a_n2146_n5888# 0.84572f
C49 drain_left.t6 a_n2146_n5888# 0.84572f
C50 drain_left.n15 a_n2146_n5888# 5.71927f
C51 drain_left.n16 a_n2146_n5888# 0.576815f
C52 plus.n0 a_n2146_n5888# 0.053864f
C53 plus.t16 a_n2146_n5888# 0.568332f
C54 plus.t9 a_n2146_n5888# 0.568332f
C55 plus.n1 a_n2146_n5888# 0.018699f
C56 plus.n2 a_n2146_n5888# 0.053864f
C57 plus.t17 a_n2146_n5888# 0.568332f
C58 plus.t19 a_n2146_n5888# 0.568332f
C59 plus.t11 a_n2146_n5888# 0.568332f
C60 plus.n3 a_n2146_n5888# 0.215106f
C61 plus.n4 a_n2146_n5888# 0.053864f
C62 plus.t15 a_n2146_n5888# 0.568332f
C63 plus.t18 a_n2146_n5888# 0.568332f
C64 plus.n5 a_n2146_n5888# 0.215106f
C65 plus.t10 a_n2146_n5888# 0.571482f
C66 plus.n6 a_n2146_n5888# 0.237378f
C67 plus.n7 a_n2146_n5888# 0.124249f
C68 plus.n8 a_n2146_n5888# 0.02285f
C69 plus.n9 a_n2146_n5888# 0.215106f
C70 plus.n10 a_n2146_n5888# 0.022019f
C71 plus.n11 a_n2146_n5888# 0.018699f
C72 plus.n12 a_n2146_n5888# 0.053864f
C73 plus.n13 a_n2146_n5888# 0.053864f
C74 plus.n14 a_n2146_n5888# 0.02285f
C75 plus.n15 a_n2146_n5888# 0.215106f
C76 plus.n16 a_n2146_n5888# 0.02285f
C77 plus.n17 a_n2146_n5888# 0.215106f
C78 plus.t14 a_n2146_n5888# 0.568332f
C79 plus.n18 a_n2146_n5888# 0.215106f
C80 plus.n19 a_n2146_n5888# 0.02285f
C81 plus.n20 a_n2146_n5888# 0.053864f
C82 plus.n21 a_n2146_n5888# 0.053864f
C83 plus.n22 a_n2146_n5888# 0.053864f
C84 plus.n23 a_n2146_n5888# 0.022019f
C85 plus.n24 a_n2146_n5888# 0.215106f
C86 plus.n25 a_n2146_n5888# 0.02285f
C87 plus.n26 a_n2146_n5888# 0.215106f
C88 plus.t13 a_n2146_n5888# 0.571482f
C89 plus.n27 a_n2146_n5888# 0.237296f
C90 plus.n28 a_n2146_n5888# 0.968898f
C91 plus.n29 a_n2146_n5888# 0.053864f
C92 plus.t0 a_n2146_n5888# 0.571482f
C93 plus.t6 a_n2146_n5888# 0.568332f
C94 plus.t3 a_n2146_n5888# 0.568332f
C95 plus.n30 a_n2146_n5888# 0.018699f
C96 plus.n31 a_n2146_n5888# 0.053864f
C97 plus.t4 a_n2146_n5888# 0.568332f
C98 plus.n32 a_n2146_n5888# 0.215106f
C99 plus.t1 a_n2146_n5888# 0.568332f
C100 plus.t8 a_n2146_n5888# 0.568332f
C101 plus.t5 a_n2146_n5888# 0.568332f
C102 plus.n33 a_n2146_n5888# 0.215106f
C103 plus.n34 a_n2146_n5888# 0.053864f
C104 plus.t2 a_n2146_n5888# 0.568332f
C105 plus.t12 a_n2146_n5888# 0.568332f
C106 plus.n35 a_n2146_n5888# 0.215106f
C107 plus.t7 a_n2146_n5888# 0.571482f
C108 plus.n36 a_n2146_n5888# 0.237378f
C109 plus.n37 a_n2146_n5888# 0.124249f
C110 plus.n38 a_n2146_n5888# 0.02285f
C111 plus.n39 a_n2146_n5888# 0.215106f
C112 plus.n40 a_n2146_n5888# 0.022019f
C113 plus.n41 a_n2146_n5888# 0.018699f
C114 plus.n42 a_n2146_n5888# 0.053864f
C115 plus.n43 a_n2146_n5888# 0.053864f
C116 plus.n44 a_n2146_n5888# 0.02285f
C117 plus.n45 a_n2146_n5888# 0.215106f
C118 plus.n46 a_n2146_n5888# 0.02285f
C119 plus.n47 a_n2146_n5888# 0.215106f
C120 plus.n48 a_n2146_n5888# 0.02285f
C121 plus.n49 a_n2146_n5888# 0.053864f
C122 plus.n50 a_n2146_n5888# 0.053864f
C123 plus.n51 a_n2146_n5888# 0.053864f
C124 plus.n52 a_n2146_n5888# 0.022019f
C125 plus.n53 a_n2146_n5888# 0.215106f
C126 plus.n54 a_n2146_n5888# 0.02285f
C127 plus.n55 a_n2146_n5888# 0.215106f
C128 plus.n56 a_n2146_n5888# 0.237296f
C129 plus.n57 a_n2146_n5888# 2.17111f
C130 drain_right.t17 a_n2146_n5888# 0.843819f
C131 drain_right.t7 a_n2146_n5888# 0.843819f
C132 drain_right.n0 a_n2146_n5888# 5.70974f
C133 drain_right.t1 a_n2146_n5888# 0.843819f
C134 drain_right.t19 a_n2146_n5888# 0.843819f
C135 drain_right.n1 a_n2146_n5888# 5.70642f
C136 drain_right.n2 a_n2146_n5888# 0.684476f
C137 drain_right.t13 a_n2146_n5888# 0.843819f
C138 drain_right.t4 a_n2146_n5888# 0.843819f
C139 drain_right.n3 a_n2146_n5888# 5.70642f
C140 drain_right.t12 a_n2146_n5888# 0.843819f
C141 drain_right.t3 a_n2146_n5888# 0.843819f
C142 drain_right.n4 a_n2146_n5888# 5.70974f
C143 drain_right.t0 a_n2146_n5888# 0.843819f
C144 drain_right.t18 a_n2146_n5888# 0.843819f
C145 drain_right.n5 a_n2146_n5888# 5.70642f
C146 drain_right.n6 a_n2146_n5888# 0.684476f
C147 drain_right.n7 a_n2146_n5888# 2.62767f
C148 drain_right.t16 a_n2146_n5888# 0.843819f
C149 drain_right.t15 a_n2146_n5888# 0.843819f
C150 drain_right.n8 a_n2146_n5888# 5.70973f
C151 drain_right.t11 a_n2146_n5888# 0.843819f
C152 drain_right.t9 a_n2146_n5888# 0.843819f
C153 drain_right.n9 a_n2146_n5888# 5.70642f
C154 drain_right.n10 a_n2146_n5888# 0.688219f
C155 drain_right.t5 a_n2146_n5888# 0.843819f
C156 drain_right.t14 a_n2146_n5888# 0.843819f
C157 drain_right.n11 a_n2146_n5888# 5.70642f
C158 drain_right.n12 a_n2146_n5888# 0.340087f
C159 drain_right.t6 a_n2146_n5888# 0.843819f
C160 drain_right.t8 a_n2146_n5888# 0.843819f
C161 drain_right.n13 a_n2146_n5888# 5.70642f
C162 drain_right.n14 a_n2146_n5888# 0.340087f
C163 drain_right.t2 a_n2146_n5888# 0.843819f
C164 drain_right.t10 a_n2146_n5888# 0.843819f
C165 drain_right.n15 a_n2146_n5888# 5.70642f
C166 drain_right.n16 a_n2146_n5888# 0.575506f
C167 source.t6 a_n2146_n5888# 5.96585f
C168 source.n0 a_n2146_n5888# 2.28282f
C169 source.t8 a_n2146_n5888# 0.723465f
C170 source.t14 a_n2146_n5888# 0.723465f
C171 source.n1 a_n2146_n5888# 4.81328f
C172 source.n2 a_n2146_n5888# 0.337964f
C173 source.t5 a_n2146_n5888# 0.723465f
C174 source.t1 a_n2146_n5888# 0.723465f
C175 source.n3 a_n2146_n5888# 4.81328f
C176 source.n4 a_n2146_n5888# 0.337964f
C177 source.t39 a_n2146_n5888# 0.723465f
C178 source.t13 a_n2146_n5888# 0.723465f
C179 source.n5 a_n2146_n5888# 4.81328f
C180 source.n6 a_n2146_n5888# 0.337964f
C181 source.t10 a_n2146_n5888# 0.723465f
C182 source.t11 a_n2146_n5888# 0.723465f
C183 source.n7 a_n2146_n5888# 4.81328f
C184 source.n8 a_n2146_n5888# 0.337964f
C185 source.t38 a_n2146_n5888# 5.96586f
C186 source.n9 a_n2146_n5888# 0.480569f
C187 source.t23 a_n2146_n5888# 5.96586f
C188 source.n10 a_n2146_n5888# 0.480569f
C189 source.t28 a_n2146_n5888# 0.723465f
C190 source.t25 a_n2146_n5888# 0.723465f
C191 source.n11 a_n2146_n5888# 4.81328f
C192 source.n12 a_n2146_n5888# 0.337964f
C193 source.t30 a_n2146_n5888# 0.723465f
C194 source.t36 a_n2146_n5888# 0.723465f
C195 source.n13 a_n2146_n5888# 4.81328f
C196 source.n14 a_n2146_n5888# 0.337964f
C197 source.t20 a_n2146_n5888# 0.723465f
C198 source.t35 a_n2146_n5888# 0.723465f
C199 source.n15 a_n2146_n5888# 4.81328f
C200 source.n16 a_n2146_n5888# 0.337964f
C201 source.t21 a_n2146_n5888# 0.723465f
C202 source.t18 a_n2146_n5888# 0.723465f
C203 source.n17 a_n2146_n5888# 4.81328f
C204 source.n18 a_n2146_n5888# 0.337964f
C205 source.t29 a_n2146_n5888# 5.96586f
C206 source.n19 a_n2146_n5888# 2.73053f
C207 source.t12 a_n2146_n5888# 5.96585f
C208 source.n20 a_n2146_n5888# 2.73055f
C209 source.t17 a_n2146_n5888# 0.723465f
C210 source.t7 a_n2146_n5888# 0.723465f
C211 source.n21 a_n2146_n5888# 4.81328f
C212 source.n22 a_n2146_n5888# 0.337966f
C213 source.t2 a_n2146_n5888# 0.723465f
C214 source.t15 a_n2146_n5888# 0.723465f
C215 source.n23 a_n2146_n5888# 4.81328f
C216 source.n24 a_n2146_n5888# 0.337966f
C217 source.t9 a_n2146_n5888# 0.723465f
C218 source.t0 a_n2146_n5888# 0.723465f
C219 source.n25 a_n2146_n5888# 4.81328f
C220 source.n26 a_n2146_n5888# 0.337966f
C221 source.t3 a_n2146_n5888# 0.723465f
C222 source.t4 a_n2146_n5888# 0.723465f
C223 source.n27 a_n2146_n5888# 4.81328f
C224 source.n28 a_n2146_n5888# 0.337966f
C225 source.t16 a_n2146_n5888# 5.96585f
C226 source.n29 a_n2146_n5888# 0.480585f
C227 source.t37 a_n2146_n5888# 5.96585f
C228 source.n30 a_n2146_n5888# 0.480585f
C229 source.t26 a_n2146_n5888# 0.723465f
C230 source.t31 a_n2146_n5888# 0.723465f
C231 source.n31 a_n2146_n5888# 4.81328f
C232 source.n32 a_n2146_n5888# 0.337966f
C233 source.t27 a_n2146_n5888# 0.723465f
C234 source.t32 a_n2146_n5888# 0.723465f
C235 source.n33 a_n2146_n5888# 4.81328f
C236 source.n34 a_n2146_n5888# 0.337966f
C237 source.t24 a_n2146_n5888# 0.723465f
C238 source.t33 a_n2146_n5888# 0.723465f
C239 source.n35 a_n2146_n5888# 4.81328f
C240 source.n36 a_n2146_n5888# 0.337966f
C241 source.t19 a_n2146_n5888# 0.723465f
C242 source.t34 a_n2146_n5888# 0.723465f
C243 source.n37 a_n2146_n5888# 4.81328f
C244 source.n38 a_n2146_n5888# 0.337966f
C245 source.t22 a_n2146_n5888# 5.96585f
C246 source.n39 a_n2146_n5888# 0.618094f
C247 source.n40 a_n2146_n5888# 2.57738f
C248 minus.n0 a_n2146_n5888# 0.052939f
C249 minus.t17 a_n2146_n5888# 0.561667f
C250 minus.t9 a_n2146_n5888# 0.55857f
C251 minus.t13 a_n2146_n5888# 0.55857f
C252 minus.n1 a_n2146_n5888# 0.018377f
C253 minus.n2 a_n2146_n5888# 0.052939f
C254 minus.t11 a_n2146_n5888# 0.55857f
C255 minus.n3 a_n2146_n5888# 0.211411f
C256 minus.t14 a_n2146_n5888# 0.55857f
C257 minus.t5 a_n2146_n5888# 0.55857f
C258 minus.t8 a_n2146_n5888# 0.55857f
C259 minus.n4 a_n2146_n5888# 0.211411f
C260 minus.n5 a_n2146_n5888# 0.052939f
C261 minus.t10 a_n2146_n5888# 0.55857f
C262 minus.t3 a_n2146_n5888# 0.55857f
C263 minus.n6 a_n2146_n5888# 0.211411f
C264 minus.t4 a_n2146_n5888# 0.561667f
C265 minus.n7 a_n2146_n5888# 0.233301f
C266 minus.n8 a_n2146_n5888# 0.122115f
C267 minus.n9 a_n2146_n5888# 0.022457f
C268 minus.n10 a_n2146_n5888# 0.211411f
C269 minus.n11 a_n2146_n5888# 0.021641f
C270 minus.n12 a_n2146_n5888# 0.018377f
C271 minus.n13 a_n2146_n5888# 0.052939f
C272 minus.n14 a_n2146_n5888# 0.052939f
C273 minus.n15 a_n2146_n5888# 0.022457f
C274 minus.n16 a_n2146_n5888# 0.211411f
C275 minus.n17 a_n2146_n5888# 0.022457f
C276 minus.n18 a_n2146_n5888# 0.211411f
C277 minus.n19 a_n2146_n5888# 0.022457f
C278 minus.n20 a_n2146_n5888# 0.052939f
C279 minus.n21 a_n2146_n5888# 0.052939f
C280 minus.n22 a_n2146_n5888# 0.052939f
C281 minus.n23 a_n2146_n5888# 0.021641f
C282 minus.n24 a_n2146_n5888# 0.211411f
C283 minus.n25 a_n2146_n5888# 0.022457f
C284 minus.n26 a_n2146_n5888# 0.211411f
C285 minus.n27 a_n2146_n5888# 0.23322f
C286 minus.n28 a_n2146_n5888# 2.77272f
C287 minus.n29 a_n2146_n5888# 0.052939f
C288 minus.t7 a_n2146_n5888# 0.55857f
C289 minus.t1 a_n2146_n5888# 0.55857f
C290 minus.n30 a_n2146_n5888# 0.018377f
C291 minus.n31 a_n2146_n5888# 0.052939f
C292 minus.t15 a_n2146_n5888# 0.55857f
C293 minus.t6 a_n2146_n5888# 0.55857f
C294 minus.t0 a_n2146_n5888# 0.55857f
C295 minus.n32 a_n2146_n5888# 0.211411f
C296 minus.n33 a_n2146_n5888# 0.052939f
C297 minus.t18 a_n2146_n5888# 0.55857f
C298 minus.t12 a_n2146_n5888# 0.55857f
C299 minus.n34 a_n2146_n5888# 0.211411f
C300 minus.t2 a_n2146_n5888# 0.561667f
C301 minus.n35 a_n2146_n5888# 0.233301f
C302 minus.n36 a_n2146_n5888# 0.122115f
C303 minus.n37 a_n2146_n5888# 0.022457f
C304 minus.n38 a_n2146_n5888# 0.211411f
C305 minus.n39 a_n2146_n5888# 0.021641f
C306 minus.n40 a_n2146_n5888# 0.018377f
C307 minus.n41 a_n2146_n5888# 0.052939f
C308 minus.n42 a_n2146_n5888# 0.052939f
C309 minus.n43 a_n2146_n5888# 0.022457f
C310 minus.n44 a_n2146_n5888# 0.211411f
C311 minus.n45 a_n2146_n5888# 0.022457f
C312 minus.n46 a_n2146_n5888# 0.211411f
C313 minus.t19 a_n2146_n5888# 0.55857f
C314 minus.n47 a_n2146_n5888# 0.211411f
C315 minus.n48 a_n2146_n5888# 0.022457f
C316 minus.n49 a_n2146_n5888# 0.052939f
C317 minus.n50 a_n2146_n5888# 0.052939f
C318 minus.n51 a_n2146_n5888# 0.052939f
C319 minus.n52 a_n2146_n5888# 0.021641f
C320 minus.n53 a_n2146_n5888# 0.211411f
C321 minus.n54 a_n2146_n5888# 0.022457f
C322 minus.n55 a_n2146_n5888# 0.211411f
C323 minus.t16 a_n2146_n5888# 0.561667f
C324 minus.n56 a_n2146_n5888# 0.23322f
C325 minus.n57 a_n2146_n5888# 0.353698f
C326 minus.n58 a_n2146_n5888# 3.26351f
.ends

