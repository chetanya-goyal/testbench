* NGSPICE file created from diffpair403.ext - technology: sky130A

.subckt diffpair403 minus drain_right drain_left source plus
X0 source.t14 minus.t0 drain_right.t6 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X1 a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X2 drain_left.t7 plus.t0 source.t4 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X3 a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X4 source.t0 plus.t1 drain_left.t6 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X5 a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X6 drain_left.t5 plus.t2 source.t15 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X7 a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X8 source.t13 minus.t1 drain_right.t5 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X9 drain_right.t4 minus.t2 source.t12 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X10 drain_right.t1 minus.t3 source.t11 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X11 source.t10 minus.t4 drain_right.t0 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X12 source.t2 plus.t3 drain_left.t4 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 source.t1 plus.t4 drain_left.t3 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X14 drain_right.t2 minus.t5 source.t9 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X15 drain_left.t2 plus.t5 source.t5 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X16 source.t8 minus.t6 drain_right.t3 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 source.t6 plus.t6 drain_left.t1 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X18 drain_left.t0 plus.t7 source.t3 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 drain_right.t7 minus.t7 source.t7 a_n1366_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
R0 minus.n5 minus.t4 2206.25
R1 minus.n1 minus.t2 2206.25
R2 minus.n12 minus.t7 2206.25
R3 minus.n8 minus.t0 2206.25
R4 minus.n4 minus.t5 2136.87
R5 minus.n2 minus.t1 2136.87
R6 minus.n11 minus.t6 2136.87
R7 minus.n9 minus.t3 2136.87
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 34.3755
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 drain_right.n5 drain_right.n3 60.1128
R28 drain_right.n2 drain_right.n1 59.7773
R29 drain_right.n2 drain_right.n0 59.7773
R30 drain_right.n5 drain_right.n4 59.5527
R31 drain_right drain_right.n2 28.7751
R32 drain_right drain_right.n5 6.21356
R33 drain_right.n1 drain_right.t3 2.5005
R34 drain_right.n1 drain_right.t7 2.5005
R35 drain_right.n0 drain_right.t6 2.5005
R36 drain_right.n0 drain_right.t1 2.5005
R37 drain_right.n3 drain_right.t5 2.5005
R38 drain_right.n3 drain_right.t4 2.5005
R39 drain_right.n4 drain_right.t0 2.5005
R40 drain_right.n4 drain_right.t2 2.5005
R41 source.n3 source.t1 45.3739
R42 source.n4 source.t12 45.3739
R43 source.n7 source.t10 45.3739
R44 source.n15 source.t7 45.3737
R45 source.n12 source.t14 45.3737
R46 source.n11 source.t15 45.3737
R47 source.n8 source.t0 45.3737
R48 source.n0 source.t5 45.3737
R49 source.n2 source.n1 42.8739
R50 source.n6 source.n5 42.8739
R51 source.n14 source.n13 42.8737
R52 source.n10 source.n9 42.8737
R53 source.n8 source.n7 21.8481
R54 source.n16 source.n0 16.305
R55 source.n16 source.n15 5.5436
R56 source.n13 source.t11 2.5005
R57 source.n13 source.t8 2.5005
R58 source.n9 source.t4 2.5005
R59 source.n9 source.t2 2.5005
R60 source.n1 source.t3 2.5005
R61 source.n1 source.t6 2.5005
R62 source.n5 source.t9 2.5005
R63 source.n5 source.t13 2.5005
R64 source.n7 source.n6 0.560845
R65 source.n6 source.n4 0.560845
R66 source.n3 source.n2 0.560845
R67 source.n2 source.n0 0.560845
R68 source.n10 source.n8 0.560845
R69 source.n11 source.n10 0.560845
R70 source.n14 source.n12 0.560845
R71 source.n15 source.n14 0.560845
R72 source.n4 source.n3 0.470328
R73 source.n12 source.n11 0.470328
R74 source source.n16 0.188
R75 plus.n1 plus.t4 2206.25
R76 plus.n5 plus.t5 2206.25
R77 plus.n8 plus.t2 2206.25
R78 plus.n12 plus.t1 2206.25
R79 plus.n2 plus.t7 2136.87
R80 plus.n4 plus.t6 2136.87
R81 plus.n9 plus.t3 2136.87
R82 plus.n11 plus.t0 2136.87
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus plus.n13 28.2566
R94 plus.n2 plus.n1 25.5611
R95 plus.n5 plus.n4 25.5611
R96 plus.n12 plus.n11 25.5611
R97 plus.n9 plus.n8 25.5611
R98 plus plus.n6 12.224
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 60.113
R102 drain_left.n2 drain_left.n1 59.7773
R103 drain_left.n2 drain_left.n0 59.7773
R104 drain_left.n5 drain_left.n4 59.5525
R105 drain_left drain_left.n2 29.3283
R106 drain_left drain_left.n5 6.21356
R107 drain_left.n1 drain_left.t4 2.5005
R108 drain_left.n1 drain_left.t5 2.5005
R109 drain_left.n0 drain_left.t6 2.5005
R110 drain_left.n0 drain_left.t7 2.5005
R111 drain_left.n4 drain_left.t1 2.5005
R112 drain_left.n4 drain_left.t2 2.5005
R113 drain_left.n3 drain_left.t3 2.5005
R114 drain_left.n3 drain_left.t0 2.5005
C0 drain_right source 16.9029f
C1 drain_right plus 0.282599f
C2 drain_right minus 2.17629f
C3 source drain_left 16.9035f
C4 drain_left plus 2.30568f
C5 drain_left minus 0.170499f
C6 source plus 1.63209f
C7 source minus 1.61805f
C8 minus plus 4.83507f
C9 drain_right drain_left 0.640281f
C10 drain_right a_n1366_n3288# 5.33636f
C11 drain_left a_n1366_n3288# 5.52971f
C12 source a_n1366_n3288# 8.554801f
C13 minus a_n1366_n3288# 4.98574f
C14 plus a_n1366_n3288# 6.74283f
C15 drain_left.t6 a_n1366_n3288# 0.402842f
C16 drain_left.t7 a_n1366_n3288# 0.402842f
C17 drain_left.n0 a_n1366_n3288# 2.64102f
C18 drain_left.t4 a_n1366_n3288# 0.402842f
C19 drain_left.t5 a_n1366_n3288# 0.402842f
C20 drain_left.n1 a_n1366_n3288# 2.64102f
C21 drain_left.n2 a_n1366_n3288# 1.87318f
C22 drain_left.t3 a_n1366_n3288# 0.402842f
C23 drain_left.t0 a_n1366_n3288# 0.402842f
C24 drain_left.n3 a_n1366_n3288# 2.64307f
C25 drain_left.t1 a_n1366_n3288# 0.402842f
C26 drain_left.t2 a_n1366_n3288# 0.402842f
C27 drain_left.n4 a_n1366_n3288# 2.63982f
C28 drain_left.n5 a_n1366_n3288# 0.915299f
C29 plus.n0 a_n1366_n3288# 0.117223f
C30 plus.t6 a_n1366_n3288# 0.251763f
C31 plus.t7 a_n1366_n3288# 0.251763f
C32 plus.t4 a_n1366_n3288# 0.255263f
C33 plus.n1 a_n1366_n3288# 0.128893f
C34 plus.n2 a_n1366_n3288# 0.107502f
C35 plus.n3 a_n1366_n3288# 0.020997f
C36 plus.n4 a_n1366_n3288# 0.107502f
C37 plus.t5 a_n1366_n3288# 0.255263f
C38 plus.n5 a_n1366_n3288# 0.128813f
C39 plus.n6 a_n1366_n3288# 0.563243f
C40 plus.n7 a_n1366_n3288# 0.117223f
C41 plus.t1 a_n1366_n3288# 0.255263f
C42 plus.t0 a_n1366_n3288# 0.251763f
C43 plus.t3 a_n1366_n3288# 0.251763f
C44 plus.t2 a_n1366_n3288# 0.255263f
C45 plus.n8 a_n1366_n3288# 0.128893f
C46 plus.n9 a_n1366_n3288# 0.107502f
C47 plus.n10 a_n1366_n3288# 0.020997f
C48 plus.n11 a_n1366_n3288# 0.107502f
C49 plus.n12 a_n1366_n3288# 0.128813f
C50 plus.n13 a_n1366_n3288# 1.36281f
C51 source.t5 a_n1366_n3288# 2.10233f
C52 source.n0 a_n1366_n3288# 1.04842f
C53 source.t3 a_n1366_n3288# 0.271689f
C54 source.t6 a_n1366_n3288# 0.271689f
C55 source.n1 a_n1366_n3288# 1.72005f
C56 source.n2 a_n1366_n3288# 0.261611f
C57 source.t1 a_n1366_n3288# 2.10234f
C58 source.n3 a_n1366_n3288# 0.362843f
C59 source.t12 a_n1366_n3288# 2.10234f
C60 source.n4 a_n1366_n3288# 0.362843f
C61 source.t9 a_n1366_n3288# 0.271689f
C62 source.t13 a_n1366_n3288# 0.271689f
C63 source.n5 a_n1366_n3288# 1.72005f
C64 source.n6 a_n1366_n3288# 0.261611f
C65 source.t10 a_n1366_n3288# 2.10234f
C66 source.n7 a_n1366_n3288# 1.34612f
C67 source.t0 a_n1366_n3288# 2.10233f
C68 source.n8 a_n1366_n3288# 1.34613f
C69 source.t4 a_n1366_n3288# 0.271689f
C70 source.t2 a_n1366_n3288# 0.271689f
C71 source.n9 a_n1366_n3288# 1.72004f
C72 source.n10 a_n1366_n3288# 0.26162f
C73 source.t15 a_n1366_n3288# 2.10233f
C74 source.n11 a_n1366_n3288# 0.362852f
C75 source.t14 a_n1366_n3288# 2.10233f
C76 source.n12 a_n1366_n3288# 0.362852f
C77 source.t11 a_n1366_n3288# 0.271689f
C78 source.t8 a_n1366_n3288# 0.271689f
C79 source.n13 a_n1366_n3288# 1.72004f
C80 source.n14 a_n1366_n3288# 0.26162f
C81 source.t7 a_n1366_n3288# 2.10233f
C82 source.n15 a_n1366_n3288# 0.470436f
C83 source.n16 a_n1366_n3288# 1.18686f
C84 drain_right.t6 a_n1366_n3288# 0.403047f
C85 drain_right.t1 a_n1366_n3288# 0.403047f
C86 drain_right.n0 a_n1366_n3288# 2.64236f
C87 drain_right.t3 a_n1366_n3288# 0.403047f
C88 drain_right.t7 a_n1366_n3288# 0.403047f
C89 drain_right.n1 a_n1366_n3288# 2.64236f
C90 drain_right.n2 a_n1366_n3288# 1.81542f
C91 drain_right.t5 a_n1366_n3288# 0.403047f
C92 drain_right.t4 a_n1366_n3288# 0.403047f
C93 drain_right.n3 a_n1366_n3288# 2.6444f
C94 drain_right.t0 a_n1366_n3288# 0.403047f
C95 drain_right.t2 a_n1366_n3288# 0.403047f
C96 drain_right.n4 a_n1366_n3288# 2.64117f
C97 drain_right.n5 a_n1366_n3288# 0.915763f
C98 minus.n0 a_n1366_n3288# 0.113966f
C99 minus.t4 a_n1366_n3288# 0.248169f
C100 minus.t5 a_n1366_n3288# 0.244766f
C101 minus.t1 a_n1366_n3288# 0.244766f
C102 minus.t2 a_n1366_n3288# 0.248169f
C103 minus.n1 a_n1366_n3288# 0.125311f
C104 minus.n2 a_n1366_n3288# 0.104515f
C105 minus.n3 a_n1366_n3288# 0.020414f
C106 minus.n4 a_n1366_n3288# 0.104515f
C107 minus.n5 a_n1366_n3288# 0.125233f
C108 minus.n6 a_n1366_n3288# 1.57066f
C109 minus.n7 a_n1366_n3288# 0.113966f
C110 minus.t6 a_n1366_n3288# 0.244766f
C111 minus.t3 a_n1366_n3288# 0.244766f
C112 minus.t0 a_n1366_n3288# 0.248169f
C113 minus.n8 a_n1366_n3288# 0.125311f
C114 minus.n9 a_n1366_n3288# 0.104515f
C115 minus.n10 a_n1366_n3288# 0.020414f
C116 minus.n11 a_n1366_n3288# 0.104515f
C117 minus.t7 a_n1366_n3288# 0.248169f
C118 minus.n12 a_n1366_n3288# 0.125233f
C119 minus.n13 a_n1366_n3288# 0.323643f
C120 minus.n14 a_n1366_n3288# 1.91445f
.ends

