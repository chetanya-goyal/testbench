* NGSPICE file created from diffpair638.ext - technology: sky130A

.subckt diffpair638 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t31 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X2 source.t5 minus.t0 drain_right.t19 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X3 source.t15 minus.t1 drain_right.t18 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X4 source.t29 plus.t1 drain_left.t18 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X5 a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X6 drain_right.t17 minus.t2 source.t16 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X7 drain_right.t16 minus.t3 source.t3 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X8 source.t19 plus.t2 drain_left.t17 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 drain_right.t15 minus.t4 source.t8 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 source.t0 minus.t5 drain_right.t14 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X11 drain_right.t13 minus.t6 source.t11 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 source.t24 plus.t3 drain_left.t16 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X13 drain_right.t12 minus.t7 source.t12 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X14 drain_left.t15 plus.t4 source.t33 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X15 a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X16 drain_left.t14 plus.t5 source.t35 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X17 source.t9 minus.t8 drain_right.t11 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X18 source.t21 plus.t6 drain_left.t13 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X19 drain_right.t10 minus.t9 source.t10 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 drain_right.t9 minus.t10 source.t39 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X21 drain_right.t8 minus.t11 source.t2 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X22 drain_left.t12 plus.t7 source.t30 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X23 source.t36 plus.t8 drain_left.t11 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X24 source.t1 minus.t12 drain_right.t7 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X25 drain_left.t10 plus.t9 source.t32 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X26 source.t38 minus.t13 drain_right.t6 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X27 drain_right.t5 minus.t14 source.t6 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X28 a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X29 drain_right.t4 minus.t15 source.t4 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X30 source.t20 plus.t10 drain_left.t9 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X31 drain_left.t8 plus.t11 source.t23 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X32 drain_left.t7 plus.t12 source.t34 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X33 source.t7 minus.t16 drain_right.t3 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X34 source.t22 plus.t13 drain_left.t6 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X35 drain_left.t5 plus.t14 source.t28 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X36 drain_left.t4 plus.t15 source.t27 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X37 source.t18 plus.t16 drain_left.t3 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X38 drain_left.t2 plus.t17 source.t25 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X39 source.t14 minus.t17 drain_right.t2 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X40 source.t37 minus.t18 drain_right.t1 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X41 source.t17 plus.t18 drain_left.t1 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X42 source.t13 minus.t19 drain_right.t0 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X43 source.t26 plus.t19 drain_left.t0 a_n3202_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n9 plus.t18 673.394
R1 plus.n39 plus.t0 673.394
R2 plus.n28 plus.t5 651.605
R3 plus.n26 plus.t8 651.605
R4 plus.n2 plus.t9 651.605
R5 plus.n21 plus.t10 651.605
R6 plus.n19 plus.t11 651.605
R7 plus.n5 plus.t16 651.605
R8 plus.n13 plus.t12 651.605
R9 plus.n12 plus.t13 651.605
R10 plus.n8 plus.t17 651.605
R11 plus.n58 plus.t19 651.605
R12 plus.n56 plus.t4 651.605
R13 plus.n32 plus.t2 651.605
R14 plus.n51 plus.t7 651.605
R15 plus.n49 plus.t1 651.605
R16 plus.n35 plus.t14 651.605
R17 plus.n43 plus.t3 651.605
R18 plus.n42 plus.t15 651.605
R19 plus.n38 plus.t6 651.605
R20 plus.n11 plus.n10 161.3
R21 plus.n15 plus.n14 161.3
R22 plus.n16 plus.n5 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n4 161.3
R25 plus.n20 plus.n3 161.3
R26 plus.n25 plus.n24 161.3
R27 plus.n26 plus.n1 161.3
R28 plus.n27 plus.n0 161.3
R29 plus.n29 plus.n28 161.3
R30 plus.n41 plus.n40 161.3
R31 plus.n45 plus.n44 161.3
R32 plus.n46 plus.n35 161.3
R33 plus.n48 plus.n47 161.3
R34 plus.n49 plus.n34 161.3
R35 plus.n50 plus.n33 161.3
R36 plus.n55 plus.n54 161.3
R37 plus.n56 plus.n31 161.3
R38 plus.n57 plus.n30 161.3
R39 plus.n59 plus.n58 161.3
R40 plus.n12 plus.n7 80.6037
R41 plus.n13 plus.n6 80.6037
R42 plus.n22 plus.n21 80.6037
R43 plus.n23 plus.n2 80.6037
R44 plus.n42 plus.n37 80.6037
R45 plus.n43 plus.n36 80.6037
R46 plus.n52 plus.n51 80.6037
R47 plus.n53 plus.n32 80.6037
R48 plus.n21 plus.n2 48.2005
R49 plus.n13 plus.n12 48.2005
R50 plus.n51 plus.n32 48.2005
R51 plus.n43 plus.n42 48.2005
R52 plus.n40 plus.n39 44.8565
R53 plus.n10 plus.n9 44.8565
R54 plus.n21 plus.n20 43.0884
R55 plus.n14 plus.n13 43.0884
R56 plus.n51 plus.n50 43.0884
R57 plus.n44 plus.n43 43.0884
R58 plus.n25 plus.n2 40.1672
R59 plus.n12 plus.n11 40.1672
R60 plus.n55 plus.n32 40.1672
R61 plus.n42 plus.n41 40.1672
R62 plus plus.n59 38.3664
R63 plus.n28 plus.n27 27.0217
R64 plus.n58 plus.n57 27.0217
R65 plus.n18 plus.n5 24.1005
R66 plus.n19 plus.n18 24.1005
R67 plus.n49 plus.n48 24.1005
R68 plus.n48 plus.n35 24.1005
R69 plus.n27 plus.n26 21.1793
R70 plus.n57 plus.n56 21.1793
R71 plus.n39 plus.n38 20.1275
R72 plus.n9 plus.n8 20.1275
R73 plus plus.n29 15.3793
R74 plus.n26 plus.n25 8.03383
R75 plus.n11 plus.n8 8.03383
R76 plus.n56 plus.n55 8.03383
R77 plus.n41 plus.n38 8.03383
R78 plus.n20 plus.n19 5.11262
R79 plus.n14 plus.n5 5.11262
R80 plus.n50 plus.n49 5.11262
R81 plus.n44 plus.n35 5.11262
R82 plus.n7 plus.n6 0.380177
R83 plus.n23 plus.n22 0.380177
R84 plus.n53 plus.n52 0.380177
R85 plus.n37 plus.n36 0.380177
R86 plus.n10 plus.n7 0.285035
R87 plus.n15 plus.n6 0.285035
R88 plus.n22 plus.n3 0.285035
R89 plus.n24 plus.n23 0.285035
R90 plus.n54 plus.n53 0.285035
R91 plus.n52 plus.n33 0.285035
R92 plus.n45 plus.n36 0.285035
R93 plus.n40 plus.n37 0.285035
R94 plus.n16 plus.n15 0.189894
R95 plus.n17 plus.n16 0.189894
R96 plus.n17 plus.n4 0.189894
R97 plus.n4 plus.n3 0.189894
R98 plus.n24 plus.n1 0.189894
R99 plus.n1 plus.n0 0.189894
R100 plus.n29 plus.n0 0.189894
R101 plus.n59 plus.n30 0.189894
R102 plus.n31 plus.n30 0.189894
R103 plus.n54 plus.n31 0.189894
R104 plus.n34 plus.n33 0.189894
R105 plus.n47 plus.n34 0.189894
R106 plus.n47 plus.n46 0.189894
R107 plus.n46 plus.n45 0.189894
R108 source.n0 source.t35 44.1297
R109 source.n9 source.t17 44.1296
R110 source.n10 source.t39 44.1296
R111 source.n19 source.t0 44.1296
R112 source.n39 source.t3 44.1295
R113 source.n30 source.t15 44.1295
R114 source.n29 source.t31 44.1295
R115 source.n20 source.t26 44.1295
R116 source.n2 source.n1 43.1397
R117 source.n4 source.n3 43.1397
R118 source.n6 source.n5 43.1397
R119 source.n8 source.n7 43.1397
R120 source.n12 source.n11 43.1397
R121 source.n14 source.n13 43.1397
R122 source.n16 source.n15 43.1397
R123 source.n18 source.n17 43.1397
R124 source.n38 source.n37 43.1396
R125 source.n36 source.n35 43.1396
R126 source.n34 source.n33 43.1396
R127 source.n32 source.n31 43.1396
R128 source.n28 source.n27 43.1396
R129 source.n26 source.n25 43.1396
R130 source.n24 source.n23 43.1396
R131 source.n22 source.n21 43.1396
R132 source.n20 source.n19 28.3225
R133 source.n40 source.n0 22.5725
R134 source.n40 source.n39 5.7505
R135 source.n37 source.t16 0.9905
R136 source.n37 source.t13 0.9905
R137 source.n35 source.t8 0.9905
R138 source.n35 source.t14 0.9905
R139 source.n33 source.t11 0.9905
R140 source.n33 source.t5 0.9905
R141 source.n31 source.t2 0.9905
R142 source.n31 source.t37 0.9905
R143 source.n27 source.t27 0.9905
R144 source.n27 source.t21 0.9905
R145 source.n25 source.t28 0.9905
R146 source.n25 source.t24 0.9905
R147 source.n23 source.t30 0.9905
R148 source.n23 source.t29 0.9905
R149 source.n21 source.t33 0.9905
R150 source.n21 source.t19 0.9905
R151 source.n1 source.t32 0.9905
R152 source.n1 source.t36 0.9905
R153 source.n3 source.t23 0.9905
R154 source.n3 source.t20 0.9905
R155 source.n5 source.t34 0.9905
R156 source.n5 source.t18 0.9905
R157 source.n7 source.t25 0.9905
R158 source.n7 source.t22 0.9905
R159 source.n11 source.t12 0.9905
R160 source.n11 source.t9 0.9905
R161 source.n13 source.t4 0.9905
R162 source.n13 source.t38 0.9905
R163 source.n15 source.t10 0.9905
R164 source.n15 source.t1 0.9905
R165 source.n17 source.t6 0.9905
R166 source.n17 source.t7 0.9905
R167 source.n19 source.n18 0.974638
R168 source.n18 source.n16 0.974638
R169 source.n16 source.n14 0.974638
R170 source.n14 source.n12 0.974638
R171 source.n12 source.n10 0.974638
R172 source.n9 source.n8 0.974638
R173 source.n8 source.n6 0.974638
R174 source.n6 source.n4 0.974638
R175 source.n4 source.n2 0.974638
R176 source.n2 source.n0 0.974638
R177 source.n22 source.n20 0.974638
R178 source.n24 source.n22 0.974638
R179 source.n26 source.n24 0.974638
R180 source.n28 source.n26 0.974638
R181 source.n29 source.n28 0.974638
R182 source.n32 source.n30 0.974638
R183 source.n34 source.n32 0.974638
R184 source.n36 source.n34 0.974638
R185 source.n38 source.n36 0.974638
R186 source.n39 source.n38 0.974638
R187 source.n10 source.n9 0.470328
R188 source.n30 source.n29 0.470328
R189 source source.n40 0.188
R190 drain_left.n10 drain_left.n8 60.7926
R191 drain_left.n6 drain_left.n4 60.7925
R192 drain_left.n2 drain_left.n0 60.7925
R193 drain_left.n16 drain_left.n15 59.8185
R194 drain_left.n14 drain_left.n13 59.8185
R195 drain_left.n12 drain_left.n11 59.8185
R196 drain_left.n10 drain_left.n9 59.8185
R197 drain_left.n7 drain_left.n3 59.8184
R198 drain_left.n6 drain_left.n5 59.8184
R199 drain_left.n2 drain_left.n1 59.8184
R200 drain_left drain_left.n7 41.2208
R201 drain_left drain_left.n16 6.62735
R202 drain_left.n3 drain_left.t18 0.9905
R203 drain_left.n3 drain_left.t5 0.9905
R204 drain_left.n4 drain_left.t13 0.9905
R205 drain_left.n4 drain_left.t19 0.9905
R206 drain_left.n5 drain_left.t16 0.9905
R207 drain_left.n5 drain_left.t4 0.9905
R208 drain_left.n1 drain_left.t17 0.9905
R209 drain_left.n1 drain_left.t12 0.9905
R210 drain_left.n0 drain_left.t0 0.9905
R211 drain_left.n0 drain_left.t15 0.9905
R212 drain_left.n15 drain_left.t11 0.9905
R213 drain_left.n15 drain_left.t14 0.9905
R214 drain_left.n13 drain_left.t9 0.9905
R215 drain_left.n13 drain_left.t10 0.9905
R216 drain_left.n11 drain_left.t3 0.9905
R217 drain_left.n11 drain_left.t8 0.9905
R218 drain_left.n9 drain_left.t6 0.9905
R219 drain_left.n9 drain_left.t7 0.9905
R220 drain_left.n8 drain_left.t1 0.9905
R221 drain_left.n8 drain_left.t2 0.9905
R222 drain_left.n12 drain_left.n10 0.974638
R223 drain_left.n14 drain_left.n12 0.974638
R224 drain_left.n16 drain_left.n14 0.974638
R225 drain_left.n7 drain_left.n6 0.919292
R226 drain_left.n7 drain_left.n2 0.919292
R227 minus.n7 minus.t10 673.394
R228 minus.n37 minus.t1 673.394
R229 minus.n8 minus.t8 651.605
R230 minus.n10 minus.t7 651.605
R231 minus.n5 minus.t13 651.605
R232 minus.n15 minus.t15 651.605
R233 minus.n3 minus.t12 651.605
R234 minus.n21 minus.t9 651.605
R235 minus.n22 minus.t16 651.605
R236 minus.n26 minus.t14 651.605
R237 minus.n28 minus.t5 651.605
R238 minus.n38 minus.t11 651.605
R239 minus.n40 minus.t18 651.605
R240 minus.n35 minus.t6 651.605
R241 minus.n45 minus.t0 651.605
R242 minus.n33 minus.t4 651.605
R243 minus.n51 minus.t17 651.605
R244 minus.n52 minus.t2 651.605
R245 minus.n56 minus.t19 651.605
R246 minus.n58 minus.t3 651.605
R247 minus.n29 minus.n28 161.3
R248 minus.n27 minus.n0 161.3
R249 minus.n26 minus.n25 161.3
R250 minus.n24 minus.n1 161.3
R251 minus.n20 minus.n19 161.3
R252 minus.n18 minus.n3 161.3
R253 minus.n17 minus.n16 161.3
R254 minus.n15 minus.n4 161.3
R255 minus.n14 minus.n13 161.3
R256 minus.n9 minus.n6 161.3
R257 minus.n59 minus.n58 161.3
R258 minus.n57 minus.n30 161.3
R259 minus.n56 minus.n55 161.3
R260 minus.n54 minus.n31 161.3
R261 minus.n50 minus.n49 161.3
R262 minus.n48 minus.n33 161.3
R263 minus.n47 minus.n46 161.3
R264 minus.n45 minus.n34 161.3
R265 minus.n44 minus.n43 161.3
R266 minus.n39 minus.n36 161.3
R267 minus.n23 minus.n22 80.6037
R268 minus.n21 minus.n2 80.6037
R269 minus.n12 minus.n5 80.6037
R270 minus.n11 minus.n10 80.6037
R271 minus.n53 minus.n52 80.6037
R272 minus.n51 minus.n32 80.6037
R273 minus.n42 minus.n35 80.6037
R274 minus.n41 minus.n40 80.6037
R275 minus.n10 minus.n5 48.2005
R276 minus.n22 minus.n21 48.2005
R277 minus.n40 minus.n35 48.2005
R278 minus.n52 minus.n51 48.2005
R279 minus.n60 minus.n29 47.5156
R280 minus.n7 minus.n6 44.8565
R281 minus.n37 minus.n36 44.8565
R282 minus.n14 minus.n5 43.0884
R283 minus.n21 minus.n20 43.0884
R284 minus.n44 minus.n35 43.0884
R285 minus.n51 minus.n50 43.0884
R286 minus.n10 minus.n9 40.1672
R287 minus.n22 minus.n1 40.1672
R288 minus.n40 minus.n39 40.1672
R289 minus.n52 minus.n31 40.1672
R290 minus.n28 minus.n27 27.0217
R291 minus.n58 minus.n57 27.0217
R292 minus.n16 minus.n3 24.1005
R293 minus.n16 minus.n15 24.1005
R294 minus.n46 minus.n45 24.1005
R295 minus.n46 minus.n33 24.1005
R296 minus.n27 minus.n26 21.1793
R297 minus.n57 minus.n56 21.1793
R298 minus.n8 minus.n7 20.1275
R299 minus.n38 minus.n37 20.1275
R300 minus.n9 minus.n8 8.03383
R301 minus.n26 minus.n1 8.03383
R302 minus.n39 minus.n38 8.03383
R303 minus.n56 minus.n31 8.03383
R304 minus.n60 minus.n59 6.70505
R305 minus.n15 minus.n14 5.11262
R306 minus.n20 minus.n3 5.11262
R307 minus.n45 minus.n44 5.11262
R308 minus.n50 minus.n33 5.11262
R309 minus.n23 minus.n2 0.380177
R310 minus.n12 minus.n11 0.380177
R311 minus.n42 minus.n41 0.380177
R312 minus.n53 minus.n32 0.380177
R313 minus.n24 minus.n23 0.285035
R314 minus.n19 minus.n2 0.285035
R315 minus.n13 minus.n12 0.285035
R316 minus.n11 minus.n6 0.285035
R317 minus.n41 minus.n36 0.285035
R318 minus.n43 minus.n42 0.285035
R319 minus.n49 minus.n32 0.285035
R320 minus.n54 minus.n53 0.285035
R321 minus.n29 minus.n0 0.189894
R322 minus.n25 minus.n0 0.189894
R323 minus.n25 minus.n24 0.189894
R324 minus.n19 minus.n18 0.189894
R325 minus.n18 minus.n17 0.189894
R326 minus.n17 minus.n4 0.189894
R327 minus.n13 minus.n4 0.189894
R328 minus.n43 minus.n34 0.189894
R329 minus.n47 minus.n34 0.189894
R330 minus.n48 minus.n47 0.189894
R331 minus.n49 minus.n48 0.189894
R332 minus.n55 minus.n54 0.189894
R333 minus.n55 minus.n30 0.189894
R334 minus.n59 minus.n30 0.189894
R335 minus minus.n60 0.188
R336 drain_right.n10 drain_right.n8 60.7926
R337 drain_right.n6 drain_right.n4 60.7925
R338 drain_right.n2 drain_right.n0 60.7925
R339 drain_right.n10 drain_right.n9 59.8185
R340 drain_right.n12 drain_right.n11 59.8185
R341 drain_right.n14 drain_right.n13 59.8185
R342 drain_right.n16 drain_right.n15 59.8185
R343 drain_right.n7 drain_right.n3 59.8184
R344 drain_right.n6 drain_right.n5 59.8184
R345 drain_right.n2 drain_right.n1 59.8184
R346 drain_right drain_right.n7 40.6676
R347 drain_right drain_right.n16 6.62735
R348 drain_right.n3 drain_right.t19 0.9905
R349 drain_right.n3 drain_right.t15 0.9905
R350 drain_right.n4 drain_right.t0 0.9905
R351 drain_right.n4 drain_right.t16 0.9905
R352 drain_right.n5 drain_right.t2 0.9905
R353 drain_right.n5 drain_right.t17 0.9905
R354 drain_right.n1 drain_right.t1 0.9905
R355 drain_right.n1 drain_right.t13 0.9905
R356 drain_right.n0 drain_right.t18 0.9905
R357 drain_right.n0 drain_right.t8 0.9905
R358 drain_right.n8 drain_right.t11 0.9905
R359 drain_right.n8 drain_right.t9 0.9905
R360 drain_right.n9 drain_right.t6 0.9905
R361 drain_right.n9 drain_right.t12 0.9905
R362 drain_right.n11 drain_right.t7 0.9905
R363 drain_right.n11 drain_right.t4 0.9905
R364 drain_right.n13 drain_right.t3 0.9905
R365 drain_right.n13 drain_right.t10 0.9905
R366 drain_right.n15 drain_right.t14 0.9905
R367 drain_right.n15 drain_right.t5 0.9905
R368 drain_right.n16 drain_right.n14 0.974638
R369 drain_right.n14 drain_right.n12 0.974638
R370 drain_right.n12 drain_right.n10 0.974638
R371 drain_right.n7 drain_right.n6 0.919292
R372 drain_right.n7 drain_right.n2 0.919292
C0 plus drain_left 22.4149f
C1 drain_left minus 0.17405f
C2 plus drain_right 0.478206f
C3 drain_right minus 22.0945f
C4 drain_right drain_left 1.72917f
C5 source plus 22.0403f
C6 source minus 22.0262f
C7 source drain_left 34.6014f
C8 source drain_right 34.6042f
C9 plus minus 8.61978f
C10 drain_right a_n3202_n4888# 8.93872f
C11 drain_left a_n3202_n4888# 9.37817f
C12 source a_n3202_n4888# 14.065453f
C13 minus a_n3202_n4888# 13.474322f
C14 plus a_n3202_n4888# 15.60424f
C15 drain_right.t18 a_n3202_n4888# 0.418953f
C16 drain_right.t8 a_n3202_n4888# 0.418953f
C17 drain_right.n0 a_n3202_n4888# 3.83659f
C18 drain_right.t1 a_n3202_n4888# 0.418953f
C19 drain_right.t13 a_n3202_n4888# 0.418953f
C20 drain_right.n1 a_n3202_n4888# 3.83016f
C21 drain_right.n2 a_n3202_n4888# 0.780407f
C22 drain_right.t19 a_n3202_n4888# 0.418953f
C23 drain_right.t15 a_n3202_n4888# 0.418953f
C24 drain_right.n3 a_n3202_n4888# 3.83016f
C25 drain_right.t0 a_n3202_n4888# 0.418953f
C26 drain_right.t16 a_n3202_n4888# 0.418953f
C27 drain_right.n4 a_n3202_n4888# 3.83659f
C28 drain_right.t2 a_n3202_n4888# 0.418953f
C29 drain_right.t17 a_n3202_n4888# 0.418953f
C30 drain_right.n5 a_n3202_n4888# 3.83016f
C31 drain_right.n6 a_n3202_n4888# 0.780407f
C32 drain_right.n7 a_n3202_n4888# 2.47721f
C33 drain_right.t11 a_n3202_n4888# 0.418953f
C34 drain_right.t9 a_n3202_n4888# 0.418953f
C35 drain_right.n8 a_n3202_n4888# 3.83658f
C36 drain_right.t6 a_n3202_n4888# 0.418953f
C37 drain_right.t12 a_n3202_n4888# 0.418953f
C38 drain_right.n9 a_n3202_n4888# 3.83016f
C39 drain_right.n10 a_n3202_n4888# 0.784477f
C40 drain_right.t7 a_n3202_n4888# 0.418953f
C41 drain_right.t4 a_n3202_n4888# 0.418953f
C42 drain_right.n11 a_n3202_n4888# 3.83016f
C43 drain_right.n12 a_n3202_n4888# 0.390111f
C44 drain_right.t3 a_n3202_n4888# 0.418953f
C45 drain_right.t10 a_n3202_n4888# 0.418953f
C46 drain_right.n13 a_n3202_n4888# 3.83016f
C47 drain_right.n14 a_n3202_n4888# 0.390111f
C48 drain_right.t14 a_n3202_n4888# 0.418953f
C49 drain_right.t5 a_n3202_n4888# 0.418953f
C50 drain_right.n15 a_n3202_n4888# 3.83016f
C51 drain_right.n16 a_n3202_n4888# 0.627809f
C52 minus.n0 a_n3202_n4888# 0.037343f
C53 minus.n1 a_n3202_n4888# 0.008474f
C54 minus.t14 a_n3202_n4888# 1.69202f
C55 minus.n2 a_n3202_n4888# 0.062199f
C56 minus.t12 a_n3202_n4888# 1.69202f
C57 minus.n3 a_n3202_n4888# 0.627536f
C58 minus.n4 a_n3202_n4888# 0.037343f
C59 minus.t13 a_n3202_n4888# 1.69202f
C60 minus.n5 a_n3202_n4888# 0.638197f
C61 minus.n6 a_n3202_n4888# 0.171889f
C62 minus.t10 a_n3202_n4888# 1.7124f
C63 minus.n7 a_n3202_n4888# 0.612942f
C64 minus.t8 a_n3202_n4888# 1.69202f
C65 minus.n8 a_n3202_n4888# 0.630674f
C66 minus.n9 a_n3202_n4888# 0.008474f
C67 minus.t7 a_n3202_n4888# 1.69202f
C68 minus.n10 a_n3202_n4888# 0.637736f
C69 minus.n11 a_n3202_n4888# 0.062199f
C70 minus.n12 a_n3202_n4888# 0.062199f
C71 minus.n13 a_n3202_n4888# 0.049829f
C72 minus.n14 a_n3202_n4888# 0.008474f
C73 minus.t15 a_n3202_n4888# 1.69202f
C74 minus.n15 a_n3202_n4888# 0.627536f
C75 minus.n16 a_n3202_n4888# 0.008474f
C76 minus.n17 a_n3202_n4888# 0.037343f
C77 minus.n18 a_n3202_n4888# 0.037343f
C78 minus.n19 a_n3202_n4888# 0.049829f
C79 minus.n20 a_n3202_n4888# 0.008474f
C80 minus.t9 a_n3202_n4888# 1.69202f
C81 minus.n21 a_n3202_n4888# 0.638197f
C82 minus.t16 a_n3202_n4888# 1.69202f
C83 minus.n22 a_n3202_n4888# 0.637736f
C84 minus.n23 a_n3202_n4888# 0.062199f
C85 minus.n24 a_n3202_n4888# 0.049829f
C86 minus.n25 a_n3202_n4888# 0.037343f
C87 minus.n26 a_n3202_n4888# 0.627536f
C88 minus.n27 a_n3202_n4888# 0.008474f
C89 minus.t5 a_n3202_n4888# 1.69202f
C90 minus.n28 a_n3202_n4888# 0.62719f
C91 minus.n29 a_n3202_n4888# 1.97989f
C92 minus.n30 a_n3202_n4888# 0.037343f
C93 minus.n31 a_n3202_n4888# 0.008474f
C94 minus.n32 a_n3202_n4888# 0.062199f
C95 minus.t4 a_n3202_n4888# 1.69202f
C96 minus.n33 a_n3202_n4888# 0.627536f
C97 minus.n34 a_n3202_n4888# 0.037343f
C98 minus.t6 a_n3202_n4888# 1.69202f
C99 minus.n35 a_n3202_n4888# 0.638197f
C100 minus.n36 a_n3202_n4888# 0.171889f
C101 minus.t1 a_n3202_n4888# 1.7124f
C102 minus.n37 a_n3202_n4888# 0.612942f
C103 minus.t11 a_n3202_n4888# 1.69202f
C104 minus.n38 a_n3202_n4888# 0.630674f
C105 minus.n39 a_n3202_n4888# 0.008474f
C106 minus.t18 a_n3202_n4888# 1.69202f
C107 minus.n40 a_n3202_n4888# 0.637736f
C108 minus.n41 a_n3202_n4888# 0.062199f
C109 minus.n42 a_n3202_n4888# 0.062199f
C110 minus.n43 a_n3202_n4888# 0.049829f
C111 minus.n44 a_n3202_n4888# 0.008474f
C112 minus.t0 a_n3202_n4888# 1.69202f
C113 minus.n45 a_n3202_n4888# 0.627536f
C114 minus.n46 a_n3202_n4888# 0.008474f
C115 minus.n47 a_n3202_n4888# 0.037343f
C116 minus.n48 a_n3202_n4888# 0.037343f
C117 minus.n49 a_n3202_n4888# 0.049829f
C118 minus.n50 a_n3202_n4888# 0.008474f
C119 minus.t17 a_n3202_n4888# 1.69202f
C120 minus.n51 a_n3202_n4888# 0.638197f
C121 minus.t2 a_n3202_n4888# 1.69202f
C122 minus.n52 a_n3202_n4888# 0.637736f
C123 minus.n53 a_n3202_n4888# 0.062199f
C124 minus.n54 a_n3202_n4888# 0.049829f
C125 minus.n55 a_n3202_n4888# 0.037343f
C126 minus.t19 a_n3202_n4888# 1.69202f
C127 minus.n56 a_n3202_n4888# 0.627536f
C128 minus.n57 a_n3202_n4888# 0.008474f
C129 minus.t3 a_n3202_n4888# 1.69202f
C130 minus.n58 a_n3202_n4888# 0.62719f
C131 minus.n59 a_n3202_n4888# 0.262007f
C132 minus.n60 a_n3202_n4888# 2.32636f
C133 drain_left.t0 a_n3202_n4888# 0.420401f
C134 drain_left.t15 a_n3202_n4888# 0.420401f
C135 drain_left.n0 a_n3202_n4888# 3.84984f
C136 drain_left.t17 a_n3202_n4888# 0.420401f
C137 drain_left.t12 a_n3202_n4888# 0.420401f
C138 drain_left.n1 a_n3202_n4888# 3.8434f
C139 drain_left.n2 a_n3202_n4888# 0.783104f
C140 drain_left.t18 a_n3202_n4888# 0.420401f
C141 drain_left.t5 a_n3202_n4888# 0.420401f
C142 drain_left.n3 a_n3202_n4888# 3.8434f
C143 drain_left.t13 a_n3202_n4888# 0.420401f
C144 drain_left.t19 a_n3202_n4888# 0.420401f
C145 drain_left.n4 a_n3202_n4888# 3.84984f
C146 drain_left.t16 a_n3202_n4888# 0.420401f
C147 drain_left.t4 a_n3202_n4888# 0.420401f
C148 drain_left.n5 a_n3202_n4888# 3.8434f
C149 drain_left.n6 a_n3202_n4888# 0.783104f
C150 drain_left.n7 a_n3202_n4888# 2.54013f
C151 drain_left.t1 a_n3202_n4888# 0.420401f
C152 drain_left.t2 a_n3202_n4888# 0.420401f
C153 drain_left.n8 a_n3202_n4888# 3.84984f
C154 drain_left.t6 a_n3202_n4888# 0.420401f
C155 drain_left.t7 a_n3202_n4888# 0.420401f
C156 drain_left.n9 a_n3202_n4888# 3.8434f
C157 drain_left.n10 a_n3202_n4888# 0.787188f
C158 drain_left.t3 a_n3202_n4888# 0.420401f
C159 drain_left.t8 a_n3202_n4888# 0.420401f
C160 drain_left.n11 a_n3202_n4888# 3.8434f
C161 drain_left.n12 a_n3202_n4888# 0.391459f
C162 drain_left.t9 a_n3202_n4888# 0.420401f
C163 drain_left.t10 a_n3202_n4888# 0.420401f
C164 drain_left.n13 a_n3202_n4888# 3.8434f
C165 drain_left.n14 a_n3202_n4888# 0.391459f
C166 drain_left.t11 a_n3202_n4888# 0.420401f
C167 drain_left.t14 a_n3202_n4888# 0.420401f
C168 drain_left.n15 a_n3202_n4888# 3.8434f
C169 drain_left.n16 a_n3202_n4888# 0.629979f
C170 source.t35 a_n3202_n4888# 4.13662f
C171 source.n0 a_n3202_n4888# 1.80956f
C172 source.t32 a_n3202_n4888# 0.36196f
C173 source.t36 a_n3202_n4888# 0.36196f
C174 source.n1 a_n3202_n4888# 3.23608f
C175 source.n2 a_n3202_n4888# 0.378949f
C176 source.t23 a_n3202_n4888# 0.36196f
C177 source.t20 a_n3202_n4888# 0.36196f
C178 source.n3 a_n3202_n4888# 3.23608f
C179 source.n4 a_n3202_n4888# 0.378949f
C180 source.t34 a_n3202_n4888# 0.36196f
C181 source.t18 a_n3202_n4888# 0.36196f
C182 source.n5 a_n3202_n4888# 3.23608f
C183 source.n6 a_n3202_n4888# 0.378949f
C184 source.t25 a_n3202_n4888# 0.36196f
C185 source.t22 a_n3202_n4888# 0.36196f
C186 source.n7 a_n3202_n4888# 3.23608f
C187 source.n8 a_n3202_n4888# 0.378949f
C188 source.t17 a_n3202_n4888# 4.13662f
C189 source.n9 a_n3202_n4888# 0.428348f
C190 source.t39 a_n3202_n4888# 4.13662f
C191 source.n10 a_n3202_n4888# 0.428348f
C192 source.t12 a_n3202_n4888# 0.36196f
C193 source.t9 a_n3202_n4888# 0.36196f
C194 source.n11 a_n3202_n4888# 3.23608f
C195 source.n12 a_n3202_n4888# 0.378949f
C196 source.t4 a_n3202_n4888# 0.36196f
C197 source.t38 a_n3202_n4888# 0.36196f
C198 source.n13 a_n3202_n4888# 3.23608f
C199 source.n14 a_n3202_n4888# 0.378949f
C200 source.t10 a_n3202_n4888# 0.36196f
C201 source.t1 a_n3202_n4888# 0.36196f
C202 source.n15 a_n3202_n4888# 3.23608f
C203 source.n16 a_n3202_n4888# 0.378949f
C204 source.t6 a_n3202_n4888# 0.36196f
C205 source.t7 a_n3202_n4888# 0.36196f
C206 source.n17 a_n3202_n4888# 3.23608f
C207 source.n18 a_n3202_n4888# 0.378949f
C208 source.t0 a_n3202_n4888# 4.13662f
C209 source.n19 a_n3202_n4888# 2.22891f
C210 source.t26 a_n3202_n4888# 4.1366f
C211 source.n20 a_n3202_n4888# 2.22894f
C212 source.t33 a_n3202_n4888# 0.36196f
C213 source.t19 a_n3202_n4888# 0.36196f
C214 source.n21 a_n3202_n4888# 3.23608f
C215 source.n22 a_n3202_n4888# 0.378942f
C216 source.t30 a_n3202_n4888# 0.36196f
C217 source.t29 a_n3202_n4888# 0.36196f
C218 source.n23 a_n3202_n4888# 3.23608f
C219 source.n24 a_n3202_n4888# 0.378942f
C220 source.t28 a_n3202_n4888# 0.36196f
C221 source.t24 a_n3202_n4888# 0.36196f
C222 source.n25 a_n3202_n4888# 3.23608f
C223 source.n26 a_n3202_n4888# 0.378942f
C224 source.t27 a_n3202_n4888# 0.36196f
C225 source.t21 a_n3202_n4888# 0.36196f
C226 source.n27 a_n3202_n4888# 3.23608f
C227 source.n28 a_n3202_n4888# 0.378942f
C228 source.t31 a_n3202_n4888# 4.1366f
C229 source.n29 a_n3202_n4888# 0.428371f
C230 source.t15 a_n3202_n4888# 4.1366f
C231 source.n30 a_n3202_n4888# 0.428371f
C232 source.t2 a_n3202_n4888# 0.36196f
C233 source.t37 a_n3202_n4888# 0.36196f
C234 source.n31 a_n3202_n4888# 3.23608f
C235 source.n32 a_n3202_n4888# 0.378942f
C236 source.t11 a_n3202_n4888# 0.36196f
C237 source.t5 a_n3202_n4888# 0.36196f
C238 source.n33 a_n3202_n4888# 3.23608f
C239 source.n34 a_n3202_n4888# 0.378942f
C240 source.t8 a_n3202_n4888# 0.36196f
C241 source.t14 a_n3202_n4888# 0.36196f
C242 source.n35 a_n3202_n4888# 3.23608f
C243 source.n36 a_n3202_n4888# 0.378942f
C244 source.t16 a_n3202_n4888# 0.36196f
C245 source.t13 a_n3202_n4888# 0.36196f
C246 source.n37 a_n3202_n4888# 3.23608f
C247 source.n38 a_n3202_n4888# 0.378942f
C248 source.t3 a_n3202_n4888# 4.1366f
C249 source.n39 a_n3202_n4888# 0.582721f
C250 source.n40 a_n3202_n4888# 2.08186f
C251 plus.n0 a_n3202_n4888# 0.037609f
C252 plus.t5 a_n3202_n4888# 1.7041f
C253 plus.t8 a_n3202_n4888# 1.7041f
C254 plus.n1 a_n3202_n4888# 0.037609f
C255 plus.t9 a_n3202_n4888# 1.7041f
C256 plus.n2 a_n3202_n4888# 0.642287f
C257 plus.n3 a_n3202_n4888# 0.050185f
C258 plus.t10 a_n3202_n4888# 1.7041f
C259 plus.t11 a_n3202_n4888# 1.7041f
C260 plus.n4 a_n3202_n4888# 0.037609f
C261 plus.t16 a_n3202_n4888# 1.7041f
C262 plus.n5 a_n3202_n4888# 0.632014f
C263 plus.n6 a_n3202_n4888# 0.062643f
C264 plus.t12 a_n3202_n4888# 1.7041f
C265 plus.t13 a_n3202_n4888# 1.7041f
C266 plus.n7 a_n3202_n4888# 0.062643f
C267 plus.t17 a_n3202_n4888# 1.7041f
C268 plus.n8 a_n3202_n4888# 0.635175f
C269 plus.t18 a_n3202_n4888# 1.72462f
C270 plus.n9 a_n3202_n4888# 0.617316f
C271 plus.n10 a_n3202_n4888# 0.173115f
C272 plus.n11 a_n3202_n4888# 0.008534f
C273 plus.n12 a_n3202_n4888# 0.642287f
C274 plus.n13 a_n3202_n4888# 0.642751f
C275 plus.n14 a_n3202_n4888# 0.008534f
C276 plus.n15 a_n3202_n4888# 0.050185f
C277 plus.n16 a_n3202_n4888# 0.037609f
C278 plus.n17 a_n3202_n4888# 0.037609f
C279 plus.n18 a_n3202_n4888# 0.008534f
C280 plus.n19 a_n3202_n4888# 0.632014f
C281 plus.n20 a_n3202_n4888# 0.008534f
C282 plus.n21 a_n3202_n4888# 0.642751f
C283 plus.n22 a_n3202_n4888# 0.062643f
C284 plus.n23 a_n3202_n4888# 0.062643f
C285 plus.n24 a_n3202_n4888# 0.050185f
C286 plus.n25 a_n3202_n4888# 0.008534f
C287 plus.n26 a_n3202_n4888# 0.632014f
C288 plus.n27 a_n3202_n4888# 0.008534f
C289 plus.n28 a_n3202_n4888# 0.631666f
C290 plus.n29 a_n3202_n4888# 0.588744f
C291 plus.n30 a_n3202_n4888# 0.037609f
C292 plus.t19 a_n3202_n4888# 1.7041f
C293 plus.n31 a_n3202_n4888# 0.037609f
C294 plus.t4 a_n3202_n4888# 1.7041f
C295 plus.t2 a_n3202_n4888# 1.7041f
C296 plus.n32 a_n3202_n4888# 0.642287f
C297 plus.n33 a_n3202_n4888# 0.050185f
C298 plus.t7 a_n3202_n4888# 1.7041f
C299 plus.n34 a_n3202_n4888# 0.037609f
C300 plus.t1 a_n3202_n4888# 1.7041f
C301 plus.t14 a_n3202_n4888# 1.7041f
C302 plus.n35 a_n3202_n4888# 0.632014f
C303 plus.n36 a_n3202_n4888# 0.062643f
C304 plus.t3 a_n3202_n4888# 1.7041f
C305 plus.n37 a_n3202_n4888# 0.062643f
C306 plus.t15 a_n3202_n4888# 1.7041f
C307 plus.t6 a_n3202_n4888# 1.7041f
C308 plus.n38 a_n3202_n4888# 0.635175f
C309 plus.t0 a_n3202_n4888# 1.72462f
C310 plus.n39 a_n3202_n4888# 0.617316f
C311 plus.n40 a_n3202_n4888# 0.173115f
C312 plus.n41 a_n3202_n4888# 0.008534f
C313 plus.n42 a_n3202_n4888# 0.642287f
C314 plus.n43 a_n3202_n4888# 0.642751f
C315 plus.n44 a_n3202_n4888# 0.008534f
C316 plus.n45 a_n3202_n4888# 0.050185f
C317 plus.n46 a_n3202_n4888# 0.037609f
C318 plus.n47 a_n3202_n4888# 0.037609f
C319 plus.n48 a_n3202_n4888# 0.008534f
C320 plus.n49 a_n3202_n4888# 0.632014f
C321 plus.n50 a_n3202_n4888# 0.008534f
C322 plus.n51 a_n3202_n4888# 0.642751f
C323 plus.n52 a_n3202_n4888# 0.062643f
C324 plus.n53 a_n3202_n4888# 0.062643f
C325 plus.n54 a_n3202_n4888# 0.050185f
C326 plus.n55 a_n3202_n4888# 0.008534f
C327 plus.n56 a_n3202_n4888# 0.632014f
C328 plus.n57 a_n3202_n4888# 0.008534f
C329 plus.n58 a_n3202_n4888# 0.631666f
C330 plus.n59 a_n3202_n4888# 1.61241f
.ends

