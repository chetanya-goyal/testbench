* NGSPICE file created from diffpair671.ext - technology: sky130A

.subckt diffpair671 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t6 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X1 source.t3 plus.t0 drain_left.t3 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X2 drain_right.t2 minus.t1 source.t4 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X3 source.t5 minus.t2 drain_right.t1 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X4 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X5 drain_left.t2 plus.t1 source.t0 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X6 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X7 source.t7 minus.t3 drain_right.t0 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X8 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X9 source.t1 plus.t2 drain_left.t1 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X10 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X11 drain_left.t0 plus.t3 source.t2 a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
R0 minus.n0 minus.t2 2158.78
R1 minus.n0 minus.t0 2158.78
R2 minus.n1 minus.t1 2158.78
R3 minus.n1 minus.t3 2158.78
R4 minus.n2 minus.n0 204.436
R5 minus.n2 minus.n1 167.809
R6 minus minus.n2 0.188
R7 source.n1114 source.n980 289.615
R8 source.n974 source.n840 289.615
R9 source.n834 source.n700 289.615
R10 source.n694 source.n560 289.615
R11 source.n134 source.n0 289.615
R12 source.n274 source.n140 289.615
R13 source.n414 source.n280 289.615
R14 source.n554 source.n420 289.615
R15 source.n1024 source.n1023 185
R16 source.n1029 source.n1028 185
R17 source.n1031 source.n1030 185
R18 source.n1020 source.n1019 185
R19 source.n1037 source.n1036 185
R20 source.n1039 source.n1038 185
R21 source.n1016 source.n1015 185
R22 source.n1046 source.n1045 185
R23 source.n1047 source.n1014 185
R24 source.n1049 source.n1048 185
R25 source.n1012 source.n1011 185
R26 source.n1055 source.n1054 185
R27 source.n1057 source.n1056 185
R28 source.n1008 source.n1007 185
R29 source.n1063 source.n1062 185
R30 source.n1065 source.n1064 185
R31 source.n1004 source.n1003 185
R32 source.n1071 source.n1070 185
R33 source.n1073 source.n1072 185
R34 source.n1000 source.n999 185
R35 source.n1079 source.n1078 185
R36 source.n1081 source.n1080 185
R37 source.n996 source.n995 185
R38 source.n1087 source.n1086 185
R39 source.n1090 source.n1089 185
R40 source.n1088 source.n992 185
R41 source.n1095 source.n991 185
R42 source.n1097 source.n1096 185
R43 source.n1099 source.n1098 185
R44 source.n988 source.n987 185
R45 source.n1105 source.n1104 185
R46 source.n1107 source.n1106 185
R47 source.n984 source.n983 185
R48 source.n1113 source.n1112 185
R49 source.n1115 source.n1114 185
R50 source.n884 source.n883 185
R51 source.n889 source.n888 185
R52 source.n891 source.n890 185
R53 source.n880 source.n879 185
R54 source.n897 source.n896 185
R55 source.n899 source.n898 185
R56 source.n876 source.n875 185
R57 source.n906 source.n905 185
R58 source.n907 source.n874 185
R59 source.n909 source.n908 185
R60 source.n872 source.n871 185
R61 source.n915 source.n914 185
R62 source.n917 source.n916 185
R63 source.n868 source.n867 185
R64 source.n923 source.n922 185
R65 source.n925 source.n924 185
R66 source.n864 source.n863 185
R67 source.n931 source.n930 185
R68 source.n933 source.n932 185
R69 source.n860 source.n859 185
R70 source.n939 source.n938 185
R71 source.n941 source.n940 185
R72 source.n856 source.n855 185
R73 source.n947 source.n946 185
R74 source.n950 source.n949 185
R75 source.n948 source.n852 185
R76 source.n955 source.n851 185
R77 source.n957 source.n956 185
R78 source.n959 source.n958 185
R79 source.n848 source.n847 185
R80 source.n965 source.n964 185
R81 source.n967 source.n966 185
R82 source.n844 source.n843 185
R83 source.n973 source.n972 185
R84 source.n975 source.n974 185
R85 source.n744 source.n743 185
R86 source.n749 source.n748 185
R87 source.n751 source.n750 185
R88 source.n740 source.n739 185
R89 source.n757 source.n756 185
R90 source.n759 source.n758 185
R91 source.n736 source.n735 185
R92 source.n766 source.n765 185
R93 source.n767 source.n734 185
R94 source.n769 source.n768 185
R95 source.n732 source.n731 185
R96 source.n775 source.n774 185
R97 source.n777 source.n776 185
R98 source.n728 source.n727 185
R99 source.n783 source.n782 185
R100 source.n785 source.n784 185
R101 source.n724 source.n723 185
R102 source.n791 source.n790 185
R103 source.n793 source.n792 185
R104 source.n720 source.n719 185
R105 source.n799 source.n798 185
R106 source.n801 source.n800 185
R107 source.n716 source.n715 185
R108 source.n807 source.n806 185
R109 source.n810 source.n809 185
R110 source.n808 source.n712 185
R111 source.n815 source.n711 185
R112 source.n817 source.n816 185
R113 source.n819 source.n818 185
R114 source.n708 source.n707 185
R115 source.n825 source.n824 185
R116 source.n827 source.n826 185
R117 source.n704 source.n703 185
R118 source.n833 source.n832 185
R119 source.n835 source.n834 185
R120 source.n604 source.n603 185
R121 source.n609 source.n608 185
R122 source.n611 source.n610 185
R123 source.n600 source.n599 185
R124 source.n617 source.n616 185
R125 source.n619 source.n618 185
R126 source.n596 source.n595 185
R127 source.n626 source.n625 185
R128 source.n627 source.n594 185
R129 source.n629 source.n628 185
R130 source.n592 source.n591 185
R131 source.n635 source.n634 185
R132 source.n637 source.n636 185
R133 source.n588 source.n587 185
R134 source.n643 source.n642 185
R135 source.n645 source.n644 185
R136 source.n584 source.n583 185
R137 source.n651 source.n650 185
R138 source.n653 source.n652 185
R139 source.n580 source.n579 185
R140 source.n659 source.n658 185
R141 source.n661 source.n660 185
R142 source.n576 source.n575 185
R143 source.n667 source.n666 185
R144 source.n670 source.n669 185
R145 source.n668 source.n572 185
R146 source.n675 source.n571 185
R147 source.n677 source.n676 185
R148 source.n679 source.n678 185
R149 source.n568 source.n567 185
R150 source.n685 source.n684 185
R151 source.n687 source.n686 185
R152 source.n564 source.n563 185
R153 source.n693 source.n692 185
R154 source.n695 source.n694 185
R155 source.n135 source.n134 185
R156 source.n133 source.n132 185
R157 source.n4 source.n3 185
R158 source.n127 source.n126 185
R159 source.n125 source.n124 185
R160 source.n8 source.n7 185
R161 source.n119 source.n118 185
R162 source.n117 source.n116 185
R163 source.n115 source.n11 185
R164 source.n15 source.n12 185
R165 source.n110 source.n109 185
R166 source.n108 source.n107 185
R167 source.n17 source.n16 185
R168 source.n102 source.n101 185
R169 source.n100 source.n99 185
R170 source.n21 source.n20 185
R171 source.n94 source.n93 185
R172 source.n92 source.n91 185
R173 source.n25 source.n24 185
R174 source.n86 source.n85 185
R175 source.n84 source.n83 185
R176 source.n29 source.n28 185
R177 source.n78 source.n77 185
R178 source.n76 source.n75 185
R179 source.n33 source.n32 185
R180 source.n70 source.n69 185
R181 source.n68 source.n35 185
R182 source.n67 source.n66 185
R183 source.n38 source.n36 185
R184 source.n61 source.n60 185
R185 source.n59 source.n58 185
R186 source.n42 source.n41 185
R187 source.n53 source.n52 185
R188 source.n51 source.n50 185
R189 source.n46 source.n45 185
R190 source.n275 source.n274 185
R191 source.n273 source.n272 185
R192 source.n144 source.n143 185
R193 source.n267 source.n266 185
R194 source.n265 source.n264 185
R195 source.n148 source.n147 185
R196 source.n259 source.n258 185
R197 source.n257 source.n256 185
R198 source.n255 source.n151 185
R199 source.n155 source.n152 185
R200 source.n250 source.n249 185
R201 source.n248 source.n247 185
R202 source.n157 source.n156 185
R203 source.n242 source.n241 185
R204 source.n240 source.n239 185
R205 source.n161 source.n160 185
R206 source.n234 source.n233 185
R207 source.n232 source.n231 185
R208 source.n165 source.n164 185
R209 source.n226 source.n225 185
R210 source.n224 source.n223 185
R211 source.n169 source.n168 185
R212 source.n218 source.n217 185
R213 source.n216 source.n215 185
R214 source.n173 source.n172 185
R215 source.n210 source.n209 185
R216 source.n208 source.n175 185
R217 source.n207 source.n206 185
R218 source.n178 source.n176 185
R219 source.n201 source.n200 185
R220 source.n199 source.n198 185
R221 source.n182 source.n181 185
R222 source.n193 source.n192 185
R223 source.n191 source.n190 185
R224 source.n186 source.n185 185
R225 source.n415 source.n414 185
R226 source.n413 source.n412 185
R227 source.n284 source.n283 185
R228 source.n407 source.n406 185
R229 source.n405 source.n404 185
R230 source.n288 source.n287 185
R231 source.n399 source.n398 185
R232 source.n397 source.n396 185
R233 source.n395 source.n291 185
R234 source.n295 source.n292 185
R235 source.n390 source.n389 185
R236 source.n388 source.n387 185
R237 source.n297 source.n296 185
R238 source.n382 source.n381 185
R239 source.n380 source.n379 185
R240 source.n301 source.n300 185
R241 source.n374 source.n373 185
R242 source.n372 source.n371 185
R243 source.n305 source.n304 185
R244 source.n366 source.n365 185
R245 source.n364 source.n363 185
R246 source.n309 source.n308 185
R247 source.n358 source.n357 185
R248 source.n356 source.n355 185
R249 source.n313 source.n312 185
R250 source.n350 source.n349 185
R251 source.n348 source.n315 185
R252 source.n347 source.n346 185
R253 source.n318 source.n316 185
R254 source.n341 source.n340 185
R255 source.n339 source.n338 185
R256 source.n322 source.n321 185
R257 source.n333 source.n332 185
R258 source.n331 source.n330 185
R259 source.n326 source.n325 185
R260 source.n555 source.n554 185
R261 source.n553 source.n552 185
R262 source.n424 source.n423 185
R263 source.n547 source.n546 185
R264 source.n545 source.n544 185
R265 source.n428 source.n427 185
R266 source.n539 source.n538 185
R267 source.n537 source.n536 185
R268 source.n535 source.n431 185
R269 source.n435 source.n432 185
R270 source.n530 source.n529 185
R271 source.n528 source.n527 185
R272 source.n437 source.n436 185
R273 source.n522 source.n521 185
R274 source.n520 source.n519 185
R275 source.n441 source.n440 185
R276 source.n514 source.n513 185
R277 source.n512 source.n511 185
R278 source.n445 source.n444 185
R279 source.n506 source.n505 185
R280 source.n504 source.n503 185
R281 source.n449 source.n448 185
R282 source.n498 source.n497 185
R283 source.n496 source.n495 185
R284 source.n453 source.n452 185
R285 source.n490 source.n489 185
R286 source.n488 source.n455 185
R287 source.n487 source.n486 185
R288 source.n458 source.n456 185
R289 source.n481 source.n480 185
R290 source.n479 source.n478 185
R291 source.n462 source.n461 185
R292 source.n473 source.n472 185
R293 source.n471 source.n470 185
R294 source.n466 source.n465 185
R295 source.n1025 source.t4 149.524
R296 source.n885 source.t7 149.524
R297 source.n745 source.t0 149.524
R298 source.n605 source.t3 149.524
R299 source.n47 source.t2 149.524
R300 source.n187 source.t1 149.524
R301 source.n327 source.t6 149.524
R302 source.n467 source.t5 149.524
R303 source.n1029 source.n1023 104.615
R304 source.n1030 source.n1029 104.615
R305 source.n1030 source.n1019 104.615
R306 source.n1037 source.n1019 104.615
R307 source.n1038 source.n1037 104.615
R308 source.n1038 source.n1015 104.615
R309 source.n1046 source.n1015 104.615
R310 source.n1047 source.n1046 104.615
R311 source.n1048 source.n1047 104.615
R312 source.n1048 source.n1011 104.615
R313 source.n1055 source.n1011 104.615
R314 source.n1056 source.n1055 104.615
R315 source.n1056 source.n1007 104.615
R316 source.n1063 source.n1007 104.615
R317 source.n1064 source.n1063 104.615
R318 source.n1064 source.n1003 104.615
R319 source.n1071 source.n1003 104.615
R320 source.n1072 source.n1071 104.615
R321 source.n1072 source.n999 104.615
R322 source.n1079 source.n999 104.615
R323 source.n1080 source.n1079 104.615
R324 source.n1080 source.n995 104.615
R325 source.n1087 source.n995 104.615
R326 source.n1089 source.n1087 104.615
R327 source.n1089 source.n1088 104.615
R328 source.n1088 source.n991 104.615
R329 source.n1097 source.n991 104.615
R330 source.n1098 source.n1097 104.615
R331 source.n1098 source.n987 104.615
R332 source.n1105 source.n987 104.615
R333 source.n1106 source.n1105 104.615
R334 source.n1106 source.n983 104.615
R335 source.n1113 source.n983 104.615
R336 source.n1114 source.n1113 104.615
R337 source.n889 source.n883 104.615
R338 source.n890 source.n889 104.615
R339 source.n890 source.n879 104.615
R340 source.n897 source.n879 104.615
R341 source.n898 source.n897 104.615
R342 source.n898 source.n875 104.615
R343 source.n906 source.n875 104.615
R344 source.n907 source.n906 104.615
R345 source.n908 source.n907 104.615
R346 source.n908 source.n871 104.615
R347 source.n915 source.n871 104.615
R348 source.n916 source.n915 104.615
R349 source.n916 source.n867 104.615
R350 source.n923 source.n867 104.615
R351 source.n924 source.n923 104.615
R352 source.n924 source.n863 104.615
R353 source.n931 source.n863 104.615
R354 source.n932 source.n931 104.615
R355 source.n932 source.n859 104.615
R356 source.n939 source.n859 104.615
R357 source.n940 source.n939 104.615
R358 source.n940 source.n855 104.615
R359 source.n947 source.n855 104.615
R360 source.n949 source.n947 104.615
R361 source.n949 source.n948 104.615
R362 source.n948 source.n851 104.615
R363 source.n957 source.n851 104.615
R364 source.n958 source.n957 104.615
R365 source.n958 source.n847 104.615
R366 source.n965 source.n847 104.615
R367 source.n966 source.n965 104.615
R368 source.n966 source.n843 104.615
R369 source.n973 source.n843 104.615
R370 source.n974 source.n973 104.615
R371 source.n749 source.n743 104.615
R372 source.n750 source.n749 104.615
R373 source.n750 source.n739 104.615
R374 source.n757 source.n739 104.615
R375 source.n758 source.n757 104.615
R376 source.n758 source.n735 104.615
R377 source.n766 source.n735 104.615
R378 source.n767 source.n766 104.615
R379 source.n768 source.n767 104.615
R380 source.n768 source.n731 104.615
R381 source.n775 source.n731 104.615
R382 source.n776 source.n775 104.615
R383 source.n776 source.n727 104.615
R384 source.n783 source.n727 104.615
R385 source.n784 source.n783 104.615
R386 source.n784 source.n723 104.615
R387 source.n791 source.n723 104.615
R388 source.n792 source.n791 104.615
R389 source.n792 source.n719 104.615
R390 source.n799 source.n719 104.615
R391 source.n800 source.n799 104.615
R392 source.n800 source.n715 104.615
R393 source.n807 source.n715 104.615
R394 source.n809 source.n807 104.615
R395 source.n809 source.n808 104.615
R396 source.n808 source.n711 104.615
R397 source.n817 source.n711 104.615
R398 source.n818 source.n817 104.615
R399 source.n818 source.n707 104.615
R400 source.n825 source.n707 104.615
R401 source.n826 source.n825 104.615
R402 source.n826 source.n703 104.615
R403 source.n833 source.n703 104.615
R404 source.n834 source.n833 104.615
R405 source.n609 source.n603 104.615
R406 source.n610 source.n609 104.615
R407 source.n610 source.n599 104.615
R408 source.n617 source.n599 104.615
R409 source.n618 source.n617 104.615
R410 source.n618 source.n595 104.615
R411 source.n626 source.n595 104.615
R412 source.n627 source.n626 104.615
R413 source.n628 source.n627 104.615
R414 source.n628 source.n591 104.615
R415 source.n635 source.n591 104.615
R416 source.n636 source.n635 104.615
R417 source.n636 source.n587 104.615
R418 source.n643 source.n587 104.615
R419 source.n644 source.n643 104.615
R420 source.n644 source.n583 104.615
R421 source.n651 source.n583 104.615
R422 source.n652 source.n651 104.615
R423 source.n652 source.n579 104.615
R424 source.n659 source.n579 104.615
R425 source.n660 source.n659 104.615
R426 source.n660 source.n575 104.615
R427 source.n667 source.n575 104.615
R428 source.n669 source.n667 104.615
R429 source.n669 source.n668 104.615
R430 source.n668 source.n571 104.615
R431 source.n677 source.n571 104.615
R432 source.n678 source.n677 104.615
R433 source.n678 source.n567 104.615
R434 source.n685 source.n567 104.615
R435 source.n686 source.n685 104.615
R436 source.n686 source.n563 104.615
R437 source.n693 source.n563 104.615
R438 source.n694 source.n693 104.615
R439 source.n134 source.n133 104.615
R440 source.n133 source.n3 104.615
R441 source.n126 source.n3 104.615
R442 source.n126 source.n125 104.615
R443 source.n125 source.n7 104.615
R444 source.n118 source.n7 104.615
R445 source.n118 source.n117 104.615
R446 source.n117 source.n11 104.615
R447 source.n15 source.n11 104.615
R448 source.n109 source.n15 104.615
R449 source.n109 source.n108 104.615
R450 source.n108 source.n16 104.615
R451 source.n101 source.n16 104.615
R452 source.n101 source.n100 104.615
R453 source.n100 source.n20 104.615
R454 source.n93 source.n20 104.615
R455 source.n93 source.n92 104.615
R456 source.n92 source.n24 104.615
R457 source.n85 source.n24 104.615
R458 source.n85 source.n84 104.615
R459 source.n84 source.n28 104.615
R460 source.n77 source.n28 104.615
R461 source.n77 source.n76 104.615
R462 source.n76 source.n32 104.615
R463 source.n69 source.n32 104.615
R464 source.n69 source.n68 104.615
R465 source.n68 source.n67 104.615
R466 source.n67 source.n36 104.615
R467 source.n60 source.n36 104.615
R468 source.n60 source.n59 104.615
R469 source.n59 source.n41 104.615
R470 source.n52 source.n41 104.615
R471 source.n52 source.n51 104.615
R472 source.n51 source.n45 104.615
R473 source.n274 source.n273 104.615
R474 source.n273 source.n143 104.615
R475 source.n266 source.n143 104.615
R476 source.n266 source.n265 104.615
R477 source.n265 source.n147 104.615
R478 source.n258 source.n147 104.615
R479 source.n258 source.n257 104.615
R480 source.n257 source.n151 104.615
R481 source.n155 source.n151 104.615
R482 source.n249 source.n155 104.615
R483 source.n249 source.n248 104.615
R484 source.n248 source.n156 104.615
R485 source.n241 source.n156 104.615
R486 source.n241 source.n240 104.615
R487 source.n240 source.n160 104.615
R488 source.n233 source.n160 104.615
R489 source.n233 source.n232 104.615
R490 source.n232 source.n164 104.615
R491 source.n225 source.n164 104.615
R492 source.n225 source.n224 104.615
R493 source.n224 source.n168 104.615
R494 source.n217 source.n168 104.615
R495 source.n217 source.n216 104.615
R496 source.n216 source.n172 104.615
R497 source.n209 source.n172 104.615
R498 source.n209 source.n208 104.615
R499 source.n208 source.n207 104.615
R500 source.n207 source.n176 104.615
R501 source.n200 source.n176 104.615
R502 source.n200 source.n199 104.615
R503 source.n199 source.n181 104.615
R504 source.n192 source.n181 104.615
R505 source.n192 source.n191 104.615
R506 source.n191 source.n185 104.615
R507 source.n414 source.n413 104.615
R508 source.n413 source.n283 104.615
R509 source.n406 source.n283 104.615
R510 source.n406 source.n405 104.615
R511 source.n405 source.n287 104.615
R512 source.n398 source.n287 104.615
R513 source.n398 source.n397 104.615
R514 source.n397 source.n291 104.615
R515 source.n295 source.n291 104.615
R516 source.n389 source.n295 104.615
R517 source.n389 source.n388 104.615
R518 source.n388 source.n296 104.615
R519 source.n381 source.n296 104.615
R520 source.n381 source.n380 104.615
R521 source.n380 source.n300 104.615
R522 source.n373 source.n300 104.615
R523 source.n373 source.n372 104.615
R524 source.n372 source.n304 104.615
R525 source.n365 source.n304 104.615
R526 source.n365 source.n364 104.615
R527 source.n364 source.n308 104.615
R528 source.n357 source.n308 104.615
R529 source.n357 source.n356 104.615
R530 source.n356 source.n312 104.615
R531 source.n349 source.n312 104.615
R532 source.n349 source.n348 104.615
R533 source.n348 source.n347 104.615
R534 source.n347 source.n316 104.615
R535 source.n340 source.n316 104.615
R536 source.n340 source.n339 104.615
R537 source.n339 source.n321 104.615
R538 source.n332 source.n321 104.615
R539 source.n332 source.n331 104.615
R540 source.n331 source.n325 104.615
R541 source.n554 source.n553 104.615
R542 source.n553 source.n423 104.615
R543 source.n546 source.n423 104.615
R544 source.n546 source.n545 104.615
R545 source.n545 source.n427 104.615
R546 source.n538 source.n427 104.615
R547 source.n538 source.n537 104.615
R548 source.n537 source.n431 104.615
R549 source.n435 source.n431 104.615
R550 source.n529 source.n435 104.615
R551 source.n529 source.n528 104.615
R552 source.n528 source.n436 104.615
R553 source.n521 source.n436 104.615
R554 source.n521 source.n520 104.615
R555 source.n520 source.n440 104.615
R556 source.n513 source.n440 104.615
R557 source.n513 source.n512 104.615
R558 source.n512 source.n444 104.615
R559 source.n505 source.n444 104.615
R560 source.n505 source.n504 104.615
R561 source.n504 source.n448 104.615
R562 source.n497 source.n448 104.615
R563 source.n497 source.n496 104.615
R564 source.n496 source.n452 104.615
R565 source.n489 source.n452 104.615
R566 source.n489 source.n488 104.615
R567 source.n488 source.n487 104.615
R568 source.n487 source.n456 104.615
R569 source.n480 source.n456 104.615
R570 source.n480 source.n479 104.615
R571 source.n479 source.n461 104.615
R572 source.n472 source.n461 104.615
R573 source.n472 source.n471 104.615
R574 source.n471 source.n465 104.615
R575 source.t4 source.n1023 52.3082
R576 source.t7 source.n883 52.3082
R577 source.t0 source.n743 52.3082
R578 source.t3 source.n603 52.3082
R579 source.t2 source.n45 52.3082
R580 source.t1 source.n185 52.3082
R581 source.t6 source.n325 52.3082
R582 source.t5 source.n465 52.3082
R583 source.n699 source.n559 31.6945
R584 source.n1119 source.n1118 30.6338
R585 source.n979 source.n978 30.6338
R586 source.n839 source.n838 30.6338
R587 source.n699 source.n698 30.6338
R588 source.n139 source.n138 30.6338
R589 source.n279 source.n278 30.6338
R590 source.n419 source.n418 30.6338
R591 source.n559 source.n558 30.6338
R592 source.n1120 source.n139 26.16
R593 source.n1049 source.n1014 13.1884
R594 source.n1096 source.n1095 13.1884
R595 source.n909 source.n874 13.1884
R596 source.n956 source.n955 13.1884
R597 source.n769 source.n734 13.1884
R598 source.n816 source.n815 13.1884
R599 source.n629 source.n594 13.1884
R600 source.n676 source.n675 13.1884
R601 source.n116 source.n115 13.1884
R602 source.n70 source.n35 13.1884
R603 source.n256 source.n255 13.1884
R604 source.n210 source.n175 13.1884
R605 source.n396 source.n395 13.1884
R606 source.n350 source.n315 13.1884
R607 source.n536 source.n535 13.1884
R608 source.n490 source.n455 13.1884
R609 source.n1045 source.n1044 12.8005
R610 source.n1050 source.n1012 12.8005
R611 source.n1094 source.n992 12.8005
R612 source.n1099 source.n990 12.8005
R613 source.n905 source.n904 12.8005
R614 source.n910 source.n872 12.8005
R615 source.n954 source.n852 12.8005
R616 source.n959 source.n850 12.8005
R617 source.n765 source.n764 12.8005
R618 source.n770 source.n732 12.8005
R619 source.n814 source.n712 12.8005
R620 source.n819 source.n710 12.8005
R621 source.n625 source.n624 12.8005
R622 source.n630 source.n592 12.8005
R623 source.n674 source.n572 12.8005
R624 source.n679 source.n570 12.8005
R625 source.n119 source.n10 12.8005
R626 source.n114 source.n12 12.8005
R627 source.n71 source.n33 12.8005
R628 source.n66 source.n37 12.8005
R629 source.n259 source.n150 12.8005
R630 source.n254 source.n152 12.8005
R631 source.n211 source.n173 12.8005
R632 source.n206 source.n177 12.8005
R633 source.n399 source.n290 12.8005
R634 source.n394 source.n292 12.8005
R635 source.n351 source.n313 12.8005
R636 source.n346 source.n317 12.8005
R637 source.n539 source.n430 12.8005
R638 source.n534 source.n432 12.8005
R639 source.n491 source.n453 12.8005
R640 source.n486 source.n457 12.8005
R641 source.n1043 source.n1016 12.0247
R642 source.n1054 source.n1053 12.0247
R643 source.n1091 source.n1090 12.0247
R644 source.n1100 source.n988 12.0247
R645 source.n903 source.n876 12.0247
R646 source.n914 source.n913 12.0247
R647 source.n951 source.n950 12.0247
R648 source.n960 source.n848 12.0247
R649 source.n763 source.n736 12.0247
R650 source.n774 source.n773 12.0247
R651 source.n811 source.n810 12.0247
R652 source.n820 source.n708 12.0247
R653 source.n623 source.n596 12.0247
R654 source.n634 source.n633 12.0247
R655 source.n671 source.n670 12.0247
R656 source.n680 source.n568 12.0247
R657 source.n120 source.n8 12.0247
R658 source.n111 source.n110 12.0247
R659 source.n75 source.n74 12.0247
R660 source.n65 source.n38 12.0247
R661 source.n260 source.n148 12.0247
R662 source.n251 source.n250 12.0247
R663 source.n215 source.n214 12.0247
R664 source.n205 source.n178 12.0247
R665 source.n400 source.n288 12.0247
R666 source.n391 source.n390 12.0247
R667 source.n355 source.n354 12.0247
R668 source.n345 source.n318 12.0247
R669 source.n540 source.n428 12.0247
R670 source.n531 source.n530 12.0247
R671 source.n495 source.n494 12.0247
R672 source.n485 source.n458 12.0247
R673 source.n1040 source.n1039 11.249
R674 source.n1057 source.n1010 11.249
R675 source.n1086 source.n994 11.249
R676 source.n1104 source.n1103 11.249
R677 source.n900 source.n899 11.249
R678 source.n917 source.n870 11.249
R679 source.n946 source.n854 11.249
R680 source.n964 source.n963 11.249
R681 source.n760 source.n759 11.249
R682 source.n777 source.n730 11.249
R683 source.n806 source.n714 11.249
R684 source.n824 source.n823 11.249
R685 source.n620 source.n619 11.249
R686 source.n637 source.n590 11.249
R687 source.n666 source.n574 11.249
R688 source.n684 source.n683 11.249
R689 source.n124 source.n123 11.249
R690 source.n107 source.n14 11.249
R691 source.n78 source.n31 11.249
R692 source.n62 source.n61 11.249
R693 source.n264 source.n263 11.249
R694 source.n247 source.n154 11.249
R695 source.n218 source.n171 11.249
R696 source.n202 source.n201 11.249
R697 source.n404 source.n403 11.249
R698 source.n387 source.n294 11.249
R699 source.n358 source.n311 11.249
R700 source.n342 source.n341 11.249
R701 source.n544 source.n543 11.249
R702 source.n527 source.n434 11.249
R703 source.n498 source.n451 11.249
R704 source.n482 source.n481 11.249
R705 source.n1036 source.n1018 10.4732
R706 source.n1058 source.n1008 10.4732
R707 source.n1085 source.n996 10.4732
R708 source.n1107 source.n986 10.4732
R709 source.n896 source.n878 10.4732
R710 source.n918 source.n868 10.4732
R711 source.n945 source.n856 10.4732
R712 source.n967 source.n846 10.4732
R713 source.n756 source.n738 10.4732
R714 source.n778 source.n728 10.4732
R715 source.n805 source.n716 10.4732
R716 source.n827 source.n706 10.4732
R717 source.n616 source.n598 10.4732
R718 source.n638 source.n588 10.4732
R719 source.n665 source.n576 10.4732
R720 source.n687 source.n566 10.4732
R721 source.n127 source.n6 10.4732
R722 source.n106 source.n17 10.4732
R723 source.n79 source.n29 10.4732
R724 source.n58 source.n40 10.4732
R725 source.n267 source.n146 10.4732
R726 source.n246 source.n157 10.4732
R727 source.n219 source.n169 10.4732
R728 source.n198 source.n180 10.4732
R729 source.n407 source.n286 10.4732
R730 source.n386 source.n297 10.4732
R731 source.n359 source.n309 10.4732
R732 source.n338 source.n320 10.4732
R733 source.n547 source.n426 10.4732
R734 source.n526 source.n437 10.4732
R735 source.n499 source.n449 10.4732
R736 source.n478 source.n460 10.4732
R737 source.n1025 source.n1024 10.2747
R738 source.n885 source.n884 10.2747
R739 source.n745 source.n744 10.2747
R740 source.n605 source.n604 10.2747
R741 source.n47 source.n46 10.2747
R742 source.n187 source.n186 10.2747
R743 source.n327 source.n326 10.2747
R744 source.n467 source.n466 10.2747
R745 source.n1035 source.n1020 9.69747
R746 source.n1062 source.n1061 9.69747
R747 source.n1082 source.n1081 9.69747
R748 source.n1108 source.n984 9.69747
R749 source.n895 source.n880 9.69747
R750 source.n922 source.n921 9.69747
R751 source.n942 source.n941 9.69747
R752 source.n968 source.n844 9.69747
R753 source.n755 source.n740 9.69747
R754 source.n782 source.n781 9.69747
R755 source.n802 source.n801 9.69747
R756 source.n828 source.n704 9.69747
R757 source.n615 source.n600 9.69747
R758 source.n642 source.n641 9.69747
R759 source.n662 source.n661 9.69747
R760 source.n688 source.n564 9.69747
R761 source.n128 source.n4 9.69747
R762 source.n103 source.n102 9.69747
R763 source.n83 source.n82 9.69747
R764 source.n57 source.n42 9.69747
R765 source.n268 source.n144 9.69747
R766 source.n243 source.n242 9.69747
R767 source.n223 source.n222 9.69747
R768 source.n197 source.n182 9.69747
R769 source.n408 source.n284 9.69747
R770 source.n383 source.n382 9.69747
R771 source.n363 source.n362 9.69747
R772 source.n337 source.n322 9.69747
R773 source.n548 source.n424 9.69747
R774 source.n523 source.n522 9.69747
R775 source.n503 source.n502 9.69747
R776 source.n477 source.n462 9.69747
R777 source.n1118 source.n1117 9.45567
R778 source.n978 source.n977 9.45567
R779 source.n838 source.n837 9.45567
R780 source.n698 source.n697 9.45567
R781 source.n138 source.n137 9.45567
R782 source.n278 source.n277 9.45567
R783 source.n418 source.n417 9.45567
R784 source.n558 source.n557 9.45567
R785 source.n982 source.n981 9.3005
R786 source.n1111 source.n1110 9.3005
R787 source.n1109 source.n1108 9.3005
R788 source.n986 source.n985 9.3005
R789 source.n1103 source.n1102 9.3005
R790 source.n1101 source.n1100 9.3005
R791 source.n990 source.n989 9.3005
R792 source.n1069 source.n1068 9.3005
R793 source.n1067 source.n1066 9.3005
R794 source.n1006 source.n1005 9.3005
R795 source.n1061 source.n1060 9.3005
R796 source.n1059 source.n1058 9.3005
R797 source.n1010 source.n1009 9.3005
R798 source.n1053 source.n1052 9.3005
R799 source.n1051 source.n1050 9.3005
R800 source.n1027 source.n1026 9.3005
R801 source.n1022 source.n1021 9.3005
R802 source.n1033 source.n1032 9.3005
R803 source.n1035 source.n1034 9.3005
R804 source.n1018 source.n1017 9.3005
R805 source.n1041 source.n1040 9.3005
R806 source.n1043 source.n1042 9.3005
R807 source.n1044 source.n1013 9.3005
R808 source.n1002 source.n1001 9.3005
R809 source.n1075 source.n1074 9.3005
R810 source.n1077 source.n1076 9.3005
R811 source.n998 source.n997 9.3005
R812 source.n1083 source.n1082 9.3005
R813 source.n1085 source.n1084 9.3005
R814 source.n994 source.n993 9.3005
R815 source.n1092 source.n1091 9.3005
R816 source.n1094 source.n1093 9.3005
R817 source.n1117 source.n1116 9.3005
R818 source.n842 source.n841 9.3005
R819 source.n971 source.n970 9.3005
R820 source.n969 source.n968 9.3005
R821 source.n846 source.n845 9.3005
R822 source.n963 source.n962 9.3005
R823 source.n961 source.n960 9.3005
R824 source.n850 source.n849 9.3005
R825 source.n929 source.n928 9.3005
R826 source.n927 source.n926 9.3005
R827 source.n866 source.n865 9.3005
R828 source.n921 source.n920 9.3005
R829 source.n919 source.n918 9.3005
R830 source.n870 source.n869 9.3005
R831 source.n913 source.n912 9.3005
R832 source.n911 source.n910 9.3005
R833 source.n887 source.n886 9.3005
R834 source.n882 source.n881 9.3005
R835 source.n893 source.n892 9.3005
R836 source.n895 source.n894 9.3005
R837 source.n878 source.n877 9.3005
R838 source.n901 source.n900 9.3005
R839 source.n903 source.n902 9.3005
R840 source.n904 source.n873 9.3005
R841 source.n862 source.n861 9.3005
R842 source.n935 source.n934 9.3005
R843 source.n937 source.n936 9.3005
R844 source.n858 source.n857 9.3005
R845 source.n943 source.n942 9.3005
R846 source.n945 source.n944 9.3005
R847 source.n854 source.n853 9.3005
R848 source.n952 source.n951 9.3005
R849 source.n954 source.n953 9.3005
R850 source.n977 source.n976 9.3005
R851 source.n702 source.n701 9.3005
R852 source.n831 source.n830 9.3005
R853 source.n829 source.n828 9.3005
R854 source.n706 source.n705 9.3005
R855 source.n823 source.n822 9.3005
R856 source.n821 source.n820 9.3005
R857 source.n710 source.n709 9.3005
R858 source.n789 source.n788 9.3005
R859 source.n787 source.n786 9.3005
R860 source.n726 source.n725 9.3005
R861 source.n781 source.n780 9.3005
R862 source.n779 source.n778 9.3005
R863 source.n730 source.n729 9.3005
R864 source.n773 source.n772 9.3005
R865 source.n771 source.n770 9.3005
R866 source.n747 source.n746 9.3005
R867 source.n742 source.n741 9.3005
R868 source.n753 source.n752 9.3005
R869 source.n755 source.n754 9.3005
R870 source.n738 source.n737 9.3005
R871 source.n761 source.n760 9.3005
R872 source.n763 source.n762 9.3005
R873 source.n764 source.n733 9.3005
R874 source.n722 source.n721 9.3005
R875 source.n795 source.n794 9.3005
R876 source.n797 source.n796 9.3005
R877 source.n718 source.n717 9.3005
R878 source.n803 source.n802 9.3005
R879 source.n805 source.n804 9.3005
R880 source.n714 source.n713 9.3005
R881 source.n812 source.n811 9.3005
R882 source.n814 source.n813 9.3005
R883 source.n837 source.n836 9.3005
R884 source.n562 source.n561 9.3005
R885 source.n691 source.n690 9.3005
R886 source.n689 source.n688 9.3005
R887 source.n566 source.n565 9.3005
R888 source.n683 source.n682 9.3005
R889 source.n681 source.n680 9.3005
R890 source.n570 source.n569 9.3005
R891 source.n649 source.n648 9.3005
R892 source.n647 source.n646 9.3005
R893 source.n586 source.n585 9.3005
R894 source.n641 source.n640 9.3005
R895 source.n639 source.n638 9.3005
R896 source.n590 source.n589 9.3005
R897 source.n633 source.n632 9.3005
R898 source.n631 source.n630 9.3005
R899 source.n607 source.n606 9.3005
R900 source.n602 source.n601 9.3005
R901 source.n613 source.n612 9.3005
R902 source.n615 source.n614 9.3005
R903 source.n598 source.n597 9.3005
R904 source.n621 source.n620 9.3005
R905 source.n623 source.n622 9.3005
R906 source.n624 source.n593 9.3005
R907 source.n582 source.n581 9.3005
R908 source.n655 source.n654 9.3005
R909 source.n657 source.n656 9.3005
R910 source.n578 source.n577 9.3005
R911 source.n663 source.n662 9.3005
R912 source.n665 source.n664 9.3005
R913 source.n574 source.n573 9.3005
R914 source.n672 source.n671 9.3005
R915 source.n674 source.n673 9.3005
R916 source.n697 source.n696 9.3005
R917 source.n49 source.n48 9.3005
R918 source.n44 source.n43 9.3005
R919 source.n55 source.n54 9.3005
R920 source.n57 source.n56 9.3005
R921 source.n40 source.n39 9.3005
R922 source.n63 source.n62 9.3005
R923 source.n65 source.n64 9.3005
R924 source.n37 source.n34 9.3005
R925 source.n96 source.n95 9.3005
R926 source.n98 source.n97 9.3005
R927 source.n19 source.n18 9.3005
R928 source.n104 source.n103 9.3005
R929 source.n106 source.n105 9.3005
R930 source.n14 source.n13 9.3005
R931 source.n112 source.n111 9.3005
R932 source.n114 source.n113 9.3005
R933 source.n137 source.n136 9.3005
R934 source.n2 source.n1 9.3005
R935 source.n131 source.n130 9.3005
R936 source.n129 source.n128 9.3005
R937 source.n6 source.n5 9.3005
R938 source.n123 source.n122 9.3005
R939 source.n121 source.n120 9.3005
R940 source.n10 source.n9 9.3005
R941 source.n23 source.n22 9.3005
R942 source.n90 source.n89 9.3005
R943 source.n88 source.n87 9.3005
R944 source.n27 source.n26 9.3005
R945 source.n82 source.n81 9.3005
R946 source.n80 source.n79 9.3005
R947 source.n31 source.n30 9.3005
R948 source.n74 source.n73 9.3005
R949 source.n72 source.n71 9.3005
R950 source.n189 source.n188 9.3005
R951 source.n184 source.n183 9.3005
R952 source.n195 source.n194 9.3005
R953 source.n197 source.n196 9.3005
R954 source.n180 source.n179 9.3005
R955 source.n203 source.n202 9.3005
R956 source.n205 source.n204 9.3005
R957 source.n177 source.n174 9.3005
R958 source.n236 source.n235 9.3005
R959 source.n238 source.n237 9.3005
R960 source.n159 source.n158 9.3005
R961 source.n244 source.n243 9.3005
R962 source.n246 source.n245 9.3005
R963 source.n154 source.n153 9.3005
R964 source.n252 source.n251 9.3005
R965 source.n254 source.n253 9.3005
R966 source.n277 source.n276 9.3005
R967 source.n142 source.n141 9.3005
R968 source.n271 source.n270 9.3005
R969 source.n269 source.n268 9.3005
R970 source.n146 source.n145 9.3005
R971 source.n263 source.n262 9.3005
R972 source.n261 source.n260 9.3005
R973 source.n150 source.n149 9.3005
R974 source.n163 source.n162 9.3005
R975 source.n230 source.n229 9.3005
R976 source.n228 source.n227 9.3005
R977 source.n167 source.n166 9.3005
R978 source.n222 source.n221 9.3005
R979 source.n220 source.n219 9.3005
R980 source.n171 source.n170 9.3005
R981 source.n214 source.n213 9.3005
R982 source.n212 source.n211 9.3005
R983 source.n329 source.n328 9.3005
R984 source.n324 source.n323 9.3005
R985 source.n335 source.n334 9.3005
R986 source.n337 source.n336 9.3005
R987 source.n320 source.n319 9.3005
R988 source.n343 source.n342 9.3005
R989 source.n345 source.n344 9.3005
R990 source.n317 source.n314 9.3005
R991 source.n376 source.n375 9.3005
R992 source.n378 source.n377 9.3005
R993 source.n299 source.n298 9.3005
R994 source.n384 source.n383 9.3005
R995 source.n386 source.n385 9.3005
R996 source.n294 source.n293 9.3005
R997 source.n392 source.n391 9.3005
R998 source.n394 source.n393 9.3005
R999 source.n417 source.n416 9.3005
R1000 source.n282 source.n281 9.3005
R1001 source.n411 source.n410 9.3005
R1002 source.n409 source.n408 9.3005
R1003 source.n286 source.n285 9.3005
R1004 source.n403 source.n402 9.3005
R1005 source.n401 source.n400 9.3005
R1006 source.n290 source.n289 9.3005
R1007 source.n303 source.n302 9.3005
R1008 source.n370 source.n369 9.3005
R1009 source.n368 source.n367 9.3005
R1010 source.n307 source.n306 9.3005
R1011 source.n362 source.n361 9.3005
R1012 source.n360 source.n359 9.3005
R1013 source.n311 source.n310 9.3005
R1014 source.n354 source.n353 9.3005
R1015 source.n352 source.n351 9.3005
R1016 source.n469 source.n468 9.3005
R1017 source.n464 source.n463 9.3005
R1018 source.n475 source.n474 9.3005
R1019 source.n477 source.n476 9.3005
R1020 source.n460 source.n459 9.3005
R1021 source.n483 source.n482 9.3005
R1022 source.n485 source.n484 9.3005
R1023 source.n457 source.n454 9.3005
R1024 source.n516 source.n515 9.3005
R1025 source.n518 source.n517 9.3005
R1026 source.n439 source.n438 9.3005
R1027 source.n524 source.n523 9.3005
R1028 source.n526 source.n525 9.3005
R1029 source.n434 source.n433 9.3005
R1030 source.n532 source.n531 9.3005
R1031 source.n534 source.n533 9.3005
R1032 source.n557 source.n556 9.3005
R1033 source.n422 source.n421 9.3005
R1034 source.n551 source.n550 9.3005
R1035 source.n549 source.n548 9.3005
R1036 source.n426 source.n425 9.3005
R1037 source.n543 source.n542 9.3005
R1038 source.n541 source.n540 9.3005
R1039 source.n430 source.n429 9.3005
R1040 source.n443 source.n442 9.3005
R1041 source.n510 source.n509 9.3005
R1042 source.n508 source.n507 9.3005
R1043 source.n447 source.n446 9.3005
R1044 source.n502 source.n501 9.3005
R1045 source.n500 source.n499 9.3005
R1046 source.n451 source.n450 9.3005
R1047 source.n494 source.n493 9.3005
R1048 source.n492 source.n491 9.3005
R1049 source.n1032 source.n1031 8.92171
R1050 source.n1065 source.n1006 8.92171
R1051 source.n1078 source.n998 8.92171
R1052 source.n1112 source.n1111 8.92171
R1053 source.n892 source.n891 8.92171
R1054 source.n925 source.n866 8.92171
R1055 source.n938 source.n858 8.92171
R1056 source.n972 source.n971 8.92171
R1057 source.n752 source.n751 8.92171
R1058 source.n785 source.n726 8.92171
R1059 source.n798 source.n718 8.92171
R1060 source.n832 source.n831 8.92171
R1061 source.n612 source.n611 8.92171
R1062 source.n645 source.n586 8.92171
R1063 source.n658 source.n578 8.92171
R1064 source.n692 source.n691 8.92171
R1065 source.n132 source.n131 8.92171
R1066 source.n99 source.n19 8.92171
R1067 source.n86 source.n27 8.92171
R1068 source.n54 source.n53 8.92171
R1069 source.n272 source.n271 8.92171
R1070 source.n239 source.n159 8.92171
R1071 source.n226 source.n167 8.92171
R1072 source.n194 source.n193 8.92171
R1073 source.n412 source.n411 8.92171
R1074 source.n379 source.n299 8.92171
R1075 source.n366 source.n307 8.92171
R1076 source.n334 source.n333 8.92171
R1077 source.n552 source.n551 8.92171
R1078 source.n519 source.n439 8.92171
R1079 source.n506 source.n447 8.92171
R1080 source.n474 source.n473 8.92171
R1081 source.n1028 source.n1022 8.14595
R1082 source.n1066 source.n1004 8.14595
R1083 source.n1077 source.n1000 8.14595
R1084 source.n1115 source.n982 8.14595
R1085 source.n888 source.n882 8.14595
R1086 source.n926 source.n864 8.14595
R1087 source.n937 source.n860 8.14595
R1088 source.n975 source.n842 8.14595
R1089 source.n748 source.n742 8.14595
R1090 source.n786 source.n724 8.14595
R1091 source.n797 source.n720 8.14595
R1092 source.n835 source.n702 8.14595
R1093 source.n608 source.n602 8.14595
R1094 source.n646 source.n584 8.14595
R1095 source.n657 source.n580 8.14595
R1096 source.n695 source.n562 8.14595
R1097 source.n135 source.n2 8.14595
R1098 source.n98 source.n21 8.14595
R1099 source.n87 source.n25 8.14595
R1100 source.n50 source.n44 8.14595
R1101 source.n275 source.n142 8.14595
R1102 source.n238 source.n161 8.14595
R1103 source.n227 source.n165 8.14595
R1104 source.n190 source.n184 8.14595
R1105 source.n415 source.n282 8.14595
R1106 source.n378 source.n301 8.14595
R1107 source.n367 source.n305 8.14595
R1108 source.n330 source.n324 8.14595
R1109 source.n555 source.n422 8.14595
R1110 source.n518 source.n441 8.14595
R1111 source.n507 source.n445 8.14595
R1112 source.n470 source.n464 8.14595
R1113 source.n1027 source.n1024 7.3702
R1114 source.n1070 source.n1069 7.3702
R1115 source.n1074 source.n1073 7.3702
R1116 source.n1116 source.n980 7.3702
R1117 source.n887 source.n884 7.3702
R1118 source.n930 source.n929 7.3702
R1119 source.n934 source.n933 7.3702
R1120 source.n976 source.n840 7.3702
R1121 source.n747 source.n744 7.3702
R1122 source.n790 source.n789 7.3702
R1123 source.n794 source.n793 7.3702
R1124 source.n836 source.n700 7.3702
R1125 source.n607 source.n604 7.3702
R1126 source.n650 source.n649 7.3702
R1127 source.n654 source.n653 7.3702
R1128 source.n696 source.n560 7.3702
R1129 source.n136 source.n0 7.3702
R1130 source.n95 source.n94 7.3702
R1131 source.n91 source.n90 7.3702
R1132 source.n49 source.n46 7.3702
R1133 source.n276 source.n140 7.3702
R1134 source.n235 source.n234 7.3702
R1135 source.n231 source.n230 7.3702
R1136 source.n189 source.n186 7.3702
R1137 source.n416 source.n280 7.3702
R1138 source.n375 source.n374 7.3702
R1139 source.n371 source.n370 7.3702
R1140 source.n329 source.n326 7.3702
R1141 source.n556 source.n420 7.3702
R1142 source.n515 source.n514 7.3702
R1143 source.n511 source.n510 7.3702
R1144 source.n469 source.n466 7.3702
R1145 source.n1070 source.n1002 6.59444
R1146 source.n1073 source.n1002 6.59444
R1147 source.n1118 source.n980 6.59444
R1148 source.n930 source.n862 6.59444
R1149 source.n933 source.n862 6.59444
R1150 source.n978 source.n840 6.59444
R1151 source.n790 source.n722 6.59444
R1152 source.n793 source.n722 6.59444
R1153 source.n838 source.n700 6.59444
R1154 source.n650 source.n582 6.59444
R1155 source.n653 source.n582 6.59444
R1156 source.n698 source.n560 6.59444
R1157 source.n138 source.n0 6.59444
R1158 source.n94 source.n23 6.59444
R1159 source.n91 source.n23 6.59444
R1160 source.n278 source.n140 6.59444
R1161 source.n234 source.n163 6.59444
R1162 source.n231 source.n163 6.59444
R1163 source.n418 source.n280 6.59444
R1164 source.n374 source.n303 6.59444
R1165 source.n371 source.n303 6.59444
R1166 source.n558 source.n420 6.59444
R1167 source.n514 source.n443 6.59444
R1168 source.n511 source.n443 6.59444
R1169 source.n1028 source.n1027 5.81868
R1170 source.n1069 source.n1004 5.81868
R1171 source.n1074 source.n1000 5.81868
R1172 source.n1116 source.n1115 5.81868
R1173 source.n888 source.n887 5.81868
R1174 source.n929 source.n864 5.81868
R1175 source.n934 source.n860 5.81868
R1176 source.n976 source.n975 5.81868
R1177 source.n748 source.n747 5.81868
R1178 source.n789 source.n724 5.81868
R1179 source.n794 source.n720 5.81868
R1180 source.n836 source.n835 5.81868
R1181 source.n608 source.n607 5.81868
R1182 source.n649 source.n584 5.81868
R1183 source.n654 source.n580 5.81868
R1184 source.n696 source.n695 5.81868
R1185 source.n136 source.n135 5.81868
R1186 source.n95 source.n21 5.81868
R1187 source.n90 source.n25 5.81868
R1188 source.n50 source.n49 5.81868
R1189 source.n276 source.n275 5.81868
R1190 source.n235 source.n161 5.81868
R1191 source.n230 source.n165 5.81868
R1192 source.n190 source.n189 5.81868
R1193 source.n416 source.n415 5.81868
R1194 source.n375 source.n301 5.81868
R1195 source.n370 source.n305 5.81868
R1196 source.n330 source.n329 5.81868
R1197 source.n556 source.n555 5.81868
R1198 source.n515 source.n441 5.81868
R1199 source.n510 source.n445 5.81868
R1200 source.n470 source.n469 5.81868
R1201 source.n1120 source.n1119 5.53498
R1202 source.n1031 source.n1022 5.04292
R1203 source.n1066 source.n1065 5.04292
R1204 source.n1078 source.n1077 5.04292
R1205 source.n1112 source.n982 5.04292
R1206 source.n891 source.n882 5.04292
R1207 source.n926 source.n925 5.04292
R1208 source.n938 source.n937 5.04292
R1209 source.n972 source.n842 5.04292
R1210 source.n751 source.n742 5.04292
R1211 source.n786 source.n785 5.04292
R1212 source.n798 source.n797 5.04292
R1213 source.n832 source.n702 5.04292
R1214 source.n611 source.n602 5.04292
R1215 source.n646 source.n645 5.04292
R1216 source.n658 source.n657 5.04292
R1217 source.n692 source.n562 5.04292
R1218 source.n132 source.n2 5.04292
R1219 source.n99 source.n98 5.04292
R1220 source.n87 source.n86 5.04292
R1221 source.n53 source.n44 5.04292
R1222 source.n272 source.n142 5.04292
R1223 source.n239 source.n238 5.04292
R1224 source.n227 source.n226 5.04292
R1225 source.n193 source.n184 5.04292
R1226 source.n412 source.n282 5.04292
R1227 source.n379 source.n378 5.04292
R1228 source.n367 source.n366 5.04292
R1229 source.n333 source.n324 5.04292
R1230 source.n552 source.n422 5.04292
R1231 source.n519 source.n518 5.04292
R1232 source.n507 source.n506 5.04292
R1233 source.n473 source.n464 5.04292
R1234 source.n1032 source.n1020 4.26717
R1235 source.n1062 source.n1006 4.26717
R1236 source.n1081 source.n998 4.26717
R1237 source.n1111 source.n984 4.26717
R1238 source.n892 source.n880 4.26717
R1239 source.n922 source.n866 4.26717
R1240 source.n941 source.n858 4.26717
R1241 source.n971 source.n844 4.26717
R1242 source.n752 source.n740 4.26717
R1243 source.n782 source.n726 4.26717
R1244 source.n801 source.n718 4.26717
R1245 source.n831 source.n704 4.26717
R1246 source.n612 source.n600 4.26717
R1247 source.n642 source.n586 4.26717
R1248 source.n661 source.n578 4.26717
R1249 source.n691 source.n564 4.26717
R1250 source.n131 source.n4 4.26717
R1251 source.n102 source.n19 4.26717
R1252 source.n83 source.n27 4.26717
R1253 source.n54 source.n42 4.26717
R1254 source.n271 source.n144 4.26717
R1255 source.n242 source.n159 4.26717
R1256 source.n223 source.n167 4.26717
R1257 source.n194 source.n182 4.26717
R1258 source.n411 source.n284 4.26717
R1259 source.n382 source.n299 4.26717
R1260 source.n363 source.n307 4.26717
R1261 source.n334 source.n322 4.26717
R1262 source.n551 source.n424 4.26717
R1263 source.n522 source.n439 4.26717
R1264 source.n503 source.n447 4.26717
R1265 source.n474 source.n462 4.26717
R1266 source.n1036 source.n1035 3.49141
R1267 source.n1061 source.n1008 3.49141
R1268 source.n1082 source.n996 3.49141
R1269 source.n1108 source.n1107 3.49141
R1270 source.n896 source.n895 3.49141
R1271 source.n921 source.n868 3.49141
R1272 source.n942 source.n856 3.49141
R1273 source.n968 source.n967 3.49141
R1274 source.n756 source.n755 3.49141
R1275 source.n781 source.n728 3.49141
R1276 source.n802 source.n716 3.49141
R1277 source.n828 source.n827 3.49141
R1278 source.n616 source.n615 3.49141
R1279 source.n641 source.n588 3.49141
R1280 source.n662 source.n576 3.49141
R1281 source.n688 source.n687 3.49141
R1282 source.n128 source.n127 3.49141
R1283 source.n103 source.n17 3.49141
R1284 source.n82 source.n29 3.49141
R1285 source.n58 source.n57 3.49141
R1286 source.n268 source.n267 3.49141
R1287 source.n243 source.n157 3.49141
R1288 source.n222 source.n169 3.49141
R1289 source.n198 source.n197 3.49141
R1290 source.n408 source.n407 3.49141
R1291 source.n383 source.n297 3.49141
R1292 source.n362 source.n309 3.49141
R1293 source.n338 source.n337 3.49141
R1294 source.n548 source.n547 3.49141
R1295 source.n523 source.n437 3.49141
R1296 source.n502 source.n449 3.49141
R1297 source.n478 source.n477 3.49141
R1298 source.n48 source.n47 2.84303
R1299 source.n188 source.n187 2.84303
R1300 source.n328 source.n327 2.84303
R1301 source.n468 source.n467 2.84303
R1302 source.n1026 source.n1025 2.84303
R1303 source.n886 source.n885 2.84303
R1304 source.n746 source.n745 2.84303
R1305 source.n606 source.n605 2.84303
R1306 source.n1039 source.n1018 2.71565
R1307 source.n1058 source.n1057 2.71565
R1308 source.n1086 source.n1085 2.71565
R1309 source.n1104 source.n986 2.71565
R1310 source.n899 source.n878 2.71565
R1311 source.n918 source.n917 2.71565
R1312 source.n946 source.n945 2.71565
R1313 source.n964 source.n846 2.71565
R1314 source.n759 source.n738 2.71565
R1315 source.n778 source.n777 2.71565
R1316 source.n806 source.n805 2.71565
R1317 source.n824 source.n706 2.71565
R1318 source.n619 source.n598 2.71565
R1319 source.n638 source.n637 2.71565
R1320 source.n666 source.n665 2.71565
R1321 source.n684 source.n566 2.71565
R1322 source.n124 source.n6 2.71565
R1323 source.n107 source.n106 2.71565
R1324 source.n79 source.n78 2.71565
R1325 source.n61 source.n40 2.71565
R1326 source.n264 source.n146 2.71565
R1327 source.n247 source.n246 2.71565
R1328 source.n219 source.n218 2.71565
R1329 source.n201 source.n180 2.71565
R1330 source.n404 source.n286 2.71565
R1331 source.n387 source.n386 2.71565
R1332 source.n359 source.n358 2.71565
R1333 source.n341 source.n320 2.71565
R1334 source.n544 source.n426 2.71565
R1335 source.n527 source.n526 2.71565
R1336 source.n499 source.n498 2.71565
R1337 source.n481 source.n460 2.71565
R1338 source.n1040 source.n1016 1.93989
R1339 source.n1054 source.n1010 1.93989
R1340 source.n1090 source.n994 1.93989
R1341 source.n1103 source.n988 1.93989
R1342 source.n900 source.n876 1.93989
R1343 source.n914 source.n870 1.93989
R1344 source.n950 source.n854 1.93989
R1345 source.n963 source.n848 1.93989
R1346 source.n760 source.n736 1.93989
R1347 source.n774 source.n730 1.93989
R1348 source.n810 source.n714 1.93989
R1349 source.n823 source.n708 1.93989
R1350 source.n620 source.n596 1.93989
R1351 source.n634 source.n590 1.93989
R1352 source.n670 source.n574 1.93989
R1353 source.n683 source.n568 1.93989
R1354 source.n123 source.n8 1.93989
R1355 source.n110 source.n14 1.93989
R1356 source.n75 source.n31 1.93989
R1357 source.n62 source.n38 1.93989
R1358 source.n263 source.n148 1.93989
R1359 source.n250 source.n154 1.93989
R1360 source.n215 source.n171 1.93989
R1361 source.n202 source.n178 1.93989
R1362 source.n403 source.n288 1.93989
R1363 source.n390 source.n294 1.93989
R1364 source.n355 source.n311 1.93989
R1365 source.n342 source.n318 1.93989
R1366 source.n543 source.n428 1.93989
R1367 source.n530 source.n434 1.93989
R1368 source.n495 source.n451 1.93989
R1369 source.n482 source.n458 1.93989
R1370 source.n1045 source.n1043 1.16414
R1371 source.n1053 source.n1012 1.16414
R1372 source.n1091 source.n992 1.16414
R1373 source.n1100 source.n1099 1.16414
R1374 source.n905 source.n903 1.16414
R1375 source.n913 source.n872 1.16414
R1376 source.n951 source.n852 1.16414
R1377 source.n960 source.n959 1.16414
R1378 source.n765 source.n763 1.16414
R1379 source.n773 source.n732 1.16414
R1380 source.n811 source.n712 1.16414
R1381 source.n820 source.n819 1.16414
R1382 source.n625 source.n623 1.16414
R1383 source.n633 source.n592 1.16414
R1384 source.n671 source.n572 1.16414
R1385 source.n680 source.n679 1.16414
R1386 source.n120 source.n119 1.16414
R1387 source.n111 source.n12 1.16414
R1388 source.n74 source.n33 1.16414
R1389 source.n66 source.n65 1.16414
R1390 source.n260 source.n259 1.16414
R1391 source.n251 source.n152 1.16414
R1392 source.n214 source.n173 1.16414
R1393 source.n206 source.n205 1.16414
R1394 source.n400 source.n399 1.16414
R1395 source.n391 source.n292 1.16414
R1396 source.n354 source.n313 1.16414
R1397 source.n346 source.n345 1.16414
R1398 source.n540 source.n539 1.16414
R1399 source.n531 source.n432 1.16414
R1400 source.n494 source.n453 1.16414
R1401 source.n486 source.n485 1.16414
R1402 source.n559 source.n419 0.543603
R1403 source.n279 source.n139 0.543603
R1404 source.n839 source.n699 0.543603
R1405 source.n1119 source.n979 0.543603
R1406 source.n419 source.n279 0.470328
R1407 source.n979 source.n839 0.470328
R1408 source.n1044 source.n1014 0.388379
R1409 source.n1050 source.n1049 0.388379
R1410 source.n1095 source.n1094 0.388379
R1411 source.n1096 source.n990 0.388379
R1412 source.n904 source.n874 0.388379
R1413 source.n910 source.n909 0.388379
R1414 source.n955 source.n954 0.388379
R1415 source.n956 source.n850 0.388379
R1416 source.n764 source.n734 0.388379
R1417 source.n770 source.n769 0.388379
R1418 source.n815 source.n814 0.388379
R1419 source.n816 source.n710 0.388379
R1420 source.n624 source.n594 0.388379
R1421 source.n630 source.n629 0.388379
R1422 source.n675 source.n674 0.388379
R1423 source.n676 source.n570 0.388379
R1424 source.n116 source.n10 0.388379
R1425 source.n115 source.n114 0.388379
R1426 source.n71 source.n70 0.388379
R1427 source.n37 source.n35 0.388379
R1428 source.n256 source.n150 0.388379
R1429 source.n255 source.n254 0.388379
R1430 source.n211 source.n210 0.388379
R1431 source.n177 source.n175 0.388379
R1432 source.n396 source.n290 0.388379
R1433 source.n395 source.n394 0.388379
R1434 source.n351 source.n350 0.388379
R1435 source.n317 source.n315 0.388379
R1436 source.n536 source.n430 0.388379
R1437 source.n535 source.n534 0.388379
R1438 source.n491 source.n490 0.388379
R1439 source.n457 source.n455 0.388379
R1440 source source.n1120 0.188
R1441 source.n1026 source.n1021 0.155672
R1442 source.n1033 source.n1021 0.155672
R1443 source.n1034 source.n1033 0.155672
R1444 source.n1034 source.n1017 0.155672
R1445 source.n1041 source.n1017 0.155672
R1446 source.n1042 source.n1041 0.155672
R1447 source.n1042 source.n1013 0.155672
R1448 source.n1051 source.n1013 0.155672
R1449 source.n1052 source.n1051 0.155672
R1450 source.n1052 source.n1009 0.155672
R1451 source.n1059 source.n1009 0.155672
R1452 source.n1060 source.n1059 0.155672
R1453 source.n1060 source.n1005 0.155672
R1454 source.n1067 source.n1005 0.155672
R1455 source.n1068 source.n1067 0.155672
R1456 source.n1068 source.n1001 0.155672
R1457 source.n1075 source.n1001 0.155672
R1458 source.n1076 source.n1075 0.155672
R1459 source.n1076 source.n997 0.155672
R1460 source.n1083 source.n997 0.155672
R1461 source.n1084 source.n1083 0.155672
R1462 source.n1084 source.n993 0.155672
R1463 source.n1092 source.n993 0.155672
R1464 source.n1093 source.n1092 0.155672
R1465 source.n1093 source.n989 0.155672
R1466 source.n1101 source.n989 0.155672
R1467 source.n1102 source.n1101 0.155672
R1468 source.n1102 source.n985 0.155672
R1469 source.n1109 source.n985 0.155672
R1470 source.n1110 source.n1109 0.155672
R1471 source.n1110 source.n981 0.155672
R1472 source.n1117 source.n981 0.155672
R1473 source.n886 source.n881 0.155672
R1474 source.n893 source.n881 0.155672
R1475 source.n894 source.n893 0.155672
R1476 source.n894 source.n877 0.155672
R1477 source.n901 source.n877 0.155672
R1478 source.n902 source.n901 0.155672
R1479 source.n902 source.n873 0.155672
R1480 source.n911 source.n873 0.155672
R1481 source.n912 source.n911 0.155672
R1482 source.n912 source.n869 0.155672
R1483 source.n919 source.n869 0.155672
R1484 source.n920 source.n919 0.155672
R1485 source.n920 source.n865 0.155672
R1486 source.n927 source.n865 0.155672
R1487 source.n928 source.n927 0.155672
R1488 source.n928 source.n861 0.155672
R1489 source.n935 source.n861 0.155672
R1490 source.n936 source.n935 0.155672
R1491 source.n936 source.n857 0.155672
R1492 source.n943 source.n857 0.155672
R1493 source.n944 source.n943 0.155672
R1494 source.n944 source.n853 0.155672
R1495 source.n952 source.n853 0.155672
R1496 source.n953 source.n952 0.155672
R1497 source.n953 source.n849 0.155672
R1498 source.n961 source.n849 0.155672
R1499 source.n962 source.n961 0.155672
R1500 source.n962 source.n845 0.155672
R1501 source.n969 source.n845 0.155672
R1502 source.n970 source.n969 0.155672
R1503 source.n970 source.n841 0.155672
R1504 source.n977 source.n841 0.155672
R1505 source.n746 source.n741 0.155672
R1506 source.n753 source.n741 0.155672
R1507 source.n754 source.n753 0.155672
R1508 source.n754 source.n737 0.155672
R1509 source.n761 source.n737 0.155672
R1510 source.n762 source.n761 0.155672
R1511 source.n762 source.n733 0.155672
R1512 source.n771 source.n733 0.155672
R1513 source.n772 source.n771 0.155672
R1514 source.n772 source.n729 0.155672
R1515 source.n779 source.n729 0.155672
R1516 source.n780 source.n779 0.155672
R1517 source.n780 source.n725 0.155672
R1518 source.n787 source.n725 0.155672
R1519 source.n788 source.n787 0.155672
R1520 source.n788 source.n721 0.155672
R1521 source.n795 source.n721 0.155672
R1522 source.n796 source.n795 0.155672
R1523 source.n796 source.n717 0.155672
R1524 source.n803 source.n717 0.155672
R1525 source.n804 source.n803 0.155672
R1526 source.n804 source.n713 0.155672
R1527 source.n812 source.n713 0.155672
R1528 source.n813 source.n812 0.155672
R1529 source.n813 source.n709 0.155672
R1530 source.n821 source.n709 0.155672
R1531 source.n822 source.n821 0.155672
R1532 source.n822 source.n705 0.155672
R1533 source.n829 source.n705 0.155672
R1534 source.n830 source.n829 0.155672
R1535 source.n830 source.n701 0.155672
R1536 source.n837 source.n701 0.155672
R1537 source.n606 source.n601 0.155672
R1538 source.n613 source.n601 0.155672
R1539 source.n614 source.n613 0.155672
R1540 source.n614 source.n597 0.155672
R1541 source.n621 source.n597 0.155672
R1542 source.n622 source.n621 0.155672
R1543 source.n622 source.n593 0.155672
R1544 source.n631 source.n593 0.155672
R1545 source.n632 source.n631 0.155672
R1546 source.n632 source.n589 0.155672
R1547 source.n639 source.n589 0.155672
R1548 source.n640 source.n639 0.155672
R1549 source.n640 source.n585 0.155672
R1550 source.n647 source.n585 0.155672
R1551 source.n648 source.n647 0.155672
R1552 source.n648 source.n581 0.155672
R1553 source.n655 source.n581 0.155672
R1554 source.n656 source.n655 0.155672
R1555 source.n656 source.n577 0.155672
R1556 source.n663 source.n577 0.155672
R1557 source.n664 source.n663 0.155672
R1558 source.n664 source.n573 0.155672
R1559 source.n672 source.n573 0.155672
R1560 source.n673 source.n672 0.155672
R1561 source.n673 source.n569 0.155672
R1562 source.n681 source.n569 0.155672
R1563 source.n682 source.n681 0.155672
R1564 source.n682 source.n565 0.155672
R1565 source.n689 source.n565 0.155672
R1566 source.n690 source.n689 0.155672
R1567 source.n690 source.n561 0.155672
R1568 source.n697 source.n561 0.155672
R1569 source.n137 source.n1 0.155672
R1570 source.n130 source.n1 0.155672
R1571 source.n130 source.n129 0.155672
R1572 source.n129 source.n5 0.155672
R1573 source.n122 source.n5 0.155672
R1574 source.n122 source.n121 0.155672
R1575 source.n121 source.n9 0.155672
R1576 source.n113 source.n9 0.155672
R1577 source.n113 source.n112 0.155672
R1578 source.n112 source.n13 0.155672
R1579 source.n105 source.n13 0.155672
R1580 source.n105 source.n104 0.155672
R1581 source.n104 source.n18 0.155672
R1582 source.n97 source.n18 0.155672
R1583 source.n97 source.n96 0.155672
R1584 source.n96 source.n22 0.155672
R1585 source.n89 source.n22 0.155672
R1586 source.n89 source.n88 0.155672
R1587 source.n88 source.n26 0.155672
R1588 source.n81 source.n26 0.155672
R1589 source.n81 source.n80 0.155672
R1590 source.n80 source.n30 0.155672
R1591 source.n73 source.n30 0.155672
R1592 source.n73 source.n72 0.155672
R1593 source.n72 source.n34 0.155672
R1594 source.n64 source.n34 0.155672
R1595 source.n64 source.n63 0.155672
R1596 source.n63 source.n39 0.155672
R1597 source.n56 source.n39 0.155672
R1598 source.n56 source.n55 0.155672
R1599 source.n55 source.n43 0.155672
R1600 source.n48 source.n43 0.155672
R1601 source.n277 source.n141 0.155672
R1602 source.n270 source.n141 0.155672
R1603 source.n270 source.n269 0.155672
R1604 source.n269 source.n145 0.155672
R1605 source.n262 source.n145 0.155672
R1606 source.n262 source.n261 0.155672
R1607 source.n261 source.n149 0.155672
R1608 source.n253 source.n149 0.155672
R1609 source.n253 source.n252 0.155672
R1610 source.n252 source.n153 0.155672
R1611 source.n245 source.n153 0.155672
R1612 source.n245 source.n244 0.155672
R1613 source.n244 source.n158 0.155672
R1614 source.n237 source.n158 0.155672
R1615 source.n237 source.n236 0.155672
R1616 source.n236 source.n162 0.155672
R1617 source.n229 source.n162 0.155672
R1618 source.n229 source.n228 0.155672
R1619 source.n228 source.n166 0.155672
R1620 source.n221 source.n166 0.155672
R1621 source.n221 source.n220 0.155672
R1622 source.n220 source.n170 0.155672
R1623 source.n213 source.n170 0.155672
R1624 source.n213 source.n212 0.155672
R1625 source.n212 source.n174 0.155672
R1626 source.n204 source.n174 0.155672
R1627 source.n204 source.n203 0.155672
R1628 source.n203 source.n179 0.155672
R1629 source.n196 source.n179 0.155672
R1630 source.n196 source.n195 0.155672
R1631 source.n195 source.n183 0.155672
R1632 source.n188 source.n183 0.155672
R1633 source.n417 source.n281 0.155672
R1634 source.n410 source.n281 0.155672
R1635 source.n410 source.n409 0.155672
R1636 source.n409 source.n285 0.155672
R1637 source.n402 source.n285 0.155672
R1638 source.n402 source.n401 0.155672
R1639 source.n401 source.n289 0.155672
R1640 source.n393 source.n289 0.155672
R1641 source.n393 source.n392 0.155672
R1642 source.n392 source.n293 0.155672
R1643 source.n385 source.n293 0.155672
R1644 source.n385 source.n384 0.155672
R1645 source.n384 source.n298 0.155672
R1646 source.n377 source.n298 0.155672
R1647 source.n377 source.n376 0.155672
R1648 source.n376 source.n302 0.155672
R1649 source.n369 source.n302 0.155672
R1650 source.n369 source.n368 0.155672
R1651 source.n368 source.n306 0.155672
R1652 source.n361 source.n306 0.155672
R1653 source.n361 source.n360 0.155672
R1654 source.n360 source.n310 0.155672
R1655 source.n353 source.n310 0.155672
R1656 source.n353 source.n352 0.155672
R1657 source.n352 source.n314 0.155672
R1658 source.n344 source.n314 0.155672
R1659 source.n344 source.n343 0.155672
R1660 source.n343 source.n319 0.155672
R1661 source.n336 source.n319 0.155672
R1662 source.n336 source.n335 0.155672
R1663 source.n335 source.n323 0.155672
R1664 source.n328 source.n323 0.155672
R1665 source.n557 source.n421 0.155672
R1666 source.n550 source.n421 0.155672
R1667 source.n550 source.n549 0.155672
R1668 source.n549 source.n425 0.155672
R1669 source.n542 source.n425 0.155672
R1670 source.n542 source.n541 0.155672
R1671 source.n541 source.n429 0.155672
R1672 source.n533 source.n429 0.155672
R1673 source.n533 source.n532 0.155672
R1674 source.n532 source.n433 0.155672
R1675 source.n525 source.n433 0.155672
R1676 source.n525 source.n524 0.155672
R1677 source.n524 source.n438 0.155672
R1678 source.n517 source.n438 0.155672
R1679 source.n517 source.n516 0.155672
R1680 source.n516 source.n442 0.155672
R1681 source.n509 source.n442 0.155672
R1682 source.n509 source.n508 0.155672
R1683 source.n508 source.n446 0.155672
R1684 source.n501 source.n446 0.155672
R1685 source.n501 source.n500 0.155672
R1686 source.n500 source.n450 0.155672
R1687 source.n493 source.n450 0.155672
R1688 source.n493 source.n492 0.155672
R1689 source.n492 source.n454 0.155672
R1690 source.n484 source.n454 0.155672
R1691 source.n484 source.n483 0.155672
R1692 source.n483 source.n459 0.155672
R1693 source.n476 source.n459 0.155672
R1694 source.n476 source.n475 0.155672
R1695 source.n475 source.n463 0.155672
R1696 source.n468 source.n463 0.155672
R1697 drain_right drain_right.n0 96.4786
R1698 drain_right drain_right.n1 64.9111
R1699 drain_right.n0 drain_right.t0 0.7925
R1700 drain_right.n0 drain_right.t2 0.7925
R1701 drain_right.n1 drain_right.t1 0.7925
R1702 drain_right.n1 drain_right.t3 0.7925
R1703 plus.n0 plus.t2 2158.78
R1704 plus.n0 plus.t3 2158.78
R1705 plus.n1 plus.t1 2158.78
R1706 plus.n1 plus.t0 2158.78
R1707 plus plus.n1 193.393
R1708 plus plus.n0 178.376
R1709 drain_left drain_left.n0 97.0318
R1710 drain_left drain_left.n1 64.9111
R1711 drain_left.n0 drain_left.t3 0.7925
R1712 drain_left.n0 drain_left.t2 0.7925
R1713 drain_left.n1 drain_left.t1 0.7925
R1714 drain_left.n1 drain_left.t0 0.7925
C0 drain_left source 18.537699f
C1 drain_right drain_left 0.477421f
C2 plus drain_left 4.1751f
C3 drain_left minus 0.171331f
C4 drain_right source 18.5362f
C5 plus source 2.96183f
C6 drain_right plus 0.255071f
C7 source minus 2.94779f
C8 drain_right minus 4.07415f
C9 plus minus 6.91591f
C10 drain_right a_n1094_n5892# 10.241549f
C11 drain_left a_n1094_n5892# 10.434311f
C12 source a_n1094_n5892# 15.877192f
C13 minus a_n1094_n5892# 5.038014f
C14 plus a_n1094_n5892# 11.137929f
C15 drain_left.t3 a_n1094_n5892# 0.656897f
C16 drain_left.t2 a_n1094_n5892# 0.656897f
C17 drain_left.n0 a_n1094_n5892# 7.08747f
C18 drain_left.t1 a_n1094_n5892# 0.656897f
C19 drain_left.t0 a_n1094_n5892# 0.656897f
C20 drain_left.n1 a_n1094_n5892# 6.11964f
C21 plus.t2 a_n1094_n5892# 1.34573f
C22 plus.t3 a_n1094_n5892# 1.34573f
C23 plus.n0 a_n1094_n5892# 1.09574f
C24 plus.t0 a_n1094_n5892# 1.34573f
C25 plus.t1 a_n1094_n5892# 1.34573f
C26 plus.n1 a_n1094_n5892# 1.35427f
C27 drain_right.t0 a_n1094_n5892# 0.657772f
C28 drain_right.t2 a_n1094_n5892# 0.657772f
C29 drain_right.n0 a_n1094_n5892# 7.06052f
C30 drain_right.t1 a_n1094_n5892# 0.657772f
C31 drain_right.t3 a_n1094_n5892# 0.657772f
C32 drain_right.n1 a_n1094_n5892# 6.12779f
C33 source.n0 a_n1094_n5892# 0.025218f
C34 source.n1 a_n1094_n5892# 0.018292f
C35 source.n2 a_n1094_n5892# 0.009829f
C36 source.n3 a_n1094_n5892# 0.023233f
C37 source.n4 a_n1094_n5892# 0.010408f
C38 source.n5 a_n1094_n5892# 0.018292f
C39 source.n6 a_n1094_n5892# 0.009829f
C40 source.n7 a_n1094_n5892# 0.023233f
C41 source.n8 a_n1094_n5892# 0.010408f
C42 source.n9 a_n1094_n5892# 0.018292f
C43 source.n10 a_n1094_n5892# 0.009829f
C44 source.n11 a_n1094_n5892# 0.023233f
C45 source.n12 a_n1094_n5892# 0.010408f
C46 source.n13 a_n1094_n5892# 0.018292f
C47 source.n14 a_n1094_n5892# 0.009829f
C48 source.n15 a_n1094_n5892# 0.023233f
C49 source.n16 a_n1094_n5892# 0.023233f
C50 source.n17 a_n1094_n5892# 0.010408f
C51 source.n18 a_n1094_n5892# 0.018292f
C52 source.n19 a_n1094_n5892# 0.009829f
C53 source.n20 a_n1094_n5892# 0.023233f
C54 source.n21 a_n1094_n5892# 0.010408f
C55 source.n22 a_n1094_n5892# 0.018292f
C56 source.n23 a_n1094_n5892# 0.009829f
C57 source.n24 a_n1094_n5892# 0.023233f
C58 source.n25 a_n1094_n5892# 0.010408f
C59 source.n26 a_n1094_n5892# 0.018292f
C60 source.n27 a_n1094_n5892# 0.009829f
C61 source.n28 a_n1094_n5892# 0.023233f
C62 source.n29 a_n1094_n5892# 0.010408f
C63 source.n30 a_n1094_n5892# 0.018292f
C64 source.n31 a_n1094_n5892# 0.009829f
C65 source.n32 a_n1094_n5892# 0.023233f
C66 source.n33 a_n1094_n5892# 0.010408f
C67 source.n34 a_n1094_n5892# 0.018292f
C68 source.n35 a_n1094_n5892# 0.010119f
C69 source.n36 a_n1094_n5892# 0.023233f
C70 source.n37 a_n1094_n5892# 0.009829f
C71 source.n38 a_n1094_n5892# 0.010408f
C72 source.n39 a_n1094_n5892# 0.018292f
C73 source.n40 a_n1094_n5892# 0.009829f
C74 source.n41 a_n1094_n5892# 0.023233f
C75 source.n42 a_n1094_n5892# 0.010408f
C76 source.n43 a_n1094_n5892# 0.018292f
C77 source.n44 a_n1094_n5892# 0.009829f
C78 source.n45 a_n1094_n5892# 0.017425f
C79 source.n46 a_n1094_n5892# 0.016424f
C80 source.t2 a_n1094_n5892# 0.04052f
C81 source.n47 a_n1094_n5892# 0.223181f
C82 source.n48 a_n1094_n5892# 1.98052f
C83 source.n49 a_n1094_n5892# 0.009829f
C84 source.n50 a_n1094_n5892# 0.010408f
C85 source.n51 a_n1094_n5892# 0.023233f
C86 source.n52 a_n1094_n5892# 0.023233f
C87 source.n53 a_n1094_n5892# 0.010408f
C88 source.n54 a_n1094_n5892# 0.009829f
C89 source.n55 a_n1094_n5892# 0.018292f
C90 source.n56 a_n1094_n5892# 0.018292f
C91 source.n57 a_n1094_n5892# 0.009829f
C92 source.n58 a_n1094_n5892# 0.010408f
C93 source.n59 a_n1094_n5892# 0.023233f
C94 source.n60 a_n1094_n5892# 0.023233f
C95 source.n61 a_n1094_n5892# 0.010408f
C96 source.n62 a_n1094_n5892# 0.009829f
C97 source.n63 a_n1094_n5892# 0.018292f
C98 source.n64 a_n1094_n5892# 0.018292f
C99 source.n65 a_n1094_n5892# 0.009829f
C100 source.n66 a_n1094_n5892# 0.010408f
C101 source.n67 a_n1094_n5892# 0.023233f
C102 source.n68 a_n1094_n5892# 0.023233f
C103 source.n69 a_n1094_n5892# 0.023233f
C104 source.n70 a_n1094_n5892# 0.010119f
C105 source.n71 a_n1094_n5892# 0.009829f
C106 source.n72 a_n1094_n5892# 0.018292f
C107 source.n73 a_n1094_n5892# 0.018292f
C108 source.n74 a_n1094_n5892# 0.009829f
C109 source.n75 a_n1094_n5892# 0.010408f
C110 source.n76 a_n1094_n5892# 0.023233f
C111 source.n77 a_n1094_n5892# 0.023233f
C112 source.n78 a_n1094_n5892# 0.010408f
C113 source.n79 a_n1094_n5892# 0.009829f
C114 source.n80 a_n1094_n5892# 0.018292f
C115 source.n81 a_n1094_n5892# 0.018292f
C116 source.n82 a_n1094_n5892# 0.009829f
C117 source.n83 a_n1094_n5892# 0.010408f
C118 source.n84 a_n1094_n5892# 0.023233f
C119 source.n85 a_n1094_n5892# 0.023233f
C120 source.n86 a_n1094_n5892# 0.010408f
C121 source.n87 a_n1094_n5892# 0.009829f
C122 source.n88 a_n1094_n5892# 0.018292f
C123 source.n89 a_n1094_n5892# 0.018292f
C124 source.n90 a_n1094_n5892# 0.009829f
C125 source.n91 a_n1094_n5892# 0.010408f
C126 source.n92 a_n1094_n5892# 0.023233f
C127 source.n93 a_n1094_n5892# 0.023233f
C128 source.n94 a_n1094_n5892# 0.010408f
C129 source.n95 a_n1094_n5892# 0.009829f
C130 source.n96 a_n1094_n5892# 0.018292f
C131 source.n97 a_n1094_n5892# 0.018292f
C132 source.n98 a_n1094_n5892# 0.009829f
C133 source.n99 a_n1094_n5892# 0.010408f
C134 source.n100 a_n1094_n5892# 0.023233f
C135 source.n101 a_n1094_n5892# 0.023233f
C136 source.n102 a_n1094_n5892# 0.010408f
C137 source.n103 a_n1094_n5892# 0.009829f
C138 source.n104 a_n1094_n5892# 0.018292f
C139 source.n105 a_n1094_n5892# 0.018292f
C140 source.n106 a_n1094_n5892# 0.009829f
C141 source.n107 a_n1094_n5892# 0.010408f
C142 source.n108 a_n1094_n5892# 0.023233f
C143 source.n109 a_n1094_n5892# 0.023233f
C144 source.n110 a_n1094_n5892# 0.010408f
C145 source.n111 a_n1094_n5892# 0.009829f
C146 source.n112 a_n1094_n5892# 0.018292f
C147 source.n113 a_n1094_n5892# 0.018292f
C148 source.n114 a_n1094_n5892# 0.009829f
C149 source.n115 a_n1094_n5892# 0.010119f
C150 source.n116 a_n1094_n5892# 0.010119f
C151 source.n117 a_n1094_n5892# 0.023233f
C152 source.n118 a_n1094_n5892# 0.023233f
C153 source.n119 a_n1094_n5892# 0.010408f
C154 source.n120 a_n1094_n5892# 0.009829f
C155 source.n121 a_n1094_n5892# 0.018292f
C156 source.n122 a_n1094_n5892# 0.018292f
C157 source.n123 a_n1094_n5892# 0.009829f
C158 source.n124 a_n1094_n5892# 0.010408f
C159 source.n125 a_n1094_n5892# 0.023233f
C160 source.n126 a_n1094_n5892# 0.023233f
C161 source.n127 a_n1094_n5892# 0.010408f
C162 source.n128 a_n1094_n5892# 0.009829f
C163 source.n129 a_n1094_n5892# 0.018292f
C164 source.n130 a_n1094_n5892# 0.018292f
C165 source.n131 a_n1094_n5892# 0.009829f
C166 source.n132 a_n1094_n5892# 0.010408f
C167 source.n133 a_n1094_n5892# 0.023233f
C168 source.n134 a_n1094_n5892# 0.049423f
C169 source.n135 a_n1094_n5892# 0.010408f
C170 source.n136 a_n1094_n5892# 0.009829f
C171 source.n137 a_n1094_n5892# 0.040283f
C172 source.n138 a_n1094_n5892# 0.027502f
C173 source.n139 a_n1094_n5892# 1.43874f
C174 source.n140 a_n1094_n5892# 0.025218f
C175 source.n141 a_n1094_n5892# 0.018292f
C176 source.n142 a_n1094_n5892# 0.009829f
C177 source.n143 a_n1094_n5892# 0.023233f
C178 source.n144 a_n1094_n5892# 0.010408f
C179 source.n145 a_n1094_n5892# 0.018292f
C180 source.n146 a_n1094_n5892# 0.009829f
C181 source.n147 a_n1094_n5892# 0.023233f
C182 source.n148 a_n1094_n5892# 0.010408f
C183 source.n149 a_n1094_n5892# 0.018292f
C184 source.n150 a_n1094_n5892# 0.009829f
C185 source.n151 a_n1094_n5892# 0.023233f
C186 source.n152 a_n1094_n5892# 0.010408f
C187 source.n153 a_n1094_n5892# 0.018292f
C188 source.n154 a_n1094_n5892# 0.009829f
C189 source.n155 a_n1094_n5892# 0.023233f
C190 source.n156 a_n1094_n5892# 0.023233f
C191 source.n157 a_n1094_n5892# 0.010408f
C192 source.n158 a_n1094_n5892# 0.018292f
C193 source.n159 a_n1094_n5892# 0.009829f
C194 source.n160 a_n1094_n5892# 0.023233f
C195 source.n161 a_n1094_n5892# 0.010408f
C196 source.n162 a_n1094_n5892# 0.018292f
C197 source.n163 a_n1094_n5892# 0.009829f
C198 source.n164 a_n1094_n5892# 0.023233f
C199 source.n165 a_n1094_n5892# 0.010408f
C200 source.n166 a_n1094_n5892# 0.018292f
C201 source.n167 a_n1094_n5892# 0.009829f
C202 source.n168 a_n1094_n5892# 0.023233f
C203 source.n169 a_n1094_n5892# 0.010408f
C204 source.n170 a_n1094_n5892# 0.018292f
C205 source.n171 a_n1094_n5892# 0.009829f
C206 source.n172 a_n1094_n5892# 0.023233f
C207 source.n173 a_n1094_n5892# 0.010408f
C208 source.n174 a_n1094_n5892# 0.018292f
C209 source.n175 a_n1094_n5892# 0.010119f
C210 source.n176 a_n1094_n5892# 0.023233f
C211 source.n177 a_n1094_n5892# 0.009829f
C212 source.n178 a_n1094_n5892# 0.010408f
C213 source.n179 a_n1094_n5892# 0.018292f
C214 source.n180 a_n1094_n5892# 0.009829f
C215 source.n181 a_n1094_n5892# 0.023233f
C216 source.n182 a_n1094_n5892# 0.010408f
C217 source.n183 a_n1094_n5892# 0.018292f
C218 source.n184 a_n1094_n5892# 0.009829f
C219 source.n185 a_n1094_n5892# 0.017425f
C220 source.n186 a_n1094_n5892# 0.016424f
C221 source.t1 a_n1094_n5892# 0.04052f
C222 source.n187 a_n1094_n5892# 0.223181f
C223 source.n188 a_n1094_n5892# 1.98052f
C224 source.n189 a_n1094_n5892# 0.009829f
C225 source.n190 a_n1094_n5892# 0.010408f
C226 source.n191 a_n1094_n5892# 0.023233f
C227 source.n192 a_n1094_n5892# 0.023233f
C228 source.n193 a_n1094_n5892# 0.010408f
C229 source.n194 a_n1094_n5892# 0.009829f
C230 source.n195 a_n1094_n5892# 0.018292f
C231 source.n196 a_n1094_n5892# 0.018292f
C232 source.n197 a_n1094_n5892# 0.009829f
C233 source.n198 a_n1094_n5892# 0.010408f
C234 source.n199 a_n1094_n5892# 0.023233f
C235 source.n200 a_n1094_n5892# 0.023233f
C236 source.n201 a_n1094_n5892# 0.010408f
C237 source.n202 a_n1094_n5892# 0.009829f
C238 source.n203 a_n1094_n5892# 0.018292f
C239 source.n204 a_n1094_n5892# 0.018292f
C240 source.n205 a_n1094_n5892# 0.009829f
C241 source.n206 a_n1094_n5892# 0.010408f
C242 source.n207 a_n1094_n5892# 0.023233f
C243 source.n208 a_n1094_n5892# 0.023233f
C244 source.n209 a_n1094_n5892# 0.023233f
C245 source.n210 a_n1094_n5892# 0.010119f
C246 source.n211 a_n1094_n5892# 0.009829f
C247 source.n212 a_n1094_n5892# 0.018292f
C248 source.n213 a_n1094_n5892# 0.018292f
C249 source.n214 a_n1094_n5892# 0.009829f
C250 source.n215 a_n1094_n5892# 0.010408f
C251 source.n216 a_n1094_n5892# 0.023233f
C252 source.n217 a_n1094_n5892# 0.023233f
C253 source.n218 a_n1094_n5892# 0.010408f
C254 source.n219 a_n1094_n5892# 0.009829f
C255 source.n220 a_n1094_n5892# 0.018292f
C256 source.n221 a_n1094_n5892# 0.018292f
C257 source.n222 a_n1094_n5892# 0.009829f
C258 source.n223 a_n1094_n5892# 0.010408f
C259 source.n224 a_n1094_n5892# 0.023233f
C260 source.n225 a_n1094_n5892# 0.023233f
C261 source.n226 a_n1094_n5892# 0.010408f
C262 source.n227 a_n1094_n5892# 0.009829f
C263 source.n228 a_n1094_n5892# 0.018292f
C264 source.n229 a_n1094_n5892# 0.018292f
C265 source.n230 a_n1094_n5892# 0.009829f
C266 source.n231 a_n1094_n5892# 0.010408f
C267 source.n232 a_n1094_n5892# 0.023233f
C268 source.n233 a_n1094_n5892# 0.023233f
C269 source.n234 a_n1094_n5892# 0.010408f
C270 source.n235 a_n1094_n5892# 0.009829f
C271 source.n236 a_n1094_n5892# 0.018292f
C272 source.n237 a_n1094_n5892# 0.018292f
C273 source.n238 a_n1094_n5892# 0.009829f
C274 source.n239 a_n1094_n5892# 0.010408f
C275 source.n240 a_n1094_n5892# 0.023233f
C276 source.n241 a_n1094_n5892# 0.023233f
C277 source.n242 a_n1094_n5892# 0.010408f
C278 source.n243 a_n1094_n5892# 0.009829f
C279 source.n244 a_n1094_n5892# 0.018292f
C280 source.n245 a_n1094_n5892# 0.018292f
C281 source.n246 a_n1094_n5892# 0.009829f
C282 source.n247 a_n1094_n5892# 0.010408f
C283 source.n248 a_n1094_n5892# 0.023233f
C284 source.n249 a_n1094_n5892# 0.023233f
C285 source.n250 a_n1094_n5892# 0.010408f
C286 source.n251 a_n1094_n5892# 0.009829f
C287 source.n252 a_n1094_n5892# 0.018292f
C288 source.n253 a_n1094_n5892# 0.018292f
C289 source.n254 a_n1094_n5892# 0.009829f
C290 source.n255 a_n1094_n5892# 0.010119f
C291 source.n256 a_n1094_n5892# 0.010119f
C292 source.n257 a_n1094_n5892# 0.023233f
C293 source.n258 a_n1094_n5892# 0.023233f
C294 source.n259 a_n1094_n5892# 0.010408f
C295 source.n260 a_n1094_n5892# 0.009829f
C296 source.n261 a_n1094_n5892# 0.018292f
C297 source.n262 a_n1094_n5892# 0.018292f
C298 source.n263 a_n1094_n5892# 0.009829f
C299 source.n264 a_n1094_n5892# 0.010408f
C300 source.n265 a_n1094_n5892# 0.023233f
C301 source.n266 a_n1094_n5892# 0.023233f
C302 source.n267 a_n1094_n5892# 0.010408f
C303 source.n268 a_n1094_n5892# 0.009829f
C304 source.n269 a_n1094_n5892# 0.018292f
C305 source.n270 a_n1094_n5892# 0.018292f
C306 source.n271 a_n1094_n5892# 0.009829f
C307 source.n272 a_n1094_n5892# 0.010408f
C308 source.n273 a_n1094_n5892# 0.023233f
C309 source.n274 a_n1094_n5892# 0.049423f
C310 source.n275 a_n1094_n5892# 0.010408f
C311 source.n276 a_n1094_n5892# 0.009829f
C312 source.n277 a_n1094_n5892# 0.040283f
C313 source.n278 a_n1094_n5892# 0.027502f
C314 source.n279 a_n1094_n5892# 0.0742f
C315 source.n280 a_n1094_n5892# 0.025218f
C316 source.n281 a_n1094_n5892# 0.018292f
C317 source.n282 a_n1094_n5892# 0.009829f
C318 source.n283 a_n1094_n5892# 0.023233f
C319 source.n284 a_n1094_n5892# 0.010408f
C320 source.n285 a_n1094_n5892# 0.018292f
C321 source.n286 a_n1094_n5892# 0.009829f
C322 source.n287 a_n1094_n5892# 0.023233f
C323 source.n288 a_n1094_n5892# 0.010408f
C324 source.n289 a_n1094_n5892# 0.018292f
C325 source.n290 a_n1094_n5892# 0.009829f
C326 source.n291 a_n1094_n5892# 0.023233f
C327 source.n292 a_n1094_n5892# 0.010408f
C328 source.n293 a_n1094_n5892# 0.018292f
C329 source.n294 a_n1094_n5892# 0.009829f
C330 source.n295 a_n1094_n5892# 0.023233f
C331 source.n296 a_n1094_n5892# 0.023233f
C332 source.n297 a_n1094_n5892# 0.010408f
C333 source.n298 a_n1094_n5892# 0.018292f
C334 source.n299 a_n1094_n5892# 0.009829f
C335 source.n300 a_n1094_n5892# 0.023233f
C336 source.n301 a_n1094_n5892# 0.010408f
C337 source.n302 a_n1094_n5892# 0.018292f
C338 source.n303 a_n1094_n5892# 0.009829f
C339 source.n304 a_n1094_n5892# 0.023233f
C340 source.n305 a_n1094_n5892# 0.010408f
C341 source.n306 a_n1094_n5892# 0.018292f
C342 source.n307 a_n1094_n5892# 0.009829f
C343 source.n308 a_n1094_n5892# 0.023233f
C344 source.n309 a_n1094_n5892# 0.010408f
C345 source.n310 a_n1094_n5892# 0.018292f
C346 source.n311 a_n1094_n5892# 0.009829f
C347 source.n312 a_n1094_n5892# 0.023233f
C348 source.n313 a_n1094_n5892# 0.010408f
C349 source.n314 a_n1094_n5892# 0.018292f
C350 source.n315 a_n1094_n5892# 0.010119f
C351 source.n316 a_n1094_n5892# 0.023233f
C352 source.n317 a_n1094_n5892# 0.009829f
C353 source.n318 a_n1094_n5892# 0.010408f
C354 source.n319 a_n1094_n5892# 0.018292f
C355 source.n320 a_n1094_n5892# 0.009829f
C356 source.n321 a_n1094_n5892# 0.023233f
C357 source.n322 a_n1094_n5892# 0.010408f
C358 source.n323 a_n1094_n5892# 0.018292f
C359 source.n324 a_n1094_n5892# 0.009829f
C360 source.n325 a_n1094_n5892# 0.017425f
C361 source.n326 a_n1094_n5892# 0.016424f
C362 source.t6 a_n1094_n5892# 0.04052f
C363 source.n327 a_n1094_n5892# 0.223181f
C364 source.n328 a_n1094_n5892# 1.98052f
C365 source.n329 a_n1094_n5892# 0.009829f
C366 source.n330 a_n1094_n5892# 0.010408f
C367 source.n331 a_n1094_n5892# 0.023233f
C368 source.n332 a_n1094_n5892# 0.023233f
C369 source.n333 a_n1094_n5892# 0.010408f
C370 source.n334 a_n1094_n5892# 0.009829f
C371 source.n335 a_n1094_n5892# 0.018292f
C372 source.n336 a_n1094_n5892# 0.018292f
C373 source.n337 a_n1094_n5892# 0.009829f
C374 source.n338 a_n1094_n5892# 0.010408f
C375 source.n339 a_n1094_n5892# 0.023233f
C376 source.n340 a_n1094_n5892# 0.023233f
C377 source.n341 a_n1094_n5892# 0.010408f
C378 source.n342 a_n1094_n5892# 0.009829f
C379 source.n343 a_n1094_n5892# 0.018292f
C380 source.n344 a_n1094_n5892# 0.018292f
C381 source.n345 a_n1094_n5892# 0.009829f
C382 source.n346 a_n1094_n5892# 0.010408f
C383 source.n347 a_n1094_n5892# 0.023233f
C384 source.n348 a_n1094_n5892# 0.023233f
C385 source.n349 a_n1094_n5892# 0.023233f
C386 source.n350 a_n1094_n5892# 0.010119f
C387 source.n351 a_n1094_n5892# 0.009829f
C388 source.n352 a_n1094_n5892# 0.018292f
C389 source.n353 a_n1094_n5892# 0.018292f
C390 source.n354 a_n1094_n5892# 0.009829f
C391 source.n355 a_n1094_n5892# 0.010408f
C392 source.n356 a_n1094_n5892# 0.023233f
C393 source.n357 a_n1094_n5892# 0.023233f
C394 source.n358 a_n1094_n5892# 0.010408f
C395 source.n359 a_n1094_n5892# 0.009829f
C396 source.n360 a_n1094_n5892# 0.018292f
C397 source.n361 a_n1094_n5892# 0.018292f
C398 source.n362 a_n1094_n5892# 0.009829f
C399 source.n363 a_n1094_n5892# 0.010408f
C400 source.n364 a_n1094_n5892# 0.023233f
C401 source.n365 a_n1094_n5892# 0.023233f
C402 source.n366 a_n1094_n5892# 0.010408f
C403 source.n367 a_n1094_n5892# 0.009829f
C404 source.n368 a_n1094_n5892# 0.018292f
C405 source.n369 a_n1094_n5892# 0.018292f
C406 source.n370 a_n1094_n5892# 0.009829f
C407 source.n371 a_n1094_n5892# 0.010408f
C408 source.n372 a_n1094_n5892# 0.023233f
C409 source.n373 a_n1094_n5892# 0.023233f
C410 source.n374 a_n1094_n5892# 0.010408f
C411 source.n375 a_n1094_n5892# 0.009829f
C412 source.n376 a_n1094_n5892# 0.018292f
C413 source.n377 a_n1094_n5892# 0.018292f
C414 source.n378 a_n1094_n5892# 0.009829f
C415 source.n379 a_n1094_n5892# 0.010408f
C416 source.n380 a_n1094_n5892# 0.023233f
C417 source.n381 a_n1094_n5892# 0.023233f
C418 source.n382 a_n1094_n5892# 0.010408f
C419 source.n383 a_n1094_n5892# 0.009829f
C420 source.n384 a_n1094_n5892# 0.018292f
C421 source.n385 a_n1094_n5892# 0.018292f
C422 source.n386 a_n1094_n5892# 0.009829f
C423 source.n387 a_n1094_n5892# 0.010408f
C424 source.n388 a_n1094_n5892# 0.023233f
C425 source.n389 a_n1094_n5892# 0.023233f
C426 source.n390 a_n1094_n5892# 0.010408f
C427 source.n391 a_n1094_n5892# 0.009829f
C428 source.n392 a_n1094_n5892# 0.018292f
C429 source.n393 a_n1094_n5892# 0.018292f
C430 source.n394 a_n1094_n5892# 0.009829f
C431 source.n395 a_n1094_n5892# 0.010119f
C432 source.n396 a_n1094_n5892# 0.010119f
C433 source.n397 a_n1094_n5892# 0.023233f
C434 source.n398 a_n1094_n5892# 0.023233f
C435 source.n399 a_n1094_n5892# 0.010408f
C436 source.n400 a_n1094_n5892# 0.009829f
C437 source.n401 a_n1094_n5892# 0.018292f
C438 source.n402 a_n1094_n5892# 0.018292f
C439 source.n403 a_n1094_n5892# 0.009829f
C440 source.n404 a_n1094_n5892# 0.010408f
C441 source.n405 a_n1094_n5892# 0.023233f
C442 source.n406 a_n1094_n5892# 0.023233f
C443 source.n407 a_n1094_n5892# 0.010408f
C444 source.n408 a_n1094_n5892# 0.009829f
C445 source.n409 a_n1094_n5892# 0.018292f
C446 source.n410 a_n1094_n5892# 0.018292f
C447 source.n411 a_n1094_n5892# 0.009829f
C448 source.n412 a_n1094_n5892# 0.010408f
C449 source.n413 a_n1094_n5892# 0.023233f
C450 source.n414 a_n1094_n5892# 0.049423f
C451 source.n415 a_n1094_n5892# 0.010408f
C452 source.n416 a_n1094_n5892# 0.009829f
C453 source.n417 a_n1094_n5892# 0.040283f
C454 source.n418 a_n1094_n5892# 0.027502f
C455 source.n419 a_n1094_n5892# 0.0742f
C456 source.n420 a_n1094_n5892# 0.025218f
C457 source.n421 a_n1094_n5892# 0.018292f
C458 source.n422 a_n1094_n5892# 0.009829f
C459 source.n423 a_n1094_n5892# 0.023233f
C460 source.n424 a_n1094_n5892# 0.010408f
C461 source.n425 a_n1094_n5892# 0.018292f
C462 source.n426 a_n1094_n5892# 0.009829f
C463 source.n427 a_n1094_n5892# 0.023233f
C464 source.n428 a_n1094_n5892# 0.010408f
C465 source.n429 a_n1094_n5892# 0.018292f
C466 source.n430 a_n1094_n5892# 0.009829f
C467 source.n431 a_n1094_n5892# 0.023233f
C468 source.n432 a_n1094_n5892# 0.010408f
C469 source.n433 a_n1094_n5892# 0.018292f
C470 source.n434 a_n1094_n5892# 0.009829f
C471 source.n435 a_n1094_n5892# 0.023233f
C472 source.n436 a_n1094_n5892# 0.023233f
C473 source.n437 a_n1094_n5892# 0.010408f
C474 source.n438 a_n1094_n5892# 0.018292f
C475 source.n439 a_n1094_n5892# 0.009829f
C476 source.n440 a_n1094_n5892# 0.023233f
C477 source.n441 a_n1094_n5892# 0.010408f
C478 source.n442 a_n1094_n5892# 0.018292f
C479 source.n443 a_n1094_n5892# 0.009829f
C480 source.n444 a_n1094_n5892# 0.023233f
C481 source.n445 a_n1094_n5892# 0.010408f
C482 source.n446 a_n1094_n5892# 0.018292f
C483 source.n447 a_n1094_n5892# 0.009829f
C484 source.n448 a_n1094_n5892# 0.023233f
C485 source.n449 a_n1094_n5892# 0.010408f
C486 source.n450 a_n1094_n5892# 0.018292f
C487 source.n451 a_n1094_n5892# 0.009829f
C488 source.n452 a_n1094_n5892# 0.023233f
C489 source.n453 a_n1094_n5892# 0.010408f
C490 source.n454 a_n1094_n5892# 0.018292f
C491 source.n455 a_n1094_n5892# 0.010119f
C492 source.n456 a_n1094_n5892# 0.023233f
C493 source.n457 a_n1094_n5892# 0.009829f
C494 source.n458 a_n1094_n5892# 0.010408f
C495 source.n459 a_n1094_n5892# 0.018292f
C496 source.n460 a_n1094_n5892# 0.009829f
C497 source.n461 a_n1094_n5892# 0.023233f
C498 source.n462 a_n1094_n5892# 0.010408f
C499 source.n463 a_n1094_n5892# 0.018292f
C500 source.n464 a_n1094_n5892# 0.009829f
C501 source.n465 a_n1094_n5892# 0.017425f
C502 source.n466 a_n1094_n5892# 0.016424f
C503 source.t5 a_n1094_n5892# 0.04052f
C504 source.n467 a_n1094_n5892# 0.223181f
C505 source.n468 a_n1094_n5892# 1.98052f
C506 source.n469 a_n1094_n5892# 0.009829f
C507 source.n470 a_n1094_n5892# 0.010408f
C508 source.n471 a_n1094_n5892# 0.023233f
C509 source.n472 a_n1094_n5892# 0.023233f
C510 source.n473 a_n1094_n5892# 0.010408f
C511 source.n474 a_n1094_n5892# 0.009829f
C512 source.n475 a_n1094_n5892# 0.018292f
C513 source.n476 a_n1094_n5892# 0.018292f
C514 source.n477 a_n1094_n5892# 0.009829f
C515 source.n478 a_n1094_n5892# 0.010408f
C516 source.n479 a_n1094_n5892# 0.023233f
C517 source.n480 a_n1094_n5892# 0.023233f
C518 source.n481 a_n1094_n5892# 0.010408f
C519 source.n482 a_n1094_n5892# 0.009829f
C520 source.n483 a_n1094_n5892# 0.018292f
C521 source.n484 a_n1094_n5892# 0.018292f
C522 source.n485 a_n1094_n5892# 0.009829f
C523 source.n486 a_n1094_n5892# 0.010408f
C524 source.n487 a_n1094_n5892# 0.023233f
C525 source.n488 a_n1094_n5892# 0.023233f
C526 source.n489 a_n1094_n5892# 0.023233f
C527 source.n490 a_n1094_n5892# 0.010119f
C528 source.n491 a_n1094_n5892# 0.009829f
C529 source.n492 a_n1094_n5892# 0.018292f
C530 source.n493 a_n1094_n5892# 0.018292f
C531 source.n494 a_n1094_n5892# 0.009829f
C532 source.n495 a_n1094_n5892# 0.010408f
C533 source.n496 a_n1094_n5892# 0.023233f
C534 source.n497 a_n1094_n5892# 0.023233f
C535 source.n498 a_n1094_n5892# 0.010408f
C536 source.n499 a_n1094_n5892# 0.009829f
C537 source.n500 a_n1094_n5892# 0.018292f
C538 source.n501 a_n1094_n5892# 0.018292f
C539 source.n502 a_n1094_n5892# 0.009829f
C540 source.n503 a_n1094_n5892# 0.010408f
C541 source.n504 a_n1094_n5892# 0.023233f
C542 source.n505 a_n1094_n5892# 0.023233f
C543 source.n506 a_n1094_n5892# 0.010408f
C544 source.n507 a_n1094_n5892# 0.009829f
C545 source.n508 a_n1094_n5892# 0.018292f
C546 source.n509 a_n1094_n5892# 0.018292f
C547 source.n510 a_n1094_n5892# 0.009829f
C548 source.n511 a_n1094_n5892# 0.010408f
C549 source.n512 a_n1094_n5892# 0.023233f
C550 source.n513 a_n1094_n5892# 0.023233f
C551 source.n514 a_n1094_n5892# 0.010408f
C552 source.n515 a_n1094_n5892# 0.009829f
C553 source.n516 a_n1094_n5892# 0.018292f
C554 source.n517 a_n1094_n5892# 0.018292f
C555 source.n518 a_n1094_n5892# 0.009829f
C556 source.n519 a_n1094_n5892# 0.010408f
C557 source.n520 a_n1094_n5892# 0.023233f
C558 source.n521 a_n1094_n5892# 0.023233f
C559 source.n522 a_n1094_n5892# 0.010408f
C560 source.n523 a_n1094_n5892# 0.009829f
C561 source.n524 a_n1094_n5892# 0.018292f
C562 source.n525 a_n1094_n5892# 0.018292f
C563 source.n526 a_n1094_n5892# 0.009829f
C564 source.n527 a_n1094_n5892# 0.010408f
C565 source.n528 a_n1094_n5892# 0.023233f
C566 source.n529 a_n1094_n5892# 0.023233f
C567 source.n530 a_n1094_n5892# 0.010408f
C568 source.n531 a_n1094_n5892# 0.009829f
C569 source.n532 a_n1094_n5892# 0.018292f
C570 source.n533 a_n1094_n5892# 0.018292f
C571 source.n534 a_n1094_n5892# 0.009829f
C572 source.n535 a_n1094_n5892# 0.010119f
C573 source.n536 a_n1094_n5892# 0.010119f
C574 source.n537 a_n1094_n5892# 0.023233f
C575 source.n538 a_n1094_n5892# 0.023233f
C576 source.n539 a_n1094_n5892# 0.010408f
C577 source.n540 a_n1094_n5892# 0.009829f
C578 source.n541 a_n1094_n5892# 0.018292f
C579 source.n542 a_n1094_n5892# 0.018292f
C580 source.n543 a_n1094_n5892# 0.009829f
C581 source.n544 a_n1094_n5892# 0.010408f
C582 source.n545 a_n1094_n5892# 0.023233f
C583 source.n546 a_n1094_n5892# 0.023233f
C584 source.n547 a_n1094_n5892# 0.010408f
C585 source.n548 a_n1094_n5892# 0.009829f
C586 source.n549 a_n1094_n5892# 0.018292f
C587 source.n550 a_n1094_n5892# 0.018292f
C588 source.n551 a_n1094_n5892# 0.009829f
C589 source.n552 a_n1094_n5892# 0.010408f
C590 source.n553 a_n1094_n5892# 0.023233f
C591 source.n554 a_n1094_n5892# 0.049423f
C592 source.n555 a_n1094_n5892# 0.010408f
C593 source.n556 a_n1094_n5892# 0.009829f
C594 source.n557 a_n1094_n5892# 0.040283f
C595 source.n558 a_n1094_n5892# 0.027502f
C596 source.n559 a_n1094_n5892# 1.77719f
C597 source.n560 a_n1094_n5892# 0.025218f
C598 source.n561 a_n1094_n5892# 0.018292f
C599 source.n562 a_n1094_n5892# 0.009829f
C600 source.n563 a_n1094_n5892# 0.023233f
C601 source.n564 a_n1094_n5892# 0.010408f
C602 source.n565 a_n1094_n5892# 0.018292f
C603 source.n566 a_n1094_n5892# 0.009829f
C604 source.n567 a_n1094_n5892# 0.023233f
C605 source.n568 a_n1094_n5892# 0.010408f
C606 source.n569 a_n1094_n5892# 0.018292f
C607 source.n570 a_n1094_n5892# 0.009829f
C608 source.n571 a_n1094_n5892# 0.023233f
C609 source.n572 a_n1094_n5892# 0.010408f
C610 source.n573 a_n1094_n5892# 0.018292f
C611 source.n574 a_n1094_n5892# 0.009829f
C612 source.n575 a_n1094_n5892# 0.023233f
C613 source.n576 a_n1094_n5892# 0.010408f
C614 source.n577 a_n1094_n5892# 0.018292f
C615 source.n578 a_n1094_n5892# 0.009829f
C616 source.n579 a_n1094_n5892# 0.023233f
C617 source.n580 a_n1094_n5892# 0.010408f
C618 source.n581 a_n1094_n5892# 0.018292f
C619 source.n582 a_n1094_n5892# 0.009829f
C620 source.n583 a_n1094_n5892# 0.023233f
C621 source.n584 a_n1094_n5892# 0.010408f
C622 source.n585 a_n1094_n5892# 0.018292f
C623 source.n586 a_n1094_n5892# 0.009829f
C624 source.n587 a_n1094_n5892# 0.023233f
C625 source.n588 a_n1094_n5892# 0.010408f
C626 source.n589 a_n1094_n5892# 0.018292f
C627 source.n590 a_n1094_n5892# 0.009829f
C628 source.n591 a_n1094_n5892# 0.023233f
C629 source.n592 a_n1094_n5892# 0.010408f
C630 source.n593 a_n1094_n5892# 0.018292f
C631 source.n594 a_n1094_n5892# 0.010119f
C632 source.n595 a_n1094_n5892# 0.023233f
C633 source.n596 a_n1094_n5892# 0.010408f
C634 source.n597 a_n1094_n5892# 0.018292f
C635 source.n598 a_n1094_n5892# 0.009829f
C636 source.n599 a_n1094_n5892# 0.023233f
C637 source.n600 a_n1094_n5892# 0.010408f
C638 source.n601 a_n1094_n5892# 0.018292f
C639 source.n602 a_n1094_n5892# 0.009829f
C640 source.n603 a_n1094_n5892# 0.017425f
C641 source.n604 a_n1094_n5892# 0.016424f
C642 source.t3 a_n1094_n5892# 0.04052f
C643 source.n605 a_n1094_n5892# 0.223181f
C644 source.n606 a_n1094_n5892# 1.98052f
C645 source.n607 a_n1094_n5892# 0.009829f
C646 source.n608 a_n1094_n5892# 0.010408f
C647 source.n609 a_n1094_n5892# 0.023233f
C648 source.n610 a_n1094_n5892# 0.023233f
C649 source.n611 a_n1094_n5892# 0.010408f
C650 source.n612 a_n1094_n5892# 0.009829f
C651 source.n613 a_n1094_n5892# 0.018292f
C652 source.n614 a_n1094_n5892# 0.018292f
C653 source.n615 a_n1094_n5892# 0.009829f
C654 source.n616 a_n1094_n5892# 0.010408f
C655 source.n617 a_n1094_n5892# 0.023233f
C656 source.n618 a_n1094_n5892# 0.023233f
C657 source.n619 a_n1094_n5892# 0.010408f
C658 source.n620 a_n1094_n5892# 0.009829f
C659 source.n621 a_n1094_n5892# 0.018292f
C660 source.n622 a_n1094_n5892# 0.018292f
C661 source.n623 a_n1094_n5892# 0.009829f
C662 source.n624 a_n1094_n5892# 0.009829f
C663 source.n625 a_n1094_n5892# 0.010408f
C664 source.n626 a_n1094_n5892# 0.023233f
C665 source.n627 a_n1094_n5892# 0.023233f
C666 source.n628 a_n1094_n5892# 0.023233f
C667 source.n629 a_n1094_n5892# 0.010119f
C668 source.n630 a_n1094_n5892# 0.009829f
C669 source.n631 a_n1094_n5892# 0.018292f
C670 source.n632 a_n1094_n5892# 0.018292f
C671 source.n633 a_n1094_n5892# 0.009829f
C672 source.n634 a_n1094_n5892# 0.010408f
C673 source.n635 a_n1094_n5892# 0.023233f
C674 source.n636 a_n1094_n5892# 0.023233f
C675 source.n637 a_n1094_n5892# 0.010408f
C676 source.n638 a_n1094_n5892# 0.009829f
C677 source.n639 a_n1094_n5892# 0.018292f
C678 source.n640 a_n1094_n5892# 0.018292f
C679 source.n641 a_n1094_n5892# 0.009829f
C680 source.n642 a_n1094_n5892# 0.010408f
C681 source.n643 a_n1094_n5892# 0.023233f
C682 source.n644 a_n1094_n5892# 0.023233f
C683 source.n645 a_n1094_n5892# 0.010408f
C684 source.n646 a_n1094_n5892# 0.009829f
C685 source.n647 a_n1094_n5892# 0.018292f
C686 source.n648 a_n1094_n5892# 0.018292f
C687 source.n649 a_n1094_n5892# 0.009829f
C688 source.n650 a_n1094_n5892# 0.010408f
C689 source.n651 a_n1094_n5892# 0.023233f
C690 source.n652 a_n1094_n5892# 0.023233f
C691 source.n653 a_n1094_n5892# 0.010408f
C692 source.n654 a_n1094_n5892# 0.009829f
C693 source.n655 a_n1094_n5892# 0.018292f
C694 source.n656 a_n1094_n5892# 0.018292f
C695 source.n657 a_n1094_n5892# 0.009829f
C696 source.n658 a_n1094_n5892# 0.010408f
C697 source.n659 a_n1094_n5892# 0.023233f
C698 source.n660 a_n1094_n5892# 0.023233f
C699 source.n661 a_n1094_n5892# 0.010408f
C700 source.n662 a_n1094_n5892# 0.009829f
C701 source.n663 a_n1094_n5892# 0.018292f
C702 source.n664 a_n1094_n5892# 0.018292f
C703 source.n665 a_n1094_n5892# 0.009829f
C704 source.n666 a_n1094_n5892# 0.010408f
C705 source.n667 a_n1094_n5892# 0.023233f
C706 source.n668 a_n1094_n5892# 0.023233f
C707 source.n669 a_n1094_n5892# 0.023233f
C708 source.n670 a_n1094_n5892# 0.010408f
C709 source.n671 a_n1094_n5892# 0.009829f
C710 source.n672 a_n1094_n5892# 0.018292f
C711 source.n673 a_n1094_n5892# 0.018292f
C712 source.n674 a_n1094_n5892# 0.009829f
C713 source.n675 a_n1094_n5892# 0.010119f
C714 source.n676 a_n1094_n5892# 0.010119f
C715 source.n677 a_n1094_n5892# 0.023233f
C716 source.n678 a_n1094_n5892# 0.023233f
C717 source.n679 a_n1094_n5892# 0.010408f
C718 source.n680 a_n1094_n5892# 0.009829f
C719 source.n681 a_n1094_n5892# 0.018292f
C720 source.n682 a_n1094_n5892# 0.018292f
C721 source.n683 a_n1094_n5892# 0.009829f
C722 source.n684 a_n1094_n5892# 0.010408f
C723 source.n685 a_n1094_n5892# 0.023233f
C724 source.n686 a_n1094_n5892# 0.023233f
C725 source.n687 a_n1094_n5892# 0.010408f
C726 source.n688 a_n1094_n5892# 0.009829f
C727 source.n689 a_n1094_n5892# 0.018292f
C728 source.n690 a_n1094_n5892# 0.018292f
C729 source.n691 a_n1094_n5892# 0.009829f
C730 source.n692 a_n1094_n5892# 0.010408f
C731 source.n693 a_n1094_n5892# 0.023233f
C732 source.n694 a_n1094_n5892# 0.049423f
C733 source.n695 a_n1094_n5892# 0.010408f
C734 source.n696 a_n1094_n5892# 0.009829f
C735 source.n697 a_n1094_n5892# 0.040283f
C736 source.n698 a_n1094_n5892# 0.027502f
C737 source.n699 a_n1094_n5892# 1.77719f
C738 source.n700 a_n1094_n5892# 0.025218f
C739 source.n701 a_n1094_n5892# 0.018292f
C740 source.n702 a_n1094_n5892# 0.009829f
C741 source.n703 a_n1094_n5892# 0.023233f
C742 source.n704 a_n1094_n5892# 0.010408f
C743 source.n705 a_n1094_n5892# 0.018292f
C744 source.n706 a_n1094_n5892# 0.009829f
C745 source.n707 a_n1094_n5892# 0.023233f
C746 source.n708 a_n1094_n5892# 0.010408f
C747 source.n709 a_n1094_n5892# 0.018292f
C748 source.n710 a_n1094_n5892# 0.009829f
C749 source.n711 a_n1094_n5892# 0.023233f
C750 source.n712 a_n1094_n5892# 0.010408f
C751 source.n713 a_n1094_n5892# 0.018292f
C752 source.n714 a_n1094_n5892# 0.009829f
C753 source.n715 a_n1094_n5892# 0.023233f
C754 source.n716 a_n1094_n5892# 0.010408f
C755 source.n717 a_n1094_n5892# 0.018292f
C756 source.n718 a_n1094_n5892# 0.009829f
C757 source.n719 a_n1094_n5892# 0.023233f
C758 source.n720 a_n1094_n5892# 0.010408f
C759 source.n721 a_n1094_n5892# 0.018292f
C760 source.n722 a_n1094_n5892# 0.009829f
C761 source.n723 a_n1094_n5892# 0.023233f
C762 source.n724 a_n1094_n5892# 0.010408f
C763 source.n725 a_n1094_n5892# 0.018292f
C764 source.n726 a_n1094_n5892# 0.009829f
C765 source.n727 a_n1094_n5892# 0.023233f
C766 source.n728 a_n1094_n5892# 0.010408f
C767 source.n729 a_n1094_n5892# 0.018292f
C768 source.n730 a_n1094_n5892# 0.009829f
C769 source.n731 a_n1094_n5892# 0.023233f
C770 source.n732 a_n1094_n5892# 0.010408f
C771 source.n733 a_n1094_n5892# 0.018292f
C772 source.n734 a_n1094_n5892# 0.010119f
C773 source.n735 a_n1094_n5892# 0.023233f
C774 source.n736 a_n1094_n5892# 0.010408f
C775 source.n737 a_n1094_n5892# 0.018292f
C776 source.n738 a_n1094_n5892# 0.009829f
C777 source.n739 a_n1094_n5892# 0.023233f
C778 source.n740 a_n1094_n5892# 0.010408f
C779 source.n741 a_n1094_n5892# 0.018292f
C780 source.n742 a_n1094_n5892# 0.009829f
C781 source.n743 a_n1094_n5892# 0.017425f
C782 source.n744 a_n1094_n5892# 0.016424f
C783 source.t0 a_n1094_n5892# 0.04052f
C784 source.n745 a_n1094_n5892# 0.223181f
C785 source.n746 a_n1094_n5892# 1.98052f
C786 source.n747 a_n1094_n5892# 0.009829f
C787 source.n748 a_n1094_n5892# 0.010408f
C788 source.n749 a_n1094_n5892# 0.023233f
C789 source.n750 a_n1094_n5892# 0.023233f
C790 source.n751 a_n1094_n5892# 0.010408f
C791 source.n752 a_n1094_n5892# 0.009829f
C792 source.n753 a_n1094_n5892# 0.018292f
C793 source.n754 a_n1094_n5892# 0.018292f
C794 source.n755 a_n1094_n5892# 0.009829f
C795 source.n756 a_n1094_n5892# 0.010408f
C796 source.n757 a_n1094_n5892# 0.023233f
C797 source.n758 a_n1094_n5892# 0.023233f
C798 source.n759 a_n1094_n5892# 0.010408f
C799 source.n760 a_n1094_n5892# 0.009829f
C800 source.n761 a_n1094_n5892# 0.018292f
C801 source.n762 a_n1094_n5892# 0.018292f
C802 source.n763 a_n1094_n5892# 0.009829f
C803 source.n764 a_n1094_n5892# 0.009829f
C804 source.n765 a_n1094_n5892# 0.010408f
C805 source.n766 a_n1094_n5892# 0.023233f
C806 source.n767 a_n1094_n5892# 0.023233f
C807 source.n768 a_n1094_n5892# 0.023233f
C808 source.n769 a_n1094_n5892# 0.010119f
C809 source.n770 a_n1094_n5892# 0.009829f
C810 source.n771 a_n1094_n5892# 0.018292f
C811 source.n772 a_n1094_n5892# 0.018292f
C812 source.n773 a_n1094_n5892# 0.009829f
C813 source.n774 a_n1094_n5892# 0.010408f
C814 source.n775 a_n1094_n5892# 0.023233f
C815 source.n776 a_n1094_n5892# 0.023233f
C816 source.n777 a_n1094_n5892# 0.010408f
C817 source.n778 a_n1094_n5892# 0.009829f
C818 source.n779 a_n1094_n5892# 0.018292f
C819 source.n780 a_n1094_n5892# 0.018292f
C820 source.n781 a_n1094_n5892# 0.009829f
C821 source.n782 a_n1094_n5892# 0.010408f
C822 source.n783 a_n1094_n5892# 0.023233f
C823 source.n784 a_n1094_n5892# 0.023233f
C824 source.n785 a_n1094_n5892# 0.010408f
C825 source.n786 a_n1094_n5892# 0.009829f
C826 source.n787 a_n1094_n5892# 0.018292f
C827 source.n788 a_n1094_n5892# 0.018292f
C828 source.n789 a_n1094_n5892# 0.009829f
C829 source.n790 a_n1094_n5892# 0.010408f
C830 source.n791 a_n1094_n5892# 0.023233f
C831 source.n792 a_n1094_n5892# 0.023233f
C832 source.n793 a_n1094_n5892# 0.010408f
C833 source.n794 a_n1094_n5892# 0.009829f
C834 source.n795 a_n1094_n5892# 0.018292f
C835 source.n796 a_n1094_n5892# 0.018292f
C836 source.n797 a_n1094_n5892# 0.009829f
C837 source.n798 a_n1094_n5892# 0.010408f
C838 source.n799 a_n1094_n5892# 0.023233f
C839 source.n800 a_n1094_n5892# 0.023233f
C840 source.n801 a_n1094_n5892# 0.010408f
C841 source.n802 a_n1094_n5892# 0.009829f
C842 source.n803 a_n1094_n5892# 0.018292f
C843 source.n804 a_n1094_n5892# 0.018292f
C844 source.n805 a_n1094_n5892# 0.009829f
C845 source.n806 a_n1094_n5892# 0.010408f
C846 source.n807 a_n1094_n5892# 0.023233f
C847 source.n808 a_n1094_n5892# 0.023233f
C848 source.n809 a_n1094_n5892# 0.023233f
C849 source.n810 a_n1094_n5892# 0.010408f
C850 source.n811 a_n1094_n5892# 0.009829f
C851 source.n812 a_n1094_n5892# 0.018292f
C852 source.n813 a_n1094_n5892# 0.018292f
C853 source.n814 a_n1094_n5892# 0.009829f
C854 source.n815 a_n1094_n5892# 0.010119f
C855 source.n816 a_n1094_n5892# 0.010119f
C856 source.n817 a_n1094_n5892# 0.023233f
C857 source.n818 a_n1094_n5892# 0.023233f
C858 source.n819 a_n1094_n5892# 0.010408f
C859 source.n820 a_n1094_n5892# 0.009829f
C860 source.n821 a_n1094_n5892# 0.018292f
C861 source.n822 a_n1094_n5892# 0.018292f
C862 source.n823 a_n1094_n5892# 0.009829f
C863 source.n824 a_n1094_n5892# 0.010408f
C864 source.n825 a_n1094_n5892# 0.023233f
C865 source.n826 a_n1094_n5892# 0.023233f
C866 source.n827 a_n1094_n5892# 0.010408f
C867 source.n828 a_n1094_n5892# 0.009829f
C868 source.n829 a_n1094_n5892# 0.018292f
C869 source.n830 a_n1094_n5892# 0.018292f
C870 source.n831 a_n1094_n5892# 0.009829f
C871 source.n832 a_n1094_n5892# 0.010408f
C872 source.n833 a_n1094_n5892# 0.023233f
C873 source.n834 a_n1094_n5892# 0.049423f
C874 source.n835 a_n1094_n5892# 0.010408f
C875 source.n836 a_n1094_n5892# 0.009829f
C876 source.n837 a_n1094_n5892# 0.040283f
C877 source.n838 a_n1094_n5892# 0.027502f
C878 source.n839 a_n1094_n5892# 0.0742f
C879 source.n840 a_n1094_n5892# 0.025218f
C880 source.n841 a_n1094_n5892# 0.018292f
C881 source.n842 a_n1094_n5892# 0.009829f
C882 source.n843 a_n1094_n5892# 0.023233f
C883 source.n844 a_n1094_n5892# 0.010408f
C884 source.n845 a_n1094_n5892# 0.018292f
C885 source.n846 a_n1094_n5892# 0.009829f
C886 source.n847 a_n1094_n5892# 0.023233f
C887 source.n848 a_n1094_n5892# 0.010408f
C888 source.n849 a_n1094_n5892# 0.018292f
C889 source.n850 a_n1094_n5892# 0.009829f
C890 source.n851 a_n1094_n5892# 0.023233f
C891 source.n852 a_n1094_n5892# 0.010408f
C892 source.n853 a_n1094_n5892# 0.018292f
C893 source.n854 a_n1094_n5892# 0.009829f
C894 source.n855 a_n1094_n5892# 0.023233f
C895 source.n856 a_n1094_n5892# 0.010408f
C896 source.n857 a_n1094_n5892# 0.018292f
C897 source.n858 a_n1094_n5892# 0.009829f
C898 source.n859 a_n1094_n5892# 0.023233f
C899 source.n860 a_n1094_n5892# 0.010408f
C900 source.n861 a_n1094_n5892# 0.018292f
C901 source.n862 a_n1094_n5892# 0.009829f
C902 source.n863 a_n1094_n5892# 0.023233f
C903 source.n864 a_n1094_n5892# 0.010408f
C904 source.n865 a_n1094_n5892# 0.018292f
C905 source.n866 a_n1094_n5892# 0.009829f
C906 source.n867 a_n1094_n5892# 0.023233f
C907 source.n868 a_n1094_n5892# 0.010408f
C908 source.n869 a_n1094_n5892# 0.018292f
C909 source.n870 a_n1094_n5892# 0.009829f
C910 source.n871 a_n1094_n5892# 0.023233f
C911 source.n872 a_n1094_n5892# 0.010408f
C912 source.n873 a_n1094_n5892# 0.018292f
C913 source.n874 a_n1094_n5892# 0.010119f
C914 source.n875 a_n1094_n5892# 0.023233f
C915 source.n876 a_n1094_n5892# 0.010408f
C916 source.n877 a_n1094_n5892# 0.018292f
C917 source.n878 a_n1094_n5892# 0.009829f
C918 source.n879 a_n1094_n5892# 0.023233f
C919 source.n880 a_n1094_n5892# 0.010408f
C920 source.n881 a_n1094_n5892# 0.018292f
C921 source.n882 a_n1094_n5892# 0.009829f
C922 source.n883 a_n1094_n5892# 0.017425f
C923 source.n884 a_n1094_n5892# 0.016424f
C924 source.t7 a_n1094_n5892# 0.04052f
C925 source.n885 a_n1094_n5892# 0.223181f
C926 source.n886 a_n1094_n5892# 1.98052f
C927 source.n887 a_n1094_n5892# 0.009829f
C928 source.n888 a_n1094_n5892# 0.010408f
C929 source.n889 a_n1094_n5892# 0.023233f
C930 source.n890 a_n1094_n5892# 0.023233f
C931 source.n891 a_n1094_n5892# 0.010408f
C932 source.n892 a_n1094_n5892# 0.009829f
C933 source.n893 a_n1094_n5892# 0.018292f
C934 source.n894 a_n1094_n5892# 0.018292f
C935 source.n895 a_n1094_n5892# 0.009829f
C936 source.n896 a_n1094_n5892# 0.010408f
C937 source.n897 a_n1094_n5892# 0.023233f
C938 source.n898 a_n1094_n5892# 0.023233f
C939 source.n899 a_n1094_n5892# 0.010408f
C940 source.n900 a_n1094_n5892# 0.009829f
C941 source.n901 a_n1094_n5892# 0.018292f
C942 source.n902 a_n1094_n5892# 0.018292f
C943 source.n903 a_n1094_n5892# 0.009829f
C944 source.n904 a_n1094_n5892# 0.009829f
C945 source.n905 a_n1094_n5892# 0.010408f
C946 source.n906 a_n1094_n5892# 0.023233f
C947 source.n907 a_n1094_n5892# 0.023233f
C948 source.n908 a_n1094_n5892# 0.023233f
C949 source.n909 a_n1094_n5892# 0.010119f
C950 source.n910 a_n1094_n5892# 0.009829f
C951 source.n911 a_n1094_n5892# 0.018292f
C952 source.n912 a_n1094_n5892# 0.018292f
C953 source.n913 a_n1094_n5892# 0.009829f
C954 source.n914 a_n1094_n5892# 0.010408f
C955 source.n915 a_n1094_n5892# 0.023233f
C956 source.n916 a_n1094_n5892# 0.023233f
C957 source.n917 a_n1094_n5892# 0.010408f
C958 source.n918 a_n1094_n5892# 0.009829f
C959 source.n919 a_n1094_n5892# 0.018292f
C960 source.n920 a_n1094_n5892# 0.018292f
C961 source.n921 a_n1094_n5892# 0.009829f
C962 source.n922 a_n1094_n5892# 0.010408f
C963 source.n923 a_n1094_n5892# 0.023233f
C964 source.n924 a_n1094_n5892# 0.023233f
C965 source.n925 a_n1094_n5892# 0.010408f
C966 source.n926 a_n1094_n5892# 0.009829f
C967 source.n927 a_n1094_n5892# 0.018292f
C968 source.n928 a_n1094_n5892# 0.018292f
C969 source.n929 a_n1094_n5892# 0.009829f
C970 source.n930 a_n1094_n5892# 0.010408f
C971 source.n931 a_n1094_n5892# 0.023233f
C972 source.n932 a_n1094_n5892# 0.023233f
C973 source.n933 a_n1094_n5892# 0.010408f
C974 source.n934 a_n1094_n5892# 0.009829f
C975 source.n935 a_n1094_n5892# 0.018292f
C976 source.n936 a_n1094_n5892# 0.018292f
C977 source.n937 a_n1094_n5892# 0.009829f
C978 source.n938 a_n1094_n5892# 0.010408f
C979 source.n939 a_n1094_n5892# 0.023233f
C980 source.n940 a_n1094_n5892# 0.023233f
C981 source.n941 a_n1094_n5892# 0.010408f
C982 source.n942 a_n1094_n5892# 0.009829f
C983 source.n943 a_n1094_n5892# 0.018292f
C984 source.n944 a_n1094_n5892# 0.018292f
C985 source.n945 a_n1094_n5892# 0.009829f
C986 source.n946 a_n1094_n5892# 0.010408f
C987 source.n947 a_n1094_n5892# 0.023233f
C988 source.n948 a_n1094_n5892# 0.023233f
C989 source.n949 a_n1094_n5892# 0.023233f
C990 source.n950 a_n1094_n5892# 0.010408f
C991 source.n951 a_n1094_n5892# 0.009829f
C992 source.n952 a_n1094_n5892# 0.018292f
C993 source.n953 a_n1094_n5892# 0.018292f
C994 source.n954 a_n1094_n5892# 0.009829f
C995 source.n955 a_n1094_n5892# 0.010119f
C996 source.n956 a_n1094_n5892# 0.010119f
C997 source.n957 a_n1094_n5892# 0.023233f
C998 source.n958 a_n1094_n5892# 0.023233f
C999 source.n959 a_n1094_n5892# 0.010408f
C1000 source.n960 a_n1094_n5892# 0.009829f
C1001 source.n961 a_n1094_n5892# 0.018292f
C1002 source.n962 a_n1094_n5892# 0.018292f
C1003 source.n963 a_n1094_n5892# 0.009829f
C1004 source.n964 a_n1094_n5892# 0.010408f
C1005 source.n965 a_n1094_n5892# 0.023233f
C1006 source.n966 a_n1094_n5892# 0.023233f
C1007 source.n967 a_n1094_n5892# 0.010408f
C1008 source.n968 a_n1094_n5892# 0.009829f
C1009 source.n969 a_n1094_n5892# 0.018292f
C1010 source.n970 a_n1094_n5892# 0.018292f
C1011 source.n971 a_n1094_n5892# 0.009829f
C1012 source.n972 a_n1094_n5892# 0.010408f
C1013 source.n973 a_n1094_n5892# 0.023233f
C1014 source.n974 a_n1094_n5892# 0.049423f
C1015 source.n975 a_n1094_n5892# 0.010408f
C1016 source.n976 a_n1094_n5892# 0.009829f
C1017 source.n977 a_n1094_n5892# 0.040283f
C1018 source.n978 a_n1094_n5892# 0.027502f
C1019 source.n979 a_n1094_n5892# 0.0742f
C1020 source.n980 a_n1094_n5892# 0.025218f
C1021 source.n981 a_n1094_n5892# 0.018292f
C1022 source.n982 a_n1094_n5892# 0.009829f
C1023 source.n983 a_n1094_n5892# 0.023233f
C1024 source.n984 a_n1094_n5892# 0.010408f
C1025 source.n985 a_n1094_n5892# 0.018292f
C1026 source.n986 a_n1094_n5892# 0.009829f
C1027 source.n987 a_n1094_n5892# 0.023233f
C1028 source.n988 a_n1094_n5892# 0.010408f
C1029 source.n989 a_n1094_n5892# 0.018292f
C1030 source.n990 a_n1094_n5892# 0.009829f
C1031 source.n991 a_n1094_n5892# 0.023233f
C1032 source.n992 a_n1094_n5892# 0.010408f
C1033 source.n993 a_n1094_n5892# 0.018292f
C1034 source.n994 a_n1094_n5892# 0.009829f
C1035 source.n995 a_n1094_n5892# 0.023233f
C1036 source.n996 a_n1094_n5892# 0.010408f
C1037 source.n997 a_n1094_n5892# 0.018292f
C1038 source.n998 a_n1094_n5892# 0.009829f
C1039 source.n999 a_n1094_n5892# 0.023233f
C1040 source.n1000 a_n1094_n5892# 0.010408f
C1041 source.n1001 a_n1094_n5892# 0.018292f
C1042 source.n1002 a_n1094_n5892# 0.009829f
C1043 source.n1003 a_n1094_n5892# 0.023233f
C1044 source.n1004 a_n1094_n5892# 0.010408f
C1045 source.n1005 a_n1094_n5892# 0.018292f
C1046 source.n1006 a_n1094_n5892# 0.009829f
C1047 source.n1007 a_n1094_n5892# 0.023233f
C1048 source.n1008 a_n1094_n5892# 0.010408f
C1049 source.n1009 a_n1094_n5892# 0.018292f
C1050 source.n1010 a_n1094_n5892# 0.009829f
C1051 source.n1011 a_n1094_n5892# 0.023233f
C1052 source.n1012 a_n1094_n5892# 0.010408f
C1053 source.n1013 a_n1094_n5892# 0.018292f
C1054 source.n1014 a_n1094_n5892# 0.010119f
C1055 source.n1015 a_n1094_n5892# 0.023233f
C1056 source.n1016 a_n1094_n5892# 0.010408f
C1057 source.n1017 a_n1094_n5892# 0.018292f
C1058 source.n1018 a_n1094_n5892# 0.009829f
C1059 source.n1019 a_n1094_n5892# 0.023233f
C1060 source.n1020 a_n1094_n5892# 0.010408f
C1061 source.n1021 a_n1094_n5892# 0.018292f
C1062 source.n1022 a_n1094_n5892# 0.009829f
C1063 source.n1023 a_n1094_n5892# 0.017425f
C1064 source.n1024 a_n1094_n5892# 0.016424f
C1065 source.t4 a_n1094_n5892# 0.04052f
C1066 source.n1025 a_n1094_n5892# 0.223181f
C1067 source.n1026 a_n1094_n5892# 1.98052f
C1068 source.n1027 a_n1094_n5892# 0.009829f
C1069 source.n1028 a_n1094_n5892# 0.010408f
C1070 source.n1029 a_n1094_n5892# 0.023233f
C1071 source.n1030 a_n1094_n5892# 0.023233f
C1072 source.n1031 a_n1094_n5892# 0.010408f
C1073 source.n1032 a_n1094_n5892# 0.009829f
C1074 source.n1033 a_n1094_n5892# 0.018292f
C1075 source.n1034 a_n1094_n5892# 0.018292f
C1076 source.n1035 a_n1094_n5892# 0.009829f
C1077 source.n1036 a_n1094_n5892# 0.010408f
C1078 source.n1037 a_n1094_n5892# 0.023233f
C1079 source.n1038 a_n1094_n5892# 0.023233f
C1080 source.n1039 a_n1094_n5892# 0.010408f
C1081 source.n1040 a_n1094_n5892# 0.009829f
C1082 source.n1041 a_n1094_n5892# 0.018292f
C1083 source.n1042 a_n1094_n5892# 0.018292f
C1084 source.n1043 a_n1094_n5892# 0.009829f
C1085 source.n1044 a_n1094_n5892# 0.009829f
C1086 source.n1045 a_n1094_n5892# 0.010408f
C1087 source.n1046 a_n1094_n5892# 0.023233f
C1088 source.n1047 a_n1094_n5892# 0.023233f
C1089 source.n1048 a_n1094_n5892# 0.023233f
C1090 source.n1049 a_n1094_n5892# 0.010119f
C1091 source.n1050 a_n1094_n5892# 0.009829f
C1092 source.n1051 a_n1094_n5892# 0.018292f
C1093 source.n1052 a_n1094_n5892# 0.018292f
C1094 source.n1053 a_n1094_n5892# 0.009829f
C1095 source.n1054 a_n1094_n5892# 0.010408f
C1096 source.n1055 a_n1094_n5892# 0.023233f
C1097 source.n1056 a_n1094_n5892# 0.023233f
C1098 source.n1057 a_n1094_n5892# 0.010408f
C1099 source.n1058 a_n1094_n5892# 0.009829f
C1100 source.n1059 a_n1094_n5892# 0.018292f
C1101 source.n1060 a_n1094_n5892# 0.018292f
C1102 source.n1061 a_n1094_n5892# 0.009829f
C1103 source.n1062 a_n1094_n5892# 0.010408f
C1104 source.n1063 a_n1094_n5892# 0.023233f
C1105 source.n1064 a_n1094_n5892# 0.023233f
C1106 source.n1065 a_n1094_n5892# 0.010408f
C1107 source.n1066 a_n1094_n5892# 0.009829f
C1108 source.n1067 a_n1094_n5892# 0.018292f
C1109 source.n1068 a_n1094_n5892# 0.018292f
C1110 source.n1069 a_n1094_n5892# 0.009829f
C1111 source.n1070 a_n1094_n5892# 0.010408f
C1112 source.n1071 a_n1094_n5892# 0.023233f
C1113 source.n1072 a_n1094_n5892# 0.023233f
C1114 source.n1073 a_n1094_n5892# 0.010408f
C1115 source.n1074 a_n1094_n5892# 0.009829f
C1116 source.n1075 a_n1094_n5892# 0.018292f
C1117 source.n1076 a_n1094_n5892# 0.018292f
C1118 source.n1077 a_n1094_n5892# 0.009829f
C1119 source.n1078 a_n1094_n5892# 0.010408f
C1120 source.n1079 a_n1094_n5892# 0.023233f
C1121 source.n1080 a_n1094_n5892# 0.023233f
C1122 source.n1081 a_n1094_n5892# 0.010408f
C1123 source.n1082 a_n1094_n5892# 0.009829f
C1124 source.n1083 a_n1094_n5892# 0.018292f
C1125 source.n1084 a_n1094_n5892# 0.018292f
C1126 source.n1085 a_n1094_n5892# 0.009829f
C1127 source.n1086 a_n1094_n5892# 0.010408f
C1128 source.n1087 a_n1094_n5892# 0.023233f
C1129 source.n1088 a_n1094_n5892# 0.023233f
C1130 source.n1089 a_n1094_n5892# 0.023233f
C1131 source.n1090 a_n1094_n5892# 0.010408f
C1132 source.n1091 a_n1094_n5892# 0.009829f
C1133 source.n1092 a_n1094_n5892# 0.018292f
C1134 source.n1093 a_n1094_n5892# 0.018292f
C1135 source.n1094 a_n1094_n5892# 0.009829f
C1136 source.n1095 a_n1094_n5892# 0.010119f
C1137 source.n1096 a_n1094_n5892# 0.010119f
C1138 source.n1097 a_n1094_n5892# 0.023233f
C1139 source.n1098 a_n1094_n5892# 0.023233f
C1140 source.n1099 a_n1094_n5892# 0.010408f
C1141 source.n1100 a_n1094_n5892# 0.009829f
C1142 source.n1101 a_n1094_n5892# 0.018292f
C1143 source.n1102 a_n1094_n5892# 0.018292f
C1144 source.n1103 a_n1094_n5892# 0.009829f
C1145 source.n1104 a_n1094_n5892# 0.010408f
C1146 source.n1105 a_n1094_n5892# 0.023233f
C1147 source.n1106 a_n1094_n5892# 0.023233f
C1148 source.n1107 a_n1094_n5892# 0.010408f
C1149 source.n1108 a_n1094_n5892# 0.009829f
C1150 source.n1109 a_n1094_n5892# 0.018292f
C1151 source.n1110 a_n1094_n5892# 0.018292f
C1152 source.n1111 a_n1094_n5892# 0.009829f
C1153 source.n1112 a_n1094_n5892# 0.010408f
C1154 source.n1113 a_n1094_n5892# 0.023233f
C1155 source.n1114 a_n1094_n5892# 0.049423f
C1156 source.n1115 a_n1094_n5892# 0.010408f
C1157 source.n1116 a_n1094_n5892# 0.009829f
C1158 source.n1117 a_n1094_n5892# 0.040283f
C1159 source.n1118 a_n1094_n5892# 0.027502f
C1160 source.n1119 a_n1094_n5892# 0.17746f
C1161 source.n1120 a_n1094_n5892# 1.95119f
C1162 minus.t2 a_n1094_n5892# 1.31471f
C1163 minus.t0 a_n1094_n5892# 1.31471f
C1164 minus.n0 a_n1094_n5892# 1.56734f
C1165 minus.t3 a_n1094_n5892# 1.31471f
C1166 minus.t1 a_n1094_n5892# 1.31471f
C1167 minus.n1 a_n1094_n5892# 0.979522f
C1168 minus.n2 a_n1094_n5892# 6.05369f
.ends

