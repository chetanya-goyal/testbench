* NGSPICE file created from diffpair197.ext - technology: sky130A

.subckt diffpair197 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t17 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 drain_left.t15 plus.t0 source.t7 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X2 source.t18 minus.t1 drain_right.t14 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X3 drain_right.t13 minus.t2 source.t23 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X4 drain_left.t14 plus.t1 source.t10 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X5 drain_right.t12 minus.t3 source.t19 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X6 a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X7 source.t26 minus.t4 drain_right.t11 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X8 source.t0 plus.t2 drain_left.t13 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X9 source.t13 plus.t3 drain_left.t12 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X10 a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X11 drain_left.t11 plus.t4 source.t2 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X12 drain_right.t10 minus.t5 source.t29 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X13 a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X14 source.t22 minus.t6 drain_right.t9 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X15 source.t1 plus.t5 drain_left.t10 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X16 source.t15 plus.t6 drain_left.t9 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X17 drain_left.t8 plus.t7 source.t4 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X18 drain_right.t8 minus.t7 source.t27 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X19 source.t28 minus.t8 drain_right.t7 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X20 drain_left.t7 plus.t8 source.t14 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X21 drain_right.t6 minus.t9 source.t20 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X22 drain_right.t5 minus.t10 source.t30 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X23 drain_left.t6 plus.t9 source.t5 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X24 a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X25 source.t21 minus.t11 drain_right.t4 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X26 source.t8 plus.t10 drain_left.t5 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X27 drain_left.t4 plus.t11 source.t11 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X28 drain_right.t3 minus.t12 source.t25 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X29 source.t16 minus.t13 drain_right.t2 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X30 source.t24 minus.t14 drain_right.t1 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X31 source.t31 minus.t15 drain_right.t0 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X32 source.t3 plus.t12 drain_left.t3 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X33 source.t12 plus.t13 drain_left.t2 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X34 source.t6 plus.t14 drain_left.t1 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X35 drain_left.t0 plus.t15 source.t9 a_n1850_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n21 minus.t14 375.377
R1 minus.n5 minus.t9 375.377
R2 minus.n44 minus.t10 375.377
R3 minus.n28 minus.t6 375.377
R4 minus.n20 minus.t5 345.433
R5 minus.n1 minus.t1 345.433
R6 minus.n14 minus.t12 345.433
R7 minus.n12 minus.t8 345.433
R8 minus.n3 minus.t3 345.433
R9 minus.n6 minus.t13 345.433
R10 minus.n43 minus.t11 345.433
R11 minus.n24 minus.t2 345.433
R12 minus.n37 minus.t4 345.433
R13 minus.n35 minus.t7 345.433
R14 minus.n26 minus.t15 345.433
R15 minus.n29 minus.t0 345.433
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 64.9975
R39 minus.n11 minus.n3 64.9975
R40 minus.n34 minus.n26 64.9975
R41 minus.n38 minus.n24 64.9975
R42 minus.n21 minus.n20 62.0763
R43 minus.n6 minus.n5 62.0763
R44 minus.n29 minus.n28 62.0763
R45 minus.n44 minus.n43 62.0763
R46 minus.n14 minus.n13 46.0096
R47 minus.n13 minus.n12 46.0096
R48 minus.n36 minus.n35 46.0096
R49 minus.n37 minus.n36 46.0096
R50 minus.n46 minus.n22 29.277
R51 minus.n15 minus.n14 27.0217
R52 minus.n12 minus.n11 27.0217
R53 minus.n35 minus.n34 27.0217
R54 minus.n38 minus.n37 27.0217
R55 minus.n20 minus.n19 10.955
R56 minus.n7 minus.n6 10.955
R57 minus.n30 minus.n29 10.955
R58 minus.n43 minus.n42 10.955
R59 minus.n18 minus.n1 8.03383
R60 minus.n8 minus.n3 8.03383
R61 minus.n31 minus.n26 8.03383
R62 minus.n41 minus.n24 8.03383
R63 minus.n46 minus.n45 6.46641
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 source.n0 source.t7 69.6943
R80 source.n7 source.t13 69.6943
R81 source.n8 source.t20 69.6943
R82 source.n15 source.t24 69.6943
R83 source.n31 source.t30 69.6942
R84 source.n24 source.t22 69.6942
R85 source.n23 source.t2 69.6942
R86 source.n16 source.t0 69.6942
R87 source.n2 source.n1 63.0943
R88 source.n4 source.n3 63.0943
R89 source.n6 source.n5 63.0943
R90 source.n10 source.n9 63.0943
R91 source.n12 source.n11 63.0943
R92 source.n14 source.n13 63.0943
R93 source.n30 source.n29 63.0942
R94 source.n28 source.n27 63.0942
R95 source.n26 source.n25 63.0942
R96 source.n22 source.n21 63.0942
R97 source.n20 source.n19 63.0942
R98 source.n18 source.n17 63.0942
R99 source.n16 source.n15 15.0126
R100 source.n32 source.n0 9.47816
R101 source.n29 source.t23 6.6005
R102 source.n29 source.t21 6.6005
R103 source.n27 source.t27 6.6005
R104 source.n27 source.t26 6.6005
R105 source.n25 source.t17 6.6005
R106 source.n25 source.t31 6.6005
R107 source.n21 source.t11 6.6005
R108 source.n21 source.t3 6.6005
R109 source.n19 source.t10 6.6005
R110 source.n19 source.t15 6.6005
R111 source.n17 source.t14 6.6005
R112 source.n17 source.t6 6.6005
R113 source.n1 source.t5 6.6005
R114 source.n1 source.t12 6.6005
R115 source.n3 source.t9 6.6005
R116 source.n3 source.t1 6.6005
R117 source.n5 source.t4 6.6005
R118 source.n5 source.t8 6.6005
R119 source.n9 source.t19 6.6005
R120 source.n9 source.t16 6.6005
R121 source.n11 source.t25 6.6005
R122 source.n11 source.t28 6.6005
R123 source.n13 source.t29 6.6005
R124 source.n13 source.t18 6.6005
R125 source.n32 source.n31 5.53498
R126 source.n15 source.n14 0.543603
R127 source.n14 source.n12 0.543603
R128 source.n12 source.n10 0.543603
R129 source.n10 source.n8 0.543603
R130 source.n7 source.n6 0.543603
R131 source.n6 source.n4 0.543603
R132 source.n4 source.n2 0.543603
R133 source.n2 source.n0 0.543603
R134 source.n18 source.n16 0.543603
R135 source.n20 source.n18 0.543603
R136 source.n22 source.n20 0.543603
R137 source.n23 source.n22 0.543603
R138 source.n26 source.n24 0.543603
R139 source.n28 source.n26 0.543603
R140 source.n30 source.n28 0.543603
R141 source.n31 source.n30 0.543603
R142 source.n8 source.n7 0.470328
R143 source.n24 source.n23 0.470328
R144 source source.n32 0.188
R145 drain_right.n9 drain_right.n7 80.3162
R146 drain_right.n5 drain_right.n3 80.3161
R147 drain_right.n2 drain_right.n0 80.3161
R148 drain_right.n9 drain_right.n8 79.7731
R149 drain_right.n11 drain_right.n10 79.7731
R150 drain_right.n13 drain_right.n12 79.7731
R151 drain_right.n5 drain_right.n4 79.773
R152 drain_right.n2 drain_right.n1 79.773
R153 drain_right drain_right.n6 23.5258
R154 drain_right.n3 drain_right.t4 6.6005
R155 drain_right.n3 drain_right.t5 6.6005
R156 drain_right.n4 drain_right.t11 6.6005
R157 drain_right.n4 drain_right.t13 6.6005
R158 drain_right.n1 drain_right.t0 6.6005
R159 drain_right.n1 drain_right.t8 6.6005
R160 drain_right.n0 drain_right.t9 6.6005
R161 drain_right.n0 drain_right.t15 6.6005
R162 drain_right.n7 drain_right.t2 6.6005
R163 drain_right.n7 drain_right.t6 6.6005
R164 drain_right.n8 drain_right.t7 6.6005
R165 drain_right.n8 drain_right.t12 6.6005
R166 drain_right.n10 drain_right.t14 6.6005
R167 drain_right.n10 drain_right.t3 6.6005
R168 drain_right.n12 drain_right.t1 6.6005
R169 drain_right.n12 drain_right.t10 6.6005
R170 drain_right drain_right.n13 6.19632
R171 drain_right.n13 drain_right.n11 0.543603
R172 drain_right.n11 drain_right.n9 0.543603
R173 drain_right.n6 drain_right.n5 0.216706
R174 drain_right.n6 drain_right.n2 0.216706
R175 plus.n5 plus.t3 375.377
R176 plus.n21 plus.t0 375.377
R177 plus.n28 plus.t4 375.377
R178 plus.n44 plus.t2 375.377
R179 plus.n6 plus.t7 345.433
R180 plus.n3 plus.t10 345.433
R181 plus.n12 plus.t15 345.433
R182 plus.n14 plus.t5 345.433
R183 plus.n1 plus.t9 345.433
R184 plus.n20 plus.t13 345.433
R185 plus.n29 plus.t12 345.433
R186 plus.n26 plus.t11 345.433
R187 plus.n35 plus.t6 345.433
R188 plus.n37 plus.t1 345.433
R189 plus.n24 plus.t14 345.433
R190 plus.n43 plus.t8 345.433
R191 plus.n5 plus.n4 161.489
R192 plus.n28 plus.n27 161.489
R193 plus.n7 plus.n4 161.3
R194 plus.n9 plus.n8 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n13 plus.n2 161.3
R197 plus.n16 plus.n15 161.3
R198 plus.n18 plus.n17 161.3
R199 plus.n19 plus.n0 161.3
R200 plus.n22 plus.n21 161.3
R201 plus.n30 plus.n27 161.3
R202 plus.n32 plus.n31 161.3
R203 plus.n34 plus.n33 161.3
R204 plus.n36 plus.n25 161.3
R205 plus.n39 plus.n38 161.3
R206 plus.n41 plus.n40 161.3
R207 plus.n42 plus.n23 161.3
R208 plus.n45 plus.n44 161.3
R209 plus.n8 plus.n7 73.0308
R210 plus.n19 plus.n18 73.0308
R211 plus.n42 plus.n41 73.0308
R212 plus.n31 plus.n30 73.0308
R213 plus.n11 plus.n3 64.9975
R214 plus.n15 plus.n1 64.9975
R215 plus.n38 plus.n24 64.9975
R216 plus.n34 plus.n26 64.9975
R217 plus.n6 plus.n5 62.0763
R218 plus.n21 plus.n20 62.0763
R219 plus.n44 plus.n43 62.0763
R220 plus.n29 plus.n28 62.0763
R221 plus.n13 plus.n12 46.0096
R222 plus.n14 plus.n13 46.0096
R223 plus.n37 plus.n36 46.0096
R224 plus.n36 plus.n35 46.0096
R225 plus.n12 plus.n11 27.0217
R226 plus.n15 plus.n14 27.0217
R227 plus.n38 plus.n37 27.0217
R228 plus.n35 plus.n34 27.0217
R229 plus plus.n45 26.5672
R230 plus.n7 plus.n6 10.955
R231 plus.n20 plus.n19 10.955
R232 plus.n43 plus.n42 10.955
R233 plus.n30 plus.n29 10.955
R234 plus plus.n22 8.70126
R235 plus.n8 plus.n3 8.03383
R236 plus.n18 plus.n1 8.03383
R237 plus.n41 plus.n24 8.03383
R238 plus.n31 plus.n26 8.03383
R239 plus.n9 plus.n4 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n2 0.189894
R242 plus.n16 plus.n2 0.189894
R243 plus.n17 plus.n16 0.189894
R244 plus.n17 plus.n0 0.189894
R245 plus.n22 plus.n0 0.189894
R246 plus.n45 plus.n23 0.189894
R247 plus.n40 plus.n23 0.189894
R248 plus.n40 plus.n39 0.189894
R249 plus.n39 plus.n25 0.189894
R250 plus.n33 plus.n25 0.189894
R251 plus.n33 plus.n32 0.189894
R252 plus.n32 plus.n27 0.189894
R253 drain_left.n9 drain_left.n7 80.3162
R254 drain_left.n5 drain_left.n3 80.3161
R255 drain_left.n2 drain_left.n0 80.3161
R256 drain_left.n13 drain_left.n12 79.7731
R257 drain_left.n11 drain_left.n10 79.7731
R258 drain_left.n9 drain_left.n8 79.7731
R259 drain_left.n5 drain_left.n4 79.773
R260 drain_left.n2 drain_left.n1 79.773
R261 drain_left drain_left.n6 24.0791
R262 drain_left.n3 drain_left.t3 6.6005
R263 drain_left.n3 drain_left.t11 6.6005
R264 drain_left.n4 drain_left.t9 6.6005
R265 drain_left.n4 drain_left.t4 6.6005
R266 drain_left.n1 drain_left.t1 6.6005
R267 drain_left.n1 drain_left.t14 6.6005
R268 drain_left.n0 drain_left.t13 6.6005
R269 drain_left.n0 drain_left.t7 6.6005
R270 drain_left.n12 drain_left.t2 6.6005
R271 drain_left.n12 drain_left.t15 6.6005
R272 drain_left.n10 drain_left.t10 6.6005
R273 drain_left.n10 drain_left.t6 6.6005
R274 drain_left.n8 drain_left.t5 6.6005
R275 drain_left.n8 drain_left.t0 6.6005
R276 drain_left.n7 drain_left.t12 6.6005
R277 drain_left.n7 drain_left.t8 6.6005
R278 drain_left drain_left.n13 6.19632
R279 drain_left.n11 drain_left.n9 0.543603
R280 drain_left.n13 drain_left.n11 0.543603
R281 drain_left.n6 drain_left.n5 0.216706
R282 drain_left.n6 drain_left.n2 0.216706
C0 drain_right drain_left 0.948737f
C1 plus minus 3.80312f
C2 plus drain_left 2.04026f
C3 drain_left minus 0.17667f
C4 drain_right source 9.73896f
C5 plus source 2.02871f
C6 minus source 2.01471f
C7 drain_right plus 0.33988f
C8 drain_left source 9.73872f
C9 drain_right minus 1.86057f
C10 drain_right a_n1850_n1488# 4.16619f
C11 drain_left a_n1850_n1488# 4.75215f
C12 source a_n1850_n1488# 3.686164f
C13 minus a_n1850_n1488# 6.513808f
C14 plus a_n1850_n1488# 7.882361f
C15 drain_left.t13 a_n1850_n1488# 0.075965f
C16 drain_left.t7 a_n1850_n1488# 0.075965f
C17 drain_left.n0 a_n1850_n1488# 0.550431f
C18 drain_left.t1 a_n1850_n1488# 0.075965f
C19 drain_left.t14 a_n1850_n1488# 0.075965f
C20 drain_left.n1 a_n1850_n1488# 0.547851f
C21 drain_left.n2 a_n1850_n1488# 0.717317f
C22 drain_left.t3 a_n1850_n1488# 0.075965f
C23 drain_left.t11 a_n1850_n1488# 0.075965f
C24 drain_left.n3 a_n1850_n1488# 0.550431f
C25 drain_left.t9 a_n1850_n1488# 0.075965f
C26 drain_left.t4 a_n1850_n1488# 0.075965f
C27 drain_left.n4 a_n1850_n1488# 0.547851f
C28 drain_left.n5 a_n1850_n1488# 0.717317f
C29 drain_left.n6 a_n1850_n1488# 0.970891f
C30 drain_left.t12 a_n1850_n1488# 0.075965f
C31 drain_left.t8 a_n1850_n1488# 0.075965f
C32 drain_left.n7 a_n1850_n1488# 0.550433f
C33 drain_left.t5 a_n1850_n1488# 0.075965f
C34 drain_left.t0 a_n1850_n1488# 0.075965f
C35 drain_left.n8 a_n1850_n1488# 0.547853f
C36 drain_left.n9 a_n1850_n1488# 0.747628f
C37 drain_left.t10 a_n1850_n1488# 0.075965f
C38 drain_left.t6 a_n1850_n1488# 0.075965f
C39 drain_left.n10 a_n1850_n1488# 0.547853f
C40 drain_left.n11 a_n1850_n1488# 0.368651f
C41 drain_left.t2 a_n1850_n1488# 0.075965f
C42 drain_left.t15 a_n1850_n1488# 0.075965f
C43 drain_left.n12 a_n1850_n1488# 0.547853f
C44 drain_left.n13 a_n1850_n1488# 0.635367f
C45 plus.n0 a_n1850_n1488# 0.051967f
C46 plus.t13 a_n1850_n1488# 0.135441f
C47 plus.t9 a_n1850_n1488# 0.135441f
C48 plus.n1 a_n1850_n1488# 0.078643f
C49 plus.n2 a_n1850_n1488# 0.051967f
C50 plus.t5 a_n1850_n1488# 0.135441f
C51 plus.t15 a_n1850_n1488# 0.135441f
C52 plus.t10 a_n1850_n1488# 0.135441f
C53 plus.n3 a_n1850_n1488# 0.078643f
C54 plus.n4 a_n1850_n1488# 0.110593f
C55 plus.t7 a_n1850_n1488# 0.135441f
C56 plus.t3 a_n1850_n1488# 0.141727f
C57 plus.n5 a_n1850_n1488# 0.093991f
C58 plus.n6 a_n1850_n1488# 0.078643f
C59 plus.n7 a_n1850_n1488# 0.019642f
C60 plus.n8 a_n1850_n1488# 0.019001f
C61 plus.n9 a_n1850_n1488# 0.051967f
C62 plus.n10 a_n1850_n1488# 0.051967f
C63 plus.n11 a_n1850_n1488# 0.021404f
C64 plus.n12 a_n1850_n1488# 0.078643f
C65 plus.n13 a_n1850_n1488# 0.021404f
C66 plus.n14 a_n1850_n1488# 0.078643f
C67 plus.n15 a_n1850_n1488# 0.021404f
C68 plus.n16 a_n1850_n1488# 0.051967f
C69 plus.n17 a_n1850_n1488# 0.051967f
C70 plus.n18 a_n1850_n1488# 0.019001f
C71 plus.n19 a_n1850_n1488# 0.019642f
C72 plus.n20 a_n1850_n1488# 0.078643f
C73 plus.t0 a_n1850_n1488# 0.141727f
C74 plus.n21 a_n1850_n1488# 0.093922f
C75 plus.n22 a_n1850_n1488# 0.383854f
C76 plus.n23 a_n1850_n1488# 0.051967f
C77 plus.t2 a_n1850_n1488# 0.141727f
C78 plus.t8 a_n1850_n1488# 0.135441f
C79 plus.t14 a_n1850_n1488# 0.135441f
C80 plus.n24 a_n1850_n1488# 0.078643f
C81 plus.n25 a_n1850_n1488# 0.051967f
C82 plus.t1 a_n1850_n1488# 0.135441f
C83 plus.t6 a_n1850_n1488# 0.135441f
C84 plus.t11 a_n1850_n1488# 0.135441f
C85 plus.n26 a_n1850_n1488# 0.078643f
C86 plus.n27 a_n1850_n1488# 0.110593f
C87 plus.t12 a_n1850_n1488# 0.135441f
C88 plus.t4 a_n1850_n1488# 0.141727f
C89 plus.n28 a_n1850_n1488# 0.093991f
C90 plus.n29 a_n1850_n1488# 0.078643f
C91 plus.n30 a_n1850_n1488# 0.019642f
C92 plus.n31 a_n1850_n1488# 0.019001f
C93 plus.n32 a_n1850_n1488# 0.051967f
C94 plus.n33 a_n1850_n1488# 0.051967f
C95 plus.n34 a_n1850_n1488# 0.021404f
C96 plus.n35 a_n1850_n1488# 0.078643f
C97 plus.n36 a_n1850_n1488# 0.021404f
C98 plus.n37 a_n1850_n1488# 0.078643f
C99 plus.n38 a_n1850_n1488# 0.021404f
C100 plus.n39 a_n1850_n1488# 0.051967f
C101 plus.n40 a_n1850_n1488# 0.051967f
C102 plus.n41 a_n1850_n1488# 0.019001f
C103 plus.n42 a_n1850_n1488# 0.019642f
C104 plus.n43 a_n1850_n1488# 0.078643f
C105 plus.n44 a_n1850_n1488# 0.093922f
C106 plus.n45 a_n1850_n1488# 1.21762f
C107 drain_right.t9 a_n1850_n1488# 0.063662f
C108 drain_right.t15 a_n1850_n1488# 0.063662f
C109 drain_right.n0 a_n1850_n1488# 0.461282f
C110 drain_right.t0 a_n1850_n1488# 0.063662f
C111 drain_right.t8 a_n1850_n1488# 0.063662f
C112 drain_right.n1 a_n1850_n1488# 0.45912f
C113 drain_right.n2 a_n1850_n1488# 0.601139f
C114 drain_right.t4 a_n1850_n1488# 0.063662f
C115 drain_right.t5 a_n1850_n1488# 0.063662f
C116 drain_right.n3 a_n1850_n1488# 0.461282f
C117 drain_right.t11 a_n1850_n1488# 0.063662f
C118 drain_right.t13 a_n1850_n1488# 0.063662f
C119 drain_right.n4 a_n1850_n1488# 0.45912f
C120 drain_right.n5 a_n1850_n1488# 0.601139f
C121 drain_right.n6 a_n1850_n1488# 0.760444f
C122 drain_right.t2 a_n1850_n1488# 0.063662f
C123 drain_right.t6 a_n1850_n1488# 0.063662f
C124 drain_right.n7 a_n1850_n1488# 0.461284f
C125 drain_right.t7 a_n1850_n1488# 0.063662f
C126 drain_right.t12 a_n1850_n1488# 0.063662f
C127 drain_right.n8 a_n1850_n1488# 0.459122f
C128 drain_right.n9 a_n1850_n1488# 0.626541f
C129 drain_right.t14 a_n1850_n1488# 0.063662f
C130 drain_right.t3 a_n1850_n1488# 0.063662f
C131 drain_right.n10 a_n1850_n1488# 0.459122f
C132 drain_right.n11 a_n1850_n1488# 0.308944f
C133 drain_right.t1 a_n1850_n1488# 0.063662f
C134 drain_right.t10 a_n1850_n1488# 0.063662f
C135 drain_right.n12 a_n1850_n1488# 0.459122f
C136 drain_right.n13 a_n1850_n1488# 0.532462f
C137 source.t7 a_n1850_n1488# 0.615869f
C138 source.n0 a_n1850_n1488# 0.840251f
C139 source.t5 a_n1850_n1488# 0.074167f
C140 source.t12 a_n1850_n1488# 0.074167f
C141 source.n1 a_n1850_n1488# 0.470261f
C142 source.n2 a_n1850_n1488# 0.382029f
C143 source.t9 a_n1850_n1488# 0.074167f
C144 source.t1 a_n1850_n1488# 0.074167f
C145 source.n3 a_n1850_n1488# 0.470261f
C146 source.n4 a_n1850_n1488# 0.382029f
C147 source.t4 a_n1850_n1488# 0.074167f
C148 source.t8 a_n1850_n1488# 0.074167f
C149 source.n5 a_n1850_n1488# 0.470261f
C150 source.n6 a_n1850_n1488# 0.382029f
C151 source.t13 a_n1850_n1488# 0.615869f
C152 source.n7 a_n1850_n1488# 0.431308f
C153 source.t20 a_n1850_n1488# 0.615869f
C154 source.n8 a_n1850_n1488# 0.431308f
C155 source.t19 a_n1850_n1488# 0.074167f
C156 source.t16 a_n1850_n1488# 0.074167f
C157 source.n9 a_n1850_n1488# 0.470261f
C158 source.n10 a_n1850_n1488# 0.382029f
C159 source.t25 a_n1850_n1488# 0.074167f
C160 source.t28 a_n1850_n1488# 0.074167f
C161 source.n11 a_n1850_n1488# 0.470261f
C162 source.n12 a_n1850_n1488# 0.382029f
C163 source.t29 a_n1850_n1488# 0.074167f
C164 source.t18 a_n1850_n1488# 0.074167f
C165 source.n13 a_n1850_n1488# 0.470261f
C166 source.n14 a_n1850_n1488# 0.382029f
C167 source.t24 a_n1850_n1488# 0.615869f
C168 source.n15 a_n1850_n1488# 1.16635f
C169 source.t0 a_n1850_n1488# 0.615866f
C170 source.n16 a_n1850_n1488# 1.16636f
C171 source.t14 a_n1850_n1488# 0.074167f
C172 source.t6 a_n1850_n1488# 0.074167f
C173 source.n17 a_n1850_n1488# 0.470257f
C174 source.n18 a_n1850_n1488# 0.382033f
C175 source.t10 a_n1850_n1488# 0.074167f
C176 source.t15 a_n1850_n1488# 0.074167f
C177 source.n19 a_n1850_n1488# 0.470257f
C178 source.n20 a_n1850_n1488# 0.382033f
C179 source.t11 a_n1850_n1488# 0.074167f
C180 source.t3 a_n1850_n1488# 0.074167f
C181 source.n21 a_n1850_n1488# 0.470257f
C182 source.n22 a_n1850_n1488# 0.382033f
C183 source.t2 a_n1850_n1488# 0.615866f
C184 source.n23 a_n1850_n1488# 0.431311f
C185 source.t22 a_n1850_n1488# 0.615866f
C186 source.n24 a_n1850_n1488# 0.431311f
C187 source.t17 a_n1850_n1488# 0.074167f
C188 source.t31 a_n1850_n1488# 0.074167f
C189 source.n25 a_n1850_n1488# 0.470257f
C190 source.n26 a_n1850_n1488# 0.382033f
C191 source.t27 a_n1850_n1488# 0.074167f
C192 source.t26 a_n1850_n1488# 0.074167f
C193 source.n27 a_n1850_n1488# 0.470257f
C194 source.n28 a_n1850_n1488# 0.382033f
C195 source.t23 a_n1850_n1488# 0.074167f
C196 source.t21 a_n1850_n1488# 0.074167f
C197 source.n29 a_n1850_n1488# 0.470257f
C198 source.n30 a_n1850_n1488# 0.382033f
C199 source.t30 a_n1850_n1488# 0.615866f
C200 source.n31 a_n1850_n1488# 0.607914f
C201 source.n32 a_n1850_n1488# 0.906799f
C202 minus.n0 a_n1850_n1488# 0.038128f
C203 minus.t14 a_n1850_n1488# 0.103986f
C204 minus.t5 a_n1850_n1488# 0.099374f
C205 minus.t1 a_n1850_n1488# 0.099374f
C206 minus.n1 a_n1850_n1488# 0.057701f
C207 minus.n2 a_n1850_n1488# 0.038128f
C208 minus.t12 a_n1850_n1488# 0.099374f
C209 minus.t8 a_n1850_n1488# 0.099374f
C210 minus.t3 a_n1850_n1488# 0.099374f
C211 minus.n3 a_n1850_n1488# 0.057701f
C212 minus.n4 a_n1850_n1488# 0.081143f
C213 minus.t13 a_n1850_n1488# 0.099374f
C214 minus.t9 a_n1850_n1488# 0.103986f
C215 minus.n5 a_n1850_n1488# 0.068962f
C216 minus.n6 a_n1850_n1488# 0.057701f
C217 minus.n7 a_n1850_n1488# 0.014411f
C218 minus.n8 a_n1850_n1488# 0.013941f
C219 minus.n9 a_n1850_n1488# 0.038128f
C220 minus.n10 a_n1850_n1488# 0.038128f
C221 minus.n11 a_n1850_n1488# 0.015704f
C222 minus.n12 a_n1850_n1488# 0.057701f
C223 minus.n13 a_n1850_n1488# 0.015704f
C224 minus.n14 a_n1850_n1488# 0.057701f
C225 minus.n15 a_n1850_n1488# 0.015704f
C226 minus.n16 a_n1850_n1488# 0.038128f
C227 minus.n17 a_n1850_n1488# 0.038128f
C228 minus.n18 a_n1850_n1488# 0.013941f
C229 minus.n19 a_n1850_n1488# 0.014411f
C230 minus.n20 a_n1850_n1488# 0.057701f
C231 minus.n21 a_n1850_n1488# 0.068911f
C232 minus.n22 a_n1850_n1488# 0.949942f
C233 minus.n23 a_n1850_n1488# 0.038128f
C234 minus.t11 a_n1850_n1488# 0.099374f
C235 minus.t2 a_n1850_n1488# 0.099374f
C236 minus.n24 a_n1850_n1488# 0.057701f
C237 minus.n25 a_n1850_n1488# 0.038128f
C238 minus.t4 a_n1850_n1488# 0.099374f
C239 minus.t7 a_n1850_n1488# 0.099374f
C240 minus.t15 a_n1850_n1488# 0.099374f
C241 minus.n26 a_n1850_n1488# 0.057701f
C242 minus.n27 a_n1850_n1488# 0.081143f
C243 minus.t0 a_n1850_n1488# 0.099374f
C244 minus.t6 a_n1850_n1488# 0.103986f
C245 minus.n28 a_n1850_n1488# 0.068962f
C246 minus.n29 a_n1850_n1488# 0.057701f
C247 minus.n30 a_n1850_n1488# 0.014411f
C248 minus.n31 a_n1850_n1488# 0.013941f
C249 minus.n32 a_n1850_n1488# 0.038128f
C250 minus.n33 a_n1850_n1488# 0.038128f
C251 minus.n34 a_n1850_n1488# 0.015704f
C252 minus.n35 a_n1850_n1488# 0.057701f
C253 minus.n36 a_n1850_n1488# 0.015704f
C254 minus.n37 a_n1850_n1488# 0.057701f
C255 minus.n38 a_n1850_n1488# 0.015704f
C256 minus.n39 a_n1850_n1488# 0.038128f
C257 minus.n40 a_n1850_n1488# 0.038128f
C258 minus.n41 a_n1850_n1488# 0.013941f
C259 minus.n42 a_n1850_n1488# 0.014411f
C260 minus.n43 a_n1850_n1488# 0.057701f
C261 minus.t10 a_n1850_n1488# 0.103986f
C262 minus.n44 a_n1850_n1488# 0.068911f
C263 minus.n45 a_n1850_n1488# 0.246251f
C264 minus.n46 a_n1850_n1488# 1.17472f
.ends

