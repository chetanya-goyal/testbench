* NGSPICE file created from diffpair389.ext - technology: sky130A

.subckt diffpair389 minus drain_right drain_left source plus
X0 a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X1 drain_left.t23 plus.t0 source.t22 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X2 source.t19 plus.t1 drain_left.t22 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X3 source.t30 plus.t2 drain_left.t21 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X4 source.t44 minus.t0 drain_right.t23 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X5 drain_right.t22 minus.t1 source.t43 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X6 drain_left.t20 plus.t3 source.t31 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X7 source.t12 plus.t4 drain_left.t19 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X8 source.t34 plus.t5 drain_left.t18 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X9 drain_right.t21 minus.t2 source.t11 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X10 a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X11 drain_right.t20 minus.t3 source.t10 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X12 source.t15 plus.t6 drain_left.t17 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X13 drain_left.t16 plus.t7 source.t26 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X14 drain_right.t19 minus.t4 source.t46 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X15 drain_right.t18 minus.t5 source.t39 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X16 drain_right.t17 minus.t6 source.t0 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X17 source.t42 minus.t7 drain_right.t16 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X18 drain_left.t15 plus.t8 source.t28 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X19 source.t23 plus.t9 drain_left.t14 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X20 drain_left.t13 plus.t10 source.t20 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X21 drain_left.t12 plus.t11 source.t17 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X22 drain_left.t11 plus.t12 source.t32 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X23 source.t13 plus.t13 drain_left.t10 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X24 drain_right.t15 minus.t8 source.t2 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X25 drain_left.t9 plus.t14 source.t35 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X26 source.t16 plus.t15 drain_left.t8 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X27 drain_left.t7 plus.t16 source.t27 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X28 a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X29 drain_right.t14 minus.t9 source.t37 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X30 drain_right.t13 minus.t10 source.t40 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X31 a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X32 source.t7 minus.t11 drain_right.t12 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X33 drain_left.t6 plus.t17 source.t29 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X34 source.t36 minus.t12 drain_right.t11 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X35 source.t24 plus.t18 drain_left.t5 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X36 drain_left.t4 plus.t19 source.t21 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X37 source.t41 minus.t13 drain_right.t10 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X38 source.t18 plus.t20 drain_left.t3 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X39 source.t3 minus.t14 drain_right.t9 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X40 drain_right.t8 minus.t15 source.t38 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X41 source.t6 minus.t16 drain_right.t7 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X42 source.t9 minus.t17 drain_right.t6 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X43 source.t8 minus.t18 drain_right.t5 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X44 drain_right.t4 minus.t19 source.t47 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X45 source.t33 plus.t21 drain_left.t2 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X46 drain_left.t1 plus.t22 source.t25 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X47 source.t1 minus.t20 drain_right.t3 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X48 source.t45 minus.t21 drain_right.t2 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X49 drain_right.t1 minus.t22 source.t5 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X50 source.t4 minus.t23 drain_right.t0 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X51 source.t14 plus.t23 drain_left.t0 a_n3394_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
R0 plus.n11 plus.t5 392.334
R1 plus.n53 plus.t19 392.334
R2 plus.n40 plus.t0 365.976
R3 plus.n38 plus.t15 365.976
R4 plus.n2 plus.t3 365.976
R5 plus.n32 plus.t23 365.976
R6 plus.n4 plus.t11 365.976
R7 plus.n26 plus.t1 365.976
R8 plus.n6 plus.t16 365.976
R9 plus.n20 plus.t4 365.976
R10 plus.n8 plus.t14 365.976
R11 plus.n14 plus.t2 365.976
R12 plus.n10 plus.t17 365.976
R13 plus.n82 plus.t13 365.976
R14 plus.n80 plus.t10 365.976
R15 plus.n44 plus.t9 365.976
R16 plus.n74 plus.t8 365.976
R17 plus.n46 plus.t18 365.976
R18 plus.n68 plus.t22 365.976
R19 plus.n48 plus.t21 365.976
R20 plus.n62 plus.t7 365.976
R21 plus.n50 plus.t6 365.976
R22 plus.n56 plus.t12 365.976
R23 plus.n52 plus.t20 365.976
R24 plus.n13 plus.n12 161.3
R25 plus.n14 plus.n9 161.3
R26 plus.n16 plus.n15 161.3
R27 plus.n17 plus.n8 161.3
R28 plus.n19 plus.n18 161.3
R29 plus.n20 plus.n7 161.3
R30 plus.n22 plus.n21 161.3
R31 plus.n23 plus.n6 161.3
R32 plus.n25 plus.n24 161.3
R33 plus.n26 plus.n5 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n4 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n32 plus.n3 161.3
R38 plus.n34 plus.n33 161.3
R39 plus.n35 plus.n2 161.3
R40 plus.n37 plus.n36 161.3
R41 plus.n38 plus.n1 161.3
R42 plus.n39 plus.n0 161.3
R43 plus.n41 plus.n40 161.3
R44 plus.n55 plus.n54 161.3
R45 plus.n56 plus.n51 161.3
R46 plus.n58 plus.n57 161.3
R47 plus.n59 plus.n50 161.3
R48 plus.n61 plus.n60 161.3
R49 plus.n62 plus.n49 161.3
R50 plus.n64 plus.n63 161.3
R51 plus.n65 plus.n48 161.3
R52 plus.n67 plus.n66 161.3
R53 plus.n68 plus.n47 161.3
R54 plus.n70 plus.n69 161.3
R55 plus.n71 plus.n46 161.3
R56 plus.n73 plus.n72 161.3
R57 plus.n74 plus.n45 161.3
R58 plus.n76 plus.n75 161.3
R59 plus.n77 plus.n44 161.3
R60 plus.n79 plus.n78 161.3
R61 plus.n80 plus.n43 161.3
R62 plus.n81 plus.n42 161.3
R63 plus.n83 plus.n82 161.3
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus.n33 plus.n2 37.246
R73 plus.n15 plus.n14 37.246
R74 plus.n75 plus.n44 37.246
R75 plus.n57 plus.n56 37.246
R76 plus plus.n83 34.9005
R77 plus.n32 plus.n31 32.8641
R78 plus.n19 plus.n8 32.8641
R79 plus.n74 plus.n73 32.8641
R80 plus.n61 plus.n50 32.8641
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus.n31 plus.n4 15.3369
R94 plus.n20 plus.n19 15.3369
R95 plus.n73 plus.n46 15.3369
R96 plus.n62 plus.n61 15.3369
R97 plus.n11 plus.n10 14.1472
R98 plus.n53 plus.n52 14.1472
R99 plus plus.n41 11.1861
R100 plus.n33 plus.n32 10.955
R101 plus.n15 plus.n8 10.955
R102 plus.n75 plus.n74 10.955
R103 plus.n57 plus.n50 10.955
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 source.n11 source.t34 51.0588
R149 source.n12 source.t40 51.0588
R150 source.n23 source.t36 51.0588
R151 source.n47 source.t47 51.0586
R152 source.n36 source.t4 51.0586
R153 source.n35 source.t21 51.0586
R154 source.n24 source.t13 51.0586
R155 source.n0 source.t22 51.0586
R156 source.n2 source.n1 48.8588
R157 source.n4 source.n3 48.8588
R158 source.n6 source.n5 48.8588
R159 source.n8 source.n7 48.8588
R160 source.n10 source.n9 48.8588
R161 source.n14 source.n13 48.8588
R162 source.n16 source.n15 48.8588
R163 source.n18 source.n17 48.8588
R164 source.n20 source.n19 48.8588
R165 source.n22 source.n21 48.8588
R166 source.n46 source.n45 48.8586
R167 source.n44 source.n43 48.8586
R168 source.n42 source.n41 48.8586
R169 source.n40 source.n39 48.8586
R170 source.n38 source.n37 48.8586
R171 source.n34 source.n33 48.8586
R172 source.n32 source.n31 48.8586
R173 source.n30 source.n29 48.8586
R174 source.n28 source.n27 48.8586
R175 source.n26 source.n25 48.8586
R176 source.n24 source.n23 19.9029
R177 source.n48 source.n0 14.196
R178 source.n48 source.n47 5.7074
R179 source.n45 source.t43 2.2005
R180 source.n45 source.t9 2.2005
R181 source.n43 source.t39 2.2005
R182 source.n43 source.t42 2.2005
R183 source.n41 source.t37 2.2005
R184 source.n41 source.t7 2.2005
R185 source.n39 source.t38 2.2005
R186 source.n39 source.t8 2.2005
R187 source.n37 source.t5 2.2005
R188 source.n37 source.t41 2.2005
R189 source.n33 source.t32 2.2005
R190 source.n33 source.t18 2.2005
R191 source.n31 source.t26 2.2005
R192 source.n31 source.t15 2.2005
R193 source.n29 source.t25 2.2005
R194 source.n29 source.t33 2.2005
R195 source.n27 source.t28 2.2005
R196 source.n27 source.t24 2.2005
R197 source.n25 source.t20 2.2005
R198 source.n25 source.t23 2.2005
R199 source.n1 source.t31 2.2005
R200 source.n1 source.t16 2.2005
R201 source.n3 source.t17 2.2005
R202 source.n3 source.t14 2.2005
R203 source.n5 source.t27 2.2005
R204 source.n5 source.t19 2.2005
R205 source.n7 source.t35 2.2005
R206 source.n7 source.t12 2.2005
R207 source.n9 source.t29 2.2005
R208 source.n9 source.t30 2.2005
R209 source.n13 source.t2 2.2005
R210 source.n13 source.t44 2.2005
R211 source.n15 source.t0 2.2005
R212 source.n15 source.t1 2.2005
R213 source.n17 source.t46 2.2005
R214 source.n17 source.t45 2.2005
R215 source.n19 source.t10 2.2005
R216 source.n19 source.t6 2.2005
R217 source.n21 source.t11 2.2005
R218 source.n21 source.t3 2.2005
R219 source.n23 source.n22 0.888431
R220 source.n22 source.n20 0.888431
R221 source.n20 source.n18 0.888431
R222 source.n18 source.n16 0.888431
R223 source.n16 source.n14 0.888431
R224 source.n14 source.n12 0.888431
R225 source.n11 source.n10 0.888431
R226 source.n10 source.n8 0.888431
R227 source.n8 source.n6 0.888431
R228 source.n6 source.n4 0.888431
R229 source.n4 source.n2 0.888431
R230 source.n2 source.n0 0.888431
R231 source.n26 source.n24 0.888431
R232 source.n28 source.n26 0.888431
R233 source.n30 source.n28 0.888431
R234 source.n32 source.n30 0.888431
R235 source.n34 source.n32 0.888431
R236 source.n35 source.n34 0.888431
R237 source.n38 source.n36 0.888431
R238 source.n40 source.n38 0.888431
R239 source.n42 source.n40 0.888431
R240 source.n44 source.n42 0.888431
R241 source.n46 source.n44 0.888431
R242 source.n47 source.n46 0.888431
R243 source.n12 source.n11 0.470328
R244 source.n36 source.n35 0.470328
R245 source source.n48 0.188
R246 drain_left.n13 drain_left.n11 66.4255
R247 drain_left.n7 drain_left.n5 66.4253
R248 drain_left.n2 drain_left.n0 66.4253
R249 drain_left.n19 drain_left.n18 65.5376
R250 drain_left.n17 drain_left.n16 65.5376
R251 drain_left.n15 drain_left.n14 65.5376
R252 drain_left.n13 drain_left.n12 65.5376
R253 drain_left.n21 drain_left.n20 65.5374
R254 drain_left.n7 drain_left.n6 65.5373
R255 drain_left.n9 drain_left.n8 65.5373
R256 drain_left.n4 drain_left.n3 65.5373
R257 drain_left.n2 drain_left.n1 65.5373
R258 drain_left drain_left.n10 33.5297
R259 drain_left drain_left.n21 6.54115
R260 drain_left.n5 drain_left.t3 2.2005
R261 drain_left.n5 drain_left.t4 2.2005
R262 drain_left.n6 drain_left.t17 2.2005
R263 drain_left.n6 drain_left.t11 2.2005
R264 drain_left.n8 drain_left.t2 2.2005
R265 drain_left.n8 drain_left.t16 2.2005
R266 drain_left.n3 drain_left.t5 2.2005
R267 drain_left.n3 drain_left.t1 2.2005
R268 drain_left.n1 drain_left.t14 2.2005
R269 drain_left.n1 drain_left.t15 2.2005
R270 drain_left.n0 drain_left.t10 2.2005
R271 drain_left.n0 drain_left.t13 2.2005
R272 drain_left.n20 drain_left.t8 2.2005
R273 drain_left.n20 drain_left.t23 2.2005
R274 drain_left.n18 drain_left.t0 2.2005
R275 drain_left.n18 drain_left.t20 2.2005
R276 drain_left.n16 drain_left.t22 2.2005
R277 drain_left.n16 drain_left.t12 2.2005
R278 drain_left.n14 drain_left.t19 2.2005
R279 drain_left.n14 drain_left.t7 2.2005
R280 drain_left.n12 drain_left.t21 2.2005
R281 drain_left.n12 drain_left.t9 2.2005
R282 drain_left.n11 drain_left.t18 2.2005
R283 drain_left.n11 drain_left.t6 2.2005
R284 drain_left.n9 drain_left.n7 0.888431
R285 drain_left.n4 drain_left.n2 0.888431
R286 drain_left.n15 drain_left.n13 0.888431
R287 drain_left.n17 drain_left.n15 0.888431
R288 drain_left.n19 drain_left.n17 0.888431
R289 drain_left.n21 drain_left.n19 0.888431
R290 drain_left.n10 drain_left.n9 0.389119
R291 drain_left.n10 drain_left.n4 0.389119
R292 minus.n11 minus.t10 392.334
R293 minus.n53 minus.t23 392.334
R294 minus.n10 minus.t0 365.976
R295 minus.n14 minus.t8 365.976
R296 minus.n16 minus.t20 365.976
R297 minus.n20 minus.t6 365.976
R298 minus.n22 minus.t21 365.976
R299 minus.n26 minus.t4 365.976
R300 minus.n28 minus.t16 365.976
R301 minus.n32 minus.t3 365.976
R302 minus.n34 minus.t14 365.976
R303 minus.n38 minus.t2 365.976
R304 minus.n40 minus.t12 365.976
R305 minus.n52 minus.t22 365.976
R306 minus.n56 minus.t13 365.976
R307 minus.n58 minus.t15 365.976
R308 minus.n62 minus.t18 365.976
R309 minus.n64 minus.t9 365.976
R310 minus.n68 minus.t11 365.976
R311 minus.n70 minus.t5 365.976
R312 minus.n74 minus.t7 365.976
R313 minus.n76 minus.t1 365.976
R314 minus.n80 minus.t17 365.976
R315 minus.n82 minus.t19 365.976
R316 minus.n41 minus.n40 161.3
R317 minus.n39 minus.n0 161.3
R318 minus.n38 minus.n37 161.3
R319 minus.n36 minus.n1 161.3
R320 minus.n35 minus.n34 161.3
R321 minus.n33 minus.n2 161.3
R322 minus.n32 minus.n31 161.3
R323 minus.n30 minus.n3 161.3
R324 minus.n29 minus.n28 161.3
R325 minus.n27 minus.n4 161.3
R326 minus.n26 minus.n25 161.3
R327 minus.n24 minus.n5 161.3
R328 minus.n23 minus.n22 161.3
R329 minus.n21 minus.n6 161.3
R330 minus.n20 minus.n19 161.3
R331 minus.n18 minus.n7 161.3
R332 minus.n17 minus.n16 161.3
R333 minus.n15 minus.n8 161.3
R334 minus.n14 minus.n13 161.3
R335 minus.n12 minus.n9 161.3
R336 minus.n83 minus.n82 161.3
R337 minus.n81 minus.n42 161.3
R338 minus.n80 minus.n79 161.3
R339 minus.n78 minus.n43 161.3
R340 minus.n77 minus.n76 161.3
R341 minus.n75 minus.n44 161.3
R342 minus.n74 minus.n73 161.3
R343 minus.n72 minus.n45 161.3
R344 minus.n71 minus.n70 161.3
R345 minus.n69 minus.n46 161.3
R346 minus.n68 minus.n67 161.3
R347 minus.n66 minus.n47 161.3
R348 minus.n65 minus.n64 161.3
R349 minus.n63 minus.n48 161.3
R350 minus.n62 minus.n61 161.3
R351 minus.n60 minus.n49 161.3
R352 minus.n59 minus.n58 161.3
R353 minus.n57 minus.n50 161.3
R354 minus.n56 minus.n55 161.3
R355 minus.n54 minus.n51 161.3
R356 minus.n40 minus.n39 46.0096
R357 minus.n82 minus.n81 46.0096
R358 minus.n12 minus.n11 45.0871
R359 minus.n54 minus.n53 45.0871
R360 minus.n10 minus.n9 41.6278
R361 minus.n38 minus.n1 41.6278
R362 minus.n52 minus.n51 41.6278
R363 minus.n80 minus.n43 41.6278
R364 minus.n84 minus.n41 39.8831
R365 minus.n15 minus.n14 37.246
R366 minus.n34 minus.n33 37.246
R367 minus.n57 minus.n56 37.246
R368 minus.n76 minus.n75 37.246
R369 minus.n16 minus.n7 32.8641
R370 minus.n32 minus.n3 32.8641
R371 minus.n58 minus.n49 32.8641
R372 minus.n74 minus.n45 32.8641
R373 minus.n21 minus.n20 28.4823
R374 minus.n28 minus.n27 28.4823
R375 minus.n63 minus.n62 28.4823
R376 minus.n70 minus.n69 28.4823
R377 minus.n26 minus.n5 24.1005
R378 minus.n22 minus.n5 24.1005
R379 minus.n64 minus.n47 24.1005
R380 minus.n68 minus.n47 24.1005
R381 minus.n22 minus.n21 19.7187
R382 minus.n27 minus.n26 19.7187
R383 minus.n64 minus.n63 19.7187
R384 minus.n69 minus.n68 19.7187
R385 minus.n20 minus.n7 15.3369
R386 minus.n28 minus.n3 15.3369
R387 minus.n62 minus.n49 15.3369
R388 minus.n70 minus.n45 15.3369
R389 minus.n11 minus.n10 14.1472
R390 minus.n53 minus.n52 14.1472
R391 minus.n16 minus.n15 10.955
R392 minus.n33 minus.n32 10.955
R393 minus.n58 minus.n57 10.955
R394 minus.n75 minus.n74 10.955
R395 minus.n84 minus.n83 6.67853
R396 minus.n14 minus.n9 6.57323
R397 minus.n34 minus.n1 6.57323
R398 minus.n56 minus.n51 6.57323
R399 minus.n76 minus.n43 6.57323
R400 minus.n39 minus.n38 2.19141
R401 minus.n81 minus.n80 2.19141
R402 minus.n41 minus.n0 0.189894
R403 minus.n37 minus.n0 0.189894
R404 minus.n37 minus.n36 0.189894
R405 minus.n36 minus.n35 0.189894
R406 minus.n35 minus.n2 0.189894
R407 minus.n31 minus.n2 0.189894
R408 minus.n31 minus.n30 0.189894
R409 minus.n30 minus.n29 0.189894
R410 minus.n29 minus.n4 0.189894
R411 minus.n25 minus.n4 0.189894
R412 minus.n25 minus.n24 0.189894
R413 minus.n24 minus.n23 0.189894
R414 minus.n23 minus.n6 0.189894
R415 minus.n19 minus.n6 0.189894
R416 minus.n19 minus.n18 0.189894
R417 minus.n18 minus.n17 0.189894
R418 minus.n17 minus.n8 0.189894
R419 minus.n13 minus.n8 0.189894
R420 minus.n13 minus.n12 0.189894
R421 minus.n55 minus.n54 0.189894
R422 minus.n55 minus.n50 0.189894
R423 minus.n59 minus.n50 0.189894
R424 minus.n60 minus.n59 0.189894
R425 minus.n61 minus.n60 0.189894
R426 minus.n61 minus.n48 0.189894
R427 minus.n65 minus.n48 0.189894
R428 minus.n66 minus.n65 0.189894
R429 minus.n67 minus.n66 0.189894
R430 minus.n67 minus.n46 0.189894
R431 minus.n71 minus.n46 0.189894
R432 minus.n72 minus.n71 0.189894
R433 minus.n73 minus.n72 0.189894
R434 minus.n73 minus.n44 0.189894
R435 minus.n77 minus.n44 0.189894
R436 minus.n78 minus.n77 0.189894
R437 minus.n79 minus.n78 0.189894
R438 minus.n79 minus.n42 0.189894
R439 minus.n83 minus.n42 0.189894
R440 minus minus.n84 0.188
R441 drain_right.n13 drain_right.n11 66.4254
R442 drain_right.n7 drain_right.n5 66.4253
R443 drain_right.n2 drain_right.n0 66.4253
R444 drain_right.n13 drain_right.n12 65.5376
R445 drain_right.n15 drain_right.n14 65.5376
R446 drain_right.n17 drain_right.n16 65.5376
R447 drain_right.n19 drain_right.n18 65.5376
R448 drain_right.n21 drain_right.n20 65.5376
R449 drain_right.n7 drain_right.n6 65.5373
R450 drain_right.n9 drain_right.n8 65.5373
R451 drain_right.n4 drain_right.n3 65.5373
R452 drain_right.n2 drain_right.n1 65.5373
R453 drain_right drain_right.n10 32.9765
R454 drain_right drain_right.n21 6.54115
R455 drain_right.n5 drain_right.t6 2.2005
R456 drain_right.n5 drain_right.t4 2.2005
R457 drain_right.n6 drain_right.t16 2.2005
R458 drain_right.n6 drain_right.t22 2.2005
R459 drain_right.n8 drain_right.t12 2.2005
R460 drain_right.n8 drain_right.t18 2.2005
R461 drain_right.n3 drain_right.t5 2.2005
R462 drain_right.n3 drain_right.t14 2.2005
R463 drain_right.n1 drain_right.t10 2.2005
R464 drain_right.n1 drain_right.t8 2.2005
R465 drain_right.n0 drain_right.t0 2.2005
R466 drain_right.n0 drain_right.t1 2.2005
R467 drain_right.n11 drain_right.t23 2.2005
R468 drain_right.n11 drain_right.t13 2.2005
R469 drain_right.n12 drain_right.t3 2.2005
R470 drain_right.n12 drain_right.t15 2.2005
R471 drain_right.n14 drain_right.t2 2.2005
R472 drain_right.n14 drain_right.t17 2.2005
R473 drain_right.n16 drain_right.t7 2.2005
R474 drain_right.n16 drain_right.t19 2.2005
R475 drain_right.n18 drain_right.t9 2.2005
R476 drain_right.n18 drain_right.t20 2.2005
R477 drain_right.n20 drain_right.t11 2.2005
R478 drain_right.n20 drain_right.t21 2.2005
R479 drain_right.n9 drain_right.n7 0.888431
R480 drain_right.n4 drain_right.n2 0.888431
R481 drain_right.n21 drain_right.n19 0.888431
R482 drain_right.n19 drain_right.n17 0.888431
R483 drain_right.n17 drain_right.n15 0.888431
R484 drain_right.n15 drain_right.n13 0.888431
R485 drain_right.n10 drain_right.n9 0.389119
R486 drain_right.n10 drain_right.n4 0.389119
C0 drain_right drain_left 1.87044f
C1 source plus 11.8215f
C2 drain_left plus 11.741f
C3 source minus 11.807401f
C4 drain_right plus 0.498726f
C5 drain_left minus 0.174517f
C6 drain_right minus 11.400599f
C7 drain_left source 22.4569f
C8 drain_right source 22.459501f
C9 minus plus 6.82534f
C10 drain_right a_n3394_n2688# 7.33929f
C11 drain_left a_n3394_n2688# 7.80975f
C12 source a_n3394_n2688# 7.915828f
C13 minus a_n3394_n2688# 13.543802f
C14 plus a_n3394_n2688# 15.28662f
C15 drain_right.t0 a_n3394_n2688# 0.19333f
C16 drain_right.t1 a_n3394_n2688# 0.19333f
C17 drain_right.n0 a_n3394_n2688# 1.69613f
C18 drain_right.t10 a_n3394_n2688# 0.19333f
C19 drain_right.t8 a_n3394_n2688# 0.19333f
C20 drain_right.n1 a_n3394_n2688# 1.69099f
C21 drain_right.n2 a_n3394_n2688# 0.752395f
C22 drain_right.t5 a_n3394_n2688# 0.19333f
C23 drain_right.t14 a_n3394_n2688# 0.19333f
C24 drain_right.n3 a_n3394_n2688# 1.69099f
C25 drain_right.n4 a_n3394_n2688# 0.331178f
C26 drain_right.t6 a_n3394_n2688# 0.19333f
C27 drain_right.t4 a_n3394_n2688# 0.19333f
C28 drain_right.n5 a_n3394_n2688# 1.69613f
C29 drain_right.t16 a_n3394_n2688# 0.19333f
C30 drain_right.t22 a_n3394_n2688# 0.19333f
C31 drain_right.n6 a_n3394_n2688# 1.69099f
C32 drain_right.n7 a_n3394_n2688# 0.752396f
C33 drain_right.t12 a_n3394_n2688# 0.19333f
C34 drain_right.t18 a_n3394_n2688# 0.19333f
C35 drain_right.n8 a_n3394_n2688# 1.69099f
C36 drain_right.n9 a_n3394_n2688# 0.331178f
C37 drain_right.n10 a_n3394_n2688# 1.55333f
C38 drain_right.t23 a_n3394_n2688# 0.19333f
C39 drain_right.t13 a_n3394_n2688# 0.19333f
C40 drain_right.n11 a_n3394_n2688# 1.69613f
C41 drain_right.t3 a_n3394_n2688# 0.19333f
C42 drain_right.t15 a_n3394_n2688# 0.19333f
C43 drain_right.n12 a_n3394_n2688# 1.691f
C44 drain_right.n13 a_n3394_n2688# 0.752396f
C45 drain_right.t2 a_n3394_n2688# 0.19333f
C46 drain_right.t17 a_n3394_n2688# 0.19333f
C47 drain_right.n14 a_n3394_n2688# 1.691f
C48 drain_right.n15 a_n3394_n2688# 0.373288f
C49 drain_right.t7 a_n3394_n2688# 0.19333f
C50 drain_right.t19 a_n3394_n2688# 0.19333f
C51 drain_right.n16 a_n3394_n2688# 1.691f
C52 drain_right.n17 a_n3394_n2688# 0.373288f
C53 drain_right.t9 a_n3394_n2688# 0.19333f
C54 drain_right.t20 a_n3394_n2688# 0.19333f
C55 drain_right.n18 a_n3394_n2688# 1.691f
C56 drain_right.n19 a_n3394_n2688# 0.373288f
C57 drain_right.t11 a_n3394_n2688# 0.19333f
C58 drain_right.t21 a_n3394_n2688# 0.19333f
C59 drain_right.n20 a_n3394_n2688# 1.691f
C60 drain_right.n21 a_n3394_n2688# 0.613727f
C61 minus.n0 a_n3394_n2688# 0.03929f
C62 minus.n1 a_n3394_n2688# 0.008916f
C63 minus.t2 a_n3394_n2688# 0.709881f
C64 minus.n2 a_n3394_n2688# 0.03929f
C65 minus.n3 a_n3394_n2688# 0.008916f
C66 minus.t3 a_n3394_n2688# 0.709881f
C67 minus.n4 a_n3394_n2688# 0.03929f
C68 minus.n5 a_n3394_n2688# 0.008916f
C69 minus.t4 a_n3394_n2688# 0.709881f
C70 minus.n6 a_n3394_n2688# 0.03929f
C71 minus.n7 a_n3394_n2688# 0.008916f
C72 minus.t6 a_n3394_n2688# 0.709881f
C73 minus.n8 a_n3394_n2688# 0.03929f
C74 minus.n9 a_n3394_n2688# 0.008916f
C75 minus.t8 a_n3394_n2688# 0.709881f
C76 minus.t10 a_n3394_n2688# 0.729965f
C77 minus.t0 a_n3394_n2688# 0.709881f
C78 minus.n10 a_n3394_n2688# 0.306297f
C79 minus.n11 a_n3394_n2688# 0.280264f
C80 minus.n12 a_n3394_n2688# 0.169147f
C81 minus.n13 a_n3394_n2688# 0.03929f
C82 minus.n14 a_n3394_n2688# 0.298256f
C83 minus.n15 a_n3394_n2688# 0.008916f
C84 minus.t20 a_n3394_n2688# 0.709881f
C85 minus.n16 a_n3394_n2688# 0.298256f
C86 minus.n17 a_n3394_n2688# 0.03929f
C87 minus.n18 a_n3394_n2688# 0.03929f
C88 minus.n19 a_n3394_n2688# 0.03929f
C89 minus.n20 a_n3394_n2688# 0.298256f
C90 minus.n21 a_n3394_n2688# 0.008916f
C91 minus.t21 a_n3394_n2688# 0.709881f
C92 minus.n22 a_n3394_n2688# 0.298256f
C93 minus.n23 a_n3394_n2688# 0.03929f
C94 minus.n24 a_n3394_n2688# 0.03929f
C95 minus.n25 a_n3394_n2688# 0.03929f
C96 minus.n26 a_n3394_n2688# 0.298256f
C97 minus.n27 a_n3394_n2688# 0.008916f
C98 minus.t16 a_n3394_n2688# 0.709881f
C99 minus.n28 a_n3394_n2688# 0.298256f
C100 minus.n29 a_n3394_n2688# 0.03929f
C101 minus.n30 a_n3394_n2688# 0.03929f
C102 minus.n31 a_n3394_n2688# 0.03929f
C103 minus.n32 a_n3394_n2688# 0.298256f
C104 minus.n33 a_n3394_n2688# 0.008916f
C105 minus.t14 a_n3394_n2688# 0.709881f
C106 minus.n34 a_n3394_n2688# 0.298256f
C107 minus.n35 a_n3394_n2688# 0.03929f
C108 minus.n36 a_n3394_n2688# 0.03929f
C109 minus.n37 a_n3394_n2688# 0.03929f
C110 minus.n38 a_n3394_n2688# 0.298256f
C111 minus.n39 a_n3394_n2688# 0.008916f
C112 minus.t12 a_n3394_n2688# 0.709881f
C113 minus.n40 a_n3394_n2688# 0.29862f
C114 minus.n41 a_n3394_n2688# 1.61613f
C115 minus.n42 a_n3394_n2688# 0.03929f
C116 minus.n43 a_n3394_n2688# 0.008916f
C117 minus.n44 a_n3394_n2688# 0.03929f
C118 minus.n45 a_n3394_n2688# 0.008916f
C119 minus.n46 a_n3394_n2688# 0.03929f
C120 minus.n47 a_n3394_n2688# 0.008916f
C121 minus.n48 a_n3394_n2688# 0.03929f
C122 minus.n49 a_n3394_n2688# 0.008916f
C123 minus.n50 a_n3394_n2688# 0.03929f
C124 minus.n51 a_n3394_n2688# 0.008916f
C125 minus.t23 a_n3394_n2688# 0.729965f
C126 minus.t22 a_n3394_n2688# 0.709881f
C127 minus.n52 a_n3394_n2688# 0.306297f
C128 minus.n53 a_n3394_n2688# 0.280264f
C129 minus.n54 a_n3394_n2688# 0.169147f
C130 minus.n55 a_n3394_n2688# 0.03929f
C131 minus.t13 a_n3394_n2688# 0.709881f
C132 minus.n56 a_n3394_n2688# 0.298256f
C133 minus.n57 a_n3394_n2688# 0.008916f
C134 minus.t15 a_n3394_n2688# 0.709881f
C135 minus.n58 a_n3394_n2688# 0.298256f
C136 minus.n59 a_n3394_n2688# 0.03929f
C137 minus.n60 a_n3394_n2688# 0.03929f
C138 minus.n61 a_n3394_n2688# 0.03929f
C139 minus.t18 a_n3394_n2688# 0.709881f
C140 minus.n62 a_n3394_n2688# 0.298256f
C141 minus.n63 a_n3394_n2688# 0.008916f
C142 minus.t9 a_n3394_n2688# 0.709881f
C143 minus.n64 a_n3394_n2688# 0.298256f
C144 minus.n65 a_n3394_n2688# 0.03929f
C145 minus.n66 a_n3394_n2688# 0.03929f
C146 minus.n67 a_n3394_n2688# 0.03929f
C147 minus.t11 a_n3394_n2688# 0.709881f
C148 minus.n68 a_n3394_n2688# 0.298256f
C149 minus.n69 a_n3394_n2688# 0.008916f
C150 minus.t5 a_n3394_n2688# 0.709881f
C151 minus.n70 a_n3394_n2688# 0.298256f
C152 minus.n71 a_n3394_n2688# 0.03929f
C153 minus.n72 a_n3394_n2688# 0.03929f
C154 minus.n73 a_n3394_n2688# 0.03929f
C155 minus.t7 a_n3394_n2688# 0.709881f
C156 minus.n74 a_n3394_n2688# 0.298256f
C157 minus.n75 a_n3394_n2688# 0.008916f
C158 minus.t1 a_n3394_n2688# 0.709881f
C159 minus.n76 a_n3394_n2688# 0.298256f
C160 minus.n77 a_n3394_n2688# 0.03929f
C161 minus.n78 a_n3394_n2688# 0.03929f
C162 minus.n79 a_n3394_n2688# 0.03929f
C163 minus.t17 a_n3394_n2688# 0.709881f
C164 minus.n80 a_n3394_n2688# 0.298256f
C165 minus.n81 a_n3394_n2688# 0.008916f
C166 minus.t19 a_n3394_n2688# 0.709881f
C167 minus.n82 a_n3394_n2688# 0.29862f
C168 minus.n83 a_n3394_n2688# 0.27326f
C169 minus.n84 a_n3394_n2688# 1.93747f
C170 drain_left.t10 a_n3394_n2688# 0.194431f
C171 drain_left.t13 a_n3394_n2688# 0.194431f
C172 drain_left.n0 a_n3394_n2688# 1.70579f
C173 drain_left.t14 a_n3394_n2688# 0.194431f
C174 drain_left.t15 a_n3394_n2688# 0.194431f
C175 drain_left.n1 a_n3394_n2688# 1.70062f
C176 drain_left.n2 a_n3394_n2688# 0.75668f
C177 drain_left.t5 a_n3394_n2688# 0.194431f
C178 drain_left.t1 a_n3394_n2688# 0.194431f
C179 drain_left.n3 a_n3394_n2688# 1.70062f
C180 drain_left.n4 a_n3394_n2688# 0.333064f
C181 drain_left.t3 a_n3394_n2688# 0.194431f
C182 drain_left.t4 a_n3394_n2688# 0.194431f
C183 drain_left.n5 a_n3394_n2688# 1.70579f
C184 drain_left.t17 a_n3394_n2688# 0.194431f
C185 drain_left.t11 a_n3394_n2688# 0.194431f
C186 drain_left.n6 a_n3394_n2688# 1.70062f
C187 drain_left.n7 a_n3394_n2688# 0.75668f
C188 drain_left.t2 a_n3394_n2688# 0.194431f
C189 drain_left.t16 a_n3394_n2688# 0.194431f
C190 drain_left.n8 a_n3394_n2688# 1.70062f
C191 drain_left.n9 a_n3394_n2688# 0.333064f
C192 drain_left.n10 a_n3394_n2688# 1.61711f
C193 drain_left.t18 a_n3394_n2688# 0.194431f
C194 drain_left.t6 a_n3394_n2688# 0.194431f
C195 drain_left.n11 a_n3394_n2688# 1.70579f
C196 drain_left.t21 a_n3394_n2688# 0.194431f
C197 drain_left.t9 a_n3394_n2688# 0.194431f
C198 drain_left.n12 a_n3394_n2688# 1.70063f
C199 drain_left.n13 a_n3394_n2688# 0.756674f
C200 drain_left.t19 a_n3394_n2688# 0.194431f
C201 drain_left.t7 a_n3394_n2688# 0.194431f
C202 drain_left.n14 a_n3394_n2688# 1.70063f
C203 drain_left.n15 a_n3394_n2688# 0.375414f
C204 drain_left.t22 a_n3394_n2688# 0.194431f
C205 drain_left.t12 a_n3394_n2688# 0.194431f
C206 drain_left.n16 a_n3394_n2688# 1.70063f
C207 drain_left.n17 a_n3394_n2688# 0.375414f
C208 drain_left.t0 a_n3394_n2688# 0.194431f
C209 drain_left.t20 a_n3394_n2688# 0.194431f
C210 drain_left.n18 a_n3394_n2688# 1.70063f
C211 drain_left.n19 a_n3394_n2688# 0.375414f
C212 drain_left.t8 a_n3394_n2688# 0.194431f
C213 drain_left.t23 a_n3394_n2688# 0.194431f
C214 drain_left.n20 a_n3394_n2688# 1.70062f
C215 drain_left.n21 a_n3394_n2688# 0.617229f
C216 source.t22 a_n3394_n2688# 1.93132f
C217 source.n0 a_n3394_n2688# 1.15787f
C218 source.t31 a_n3394_n2688# 0.181115f
C219 source.t16 a_n3394_n2688# 0.181115f
C220 source.n1 a_n3394_n2688# 1.51618f
C221 source.n2 a_n3394_n2688# 0.383068f
C222 source.t17 a_n3394_n2688# 0.181115f
C223 source.t14 a_n3394_n2688# 0.181115f
C224 source.n3 a_n3394_n2688# 1.51618f
C225 source.n4 a_n3394_n2688# 0.383068f
C226 source.t27 a_n3394_n2688# 0.181115f
C227 source.t19 a_n3394_n2688# 0.181115f
C228 source.n5 a_n3394_n2688# 1.51618f
C229 source.n6 a_n3394_n2688# 0.383068f
C230 source.t35 a_n3394_n2688# 0.181115f
C231 source.t12 a_n3394_n2688# 0.181115f
C232 source.n7 a_n3394_n2688# 1.51618f
C233 source.n8 a_n3394_n2688# 0.383068f
C234 source.t29 a_n3394_n2688# 0.181115f
C235 source.t30 a_n3394_n2688# 0.181115f
C236 source.n9 a_n3394_n2688# 1.51618f
C237 source.n10 a_n3394_n2688# 0.383068f
C238 source.t34 a_n3394_n2688# 1.93132f
C239 source.n11 a_n3394_n2688# 0.427568f
C240 source.t40 a_n3394_n2688# 1.93132f
C241 source.n12 a_n3394_n2688# 0.427568f
C242 source.t2 a_n3394_n2688# 0.181115f
C243 source.t44 a_n3394_n2688# 0.181115f
C244 source.n13 a_n3394_n2688# 1.51618f
C245 source.n14 a_n3394_n2688# 0.383068f
C246 source.t0 a_n3394_n2688# 0.181115f
C247 source.t1 a_n3394_n2688# 0.181115f
C248 source.n15 a_n3394_n2688# 1.51618f
C249 source.n16 a_n3394_n2688# 0.383068f
C250 source.t46 a_n3394_n2688# 0.181115f
C251 source.t45 a_n3394_n2688# 0.181115f
C252 source.n17 a_n3394_n2688# 1.51618f
C253 source.n18 a_n3394_n2688# 0.383068f
C254 source.t10 a_n3394_n2688# 0.181115f
C255 source.t6 a_n3394_n2688# 0.181115f
C256 source.n19 a_n3394_n2688# 1.51618f
C257 source.n20 a_n3394_n2688# 0.383068f
C258 source.t11 a_n3394_n2688# 0.181115f
C259 source.t3 a_n3394_n2688# 0.181115f
C260 source.n21 a_n3394_n2688# 1.51618f
C261 source.n22 a_n3394_n2688# 0.383068f
C262 source.t36 a_n3394_n2688# 1.93132f
C263 source.n23 a_n3394_n2688# 1.53716f
C264 source.t13 a_n3394_n2688# 1.93132f
C265 source.n24 a_n3394_n2688# 1.53717f
C266 source.t20 a_n3394_n2688# 0.181115f
C267 source.t23 a_n3394_n2688# 0.181115f
C268 source.n25 a_n3394_n2688# 1.51617f
C269 source.n26 a_n3394_n2688# 0.383072f
C270 source.t28 a_n3394_n2688# 0.181115f
C271 source.t24 a_n3394_n2688# 0.181115f
C272 source.n27 a_n3394_n2688# 1.51617f
C273 source.n28 a_n3394_n2688# 0.383072f
C274 source.t25 a_n3394_n2688# 0.181115f
C275 source.t33 a_n3394_n2688# 0.181115f
C276 source.n29 a_n3394_n2688# 1.51617f
C277 source.n30 a_n3394_n2688# 0.383072f
C278 source.t26 a_n3394_n2688# 0.181115f
C279 source.t15 a_n3394_n2688# 0.181115f
C280 source.n31 a_n3394_n2688# 1.51617f
C281 source.n32 a_n3394_n2688# 0.383072f
C282 source.t32 a_n3394_n2688# 0.181115f
C283 source.t18 a_n3394_n2688# 0.181115f
C284 source.n33 a_n3394_n2688# 1.51617f
C285 source.n34 a_n3394_n2688# 0.383072f
C286 source.t21 a_n3394_n2688# 1.93132f
C287 source.n35 a_n3394_n2688# 0.427573f
C288 source.t4 a_n3394_n2688# 1.93132f
C289 source.n36 a_n3394_n2688# 0.427573f
C290 source.t5 a_n3394_n2688# 0.181115f
C291 source.t41 a_n3394_n2688# 0.181115f
C292 source.n37 a_n3394_n2688# 1.51617f
C293 source.n38 a_n3394_n2688# 0.383072f
C294 source.t38 a_n3394_n2688# 0.181115f
C295 source.t8 a_n3394_n2688# 0.181115f
C296 source.n39 a_n3394_n2688# 1.51617f
C297 source.n40 a_n3394_n2688# 0.383072f
C298 source.t37 a_n3394_n2688# 0.181115f
C299 source.t7 a_n3394_n2688# 0.181115f
C300 source.n41 a_n3394_n2688# 1.51617f
C301 source.n42 a_n3394_n2688# 0.383072f
C302 source.t39 a_n3394_n2688# 0.181115f
C303 source.t42 a_n3394_n2688# 0.181115f
C304 source.n43 a_n3394_n2688# 1.51617f
C305 source.n44 a_n3394_n2688# 0.383072f
C306 source.t43 a_n3394_n2688# 0.181115f
C307 source.t9 a_n3394_n2688# 0.181115f
C308 source.n45 a_n3394_n2688# 1.51617f
C309 source.n46 a_n3394_n2688# 0.383072f
C310 source.t47 a_n3394_n2688# 1.93132f
C311 source.n47 a_n3394_n2688# 0.593688f
C312 source.n48 a_n3394_n2688# 1.34089f
C313 plus.n0 a_n3394_n2688# 0.039789f
C314 plus.t0 a_n3394_n2688# 0.718883f
C315 plus.t15 a_n3394_n2688# 0.718883f
C316 plus.n1 a_n3394_n2688# 0.039789f
C317 plus.t3 a_n3394_n2688# 0.718883f
C318 plus.n2 a_n3394_n2688# 0.302039f
C319 plus.n3 a_n3394_n2688# 0.039789f
C320 plus.t23 a_n3394_n2688# 0.718883f
C321 plus.t11 a_n3394_n2688# 0.718883f
C322 plus.n4 a_n3394_n2688# 0.302039f
C323 plus.n5 a_n3394_n2688# 0.039789f
C324 plus.t1 a_n3394_n2688# 0.718883f
C325 plus.t16 a_n3394_n2688# 0.718883f
C326 plus.n6 a_n3394_n2688# 0.302039f
C327 plus.n7 a_n3394_n2688# 0.039789f
C328 plus.t4 a_n3394_n2688# 0.718883f
C329 plus.t14 a_n3394_n2688# 0.718883f
C330 plus.n8 a_n3394_n2688# 0.302039f
C331 plus.n9 a_n3394_n2688# 0.039789f
C332 plus.t2 a_n3394_n2688# 0.718883f
C333 plus.t17 a_n3394_n2688# 0.718883f
C334 plus.n10 a_n3394_n2688# 0.310181f
C335 plus.t5 a_n3394_n2688# 0.739222f
C336 plus.n11 a_n3394_n2688# 0.283818f
C337 plus.n12 a_n3394_n2688# 0.171293f
C338 plus.n13 a_n3394_n2688# 0.009029f
C339 plus.n14 a_n3394_n2688# 0.302039f
C340 plus.n15 a_n3394_n2688# 0.009029f
C341 plus.n16 a_n3394_n2688# 0.039789f
C342 plus.n17 a_n3394_n2688# 0.039789f
C343 plus.n18 a_n3394_n2688# 0.039789f
C344 plus.n19 a_n3394_n2688# 0.009029f
C345 plus.n20 a_n3394_n2688# 0.302039f
C346 plus.n21 a_n3394_n2688# 0.009029f
C347 plus.n22 a_n3394_n2688# 0.039789f
C348 plus.n23 a_n3394_n2688# 0.039789f
C349 plus.n24 a_n3394_n2688# 0.039789f
C350 plus.n25 a_n3394_n2688# 0.009029f
C351 plus.n26 a_n3394_n2688# 0.302039f
C352 plus.n27 a_n3394_n2688# 0.009029f
C353 plus.n28 a_n3394_n2688# 0.039789f
C354 plus.n29 a_n3394_n2688# 0.039789f
C355 plus.n30 a_n3394_n2688# 0.039789f
C356 plus.n31 a_n3394_n2688# 0.009029f
C357 plus.n32 a_n3394_n2688# 0.302039f
C358 plus.n33 a_n3394_n2688# 0.009029f
C359 plus.n34 a_n3394_n2688# 0.039789f
C360 plus.n35 a_n3394_n2688# 0.039789f
C361 plus.n36 a_n3394_n2688# 0.039789f
C362 plus.n37 a_n3394_n2688# 0.009029f
C363 plus.n38 a_n3394_n2688# 0.302039f
C364 plus.n39 a_n3394_n2688# 0.009029f
C365 plus.n40 a_n3394_n2688# 0.302407f
C366 plus.n41 a_n3394_n2688# 0.407985f
C367 plus.n42 a_n3394_n2688# 0.039789f
C368 plus.t13 a_n3394_n2688# 0.718883f
C369 plus.n43 a_n3394_n2688# 0.039789f
C370 plus.t10 a_n3394_n2688# 0.718883f
C371 plus.t9 a_n3394_n2688# 0.718883f
C372 plus.n44 a_n3394_n2688# 0.302039f
C373 plus.n45 a_n3394_n2688# 0.039789f
C374 plus.t8 a_n3394_n2688# 0.718883f
C375 plus.t18 a_n3394_n2688# 0.718883f
C376 plus.n46 a_n3394_n2688# 0.302039f
C377 plus.n47 a_n3394_n2688# 0.039789f
C378 plus.t22 a_n3394_n2688# 0.718883f
C379 plus.t21 a_n3394_n2688# 0.718883f
C380 plus.n48 a_n3394_n2688# 0.302039f
C381 plus.n49 a_n3394_n2688# 0.039789f
C382 plus.t7 a_n3394_n2688# 0.718883f
C383 plus.t6 a_n3394_n2688# 0.718883f
C384 plus.n50 a_n3394_n2688# 0.302039f
C385 plus.n51 a_n3394_n2688# 0.039789f
C386 plus.t12 a_n3394_n2688# 0.718883f
C387 plus.t20 a_n3394_n2688# 0.718883f
C388 plus.n52 a_n3394_n2688# 0.310181f
C389 plus.t19 a_n3394_n2688# 0.739222f
C390 plus.n53 a_n3394_n2688# 0.283818f
C391 plus.n54 a_n3394_n2688# 0.171293f
C392 plus.n55 a_n3394_n2688# 0.009029f
C393 plus.n56 a_n3394_n2688# 0.302039f
C394 plus.n57 a_n3394_n2688# 0.009029f
C395 plus.n58 a_n3394_n2688# 0.039789f
C396 plus.n59 a_n3394_n2688# 0.039789f
C397 plus.n60 a_n3394_n2688# 0.039789f
C398 plus.n61 a_n3394_n2688# 0.009029f
C399 plus.n62 a_n3394_n2688# 0.302039f
C400 plus.n63 a_n3394_n2688# 0.009029f
C401 plus.n64 a_n3394_n2688# 0.039789f
C402 plus.n65 a_n3394_n2688# 0.039789f
C403 plus.n66 a_n3394_n2688# 0.039789f
C404 plus.n67 a_n3394_n2688# 0.009029f
C405 plus.n68 a_n3394_n2688# 0.302039f
C406 plus.n69 a_n3394_n2688# 0.009029f
C407 plus.n70 a_n3394_n2688# 0.039789f
C408 plus.n71 a_n3394_n2688# 0.039789f
C409 plus.n72 a_n3394_n2688# 0.039789f
C410 plus.n73 a_n3394_n2688# 0.009029f
C411 plus.n74 a_n3394_n2688# 0.302039f
C412 plus.n75 a_n3394_n2688# 0.009029f
C413 plus.n76 a_n3394_n2688# 0.039789f
C414 plus.n77 a_n3394_n2688# 0.039789f
C415 plus.n78 a_n3394_n2688# 0.039789f
C416 plus.n79 a_n3394_n2688# 0.009029f
C417 plus.n80 a_n3394_n2688# 0.302039f
C418 plus.n81 a_n3394_n2688# 0.009029f
C419 plus.n82 a_n3394_n2688# 0.302407f
C420 plus.n83 a_n3394_n2688# 1.44445f
.ends

