* NGSPICE file created from diffpair332.ext - technology: sky130A

.subckt diffpair332 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t6 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X1 drain_right.t4 minus.t1 source.t7 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 drain_right.t3 minus.t2 source.t8 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X3 source.t9 minus.t3 drain_right.t2 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 source.t4 plus.t0 drain_left.t5 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 source.t10 minus.t4 drain_right.t1 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X6 a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X7 a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X8 drain_left.t4 plus.t1 source.t5 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X9 a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X10 drain_right.t0 minus.t5 source.t11 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X11 drain_left.t3 plus.t2 source.t1 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X12 drain_left.t2 plus.t3 source.t3 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X13 a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X14 source.t2 plus.t4 drain_left.t1 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X15 drain_left.t0 plus.t5 source.t0 a_n1140_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
R0 minus.n2 minus.t2 1282.05
R1 minus.n0 minus.t5 1282.05
R2 minus.n6 minus.t0 1282.05
R3 minus.n4 minus.t1 1282.05
R4 minus.n1 minus.t4 1241.15
R5 minus.n5 minus.t3 1241.15
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 31.1047
R15 minus.n8 minus.n7 6.438
R16 minus minus.n8 0.188
R17 source.n3 source.t11 51.0588
R18 source.n11 source.t6 51.0586
R19 source.n8 source.t1 51.0586
R20 source.n0 source.t0 51.0586
R21 source.n2 source.n1 48.8588
R22 source.n5 source.n4 48.8588
R23 source.n10 source.n9 48.8586
R24 source.n7 source.n6 48.8586
R25 source.n7 source.n5 19.9288
R26 source.n12 source.n0 13.9805
R27 source.n12 source.n11 5.49188
R28 source.n9 source.t7 2.2005
R29 source.n9 source.t9 2.2005
R30 source.n6 source.t3 2.2005
R31 source.n6 source.t2 2.2005
R32 source.n1 source.t5 2.2005
R33 source.n1 source.t4 2.2005
R34 source.n4 source.t8 2.2005
R35 source.n4 source.t10 2.2005
R36 source.n3 source.n2 0.698776
R37 source.n10 source.n8 0.698776
R38 source.n5 source.n3 0.457397
R39 source.n2 source.n0 0.457397
R40 source.n8 source.n7 0.457397
R41 source.n11 source.n10 0.457397
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t4 68.0247
R44 drain_right.n3 drain_right.t3 67.7376
R45 drain_right.n3 drain_right.n2 65.9943
R46 drain_right.n1 drain_right.n0 65.5962
R47 drain_right drain_right.n1 25.7976
R48 drain_right drain_right.n3 5.88166
R49 drain_right.n0 drain_right.t2 2.2005
R50 drain_right.n0 drain_right.t5 2.2005
R51 drain_right.n2 drain_right.t1 2.2005
R52 drain_right.n2 drain_right.t0 2.2005
R53 plus.n0 plus.t1 1282.05
R54 plus.n2 plus.t5 1282.05
R55 plus.n4 plus.t2 1282.05
R56 plus.n6 plus.t3 1282.05
R57 plus.n1 plus.t0 1241.15
R58 plus.n5 plus.t4 1241.15
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 26.1221
R68 plus plus.n3 10.9456
R69 drain_left.n3 drain_left.t4 68.1945
R70 drain_left.n1 drain_left.t2 68.0247
R71 drain_left.n1 drain_left.n0 65.5962
R72 drain_left.n3 drain_left.n2 65.5374
R73 drain_left drain_left.n1 26.3508
R74 drain_left drain_left.n3 6.11011
R75 drain_left.n0 drain_left.t1 2.2005
R76 drain_left.n0 drain_left.t3 2.2005
R77 drain_left.n2 drain_left.t5 2.2005
R78 drain_left.n2 drain_left.t0 2.2005
C0 minus source 1.31729f
C1 drain_left plus 1.80806f
C2 drain_left drain_right 0.533726f
C3 drain_left source 12.704401f
C4 drain_right plus 0.26071f
C5 minus drain_left 0.170484f
C6 source plus 1.33186f
C7 minus plus 4.02058f
C8 source drain_right 12.694f
C9 minus drain_right 1.70445f
C10 drain_right a_n1140_n2688# 5.30698f
C11 drain_left a_n1140_n2688# 5.46525f
C12 source a_n1140_n2688# 4.927135f
C13 minus a_n1140_n2688# 4.152953f
C14 plus a_n1140_n2688# 5.15616f
C15 drain_left.t2 a_n1140_n2688# 2.10374f
C16 drain_left.t1 a_n1140_n2688# 0.188832f
C17 drain_left.t3 a_n1140_n2688# 0.188832f
C18 drain_left.n0 a_n1140_n2688# 1.6519f
C19 drain_left.n1 a_n1140_n2688# 1.5059f
C20 drain_left.t4 a_n1140_n2688# 2.1046f
C21 drain_left.t5 a_n1140_n2688# 0.188832f
C22 drain_left.t0 a_n1140_n2688# 0.188832f
C23 drain_left.n2 a_n1140_n2688# 1.65165f
C24 drain_left.n3 a_n1140_n2688# 0.832654f
C25 plus.t1 a_n1140_n2688# 0.180903f
C26 plus.n0 a_n1140_n2688# 0.087492f
C27 plus.t0 a_n1140_n2688# 0.178425f
C28 plus.n1 a_n1140_n2688# 0.078102f
C29 plus.t5 a_n1140_n2688# 0.180903f
C30 plus.n2 a_n1140_n2688# 0.087444f
C31 plus.n3 a_n1140_n2688# 0.378897f
C32 plus.t2 a_n1140_n2688# 0.180903f
C33 plus.n4 a_n1140_n2688# 0.087492f
C34 plus.t3 a_n1140_n2688# 0.180903f
C35 plus.t4 a_n1140_n2688# 0.178425f
C36 plus.n5 a_n1140_n2688# 0.078102f
C37 plus.n6 a_n1140_n2688# 0.087444f
C38 plus.n7 a_n1140_n2688# 0.880689f
C39 drain_right.t4 a_n1140_n2688# 2.12108f
C40 drain_right.t2 a_n1140_n2688# 0.190389f
C41 drain_right.t5 a_n1140_n2688# 0.190389f
C42 drain_right.n0 a_n1140_n2688# 1.66552f
C43 drain_right.n1 a_n1140_n2688# 1.46246f
C44 drain_right.t1 a_n1140_n2688# 0.190389f
C45 drain_right.t0 a_n1140_n2688# 0.190389f
C46 drain_right.n2 a_n1140_n2688# 1.66737f
C47 drain_right.t3 a_n1140_n2688# 2.11975f
C48 drain_right.n3 a_n1140_n2688# 0.848898f
C49 source.t0 a_n1140_n2688# 2.17356f
C50 source.n0 a_n1140_n2688# 1.23652f
C51 source.t5 a_n1140_n2688# 0.203833f
C52 source.t4 a_n1140_n2688# 0.203833f
C53 source.n1 a_n1140_n2688# 1.70635f
C54 source.n2 a_n1140_n2688# 0.373796f
C55 source.t11 a_n1140_n2688# 2.17357f
C56 source.n3 a_n1140_n2688# 0.46249f
C57 source.t8 a_n1140_n2688# 0.203833f
C58 source.t10 a_n1140_n2688# 0.203833f
C59 source.n4 a_n1140_n2688# 1.70635f
C60 source.n5 a_n1140_n2688# 1.60386f
C61 source.t3 a_n1140_n2688# 0.203833f
C62 source.t2 a_n1140_n2688# 0.203833f
C63 source.n6 a_n1140_n2688# 1.70635f
C64 source.n7 a_n1140_n2688# 1.60387f
C65 source.t1 a_n1140_n2688# 2.17356f
C66 source.n8 a_n1140_n2688# 0.462495f
C67 source.t7 a_n1140_n2688# 0.203833f
C68 source.t9 a_n1140_n2688# 0.203833f
C69 source.n9 a_n1140_n2688# 1.70635f
C70 source.n10 a_n1140_n2688# 0.373801f
C71 source.t6 a_n1140_n2688# 2.17356f
C72 source.n11 a_n1140_n2688# 0.596802f
C73 source.n12 a_n1140_n2688# 1.48779f
C74 minus.t5 a_n1140_n2688# 0.177759f
C75 minus.n0 a_n1140_n2688# 0.085972f
C76 minus.t2 a_n1140_n2688# 0.177759f
C77 minus.t4 a_n1140_n2688# 0.175324f
C78 minus.n1 a_n1140_n2688# 0.076744f
C79 minus.n2 a_n1140_n2688# 0.085925f
C80 minus.n3 a_n1140_n2688# 0.98856f
C81 minus.t1 a_n1140_n2688# 0.177759f
C82 minus.n4 a_n1140_n2688# 0.085972f
C83 minus.t3 a_n1140_n2688# 0.175324f
C84 minus.n5 a_n1140_n2688# 0.076744f
C85 minus.t0 a_n1140_n2688# 0.177759f
C86 minus.n6 a_n1140_n2688# 0.085925f
C87 minus.n7 a_n1140_n2688# 0.25953f
C88 minus.n8 a_n1140_n2688# 1.17037f
.ends

