* NGSPICE file created from diffpair353.ext - technology: sky130A

.subckt diffpair353 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t9 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X1 a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X2 source.t3 plus.t0 drain_left.t7 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X3 source.t2 plus.t1 drain_left.t6 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X5 source.t7 plus.t2 drain_left.t5 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X6 drain_left.t4 plus.t3 source.t6 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X7 drain_right.t6 minus.t1 source.t10 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X8 drain_right.t5 minus.t2 source.t14 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 source.t11 minus.t3 drain_right.t4 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X10 drain_right.t3 minus.t4 source.t15 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X11 drain_left.t3 plus.t4 source.t0 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X12 source.t5 plus.t5 drain_left.t2 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X13 drain_left.t1 plus.t6 source.t4 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X14 source.t12 minus.t5 drain_right.t2 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 source.t13 minus.t6 drain_right.t1 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X16 source.t8 minus.t7 drain_right.t0 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X17 a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X18 drain_left.t0 plus.t7 source.t1 a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X19 a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# a_n1346_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
R0 minus.n7 minus.t3 855.915
R1 minus.n2 minus.t4 855.915
R2 minus.n16 minus.t1 855.915
R3 minus.n11 minus.t7 855.915
R4 minus.n6 minus.t0 827.433
R5 minus.n1 minus.t5 827.433
R6 minus.n15 minus.t6 827.433
R7 minus.n10 minus.t2 827.433
R8 minus.n3 minus.n2 161.489
R9 minus.n12 minus.n11 161.489
R10 minus.n8 minus.n7 161.3
R11 minus.n5 minus.n0 161.3
R12 minus.n4 minus.n3 161.3
R13 minus.n17 minus.n16 161.3
R14 minus.n14 minus.n9 161.3
R15 minus.n13 minus.n12 161.3
R16 minus.n5 minus.n4 73.0308
R17 minus.n14 minus.n13 73.0308
R18 minus.n7 minus.n6 63.5369
R19 minus.n2 minus.n1 63.5369
R20 minus.n11 minus.n10 63.5369
R21 minus.n16 minus.n15 63.5369
R22 minus.n18 minus.n8 31.9096
R23 minus.n6 minus.n5 9.49444
R24 minus.n4 minus.n1 9.49444
R25 minus.n13 minus.n10 9.49444
R26 minus.n15 minus.n14 9.49444
R27 minus.n18 minus.n17 6.46262
R28 minus.n8 minus.n0 0.189894
R29 minus.n3 minus.n0 0.189894
R30 minus.n12 minus.n9 0.189894
R31 minus.n17 minus.n9 0.189894
R32 minus minus.n18 0.188
R33 source.n3 source.t3 51.0588
R34 source.n4 source.t15 51.0588
R35 source.n7 source.t11 51.0588
R36 source.n15 source.t10 51.0586
R37 source.n12 source.t8 51.0586
R38 source.n11 source.t0 51.0586
R39 source.n8 source.t7 51.0586
R40 source.n0 source.t1 51.0586
R41 source.n2 source.n1 48.8588
R42 source.n6 source.n5 48.8588
R43 source.n14 source.n13 48.8586
R44 source.n10 source.n9 48.8586
R45 source.n8 source.n7 19.5581
R46 source.n16 source.n0 14.0236
R47 source.n16 source.n15 5.53498
R48 source.n13 source.t14 2.2005
R49 source.n13 source.t13 2.2005
R50 source.n9 source.t4 2.2005
R51 source.n9 source.t2 2.2005
R52 source.n1 source.t6 2.2005
R53 source.n1 source.t5 2.2005
R54 source.n5 source.t9 2.2005
R55 source.n5 source.t12 2.2005
R56 source.n7 source.n6 0.543603
R57 source.n6 source.n4 0.543603
R58 source.n3 source.n2 0.543603
R59 source.n2 source.n0 0.543603
R60 source.n10 source.n8 0.543603
R61 source.n11 source.n10 0.543603
R62 source.n14 source.n12 0.543603
R63 source.n15 source.n14 0.543603
R64 source.n4 source.n3 0.470328
R65 source.n12 source.n11 0.470328
R66 source source.n16 0.188
R67 drain_right.n5 drain_right.n3 66.0805
R68 drain_right.n2 drain_right.n1 65.7535
R69 drain_right.n2 drain_right.n0 65.7535
R70 drain_right.n5 drain_right.n4 65.5376
R71 drain_right drain_right.n2 26.442
R72 drain_right drain_right.n5 6.19632
R73 drain_right.n1 drain_right.t1 2.2005
R74 drain_right.n1 drain_right.t6 2.2005
R75 drain_right.n0 drain_right.t0 2.2005
R76 drain_right.n0 drain_right.t5 2.2005
R77 drain_right.n3 drain_right.t2 2.2005
R78 drain_right.n3 drain_right.t3 2.2005
R79 drain_right.n4 drain_right.t4 2.2005
R80 drain_right.n4 drain_right.t7 2.2005
R81 plus.n2 plus.t0 855.915
R82 plus.n7 plus.t7 855.915
R83 plus.n11 plus.t4 855.915
R84 plus.n16 plus.t2 855.915
R85 plus.n1 plus.t3 827.433
R86 plus.n6 plus.t5 827.433
R87 plus.n10 plus.t1 827.433
R88 plus.n15 plus.t6 827.433
R89 plus.n3 plus.n2 161.489
R90 plus.n12 plus.n11 161.489
R91 plus.n4 plus.n3 161.3
R92 plus.n5 plus.n0 161.3
R93 plus.n8 plus.n7 161.3
R94 plus.n13 plus.n12 161.3
R95 plus.n14 plus.n9 161.3
R96 plus.n17 plus.n16 161.3
R97 plus.n5 plus.n4 73.0308
R98 plus.n14 plus.n13 73.0308
R99 plus.n2 plus.n1 63.5369
R100 plus.n7 plus.n6 63.5369
R101 plus.n16 plus.n15 63.5369
R102 plus.n11 plus.n10 63.5369
R103 plus plus.n17 26.9271
R104 plus plus.n8 10.9702
R105 plus.n4 plus.n1 9.49444
R106 plus.n6 plus.n5 9.49444
R107 plus.n15 plus.n14 9.49444
R108 plus.n13 plus.n10 9.49444
R109 plus.n3 plus.n0 0.189894
R110 plus.n8 plus.n0 0.189894
R111 plus.n17 plus.n9 0.189894
R112 plus.n12 plus.n9 0.189894
R113 drain_left.n5 drain_left.n3 66.0807
R114 drain_left.n2 drain_left.n1 65.7535
R115 drain_left.n2 drain_left.n0 65.7535
R116 drain_left.n5 drain_left.n4 65.5374
R117 drain_left drain_left.n2 26.9952
R118 drain_left drain_left.n5 6.19632
R119 drain_left.n1 drain_left.t6 2.2005
R120 drain_left.n1 drain_left.t3 2.2005
R121 drain_left.n0 drain_left.t5 2.2005
R122 drain_left.n0 drain_left.t1 2.2005
R123 drain_left.n4 drain_left.t2 2.2005
R124 drain_left.n4 drain_left.t0 2.2005
R125 drain_left.n3 drain_left.t7 2.2005
R126 drain_left.n3 drain_left.t4 2.2005
C0 source minus 2.29886f
C1 drain_left minus 0.170671f
C2 drain_right minus 2.6061f
C3 plus source 2.3129f
C4 plus drain_left 2.7333f
C5 drain_left source 12.8799f
C6 plus drain_right 0.280736f
C7 drain_right source 12.8791f
C8 drain_right drain_left 0.630082f
C9 plus minus 4.27661f
C10 drain_right a_n1346_n2688# 5.08925f
C11 drain_left a_n1346_n2688# 5.28602f
C12 source a_n1346_n2688# 6.888966f
C13 minus a_n1346_n2688# 4.984105f
C14 plus a_n1346_n2688# 6.75499f
C15 drain_left.t5 a_n1346_n2688# 0.232314f
C16 drain_left.t1 a_n1346_n2688# 0.232314f
C17 drain_left.n0 a_n1346_n2688# 2.03315f
C18 drain_left.t6 a_n1346_n2688# 0.232314f
C19 drain_left.t3 a_n1346_n2688# 0.232314f
C20 drain_left.n1 a_n1346_n2688# 2.03315f
C21 drain_left.n2 a_n1346_n2688# 1.92472f
C22 drain_left.t7 a_n1346_n2688# 0.232314f
C23 drain_left.t4 a_n1346_n2688# 0.232314f
C24 drain_left.n3 a_n1346_n2688# 2.03518f
C25 drain_left.t2 a_n1346_n2688# 0.232314f
C26 drain_left.t0 a_n1346_n2688# 0.232314f
C27 drain_left.n4 a_n1346_n2688# 2.03197f
C28 drain_left.n5 a_n1346_n2688# 1.0338f
C29 plus.n0 a_n1346_n2688# 0.056195f
C30 plus.t5 a_n1346_n2688# 0.429932f
C31 plus.t3 a_n1346_n2688# 0.429932f
C32 plus.n1 a_n1346_n2688# 0.179532f
C33 plus.t0 a_n1346_n2688# 0.435901f
C34 plus.n2 a_n1346_n2688# 0.19661f
C35 plus.n3 a_n1346_n2688# 0.118899f
C36 plus.n4 a_n1346_n2688# 0.020894f
C37 plus.n5 a_n1346_n2688# 0.020894f
C38 plus.n6 a_n1346_n2688# 0.179532f
C39 plus.t7 a_n1346_n2688# 0.435901f
C40 plus.n7 a_n1346_n2688# 0.196536f
C41 plus.n8 a_n1346_n2688# 0.5469f
C42 plus.n9 a_n1346_n2688# 0.056195f
C43 plus.t2 a_n1346_n2688# 0.435901f
C44 plus.t6 a_n1346_n2688# 0.429932f
C45 plus.t1 a_n1346_n2688# 0.429932f
C46 plus.n10 a_n1346_n2688# 0.179532f
C47 plus.t4 a_n1346_n2688# 0.435901f
C48 plus.n11 a_n1346_n2688# 0.19661f
C49 plus.n12 a_n1346_n2688# 0.118899f
C50 plus.n13 a_n1346_n2688# 0.020894f
C51 plus.n14 a_n1346_n2688# 0.020894f
C52 plus.n15 a_n1346_n2688# 0.179532f
C53 plus.n16 a_n1346_n2688# 0.196536f
C54 plus.n17 a_n1346_n2688# 1.41001f
C55 drain_right.t0 a_n1346_n2688# 0.232731f
C56 drain_right.t5 a_n1346_n2688# 0.232731f
C57 drain_right.n0 a_n1346_n2688# 2.0368f
C58 drain_right.t1 a_n1346_n2688# 0.232731f
C59 drain_right.t6 a_n1346_n2688# 0.232731f
C60 drain_right.n1 a_n1346_n2688# 2.0368f
C61 drain_right.n2 a_n1346_n2688# 1.86018f
C62 drain_right.t2 a_n1346_n2688# 0.232731f
C63 drain_right.t3 a_n1346_n2688# 0.232731f
C64 drain_right.n3 a_n1346_n2688# 2.03882f
C65 drain_right.t4 a_n1346_n2688# 0.232731f
C66 drain_right.t7 a_n1346_n2688# 0.232731f
C67 drain_right.n4 a_n1346_n2688# 2.03563f
C68 drain_right.n5 a_n1346_n2688# 1.03565f
C69 source.t1 a_n1346_n2688# 1.84336f
C70 source.n0 a_n1346_n2688# 1.05998f
C71 source.t6 a_n1346_n2688# 0.172867f
C72 source.t5 a_n1346_n2688# 0.172867f
C73 source.n1 a_n1346_n2688# 1.44713f
C74 source.n2 a_n1346_n2688# 0.311609f
C75 source.t3 a_n1346_n2688# 1.84337f
C76 source.n3 a_n1346_n2688# 0.38109f
C77 source.t15 a_n1346_n2688# 1.84337f
C78 source.n4 a_n1346_n2688# 0.38109f
C79 source.t9 a_n1346_n2688# 0.172867f
C80 source.t12 a_n1346_n2688# 0.172867f
C81 source.n5 a_n1346_n2688# 1.44713f
C82 source.n6 a_n1346_n2688# 0.311609f
C83 source.t11 a_n1346_n2688# 1.84337f
C84 source.n7 a_n1346_n2688# 1.41315f
C85 source.t7 a_n1346_n2688# 1.84336f
C86 source.n8 a_n1346_n2688# 1.41315f
C87 source.t4 a_n1346_n2688# 0.172867f
C88 source.t2 a_n1346_n2688# 0.172867f
C89 source.n9 a_n1346_n2688# 1.44713f
C90 source.n10 a_n1346_n2688# 0.311614f
C91 source.t0 a_n1346_n2688# 1.84336f
C92 source.n11 a_n1346_n2688# 0.381094f
C93 source.t8 a_n1346_n2688# 1.84336f
C94 source.n12 a_n1346_n2688# 0.381094f
C95 source.t14 a_n1346_n2688# 0.172867f
C96 source.t13 a_n1346_n2688# 0.172867f
C97 source.n13 a_n1346_n2688# 1.44713f
C98 source.n14 a_n1346_n2688# 0.311614f
C99 source.t10 a_n1346_n2688# 1.84336f
C100 source.n15 a_n1346_n2688# 0.518302f
C101 source.n16 a_n1346_n2688# 1.26531f
C102 minus.n0 a_n1346_n2688# 0.05492f
C103 minus.t3 a_n1346_n2688# 0.426008f
C104 minus.t0 a_n1346_n2688# 0.420175f
C105 minus.t5 a_n1346_n2688# 0.420175f
C106 minus.n1 a_n1346_n2688# 0.175458f
C107 minus.t4 a_n1346_n2688# 0.426008f
C108 minus.n2 a_n1346_n2688# 0.192148f
C109 minus.n3 a_n1346_n2688# 0.116201f
C110 minus.n4 a_n1346_n2688# 0.02042f
C111 minus.n5 a_n1346_n2688# 0.02042f
C112 minus.n6 a_n1346_n2688# 0.175458f
C113 minus.n7 a_n1346_n2688# 0.192076f
C114 minus.n8 a_n1346_n2688# 1.5831f
C115 minus.n9 a_n1346_n2688# 0.05492f
C116 minus.t6 a_n1346_n2688# 0.420175f
C117 minus.t2 a_n1346_n2688# 0.420175f
C118 minus.n10 a_n1346_n2688# 0.175458f
C119 minus.t7 a_n1346_n2688# 0.426008f
C120 minus.n11 a_n1346_n2688# 0.192148f
C121 minus.n12 a_n1346_n2688# 0.116201f
C122 minus.n13 a_n1346_n2688# 0.02042f
C123 minus.n14 a_n1346_n2688# 0.02042f
C124 minus.n15 a_n1346_n2688# 0.175458f
C125 minus.t1 a_n1346_n2688# 0.426008f
C126 minus.n16 a_n1346_n2688# 0.192076f
C127 minus.n17 a_n1346_n2688# 0.354205f
C128 minus.n18 a_n1346_n2688# 1.9477f
.ends

