* NGSPICE file created from diffpair577.ext - technology: sky130A

.subckt diffpair577 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t27 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t14 plus.t1 source.t26 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X3 drain_right.t15 minus.t0 source.t8 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 drain_right.t14 minus.t1 source.t7 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 source.t18 plus.t2 drain_left.t13 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X7 source.t29 plus.t3 drain_left.t12 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X8 drain_left.t11 plus.t4 source.t21 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X9 source.t30 minus.t2 drain_right.t13 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X10 source.t31 minus.t3 drain_right.t12 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 source.t2 minus.t4 drain_right.t11 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X12 source.t6 minus.t5 drain_right.t10 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X13 drain_right.t9 minus.t6 source.t1 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X14 drain_right.t8 minus.t7 source.t10 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X15 drain_left.t10 plus.t5 source.t23 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X16 source.t14 plus.t6 drain_left.t9 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X17 drain_right.t7 minus.t8 source.t12 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X18 a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X19 a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X20 drain_right.t6 minus.t9 source.t5 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 source.t9 minus.t10 drain_right.t5 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X22 drain_right.t4 minus.t11 source.t11 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X23 drain_right.t3 minus.t12 source.t4 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X24 source.t13 minus.t13 drain_right.t2 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X25 source.t25 plus.t7 drain_left.t8 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X26 drain_left.t7 plus.t8 source.t19 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X27 source.t28 plus.t9 drain_left.t6 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X28 source.t3 minus.t14 drain_right.t1 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X29 source.t0 minus.t15 drain_right.t0 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X30 source.t17 plus.t10 drain_left.t5 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X31 source.t20 plus.t11 drain_left.t4 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X32 drain_left.t3 plus.t12 source.t16 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X33 drain_left.t2 plus.t13 source.t22 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X34 source.t15 plus.t14 drain_left.t1 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X35 drain_left.t0 plus.t15 source.t24 a_n1670_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n4 plus.t6 2618.5
R1 plus.n17 plus.t13 2618.5
R2 plus.n23 plus.t0 2618.5
R3 plus.n36 plus.t9 2618.5
R4 plus.n3 plus.t4 2566.65
R5 plus.n7 plus.t14 2566.65
R6 plus.n9 plus.t8 2566.65
R7 plus.n1 plus.t7 2566.65
R8 plus.n14 plus.t5 2566.65
R9 plus.n16 plus.t3 2566.65
R10 plus.n22 plus.t2 2566.65
R11 plus.n26 plus.t1 2566.65
R12 plus.n28 plus.t10 2566.65
R13 plus.n20 plus.t15 2566.65
R14 plus.n33 plus.t11 2566.65
R15 plus.n35 plus.t12 2566.65
R16 plus.n5 plus.n4 161.489
R17 plus.n24 plus.n23 161.489
R18 plus.n6 plus.n5 161.3
R19 plus.n8 plus.n2 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n0 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n25 plus.n24 161.3
R25 plus.n27 plus.n21 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n19 161.3
R29 plus.n37 plus.n36 161.3
R30 plus.n6 plus.n3 47.4702
R31 plus.n16 plus.n15 47.4702
R32 plus.n35 plus.n34 47.4702
R33 plus.n25 plus.n22 47.4702
R34 plus.n8 plus.n7 43.0884
R35 plus.n14 plus.n13 43.0884
R36 plus.n33 plus.n32 43.0884
R37 plus.n27 plus.n26 43.0884
R38 plus.n10 plus.n9 38.7066
R39 plus.n10 plus.n1 38.7066
R40 plus.n29 plus.n20 38.7066
R41 plus.n29 plus.n28 38.7066
R42 plus.n9 plus.n8 34.3247
R43 plus.n13 plus.n1 34.3247
R44 plus.n32 plus.n20 34.3247
R45 plus.n28 plus.n27 34.3247
R46 plus plus.n37 32.3248
R47 plus.n7 plus.n6 29.9429
R48 plus.n15 plus.n14 29.9429
R49 plus.n34 plus.n33 29.9429
R50 plus.n26 plus.n25 29.9429
R51 plus.n4 plus.n3 25.5611
R52 plus.n17 plus.n16 25.5611
R53 plus.n36 plus.n35 25.5611
R54 plus.n23 plus.n22 25.5611
R55 plus plus.n18 15.1407
R56 plus.n5 plus.n2 0.189894
R57 plus.n11 plus.n2 0.189894
R58 plus.n12 plus.n11 0.189894
R59 plus.n12 plus.n0 0.189894
R60 plus.n18 plus.n0 0.189894
R61 plus.n37 plus.n19 0.189894
R62 plus.n31 plus.n19 0.189894
R63 plus.n31 plus.n30 0.189894
R64 plus.n30 plus.n21 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n0 source.t22 44.1297
R67 source.n7 source.t14 44.1296
R68 source.n8 source.t11 44.1296
R69 source.n15 source.t0 44.1296
R70 source.n31 source.t12 44.1295
R71 source.n24 source.t2 44.1295
R72 source.n23 source.t27 44.1295
R73 source.n16 source.t28 44.1295
R74 source.n2 source.n1 43.1397
R75 source.n4 source.n3 43.1397
R76 source.n6 source.n5 43.1397
R77 source.n10 source.n9 43.1397
R78 source.n12 source.n11 43.1397
R79 source.n14 source.n13 43.1397
R80 source.n30 source.n29 43.1396
R81 source.n28 source.n27 43.1396
R82 source.n26 source.n25 43.1396
R83 source.n22 source.n21 43.1396
R84 source.n20 source.n19 43.1396
R85 source.n18 source.n17 43.1396
R86 source.n16 source.n15 27.8052
R87 source.n32 source.n0 22.3138
R88 source.n32 source.n31 5.49188
R89 source.n29 source.t5 0.9905
R90 source.n29 source.t9 0.9905
R91 source.n27 source.t1 0.9905
R92 source.n27 source.t13 0.9905
R93 source.n25 source.t10 0.9905
R94 source.n25 source.t30 0.9905
R95 source.n21 source.t26 0.9905
R96 source.n21 source.t18 0.9905
R97 source.n19 source.t24 0.9905
R98 source.n19 source.t17 0.9905
R99 source.n17 source.t16 0.9905
R100 source.n17 source.t20 0.9905
R101 source.n1 source.t23 0.9905
R102 source.n1 source.t29 0.9905
R103 source.n3 source.t19 0.9905
R104 source.n3 source.t25 0.9905
R105 source.n5 source.t21 0.9905
R106 source.n5 source.t15 0.9905
R107 source.n9 source.t8 0.9905
R108 source.n9 source.t6 0.9905
R109 source.n11 source.t4 0.9905
R110 source.n11 source.t3 0.9905
R111 source.n13 source.t7 0.9905
R112 source.n13 source.t31 0.9905
R113 source.n8 source.n7 0.470328
R114 source.n24 source.n23 0.470328
R115 source.n15 source.n14 0.457397
R116 source.n14 source.n12 0.457397
R117 source.n12 source.n10 0.457397
R118 source.n10 source.n8 0.457397
R119 source.n7 source.n6 0.457397
R120 source.n6 source.n4 0.457397
R121 source.n4 source.n2 0.457397
R122 source.n2 source.n0 0.457397
R123 source.n18 source.n16 0.457397
R124 source.n20 source.n18 0.457397
R125 source.n22 source.n20 0.457397
R126 source.n23 source.n22 0.457397
R127 source.n26 source.n24 0.457397
R128 source.n28 source.n26 0.457397
R129 source.n30 source.n28 0.457397
R130 source.n31 source.n30 0.457397
R131 source source.n32 0.188
R132 drain_left.n9 drain_left.n7 60.2753
R133 drain_left.n5 drain_left.n3 60.2753
R134 drain_left.n2 drain_left.n0 60.2753
R135 drain_left.n13 drain_left.n12 59.8185
R136 drain_left.n11 drain_left.n10 59.8185
R137 drain_left.n9 drain_left.n8 59.8185
R138 drain_left.n5 drain_left.n4 59.8184
R139 drain_left.n2 drain_left.n1 59.8184
R140 drain_left drain_left.n6 36.3975
R141 drain_left drain_left.n13 6.11011
R142 drain_left.n3 drain_left.t13 0.9905
R143 drain_left.n3 drain_left.t15 0.9905
R144 drain_left.n4 drain_left.t5 0.9905
R145 drain_left.n4 drain_left.t14 0.9905
R146 drain_left.n1 drain_left.t4 0.9905
R147 drain_left.n1 drain_left.t0 0.9905
R148 drain_left.n0 drain_left.t6 0.9905
R149 drain_left.n0 drain_left.t3 0.9905
R150 drain_left.n12 drain_left.t12 0.9905
R151 drain_left.n12 drain_left.t2 0.9905
R152 drain_left.n10 drain_left.t8 0.9905
R153 drain_left.n10 drain_left.t10 0.9905
R154 drain_left.n8 drain_left.t1 0.9905
R155 drain_left.n8 drain_left.t7 0.9905
R156 drain_left.n7 drain_left.t9 0.9905
R157 drain_left.n7 drain_left.t11 0.9905
R158 drain_left.n11 drain_left.n9 0.457397
R159 drain_left.n13 drain_left.n11 0.457397
R160 drain_left.n6 drain_left.n5 0.173602
R161 drain_left.n6 drain_left.n2 0.173602
R162 minus.n17 minus.t15 2618.5
R163 minus.n4 minus.t11 2618.5
R164 minus.n36 minus.t8 2618.5
R165 minus.n23 minus.t4 2618.5
R166 minus.n16 minus.t1 2566.65
R167 minus.n14 minus.t3 2566.65
R168 minus.n1 minus.t12 2566.65
R169 minus.n9 minus.t14 2566.65
R170 minus.n7 minus.t0 2566.65
R171 minus.n3 minus.t5 2566.65
R172 minus.n35 minus.t10 2566.65
R173 minus.n33 minus.t9 2566.65
R174 minus.n20 minus.t13 2566.65
R175 minus.n28 minus.t6 2566.65
R176 minus.n26 minus.t2 2566.65
R177 minus.n22 minus.t7 2566.65
R178 minus.n5 minus.n4 161.489
R179 minus.n24 minus.n23 161.489
R180 minus.n18 minus.n17 161.3
R181 minus.n15 minus.n0 161.3
R182 minus.n13 minus.n12 161.3
R183 minus.n11 minus.n10 161.3
R184 minus.n8 minus.n2 161.3
R185 minus.n6 minus.n5 161.3
R186 minus.n37 minus.n36 161.3
R187 minus.n34 minus.n19 161.3
R188 minus.n32 minus.n31 161.3
R189 minus.n30 minus.n29 161.3
R190 minus.n27 minus.n21 161.3
R191 minus.n25 minus.n24 161.3
R192 minus.n16 minus.n15 47.4702
R193 minus.n6 minus.n3 47.4702
R194 minus.n25 minus.n22 47.4702
R195 minus.n35 minus.n34 47.4702
R196 minus.n14 minus.n13 43.0884
R197 minus.n8 minus.n7 43.0884
R198 minus.n27 minus.n26 43.0884
R199 minus.n33 minus.n32 43.0884
R200 minus.n38 minus.n18 41.474
R201 minus.n10 minus.n1 38.7066
R202 minus.n10 minus.n9 38.7066
R203 minus.n29 minus.n28 38.7066
R204 minus.n29 minus.n20 38.7066
R205 minus.n13 minus.n1 34.3247
R206 minus.n9 minus.n8 34.3247
R207 minus.n28 minus.n27 34.3247
R208 minus.n32 minus.n20 34.3247
R209 minus.n15 minus.n14 29.9429
R210 minus.n7 minus.n6 29.9429
R211 minus.n26 minus.n25 29.9429
R212 minus.n34 minus.n33 29.9429
R213 minus.n17 minus.n16 25.5611
R214 minus.n4 minus.n3 25.5611
R215 minus.n23 minus.n22 25.5611
R216 minus.n36 minus.n35 25.5611
R217 minus.n38 minus.n37 6.46641
R218 minus.n18 minus.n0 0.189894
R219 minus.n12 minus.n0 0.189894
R220 minus.n12 minus.n11 0.189894
R221 minus.n11 minus.n2 0.189894
R222 minus.n5 minus.n2 0.189894
R223 minus.n24 minus.n21 0.189894
R224 minus.n30 minus.n21 0.189894
R225 minus.n31 minus.n30 0.189894
R226 minus.n31 minus.n19 0.189894
R227 minus.n37 minus.n19 0.189894
R228 minus minus.n38 0.188
R229 drain_right.n9 drain_right.n7 60.2753
R230 drain_right.n5 drain_right.n3 60.2753
R231 drain_right.n2 drain_right.n0 60.2753
R232 drain_right.n9 drain_right.n8 59.8185
R233 drain_right.n11 drain_right.n10 59.8185
R234 drain_right.n13 drain_right.n12 59.8185
R235 drain_right.n5 drain_right.n4 59.8184
R236 drain_right.n2 drain_right.n1 59.8184
R237 drain_right drain_right.n6 35.8443
R238 drain_right drain_right.n13 6.11011
R239 drain_right.n3 drain_right.t5 0.9905
R240 drain_right.n3 drain_right.t7 0.9905
R241 drain_right.n4 drain_right.t2 0.9905
R242 drain_right.n4 drain_right.t6 0.9905
R243 drain_right.n1 drain_right.t13 0.9905
R244 drain_right.n1 drain_right.t9 0.9905
R245 drain_right.n0 drain_right.t11 0.9905
R246 drain_right.n0 drain_right.t8 0.9905
R247 drain_right.n7 drain_right.t10 0.9905
R248 drain_right.n7 drain_right.t4 0.9905
R249 drain_right.n8 drain_right.t1 0.9905
R250 drain_right.n8 drain_right.t15 0.9905
R251 drain_right.n10 drain_right.t12 0.9905
R252 drain_right.n10 drain_right.t3 0.9905
R253 drain_right.n12 drain_right.t0 0.9905
R254 drain_right.n12 drain_right.t14 0.9905
R255 drain_right.n13 drain_right.n11 0.457397
R256 drain_right.n11 drain_right.n9 0.457397
R257 drain_right.n6 drain_right.n5 0.173602
R258 drain_right.n6 drain_right.n2 0.173602
C0 drain_right plus 0.314737f
C1 drain_left minus 0.170856f
C2 source minus 6.28667f
C3 drain_left plus 7.206201f
C4 source plus 6.30071f
C5 plus minus 6.71871f
C6 drain_right drain_left 0.846053f
C7 drain_right source 59.341503f
C8 drain_right minus 7.04523f
C9 source drain_left 59.341904f
C10 drain_right a_n1670_n4888# 8.644311f
C11 drain_left a_n1670_n4888# 8.9189f
C12 source a_n1670_n4888# 12.804441f
C13 minus a_n1670_n4888# 7.011878f
C14 plus a_n1670_n4888# 9.647321f
C15 drain_right.t11 a_n1670_n4888# 0.61714f
C16 drain_right.t8 a_n1670_n4888# 0.61714f
C17 drain_right.n0 a_n1670_n4888# 5.64552f
C18 drain_right.t13 a_n1670_n4888# 0.61714f
C19 drain_right.t9 a_n1670_n4888# 0.61714f
C20 drain_right.n1 a_n1670_n4888# 5.64203f
C21 drain_right.n2 a_n1670_n4888# 0.870732f
C22 drain_right.t5 a_n1670_n4888# 0.61714f
C23 drain_right.t7 a_n1670_n4888# 0.61714f
C24 drain_right.n3 a_n1670_n4888# 5.64552f
C25 drain_right.t2 a_n1670_n4888# 0.61714f
C26 drain_right.t6 a_n1670_n4888# 0.61714f
C27 drain_right.n4 a_n1670_n4888# 5.64203f
C28 drain_right.n5 a_n1670_n4888# 0.870732f
C29 drain_right.n6 a_n1670_n4888# 2.51664f
C30 drain_right.t10 a_n1670_n4888# 0.61714f
C31 drain_right.t4 a_n1670_n4888# 0.61714f
C32 drain_right.n7 a_n1670_n4888# 5.64551f
C33 drain_right.t1 a_n1670_n4888# 0.61714f
C34 drain_right.t15 a_n1670_n4888# 0.61714f
C35 drain_right.n8 a_n1670_n4888# 5.64202f
C36 drain_right.n9 a_n1670_n4888# 0.901226f
C37 drain_right.t12 a_n1670_n4888# 0.61714f
C38 drain_right.t3 a_n1670_n4888# 0.61714f
C39 drain_right.n10 a_n1670_n4888# 5.64202f
C40 drain_right.n11 a_n1670_n4888# 0.444493f
C41 drain_right.t0 a_n1670_n4888# 0.61714f
C42 drain_right.t14 a_n1670_n4888# 0.61714f
C43 drain_right.n12 a_n1670_n4888# 5.64202f
C44 drain_right.n13 a_n1670_n4888# 0.764065f
C45 minus.n0 a_n1670_n4888# 0.054208f
C46 minus.t15 a_n1670_n4888# 0.615344f
C47 minus.t1 a_n1670_n4888# 0.610705f
C48 minus.t3 a_n1670_n4888# 0.610705f
C49 minus.t12 a_n1670_n4888# 0.610705f
C50 minus.n1 a_n1670_n4888# 0.232433f
C51 minus.n2 a_n1670_n4888# 0.054208f
C52 minus.t14 a_n1670_n4888# 0.610705f
C53 minus.t0 a_n1670_n4888# 0.610705f
C54 minus.t5 a_n1670_n4888# 0.610705f
C55 minus.n3 a_n1670_n4888# 0.232433f
C56 minus.t11 a_n1670_n4888# 0.615344f
C57 minus.n4 a_n1670_n4888# 0.248697f
C58 minus.n5 a_n1670_n4888# 0.12204f
C59 minus.n6 a_n1670_n4888# 0.018985f
C60 minus.n7 a_n1670_n4888# 0.232433f
C61 minus.n8 a_n1670_n4888# 0.018985f
C62 minus.n9 a_n1670_n4888# 0.232433f
C63 minus.n10 a_n1670_n4888# 0.018985f
C64 minus.n11 a_n1670_n4888# 0.054208f
C65 minus.n12 a_n1670_n4888# 0.054208f
C66 minus.n13 a_n1670_n4888# 0.018985f
C67 minus.n14 a_n1670_n4888# 0.232433f
C68 minus.n15 a_n1670_n4888# 0.018985f
C69 minus.n16 a_n1670_n4888# 0.232433f
C70 minus.n17 a_n1670_n4888# 0.248617f
C71 minus.n18 a_n1670_n4888# 2.35522f
C72 minus.n19 a_n1670_n4888# 0.054208f
C73 minus.t10 a_n1670_n4888# 0.610705f
C74 minus.t9 a_n1670_n4888# 0.610705f
C75 minus.t13 a_n1670_n4888# 0.610705f
C76 minus.n20 a_n1670_n4888# 0.232433f
C77 minus.n21 a_n1670_n4888# 0.054208f
C78 minus.t6 a_n1670_n4888# 0.610705f
C79 minus.t2 a_n1670_n4888# 0.610705f
C80 minus.t7 a_n1670_n4888# 0.610705f
C81 minus.n22 a_n1670_n4888# 0.232433f
C82 minus.t4 a_n1670_n4888# 0.615344f
C83 minus.n23 a_n1670_n4888# 0.248697f
C84 minus.n24 a_n1670_n4888# 0.12204f
C85 minus.n25 a_n1670_n4888# 0.018985f
C86 minus.n26 a_n1670_n4888# 0.232433f
C87 minus.n27 a_n1670_n4888# 0.018985f
C88 minus.n28 a_n1670_n4888# 0.232433f
C89 minus.n29 a_n1670_n4888# 0.018985f
C90 minus.n30 a_n1670_n4888# 0.054208f
C91 minus.n31 a_n1670_n4888# 0.054208f
C92 minus.n32 a_n1670_n4888# 0.018985f
C93 minus.n33 a_n1670_n4888# 0.232433f
C94 minus.n34 a_n1670_n4888# 0.018985f
C95 minus.n35 a_n1670_n4888# 0.232433f
C96 minus.t8 a_n1670_n4888# 0.615344f
C97 minus.n36 a_n1670_n4888# 0.248617f
C98 minus.n37 a_n1670_n4888# 0.350102f
C99 minus.n38 a_n1670_n4888# 2.81783f
C100 drain_left.t6 a_n1670_n4888# 0.617579f
C101 drain_left.t3 a_n1670_n4888# 0.617579f
C102 drain_left.n0 a_n1670_n4888# 5.64953f
C103 drain_left.t4 a_n1670_n4888# 0.617579f
C104 drain_left.t0 a_n1670_n4888# 0.617579f
C105 drain_left.n1 a_n1670_n4888# 5.64604f
C106 drain_left.n2 a_n1670_n4888# 0.871351f
C107 drain_left.t13 a_n1670_n4888# 0.617579f
C108 drain_left.t15 a_n1670_n4888# 0.617579f
C109 drain_left.n3 a_n1670_n4888# 5.64953f
C110 drain_left.t5 a_n1670_n4888# 0.617579f
C111 drain_left.t14 a_n1670_n4888# 0.617579f
C112 drain_left.n4 a_n1670_n4888# 5.64604f
C113 drain_left.n5 a_n1670_n4888# 0.871351f
C114 drain_left.n6 a_n1670_n4888# 2.59997f
C115 drain_left.t9 a_n1670_n4888# 0.617579f
C116 drain_left.t11 a_n1670_n4888# 0.617579f
C117 drain_left.n7 a_n1670_n4888# 5.64953f
C118 drain_left.t1 a_n1670_n4888# 0.617579f
C119 drain_left.t7 a_n1670_n4888# 0.617579f
C120 drain_left.n8 a_n1670_n4888# 5.64604f
C121 drain_left.n9 a_n1670_n4888# 0.901866f
C122 drain_left.t8 a_n1670_n4888# 0.617579f
C123 drain_left.t10 a_n1670_n4888# 0.617579f
C124 drain_left.n10 a_n1670_n4888# 5.64604f
C125 drain_left.n11 a_n1670_n4888# 0.444809f
C126 drain_left.t12 a_n1670_n4888# 0.617579f
C127 drain_left.t2 a_n1670_n4888# 0.617579f
C128 drain_left.n12 a_n1670_n4888# 5.64604f
C129 drain_left.n13 a_n1670_n4888# 0.764608f
C130 source.t22 a_n1670_n4888# 5.74493f
C131 source.n0 a_n1670_n4888# 2.42958f
C132 source.t23 a_n1670_n4888# 0.50269f
C133 source.t29 a_n1670_n4888# 0.50269f
C134 source.n1 a_n1670_n4888# 4.49426f
C135 source.n2 a_n1670_n4888# 0.420262f
C136 source.t19 a_n1670_n4888# 0.50269f
C137 source.t25 a_n1670_n4888# 0.50269f
C138 source.n3 a_n1670_n4888# 4.49426f
C139 source.n4 a_n1670_n4888# 0.420262f
C140 source.t21 a_n1670_n4888# 0.50269f
C141 source.t15 a_n1670_n4888# 0.50269f
C142 source.n5 a_n1670_n4888# 4.49426f
C143 source.n6 a_n1670_n4888# 0.420262f
C144 source.t14 a_n1670_n4888# 5.74494f
C145 source.n7 a_n1670_n4888# 0.541879f
C146 source.t11 a_n1670_n4888# 5.74494f
C147 source.n8 a_n1670_n4888# 0.541879f
C148 source.t8 a_n1670_n4888# 0.50269f
C149 source.t6 a_n1670_n4888# 0.50269f
C150 source.n9 a_n1670_n4888# 4.49426f
C151 source.n10 a_n1670_n4888# 0.420262f
C152 source.t4 a_n1670_n4888# 0.50269f
C153 source.t3 a_n1670_n4888# 0.50269f
C154 source.n11 a_n1670_n4888# 4.49426f
C155 source.n12 a_n1670_n4888# 0.420262f
C156 source.t7 a_n1670_n4888# 0.50269f
C157 source.t31 a_n1670_n4888# 0.50269f
C158 source.n13 a_n1670_n4888# 4.49426f
C159 source.n14 a_n1670_n4888# 0.420262f
C160 source.t0 a_n1670_n4888# 5.74494f
C161 source.n15 a_n1670_n4888# 2.98949f
C162 source.t28 a_n1670_n4888# 5.74491f
C163 source.n16 a_n1670_n4888# 2.98952f
C164 source.t16 a_n1670_n4888# 0.50269f
C165 source.t20 a_n1670_n4888# 0.50269f
C166 source.n17 a_n1670_n4888# 4.49427f
C167 source.n18 a_n1670_n4888# 0.420253f
C168 source.t24 a_n1670_n4888# 0.50269f
C169 source.t17 a_n1670_n4888# 0.50269f
C170 source.n19 a_n1670_n4888# 4.49427f
C171 source.n20 a_n1670_n4888# 0.420253f
C172 source.t26 a_n1670_n4888# 0.50269f
C173 source.t18 a_n1670_n4888# 0.50269f
C174 source.n21 a_n1670_n4888# 4.49427f
C175 source.n22 a_n1670_n4888# 0.420253f
C176 source.t27 a_n1670_n4888# 5.74491f
C177 source.n23 a_n1670_n4888# 0.541911f
C178 source.t2 a_n1670_n4888# 5.74491f
C179 source.n24 a_n1670_n4888# 0.541911f
C180 source.t10 a_n1670_n4888# 0.50269f
C181 source.t30 a_n1670_n4888# 0.50269f
C182 source.n25 a_n1670_n4888# 4.49427f
C183 source.n26 a_n1670_n4888# 0.420253f
C184 source.t1 a_n1670_n4888# 0.50269f
C185 source.t13 a_n1670_n4888# 0.50269f
C186 source.n27 a_n1670_n4888# 4.49427f
C187 source.n28 a_n1670_n4888# 0.420253f
C188 source.t5 a_n1670_n4888# 0.50269f
C189 source.t9 a_n1670_n4888# 0.50269f
C190 source.n29 a_n1670_n4888# 4.49427f
C191 source.n30 a_n1670_n4888# 0.420253f
C192 source.t12 a_n1670_n4888# 5.74491f
C193 source.n31 a_n1670_n4888# 0.714376f
C194 source.n32 a_n1670_n4888# 2.85769f
C195 plus.n0 a_n1670_n4888# 0.055052f
C196 plus.t3 a_n1670_n4888# 0.620212f
C197 plus.t5 a_n1670_n4888# 0.620212f
C198 plus.t7 a_n1670_n4888# 0.620212f
C199 plus.n1 a_n1670_n4888# 0.236051f
C200 plus.n2 a_n1670_n4888# 0.055052f
C201 plus.t8 a_n1670_n4888# 0.620212f
C202 plus.t14 a_n1670_n4888# 0.620212f
C203 plus.t4 a_n1670_n4888# 0.620212f
C204 plus.n3 a_n1670_n4888# 0.236051f
C205 plus.t6 a_n1670_n4888# 0.624923f
C206 plus.n4 a_n1670_n4888# 0.252568f
C207 plus.n5 a_n1670_n4888# 0.123939f
C208 plus.n6 a_n1670_n4888# 0.019281f
C209 plus.n7 a_n1670_n4888# 0.236051f
C210 plus.n8 a_n1670_n4888# 0.019281f
C211 plus.n9 a_n1670_n4888# 0.236051f
C212 plus.n10 a_n1670_n4888# 0.019281f
C213 plus.n11 a_n1670_n4888# 0.055052f
C214 plus.n12 a_n1670_n4888# 0.055052f
C215 plus.n13 a_n1670_n4888# 0.019281f
C216 plus.n14 a_n1670_n4888# 0.236051f
C217 plus.n15 a_n1670_n4888# 0.019281f
C218 plus.n16 a_n1670_n4888# 0.236051f
C219 plus.t13 a_n1670_n4888# 0.624923f
C220 plus.n17 a_n1670_n4888# 0.252487f
C221 plus.n18 a_n1670_n4888# 0.831671f
C222 plus.n19 a_n1670_n4888# 0.055052f
C223 plus.t9 a_n1670_n4888# 0.624923f
C224 plus.t12 a_n1670_n4888# 0.620212f
C225 plus.t11 a_n1670_n4888# 0.620212f
C226 plus.t15 a_n1670_n4888# 0.620212f
C227 plus.n20 a_n1670_n4888# 0.236051f
C228 plus.n21 a_n1670_n4888# 0.055052f
C229 plus.t10 a_n1670_n4888# 0.620212f
C230 plus.t1 a_n1670_n4888# 0.620212f
C231 plus.t2 a_n1670_n4888# 0.620212f
C232 plus.n22 a_n1670_n4888# 0.236051f
C233 plus.t0 a_n1670_n4888# 0.624923f
C234 plus.n23 a_n1670_n4888# 0.252568f
C235 plus.n24 a_n1670_n4888# 0.123939f
C236 plus.n25 a_n1670_n4888# 0.019281f
C237 plus.n26 a_n1670_n4888# 0.236051f
C238 plus.n27 a_n1670_n4888# 0.019281f
C239 plus.n28 a_n1670_n4888# 0.236051f
C240 plus.n29 a_n1670_n4888# 0.019281f
C241 plus.n30 a_n1670_n4888# 0.055052f
C242 plus.n31 a_n1670_n4888# 0.055052f
C243 plus.n32 a_n1670_n4888# 0.019281f
C244 plus.n33 a_n1670_n4888# 0.236051f
C245 plus.n34 a_n1670_n4888# 0.019281f
C246 plus.n35 a_n1670_n4888# 0.236051f
C247 plus.n36 a_n1670_n4888# 0.252487f
C248 plus.n37 a_n1670_n4888# 1.88621f
.ends

