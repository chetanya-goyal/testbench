* NGSPICE file created from diffpair395.ext - technology: sky130A

.subckt diffpair395 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t15 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X1 drain_right.t10 minus.t1 source.t19 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X2 source.t23 plus.t0 drain_left.t11 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X3 source.t22 plus.t1 drain_left.t10 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X5 drain_right.t9 minus.t2 source.t10 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X7 drain_right.t8 minus.t3 source.t12 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X9 drain_left.t9 plus.t2 source.t5 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 drain_left.t8 plus.t3 source.t8 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 source.t20 minus.t4 drain_right.t7 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X12 source.t18 minus.t5 drain_right.t6 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X13 a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X14 drain_right.t5 minus.t6 source.t17 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X15 source.t14 minus.t7 drain_right.t4 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X16 source.t13 minus.t8 drain_right.t3 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X17 drain_left.t7 plus.t4 source.t4 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X18 drain_right.t2 minus.t9 source.t11 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 source.t16 minus.t10 drain_right.t1 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X20 drain_left.t6 plus.t5 source.t7 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X21 drain_left.t5 plus.t6 source.t9 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X22 source.t21 minus.t11 drain_right.t0 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X23 source.t3 plus.t7 drain_left.t4 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X24 source.t2 plus.t8 drain_left.t3 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X25 source.t0 plus.t9 drain_left.t2 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X26 drain_left.t1 plus.t10 source.t6 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X27 source.t1 plus.t11 drain_left.t0 a_n2298_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n4 minus.t6 341.625
R1 minus.n20 minus.t11 341.625
R2 minus.n3 minus.t4 320.229
R3 minus.n7 minus.t3 320.229
R4 minus.n8 minus.t8 320.229
R5 minus.n12 minus.t9 320.229
R6 minus.n14 minus.t7 320.229
R7 minus.n19 minus.t2 320.229
R8 minus.n23 minus.t5 320.229
R9 minus.n24 minus.t1 320.229
R10 minus.n28 minus.t10 320.229
R11 minus.n30 minus.t0 320.229
R12 minus.n15 minus.n14 161.3
R13 minus.n13 minus.n0 161.3
R14 minus.n12 minus.n11 161.3
R15 minus.n10 minus.n1 161.3
R16 minus.n6 minus.n5 161.3
R17 minus.n31 minus.n30 161.3
R18 minus.n29 minus.n16 161.3
R19 minus.n28 minus.n27 161.3
R20 minus.n26 minus.n17 161.3
R21 minus.n22 minus.n21 161.3
R22 minus.n9 minus.n8 80.6037
R23 minus.n7 minus.n2 80.6037
R24 minus.n25 minus.n24 80.6037
R25 minus.n23 minus.n18 80.6037
R26 minus.n8 minus.n7 48.2005
R27 minus.n24 minus.n23 48.2005
R28 minus.n5 minus.n4 44.853
R29 minus.n21 minus.n20 44.853
R30 minus.n7 minus.n6 41.6278
R31 minus.n8 minus.n1 41.6278
R32 minus.n23 minus.n22 41.6278
R33 minus.n24 minus.n17 41.6278
R34 minus.n32 minus.n15 35.7543
R35 minus.n14 minus.n13 25.5611
R36 minus.n30 minus.n29 25.5611
R37 minus.n13 minus.n12 22.6399
R38 minus.n29 minus.n28 22.6399
R39 minus.n4 minus.n3 20.5405
R40 minus.n20 minus.n19 20.5405
R41 minus.n32 minus.n31 6.70126
R42 minus.n6 minus.n3 6.57323
R43 minus.n12 minus.n1 6.57323
R44 minus.n22 minus.n19 6.57323
R45 minus.n28 minus.n17 6.57323
R46 minus.n9 minus.n2 0.380177
R47 minus.n25 minus.n18 0.380177
R48 minus.n10 minus.n9 0.285035
R49 minus.n5 minus.n2 0.285035
R50 minus.n21 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n27 minus.n26 0.189894
R56 minus.n27 minus.n16 0.189894
R57 minus.n31 minus.n16 0.189894
R58 minus minus.n32 0.188
R59 source.n5 source.t1 51.0588
R60 source.n6 source.t17 51.0588
R61 source.n11 source.t14 51.0588
R62 source.n23 source.t15 51.0586
R63 source.n18 source.t21 51.0586
R64 source.n17 source.t4 51.0586
R65 source.n12 source.t3 51.0586
R66 source.n0 source.t7 51.0586
R67 source.n2 source.n1 48.8588
R68 source.n4 source.n3 48.8588
R69 source.n8 source.n7 48.8588
R70 source.n10 source.n9 48.8588
R71 source.n22 source.n21 48.8586
R72 source.n20 source.n19 48.8586
R73 source.n16 source.n15 48.8586
R74 source.n14 source.n13 48.8586
R75 source.n12 source.n11 19.9891
R76 source.n24 source.n0 14.2391
R77 source.n24 source.n23 5.7505
R78 source.n21 source.t19 2.2005
R79 source.n21 source.t16 2.2005
R80 source.n19 source.t10 2.2005
R81 source.n19 source.t18 2.2005
R82 source.n15 source.t8 2.2005
R83 source.n15 source.t22 2.2005
R84 source.n13 source.t5 2.2005
R85 source.n13 source.t23 2.2005
R86 source.n1 source.t9 2.2005
R87 source.n1 source.t0 2.2005
R88 source.n3 source.t6 2.2005
R89 source.n3 source.t2 2.2005
R90 source.n7 source.t12 2.2005
R91 source.n7 source.t20 2.2005
R92 source.n9 source.t11 2.2005
R93 source.n9 source.t13 2.2005
R94 source.n11 source.n10 0.974638
R95 source.n10 source.n8 0.974638
R96 source.n8 source.n6 0.974638
R97 source.n5 source.n4 0.974638
R98 source.n4 source.n2 0.974638
R99 source.n2 source.n0 0.974638
R100 source.n14 source.n12 0.974638
R101 source.n16 source.n14 0.974638
R102 source.n17 source.n16 0.974638
R103 source.n20 source.n18 0.974638
R104 source.n22 source.n20 0.974638
R105 source.n23 source.n22 0.974638
R106 source.n6 source.n5 0.470328
R107 source.n18 source.n17 0.470328
R108 source source.n24 0.188
R109 drain_right.n6 drain_right.n4 66.5116
R110 drain_right.n3 drain_right.n2 66.4561
R111 drain_right.n3 drain_right.n0 66.4561
R112 drain_right.n6 drain_right.n5 65.5376
R113 drain_right.n8 drain_right.n7 65.5376
R114 drain_right.n3 drain_right.n1 65.5373
R115 drain_right drain_right.n3 29.4118
R116 drain_right drain_right.n8 6.62735
R117 drain_right.n1 drain_right.t6 2.2005
R118 drain_right.n1 drain_right.t10 2.2005
R119 drain_right.n2 drain_right.t1 2.2005
R120 drain_right.n2 drain_right.t11 2.2005
R121 drain_right.n0 drain_right.t0 2.2005
R122 drain_right.n0 drain_right.t9 2.2005
R123 drain_right.n4 drain_right.t7 2.2005
R124 drain_right.n4 drain_right.t5 2.2005
R125 drain_right.n5 drain_right.t3 2.2005
R126 drain_right.n5 drain_right.t8 2.2005
R127 drain_right.n7 drain_right.t4 2.2005
R128 drain_right.n7 drain_right.t2 2.2005
R129 drain_right.n8 drain_right.n6 0.974638
R130 plus.n4 plus.t11 341.625
R131 plus.n20 plus.t4 341.625
R132 plus.n14 plus.t5 320.229
R133 plus.n12 plus.t9 320.229
R134 plus.n2 plus.t6 320.229
R135 plus.n7 plus.t8 320.229
R136 plus.n5 plus.t10 320.229
R137 plus.n30 plus.t7 320.229
R138 plus.n28 plus.t2 320.229
R139 plus.n18 plus.t0 320.229
R140 plus.n23 plus.t3 320.229
R141 plus.n21 plus.t1 320.229
R142 plus.n6 plus.n3 161.3
R143 plus.n11 plus.n10 161.3
R144 plus.n12 plus.n1 161.3
R145 plus.n13 plus.n0 161.3
R146 plus.n15 plus.n14 161.3
R147 plus.n22 plus.n19 161.3
R148 plus.n27 plus.n26 161.3
R149 plus.n28 plus.n17 161.3
R150 plus.n29 plus.n16 161.3
R151 plus.n31 plus.n30 161.3
R152 plus.n8 plus.n7 80.6037
R153 plus.n9 plus.n2 80.6037
R154 plus.n24 plus.n23 80.6037
R155 plus.n25 plus.n18 80.6037
R156 plus.n7 plus.n2 48.2005
R157 plus.n23 plus.n18 48.2005
R158 plus.n4 plus.n3 44.853
R159 plus.n20 plus.n19 44.853
R160 plus.n11 plus.n2 41.6278
R161 plus.n7 plus.n6 41.6278
R162 plus.n27 plus.n18 41.6278
R163 plus.n23 plus.n22 41.6278
R164 plus plus.n31 30.7717
R165 plus.n14 plus.n13 25.5611
R166 plus.n30 plus.n29 25.5611
R167 plus.n13 plus.n12 22.6399
R168 plus.n29 plus.n28 22.6399
R169 plus.n5 plus.n4 20.5405
R170 plus.n21 plus.n20 20.5405
R171 plus plus.n15 11.2088
R172 plus.n12 plus.n11 6.57323
R173 plus.n6 plus.n5 6.57323
R174 plus.n28 plus.n27 6.57323
R175 plus.n22 plus.n21 6.57323
R176 plus.n9 plus.n8 0.380177
R177 plus.n25 plus.n24 0.380177
R178 plus.n8 plus.n3 0.285035
R179 plus.n10 plus.n9 0.285035
R180 plus.n26 plus.n25 0.285035
R181 plus.n24 plus.n19 0.285035
R182 plus.n10 plus.n1 0.189894
R183 plus.n1 plus.n0 0.189894
R184 plus.n15 plus.n0 0.189894
R185 plus.n31 plus.n16 0.189894
R186 plus.n17 plus.n16 0.189894
R187 plus.n26 plus.n17 0.189894
R188 drain_left.n6 drain_left.n4 66.5117
R189 drain_left.n3 drain_left.n2 66.4561
R190 drain_left.n3 drain_left.n0 66.4561
R191 drain_left.n6 drain_left.n5 65.5376
R192 drain_left.n8 drain_left.n7 65.5374
R193 drain_left.n3 drain_left.n1 65.5373
R194 drain_left drain_left.n3 29.965
R195 drain_left drain_left.n8 6.62735
R196 drain_left.n1 drain_left.t11 2.2005
R197 drain_left.n1 drain_left.t8 2.2005
R198 drain_left.n2 drain_left.t10 2.2005
R199 drain_left.n2 drain_left.t7 2.2005
R200 drain_left.n0 drain_left.t4 2.2005
R201 drain_left.n0 drain_left.t9 2.2005
R202 drain_left.n7 drain_left.t2 2.2005
R203 drain_left.n7 drain_left.t6 2.2005
R204 drain_left.n5 drain_left.t3 2.2005
R205 drain_left.n5 drain_left.t5 2.2005
R206 drain_left.n4 drain_left.t0 2.2005
R207 drain_left.n4 drain_left.t1 2.2005
R208 drain_left.n8 drain_left.n6 0.974638
C0 drain_left drain_right 1.16185f
C1 minus source 6.52572f
C2 minus plus 5.44999f
C3 source drain_left 11.6601f
C4 drain_left plus 6.68972f
C5 source drain_right 11.6627f
C6 drain_right plus 0.381869f
C7 minus drain_left 0.17224f
C8 source plus 6.53976f
C9 minus drain_right 6.46341f
C10 drain_right a_n2298_n2688# 5.75739f
C11 drain_left a_n2298_n2688# 6.08396f
C12 source a_n2298_n2688# 7.517985f
C13 minus a_n2298_n2688# 8.874605f
C14 plus a_n2298_n2688# 10.3799f
C15 drain_left.t4 a_n2298_n2688# 0.189475f
C16 drain_left.t9 a_n2298_n2688# 0.189475f
C17 drain_left.n0 a_n2298_n2688# 1.66263f
C18 drain_left.t11 a_n2298_n2688# 0.189475f
C19 drain_left.t8 a_n2298_n2688# 0.189475f
C20 drain_left.n1 a_n2298_n2688# 1.65728f
C21 drain_left.t10 a_n2298_n2688# 0.189475f
C22 drain_left.t7 a_n2298_n2688# 0.189475f
C23 drain_left.n2 a_n2298_n2688# 1.66263f
C24 drain_left.n3 a_n2298_n2688# 2.34229f
C25 drain_left.t0 a_n2298_n2688# 0.189475f
C26 drain_left.t1 a_n2298_n2688# 0.189475f
C27 drain_left.n4 a_n2298_n2688# 1.66301f
C28 drain_left.t3 a_n2298_n2688# 0.189475f
C29 drain_left.t5 a_n2298_n2688# 0.189475f
C30 drain_left.n5 a_n2298_n2688# 1.65728f
C31 drain_left.n6 a_n2298_n2688# 0.766289f
C32 drain_left.t2 a_n2298_n2688# 0.189475f
C33 drain_left.t6 a_n2298_n2688# 0.189475f
C34 drain_left.n7 a_n2298_n2688# 1.65727f
C35 drain_left.n8 a_n2298_n2688# 0.619544f
C36 plus.n0 a_n2298_n2688# 0.040533f
C37 plus.t5 a_n2298_n2688# 0.83695f
C38 plus.t9 a_n2298_n2688# 0.83695f
C39 plus.n1 a_n2298_n2688# 0.040533f
C40 plus.t6 a_n2298_n2688# 0.83695f
C41 plus.n2 a_n2298_n2688# 0.35926f
C42 plus.n3 a_n2298_n2688# 0.186078f
C43 plus.t8 a_n2298_n2688# 0.83695f
C44 plus.t10 a_n2298_n2688# 0.83695f
C45 plus.t11 a_n2298_n2688# 0.858882f
C46 plus.n4 a_n2298_n2688# 0.332275f
C47 plus.n5 a_n2298_n2688# 0.351096f
C48 plus.n6 a_n2298_n2688# 0.009198f
C49 plus.n7 a_n2298_n2688# 0.35926f
C50 plus.n8 a_n2298_n2688# 0.067513f
C51 plus.n9 a_n2298_n2688# 0.067513f
C52 plus.n10 a_n2298_n2688# 0.054086f
C53 plus.n11 a_n2298_n2688# 0.009198f
C54 plus.n12 a_n2298_n2688# 0.347938f
C55 plus.n13 a_n2298_n2688# 0.009198f
C56 plus.n14 a_n2298_n2688# 0.347314f
C57 plus.n15 a_n2298_n2688# 0.417827f
C58 plus.n16 a_n2298_n2688# 0.040533f
C59 plus.t7 a_n2298_n2688# 0.83695f
C60 plus.n17 a_n2298_n2688# 0.040533f
C61 plus.t2 a_n2298_n2688# 0.83695f
C62 plus.t0 a_n2298_n2688# 0.83695f
C63 plus.n18 a_n2298_n2688# 0.35926f
C64 plus.n19 a_n2298_n2688# 0.186078f
C65 plus.t3 a_n2298_n2688# 0.83695f
C66 plus.t4 a_n2298_n2688# 0.858882f
C67 plus.n20 a_n2298_n2688# 0.332275f
C68 plus.t1 a_n2298_n2688# 0.83695f
C69 plus.n21 a_n2298_n2688# 0.351096f
C70 plus.n22 a_n2298_n2688# 0.009198f
C71 plus.n23 a_n2298_n2688# 0.35926f
C72 plus.n24 a_n2298_n2688# 0.067513f
C73 plus.n25 a_n2298_n2688# 0.067513f
C74 plus.n26 a_n2298_n2688# 0.054086f
C75 plus.n27 a_n2298_n2688# 0.009198f
C76 plus.n28 a_n2298_n2688# 0.347938f
C77 plus.n29 a_n2298_n2688# 0.009198f
C78 plus.n30 a_n2298_n2688# 0.347314f
C79 plus.n31 a_n2298_n2688# 1.23647f
C80 drain_right.t0 a_n2298_n2688# 0.188483f
C81 drain_right.t9 a_n2298_n2688# 0.188483f
C82 drain_right.n0 a_n2298_n2688# 1.65393f
C83 drain_right.t6 a_n2298_n2688# 0.188483f
C84 drain_right.t10 a_n2298_n2688# 0.188483f
C85 drain_right.n1 a_n2298_n2688# 1.6486f
C86 drain_right.t1 a_n2298_n2688# 0.188483f
C87 drain_right.t11 a_n2298_n2688# 0.188483f
C88 drain_right.n2 a_n2298_n2688# 1.65393f
C89 drain_right.n3 a_n2298_n2688# 2.27587f
C90 drain_right.t7 a_n2298_n2688# 0.188483f
C91 drain_right.t5 a_n2298_n2688# 0.188483f
C92 drain_right.n4 a_n2298_n2688# 1.6543f
C93 drain_right.t3 a_n2298_n2688# 0.188483f
C94 drain_right.t8 a_n2298_n2688# 0.188483f
C95 drain_right.n5 a_n2298_n2688# 1.6486f
C96 drain_right.n6 a_n2298_n2688# 0.762285f
C97 drain_right.t4 a_n2298_n2688# 0.188483f
C98 drain_right.t2 a_n2298_n2688# 0.188483f
C99 drain_right.n7 a_n2298_n2688# 1.6486f
C100 drain_right.n8 a_n2298_n2688# 0.616294f
C101 source.t7 a_n2298_n2688# 1.68745f
C102 source.n0 a_n2298_n2688# 1.02199f
C103 source.t9 a_n2298_n2688# 0.158246f
C104 source.t0 a_n2298_n2688# 0.158246f
C105 source.n1 a_n2298_n2688# 1.32473f
C106 source.n2 a_n2298_n2688# 0.34706f
C107 source.t6 a_n2298_n2688# 0.158246f
C108 source.t2 a_n2298_n2688# 0.158246f
C109 source.n3 a_n2298_n2688# 1.32473f
C110 source.n4 a_n2298_n2688# 0.34706f
C111 source.t1 a_n2298_n2688# 1.68746f
C112 source.n5 a_n2298_n2688# 0.379761f
C113 source.t17 a_n2298_n2688# 1.68746f
C114 source.n6 a_n2298_n2688# 0.379761f
C115 source.t12 a_n2298_n2688# 0.158246f
C116 source.t20 a_n2298_n2688# 0.158246f
C117 source.n7 a_n2298_n2688# 1.32473f
C118 source.n8 a_n2298_n2688# 0.34706f
C119 source.t11 a_n2298_n2688# 0.158246f
C120 source.t13 a_n2298_n2688# 0.158246f
C121 source.n9 a_n2298_n2688# 1.32473f
C122 source.n10 a_n2298_n2688# 0.34706f
C123 source.t14 a_n2298_n2688# 1.68746f
C124 source.n11 a_n2298_n2688# 1.35543f
C125 source.t3 a_n2298_n2688# 1.68745f
C126 source.n12 a_n2298_n2688# 1.35544f
C127 source.t5 a_n2298_n2688# 0.158246f
C128 source.t23 a_n2298_n2688# 0.158246f
C129 source.n13 a_n2298_n2688# 1.32473f
C130 source.n14 a_n2298_n2688# 0.347064f
C131 source.t8 a_n2298_n2688# 0.158246f
C132 source.t22 a_n2298_n2688# 0.158246f
C133 source.n15 a_n2298_n2688# 1.32473f
C134 source.n16 a_n2298_n2688# 0.347064f
C135 source.t4 a_n2298_n2688# 1.68745f
C136 source.n17 a_n2298_n2688# 0.379765f
C137 source.t21 a_n2298_n2688# 1.68745f
C138 source.n18 a_n2298_n2688# 0.379765f
C139 source.t10 a_n2298_n2688# 0.158246f
C140 source.t18 a_n2298_n2688# 0.158246f
C141 source.n19 a_n2298_n2688# 1.32473f
C142 source.n20 a_n2298_n2688# 0.347064f
C143 source.t19 a_n2298_n2688# 0.158246f
C144 source.t16 a_n2298_n2688# 0.158246f
C145 source.n21 a_n2298_n2688# 1.32473f
C146 source.n22 a_n2298_n2688# 0.347064f
C147 source.t15 a_n2298_n2688# 1.68745f
C148 source.n23 a_n2298_n2688# 0.529722f
C149 source.n24 a_n2298_n2688# 1.17499f
C150 minus.n0 a_n2298_n2688# 0.039921f
C151 minus.n1 a_n2298_n2688# 0.009059f
C152 minus.t9 a_n2298_n2688# 0.824318f
C153 minus.n2 a_n2298_n2688# 0.066494f
C154 minus.t4 a_n2298_n2688# 0.824318f
C155 minus.n3 a_n2298_n2688# 0.345797f
C156 minus.t6 a_n2298_n2688# 0.845919f
C157 minus.n4 a_n2298_n2688# 0.32726f
C158 minus.n5 a_n2298_n2688# 0.183269f
C159 minus.n6 a_n2298_n2688# 0.009059f
C160 minus.t3 a_n2298_n2688# 0.824318f
C161 minus.n7 a_n2298_n2688# 0.353838f
C162 minus.t8 a_n2298_n2688# 0.824318f
C163 minus.n8 a_n2298_n2688# 0.353838f
C164 minus.n9 a_n2298_n2688# 0.066494f
C165 minus.n10 a_n2298_n2688# 0.05327f
C166 minus.n11 a_n2298_n2688# 0.039921f
C167 minus.n12 a_n2298_n2688# 0.342687f
C168 minus.n13 a_n2298_n2688# 0.009059f
C169 minus.t7 a_n2298_n2688# 0.824318f
C170 minus.n14 a_n2298_n2688# 0.342072f
C171 minus.n15 a_n2298_n2688# 1.39037f
C172 minus.n16 a_n2298_n2688# 0.039921f
C173 minus.n17 a_n2298_n2688# 0.009059f
C174 minus.n18 a_n2298_n2688# 0.066494f
C175 minus.t2 a_n2298_n2688# 0.824318f
C176 minus.n19 a_n2298_n2688# 0.345797f
C177 minus.t11 a_n2298_n2688# 0.845919f
C178 minus.n20 a_n2298_n2688# 0.32726f
C179 minus.n21 a_n2298_n2688# 0.183269f
C180 minus.n22 a_n2298_n2688# 0.009059f
C181 minus.t5 a_n2298_n2688# 0.824318f
C182 minus.n23 a_n2298_n2688# 0.353838f
C183 minus.t1 a_n2298_n2688# 0.824318f
C184 minus.n24 a_n2298_n2688# 0.353838f
C185 minus.n25 a_n2298_n2688# 0.066494f
C186 minus.n26 a_n2298_n2688# 0.05327f
C187 minus.n27 a_n2298_n2688# 0.039921f
C188 minus.t10 a_n2298_n2688# 0.824318f
C189 minus.n28 a_n2298_n2688# 0.342687f
C190 minus.n29 a_n2298_n2688# 0.009059f
C191 minus.t0 a_n2298_n2688# 0.824318f
C192 minus.n30 a_n2298_n2688# 0.342072f
C193 minus.n31 a_n2298_n2688# 0.279748f
C194 minus.n32 a_n2298_n2688# 1.68457f
.ends

