* NGSPICE file created from diffpair526.ext - technology: sky130A

.subckt diffpair526 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t26 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X1 a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X2 source.t3 plus.t0 drain_left.t13 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X3 drain_left.t12 plus.t1 source.t8 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X4 a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X5 source.t25 minus.t1 drain_right.t12 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X6 drain_left.t11 plus.t2 source.t4 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X7 source.t7 plus.t3 drain_left.t10 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X8 drain_left.t9 plus.t4 source.t9 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X9 drain_right.t11 minus.t2 source.t24 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X10 source.t19 minus.t3 drain_right.t10 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X11 drain_right.t9 minus.t4 source.t20 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X12 drain_right.t8 minus.t5 source.t27 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X13 source.t0 plus.t5 drain_left.t8 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X14 drain_right.t7 minus.t6 source.t14 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 drain_left.t7 plus.t6 source.t11 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X16 a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X17 a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X18 drain_left.t6 plus.t7 source.t1 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 drain_left.t5 plus.t8 source.t6 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X20 source.t16 minus.t7 drain_right.t6 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X21 source.t2 plus.t9 drain_left.t4 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X22 drain_right.t5 minus.t8 source.t18 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X23 source.t22 minus.t9 drain_right.t4 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X24 drain_right.t3 minus.t10 source.t15 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X25 source.t10 plus.t10 drain_left.t3 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X26 source.t17 minus.t11 drain_right.t2 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X27 drain_right.t1 minus.t12 source.t23 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X28 source.t21 minus.t13 drain_right.t0 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X29 drain_left.t2 plus.t11 source.t13 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X30 drain_left.t1 plus.t12 source.t12 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X31 source.t5 plus.t13 drain_left.t0 a_n2044_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
R0 minus.n4 minus.t8 822.548
R1 minus.n20 minus.t4 822.548
R2 minus.n3 minus.t1 801.567
R3 minus.n7 minus.t5 801.567
R4 minus.n8 minus.t11 801.567
R5 minus.n1 minus.t2 801.567
R6 minus.n13 minus.t7 801.567
R7 minus.n14 minus.t0 801.567
R8 minus.n19 minus.t3 801.567
R9 minus.n23 minus.t10 801.567
R10 minus.n24 minus.t9 801.567
R11 minus.n17 minus.t6 801.567
R12 minus.n29 minus.t13 801.567
R13 minus.n30 minus.t12 801.567
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n0 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n1 161.3
R18 minus.n7 minus.n2 161.3
R19 minus.n6 minus.n5 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n16 161.3
R22 minus.n28 minus.n27 161.3
R23 minus.n26 minus.n17 161.3
R24 minus.n23 minus.n18 161.3
R25 minus.n22 minus.n21 161.3
R26 minus.n9 minus.n8 80.6037
R27 minus.n25 minus.n24 80.6037
R28 minus.n5 minus.n4 70.4033
R29 minus.n21 minus.n20 70.4033
R30 minus.n8 minus.n7 48.2005
R31 minus.n8 minus.n1 48.2005
R32 minus.n14 minus.n13 48.2005
R33 minus.n24 minus.n23 48.2005
R34 minus.n24 minus.n17 48.2005
R35 minus.n30 minus.n29 48.2005
R36 minus.n32 minus.n15 39.2297
R37 minus.n7 minus.n6 24.8308
R38 minus.n12 minus.n1 24.8308
R39 minus.n23 minus.n22 24.8308
R40 minus.n28 minus.n17 24.8308
R41 minus.n6 minus.n3 23.3702
R42 minus.n13 minus.n12 23.3702
R43 minus.n22 minus.n19 23.3702
R44 minus.n29 minus.n28 23.3702
R45 minus.n4 minus.n3 20.9576
R46 minus.n20 minus.n19 20.9576
R47 minus.n32 minus.n31 6.5933
R48 minus.n10 minus.n9 0.285035
R49 minus.n9 minus.n2 0.285035
R50 minus.n25 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n5 minus.n2 0.189894
R56 minus.n21 minus.n18 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n16 0.189894
R59 minus.n31 minus.n16 0.189894
R60 minus minus.n32 0.188
R61 source.n7 source.t18 45.521
R62 source.n27 source.t23 45.5208
R63 source.n20 source.t8 45.5208
R64 source.n0 source.t6 45.5208
R65 source.n2 source.n1 44.201
R66 source.n4 source.n3 44.201
R67 source.n6 source.n5 44.201
R68 source.n9 source.n8 44.201
R69 source.n11 source.n10 44.201
R70 source.n13 source.n12 44.201
R71 source.n26 source.n25 44.2008
R72 source.n24 source.n23 44.2008
R73 source.n22 source.n21 44.2008
R74 source.n19 source.n18 44.2008
R75 source.n17 source.n16 44.2008
R76 source.n15 source.n14 44.2008
R77 source.n15 source.n13 24.9915
R78 source.n28 source.n0 18.6553
R79 source.n28 source.n27 5.62119
R80 source.n25 source.t14 1.3205
R81 source.n25 source.t21 1.3205
R82 source.n23 source.t15 1.3205
R83 source.n23 source.t22 1.3205
R84 source.n21 source.t20 1.3205
R85 source.n21 source.t19 1.3205
R86 source.n18 source.t1 1.3205
R87 source.n18 source.t3 1.3205
R88 source.n16 source.t9 1.3205
R89 source.n16 source.t7 1.3205
R90 source.n14 source.t11 1.3205
R91 source.n14 source.t2 1.3205
R92 source.n1 source.t13 1.3205
R93 source.n1 source.t5 1.3205
R94 source.n3 source.t12 1.3205
R95 source.n3 source.t0 1.3205
R96 source.n5 source.t4 1.3205
R97 source.n5 source.t10 1.3205
R98 source.n8 source.t27 1.3205
R99 source.n8 source.t25 1.3205
R100 source.n10 source.t24 1.3205
R101 source.n10 source.t17 1.3205
R102 source.n12 source.t26 1.3205
R103 source.n12 source.t16 1.3205
R104 source.n7 source.n6 0.828086
R105 source.n22 source.n20 0.828086
R106 source.n13 source.n11 0.716017
R107 source.n11 source.n9 0.716017
R108 source.n9 source.n7 0.716017
R109 source.n6 source.n4 0.716017
R110 source.n4 source.n2 0.716017
R111 source.n2 source.n0 0.716017
R112 source.n17 source.n15 0.716017
R113 source.n19 source.n17 0.716017
R114 source.n20 source.n19 0.716017
R115 source.n24 source.n22 0.716017
R116 source.n26 source.n24 0.716017
R117 source.n27 source.n26 0.716017
R118 source source.n28 0.188
R119 drain_right.n1 drain_right.t9 62.9151
R120 drain_right.n11 drain_right.t13 62.1998
R121 drain_right.n8 drain_right.n6 61.5952
R122 drain_right.n4 drain_right.n2 61.5951
R123 drain_right.n8 drain_right.n7 60.8798
R124 drain_right.n10 drain_right.n9 60.8798
R125 drain_right.n4 drain_right.n3 60.8796
R126 drain_right.n1 drain_right.n0 60.8796
R127 drain_right drain_right.n5 33.2008
R128 drain_right drain_right.n11 6.01097
R129 drain_right.n2 drain_right.t0 1.3205
R130 drain_right.n2 drain_right.t1 1.3205
R131 drain_right.n3 drain_right.t4 1.3205
R132 drain_right.n3 drain_right.t7 1.3205
R133 drain_right.n0 drain_right.t10 1.3205
R134 drain_right.n0 drain_right.t3 1.3205
R135 drain_right.n6 drain_right.t12 1.3205
R136 drain_right.n6 drain_right.t5 1.3205
R137 drain_right.n7 drain_right.t2 1.3205
R138 drain_right.n7 drain_right.t8 1.3205
R139 drain_right.n9 drain_right.t6 1.3205
R140 drain_right.n9 drain_right.t11 1.3205
R141 drain_right.n11 drain_right.n10 0.716017
R142 drain_right.n10 drain_right.n8 0.716017
R143 drain_right.n5 drain_right.n1 0.481792
R144 drain_right.n5 drain_right.n4 0.124033
R145 plus.n4 plus.t2 822.548
R146 plus.n20 plus.t1 822.548
R147 plus.n14 plus.t8 801.567
R148 plus.n13 plus.t13 801.567
R149 plus.n1 plus.t11 801.567
R150 plus.n8 plus.t5 801.567
R151 plus.n7 plus.t12 801.567
R152 plus.n3 plus.t10 801.567
R153 plus.n30 plus.t6 801.567
R154 plus.n29 plus.t9 801.567
R155 plus.n17 plus.t4 801.567
R156 plus.n24 plus.t3 801.567
R157 plus.n23 plus.t7 801.567
R158 plus.n19 plus.t0 801.567
R159 plus.n6 plus.n5 161.3
R160 plus.n7 plus.n2 161.3
R161 plus.n10 plus.n1 161.3
R162 plus.n12 plus.n11 161.3
R163 plus.n13 plus.n0 161.3
R164 plus.n15 plus.n14 161.3
R165 plus.n22 plus.n21 161.3
R166 plus.n23 plus.n18 161.3
R167 plus.n26 plus.n17 161.3
R168 plus.n28 plus.n27 161.3
R169 plus.n29 plus.n16 161.3
R170 plus.n31 plus.n30 161.3
R171 plus.n9 plus.n8 80.6037
R172 plus.n25 plus.n24 80.6037
R173 plus.n5 plus.n4 70.4033
R174 plus.n21 plus.n20 70.4033
R175 plus.n14 plus.n13 48.2005
R176 plus.n8 plus.n1 48.2005
R177 plus.n8 plus.n7 48.2005
R178 plus.n30 plus.n29 48.2005
R179 plus.n24 plus.n17 48.2005
R180 plus.n24 plus.n23 48.2005
R181 plus plus.n31 31.9744
R182 plus.n12 plus.n1 24.8308
R183 plus.n7 plus.n6 24.8308
R184 plus.n28 plus.n17 24.8308
R185 plus.n23 plus.n22 24.8308
R186 plus.n13 plus.n12 23.3702
R187 plus.n6 plus.n3 23.3702
R188 plus.n29 plus.n28 23.3702
R189 plus.n22 plus.n19 23.3702
R190 plus.n4 plus.n3 20.9576
R191 plus.n20 plus.n19 20.9576
R192 plus plus.n15 13.3736
R193 plus.n9 plus.n2 0.285035
R194 plus.n10 plus.n9 0.285035
R195 plus.n26 plus.n25 0.285035
R196 plus.n25 plus.n18 0.285035
R197 plus.n5 plus.n2 0.189894
R198 plus.n11 plus.n10 0.189894
R199 plus.n11 plus.n0 0.189894
R200 plus.n15 plus.n0 0.189894
R201 plus.n31 plus.n16 0.189894
R202 plus.n27 plus.n16 0.189894
R203 plus.n27 plus.n26 0.189894
R204 plus.n21 plus.n18 0.189894
R205 drain_left.n7 drain_left.t11 62.9153
R206 drain_left.n1 drain_left.t7 62.9151
R207 drain_left.n4 drain_left.n2 61.5951
R208 drain_left.n9 drain_left.n8 60.8798
R209 drain_left.n7 drain_left.n6 60.8798
R210 drain_left.n11 drain_left.n10 60.8796
R211 drain_left.n4 drain_left.n3 60.8796
R212 drain_left.n1 drain_left.n0 60.8796
R213 drain_left drain_left.n5 33.754
R214 drain_left drain_left.n11 6.36873
R215 drain_left.n2 drain_left.t13 1.3205
R216 drain_left.n2 drain_left.t12 1.3205
R217 drain_left.n3 drain_left.t10 1.3205
R218 drain_left.n3 drain_left.t6 1.3205
R219 drain_left.n0 drain_left.t4 1.3205
R220 drain_left.n0 drain_left.t9 1.3205
R221 drain_left.n10 drain_left.t0 1.3205
R222 drain_left.n10 drain_left.t5 1.3205
R223 drain_left.n8 drain_left.t8 1.3205
R224 drain_left.n8 drain_left.t2 1.3205
R225 drain_left.n6 drain_left.t3 1.3205
R226 drain_left.n6 drain_left.t1 1.3205
R227 drain_left.n9 drain_left.n7 0.716017
R228 drain_left.n11 drain_left.n9 0.716017
R229 drain_left.n5 drain_left.n1 0.481792
R230 drain_left.n5 drain_left.n4 0.124033
C0 drain_right drain_left 1.06037f
C1 drain_right minus 9.15322f
C2 drain_left minus 0.172393f
C3 drain_right source 26.6556f
C4 drain_left source 26.6661f
C5 source minus 8.864841f
C6 drain_right plus 0.357905f
C7 drain_left plus 9.34989f
C8 plus minus 6.25139f
C9 plus source 8.879589f
C10 drain_right a_n2044_n3888# 8.232901f
C11 drain_left a_n2044_n3888# 8.537509f
C12 source a_n2044_n3888# 7.501649f
C13 minus a_n2044_n3888# 8.242093f
C14 plus a_n2044_n3888# 10.26408f
C15 drain_left.t7 a_n2044_n3888# 3.67724f
C16 drain_left.t4 a_n2044_n3888# 0.318357f
C17 drain_left.t9 a_n2044_n3888# 0.318357f
C18 drain_left.n0 a_n2044_n3888# 2.87758f
C19 drain_left.n1 a_n2044_n3888# 0.686152f
C20 drain_left.t13 a_n2044_n3888# 0.318357f
C21 drain_left.t12 a_n2044_n3888# 0.318357f
C22 drain_left.n2 a_n2044_n3888# 2.8817f
C23 drain_left.t10 a_n2044_n3888# 0.318357f
C24 drain_left.t6 a_n2044_n3888# 0.318357f
C25 drain_left.n3 a_n2044_n3888# 2.87758f
C26 drain_left.n4 a_n2044_n3888# 0.648158f
C27 drain_left.n5 a_n2044_n3888# 1.57275f
C28 drain_left.t11 a_n2044_n3888# 3.67724f
C29 drain_left.t3 a_n2044_n3888# 0.318357f
C30 drain_left.t1 a_n2044_n3888# 0.318357f
C31 drain_left.n6 a_n2044_n3888# 2.87758f
C32 drain_left.n7 a_n2044_n3888# 0.705124f
C33 drain_left.t8 a_n2044_n3888# 0.318357f
C34 drain_left.t2 a_n2044_n3888# 0.318357f
C35 drain_left.n8 a_n2044_n3888# 2.87758f
C36 drain_left.n9 a_n2044_n3888# 0.343823f
C37 drain_left.t0 a_n2044_n3888# 0.318357f
C38 drain_left.t5 a_n2044_n3888# 0.318357f
C39 drain_left.n10 a_n2044_n3888# 2.87757f
C40 drain_left.n11 a_n2044_n3888# 0.574579f
C41 plus.n0 a_n2044_n3888# 0.046313f
C42 plus.t8 a_n2044_n3888# 0.987051f
C43 plus.t13 a_n2044_n3888# 0.987051f
C44 plus.t11 a_n2044_n3888# 0.987051f
C45 plus.n1 a_n2044_n3888# 0.389374f
C46 plus.n2 a_n2044_n3888# 0.061798f
C47 plus.t5 a_n2044_n3888# 0.987051f
C48 plus.t12 a_n2044_n3888# 0.987051f
C49 plus.t10 a_n2044_n3888# 0.987051f
C50 plus.n3 a_n2044_n3888# 0.389089f
C51 plus.t2 a_n2044_n3888# 0.996862f
C52 plus.n4 a_n2044_n3888# 0.375066f
C53 plus.n5 a_n2044_n3888# 0.152288f
C54 plus.n6 a_n2044_n3888# 0.010509f
C55 plus.n7 a_n2044_n3888# 0.389374f
C56 plus.n8 a_n2044_n3888# 0.39503f
C57 plus.n9 a_n2044_n3888# 0.061654f
C58 plus.n10 a_n2044_n3888# 0.061798f
C59 plus.n11 a_n2044_n3888# 0.046313f
C60 plus.n12 a_n2044_n3888# 0.010509f
C61 plus.n13 a_n2044_n3888# 0.389089f
C62 plus.n14 a_n2044_n3888# 0.38452f
C63 plus.n15 a_n2044_n3888# 0.595404f
C64 plus.n16 a_n2044_n3888# 0.046313f
C65 plus.t6 a_n2044_n3888# 0.987051f
C66 plus.t9 a_n2044_n3888# 0.987051f
C67 plus.t4 a_n2044_n3888# 0.987051f
C68 plus.n17 a_n2044_n3888# 0.389374f
C69 plus.n18 a_n2044_n3888# 0.061798f
C70 plus.t3 a_n2044_n3888# 0.987051f
C71 plus.t7 a_n2044_n3888# 0.987051f
C72 plus.t0 a_n2044_n3888# 0.987051f
C73 plus.n19 a_n2044_n3888# 0.389089f
C74 plus.t1 a_n2044_n3888# 0.996862f
C75 plus.n20 a_n2044_n3888# 0.375066f
C76 plus.n21 a_n2044_n3888# 0.152288f
C77 plus.n22 a_n2044_n3888# 0.010509f
C78 plus.n23 a_n2044_n3888# 0.389374f
C79 plus.n24 a_n2044_n3888# 0.395029f
C80 plus.n25 a_n2044_n3888# 0.061654f
C81 plus.n26 a_n2044_n3888# 0.061798f
C82 plus.n27 a_n2044_n3888# 0.046313f
C83 plus.n28 a_n2044_n3888# 0.010509f
C84 plus.n29 a_n2044_n3888# 0.389089f
C85 plus.n30 a_n2044_n3888# 0.38452f
C86 plus.n31 a_n2044_n3888# 1.53171f
C87 drain_right.t9 a_n2044_n3888# 3.67776f
C88 drain_right.t10 a_n2044_n3888# 0.318402f
C89 drain_right.t3 a_n2044_n3888# 0.318402f
C90 drain_right.n0 a_n2044_n3888# 2.87798f
C91 drain_right.n1 a_n2044_n3888# 0.686249f
C92 drain_right.t0 a_n2044_n3888# 0.318402f
C93 drain_right.t1 a_n2044_n3888# 0.318402f
C94 drain_right.n2 a_n2044_n3888# 2.8821f
C95 drain_right.t4 a_n2044_n3888# 0.318402f
C96 drain_right.t7 a_n2044_n3888# 0.318402f
C97 drain_right.n3 a_n2044_n3888# 2.87798f
C98 drain_right.n4 a_n2044_n3888# 0.648249f
C99 drain_right.n5 a_n2044_n3888# 1.51725f
C100 drain_right.t12 a_n2044_n3888# 0.318402f
C101 drain_right.t5 a_n2044_n3888# 0.318402f
C102 drain_right.n6 a_n2044_n3888# 2.88209f
C103 drain_right.t2 a_n2044_n3888# 0.318402f
C104 drain_right.t8 a_n2044_n3888# 0.318402f
C105 drain_right.n7 a_n2044_n3888# 2.87798f
C106 drain_right.n8 a_n2044_n3888# 0.694452f
C107 drain_right.t6 a_n2044_n3888# 0.318402f
C108 drain_right.t11 a_n2044_n3888# 0.318402f
C109 drain_right.n9 a_n2044_n3888# 2.87798f
C110 drain_right.n10 a_n2044_n3888# 0.343872f
C111 drain_right.t13 a_n2044_n3888# 3.67361f
C112 drain_right.n11 a_n2044_n3888# 0.601047f
C113 source.t6 a_n2044_n3888# 3.68827f
C114 source.n0 a_n2044_n3888# 1.73321f
C115 source.t13 a_n2044_n3888# 0.329115f
C116 source.t5 a_n2044_n3888# 0.329115f
C117 source.n1 a_n2044_n3888# 2.891f
C118 source.n2 a_n2044_n3888# 0.401521f
C119 source.t12 a_n2044_n3888# 0.329115f
C120 source.t0 a_n2044_n3888# 0.329115f
C121 source.n3 a_n2044_n3888# 2.891f
C122 source.n4 a_n2044_n3888# 0.401521f
C123 source.t4 a_n2044_n3888# 0.329115f
C124 source.t10 a_n2044_n3888# 0.329115f
C125 source.n5 a_n2044_n3888# 2.891f
C126 source.n6 a_n2044_n3888# 0.411548f
C127 source.t18 a_n2044_n3888# 3.68827f
C128 source.n7 a_n2044_n3888# 0.511865f
C129 source.t27 a_n2044_n3888# 0.329115f
C130 source.t25 a_n2044_n3888# 0.329115f
C131 source.n8 a_n2044_n3888# 2.891f
C132 source.n9 a_n2044_n3888# 0.401521f
C133 source.t24 a_n2044_n3888# 0.329115f
C134 source.t17 a_n2044_n3888# 0.329115f
C135 source.n10 a_n2044_n3888# 2.891f
C136 source.n11 a_n2044_n3888# 0.401521f
C137 source.t26 a_n2044_n3888# 0.329115f
C138 source.t16 a_n2044_n3888# 0.329115f
C139 source.n12 a_n2044_n3888# 2.891f
C140 source.n13 a_n2044_n3888# 2.1645f
C141 source.t11 a_n2044_n3888# 0.329115f
C142 source.t2 a_n2044_n3888# 0.329115f
C143 source.n14 a_n2044_n3888# 2.891f
C144 source.n15 a_n2044_n3888# 2.16451f
C145 source.t9 a_n2044_n3888# 0.329115f
C146 source.t7 a_n2044_n3888# 0.329115f
C147 source.n16 a_n2044_n3888# 2.891f
C148 source.n17 a_n2044_n3888# 0.401525f
C149 source.t1 a_n2044_n3888# 0.329115f
C150 source.t3 a_n2044_n3888# 0.329115f
C151 source.n18 a_n2044_n3888# 2.891f
C152 source.n19 a_n2044_n3888# 0.401525f
C153 source.t8 a_n2044_n3888# 3.68827f
C154 source.n20 a_n2044_n3888# 0.51187f
C155 source.t20 a_n2044_n3888# 0.329115f
C156 source.t19 a_n2044_n3888# 0.329115f
C157 source.n21 a_n2044_n3888# 2.891f
C158 source.n22 a_n2044_n3888# 0.411552f
C159 source.t15 a_n2044_n3888# 0.329115f
C160 source.t22 a_n2044_n3888# 0.329115f
C161 source.n23 a_n2044_n3888# 2.891f
C162 source.n24 a_n2044_n3888# 0.401525f
C163 source.t14 a_n2044_n3888# 0.329115f
C164 source.t21 a_n2044_n3888# 0.329115f
C165 source.n25 a_n2044_n3888# 2.891f
C166 source.n26 a_n2044_n3888# 0.401525f
C167 source.t23 a_n2044_n3888# 3.68827f
C168 source.n27 a_n2044_n3888# 0.648856f
C169 source.n28 a_n2044_n3888# 2.03931f
C170 minus.n0 a_n2044_n3888# 0.045948f
C171 minus.t2 a_n2044_n3888# 0.979279f
C172 minus.n1 a_n2044_n3888# 0.386308f
C173 minus.n2 a_n2044_n3888# 0.061312f
C174 minus.t1 a_n2044_n3888# 0.979279f
C175 minus.n3 a_n2044_n3888# 0.386025f
C176 minus.t8 a_n2044_n3888# 0.989012f
C177 minus.n4 a_n2044_n3888# 0.372113f
C178 minus.n5 a_n2044_n3888# 0.151088f
C179 minus.n6 a_n2044_n3888# 0.010426f
C180 minus.t5 a_n2044_n3888# 0.979279f
C181 minus.n7 a_n2044_n3888# 0.386308f
C182 minus.t11 a_n2044_n3888# 0.979279f
C183 minus.n8 a_n2044_n3888# 0.391919f
C184 minus.n9 a_n2044_n3888# 0.061168f
C185 minus.n10 a_n2044_n3888# 0.061312f
C186 minus.n11 a_n2044_n3888# 0.045948f
C187 minus.n12 a_n2044_n3888# 0.010426f
C188 minus.t7 a_n2044_n3888# 0.979279f
C189 minus.n13 a_n2044_n3888# 0.386025f
C190 minus.t0 a_n2044_n3888# 0.979279f
C191 minus.n14 a_n2044_n3888# 0.381492f
C192 minus.n15 a_n2044_n3888# 1.84096f
C193 minus.n16 a_n2044_n3888# 0.045948f
C194 minus.t6 a_n2044_n3888# 0.979279f
C195 minus.n17 a_n2044_n3888# 0.386308f
C196 minus.n18 a_n2044_n3888# 0.061312f
C197 minus.t3 a_n2044_n3888# 0.979279f
C198 minus.n19 a_n2044_n3888# 0.386025f
C199 minus.t4 a_n2044_n3888# 0.989012f
C200 minus.n20 a_n2044_n3888# 0.372113f
C201 minus.n21 a_n2044_n3888# 0.151088f
C202 minus.n22 a_n2044_n3888# 0.010426f
C203 minus.t10 a_n2044_n3888# 0.979279f
C204 minus.n23 a_n2044_n3888# 0.386308f
C205 minus.t9 a_n2044_n3888# 0.979279f
C206 minus.n24 a_n2044_n3888# 0.391919f
C207 minus.n25 a_n2044_n3888# 0.061168f
C208 minus.n26 a_n2044_n3888# 0.061312f
C209 minus.n27 a_n2044_n3888# 0.045948f
C210 minus.n28 a_n2044_n3888# 0.010426f
C211 minus.t13 a_n2044_n3888# 0.979279f
C212 minus.n29 a_n2044_n3888# 0.386025f
C213 minus.t12 a_n2044_n3888# 0.979279f
C214 minus.n30 a_n2044_n3888# 0.381492f
C215 minus.n31 a_n2044_n3888# 0.310452f
C216 minus.n32 a_n2044_n3888# 2.21341f
.ends

