* NGSPICE file created from diffpair494.ext - technology: sky130A

.subckt diffpair494 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t14 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X1 a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X2 drain_left.t8 plus.t1 source.t13 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X3 drain_left.t7 plus.t2 source.t19 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X4 drain_right.t9 minus.t0 source.t4 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 source.t12 plus.t3 drain_left.t6 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 source.t16 plus.t4 drain_left.t5 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X7 drain_right.t8 minus.t1 source.t1 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 source.t7 minus.t2 drain_right.t7 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 drain_right.t6 minus.t3 source.t9 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X10 drain_left.t4 plus.t5 source.t10 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X11 source.t8 minus.t4 drain_right.t5 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X12 source.t2 minus.t5 drain_right.t4 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X13 drain_right.t3 minus.t6 source.t5 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X14 drain_right.t2 minus.t7 source.t6 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X15 drain_right.t1 minus.t8 source.t0 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X16 a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X17 drain_left.t3 plus.t6 source.t15 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X18 source.t17 plus.t7 drain_left.t2 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X19 a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X20 source.t3 minus.t9 drain_right.t0 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X21 a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X22 source.t11 plus.t8 drain_left.t1 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X23 drain_left.t0 plus.t9 source.t18 a_n1352_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n2 plus.t5 2009.43
R1 plus.n8 plus.t6 2009.43
R2 plus.n12 plus.t2 2009.43
R3 plus.n18 plus.t0 2009.43
R4 plus.n1 plus.t4 1964.15
R5 plus.n5 plus.t9 1964.15
R6 plus.n7 plus.t7 1964.15
R7 plus.n11 plus.t3 1964.15
R8 plus.n15 plus.t1 1964.15
R9 plus.n17 plus.t8 1964.15
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 40.8975
R19 plus.n7 plus.n6 40.8975
R20 plus.n17 plus.n16 40.8975
R21 plus.n14 plus.n11 40.8975
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus.n2 plus.n1 32.1338
R27 plus.n8 plus.n7 32.1338
R28 plus.n18 plus.n17 32.1338
R29 plus.n12 plus.n11 32.1338
R30 plus plus.n19 29.2092
R31 plus plus.n9 13.2297
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 source.n5 source.t5 45.521
R37 source.n19 source.t0 45.5208
R38 source.n14 source.t19 45.5208
R39 source.n0 source.t15 45.5208
R40 source.n2 source.n1 44.201
R41 source.n4 source.n3 44.201
R42 source.n7 source.n6 44.201
R43 source.n9 source.n8 44.201
R44 source.n18 source.n17 44.2008
R45 source.n16 source.n15 44.2008
R46 source.n13 source.n12 44.2008
R47 source.n11 source.n10 44.2008
R48 source.n11 source.n9 24.4742
R49 source.n20 source.n0 18.526
R50 source.n20 source.n19 5.49188
R51 source.n17 source.t1 1.3205
R52 source.n17 source.t8 1.3205
R53 source.n15 source.t9 1.3205
R54 source.n15 source.t2 1.3205
R55 source.n12 source.t13 1.3205
R56 source.n12 source.t12 1.3205
R57 source.n10 source.t14 1.3205
R58 source.n10 source.t11 1.3205
R59 source.n1 source.t18 1.3205
R60 source.n1 source.t17 1.3205
R61 source.n3 source.t10 1.3205
R62 source.n3 source.t16 1.3205
R63 source.n6 source.t4 1.3205
R64 source.n6 source.t7 1.3205
R65 source.n8 source.t6 1.3205
R66 source.n8 source.t3 1.3205
R67 source.n5 source.n4 0.698776
R68 source.n16 source.n14 0.698776
R69 source.n9 source.n7 0.457397
R70 source.n7 source.n5 0.457397
R71 source.n4 source.n2 0.457397
R72 source.n2 source.n0 0.457397
R73 source.n13 source.n11 0.457397
R74 source.n14 source.n13 0.457397
R75 source.n18 source.n16 0.457397
R76 source.n19 source.n18 0.457397
R77 source source.n20 0.188
R78 drain_left.n5 drain_left.t4 62.6567
R79 drain_left.n1 drain_left.t9 62.6565
R80 drain_left.n3 drain_left.n2 61.1669
R81 drain_left.n5 drain_left.n4 60.8798
R82 drain_left.n7 drain_left.n6 60.8796
R83 drain_left.n1 drain_left.n0 60.8796
R84 drain_left drain_left.n3 31.5816
R85 drain_left drain_left.n7 6.11011
R86 drain_left.n2 drain_left.t6 1.3205
R87 drain_left.n2 drain_left.t7 1.3205
R88 drain_left.n0 drain_left.t1 1.3205
R89 drain_left.n0 drain_left.t8 1.3205
R90 drain_left.n6 drain_left.t2 1.3205
R91 drain_left.n6 drain_left.t3 1.3205
R92 drain_left.n4 drain_left.t5 1.3205
R93 drain_left.n4 drain_left.t0 1.3205
R94 drain_left.n7 drain_left.n5 0.457397
R95 drain_left.n3 drain_left.n1 0.0593781
R96 minus.n8 minus.t7 2009.43
R97 minus.n2 minus.t6 2009.43
R98 minus.n18 minus.t8 2009.43
R99 minus.n12 minus.t3 2009.43
R100 minus.n7 minus.t9 1964.15
R101 minus.n5 minus.t0 1964.15
R102 minus.n1 minus.t2 1964.15
R103 minus.n17 minus.t4 1964.15
R104 minus.n15 minus.t1 1964.15
R105 minus.n11 minus.t5 1964.15
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 40.8975
R115 minus.n4 minus.n1 40.8975
R116 minus.n14 minus.n11 40.8975
R117 minus.n17 minus.n16 40.8975
R118 minus.n6 minus.n5 36.5157
R119 minus.n5 minus.n4 36.5157
R120 minus.n15 minus.n14 36.5157
R121 minus.n16 minus.n15 36.5157
R122 minus.n20 minus.n9 36.4645
R123 minus.n8 minus.n7 32.1338
R124 minus.n2 minus.n1 32.1338
R125 minus.n12 minus.n11 32.1338
R126 minus.n18 minus.n17 32.1338
R127 minus.n20 minus.n19 6.44936
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t6 62.6565
R134 drain_right.n7 drain_right.t2 62.1998
R135 drain_right.n6 drain_right.n4 61.3365
R136 drain_right.n3 drain_right.n2 61.1669
R137 drain_right.n6 drain_right.n5 60.8798
R138 drain_right.n1 drain_right.n0 60.8796
R139 drain_right drain_right.n3 31.0284
R140 drain_right drain_right.n7 5.88166
R141 drain_right.n2 drain_right.t5 1.3205
R142 drain_right.n2 drain_right.t1 1.3205
R143 drain_right.n0 drain_right.t4 1.3205
R144 drain_right.n0 drain_right.t8 1.3205
R145 drain_right.n4 drain_right.t7 1.3205
R146 drain_right.n4 drain_right.t3 1.3205
R147 drain_right.n5 drain_right.t0 1.3205
R148 drain_right.n5 drain_right.t9 1.3205
R149 drain_right.n7 drain_right.n6 0.457397
R150 drain_right.n3 drain_right.n1 0.0593781
C0 drain_left drain_right 0.664257f
C1 minus source 3.14907f
C2 plus minus 5.39611f
C3 plus source 3.16398f
C4 drain_left minus 0.170748f
C5 drain_right minus 3.74972f
C6 drain_left source 30.6323f
C7 drain_right source 30.6173f
C8 drain_left plus 3.87394f
C9 drain_right plus 0.284239f
C10 drain_right a_n1352_n3888# 8.02153f
C11 drain_left a_n1352_n3888# 8.24615f
C12 source a_n1352_n3888# 6.985667f
C13 minus a_n1352_n3888# 5.415092f
C14 plus a_n1352_n3888# 7.74949f
C15 drain_right.t6 a_n1352_n3888# 4.57506f
C16 drain_right.t4 a_n1352_n3888# 0.396264f
C17 drain_right.t8 a_n1352_n3888# 0.396264f
C18 drain_right.n0 a_n1352_n3888# 3.58176f
C19 drain_right.n1 a_n1352_n3888# 0.766457f
C20 drain_right.t5 a_n1352_n3888# 0.396264f
C21 drain_right.t1 a_n1352_n3888# 0.396264f
C22 drain_right.n2 a_n1352_n3888# 3.5835f
C23 drain_right.n3 a_n1352_n3888# 1.98616f
C24 drain_right.t7 a_n1352_n3888# 0.396264f
C25 drain_right.t3 a_n1352_n3888# 0.396264f
C26 drain_right.n4 a_n1352_n3888# 3.58463f
C27 drain_right.t0 a_n1352_n3888# 0.396264f
C28 drain_right.t9 a_n1352_n3888# 0.396264f
C29 drain_right.n5 a_n1352_n3888# 3.58177f
C30 drain_right.n6 a_n1352_n3888# 0.755094f
C31 drain_right.t2 a_n1352_n3888# 4.57195f
C32 drain_right.n7 a_n1352_n3888# 0.698745f
C33 minus.n0 a_n1352_n3888# 0.057123f
C34 minus.t7 a_n1352_n3888# 0.487785f
C35 minus.t9 a_n1352_n3888# 0.48346f
C36 minus.t0 a_n1352_n3888# 0.48346f
C37 minus.t2 a_n1352_n3888# 0.48346f
C38 minus.n1 a_n1352_n3888# 0.19157f
C39 minus.t6 a_n1352_n3888# 0.487785f
C40 minus.n2 a_n1352_n3888# 0.207684f
C41 minus.n3 a_n1352_n3888# 0.125436f
C42 minus.n4 a_n1352_n3888# 0.020006f
C43 minus.n5 a_n1352_n3888# 0.19157f
C44 minus.n6 a_n1352_n3888# 0.020006f
C45 minus.n7 a_n1352_n3888# 0.19157f
C46 minus.n8 a_n1352_n3888# 0.207604f
C47 minus.n9 a_n1352_n3888# 2.04021f
C48 minus.n10 a_n1352_n3888# 0.057123f
C49 minus.t4 a_n1352_n3888# 0.48346f
C50 minus.t1 a_n1352_n3888# 0.48346f
C51 minus.t5 a_n1352_n3888# 0.48346f
C52 minus.n11 a_n1352_n3888# 0.19157f
C53 minus.t3 a_n1352_n3888# 0.487785f
C54 minus.n12 a_n1352_n3888# 0.207684f
C55 minus.n13 a_n1352_n3888# 0.125436f
C56 minus.n14 a_n1352_n3888# 0.020006f
C57 minus.n15 a_n1352_n3888# 0.19157f
C58 minus.n16 a_n1352_n3888# 0.020006f
C59 minus.n17 a_n1352_n3888# 0.19157f
C60 minus.t8 a_n1352_n3888# 0.487785f
C61 minus.n18 a_n1352_n3888# 0.207604f
C62 minus.n19 a_n1352_n3888# 0.366626f
C63 minus.n20 a_n1352_n3888# 2.47861f
C64 drain_left.t9 a_n1352_n3888# 4.58426f
C65 drain_left.t1 a_n1352_n3888# 0.397061f
C66 drain_left.t8 a_n1352_n3888# 0.397061f
C67 drain_left.n0 a_n1352_n3888# 3.58897f
C68 drain_left.n1 a_n1352_n3888# 0.767998f
C69 drain_left.t6 a_n1352_n3888# 0.397061f
C70 drain_left.t7 a_n1352_n3888# 0.397061f
C71 drain_left.n2 a_n1352_n3888# 3.59071f
C72 drain_left.n3 a_n1352_n3888# 2.06048f
C73 drain_left.t4 a_n1352_n3888# 4.58426f
C74 drain_left.t5 a_n1352_n3888# 0.397061f
C75 drain_left.t0 a_n1352_n3888# 0.397061f
C76 drain_left.n4 a_n1352_n3888# 3.58897f
C77 drain_left.n5 a_n1352_n3888# 0.797763f
C78 drain_left.t2 a_n1352_n3888# 0.397061f
C79 drain_left.t3 a_n1352_n3888# 0.397061f
C80 drain_left.n6 a_n1352_n3888# 3.58896f
C81 drain_left.n7 a_n1352_n3888# 0.647151f
C82 source.t15 a_n1352_n3888# 4.53958f
C83 source.n0 a_n1352_n3888# 2.08733f
C84 source.t18 a_n1352_n3888# 0.405081f
C85 source.t17 a_n1352_n3888# 0.405081f
C86 source.n1 a_n1352_n3888# 3.55829f
C87 source.n2 a_n1352_n3888# 0.437242f
C88 source.t10 a_n1352_n3888# 0.405081f
C89 source.t16 a_n1352_n3888# 0.405081f
C90 source.n3 a_n1352_n3888# 3.55829f
C91 source.n4 a_n1352_n3888# 0.463822f
C92 source.t5 a_n1352_n3888# 4.53958f
C93 source.n5 a_n1352_n3888# 0.587294f
C94 source.t4 a_n1352_n3888# 0.405081f
C95 source.t7 a_n1352_n3888# 0.405081f
C96 source.n6 a_n1352_n3888# 3.55829f
C97 source.n7 a_n1352_n3888# 0.437242f
C98 source.t6 a_n1352_n3888# 0.405081f
C99 source.t3 a_n1352_n3888# 0.405081f
C100 source.n8 a_n1352_n3888# 3.55829f
C101 source.n9 a_n1352_n3888# 2.57867f
C102 source.t14 a_n1352_n3888# 0.405081f
C103 source.t11 a_n1352_n3888# 0.405081f
C104 source.n10 a_n1352_n3888# 3.55829f
C105 source.n11 a_n1352_n3888# 2.57867f
C106 source.t13 a_n1352_n3888# 0.405081f
C107 source.t12 a_n1352_n3888# 0.405081f
C108 source.n12 a_n1352_n3888# 3.55829f
C109 source.n13 a_n1352_n3888# 0.437247f
C110 source.t19 a_n1352_n3888# 4.53958f
C111 source.n14 a_n1352_n3888# 0.5873f
C112 source.t9 a_n1352_n3888# 0.405081f
C113 source.t2 a_n1352_n3888# 0.405081f
C114 source.n15 a_n1352_n3888# 3.55829f
C115 source.n16 a_n1352_n3888# 0.463827f
C116 source.t1 a_n1352_n3888# 0.405081f
C117 source.t8 a_n1352_n3888# 0.405081f
C118 source.n17 a_n1352_n3888# 3.55829f
C119 source.n18 a_n1352_n3888# 0.437247f
C120 source.t0 a_n1352_n3888# 4.53958f
C121 source.n19 a_n1352_n3888# 0.747446f
C122 source.n20 a_n1352_n3888# 2.4932f
C123 plus.n0 a_n1352_n3888# 0.059087f
C124 plus.t7 a_n1352_n3888# 0.500084f
C125 plus.t9 a_n1352_n3888# 0.500084f
C126 plus.t4 a_n1352_n3888# 0.500084f
C127 plus.n1 a_n1352_n3888# 0.198157f
C128 plus.t5 a_n1352_n3888# 0.504557f
C129 plus.n2 a_n1352_n3888# 0.214825f
C130 plus.n3 a_n1352_n3888# 0.12975f
C131 plus.n4 a_n1352_n3888# 0.020694f
C132 plus.n5 a_n1352_n3888# 0.198157f
C133 plus.n6 a_n1352_n3888# 0.020694f
C134 plus.n7 a_n1352_n3888# 0.198157f
C135 plus.t6 a_n1352_n3888# 0.504557f
C136 plus.n8 a_n1352_n3888# 0.214742f
C137 plus.n9 a_n1352_n3888# 0.739622f
C138 plus.n10 a_n1352_n3888# 0.059087f
C139 plus.t0 a_n1352_n3888# 0.504557f
C140 plus.t8 a_n1352_n3888# 0.500084f
C141 plus.t1 a_n1352_n3888# 0.500084f
C142 plus.t3 a_n1352_n3888# 0.500084f
C143 plus.n11 a_n1352_n3888# 0.198157f
C144 plus.t2 a_n1352_n3888# 0.504557f
C145 plus.n12 a_n1352_n3888# 0.214825f
C146 plus.n13 a_n1352_n3888# 0.12975f
C147 plus.n14 a_n1352_n3888# 0.020694f
C148 plus.n15 a_n1352_n3888# 0.198157f
C149 plus.n16 a_n1352_n3888# 0.020694f
C150 plus.n17 a_n1352_n3888# 0.198157f
C151 plus.n18 a_n1352_n3888# 0.214742f
C152 plus.n19 a_n1352_n3888# 1.72632f
.ends

