* NGSPICE file created from diffpair320.ext - technology: sky130A

.subckt diffpair320 minus drain_right drain_left source plus
X0 drain_right minus source a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=4.275 ps=18.95 w=9 l=0.15
X1 drain_left plus source a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=4.275 ps=18.95 w=9 l=0.15
X2 a_n976_n2692# a_n976_n2692# a_n976_n2692# a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X3 drain_right minus source a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=4.275 ps=18.95 w=9 l=0.15
X4 a_n976_n2692# a_n976_n2692# a_n976_n2692# a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X5 a_n976_n2692# a_n976_n2692# a_n976_n2692# a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X6 drain_left plus source a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=4.275 ps=18.95 w=9 l=0.15
X7 a_n976_n2692# a_n976_n2692# a_n976_n2692# a_n976_n2692# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
.ends

