* NGSPICE file created from diffpair57.ext - technology: sky130A

.subckt diffpair57 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t16 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X1 drain_left.t14 plus.t1 source.t23 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X2 source.t18 plus.t2 drain_left.t13 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X3 source.t17 plus.t3 drain_left.t12 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X4 drain_left.t11 plus.t4 source.t19 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 source.t15 minus.t0 drain_right.t15 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X6 drain_right.t14 minus.t1 source.t14 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X7 drain_right.t13 minus.t2 source.t7 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 drain_right.t12 minus.t3 source.t6 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X9 source.t13 minus.t4 drain_right.t11 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X10 a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X11 source.t10 minus.t5 drain_right.t10 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X12 source.t9 minus.t6 drain_right.t9 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 drain_right.t8 minus.t7 source.t8 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 source.t24 plus.t5 drain_left.t10 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 source.t28 plus.t6 drain_left.t9 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X16 source.t3 minus.t8 drain_right.t7 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X17 drain_right.t6 minus.t9 source.t5 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X18 drain_left.t8 plus.t7 source.t20 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X19 a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X20 drain_left.t7 plus.t8 source.t26 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 source.t4 minus.t10 drain_right.t5 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X22 drain_left.t6 plus.t9 source.t27 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X23 source.t21 plus.t10 drain_left.t5 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X24 drain_right.t4 minus.t11 source.t12 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X25 drain_left.t4 plus.t11 source.t25 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X26 source.t22 plus.t12 drain_left.t3 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X27 a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X28 source.t2 minus.t12 drain_right.t3 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X29 source.t31 plus.t13 drain_left.t2 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X30 drain_right.t2 minus.t13 source.t1 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X31 source.t30 plus.t14 drain_left.t1 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X32 drain_right.t1 minus.t14 source.t0 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X33 source.t11 minus.t15 drain_right.t0 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X34 a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X35 drain_left.t0 plus.t15 source.t29 a_n2390_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n8 plus.n7 161.3
R1 plus.n9 plus.n4 161.3
R2 plus.n11 plus.n10 161.3
R3 plus.n12 plus.n3 161.3
R4 plus.n14 plus.n13 161.3
R5 plus.n15 plus.n2 161.3
R6 plus.n17 plus.n16 161.3
R7 plus.n18 plus.n1 161.3
R8 plus.n20 plus.n19 161.3
R9 plus.n21 plus.n0 161.3
R10 plus.n23 plus.n22 161.3
R11 plus.n32 plus.n31 161.3
R12 plus.n33 plus.n28 161.3
R13 plus.n35 plus.n34 161.3
R14 plus.n36 plus.n27 161.3
R15 plus.n38 plus.n37 161.3
R16 plus.n39 plus.n26 161.3
R17 plus.n41 plus.n40 161.3
R18 plus.n42 plus.n25 161.3
R19 plus.n44 plus.n43 161.3
R20 plus.n45 plus.n24 161.3
R21 plus.n47 plus.n46 161.3
R22 plus.n6 plus.t12 126.621
R23 plus.n30 plus.t7 126.621
R24 plus.n22 plus.t1 105.638
R25 plus.n21 plus.t3 105.638
R26 plus.n1 plus.t4 105.638
R27 plus.n15 plus.t6 105.638
R28 plus.n3 plus.t8 105.638
R29 plus.n9 plus.t10 105.638
R30 plus.n5 plus.t11 105.638
R31 plus.n46 plus.t14 105.638
R32 plus.n45 plus.t0 105.638
R33 plus.n25 plus.t5 105.638
R34 plus.n39 plus.t9 105.638
R35 plus.n27 plus.t13 105.638
R36 plus.n33 plus.t15 105.638
R37 plus.n29 plus.t2 105.638
R38 plus.n7 plus.n6 70.4033
R39 plus.n31 plus.n30 70.4033
R40 plus.n22 plus.n21 48.2005
R41 plus.n46 plus.n45 48.2005
R42 plus.n20 plus.n1 44.549
R43 plus.n9 plus.n8 44.549
R44 plus.n44 plus.n25 44.549
R45 plus.n33 plus.n32 44.549
R46 plus.n16 plus.n15 34.3247
R47 plus.n10 plus.n3 34.3247
R48 plus.n40 plus.n39 34.3247
R49 plus.n34 plus.n27 34.3247
R50 plus plus.n47 28.0445
R51 plus.n14 plus.n3 24.1005
R52 plus.n15 plus.n14 24.1005
R53 plus.n39 plus.n38 24.1005
R54 plus.n38 plus.n27 24.1005
R55 plus.n6 plus.n5 20.9576
R56 plus.n30 plus.n29 20.9576
R57 plus.n16 plus.n1 13.8763
R58 plus.n10 plus.n9 13.8763
R59 plus.n40 plus.n25 13.8763
R60 plus.n34 plus.n33 13.8763
R61 plus plus.n23 8.13308
R62 plus.n21 plus.n20 3.65202
R63 plus.n8 plus.n5 3.65202
R64 plus.n45 plus.n44 3.65202
R65 plus.n32 plus.n29 3.65202
R66 plus.n7 plus.n4 0.189894
R67 plus.n11 plus.n4 0.189894
R68 plus.n12 plus.n11 0.189894
R69 plus.n13 plus.n12 0.189894
R70 plus.n13 plus.n2 0.189894
R71 plus.n17 plus.n2 0.189894
R72 plus.n18 plus.n17 0.189894
R73 plus.n19 plus.n18 0.189894
R74 plus.n19 plus.n0 0.189894
R75 plus.n23 plus.n0 0.189894
R76 plus.n47 plus.n24 0.189894
R77 plus.n43 plus.n24 0.189894
R78 plus.n43 plus.n42 0.189894
R79 plus.n42 plus.n41 0.189894
R80 plus.n41 plus.n26 0.189894
R81 plus.n37 plus.n26 0.189894
R82 plus.n37 plus.n36 0.189894
R83 plus.n36 plus.n35 0.189894
R84 plus.n35 plus.n28 0.189894
R85 plus.n31 plus.n28 0.189894
R86 source.n0 source.t23 243.255
R87 source.n7 source.t22 243.255
R88 source.n8 source.t12 243.255
R89 source.n15 source.t15 243.255
R90 source.n31 source.t6 243.254
R91 source.n24 source.t11 243.254
R92 source.n23 source.t20 243.254
R93 source.n16 source.t30 243.254
R94 source.n2 source.n1 223.454
R95 source.n4 source.n3 223.454
R96 source.n6 source.n5 223.454
R97 source.n10 source.n9 223.454
R98 source.n12 source.n11 223.454
R99 source.n14 source.n13 223.454
R100 source.n30 source.n29 223.453
R101 source.n28 source.n27 223.453
R102 source.n26 source.n25 223.453
R103 source.n22 source.n21 223.453
R104 source.n20 source.n19 223.453
R105 source.n18 source.n17 223.453
R106 source.n29 source.t1 19.8005
R107 source.n29 source.t9 19.8005
R108 source.n27 source.t0 19.8005
R109 source.n27 source.t2 19.8005
R110 source.n25 source.t8 19.8005
R111 source.n25 source.t10 19.8005
R112 source.n21 source.t29 19.8005
R113 source.n21 source.t18 19.8005
R114 source.n19 source.t27 19.8005
R115 source.n19 source.t31 19.8005
R116 source.n17 source.t16 19.8005
R117 source.n17 source.t24 19.8005
R118 source.n1 source.t19 19.8005
R119 source.n1 source.t17 19.8005
R120 source.n3 source.t26 19.8005
R121 source.n3 source.t28 19.8005
R122 source.n5 source.t25 19.8005
R123 source.n5 source.t21 19.8005
R124 source.n9 source.t5 19.8005
R125 source.n9 source.t4 19.8005
R126 source.n11 source.t14 19.8005
R127 source.n11 source.t3 19.8005
R128 source.n13 source.t7 19.8005
R129 source.n13 source.t13 19.8005
R130 source.n16 source.n15 13.7561
R131 source.n32 source.n0 8.09232
R132 source.n32 source.n31 5.66429
R133 source.n15 source.n14 0.802224
R134 source.n14 source.n12 0.802224
R135 source.n12 source.n10 0.802224
R136 source.n10 source.n8 0.802224
R137 source.n7 source.n6 0.802224
R138 source.n6 source.n4 0.802224
R139 source.n4 source.n2 0.802224
R140 source.n2 source.n0 0.802224
R141 source.n18 source.n16 0.802224
R142 source.n20 source.n18 0.802224
R143 source.n22 source.n20 0.802224
R144 source.n23 source.n22 0.802224
R145 source.n26 source.n24 0.802224
R146 source.n28 source.n26 0.802224
R147 source.n30 source.n28 0.802224
R148 source.n31 source.n30 0.802224
R149 source.n8 source.n7 0.470328
R150 source.n24 source.n23 0.470328
R151 source source.n32 0.188
R152 drain_left.n9 drain_left.n7 240.935
R153 drain_left.n5 drain_left.n3 240.934
R154 drain_left.n2 drain_left.n0 240.934
R155 drain_left.n13 drain_left.n12 240.132
R156 drain_left.n11 drain_left.n10 240.132
R157 drain_left.n9 drain_left.n8 240.132
R158 drain_left.n5 drain_left.n4 240.131
R159 drain_left.n2 drain_left.n1 240.131
R160 drain_left drain_left.n6 24.2449
R161 drain_left.n3 drain_left.t13 19.8005
R162 drain_left.n3 drain_left.t8 19.8005
R163 drain_left.n4 drain_left.t2 19.8005
R164 drain_left.n4 drain_left.t0 19.8005
R165 drain_left.n1 drain_left.t10 19.8005
R166 drain_left.n1 drain_left.t6 19.8005
R167 drain_left.n0 drain_left.t1 19.8005
R168 drain_left.n0 drain_left.t15 19.8005
R169 drain_left.n12 drain_left.t12 19.8005
R170 drain_left.n12 drain_left.t14 19.8005
R171 drain_left.n10 drain_left.t9 19.8005
R172 drain_left.n10 drain_left.t11 19.8005
R173 drain_left.n8 drain_left.t5 19.8005
R174 drain_left.n8 drain_left.t7 19.8005
R175 drain_left.n7 drain_left.t3 19.8005
R176 drain_left.n7 drain_left.t4 19.8005
R177 drain_left drain_left.n13 6.45494
R178 drain_left.n11 drain_left.n9 0.802224
R179 drain_left.n13 drain_left.n11 0.802224
R180 drain_left.n6 drain_left.n5 0.346016
R181 drain_left.n6 drain_left.n2 0.346016
R182 minus.n23 minus.n22 161.3
R183 minus.n21 minus.n0 161.3
R184 minus.n20 minus.n19 161.3
R185 minus.n18 minus.n1 161.3
R186 minus.n17 minus.n16 161.3
R187 minus.n15 minus.n2 161.3
R188 minus.n14 minus.n13 161.3
R189 minus.n12 minus.n3 161.3
R190 minus.n11 minus.n10 161.3
R191 minus.n9 minus.n4 161.3
R192 minus.n8 minus.n7 161.3
R193 minus.n47 minus.n46 161.3
R194 minus.n45 minus.n24 161.3
R195 minus.n44 minus.n43 161.3
R196 minus.n42 minus.n25 161.3
R197 minus.n41 minus.n40 161.3
R198 minus.n39 minus.n26 161.3
R199 minus.n38 minus.n37 161.3
R200 minus.n36 minus.n27 161.3
R201 minus.n35 minus.n34 161.3
R202 minus.n33 minus.n28 161.3
R203 minus.n32 minus.n31 161.3
R204 minus.n6 minus.t11 126.621
R205 minus.n30 minus.t15 126.621
R206 minus.n5 minus.t10 105.638
R207 minus.n9 minus.t9 105.638
R208 minus.n3 minus.t8 105.638
R209 minus.n15 minus.t1 105.638
R210 minus.n1 minus.t4 105.638
R211 minus.n21 minus.t2 105.638
R212 minus.n22 minus.t0 105.638
R213 minus.n29 minus.t7 105.638
R214 minus.n33 minus.t5 105.638
R215 minus.n27 minus.t14 105.638
R216 minus.n39 minus.t12 105.638
R217 minus.n25 minus.t13 105.638
R218 minus.n45 minus.t6 105.638
R219 minus.n46 minus.t3 105.638
R220 minus.n7 minus.n6 70.4033
R221 minus.n31 minus.n30 70.4033
R222 minus.n22 minus.n21 48.2005
R223 minus.n46 minus.n45 48.2005
R224 minus.n9 minus.n8 44.549
R225 minus.n20 minus.n1 44.549
R226 minus.n33 minus.n32 44.549
R227 minus.n44 minus.n25 44.549
R228 minus.n10 minus.n3 34.3247
R229 minus.n16 minus.n15 34.3247
R230 minus.n34 minus.n27 34.3247
R231 minus.n40 minus.n39 34.3247
R232 minus.n48 minus.n23 29.9967
R233 minus.n15 minus.n14 24.1005
R234 minus.n14 minus.n3 24.1005
R235 minus.n38 minus.n27 24.1005
R236 minus.n39 minus.n38 24.1005
R237 minus.n6 minus.n5 20.9576
R238 minus.n30 minus.n29 20.9576
R239 minus.n10 minus.n9 13.8763
R240 minus.n16 minus.n1 13.8763
R241 minus.n34 minus.n33 13.8763
R242 minus.n40 minus.n25 13.8763
R243 minus.n48 minus.n47 6.6558
R244 minus.n8 minus.n5 3.65202
R245 minus.n21 minus.n20 3.65202
R246 minus.n32 minus.n29 3.65202
R247 minus.n45 minus.n44 3.65202
R248 minus.n23 minus.n0 0.189894
R249 minus.n19 minus.n0 0.189894
R250 minus.n19 minus.n18 0.189894
R251 minus.n18 minus.n17 0.189894
R252 minus.n17 minus.n2 0.189894
R253 minus.n13 minus.n2 0.189894
R254 minus.n13 minus.n12 0.189894
R255 minus.n12 minus.n11 0.189894
R256 minus.n11 minus.n4 0.189894
R257 minus.n7 minus.n4 0.189894
R258 minus.n31 minus.n28 0.189894
R259 minus.n35 minus.n28 0.189894
R260 minus.n36 minus.n35 0.189894
R261 minus.n37 minus.n36 0.189894
R262 minus.n37 minus.n26 0.189894
R263 minus.n41 minus.n26 0.189894
R264 minus.n42 minus.n41 0.189894
R265 minus.n43 minus.n42 0.189894
R266 minus.n43 minus.n24 0.189894
R267 minus.n47 minus.n24 0.189894
R268 minus minus.n48 0.188
R269 drain_right.n9 drain_right.n7 240.935
R270 drain_right.n5 drain_right.n3 240.934
R271 drain_right.n2 drain_right.n0 240.934
R272 drain_right.n9 drain_right.n8 240.132
R273 drain_right.n11 drain_right.n10 240.132
R274 drain_right.n13 drain_right.n12 240.132
R275 drain_right.n5 drain_right.n4 240.131
R276 drain_right.n2 drain_right.n1 240.131
R277 drain_right drain_right.n6 23.6917
R278 drain_right.n3 drain_right.t9 19.8005
R279 drain_right.n3 drain_right.t12 19.8005
R280 drain_right.n4 drain_right.t3 19.8005
R281 drain_right.n4 drain_right.t2 19.8005
R282 drain_right.n1 drain_right.t10 19.8005
R283 drain_right.n1 drain_right.t1 19.8005
R284 drain_right.n0 drain_right.t0 19.8005
R285 drain_right.n0 drain_right.t8 19.8005
R286 drain_right.n7 drain_right.t5 19.8005
R287 drain_right.n7 drain_right.t4 19.8005
R288 drain_right.n8 drain_right.t7 19.8005
R289 drain_right.n8 drain_right.t6 19.8005
R290 drain_right.n10 drain_right.t11 19.8005
R291 drain_right.n10 drain_right.t14 19.8005
R292 drain_right.n12 drain_right.t15 19.8005
R293 drain_right.n12 drain_right.t13 19.8005
R294 drain_right drain_right.n13 6.45494
R295 drain_right.n13 drain_right.n11 0.802224
R296 drain_right.n11 drain_right.n9 0.802224
R297 drain_right.n6 drain_right.n5 0.346016
R298 drain_right.n6 drain_right.n2 0.346016
C0 drain_left source 4.79536f
C1 drain_left drain_right 1.24378f
C2 plus minus 4.09681f
C3 source drain_right 4.79706f
C4 drain_left minus 0.180003f
C5 drain_left plus 1.54076f
C6 source minus 1.89557f
C7 drain_right minus 1.30502f
C8 source plus 1.90944f
C9 drain_right plus 0.40055f
C10 drain_right a_n2390_n1088# 4.0997f
C11 drain_left a_n2390_n1088# 4.40217f
C12 source a_n2390_n1088# 2.686463f
C13 minus a_n2390_n1088# 8.561111f
C14 plus a_n2390_n1088# 9.172887f
C15 drain_right.t0 a_n2390_n1088# 0.016638f
C16 drain_right.t8 a_n2390_n1088# 0.016638f
C17 drain_right.n0 a_n2390_n1088# 0.06553f
C18 drain_right.t10 a_n2390_n1088# 0.016638f
C19 drain_right.t1 a_n2390_n1088# 0.016638f
C20 drain_right.n1 a_n2390_n1088# 0.06465f
C21 drain_right.n2 a_n2390_n1088# 0.490096f
C22 drain_right.t9 a_n2390_n1088# 0.016638f
C23 drain_right.t12 a_n2390_n1088# 0.016638f
C24 drain_right.n3 a_n2390_n1088# 0.06553f
C25 drain_right.t3 a_n2390_n1088# 0.016638f
C26 drain_right.t2 a_n2390_n1088# 0.016638f
C27 drain_right.n4 a_n2390_n1088# 0.06465f
C28 drain_right.n5 a_n2390_n1088# 0.490096f
C29 drain_right.n6 a_n2390_n1088# 0.652564f
C30 drain_right.t5 a_n2390_n1088# 0.016638f
C31 drain_right.t4 a_n2390_n1088# 0.016638f
C32 drain_right.n7 a_n2390_n1088# 0.06553f
C33 drain_right.t7 a_n2390_n1088# 0.016638f
C34 drain_right.t6 a_n2390_n1088# 0.016638f
C35 drain_right.n8 a_n2390_n1088# 0.06465f
C36 drain_right.n9 a_n2390_n1088# 0.519633f
C37 drain_right.t11 a_n2390_n1088# 0.016638f
C38 drain_right.t14 a_n2390_n1088# 0.016638f
C39 drain_right.n10 a_n2390_n1088# 0.06465f
C40 drain_right.n11 a_n2390_n1088# 0.256017f
C41 drain_right.t15 a_n2390_n1088# 0.016638f
C42 drain_right.t13 a_n2390_n1088# 0.016638f
C43 drain_right.n12 a_n2390_n1088# 0.06465f
C44 drain_right.n13 a_n2390_n1088# 0.439609f
C45 minus.n0 a_n2390_n1088# 0.0258f
C46 minus.t4 a_n2390_n1088# 0.052492f
C47 minus.n1 a_n2390_n1088# 0.054544f
C48 minus.n2 a_n2390_n1088# 0.0258f
C49 minus.t8 a_n2390_n1088# 0.052492f
C50 minus.n3 a_n2390_n1088# 0.054544f
C51 minus.n4 a_n2390_n1088# 0.0258f
C52 minus.t10 a_n2390_n1088# 0.052492f
C53 minus.n5 a_n2390_n1088# 0.053828f
C54 minus.t11 a_n2390_n1088# 0.061353f
C55 minus.n6 a_n2390_n1088# 0.044776f
C56 minus.n7 a_n2390_n1088# 0.086896f
C57 minus.n8 a_n2390_n1088# 0.005855f
C58 minus.t9 a_n2390_n1088# 0.052492f
C59 minus.n9 a_n2390_n1088# 0.054544f
C60 minus.n10 a_n2390_n1088# 0.005855f
C61 minus.n11 a_n2390_n1088# 0.0258f
C62 minus.n12 a_n2390_n1088# 0.0258f
C63 minus.n13 a_n2390_n1088# 0.0258f
C64 minus.n14 a_n2390_n1088# 0.005855f
C65 minus.t1 a_n2390_n1088# 0.052492f
C66 minus.n15 a_n2390_n1088# 0.054544f
C67 minus.n16 a_n2390_n1088# 0.005855f
C68 minus.n17 a_n2390_n1088# 0.0258f
C69 minus.n18 a_n2390_n1088# 0.0258f
C70 minus.n19 a_n2390_n1088# 0.0258f
C71 minus.n20 a_n2390_n1088# 0.005855f
C72 minus.t2 a_n2390_n1088# 0.052492f
C73 minus.n21 a_n2390_n1088# 0.053828f
C74 minus.t0 a_n2390_n1088# 0.052492f
C75 minus.n22 a_n2390_n1088# 0.05343f
C76 minus.n23 a_n2390_n1088# 0.67478f
C77 minus.n24 a_n2390_n1088# 0.0258f
C78 minus.t13 a_n2390_n1088# 0.052492f
C79 minus.n25 a_n2390_n1088# 0.054544f
C80 minus.n26 a_n2390_n1088# 0.0258f
C81 minus.t14 a_n2390_n1088# 0.052492f
C82 minus.n27 a_n2390_n1088# 0.054544f
C83 minus.n28 a_n2390_n1088# 0.0258f
C84 minus.t7 a_n2390_n1088# 0.052492f
C85 minus.n29 a_n2390_n1088# 0.053828f
C86 minus.t15 a_n2390_n1088# 0.061353f
C87 minus.n30 a_n2390_n1088# 0.044776f
C88 minus.n31 a_n2390_n1088# 0.086896f
C89 minus.n32 a_n2390_n1088# 0.005855f
C90 minus.t5 a_n2390_n1088# 0.052492f
C91 minus.n33 a_n2390_n1088# 0.054544f
C92 minus.n34 a_n2390_n1088# 0.005855f
C93 minus.n35 a_n2390_n1088# 0.0258f
C94 minus.n36 a_n2390_n1088# 0.0258f
C95 minus.n37 a_n2390_n1088# 0.0258f
C96 minus.n38 a_n2390_n1088# 0.005855f
C97 minus.t12 a_n2390_n1088# 0.052492f
C98 minus.n39 a_n2390_n1088# 0.054544f
C99 minus.n40 a_n2390_n1088# 0.005855f
C100 minus.n41 a_n2390_n1088# 0.0258f
C101 minus.n42 a_n2390_n1088# 0.0258f
C102 minus.n43 a_n2390_n1088# 0.0258f
C103 minus.n44 a_n2390_n1088# 0.005855f
C104 minus.t6 a_n2390_n1088# 0.052492f
C105 minus.n45 a_n2390_n1088# 0.053828f
C106 minus.t3 a_n2390_n1088# 0.052492f
C107 minus.n46 a_n2390_n1088# 0.05343f
C108 minus.n47 a_n2390_n1088# 0.178075f
C109 minus.n48 a_n2390_n1088# 0.827795f
C110 drain_left.t1 a_n2390_n1088# 0.016357f
C111 drain_left.t15 a_n2390_n1088# 0.016357f
C112 drain_left.n0 a_n2390_n1088# 0.064424f
C113 drain_left.t10 a_n2390_n1088# 0.016357f
C114 drain_left.t6 a_n2390_n1088# 0.016357f
C115 drain_left.n1 a_n2390_n1088# 0.063559f
C116 drain_left.n2 a_n2390_n1088# 0.481828f
C117 drain_left.t13 a_n2390_n1088# 0.016357f
C118 drain_left.t8 a_n2390_n1088# 0.016357f
C119 drain_left.n3 a_n2390_n1088# 0.064424f
C120 drain_left.t2 a_n2390_n1088# 0.016357f
C121 drain_left.t0 a_n2390_n1088# 0.016357f
C122 drain_left.n4 a_n2390_n1088# 0.063559f
C123 drain_left.n5 a_n2390_n1088# 0.481828f
C124 drain_left.n6 a_n2390_n1088# 0.681415f
C125 drain_left.t3 a_n2390_n1088# 0.016357f
C126 drain_left.t4 a_n2390_n1088# 0.016357f
C127 drain_left.n7 a_n2390_n1088# 0.064424f
C128 drain_left.t5 a_n2390_n1088# 0.016357f
C129 drain_left.t7 a_n2390_n1088# 0.016357f
C130 drain_left.n8 a_n2390_n1088# 0.063559f
C131 drain_left.n9 a_n2390_n1088# 0.510867f
C132 drain_left.t9 a_n2390_n1088# 0.016357f
C133 drain_left.t11 a_n2390_n1088# 0.016357f
C134 drain_left.n10 a_n2390_n1088# 0.063559f
C135 drain_left.n11 a_n2390_n1088# 0.251698f
C136 drain_left.t12 a_n2390_n1088# 0.016357f
C137 drain_left.t14 a_n2390_n1088# 0.016357f
C138 drain_left.n12 a_n2390_n1088# 0.063559f
C139 drain_left.n13 a_n2390_n1088# 0.432193f
C140 source.t23 a_n2390_n1088# 0.111263f
C141 source.n0 a_n2390_n1088# 0.515422f
C142 source.t19 a_n2390_n1088# 0.01999f
C143 source.t17 a_n2390_n1088# 0.01999f
C144 source.n1 a_n2390_n1088# 0.064831f
C145 source.n2 a_n2390_n1088# 0.286063f
C146 source.t26 a_n2390_n1088# 0.01999f
C147 source.t28 a_n2390_n1088# 0.01999f
C148 source.n3 a_n2390_n1088# 0.064831f
C149 source.n4 a_n2390_n1088# 0.286063f
C150 source.t25 a_n2390_n1088# 0.01999f
C151 source.t21 a_n2390_n1088# 0.01999f
C152 source.n5 a_n2390_n1088# 0.064831f
C153 source.n6 a_n2390_n1088# 0.286063f
C154 source.t22 a_n2390_n1088# 0.111263f
C155 source.n7 a_n2390_n1088# 0.267097f
C156 source.t12 a_n2390_n1088# 0.111263f
C157 source.n8 a_n2390_n1088# 0.267097f
C158 source.t5 a_n2390_n1088# 0.01999f
C159 source.t4 a_n2390_n1088# 0.01999f
C160 source.n9 a_n2390_n1088# 0.064831f
C161 source.n10 a_n2390_n1088# 0.286063f
C162 source.t14 a_n2390_n1088# 0.01999f
C163 source.t3 a_n2390_n1088# 0.01999f
C164 source.n11 a_n2390_n1088# 0.064831f
C165 source.n12 a_n2390_n1088# 0.286063f
C166 source.t7 a_n2390_n1088# 0.01999f
C167 source.t13 a_n2390_n1088# 0.01999f
C168 source.n13 a_n2390_n1088# 0.064831f
C169 source.n14 a_n2390_n1088# 0.286063f
C170 source.t15 a_n2390_n1088# 0.111263f
C171 source.n15 a_n2390_n1088# 0.722608f
C172 source.t30 a_n2390_n1088# 0.111262f
C173 source.n16 a_n2390_n1088# 0.722608f
C174 source.t16 a_n2390_n1088# 0.01999f
C175 source.t24 a_n2390_n1088# 0.01999f
C176 source.n17 a_n2390_n1088# 0.064831f
C177 source.n18 a_n2390_n1088# 0.286063f
C178 source.t27 a_n2390_n1088# 0.01999f
C179 source.t31 a_n2390_n1088# 0.01999f
C180 source.n19 a_n2390_n1088# 0.064831f
C181 source.n20 a_n2390_n1088# 0.286063f
C182 source.t29 a_n2390_n1088# 0.01999f
C183 source.t18 a_n2390_n1088# 0.01999f
C184 source.n21 a_n2390_n1088# 0.064831f
C185 source.n22 a_n2390_n1088# 0.286063f
C186 source.t20 a_n2390_n1088# 0.111262f
C187 source.n23 a_n2390_n1088# 0.267098f
C188 source.t11 a_n2390_n1088# 0.111262f
C189 source.n24 a_n2390_n1088# 0.267098f
C190 source.t8 a_n2390_n1088# 0.01999f
C191 source.t10 a_n2390_n1088# 0.01999f
C192 source.n25 a_n2390_n1088# 0.064831f
C193 source.n26 a_n2390_n1088# 0.286063f
C194 source.t0 a_n2390_n1088# 0.01999f
C195 source.t2 a_n2390_n1088# 0.01999f
C196 source.n27 a_n2390_n1088# 0.064831f
C197 source.n28 a_n2390_n1088# 0.286063f
C198 source.t1 a_n2390_n1088# 0.01999f
C199 source.t9 a_n2390_n1088# 0.01999f
C200 source.n29 a_n2390_n1088# 0.064831f
C201 source.n30 a_n2390_n1088# 0.286063f
C202 source.t6 a_n2390_n1088# 0.111262f
C203 source.n31 a_n2390_n1088# 0.426602f
C204 source.n32 a_n2390_n1088# 0.521184f
C205 plus.n0 a_n2390_n1088# 0.026132f
C206 plus.t1 a_n2390_n1088# 0.053169f
C207 plus.t3 a_n2390_n1088# 0.053169f
C208 plus.t4 a_n2390_n1088# 0.053169f
C209 plus.n1 a_n2390_n1088# 0.055247f
C210 plus.n2 a_n2390_n1088# 0.026132f
C211 plus.t6 a_n2390_n1088# 0.053169f
C212 plus.t8 a_n2390_n1088# 0.053169f
C213 plus.n3 a_n2390_n1088# 0.055247f
C214 plus.n4 a_n2390_n1088# 0.026132f
C215 plus.t10 a_n2390_n1088# 0.053169f
C216 plus.t11 a_n2390_n1088# 0.053169f
C217 plus.n5 a_n2390_n1088# 0.054522f
C218 plus.t12 a_n2390_n1088# 0.062144f
C219 plus.n6 a_n2390_n1088# 0.045353f
C220 plus.n7 a_n2390_n1088# 0.088017f
C221 plus.n8 a_n2390_n1088# 0.00593f
C222 plus.n9 a_n2390_n1088# 0.055247f
C223 plus.n10 a_n2390_n1088# 0.00593f
C224 plus.n11 a_n2390_n1088# 0.026132f
C225 plus.n12 a_n2390_n1088# 0.026132f
C226 plus.n13 a_n2390_n1088# 0.026132f
C227 plus.n14 a_n2390_n1088# 0.00593f
C228 plus.n15 a_n2390_n1088# 0.055247f
C229 plus.n16 a_n2390_n1088# 0.00593f
C230 plus.n17 a_n2390_n1088# 0.026132f
C231 plus.n18 a_n2390_n1088# 0.026132f
C232 plus.n19 a_n2390_n1088# 0.026132f
C233 plus.n20 a_n2390_n1088# 0.00593f
C234 plus.n21 a_n2390_n1088# 0.054522f
C235 plus.n22 a_n2390_n1088# 0.054119f
C236 plus.n23 a_n2390_n1088# 0.189205f
C237 plus.n24 a_n2390_n1088# 0.026132f
C238 plus.t14 a_n2390_n1088# 0.053169f
C239 plus.t0 a_n2390_n1088# 0.053169f
C240 plus.t5 a_n2390_n1088# 0.053169f
C241 plus.n25 a_n2390_n1088# 0.055247f
C242 plus.n26 a_n2390_n1088# 0.026132f
C243 plus.t9 a_n2390_n1088# 0.053169f
C244 plus.t13 a_n2390_n1088# 0.053169f
C245 plus.n27 a_n2390_n1088# 0.055247f
C246 plus.n28 a_n2390_n1088# 0.026132f
C247 plus.t15 a_n2390_n1088# 0.053169f
C248 plus.t2 a_n2390_n1088# 0.053169f
C249 plus.n29 a_n2390_n1088# 0.054522f
C250 plus.t7 a_n2390_n1088# 0.062144f
C251 plus.n30 a_n2390_n1088# 0.045353f
C252 plus.n31 a_n2390_n1088# 0.088017f
C253 plus.n32 a_n2390_n1088# 0.00593f
C254 plus.n33 a_n2390_n1088# 0.055247f
C255 plus.n34 a_n2390_n1088# 0.00593f
C256 plus.n35 a_n2390_n1088# 0.026132f
C257 plus.n36 a_n2390_n1088# 0.026132f
C258 plus.n37 a_n2390_n1088# 0.026132f
C259 plus.n38 a_n2390_n1088# 0.00593f
C260 plus.n39 a_n2390_n1088# 0.055247f
C261 plus.n40 a_n2390_n1088# 0.00593f
C262 plus.n41 a_n2390_n1088# 0.026132f
C263 plus.n42 a_n2390_n1088# 0.026132f
C264 plus.n43 a_n2390_n1088# 0.026132f
C265 plus.n44 a_n2390_n1088# 0.00593f
C266 plus.n45 a_n2390_n1088# 0.054522f
C267 plus.n46 a_n2390_n1088# 0.054119f
C268 plus.n47 a_n2390_n1088# 0.660005f
.ends

