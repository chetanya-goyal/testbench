* NGSPICE file created from diffpair468.ext - technology: sky130A

.subckt diffpair468 minus drain_right drain_left source plus
X0 source.t38 plus.t0 drain_left.t7 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X1 drain_left.t0 plus.t1 source.t37 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X2 source.t36 plus.t2 drain_left.t18 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X3 source.t9 minus.t0 drain_right.t19 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X4 source.t35 plus.t3 drain_left.t11 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X5 source.t11 minus.t1 drain_right.t18 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X6 drain_right.t17 minus.t2 source.t4 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X7 a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X8 drain_left.t19 plus.t4 source.t34 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X9 source.t33 plus.t5 drain_left.t6 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X10 source.t32 plus.t6 drain_left.t8 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X11 a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X12 drain_right.t16 minus.t3 source.t0 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X13 drain_right.t15 minus.t4 source.t1 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X14 drain_right.t14 minus.t5 source.t5 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X15 source.t31 plus.t7 drain_left.t5 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X16 drain_right.t13 minus.t6 source.t10 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X17 drain_left.t10 plus.t8 source.t30 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X18 drain_left.t9 plus.t9 source.t29 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X19 drain_right.t12 minus.t7 source.t8 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X20 a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X21 drain_left.t4 plus.t10 source.t28 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X22 source.t17 minus.t8 drain_right.t11 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X23 drain_right.t10 minus.t9 source.t18 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X24 drain_left.t17 plus.t11 source.t27 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X25 drain_left.t16 plus.t12 source.t26 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X26 drain_right.t9 minus.t10 source.t6 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X27 source.t25 plus.t13 drain_left.t14 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X28 drain_left.t1 plus.t14 source.t24 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X29 drain_left.t13 plus.t15 source.t23 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X30 a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X31 source.t12 minus.t11 drain_right.t8 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X32 drain_right.t7 minus.t12 source.t15 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X33 source.t14 minus.t13 drain_right.t6 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X34 source.t22 plus.t16 drain_left.t12 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X35 source.t13 minus.t14 drain_right.t5 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X36 drain_left.t2 plus.t17 source.t21 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X37 source.t7 minus.t15 drain_right.t4 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X38 source.t20 plus.t18 drain_left.t15 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X39 drain_right.t3 minus.t16 source.t3 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X40 source.t16 minus.t17 drain_right.t2 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X41 source.t2 minus.t18 drain_right.t1 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X42 source.t19 plus.t19 drain_left.t3 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X43 source.t39 minus.t19 drain_right.t0 a_n2982_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
R0 plus.n9 plus.t6 494.654
R1 plus.n43 plus.t17 494.654
R2 plus.n32 plus.t4 469.262
R3 plus.n30 plus.t19 469.262
R4 plus.n2 plus.t9 469.262
R5 plus.n24 plus.t2 469.262
R6 plus.n4 plus.t11 469.262
R7 plus.n18 plus.t5 469.262
R8 plus.n6 plus.t10 469.262
R9 plus.n12 plus.t3 469.262
R10 plus.n8 plus.t14 469.262
R11 plus.n66 plus.t13 469.262
R12 plus.n64 plus.t12 469.262
R13 plus.n36 plus.t16 469.262
R14 plus.n58 plus.t1 469.262
R15 plus.n38 plus.t0 469.262
R16 plus.n52 plus.t8 469.262
R17 plus.n40 plus.t7 469.262
R18 plus.n46 plus.t15 469.262
R19 plus.n42 plus.t18 469.262
R20 plus.n11 plus.n10 161.3
R21 plus.n12 plus.n7 161.3
R22 plus.n14 plus.n13 161.3
R23 plus.n15 plus.n6 161.3
R24 plus.n17 plus.n16 161.3
R25 plus.n18 plus.n5 161.3
R26 plus.n20 plus.n19 161.3
R27 plus.n21 plus.n4 161.3
R28 plus.n23 plus.n22 161.3
R29 plus.n24 plus.n3 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n27 plus.n2 161.3
R32 plus.n29 plus.n28 161.3
R33 plus.n30 plus.n1 161.3
R34 plus.n31 plus.n0 161.3
R35 plus.n33 plus.n32 161.3
R36 plus.n45 plus.n44 161.3
R37 plus.n46 plus.n41 161.3
R38 plus.n48 plus.n47 161.3
R39 plus.n49 plus.n40 161.3
R40 plus.n51 plus.n50 161.3
R41 plus.n52 plus.n39 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n55 plus.n38 161.3
R44 plus.n57 plus.n56 161.3
R45 plus.n58 plus.n37 161.3
R46 plus.n60 plus.n59 161.3
R47 plus.n61 plus.n36 161.3
R48 plus.n63 plus.n62 161.3
R49 plus.n64 plus.n35 161.3
R50 plus.n65 plus.n34 161.3
R51 plus.n67 plus.n66 161.3
R52 plus.n10 plus.n9 45.0031
R53 plus.n44 plus.n43 45.0031
R54 plus.n32 plus.n31 41.6278
R55 plus.n66 plus.n65 41.6278
R56 plus.n30 plus.n29 37.246
R57 plus.n11 plus.n8 37.246
R58 plus.n64 plus.n63 37.246
R59 plus.n45 plus.n42 37.246
R60 plus plus.n67 34.4649
R61 plus.n25 plus.n2 32.8641
R62 plus.n13 plus.n12 32.8641
R63 plus.n59 plus.n36 32.8641
R64 plus.n47 plus.n46 32.8641
R65 plus.n24 plus.n23 28.4823
R66 plus.n17 plus.n6 28.4823
R67 plus.n58 plus.n57 28.4823
R68 plus.n51 plus.n40 28.4823
R69 plus.n19 plus.n18 24.1005
R70 plus.n19 plus.n4 24.1005
R71 plus.n53 plus.n38 24.1005
R72 plus.n53 plus.n52 24.1005
R73 plus.n23 plus.n4 19.7187
R74 plus.n18 plus.n17 19.7187
R75 plus.n57 plus.n38 19.7187
R76 plus.n52 plus.n51 19.7187
R77 plus.n9 plus.n8 15.6319
R78 plus.n43 plus.n42 15.6319
R79 plus.n25 plus.n24 15.3369
R80 plus.n13 plus.n6 15.3369
R81 plus.n59 plus.n58 15.3369
R82 plus.n47 plus.n40 15.3369
R83 plus plus.n33 12.3111
R84 plus.n29 plus.n2 10.955
R85 plus.n12 plus.n11 10.955
R86 plus.n63 plus.n36 10.955
R87 plus.n46 plus.n45 10.955
R88 plus.n31 plus.n30 6.57323
R89 plus.n65 plus.n64 6.57323
R90 plus.n10 plus.n7 0.189894
R91 plus.n14 plus.n7 0.189894
R92 plus.n15 plus.n14 0.189894
R93 plus.n16 plus.n15 0.189894
R94 plus.n16 plus.n5 0.189894
R95 plus.n20 plus.n5 0.189894
R96 plus.n21 plus.n20 0.189894
R97 plus.n22 plus.n21 0.189894
R98 plus.n22 plus.n3 0.189894
R99 plus.n26 plus.n3 0.189894
R100 plus.n27 plus.n26 0.189894
R101 plus.n28 plus.n27 0.189894
R102 plus.n28 plus.n1 0.189894
R103 plus.n1 plus.n0 0.189894
R104 plus.n33 plus.n0 0.189894
R105 plus.n67 plus.n34 0.189894
R106 plus.n35 plus.n34 0.189894
R107 plus.n62 plus.n35 0.189894
R108 plus.n62 plus.n61 0.189894
R109 plus.n61 plus.n60 0.189894
R110 plus.n60 plus.n37 0.189894
R111 plus.n56 plus.n37 0.189894
R112 plus.n56 plus.n55 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n39 0.189894
R115 plus.n50 plus.n39 0.189894
R116 plus.n50 plus.n49 0.189894
R117 plus.n49 plus.n48 0.189894
R118 plus.n48 plus.n41 0.189894
R119 plus.n44 plus.n41 0.189894
R120 drain_left.n10 drain_left.n8 60.4406
R121 drain_left.n6 drain_left.n4 60.4404
R122 drain_left.n2 drain_left.n0 60.4404
R123 drain_left.n14 drain_left.n13 59.5527
R124 drain_left.n12 drain_left.n11 59.5527
R125 drain_left.n10 drain_left.n9 59.5527
R126 drain_left.n7 drain_left.n3 59.5525
R127 drain_left.n6 drain_left.n5 59.5525
R128 drain_left.n2 drain_left.n1 59.5525
R129 drain_left.n16 drain_left.n15 59.5525
R130 drain_left drain_left.n7 34.4705
R131 drain_left drain_left.n16 6.54115
R132 drain_left.n3 drain_left.t7 1.6505
R133 drain_left.n3 drain_left.t10 1.6505
R134 drain_left.n4 drain_left.t15 1.6505
R135 drain_left.n4 drain_left.t2 1.6505
R136 drain_left.n5 drain_left.t5 1.6505
R137 drain_left.n5 drain_left.t13 1.6505
R138 drain_left.n1 drain_left.t12 1.6505
R139 drain_left.n1 drain_left.t0 1.6505
R140 drain_left.n0 drain_left.t14 1.6505
R141 drain_left.n0 drain_left.t16 1.6505
R142 drain_left.n15 drain_left.t3 1.6505
R143 drain_left.n15 drain_left.t19 1.6505
R144 drain_left.n13 drain_left.t18 1.6505
R145 drain_left.n13 drain_left.t9 1.6505
R146 drain_left.n11 drain_left.t6 1.6505
R147 drain_left.n11 drain_left.t17 1.6505
R148 drain_left.n9 drain_left.t11 1.6505
R149 drain_left.n9 drain_left.t4 1.6505
R150 drain_left.n8 drain_left.t8 1.6505
R151 drain_left.n8 drain_left.t1 1.6505
R152 drain_left.n12 drain_left.n10 0.888431
R153 drain_left.n14 drain_left.n12 0.888431
R154 drain_left.n16 drain_left.n14 0.888431
R155 drain_left.n7 drain_left.n6 0.833085
R156 drain_left.n7 drain_left.n2 0.833085
R157 source.n554 source.n494 289.615
R158 source.n480 source.n420 289.615
R159 source.n414 source.n354 289.615
R160 source.n340 source.n280 289.615
R161 source.n60 source.n0 289.615
R162 source.n134 source.n74 289.615
R163 source.n200 source.n140 289.615
R164 source.n274 source.n214 289.615
R165 source.n514 source.n513 185
R166 source.n519 source.n518 185
R167 source.n521 source.n520 185
R168 source.n510 source.n509 185
R169 source.n527 source.n526 185
R170 source.n529 source.n528 185
R171 source.n506 source.n505 185
R172 source.n536 source.n535 185
R173 source.n537 source.n504 185
R174 source.n539 source.n538 185
R175 source.n502 source.n501 185
R176 source.n545 source.n544 185
R177 source.n547 source.n546 185
R178 source.n498 source.n497 185
R179 source.n553 source.n552 185
R180 source.n555 source.n554 185
R181 source.n440 source.n439 185
R182 source.n445 source.n444 185
R183 source.n447 source.n446 185
R184 source.n436 source.n435 185
R185 source.n453 source.n452 185
R186 source.n455 source.n454 185
R187 source.n432 source.n431 185
R188 source.n462 source.n461 185
R189 source.n463 source.n430 185
R190 source.n465 source.n464 185
R191 source.n428 source.n427 185
R192 source.n471 source.n470 185
R193 source.n473 source.n472 185
R194 source.n424 source.n423 185
R195 source.n479 source.n478 185
R196 source.n481 source.n480 185
R197 source.n374 source.n373 185
R198 source.n379 source.n378 185
R199 source.n381 source.n380 185
R200 source.n370 source.n369 185
R201 source.n387 source.n386 185
R202 source.n389 source.n388 185
R203 source.n366 source.n365 185
R204 source.n396 source.n395 185
R205 source.n397 source.n364 185
R206 source.n399 source.n398 185
R207 source.n362 source.n361 185
R208 source.n405 source.n404 185
R209 source.n407 source.n406 185
R210 source.n358 source.n357 185
R211 source.n413 source.n412 185
R212 source.n415 source.n414 185
R213 source.n300 source.n299 185
R214 source.n305 source.n304 185
R215 source.n307 source.n306 185
R216 source.n296 source.n295 185
R217 source.n313 source.n312 185
R218 source.n315 source.n314 185
R219 source.n292 source.n291 185
R220 source.n322 source.n321 185
R221 source.n323 source.n290 185
R222 source.n325 source.n324 185
R223 source.n288 source.n287 185
R224 source.n331 source.n330 185
R225 source.n333 source.n332 185
R226 source.n284 source.n283 185
R227 source.n339 source.n338 185
R228 source.n341 source.n340 185
R229 source.n61 source.n60 185
R230 source.n59 source.n58 185
R231 source.n4 source.n3 185
R232 source.n53 source.n52 185
R233 source.n51 source.n50 185
R234 source.n8 source.n7 185
R235 source.n45 source.n44 185
R236 source.n43 source.n10 185
R237 source.n42 source.n41 185
R238 source.n13 source.n11 185
R239 source.n36 source.n35 185
R240 source.n34 source.n33 185
R241 source.n17 source.n16 185
R242 source.n28 source.n27 185
R243 source.n26 source.n25 185
R244 source.n21 source.n20 185
R245 source.n135 source.n134 185
R246 source.n133 source.n132 185
R247 source.n78 source.n77 185
R248 source.n127 source.n126 185
R249 source.n125 source.n124 185
R250 source.n82 source.n81 185
R251 source.n119 source.n118 185
R252 source.n117 source.n84 185
R253 source.n116 source.n115 185
R254 source.n87 source.n85 185
R255 source.n110 source.n109 185
R256 source.n108 source.n107 185
R257 source.n91 source.n90 185
R258 source.n102 source.n101 185
R259 source.n100 source.n99 185
R260 source.n95 source.n94 185
R261 source.n201 source.n200 185
R262 source.n199 source.n198 185
R263 source.n144 source.n143 185
R264 source.n193 source.n192 185
R265 source.n191 source.n190 185
R266 source.n148 source.n147 185
R267 source.n185 source.n184 185
R268 source.n183 source.n150 185
R269 source.n182 source.n181 185
R270 source.n153 source.n151 185
R271 source.n176 source.n175 185
R272 source.n174 source.n173 185
R273 source.n157 source.n156 185
R274 source.n168 source.n167 185
R275 source.n166 source.n165 185
R276 source.n161 source.n160 185
R277 source.n275 source.n274 185
R278 source.n273 source.n272 185
R279 source.n218 source.n217 185
R280 source.n267 source.n266 185
R281 source.n265 source.n264 185
R282 source.n222 source.n221 185
R283 source.n259 source.n258 185
R284 source.n257 source.n224 185
R285 source.n256 source.n255 185
R286 source.n227 source.n225 185
R287 source.n250 source.n249 185
R288 source.n248 source.n247 185
R289 source.n231 source.n230 185
R290 source.n242 source.n241 185
R291 source.n240 source.n239 185
R292 source.n235 source.n234 185
R293 source.n515 source.t0 149.524
R294 source.n441 source.t9 149.524
R295 source.n375 source.t21 149.524
R296 source.n301 source.t25 149.524
R297 source.n22 source.t34 149.524
R298 source.n96 source.t32 149.524
R299 source.n162 source.t6 149.524
R300 source.n236 source.t12 149.524
R301 source.n519 source.n513 104.615
R302 source.n520 source.n519 104.615
R303 source.n520 source.n509 104.615
R304 source.n527 source.n509 104.615
R305 source.n528 source.n527 104.615
R306 source.n528 source.n505 104.615
R307 source.n536 source.n505 104.615
R308 source.n537 source.n536 104.615
R309 source.n538 source.n537 104.615
R310 source.n538 source.n501 104.615
R311 source.n545 source.n501 104.615
R312 source.n546 source.n545 104.615
R313 source.n546 source.n497 104.615
R314 source.n553 source.n497 104.615
R315 source.n554 source.n553 104.615
R316 source.n445 source.n439 104.615
R317 source.n446 source.n445 104.615
R318 source.n446 source.n435 104.615
R319 source.n453 source.n435 104.615
R320 source.n454 source.n453 104.615
R321 source.n454 source.n431 104.615
R322 source.n462 source.n431 104.615
R323 source.n463 source.n462 104.615
R324 source.n464 source.n463 104.615
R325 source.n464 source.n427 104.615
R326 source.n471 source.n427 104.615
R327 source.n472 source.n471 104.615
R328 source.n472 source.n423 104.615
R329 source.n479 source.n423 104.615
R330 source.n480 source.n479 104.615
R331 source.n379 source.n373 104.615
R332 source.n380 source.n379 104.615
R333 source.n380 source.n369 104.615
R334 source.n387 source.n369 104.615
R335 source.n388 source.n387 104.615
R336 source.n388 source.n365 104.615
R337 source.n396 source.n365 104.615
R338 source.n397 source.n396 104.615
R339 source.n398 source.n397 104.615
R340 source.n398 source.n361 104.615
R341 source.n405 source.n361 104.615
R342 source.n406 source.n405 104.615
R343 source.n406 source.n357 104.615
R344 source.n413 source.n357 104.615
R345 source.n414 source.n413 104.615
R346 source.n305 source.n299 104.615
R347 source.n306 source.n305 104.615
R348 source.n306 source.n295 104.615
R349 source.n313 source.n295 104.615
R350 source.n314 source.n313 104.615
R351 source.n314 source.n291 104.615
R352 source.n322 source.n291 104.615
R353 source.n323 source.n322 104.615
R354 source.n324 source.n323 104.615
R355 source.n324 source.n287 104.615
R356 source.n331 source.n287 104.615
R357 source.n332 source.n331 104.615
R358 source.n332 source.n283 104.615
R359 source.n339 source.n283 104.615
R360 source.n340 source.n339 104.615
R361 source.n60 source.n59 104.615
R362 source.n59 source.n3 104.615
R363 source.n52 source.n3 104.615
R364 source.n52 source.n51 104.615
R365 source.n51 source.n7 104.615
R366 source.n44 source.n7 104.615
R367 source.n44 source.n43 104.615
R368 source.n43 source.n42 104.615
R369 source.n42 source.n11 104.615
R370 source.n35 source.n11 104.615
R371 source.n35 source.n34 104.615
R372 source.n34 source.n16 104.615
R373 source.n27 source.n16 104.615
R374 source.n27 source.n26 104.615
R375 source.n26 source.n20 104.615
R376 source.n134 source.n133 104.615
R377 source.n133 source.n77 104.615
R378 source.n126 source.n77 104.615
R379 source.n126 source.n125 104.615
R380 source.n125 source.n81 104.615
R381 source.n118 source.n81 104.615
R382 source.n118 source.n117 104.615
R383 source.n117 source.n116 104.615
R384 source.n116 source.n85 104.615
R385 source.n109 source.n85 104.615
R386 source.n109 source.n108 104.615
R387 source.n108 source.n90 104.615
R388 source.n101 source.n90 104.615
R389 source.n101 source.n100 104.615
R390 source.n100 source.n94 104.615
R391 source.n200 source.n199 104.615
R392 source.n199 source.n143 104.615
R393 source.n192 source.n143 104.615
R394 source.n192 source.n191 104.615
R395 source.n191 source.n147 104.615
R396 source.n184 source.n147 104.615
R397 source.n184 source.n183 104.615
R398 source.n183 source.n182 104.615
R399 source.n182 source.n151 104.615
R400 source.n175 source.n151 104.615
R401 source.n175 source.n174 104.615
R402 source.n174 source.n156 104.615
R403 source.n167 source.n156 104.615
R404 source.n167 source.n166 104.615
R405 source.n166 source.n160 104.615
R406 source.n274 source.n273 104.615
R407 source.n273 source.n217 104.615
R408 source.n266 source.n217 104.615
R409 source.n266 source.n265 104.615
R410 source.n265 source.n221 104.615
R411 source.n258 source.n221 104.615
R412 source.n258 source.n257 104.615
R413 source.n257 source.n256 104.615
R414 source.n256 source.n225 104.615
R415 source.n249 source.n225 104.615
R416 source.n249 source.n248 104.615
R417 source.n248 source.n230 104.615
R418 source.n241 source.n230 104.615
R419 source.n241 source.n240 104.615
R420 source.n240 source.n234 104.615
R421 source.t0 source.n513 52.3082
R422 source.t9 source.n439 52.3082
R423 source.t21 source.n373 52.3082
R424 source.t25 source.n299 52.3082
R425 source.t34 source.n20 52.3082
R426 source.t32 source.n94 52.3082
R427 source.t6 source.n160 52.3082
R428 source.t12 source.n234 52.3082
R429 source.n67 source.n66 42.8739
R430 source.n69 source.n68 42.8739
R431 source.n71 source.n70 42.8739
R432 source.n73 source.n72 42.8739
R433 source.n207 source.n206 42.8739
R434 source.n209 source.n208 42.8739
R435 source.n211 source.n210 42.8739
R436 source.n213 source.n212 42.8739
R437 source.n493 source.n492 42.8737
R438 source.n491 source.n490 42.8737
R439 source.n489 source.n488 42.8737
R440 source.n487 source.n486 42.8737
R441 source.n353 source.n352 42.8737
R442 source.n351 source.n350 42.8737
R443 source.n349 source.n348 42.8737
R444 source.n347 source.n346 42.8737
R445 source.n559 source.n558 29.8581
R446 source.n485 source.n484 29.8581
R447 source.n419 source.n418 29.8581
R448 source.n345 source.n344 29.8581
R449 source.n65 source.n64 29.8581
R450 source.n139 source.n138 29.8581
R451 source.n205 source.n204 29.8581
R452 source.n279 source.n278 29.8581
R453 source.n345 source.n279 22.1757
R454 source.n560 source.n65 16.4688
R455 source.n539 source.n504 13.1884
R456 source.n465 source.n430 13.1884
R457 source.n399 source.n364 13.1884
R458 source.n325 source.n290 13.1884
R459 source.n45 source.n10 13.1884
R460 source.n119 source.n84 13.1884
R461 source.n185 source.n150 13.1884
R462 source.n259 source.n224 13.1884
R463 source.n535 source.n534 12.8005
R464 source.n540 source.n502 12.8005
R465 source.n461 source.n460 12.8005
R466 source.n466 source.n428 12.8005
R467 source.n395 source.n394 12.8005
R468 source.n400 source.n362 12.8005
R469 source.n321 source.n320 12.8005
R470 source.n326 source.n288 12.8005
R471 source.n46 source.n8 12.8005
R472 source.n41 source.n12 12.8005
R473 source.n120 source.n82 12.8005
R474 source.n115 source.n86 12.8005
R475 source.n186 source.n148 12.8005
R476 source.n181 source.n152 12.8005
R477 source.n260 source.n222 12.8005
R478 source.n255 source.n226 12.8005
R479 source.n533 source.n506 12.0247
R480 source.n544 source.n543 12.0247
R481 source.n459 source.n432 12.0247
R482 source.n470 source.n469 12.0247
R483 source.n393 source.n366 12.0247
R484 source.n404 source.n403 12.0247
R485 source.n319 source.n292 12.0247
R486 source.n330 source.n329 12.0247
R487 source.n50 source.n49 12.0247
R488 source.n40 source.n13 12.0247
R489 source.n124 source.n123 12.0247
R490 source.n114 source.n87 12.0247
R491 source.n190 source.n189 12.0247
R492 source.n180 source.n153 12.0247
R493 source.n264 source.n263 12.0247
R494 source.n254 source.n227 12.0247
R495 source.n530 source.n529 11.249
R496 source.n547 source.n500 11.249
R497 source.n456 source.n455 11.249
R498 source.n473 source.n426 11.249
R499 source.n390 source.n389 11.249
R500 source.n407 source.n360 11.249
R501 source.n316 source.n315 11.249
R502 source.n333 source.n286 11.249
R503 source.n53 source.n6 11.249
R504 source.n37 source.n36 11.249
R505 source.n127 source.n80 11.249
R506 source.n111 source.n110 11.249
R507 source.n193 source.n146 11.249
R508 source.n177 source.n176 11.249
R509 source.n267 source.n220 11.249
R510 source.n251 source.n250 11.249
R511 source.n526 source.n508 10.4732
R512 source.n548 source.n498 10.4732
R513 source.n452 source.n434 10.4732
R514 source.n474 source.n424 10.4732
R515 source.n386 source.n368 10.4732
R516 source.n408 source.n358 10.4732
R517 source.n312 source.n294 10.4732
R518 source.n334 source.n284 10.4732
R519 source.n54 source.n4 10.4732
R520 source.n33 source.n15 10.4732
R521 source.n128 source.n78 10.4732
R522 source.n107 source.n89 10.4732
R523 source.n194 source.n144 10.4732
R524 source.n173 source.n155 10.4732
R525 source.n268 source.n218 10.4732
R526 source.n247 source.n229 10.4732
R527 source.n515 source.n514 10.2747
R528 source.n441 source.n440 10.2747
R529 source.n375 source.n374 10.2747
R530 source.n301 source.n300 10.2747
R531 source.n22 source.n21 10.2747
R532 source.n96 source.n95 10.2747
R533 source.n162 source.n161 10.2747
R534 source.n236 source.n235 10.2747
R535 source.n525 source.n510 9.69747
R536 source.n552 source.n551 9.69747
R537 source.n451 source.n436 9.69747
R538 source.n478 source.n477 9.69747
R539 source.n385 source.n370 9.69747
R540 source.n412 source.n411 9.69747
R541 source.n311 source.n296 9.69747
R542 source.n338 source.n337 9.69747
R543 source.n58 source.n57 9.69747
R544 source.n32 source.n17 9.69747
R545 source.n132 source.n131 9.69747
R546 source.n106 source.n91 9.69747
R547 source.n198 source.n197 9.69747
R548 source.n172 source.n157 9.69747
R549 source.n272 source.n271 9.69747
R550 source.n246 source.n231 9.69747
R551 source.n558 source.n557 9.45567
R552 source.n484 source.n483 9.45567
R553 source.n418 source.n417 9.45567
R554 source.n344 source.n343 9.45567
R555 source.n64 source.n63 9.45567
R556 source.n138 source.n137 9.45567
R557 source.n204 source.n203 9.45567
R558 source.n278 source.n277 9.45567
R559 source.n557 source.n556 9.3005
R560 source.n496 source.n495 9.3005
R561 source.n551 source.n550 9.3005
R562 source.n549 source.n548 9.3005
R563 source.n500 source.n499 9.3005
R564 source.n543 source.n542 9.3005
R565 source.n541 source.n540 9.3005
R566 source.n517 source.n516 9.3005
R567 source.n512 source.n511 9.3005
R568 source.n523 source.n522 9.3005
R569 source.n525 source.n524 9.3005
R570 source.n508 source.n507 9.3005
R571 source.n531 source.n530 9.3005
R572 source.n533 source.n532 9.3005
R573 source.n534 source.n503 9.3005
R574 source.n483 source.n482 9.3005
R575 source.n422 source.n421 9.3005
R576 source.n477 source.n476 9.3005
R577 source.n475 source.n474 9.3005
R578 source.n426 source.n425 9.3005
R579 source.n469 source.n468 9.3005
R580 source.n467 source.n466 9.3005
R581 source.n443 source.n442 9.3005
R582 source.n438 source.n437 9.3005
R583 source.n449 source.n448 9.3005
R584 source.n451 source.n450 9.3005
R585 source.n434 source.n433 9.3005
R586 source.n457 source.n456 9.3005
R587 source.n459 source.n458 9.3005
R588 source.n460 source.n429 9.3005
R589 source.n417 source.n416 9.3005
R590 source.n356 source.n355 9.3005
R591 source.n411 source.n410 9.3005
R592 source.n409 source.n408 9.3005
R593 source.n360 source.n359 9.3005
R594 source.n403 source.n402 9.3005
R595 source.n401 source.n400 9.3005
R596 source.n377 source.n376 9.3005
R597 source.n372 source.n371 9.3005
R598 source.n383 source.n382 9.3005
R599 source.n385 source.n384 9.3005
R600 source.n368 source.n367 9.3005
R601 source.n391 source.n390 9.3005
R602 source.n393 source.n392 9.3005
R603 source.n394 source.n363 9.3005
R604 source.n343 source.n342 9.3005
R605 source.n282 source.n281 9.3005
R606 source.n337 source.n336 9.3005
R607 source.n335 source.n334 9.3005
R608 source.n286 source.n285 9.3005
R609 source.n329 source.n328 9.3005
R610 source.n327 source.n326 9.3005
R611 source.n303 source.n302 9.3005
R612 source.n298 source.n297 9.3005
R613 source.n309 source.n308 9.3005
R614 source.n311 source.n310 9.3005
R615 source.n294 source.n293 9.3005
R616 source.n317 source.n316 9.3005
R617 source.n319 source.n318 9.3005
R618 source.n320 source.n289 9.3005
R619 source.n24 source.n23 9.3005
R620 source.n19 source.n18 9.3005
R621 source.n30 source.n29 9.3005
R622 source.n32 source.n31 9.3005
R623 source.n15 source.n14 9.3005
R624 source.n38 source.n37 9.3005
R625 source.n40 source.n39 9.3005
R626 source.n12 source.n9 9.3005
R627 source.n63 source.n62 9.3005
R628 source.n2 source.n1 9.3005
R629 source.n57 source.n56 9.3005
R630 source.n55 source.n54 9.3005
R631 source.n6 source.n5 9.3005
R632 source.n49 source.n48 9.3005
R633 source.n47 source.n46 9.3005
R634 source.n98 source.n97 9.3005
R635 source.n93 source.n92 9.3005
R636 source.n104 source.n103 9.3005
R637 source.n106 source.n105 9.3005
R638 source.n89 source.n88 9.3005
R639 source.n112 source.n111 9.3005
R640 source.n114 source.n113 9.3005
R641 source.n86 source.n83 9.3005
R642 source.n137 source.n136 9.3005
R643 source.n76 source.n75 9.3005
R644 source.n131 source.n130 9.3005
R645 source.n129 source.n128 9.3005
R646 source.n80 source.n79 9.3005
R647 source.n123 source.n122 9.3005
R648 source.n121 source.n120 9.3005
R649 source.n164 source.n163 9.3005
R650 source.n159 source.n158 9.3005
R651 source.n170 source.n169 9.3005
R652 source.n172 source.n171 9.3005
R653 source.n155 source.n154 9.3005
R654 source.n178 source.n177 9.3005
R655 source.n180 source.n179 9.3005
R656 source.n152 source.n149 9.3005
R657 source.n203 source.n202 9.3005
R658 source.n142 source.n141 9.3005
R659 source.n197 source.n196 9.3005
R660 source.n195 source.n194 9.3005
R661 source.n146 source.n145 9.3005
R662 source.n189 source.n188 9.3005
R663 source.n187 source.n186 9.3005
R664 source.n238 source.n237 9.3005
R665 source.n233 source.n232 9.3005
R666 source.n244 source.n243 9.3005
R667 source.n246 source.n245 9.3005
R668 source.n229 source.n228 9.3005
R669 source.n252 source.n251 9.3005
R670 source.n254 source.n253 9.3005
R671 source.n226 source.n223 9.3005
R672 source.n277 source.n276 9.3005
R673 source.n216 source.n215 9.3005
R674 source.n271 source.n270 9.3005
R675 source.n269 source.n268 9.3005
R676 source.n220 source.n219 9.3005
R677 source.n263 source.n262 9.3005
R678 source.n261 source.n260 9.3005
R679 source.n522 source.n521 8.92171
R680 source.n555 source.n496 8.92171
R681 source.n448 source.n447 8.92171
R682 source.n481 source.n422 8.92171
R683 source.n382 source.n381 8.92171
R684 source.n415 source.n356 8.92171
R685 source.n308 source.n307 8.92171
R686 source.n341 source.n282 8.92171
R687 source.n61 source.n2 8.92171
R688 source.n29 source.n28 8.92171
R689 source.n135 source.n76 8.92171
R690 source.n103 source.n102 8.92171
R691 source.n201 source.n142 8.92171
R692 source.n169 source.n168 8.92171
R693 source.n275 source.n216 8.92171
R694 source.n243 source.n242 8.92171
R695 source.n518 source.n512 8.14595
R696 source.n556 source.n494 8.14595
R697 source.n444 source.n438 8.14595
R698 source.n482 source.n420 8.14595
R699 source.n378 source.n372 8.14595
R700 source.n416 source.n354 8.14595
R701 source.n304 source.n298 8.14595
R702 source.n342 source.n280 8.14595
R703 source.n62 source.n0 8.14595
R704 source.n25 source.n19 8.14595
R705 source.n136 source.n74 8.14595
R706 source.n99 source.n93 8.14595
R707 source.n202 source.n140 8.14595
R708 source.n165 source.n159 8.14595
R709 source.n276 source.n214 8.14595
R710 source.n239 source.n233 8.14595
R711 source.n517 source.n514 7.3702
R712 source.n443 source.n440 7.3702
R713 source.n377 source.n374 7.3702
R714 source.n303 source.n300 7.3702
R715 source.n24 source.n21 7.3702
R716 source.n98 source.n95 7.3702
R717 source.n164 source.n161 7.3702
R718 source.n238 source.n235 7.3702
R719 source.n518 source.n517 5.81868
R720 source.n558 source.n494 5.81868
R721 source.n444 source.n443 5.81868
R722 source.n484 source.n420 5.81868
R723 source.n378 source.n377 5.81868
R724 source.n418 source.n354 5.81868
R725 source.n304 source.n303 5.81868
R726 source.n344 source.n280 5.81868
R727 source.n64 source.n0 5.81868
R728 source.n25 source.n24 5.81868
R729 source.n138 source.n74 5.81868
R730 source.n99 source.n98 5.81868
R731 source.n204 source.n140 5.81868
R732 source.n165 source.n164 5.81868
R733 source.n278 source.n214 5.81868
R734 source.n239 source.n238 5.81868
R735 source.n560 source.n559 5.7074
R736 source.n521 source.n512 5.04292
R737 source.n556 source.n555 5.04292
R738 source.n447 source.n438 5.04292
R739 source.n482 source.n481 5.04292
R740 source.n381 source.n372 5.04292
R741 source.n416 source.n415 5.04292
R742 source.n307 source.n298 5.04292
R743 source.n342 source.n341 5.04292
R744 source.n62 source.n61 5.04292
R745 source.n28 source.n19 5.04292
R746 source.n136 source.n135 5.04292
R747 source.n102 source.n93 5.04292
R748 source.n202 source.n201 5.04292
R749 source.n168 source.n159 5.04292
R750 source.n276 source.n275 5.04292
R751 source.n242 source.n233 5.04292
R752 source.n522 source.n510 4.26717
R753 source.n552 source.n496 4.26717
R754 source.n448 source.n436 4.26717
R755 source.n478 source.n422 4.26717
R756 source.n382 source.n370 4.26717
R757 source.n412 source.n356 4.26717
R758 source.n308 source.n296 4.26717
R759 source.n338 source.n282 4.26717
R760 source.n58 source.n2 4.26717
R761 source.n29 source.n17 4.26717
R762 source.n132 source.n76 4.26717
R763 source.n103 source.n91 4.26717
R764 source.n198 source.n142 4.26717
R765 source.n169 source.n157 4.26717
R766 source.n272 source.n216 4.26717
R767 source.n243 source.n231 4.26717
R768 source.n526 source.n525 3.49141
R769 source.n551 source.n498 3.49141
R770 source.n452 source.n451 3.49141
R771 source.n477 source.n424 3.49141
R772 source.n386 source.n385 3.49141
R773 source.n411 source.n358 3.49141
R774 source.n312 source.n311 3.49141
R775 source.n337 source.n284 3.49141
R776 source.n57 source.n4 3.49141
R777 source.n33 source.n32 3.49141
R778 source.n131 source.n78 3.49141
R779 source.n107 source.n106 3.49141
R780 source.n197 source.n144 3.49141
R781 source.n173 source.n172 3.49141
R782 source.n271 source.n218 3.49141
R783 source.n247 source.n246 3.49141
R784 source.n516 source.n515 2.84303
R785 source.n442 source.n441 2.84303
R786 source.n376 source.n375 2.84303
R787 source.n302 source.n301 2.84303
R788 source.n23 source.n22 2.84303
R789 source.n97 source.n96 2.84303
R790 source.n163 source.n162 2.84303
R791 source.n237 source.n236 2.84303
R792 source.n529 source.n508 2.71565
R793 source.n548 source.n547 2.71565
R794 source.n455 source.n434 2.71565
R795 source.n474 source.n473 2.71565
R796 source.n389 source.n368 2.71565
R797 source.n408 source.n407 2.71565
R798 source.n315 source.n294 2.71565
R799 source.n334 source.n333 2.71565
R800 source.n54 source.n53 2.71565
R801 source.n36 source.n15 2.71565
R802 source.n128 source.n127 2.71565
R803 source.n110 source.n89 2.71565
R804 source.n194 source.n193 2.71565
R805 source.n176 source.n155 2.71565
R806 source.n268 source.n267 2.71565
R807 source.n250 source.n229 2.71565
R808 source.n530 source.n506 1.93989
R809 source.n544 source.n500 1.93989
R810 source.n456 source.n432 1.93989
R811 source.n470 source.n426 1.93989
R812 source.n390 source.n366 1.93989
R813 source.n404 source.n360 1.93989
R814 source.n316 source.n292 1.93989
R815 source.n330 source.n286 1.93989
R816 source.n50 source.n6 1.93989
R817 source.n37 source.n13 1.93989
R818 source.n124 source.n80 1.93989
R819 source.n111 source.n87 1.93989
R820 source.n190 source.n146 1.93989
R821 source.n177 source.n153 1.93989
R822 source.n264 source.n220 1.93989
R823 source.n251 source.n227 1.93989
R824 source.n492 source.t18 1.6505
R825 source.n492 source.t17 1.6505
R826 source.n490 source.t15 1.6505
R827 source.n490 source.t14 1.6505
R828 source.n488 source.t3 1.6505
R829 source.n488 source.t39 1.6505
R830 source.n486 source.t4 1.6505
R831 source.n486 source.t7 1.6505
R832 source.n352 source.t23 1.6505
R833 source.n352 source.t20 1.6505
R834 source.n350 source.t30 1.6505
R835 source.n350 source.t31 1.6505
R836 source.n348 source.t37 1.6505
R837 source.n348 source.t38 1.6505
R838 source.n346 source.t26 1.6505
R839 source.n346 source.t22 1.6505
R840 source.n66 source.t29 1.6505
R841 source.n66 source.t19 1.6505
R842 source.n68 source.t27 1.6505
R843 source.n68 source.t36 1.6505
R844 source.n70 source.t28 1.6505
R845 source.n70 source.t33 1.6505
R846 source.n72 source.t24 1.6505
R847 source.n72 source.t35 1.6505
R848 source.n206 source.t8 1.6505
R849 source.n206 source.t11 1.6505
R850 source.n208 source.t10 1.6505
R851 source.n208 source.t16 1.6505
R852 source.n210 source.t5 1.6505
R853 source.n210 source.t2 1.6505
R854 source.n212 source.t1 1.6505
R855 source.n212 source.t13 1.6505
R856 source.n535 source.n533 1.16414
R857 source.n543 source.n502 1.16414
R858 source.n461 source.n459 1.16414
R859 source.n469 source.n428 1.16414
R860 source.n395 source.n393 1.16414
R861 source.n403 source.n362 1.16414
R862 source.n321 source.n319 1.16414
R863 source.n329 source.n288 1.16414
R864 source.n49 source.n8 1.16414
R865 source.n41 source.n40 1.16414
R866 source.n123 source.n82 1.16414
R867 source.n115 source.n114 1.16414
R868 source.n189 source.n148 1.16414
R869 source.n181 source.n180 1.16414
R870 source.n263 source.n222 1.16414
R871 source.n255 source.n254 1.16414
R872 source.n279 source.n213 0.888431
R873 source.n213 source.n211 0.888431
R874 source.n211 source.n209 0.888431
R875 source.n209 source.n207 0.888431
R876 source.n207 source.n205 0.888431
R877 source.n139 source.n73 0.888431
R878 source.n73 source.n71 0.888431
R879 source.n71 source.n69 0.888431
R880 source.n69 source.n67 0.888431
R881 source.n67 source.n65 0.888431
R882 source.n347 source.n345 0.888431
R883 source.n349 source.n347 0.888431
R884 source.n351 source.n349 0.888431
R885 source.n353 source.n351 0.888431
R886 source.n419 source.n353 0.888431
R887 source.n487 source.n485 0.888431
R888 source.n489 source.n487 0.888431
R889 source.n491 source.n489 0.888431
R890 source.n493 source.n491 0.888431
R891 source.n559 source.n493 0.888431
R892 source.n205 source.n139 0.470328
R893 source.n485 source.n419 0.470328
R894 source.n534 source.n504 0.388379
R895 source.n540 source.n539 0.388379
R896 source.n460 source.n430 0.388379
R897 source.n466 source.n465 0.388379
R898 source.n394 source.n364 0.388379
R899 source.n400 source.n399 0.388379
R900 source.n320 source.n290 0.388379
R901 source.n326 source.n325 0.388379
R902 source.n46 source.n45 0.388379
R903 source.n12 source.n10 0.388379
R904 source.n120 source.n119 0.388379
R905 source.n86 source.n84 0.388379
R906 source.n186 source.n185 0.388379
R907 source.n152 source.n150 0.388379
R908 source.n260 source.n259 0.388379
R909 source.n226 source.n224 0.388379
R910 source source.n560 0.188
R911 source.n516 source.n511 0.155672
R912 source.n523 source.n511 0.155672
R913 source.n524 source.n523 0.155672
R914 source.n524 source.n507 0.155672
R915 source.n531 source.n507 0.155672
R916 source.n532 source.n531 0.155672
R917 source.n532 source.n503 0.155672
R918 source.n541 source.n503 0.155672
R919 source.n542 source.n541 0.155672
R920 source.n542 source.n499 0.155672
R921 source.n549 source.n499 0.155672
R922 source.n550 source.n549 0.155672
R923 source.n550 source.n495 0.155672
R924 source.n557 source.n495 0.155672
R925 source.n442 source.n437 0.155672
R926 source.n449 source.n437 0.155672
R927 source.n450 source.n449 0.155672
R928 source.n450 source.n433 0.155672
R929 source.n457 source.n433 0.155672
R930 source.n458 source.n457 0.155672
R931 source.n458 source.n429 0.155672
R932 source.n467 source.n429 0.155672
R933 source.n468 source.n467 0.155672
R934 source.n468 source.n425 0.155672
R935 source.n475 source.n425 0.155672
R936 source.n476 source.n475 0.155672
R937 source.n476 source.n421 0.155672
R938 source.n483 source.n421 0.155672
R939 source.n376 source.n371 0.155672
R940 source.n383 source.n371 0.155672
R941 source.n384 source.n383 0.155672
R942 source.n384 source.n367 0.155672
R943 source.n391 source.n367 0.155672
R944 source.n392 source.n391 0.155672
R945 source.n392 source.n363 0.155672
R946 source.n401 source.n363 0.155672
R947 source.n402 source.n401 0.155672
R948 source.n402 source.n359 0.155672
R949 source.n409 source.n359 0.155672
R950 source.n410 source.n409 0.155672
R951 source.n410 source.n355 0.155672
R952 source.n417 source.n355 0.155672
R953 source.n302 source.n297 0.155672
R954 source.n309 source.n297 0.155672
R955 source.n310 source.n309 0.155672
R956 source.n310 source.n293 0.155672
R957 source.n317 source.n293 0.155672
R958 source.n318 source.n317 0.155672
R959 source.n318 source.n289 0.155672
R960 source.n327 source.n289 0.155672
R961 source.n328 source.n327 0.155672
R962 source.n328 source.n285 0.155672
R963 source.n335 source.n285 0.155672
R964 source.n336 source.n335 0.155672
R965 source.n336 source.n281 0.155672
R966 source.n343 source.n281 0.155672
R967 source.n63 source.n1 0.155672
R968 source.n56 source.n1 0.155672
R969 source.n56 source.n55 0.155672
R970 source.n55 source.n5 0.155672
R971 source.n48 source.n5 0.155672
R972 source.n48 source.n47 0.155672
R973 source.n47 source.n9 0.155672
R974 source.n39 source.n9 0.155672
R975 source.n39 source.n38 0.155672
R976 source.n38 source.n14 0.155672
R977 source.n31 source.n14 0.155672
R978 source.n31 source.n30 0.155672
R979 source.n30 source.n18 0.155672
R980 source.n23 source.n18 0.155672
R981 source.n137 source.n75 0.155672
R982 source.n130 source.n75 0.155672
R983 source.n130 source.n129 0.155672
R984 source.n129 source.n79 0.155672
R985 source.n122 source.n79 0.155672
R986 source.n122 source.n121 0.155672
R987 source.n121 source.n83 0.155672
R988 source.n113 source.n83 0.155672
R989 source.n113 source.n112 0.155672
R990 source.n112 source.n88 0.155672
R991 source.n105 source.n88 0.155672
R992 source.n105 source.n104 0.155672
R993 source.n104 source.n92 0.155672
R994 source.n97 source.n92 0.155672
R995 source.n203 source.n141 0.155672
R996 source.n196 source.n141 0.155672
R997 source.n196 source.n195 0.155672
R998 source.n195 source.n145 0.155672
R999 source.n188 source.n145 0.155672
R1000 source.n188 source.n187 0.155672
R1001 source.n187 source.n149 0.155672
R1002 source.n179 source.n149 0.155672
R1003 source.n179 source.n178 0.155672
R1004 source.n178 source.n154 0.155672
R1005 source.n171 source.n154 0.155672
R1006 source.n171 source.n170 0.155672
R1007 source.n170 source.n158 0.155672
R1008 source.n163 source.n158 0.155672
R1009 source.n277 source.n215 0.155672
R1010 source.n270 source.n215 0.155672
R1011 source.n270 source.n269 0.155672
R1012 source.n269 source.n219 0.155672
R1013 source.n262 source.n219 0.155672
R1014 source.n262 source.n261 0.155672
R1015 source.n261 source.n223 0.155672
R1016 source.n253 source.n223 0.155672
R1017 source.n253 source.n252 0.155672
R1018 source.n252 source.n228 0.155672
R1019 source.n245 source.n228 0.155672
R1020 source.n245 source.n244 0.155672
R1021 source.n244 source.n232 0.155672
R1022 source.n237 source.n232 0.155672
R1023 minus.n9 minus.t10 494.654
R1024 minus.n43 minus.t0 494.654
R1025 minus.n8 minus.t1 469.262
R1026 minus.n12 minus.t7 469.262
R1027 minus.n14 minus.t17 469.262
R1028 minus.n18 minus.t6 469.262
R1029 minus.n20 minus.t18 469.262
R1030 minus.n24 minus.t5 469.262
R1031 minus.n26 minus.t14 469.262
R1032 minus.n30 minus.t4 469.262
R1033 minus.n32 minus.t11 469.262
R1034 minus.n42 minus.t2 469.262
R1035 minus.n46 minus.t15 469.262
R1036 minus.n48 minus.t16 469.262
R1037 minus.n52 minus.t19 469.262
R1038 minus.n54 minus.t12 469.262
R1039 minus.n58 minus.t13 469.262
R1040 minus.n60 minus.t9 469.262
R1041 minus.n64 minus.t8 469.262
R1042 minus.n66 minus.t3 469.262
R1043 minus.n33 minus.n32 161.3
R1044 minus.n31 minus.n0 161.3
R1045 minus.n30 minus.n29 161.3
R1046 minus.n28 minus.n1 161.3
R1047 minus.n27 minus.n26 161.3
R1048 minus.n25 minus.n2 161.3
R1049 minus.n24 minus.n23 161.3
R1050 minus.n22 minus.n3 161.3
R1051 minus.n21 minus.n20 161.3
R1052 minus.n19 minus.n4 161.3
R1053 minus.n18 minus.n17 161.3
R1054 minus.n16 minus.n5 161.3
R1055 minus.n15 minus.n14 161.3
R1056 minus.n13 minus.n6 161.3
R1057 minus.n12 minus.n11 161.3
R1058 minus.n10 minus.n7 161.3
R1059 minus.n67 minus.n66 161.3
R1060 minus.n65 minus.n34 161.3
R1061 minus.n64 minus.n63 161.3
R1062 minus.n62 minus.n35 161.3
R1063 minus.n61 minus.n60 161.3
R1064 minus.n59 minus.n36 161.3
R1065 minus.n58 minus.n57 161.3
R1066 minus.n56 minus.n37 161.3
R1067 minus.n55 minus.n54 161.3
R1068 minus.n53 minus.n38 161.3
R1069 minus.n52 minus.n51 161.3
R1070 minus.n50 minus.n39 161.3
R1071 minus.n49 minus.n48 161.3
R1072 minus.n47 minus.n40 161.3
R1073 minus.n46 minus.n45 161.3
R1074 minus.n44 minus.n41 161.3
R1075 minus.n10 minus.n9 45.0031
R1076 minus.n44 minus.n43 45.0031
R1077 minus.n32 minus.n31 41.6278
R1078 minus.n66 minus.n65 41.6278
R1079 minus.n68 minus.n33 40.5838
R1080 minus.n8 minus.n7 37.246
R1081 minus.n30 minus.n1 37.246
R1082 minus.n42 minus.n41 37.246
R1083 minus.n64 minus.n35 37.246
R1084 minus.n13 minus.n12 32.8641
R1085 minus.n26 minus.n25 32.8641
R1086 minus.n47 minus.n46 32.8641
R1087 minus.n60 minus.n59 32.8641
R1088 minus.n14 minus.n5 28.4823
R1089 minus.n24 minus.n3 28.4823
R1090 minus.n48 minus.n39 28.4823
R1091 minus.n58 minus.n37 28.4823
R1092 minus.n20 minus.n19 24.1005
R1093 minus.n19 minus.n18 24.1005
R1094 minus.n53 minus.n52 24.1005
R1095 minus.n54 minus.n53 24.1005
R1096 minus.n18 minus.n5 19.7187
R1097 minus.n20 minus.n3 19.7187
R1098 minus.n52 minus.n39 19.7187
R1099 minus.n54 minus.n37 19.7187
R1100 minus.n9 minus.n8 15.6319
R1101 minus.n43 minus.n42 15.6319
R1102 minus.n14 minus.n13 15.3369
R1103 minus.n25 minus.n24 15.3369
R1104 minus.n48 minus.n47 15.3369
R1105 minus.n59 minus.n58 15.3369
R1106 minus.n12 minus.n7 10.955
R1107 minus.n26 minus.n1 10.955
R1108 minus.n46 minus.n41 10.955
R1109 minus.n60 minus.n35 10.955
R1110 minus.n68 minus.n67 6.66717
R1111 minus.n31 minus.n30 6.57323
R1112 minus.n65 minus.n64 6.57323
R1113 minus.n33 minus.n0 0.189894
R1114 minus.n29 minus.n0 0.189894
R1115 minus.n29 minus.n28 0.189894
R1116 minus.n28 minus.n27 0.189894
R1117 minus.n27 minus.n2 0.189894
R1118 minus.n23 minus.n2 0.189894
R1119 minus.n23 minus.n22 0.189894
R1120 minus.n22 minus.n21 0.189894
R1121 minus.n21 minus.n4 0.189894
R1122 minus.n17 minus.n4 0.189894
R1123 minus.n17 minus.n16 0.189894
R1124 minus.n16 minus.n15 0.189894
R1125 minus.n15 minus.n6 0.189894
R1126 minus.n11 minus.n6 0.189894
R1127 minus.n11 minus.n10 0.189894
R1128 minus.n45 minus.n44 0.189894
R1129 minus.n45 minus.n40 0.189894
R1130 minus.n49 minus.n40 0.189894
R1131 minus.n50 minus.n49 0.189894
R1132 minus.n51 minus.n50 0.189894
R1133 minus.n51 minus.n38 0.189894
R1134 minus.n55 minus.n38 0.189894
R1135 minus.n56 minus.n55 0.189894
R1136 minus.n57 minus.n56 0.189894
R1137 minus.n57 minus.n36 0.189894
R1138 minus.n61 minus.n36 0.189894
R1139 minus.n62 minus.n61 0.189894
R1140 minus.n63 minus.n62 0.189894
R1141 minus.n63 minus.n34 0.189894
R1142 minus.n67 minus.n34 0.189894
R1143 minus minus.n68 0.188
R1144 drain_right.n6 drain_right.n4 60.4404
R1145 drain_right.n2 drain_right.n0 60.4404
R1146 drain_right.n10 drain_right.n8 60.4404
R1147 drain_right.n10 drain_right.n9 59.5527
R1148 drain_right.n12 drain_right.n11 59.5527
R1149 drain_right.n14 drain_right.n13 59.5527
R1150 drain_right.n16 drain_right.n15 59.5527
R1151 drain_right.n7 drain_right.n3 59.5525
R1152 drain_right.n6 drain_right.n5 59.5525
R1153 drain_right.n2 drain_right.n1 59.5525
R1154 drain_right drain_right.n7 33.9173
R1155 drain_right drain_right.n16 6.54115
R1156 drain_right.n3 drain_right.t0 1.6505
R1157 drain_right.n3 drain_right.t7 1.6505
R1158 drain_right.n4 drain_right.t11 1.6505
R1159 drain_right.n4 drain_right.t16 1.6505
R1160 drain_right.n5 drain_right.t6 1.6505
R1161 drain_right.n5 drain_right.t10 1.6505
R1162 drain_right.n1 drain_right.t4 1.6505
R1163 drain_right.n1 drain_right.t3 1.6505
R1164 drain_right.n0 drain_right.t19 1.6505
R1165 drain_right.n0 drain_right.t17 1.6505
R1166 drain_right.n8 drain_right.t18 1.6505
R1167 drain_right.n8 drain_right.t9 1.6505
R1168 drain_right.n9 drain_right.t2 1.6505
R1169 drain_right.n9 drain_right.t12 1.6505
R1170 drain_right.n11 drain_right.t1 1.6505
R1171 drain_right.n11 drain_right.t13 1.6505
R1172 drain_right.n13 drain_right.t5 1.6505
R1173 drain_right.n13 drain_right.t14 1.6505
R1174 drain_right.n15 drain_right.t8 1.6505
R1175 drain_right.n15 drain_right.t15 1.6505
R1176 drain_right.n16 drain_right.n14 0.888431
R1177 drain_right.n14 drain_right.n12 0.888431
R1178 drain_right.n12 drain_right.n10 0.888431
R1179 drain_right.n7 drain_right.n6 0.833085
R1180 drain_right.n7 drain_right.n2 0.833085
C0 drain_left minus 0.173554f
C1 minus plus 6.86553f
C2 source drain_right 24.0697f
C3 source drain_left 24.0673f
C4 source plus 12.7614f
C5 drain_left drain_right 1.59885f
C6 source minus 12.7474f
C7 drain_right plus 0.454687f
C8 drain_left plus 12.8881f
C9 drain_right minus 12.590599f
C10 drain_right a_n2982_n3288# 7.33447f
C11 drain_left a_n2982_n3288# 7.75292f
C12 source a_n2982_n3288# 9.423556f
C13 minus a_n2982_n3288# 12.001272f
C14 plus a_n2982_n3288# 13.82572f
C15 drain_right.t19 a_n2982_n3288# 0.257766f
C16 drain_right.t17 a_n2982_n3288# 0.257766f
C17 drain_right.n0 a_n2982_n3288# 2.29952f
C18 drain_right.t4 a_n2982_n3288# 0.257766f
C19 drain_right.t3 a_n2982_n3288# 0.257766f
C20 drain_right.n1 a_n2982_n3288# 2.29372f
C21 drain_right.n2 a_n2982_n3288# 0.768413f
C22 drain_right.t0 a_n2982_n3288# 0.257766f
C23 drain_right.t7 a_n2982_n3288# 0.257766f
C24 drain_right.n3 a_n2982_n3288# 2.29372f
C25 drain_right.t11 a_n2982_n3288# 0.257766f
C26 drain_right.t16 a_n2982_n3288# 0.257766f
C27 drain_right.n4 a_n2982_n3288# 2.29952f
C28 drain_right.t6 a_n2982_n3288# 0.257766f
C29 drain_right.t10 a_n2982_n3288# 0.257766f
C30 drain_right.n5 a_n2982_n3288# 2.29372f
C31 drain_right.n6 a_n2982_n3288# 0.768413f
C32 drain_right.n7 a_n2982_n3288# 1.92967f
C33 drain_right.t18 a_n2982_n3288# 0.257766f
C34 drain_right.t9 a_n2982_n3288# 0.257766f
C35 drain_right.n8 a_n2982_n3288# 2.29952f
C36 drain_right.t2 a_n2982_n3288# 0.257766f
C37 drain_right.t12 a_n2982_n3288# 0.257766f
C38 drain_right.n9 a_n2982_n3288# 2.29373f
C39 drain_right.n10 a_n2982_n3288# 0.772494f
C40 drain_right.t1 a_n2982_n3288# 0.257766f
C41 drain_right.t13 a_n2982_n3288# 0.257766f
C42 drain_right.n11 a_n2982_n3288# 2.29373f
C43 drain_right.n12 a_n2982_n3288# 0.383667f
C44 drain_right.t5 a_n2982_n3288# 0.257766f
C45 drain_right.t14 a_n2982_n3288# 0.257766f
C46 drain_right.n13 a_n2982_n3288# 2.29373f
C47 drain_right.n14 a_n2982_n3288# 0.383667f
C48 drain_right.t8 a_n2982_n3288# 0.257766f
C49 drain_right.t15 a_n2982_n3288# 0.257766f
C50 drain_right.n15 a_n2982_n3288# 2.29373f
C51 drain_right.n16 a_n2982_n3288# 0.624098f
C52 minus.n0 a_n2982_n3288# 0.039702f
C53 minus.n1 a_n2982_n3288# 0.009009f
C54 minus.t4 a_n2982_n3288# 0.950976f
C55 minus.n2 a_n2982_n3288# 0.039702f
C56 minus.n3 a_n2982_n3288# 0.009009f
C57 minus.t5 a_n2982_n3288# 0.950976f
C58 minus.n4 a_n2982_n3288# 0.039702f
C59 minus.n5 a_n2982_n3288# 0.009009f
C60 minus.t6 a_n2982_n3288# 0.950976f
C61 minus.n6 a_n2982_n3288# 0.039702f
C62 minus.n7 a_n2982_n3288# 0.009009f
C63 minus.t7 a_n2982_n3288# 0.950976f
C64 minus.t10 a_n2982_n3288# 0.970467f
C65 minus.t1 a_n2982_n3288# 0.950976f
C66 minus.n8 a_n2982_n3288# 0.385908f
C67 minus.n9 a_n2982_n3288# 0.362627f
C68 minus.n10 a_n2982_n3288# 0.169465f
C69 minus.n11 a_n2982_n3288# 0.039702f
C70 minus.n12 a_n2982_n3288# 0.379267f
C71 minus.n13 a_n2982_n3288# 0.009009f
C72 minus.t17 a_n2982_n3288# 0.950976f
C73 minus.n14 a_n2982_n3288# 0.379267f
C74 minus.n15 a_n2982_n3288# 0.039702f
C75 minus.n16 a_n2982_n3288# 0.039702f
C76 minus.n17 a_n2982_n3288# 0.039702f
C77 minus.n18 a_n2982_n3288# 0.379267f
C78 minus.n19 a_n2982_n3288# 0.009009f
C79 minus.t18 a_n2982_n3288# 0.950976f
C80 minus.n20 a_n2982_n3288# 0.379267f
C81 minus.n21 a_n2982_n3288# 0.039702f
C82 minus.n22 a_n2982_n3288# 0.039702f
C83 minus.n23 a_n2982_n3288# 0.039702f
C84 minus.n24 a_n2982_n3288# 0.379267f
C85 minus.n25 a_n2982_n3288# 0.009009f
C86 minus.t14 a_n2982_n3288# 0.950976f
C87 minus.n26 a_n2982_n3288# 0.379267f
C88 minus.n27 a_n2982_n3288# 0.039702f
C89 minus.n28 a_n2982_n3288# 0.039702f
C90 minus.n29 a_n2982_n3288# 0.039702f
C91 minus.n30 a_n2982_n3288# 0.379267f
C92 minus.n31 a_n2982_n3288# 0.009009f
C93 minus.t11 a_n2982_n3288# 0.950976f
C94 minus.n32 a_n2982_n3288# 0.3789f
C95 minus.n33 a_n2982_n3288# 1.67569f
C96 minus.n34 a_n2982_n3288# 0.039702f
C97 minus.n35 a_n2982_n3288# 0.009009f
C98 minus.n36 a_n2982_n3288# 0.039702f
C99 minus.n37 a_n2982_n3288# 0.009009f
C100 minus.n38 a_n2982_n3288# 0.039702f
C101 minus.n39 a_n2982_n3288# 0.009009f
C102 minus.n40 a_n2982_n3288# 0.039702f
C103 minus.n41 a_n2982_n3288# 0.009009f
C104 minus.t0 a_n2982_n3288# 0.970467f
C105 minus.t2 a_n2982_n3288# 0.950976f
C106 minus.n42 a_n2982_n3288# 0.385908f
C107 minus.n43 a_n2982_n3288# 0.362627f
C108 minus.n44 a_n2982_n3288# 0.169465f
C109 minus.n45 a_n2982_n3288# 0.039702f
C110 minus.t15 a_n2982_n3288# 0.950976f
C111 minus.n46 a_n2982_n3288# 0.379267f
C112 minus.n47 a_n2982_n3288# 0.009009f
C113 minus.t16 a_n2982_n3288# 0.950976f
C114 minus.n48 a_n2982_n3288# 0.379267f
C115 minus.n49 a_n2982_n3288# 0.039702f
C116 minus.n50 a_n2982_n3288# 0.039702f
C117 minus.n51 a_n2982_n3288# 0.039702f
C118 minus.t19 a_n2982_n3288# 0.950976f
C119 minus.n52 a_n2982_n3288# 0.379267f
C120 minus.n53 a_n2982_n3288# 0.009009f
C121 minus.t12 a_n2982_n3288# 0.950976f
C122 minus.n54 a_n2982_n3288# 0.379267f
C123 minus.n55 a_n2982_n3288# 0.039702f
C124 minus.n56 a_n2982_n3288# 0.039702f
C125 minus.n57 a_n2982_n3288# 0.039702f
C126 minus.t13 a_n2982_n3288# 0.950976f
C127 minus.n58 a_n2982_n3288# 0.379267f
C128 minus.n59 a_n2982_n3288# 0.009009f
C129 minus.t9 a_n2982_n3288# 0.950976f
C130 minus.n60 a_n2982_n3288# 0.379267f
C131 minus.n61 a_n2982_n3288# 0.039702f
C132 minus.n62 a_n2982_n3288# 0.039702f
C133 minus.n63 a_n2982_n3288# 0.039702f
C134 minus.t8 a_n2982_n3288# 0.950976f
C135 minus.n64 a_n2982_n3288# 0.379267f
C136 minus.n65 a_n2982_n3288# 0.009009f
C137 minus.t3 a_n2982_n3288# 0.950976f
C138 minus.n66 a_n2982_n3288# 0.3789f
C139 minus.n67 a_n2982_n3288# 0.275078f
C140 minus.n68 a_n2982_n3288# 2.00531f
C141 source.n0 a_n2982_n3288# 0.032056f
C142 source.n1 a_n2982_n3288# 0.0242f
C143 source.n2 a_n2982_n3288# 0.013004f
C144 source.n3 a_n2982_n3288# 0.030737f
C145 source.n4 a_n2982_n3288# 0.013769f
C146 source.n5 a_n2982_n3288# 0.0242f
C147 source.n6 a_n2982_n3288# 0.013004f
C148 source.n7 a_n2982_n3288# 0.030737f
C149 source.n8 a_n2982_n3288# 0.013769f
C150 source.n9 a_n2982_n3288# 0.0242f
C151 source.n10 a_n2982_n3288# 0.013386f
C152 source.n11 a_n2982_n3288# 0.030737f
C153 source.n12 a_n2982_n3288# 0.013004f
C154 source.n13 a_n2982_n3288# 0.013769f
C155 source.n14 a_n2982_n3288# 0.0242f
C156 source.n15 a_n2982_n3288# 0.013004f
C157 source.n16 a_n2982_n3288# 0.030737f
C158 source.n17 a_n2982_n3288# 0.013769f
C159 source.n18 a_n2982_n3288# 0.0242f
C160 source.n19 a_n2982_n3288# 0.013004f
C161 source.n20 a_n2982_n3288# 0.023052f
C162 source.n21 a_n2982_n3288# 0.021728f
C163 source.t34 a_n2982_n3288# 0.051912f
C164 source.n22 a_n2982_n3288# 0.174478f
C165 source.n23 a_n2982_n3288# 1.22084f
C166 source.n24 a_n2982_n3288# 0.013004f
C167 source.n25 a_n2982_n3288# 0.013769f
C168 source.n26 a_n2982_n3288# 0.030737f
C169 source.n27 a_n2982_n3288# 0.030737f
C170 source.n28 a_n2982_n3288# 0.013769f
C171 source.n29 a_n2982_n3288# 0.013004f
C172 source.n30 a_n2982_n3288# 0.0242f
C173 source.n31 a_n2982_n3288# 0.0242f
C174 source.n32 a_n2982_n3288# 0.013004f
C175 source.n33 a_n2982_n3288# 0.013769f
C176 source.n34 a_n2982_n3288# 0.030737f
C177 source.n35 a_n2982_n3288# 0.030737f
C178 source.n36 a_n2982_n3288# 0.013769f
C179 source.n37 a_n2982_n3288# 0.013004f
C180 source.n38 a_n2982_n3288# 0.0242f
C181 source.n39 a_n2982_n3288# 0.0242f
C182 source.n40 a_n2982_n3288# 0.013004f
C183 source.n41 a_n2982_n3288# 0.013769f
C184 source.n42 a_n2982_n3288# 0.030737f
C185 source.n43 a_n2982_n3288# 0.030737f
C186 source.n44 a_n2982_n3288# 0.030737f
C187 source.n45 a_n2982_n3288# 0.013386f
C188 source.n46 a_n2982_n3288# 0.013004f
C189 source.n47 a_n2982_n3288# 0.0242f
C190 source.n48 a_n2982_n3288# 0.0242f
C191 source.n49 a_n2982_n3288# 0.013004f
C192 source.n50 a_n2982_n3288# 0.013769f
C193 source.n51 a_n2982_n3288# 0.030737f
C194 source.n52 a_n2982_n3288# 0.030737f
C195 source.n53 a_n2982_n3288# 0.013769f
C196 source.n54 a_n2982_n3288# 0.013004f
C197 source.n55 a_n2982_n3288# 0.0242f
C198 source.n56 a_n2982_n3288# 0.0242f
C199 source.n57 a_n2982_n3288# 0.013004f
C200 source.n58 a_n2982_n3288# 0.013769f
C201 source.n59 a_n2982_n3288# 0.030737f
C202 source.n60 a_n2982_n3288# 0.063075f
C203 source.n61 a_n2982_n3288# 0.013769f
C204 source.n62 a_n2982_n3288# 0.013004f
C205 source.n63 a_n2982_n3288# 0.05197f
C206 source.n64 a_n2982_n3288# 0.03481f
C207 source.n65 a_n2982_n3288# 1.018f
C208 source.t29 a_n2982_n3288# 0.229481f
C209 source.t19 a_n2982_n3288# 0.229481f
C210 source.n66 a_n2982_n3288# 1.96482f
C211 source.n67 a_n2982_n3288# 0.385889f
C212 source.t27 a_n2982_n3288# 0.229481f
C213 source.t36 a_n2982_n3288# 0.229481f
C214 source.n68 a_n2982_n3288# 1.96482f
C215 source.n69 a_n2982_n3288# 0.385889f
C216 source.t28 a_n2982_n3288# 0.229481f
C217 source.t33 a_n2982_n3288# 0.229481f
C218 source.n70 a_n2982_n3288# 1.96482f
C219 source.n71 a_n2982_n3288# 0.385889f
C220 source.t24 a_n2982_n3288# 0.229481f
C221 source.t35 a_n2982_n3288# 0.229481f
C222 source.n72 a_n2982_n3288# 1.96482f
C223 source.n73 a_n2982_n3288# 0.385889f
C224 source.n74 a_n2982_n3288# 0.032056f
C225 source.n75 a_n2982_n3288# 0.0242f
C226 source.n76 a_n2982_n3288# 0.013004f
C227 source.n77 a_n2982_n3288# 0.030737f
C228 source.n78 a_n2982_n3288# 0.013769f
C229 source.n79 a_n2982_n3288# 0.0242f
C230 source.n80 a_n2982_n3288# 0.013004f
C231 source.n81 a_n2982_n3288# 0.030737f
C232 source.n82 a_n2982_n3288# 0.013769f
C233 source.n83 a_n2982_n3288# 0.0242f
C234 source.n84 a_n2982_n3288# 0.013386f
C235 source.n85 a_n2982_n3288# 0.030737f
C236 source.n86 a_n2982_n3288# 0.013004f
C237 source.n87 a_n2982_n3288# 0.013769f
C238 source.n88 a_n2982_n3288# 0.0242f
C239 source.n89 a_n2982_n3288# 0.013004f
C240 source.n90 a_n2982_n3288# 0.030737f
C241 source.n91 a_n2982_n3288# 0.013769f
C242 source.n92 a_n2982_n3288# 0.0242f
C243 source.n93 a_n2982_n3288# 0.013004f
C244 source.n94 a_n2982_n3288# 0.023052f
C245 source.n95 a_n2982_n3288# 0.021728f
C246 source.t32 a_n2982_n3288# 0.051912f
C247 source.n96 a_n2982_n3288# 0.174478f
C248 source.n97 a_n2982_n3288# 1.22084f
C249 source.n98 a_n2982_n3288# 0.013004f
C250 source.n99 a_n2982_n3288# 0.013769f
C251 source.n100 a_n2982_n3288# 0.030737f
C252 source.n101 a_n2982_n3288# 0.030737f
C253 source.n102 a_n2982_n3288# 0.013769f
C254 source.n103 a_n2982_n3288# 0.013004f
C255 source.n104 a_n2982_n3288# 0.0242f
C256 source.n105 a_n2982_n3288# 0.0242f
C257 source.n106 a_n2982_n3288# 0.013004f
C258 source.n107 a_n2982_n3288# 0.013769f
C259 source.n108 a_n2982_n3288# 0.030737f
C260 source.n109 a_n2982_n3288# 0.030737f
C261 source.n110 a_n2982_n3288# 0.013769f
C262 source.n111 a_n2982_n3288# 0.013004f
C263 source.n112 a_n2982_n3288# 0.0242f
C264 source.n113 a_n2982_n3288# 0.0242f
C265 source.n114 a_n2982_n3288# 0.013004f
C266 source.n115 a_n2982_n3288# 0.013769f
C267 source.n116 a_n2982_n3288# 0.030737f
C268 source.n117 a_n2982_n3288# 0.030737f
C269 source.n118 a_n2982_n3288# 0.030737f
C270 source.n119 a_n2982_n3288# 0.013386f
C271 source.n120 a_n2982_n3288# 0.013004f
C272 source.n121 a_n2982_n3288# 0.0242f
C273 source.n122 a_n2982_n3288# 0.0242f
C274 source.n123 a_n2982_n3288# 0.013004f
C275 source.n124 a_n2982_n3288# 0.013769f
C276 source.n125 a_n2982_n3288# 0.030737f
C277 source.n126 a_n2982_n3288# 0.030737f
C278 source.n127 a_n2982_n3288# 0.013769f
C279 source.n128 a_n2982_n3288# 0.013004f
C280 source.n129 a_n2982_n3288# 0.0242f
C281 source.n130 a_n2982_n3288# 0.0242f
C282 source.n131 a_n2982_n3288# 0.013004f
C283 source.n132 a_n2982_n3288# 0.013769f
C284 source.n133 a_n2982_n3288# 0.030737f
C285 source.n134 a_n2982_n3288# 0.063075f
C286 source.n135 a_n2982_n3288# 0.013769f
C287 source.n136 a_n2982_n3288# 0.013004f
C288 source.n137 a_n2982_n3288# 0.05197f
C289 source.n138 a_n2982_n3288# 0.03481f
C290 source.n139 a_n2982_n3288# 0.124308f
C291 source.n140 a_n2982_n3288# 0.032056f
C292 source.n141 a_n2982_n3288# 0.0242f
C293 source.n142 a_n2982_n3288# 0.013004f
C294 source.n143 a_n2982_n3288# 0.030737f
C295 source.n144 a_n2982_n3288# 0.013769f
C296 source.n145 a_n2982_n3288# 0.0242f
C297 source.n146 a_n2982_n3288# 0.013004f
C298 source.n147 a_n2982_n3288# 0.030737f
C299 source.n148 a_n2982_n3288# 0.013769f
C300 source.n149 a_n2982_n3288# 0.0242f
C301 source.n150 a_n2982_n3288# 0.013386f
C302 source.n151 a_n2982_n3288# 0.030737f
C303 source.n152 a_n2982_n3288# 0.013004f
C304 source.n153 a_n2982_n3288# 0.013769f
C305 source.n154 a_n2982_n3288# 0.0242f
C306 source.n155 a_n2982_n3288# 0.013004f
C307 source.n156 a_n2982_n3288# 0.030737f
C308 source.n157 a_n2982_n3288# 0.013769f
C309 source.n158 a_n2982_n3288# 0.0242f
C310 source.n159 a_n2982_n3288# 0.013004f
C311 source.n160 a_n2982_n3288# 0.023052f
C312 source.n161 a_n2982_n3288# 0.021728f
C313 source.t6 a_n2982_n3288# 0.051912f
C314 source.n162 a_n2982_n3288# 0.174478f
C315 source.n163 a_n2982_n3288# 1.22084f
C316 source.n164 a_n2982_n3288# 0.013004f
C317 source.n165 a_n2982_n3288# 0.013769f
C318 source.n166 a_n2982_n3288# 0.030737f
C319 source.n167 a_n2982_n3288# 0.030737f
C320 source.n168 a_n2982_n3288# 0.013769f
C321 source.n169 a_n2982_n3288# 0.013004f
C322 source.n170 a_n2982_n3288# 0.0242f
C323 source.n171 a_n2982_n3288# 0.0242f
C324 source.n172 a_n2982_n3288# 0.013004f
C325 source.n173 a_n2982_n3288# 0.013769f
C326 source.n174 a_n2982_n3288# 0.030737f
C327 source.n175 a_n2982_n3288# 0.030737f
C328 source.n176 a_n2982_n3288# 0.013769f
C329 source.n177 a_n2982_n3288# 0.013004f
C330 source.n178 a_n2982_n3288# 0.0242f
C331 source.n179 a_n2982_n3288# 0.0242f
C332 source.n180 a_n2982_n3288# 0.013004f
C333 source.n181 a_n2982_n3288# 0.013769f
C334 source.n182 a_n2982_n3288# 0.030737f
C335 source.n183 a_n2982_n3288# 0.030737f
C336 source.n184 a_n2982_n3288# 0.030737f
C337 source.n185 a_n2982_n3288# 0.013386f
C338 source.n186 a_n2982_n3288# 0.013004f
C339 source.n187 a_n2982_n3288# 0.0242f
C340 source.n188 a_n2982_n3288# 0.0242f
C341 source.n189 a_n2982_n3288# 0.013004f
C342 source.n190 a_n2982_n3288# 0.013769f
C343 source.n191 a_n2982_n3288# 0.030737f
C344 source.n192 a_n2982_n3288# 0.030737f
C345 source.n193 a_n2982_n3288# 0.013769f
C346 source.n194 a_n2982_n3288# 0.013004f
C347 source.n195 a_n2982_n3288# 0.0242f
C348 source.n196 a_n2982_n3288# 0.0242f
C349 source.n197 a_n2982_n3288# 0.013004f
C350 source.n198 a_n2982_n3288# 0.013769f
C351 source.n199 a_n2982_n3288# 0.030737f
C352 source.n200 a_n2982_n3288# 0.063075f
C353 source.n201 a_n2982_n3288# 0.013769f
C354 source.n202 a_n2982_n3288# 0.013004f
C355 source.n203 a_n2982_n3288# 0.05197f
C356 source.n204 a_n2982_n3288# 0.03481f
C357 source.n205 a_n2982_n3288# 0.124308f
C358 source.t8 a_n2982_n3288# 0.229481f
C359 source.t11 a_n2982_n3288# 0.229481f
C360 source.n206 a_n2982_n3288# 1.96482f
C361 source.n207 a_n2982_n3288# 0.385889f
C362 source.t10 a_n2982_n3288# 0.229481f
C363 source.t16 a_n2982_n3288# 0.229481f
C364 source.n208 a_n2982_n3288# 1.96482f
C365 source.n209 a_n2982_n3288# 0.385889f
C366 source.t5 a_n2982_n3288# 0.229481f
C367 source.t2 a_n2982_n3288# 0.229481f
C368 source.n210 a_n2982_n3288# 1.96482f
C369 source.n211 a_n2982_n3288# 0.385889f
C370 source.t1 a_n2982_n3288# 0.229481f
C371 source.t13 a_n2982_n3288# 0.229481f
C372 source.n212 a_n2982_n3288# 1.96482f
C373 source.n213 a_n2982_n3288# 0.385889f
C374 source.n214 a_n2982_n3288# 0.032056f
C375 source.n215 a_n2982_n3288# 0.0242f
C376 source.n216 a_n2982_n3288# 0.013004f
C377 source.n217 a_n2982_n3288# 0.030737f
C378 source.n218 a_n2982_n3288# 0.013769f
C379 source.n219 a_n2982_n3288# 0.0242f
C380 source.n220 a_n2982_n3288# 0.013004f
C381 source.n221 a_n2982_n3288# 0.030737f
C382 source.n222 a_n2982_n3288# 0.013769f
C383 source.n223 a_n2982_n3288# 0.0242f
C384 source.n224 a_n2982_n3288# 0.013386f
C385 source.n225 a_n2982_n3288# 0.030737f
C386 source.n226 a_n2982_n3288# 0.013004f
C387 source.n227 a_n2982_n3288# 0.013769f
C388 source.n228 a_n2982_n3288# 0.0242f
C389 source.n229 a_n2982_n3288# 0.013004f
C390 source.n230 a_n2982_n3288# 0.030737f
C391 source.n231 a_n2982_n3288# 0.013769f
C392 source.n232 a_n2982_n3288# 0.0242f
C393 source.n233 a_n2982_n3288# 0.013004f
C394 source.n234 a_n2982_n3288# 0.023052f
C395 source.n235 a_n2982_n3288# 0.021728f
C396 source.t12 a_n2982_n3288# 0.051912f
C397 source.n236 a_n2982_n3288# 0.174478f
C398 source.n237 a_n2982_n3288# 1.22084f
C399 source.n238 a_n2982_n3288# 0.013004f
C400 source.n239 a_n2982_n3288# 0.013769f
C401 source.n240 a_n2982_n3288# 0.030737f
C402 source.n241 a_n2982_n3288# 0.030737f
C403 source.n242 a_n2982_n3288# 0.013769f
C404 source.n243 a_n2982_n3288# 0.013004f
C405 source.n244 a_n2982_n3288# 0.0242f
C406 source.n245 a_n2982_n3288# 0.0242f
C407 source.n246 a_n2982_n3288# 0.013004f
C408 source.n247 a_n2982_n3288# 0.013769f
C409 source.n248 a_n2982_n3288# 0.030737f
C410 source.n249 a_n2982_n3288# 0.030737f
C411 source.n250 a_n2982_n3288# 0.013769f
C412 source.n251 a_n2982_n3288# 0.013004f
C413 source.n252 a_n2982_n3288# 0.0242f
C414 source.n253 a_n2982_n3288# 0.0242f
C415 source.n254 a_n2982_n3288# 0.013004f
C416 source.n255 a_n2982_n3288# 0.013769f
C417 source.n256 a_n2982_n3288# 0.030737f
C418 source.n257 a_n2982_n3288# 0.030737f
C419 source.n258 a_n2982_n3288# 0.030737f
C420 source.n259 a_n2982_n3288# 0.013386f
C421 source.n260 a_n2982_n3288# 0.013004f
C422 source.n261 a_n2982_n3288# 0.0242f
C423 source.n262 a_n2982_n3288# 0.0242f
C424 source.n263 a_n2982_n3288# 0.013004f
C425 source.n264 a_n2982_n3288# 0.013769f
C426 source.n265 a_n2982_n3288# 0.030737f
C427 source.n266 a_n2982_n3288# 0.030737f
C428 source.n267 a_n2982_n3288# 0.013769f
C429 source.n268 a_n2982_n3288# 0.013004f
C430 source.n269 a_n2982_n3288# 0.0242f
C431 source.n270 a_n2982_n3288# 0.0242f
C432 source.n271 a_n2982_n3288# 0.013004f
C433 source.n272 a_n2982_n3288# 0.013769f
C434 source.n273 a_n2982_n3288# 0.030737f
C435 source.n274 a_n2982_n3288# 0.063075f
C436 source.n275 a_n2982_n3288# 0.013769f
C437 source.n276 a_n2982_n3288# 0.013004f
C438 source.n277 a_n2982_n3288# 0.05197f
C439 source.n278 a_n2982_n3288# 0.03481f
C440 source.n279 a_n2982_n3288# 1.40822f
C441 source.n280 a_n2982_n3288# 0.032056f
C442 source.n281 a_n2982_n3288# 0.0242f
C443 source.n282 a_n2982_n3288# 0.013004f
C444 source.n283 a_n2982_n3288# 0.030737f
C445 source.n284 a_n2982_n3288# 0.013769f
C446 source.n285 a_n2982_n3288# 0.0242f
C447 source.n286 a_n2982_n3288# 0.013004f
C448 source.n287 a_n2982_n3288# 0.030737f
C449 source.n288 a_n2982_n3288# 0.013769f
C450 source.n289 a_n2982_n3288# 0.0242f
C451 source.n290 a_n2982_n3288# 0.013386f
C452 source.n291 a_n2982_n3288# 0.030737f
C453 source.n292 a_n2982_n3288# 0.013769f
C454 source.n293 a_n2982_n3288# 0.0242f
C455 source.n294 a_n2982_n3288# 0.013004f
C456 source.n295 a_n2982_n3288# 0.030737f
C457 source.n296 a_n2982_n3288# 0.013769f
C458 source.n297 a_n2982_n3288# 0.0242f
C459 source.n298 a_n2982_n3288# 0.013004f
C460 source.n299 a_n2982_n3288# 0.023052f
C461 source.n300 a_n2982_n3288# 0.021728f
C462 source.t25 a_n2982_n3288# 0.051912f
C463 source.n301 a_n2982_n3288# 0.174478f
C464 source.n302 a_n2982_n3288# 1.22084f
C465 source.n303 a_n2982_n3288# 0.013004f
C466 source.n304 a_n2982_n3288# 0.013769f
C467 source.n305 a_n2982_n3288# 0.030737f
C468 source.n306 a_n2982_n3288# 0.030737f
C469 source.n307 a_n2982_n3288# 0.013769f
C470 source.n308 a_n2982_n3288# 0.013004f
C471 source.n309 a_n2982_n3288# 0.0242f
C472 source.n310 a_n2982_n3288# 0.0242f
C473 source.n311 a_n2982_n3288# 0.013004f
C474 source.n312 a_n2982_n3288# 0.013769f
C475 source.n313 a_n2982_n3288# 0.030737f
C476 source.n314 a_n2982_n3288# 0.030737f
C477 source.n315 a_n2982_n3288# 0.013769f
C478 source.n316 a_n2982_n3288# 0.013004f
C479 source.n317 a_n2982_n3288# 0.0242f
C480 source.n318 a_n2982_n3288# 0.0242f
C481 source.n319 a_n2982_n3288# 0.013004f
C482 source.n320 a_n2982_n3288# 0.013004f
C483 source.n321 a_n2982_n3288# 0.013769f
C484 source.n322 a_n2982_n3288# 0.030737f
C485 source.n323 a_n2982_n3288# 0.030737f
C486 source.n324 a_n2982_n3288# 0.030737f
C487 source.n325 a_n2982_n3288# 0.013386f
C488 source.n326 a_n2982_n3288# 0.013004f
C489 source.n327 a_n2982_n3288# 0.0242f
C490 source.n328 a_n2982_n3288# 0.0242f
C491 source.n329 a_n2982_n3288# 0.013004f
C492 source.n330 a_n2982_n3288# 0.013769f
C493 source.n331 a_n2982_n3288# 0.030737f
C494 source.n332 a_n2982_n3288# 0.030737f
C495 source.n333 a_n2982_n3288# 0.013769f
C496 source.n334 a_n2982_n3288# 0.013004f
C497 source.n335 a_n2982_n3288# 0.0242f
C498 source.n336 a_n2982_n3288# 0.0242f
C499 source.n337 a_n2982_n3288# 0.013004f
C500 source.n338 a_n2982_n3288# 0.013769f
C501 source.n339 a_n2982_n3288# 0.030737f
C502 source.n340 a_n2982_n3288# 0.063075f
C503 source.n341 a_n2982_n3288# 0.013769f
C504 source.n342 a_n2982_n3288# 0.013004f
C505 source.n343 a_n2982_n3288# 0.05197f
C506 source.n344 a_n2982_n3288# 0.03481f
C507 source.n345 a_n2982_n3288# 1.40822f
C508 source.t26 a_n2982_n3288# 0.229481f
C509 source.t22 a_n2982_n3288# 0.229481f
C510 source.n346 a_n2982_n3288# 1.96481f
C511 source.n347 a_n2982_n3288# 0.385901f
C512 source.t37 a_n2982_n3288# 0.229481f
C513 source.t38 a_n2982_n3288# 0.229481f
C514 source.n348 a_n2982_n3288# 1.96481f
C515 source.n349 a_n2982_n3288# 0.385901f
C516 source.t30 a_n2982_n3288# 0.229481f
C517 source.t31 a_n2982_n3288# 0.229481f
C518 source.n350 a_n2982_n3288# 1.96481f
C519 source.n351 a_n2982_n3288# 0.385901f
C520 source.t23 a_n2982_n3288# 0.229481f
C521 source.t20 a_n2982_n3288# 0.229481f
C522 source.n352 a_n2982_n3288# 1.96481f
C523 source.n353 a_n2982_n3288# 0.385901f
C524 source.n354 a_n2982_n3288# 0.032056f
C525 source.n355 a_n2982_n3288# 0.0242f
C526 source.n356 a_n2982_n3288# 0.013004f
C527 source.n357 a_n2982_n3288# 0.030737f
C528 source.n358 a_n2982_n3288# 0.013769f
C529 source.n359 a_n2982_n3288# 0.0242f
C530 source.n360 a_n2982_n3288# 0.013004f
C531 source.n361 a_n2982_n3288# 0.030737f
C532 source.n362 a_n2982_n3288# 0.013769f
C533 source.n363 a_n2982_n3288# 0.0242f
C534 source.n364 a_n2982_n3288# 0.013386f
C535 source.n365 a_n2982_n3288# 0.030737f
C536 source.n366 a_n2982_n3288# 0.013769f
C537 source.n367 a_n2982_n3288# 0.0242f
C538 source.n368 a_n2982_n3288# 0.013004f
C539 source.n369 a_n2982_n3288# 0.030737f
C540 source.n370 a_n2982_n3288# 0.013769f
C541 source.n371 a_n2982_n3288# 0.0242f
C542 source.n372 a_n2982_n3288# 0.013004f
C543 source.n373 a_n2982_n3288# 0.023052f
C544 source.n374 a_n2982_n3288# 0.021728f
C545 source.t21 a_n2982_n3288# 0.051912f
C546 source.n375 a_n2982_n3288# 0.174478f
C547 source.n376 a_n2982_n3288# 1.22084f
C548 source.n377 a_n2982_n3288# 0.013004f
C549 source.n378 a_n2982_n3288# 0.013769f
C550 source.n379 a_n2982_n3288# 0.030737f
C551 source.n380 a_n2982_n3288# 0.030737f
C552 source.n381 a_n2982_n3288# 0.013769f
C553 source.n382 a_n2982_n3288# 0.013004f
C554 source.n383 a_n2982_n3288# 0.0242f
C555 source.n384 a_n2982_n3288# 0.0242f
C556 source.n385 a_n2982_n3288# 0.013004f
C557 source.n386 a_n2982_n3288# 0.013769f
C558 source.n387 a_n2982_n3288# 0.030737f
C559 source.n388 a_n2982_n3288# 0.030737f
C560 source.n389 a_n2982_n3288# 0.013769f
C561 source.n390 a_n2982_n3288# 0.013004f
C562 source.n391 a_n2982_n3288# 0.0242f
C563 source.n392 a_n2982_n3288# 0.0242f
C564 source.n393 a_n2982_n3288# 0.013004f
C565 source.n394 a_n2982_n3288# 0.013004f
C566 source.n395 a_n2982_n3288# 0.013769f
C567 source.n396 a_n2982_n3288# 0.030737f
C568 source.n397 a_n2982_n3288# 0.030737f
C569 source.n398 a_n2982_n3288# 0.030737f
C570 source.n399 a_n2982_n3288# 0.013386f
C571 source.n400 a_n2982_n3288# 0.013004f
C572 source.n401 a_n2982_n3288# 0.0242f
C573 source.n402 a_n2982_n3288# 0.0242f
C574 source.n403 a_n2982_n3288# 0.013004f
C575 source.n404 a_n2982_n3288# 0.013769f
C576 source.n405 a_n2982_n3288# 0.030737f
C577 source.n406 a_n2982_n3288# 0.030737f
C578 source.n407 a_n2982_n3288# 0.013769f
C579 source.n408 a_n2982_n3288# 0.013004f
C580 source.n409 a_n2982_n3288# 0.0242f
C581 source.n410 a_n2982_n3288# 0.0242f
C582 source.n411 a_n2982_n3288# 0.013004f
C583 source.n412 a_n2982_n3288# 0.013769f
C584 source.n413 a_n2982_n3288# 0.030737f
C585 source.n414 a_n2982_n3288# 0.063075f
C586 source.n415 a_n2982_n3288# 0.013769f
C587 source.n416 a_n2982_n3288# 0.013004f
C588 source.n417 a_n2982_n3288# 0.05197f
C589 source.n418 a_n2982_n3288# 0.03481f
C590 source.n419 a_n2982_n3288# 0.124308f
C591 source.n420 a_n2982_n3288# 0.032056f
C592 source.n421 a_n2982_n3288# 0.0242f
C593 source.n422 a_n2982_n3288# 0.013004f
C594 source.n423 a_n2982_n3288# 0.030737f
C595 source.n424 a_n2982_n3288# 0.013769f
C596 source.n425 a_n2982_n3288# 0.0242f
C597 source.n426 a_n2982_n3288# 0.013004f
C598 source.n427 a_n2982_n3288# 0.030737f
C599 source.n428 a_n2982_n3288# 0.013769f
C600 source.n429 a_n2982_n3288# 0.0242f
C601 source.n430 a_n2982_n3288# 0.013386f
C602 source.n431 a_n2982_n3288# 0.030737f
C603 source.n432 a_n2982_n3288# 0.013769f
C604 source.n433 a_n2982_n3288# 0.0242f
C605 source.n434 a_n2982_n3288# 0.013004f
C606 source.n435 a_n2982_n3288# 0.030737f
C607 source.n436 a_n2982_n3288# 0.013769f
C608 source.n437 a_n2982_n3288# 0.0242f
C609 source.n438 a_n2982_n3288# 0.013004f
C610 source.n439 a_n2982_n3288# 0.023052f
C611 source.n440 a_n2982_n3288# 0.021728f
C612 source.t9 a_n2982_n3288# 0.051912f
C613 source.n441 a_n2982_n3288# 0.174478f
C614 source.n442 a_n2982_n3288# 1.22084f
C615 source.n443 a_n2982_n3288# 0.013004f
C616 source.n444 a_n2982_n3288# 0.013769f
C617 source.n445 a_n2982_n3288# 0.030737f
C618 source.n446 a_n2982_n3288# 0.030737f
C619 source.n447 a_n2982_n3288# 0.013769f
C620 source.n448 a_n2982_n3288# 0.013004f
C621 source.n449 a_n2982_n3288# 0.0242f
C622 source.n450 a_n2982_n3288# 0.0242f
C623 source.n451 a_n2982_n3288# 0.013004f
C624 source.n452 a_n2982_n3288# 0.013769f
C625 source.n453 a_n2982_n3288# 0.030737f
C626 source.n454 a_n2982_n3288# 0.030737f
C627 source.n455 a_n2982_n3288# 0.013769f
C628 source.n456 a_n2982_n3288# 0.013004f
C629 source.n457 a_n2982_n3288# 0.0242f
C630 source.n458 a_n2982_n3288# 0.0242f
C631 source.n459 a_n2982_n3288# 0.013004f
C632 source.n460 a_n2982_n3288# 0.013004f
C633 source.n461 a_n2982_n3288# 0.013769f
C634 source.n462 a_n2982_n3288# 0.030737f
C635 source.n463 a_n2982_n3288# 0.030737f
C636 source.n464 a_n2982_n3288# 0.030737f
C637 source.n465 a_n2982_n3288# 0.013386f
C638 source.n466 a_n2982_n3288# 0.013004f
C639 source.n467 a_n2982_n3288# 0.0242f
C640 source.n468 a_n2982_n3288# 0.0242f
C641 source.n469 a_n2982_n3288# 0.013004f
C642 source.n470 a_n2982_n3288# 0.013769f
C643 source.n471 a_n2982_n3288# 0.030737f
C644 source.n472 a_n2982_n3288# 0.030737f
C645 source.n473 a_n2982_n3288# 0.013769f
C646 source.n474 a_n2982_n3288# 0.013004f
C647 source.n475 a_n2982_n3288# 0.0242f
C648 source.n476 a_n2982_n3288# 0.0242f
C649 source.n477 a_n2982_n3288# 0.013004f
C650 source.n478 a_n2982_n3288# 0.013769f
C651 source.n479 a_n2982_n3288# 0.030737f
C652 source.n480 a_n2982_n3288# 0.063075f
C653 source.n481 a_n2982_n3288# 0.013769f
C654 source.n482 a_n2982_n3288# 0.013004f
C655 source.n483 a_n2982_n3288# 0.05197f
C656 source.n484 a_n2982_n3288# 0.03481f
C657 source.n485 a_n2982_n3288# 0.124308f
C658 source.t4 a_n2982_n3288# 0.229481f
C659 source.t7 a_n2982_n3288# 0.229481f
C660 source.n486 a_n2982_n3288# 1.96481f
C661 source.n487 a_n2982_n3288# 0.385901f
C662 source.t3 a_n2982_n3288# 0.229481f
C663 source.t39 a_n2982_n3288# 0.229481f
C664 source.n488 a_n2982_n3288# 1.96481f
C665 source.n489 a_n2982_n3288# 0.385901f
C666 source.t15 a_n2982_n3288# 0.229481f
C667 source.t14 a_n2982_n3288# 0.229481f
C668 source.n490 a_n2982_n3288# 1.96481f
C669 source.n491 a_n2982_n3288# 0.385901f
C670 source.t18 a_n2982_n3288# 0.229481f
C671 source.t17 a_n2982_n3288# 0.229481f
C672 source.n492 a_n2982_n3288# 1.96481f
C673 source.n493 a_n2982_n3288# 0.385901f
C674 source.n494 a_n2982_n3288# 0.032056f
C675 source.n495 a_n2982_n3288# 0.0242f
C676 source.n496 a_n2982_n3288# 0.013004f
C677 source.n497 a_n2982_n3288# 0.030737f
C678 source.n498 a_n2982_n3288# 0.013769f
C679 source.n499 a_n2982_n3288# 0.0242f
C680 source.n500 a_n2982_n3288# 0.013004f
C681 source.n501 a_n2982_n3288# 0.030737f
C682 source.n502 a_n2982_n3288# 0.013769f
C683 source.n503 a_n2982_n3288# 0.0242f
C684 source.n504 a_n2982_n3288# 0.013386f
C685 source.n505 a_n2982_n3288# 0.030737f
C686 source.n506 a_n2982_n3288# 0.013769f
C687 source.n507 a_n2982_n3288# 0.0242f
C688 source.n508 a_n2982_n3288# 0.013004f
C689 source.n509 a_n2982_n3288# 0.030737f
C690 source.n510 a_n2982_n3288# 0.013769f
C691 source.n511 a_n2982_n3288# 0.0242f
C692 source.n512 a_n2982_n3288# 0.013004f
C693 source.n513 a_n2982_n3288# 0.023052f
C694 source.n514 a_n2982_n3288# 0.021728f
C695 source.t0 a_n2982_n3288# 0.051912f
C696 source.n515 a_n2982_n3288# 0.174478f
C697 source.n516 a_n2982_n3288# 1.22084f
C698 source.n517 a_n2982_n3288# 0.013004f
C699 source.n518 a_n2982_n3288# 0.013769f
C700 source.n519 a_n2982_n3288# 0.030737f
C701 source.n520 a_n2982_n3288# 0.030737f
C702 source.n521 a_n2982_n3288# 0.013769f
C703 source.n522 a_n2982_n3288# 0.013004f
C704 source.n523 a_n2982_n3288# 0.0242f
C705 source.n524 a_n2982_n3288# 0.0242f
C706 source.n525 a_n2982_n3288# 0.013004f
C707 source.n526 a_n2982_n3288# 0.013769f
C708 source.n527 a_n2982_n3288# 0.030737f
C709 source.n528 a_n2982_n3288# 0.030737f
C710 source.n529 a_n2982_n3288# 0.013769f
C711 source.n530 a_n2982_n3288# 0.013004f
C712 source.n531 a_n2982_n3288# 0.0242f
C713 source.n532 a_n2982_n3288# 0.0242f
C714 source.n533 a_n2982_n3288# 0.013004f
C715 source.n534 a_n2982_n3288# 0.013004f
C716 source.n535 a_n2982_n3288# 0.013769f
C717 source.n536 a_n2982_n3288# 0.030737f
C718 source.n537 a_n2982_n3288# 0.030737f
C719 source.n538 a_n2982_n3288# 0.030737f
C720 source.n539 a_n2982_n3288# 0.013386f
C721 source.n540 a_n2982_n3288# 0.013004f
C722 source.n541 a_n2982_n3288# 0.0242f
C723 source.n542 a_n2982_n3288# 0.0242f
C724 source.n543 a_n2982_n3288# 0.013004f
C725 source.n544 a_n2982_n3288# 0.013769f
C726 source.n545 a_n2982_n3288# 0.030737f
C727 source.n546 a_n2982_n3288# 0.030737f
C728 source.n547 a_n2982_n3288# 0.013769f
C729 source.n548 a_n2982_n3288# 0.013004f
C730 source.n549 a_n2982_n3288# 0.0242f
C731 source.n550 a_n2982_n3288# 0.0242f
C732 source.n551 a_n2982_n3288# 0.013004f
C733 source.n552 a_n2982_n3288# 0.013769f
C734 source.n553 a_n2982_n3288# 0.030737f
C735 source.n554 a_n2982_n3288# 0.063075f
C736 source.n555 a_n2982_n3288# 0.013769f
C737 source.n556 a_n2982_n3288# 0.013004f
C738 source.n557 a_n2982_n3288# 0.05197f
C739 source.n558 a_n2982_n3288# 0.03481f
C740 source.n559 a_n2982_n3288# 0.282164f
C741 source.n560 a_n2982_n3288# 1.53349f
C742 drain_left.t14 a_n2982_n3288# 0.259122f
C743 drain_left.t16 a_n2982_n3288# 0.259122f
C744 drain_left.n0 a_n2982_n3288# 2.31162f
C745 drain_left.t12 a_n2982_n3288# 0.259122f
C746 drain_left.t0 a_n2982_n3288# 0.259122f
C747 drain_left.n1 a_n2982_n3288# 2.30579f
C748 drain_left.n2 a_n2982_n3288# 0.772456f
C749 drain_left.t7 a_n2982_n3288# 0.259122f
C750 drain_left.t10 a_n2982_n3288# 0.259122f
C751 drain_left.n3 a_n2982_n3288# 2.30579f
C752 drain_left.t15 a_n2982_n3288# 0.259122f
C753 drain_left.t2 a_n2982_n3288# 0.259122f
C754 drain_left.n4 a_n2982_n3288# 2.31162f
C755 drain_left.t5 a_n2982_n3288# 0.259122f
C756 drain_left.t13 a_n2982_n3288# 0.259122f
C757 drain_left.n5 a_n2982_n3288# 2.30579f
C758 drain_left.n6 a_n2982_n3288# 0.772456f
C759 drain_left.n7 a_n2982_n3288# 1.99548f
C760 drain_left.t8 a_n2982_n3288# 0.259122f
C761 drain_left.t1 a_n2982_n3288# 0.259122f
C762 drain_left.n8 a_n2982_n3288# 2.31163f
C763 drain_left.t11 a_n2982_n3288# 0.259122f
C764 drain_left.t4 a_n2982_n3288# 0.259122f
C765 drain_left.n9 a_n2982_n3288# 2.3058f
C766 drain_left.n10 a_n2982_n3288# 0.776549f
C767 drain_left.t6 a_n2982_n3288# 0.259122f
C768 drain_left.t17 a_n2982_n3288# 0.259122f
C769 drain_left.n11 a_n2982_n3288# 2.3058f
C770 drain_left.n12 a_n2982_n3288# 0.385686f
C771 drain_left.t18 a_n2982_n3288# 0.259122f
C772 drain_left.t9 a_n2982_n3288# 0.259122f
C773 drain_left.n13 a_n2982_n3288# 2.3058f
C774 drain_left.n14 a_n2982_n3288# 0.385686f
C775 drain_left.t3 a_n2982_n3288# 0.259122f
C776 drain_left.t19 a_n2982_n3288# 0.259122f
C777 drain_left.n15 a_n2982_n3288# 2.30579f
C778 drain_left.n16 a_n2982_n3288# 0.627392f
C779 plus.n0 a_n2982_n3288# 0.040296f
C780 plus.t4 a_n2982_n3288# 0.965196f
C781 plus.t19 a_n2982_n3288# 0.965196f
C782 plus.n1 a_n2982_n3288# 0.040296f
C783 plus.t9 a_n2982_n3288# 0.965196f
C784 plus.n2 a_n2982_n3288# 0.384939f
C785 plus.n3 a_n2982_n3288# 0.040296f
C786 plus.t2 a_n2982_n3288# 0.965196f
C787 plus.t11 a_n2982_n3288# 0.965196f
C788 plus.n4 a_n2982_n3288# 0.384939f
C789 plus.n5 a_n2982_n3288# 0.040296f
C790 plus.t5 a_n2982_n3288# 0.965196f
C791 plus.t10 a_n2982_n3288# 0.965196f
C792 plus.n6 a_n2982_n3288# 0.384939f
C793 plus.n7 a_n2982_n3288# 0.040296f
C794 plus.t3 a_n2982_n3288# 0.965196f
C795 plus.t14 a_n2982_n3288# 0.965196f
C796 plus.n8 a_n2982_n3288# 0.391678f
C797 plus.t6 a_n2982_n3288# 0.984978f
C798 plus.n9 a_n2982_n3288# 0.368049f
C799 plus.n10 a_n2982_n3288# 0.171999f
C800 plus.n11 a_n2982_n3288# 0.009144f
C801 plus.n12 a_n2982_n3288# 0.384939f
C802 plus.n13 a_n2982_n3288# 0.009144f
C803 plus.n14 a_n2982_n3288# 0.040296f
C804 plus.n15 a_n2982_n3288# 0.040296f
C805 plus.n16 a_n2982_n3288# 0.040296f
C806 plus.n17 a_n2982_n3288# 0.009144f
C807 plus.n18 a_n2982_n3288# 0.384939f
C808 plus.n19 a_n2982_n3288# 0.009144f
C809 plus.n20 a_n2982_n3288# 0.040296f
C810 plus.n21 a_n2982_n3288# 0.040296f
C811 plus.n22 a_n2982_n3288# 0.040296f
C812 plus.n23 a_n2982_n3288# 0.009144f
C813 plus.n24 a_n2982_n3288# 0.384939f
C814 plus.n25 a_n2982_n3288# 0.009144f
C815 plus.n26 a_n2982_n3288# 0.040296f
C816 plus.n27 a_n2982_n3288# 0.040296f
C817 plus.n28 a_n2982_n3288# 0.040296f
C818 plus.n29 a_n2982_n3288# 0.009144f
C819 plus.n30 a_n2982_n3288# 0.384939f
C820 plus.n31 a_n2982_n3288# 0.009144f
C821 plus.n32 a_n2982_n3288# 0.384566f
C822 plus.n33 a_n2982_n3288# 0.466886f
C823 plus.n34 a_n2982_n3288# 0.040296f
C824 plus.t13 a_n2982_n3288# 0.965196f
C825 plus.n35 a_n2982_n3288# 0.040296f
C826 plus.t12 a_n2982_n3288# 0.965196f
C827 plus.t16 a_n2982_n3288# 0.965196f
C828 plus.n36 a_n2982_n3288# 0.384939f
C829 plus.n37 a_n2982_n3288# 0.040296f
C830 plus.t1 a_n2982_n3288# 0.965196f
C831 plus.t0 a_n2982_n3288# 0.965196f
C832 plus.n38 a_n2982_n3288# 0.384939f
C833 plus.n39 a_n2982_n3288# 0.040296f
C834 plus.t8 a_n2982_n3288# 0.965196f
C835 plus.t7 a_n2982_n3288# 0.965196f
C836 plus.n40 a_n2982_n3288# 0.384939f
C837 plus.n41 a_n2982_n3288# 0.040296f
C838 plus.t15 a_n2982_n3288# 0.965196f
C839 plus.t18 a_n2982_n3288# 0.965196f
C840 plus.n42 a_n2982_n3288# 0.391678f
C841 plus.t17 a_n2982_n3288# 0.984978f
C842 plus.n43 a_n2982_n3288# 0.368049f
C843 plus.n44 a_n2982_n3288# 0.171999f
C844 plus.n45 a_n2982_n3288# 0.009144f
C845 plus.n46 a_n2982_n3288# 0.384939f
C846 plus.n47 a_n2982_n3288# 0.009144f
C847 plus.n48 a_n2982_n3288# 0.040296f
C848 plus.n49 a_n2982_n3288# 0.040296f
C849 plus.n50 a_n2982_n3288# 0.040296f
C850 plus.n51 a_n2982_n3288# 0.009144f
C851 plus.n52 a_n2982_n3288# 0.384939f
C852 plus.n53 a_n2982_n3288# 0.009144f
C853 plus.n54 a_n2982_n3288# 0.040296f
C854 plus.n55 a_n2982_n3288# 0.040296f
C855 plus.n56 a_n2982_n3288# 0.040296f
C856 plus.n57 a_n2982_n3288# 0.009144f
C857 plus.n58 a_n2982_n3288# 0.384939f
C858 plus.n59 a_n2982_n3288# 0.009144f
C859 plus.n60 a_n2982_n3288# 0.040296f
C860 plus.n61 a_n2982_n3288# 0.040296f
C861 plus.n62 a_n2982_n3288# 0.040296f
C862 plus.n63 a_n2982_n3288# 0.009144f
C863 plus.n64 a_n2982_n3288# 0.384939f
C864 plus.n65 a_n2982_n3288# 0.009144f
C865 plus.n66 a_n2982_n3288# 0.384566f
C866 plus.n67 a_n2982_n3288# 1.4559f
.ends

