* NGSPICE file created from diffpair51.ext - technology: sky130A

.subckt diffpair51 minus drain_right drain_left source plus
X0 a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X1 source plus drain_left a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X2 a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X3 a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X4 drain_right minus source a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X5 drain_left plus source a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X6 source minus drain_right a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X7 drain_right minus source a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X8 drain_left plus source a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X9 source plus drain_left a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X10 a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X11 source minus drain_right a_n1274_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
.ends

