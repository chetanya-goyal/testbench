* NGSPICE file created from diffpair257.ext - technology: sky130A

.subckt diffpair257 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t1 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X1 drain_right.t10 minus.t1 source.t30 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 drain_right.t8 minus.t2 source.t29 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X3 source.t28 minus.t3 drain_right.t7 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X5 source.t4 plus.t0 drain_left.t15 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X6 drain_left.t14 plus.t1 source.t15 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 source.t14 plus.t2 drain_left.t13 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X8 source.t6 plus.t3 drain_left.t12 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X9 source.t27 minus.t4 drain_right.t3 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X10 source.t5 plus.t4 drain_left.t11 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X11 source.t26 minus.t5 drain_right.t2 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X12 drain_left.t10 plus.t5 source.t7 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X13 drain_left.t9 plus.t6 source.t12 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X14 source.t0 plus.t7 drain_left.t8 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X15 drain_left.t7 plus.t8 source.t13 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X16 drain_left.t6 plus.t9 source.t1 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X17 a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X18 drain_left.t5 plus.t10 source.t8 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X19 a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X20 drain_right.t0 minus.t6 source.t25 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X21 drain_right.t6 minus.t7 source.t24 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X22 source.t11 plus.t11 drain_left.t4 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X23 source.t3 plus.t12 drain_left.t3 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X24 drain_left.t2 plus.t13 source.t9 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X25 source.t23 minus.t8 drain_right.t14 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X26 source.t22 minus.t9 drain_right.t13 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X27 source.t21 minus.t10 drain_right.t12 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X28 source.t20 minus.t11 drain_right.t5 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X29 drain_right.t15 minus.t12 source.t19 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X30 drain_right.t11 minus.t13 source.t18 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X31 drain_left.t1 plus.t14 source.t2 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X32 source.t10 plus.t15 drain_left.t0 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X33 a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X34 drain_right.t9 minus.t14 source.t17 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X35 drain_right.t4 minus.t15 source.t16 a_n1670_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n17 minus.t11 931.503
R1 minus.n4 minus.t6 931.503
R2 minus.n36 minus.t14 931.503
R3 minus.n23 minus.t9 931.503
R4 minus.n16 minus.t2 879.65
R5 minus.n14 minus.t4 879.65
R6 minus.n1 minus.t7 879.65
R7 minus.n9 minus.t10 879.65
R8 minus.n7 minus.t1 879.65
R9 minus.n3 minus.t5 879.65
R10 minus.n35 minus.t0 879.65
R11 minus.n33 minus.t15 879.65
R12 minus.n20 minus.t3 879.65
R13 minus.n28 minus.t12 879.65
R14 minus.n26 minus.t8 879.65
R15 minus.n22 minus.t13 879.65
R16 minus.n5 minus.n4 161.489
R17 minus.n24 minus.n23 161.489
R18 minus.n18 minus.n17 161.3
R19 minus.n15 minus.n0 161.3
R20 minus.n13 minus.n12 161.3
R21 minus.n11 minus.n10 161.3
R22 minus.n8 minus.n2 161.3
R23 minus.n6 minus.n5 161.3
R24 minus.n37 minus.n36 161.3
R25 minus.n34 minus.n19 161.3
R26 minus.n32 minus.n31 161.3
R27 minus.n30 minus.n29 161.3
R28 minus.n27 minus.n21 161.3
R29 minus.n25 minus.n24 161.3
R30 minus.n16 minus.n15 47.4702
R31 minus.n6 minus.n3 47.4702
R32 minus.n25 minus.n22 47.4702
R33 minus.n35 minus.n34 47.4702
R34 minus.n14 minus.n13 43.0884
R35 minus.n8 minus.n7 43.0884
R36 minus.n27 minus.n26 43.0884
R37 minus.n33 minus.n32 43.0884
R38 minus.n10 minus.n1 38.7066
R39 minus.n10 minus.n9 38.7066
R40 minus.n29 minus.n28 38.7066
R41 minus.n29 minus.n20 38.7066
R42 minus.n13 minus.n1 34.3247
R43 minus.n9 minus.n8 34.3247
R44 minus.n28 minus.n27 34.3247
R45 minus.n32 minus.n20 34.3247
R46 minus.n38 minus.n18 30.8679
R47 minus.n15 minus.n14 29.9429
R48 minus.n7 minus.n6 29.9429
R49 minus.n26 minus.n25 29.9429
R50 minus.n34 minus.n33 29.9429
R51 minus.n17 minus.n16 25.5611
R52 minus.n4 minus.n3 25.5611
R53 minus.n23 minus.n22 25.5611
R54 minus.n36 minus.n35 25.5611
R55 minus.n38 minus.n37 6.46641
R56 minus.n18 minus.n0 0.189894
R57 minus.n12 minus.n0 0.189894
R58 minus.n12 minus.n11 0.189894
R59 minus.n11 minus.n2 0.189894
R60 minus.n5 minus.n2 0.189894
R61 minus.n24 minus.n21 0.189894
R62 minus.n30 minus.n21 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n19 0.189894
R65 minus.n37 minus.n19 0.189894
R66 minus minus.n38 0.188
R67 drain_right.n5 drain_right.n3 67.6476
R68 drain_right.n2 drain_right.n0 67.6476
R69 drain_right.n9 drain_right.n7 67.6476
R70 drain_right.n9 drain_right.n8 67.1908
R71 drain_right.n11 drain_right.n10 67.1908
R72 drain_right.n13 drain_right.n12 67.1908
R73 drain_right.n5 drain_right.n4 67.1907
R74 drain_right.n2 drain_right.n1 67.1907
R75 drain_right drain_right.n6 25.2382
R76 drain_right drain_right.n13 6.11011
R77 drain_right.n3 drain_right.t1 3.3005
R78 drain_right.n3 drain_right.t9 3.3005
R79 drain_right.n4 drain_right.t7 3.3005
R80 drain_right.n4 drain_right.t4 3.3005
R81 drain_right.n1 drain_right.t14 3.3005
R82 drain_right.n1 drain_right.t15 3.3005
R83 drain_right.n0 drain_right.t13 3.3005
R84 drain_right.n0 drain_right.t11 3.3005
R85 drain_right.n7 drain_right.t2 3.3005
R86 drain_right.n7 drain_right.t0 3.3005
R87 drain_right.n8 drain_right.t12 3.3005
R88 drain_right.n8 drain_right.t10 3.3005
R89 drain_right.n10 drain_right.t3 3.3005
R90 drain_right.n10 drain_right.t6 3.3005
R91 drain_right.n12 drain_right.t5 3.3005
R92 drain_right.n12 drain_right.t8 3.3005
R93 drain_right.n13 drain_right.n11 0.457397
R94 drain_right.n11 drain_right.n9 0.457397
R95 drain_right.n6 drain_right.n5 0.173602
R96 drain_right.n6 drain_right.n2 0.173602
R97 source.n274 source.n248 289.615
R98 source.n236 source.n210 289.615
R99 source.n204 source.n178 289.615
R100 source.n166 source.n140 289.615
R101 source.n26 source.n0 289.615
R102 source.n64 source.n38 289.615
R103 source.n96 source.n70 289.615
R104 source.n134 source.n108 289.615
R105 source.n259 source.n258 185
R106 source.n256 source.n255 185
R107 source.n265 source.n264 185
R108 source.n267 source.n266 185
R109 source.n252 source.n251 185
R110 source.n273 source.n272 185
R111 source.n275 source.n274 185
R112 source.n221 source.n220 185
R113 source.n218 source.n217 185
R114 source.n227 source.n226 185
R115 source.n229 source.n228 185
R116 source.n214 source.n213 185
R117 source.n235 source.n234 185
R118 source.n237 source.n236 185
R119 source.n189 source.n188 185
R120 source.n186 source.n185 185
R121 source.n195 source.n194 185
R122 source.n197 source.n196 185
R123 source.n182 source.n181 185
R124 source.n203 source.n202 185
R125 source.n205 source.n204 185
R126 source.n151 source.n150 185
R127 source.n148 source.n147 185
R128 source.n157 source.n156 185
R129 source.n159 source.n158 185
R130 source.n144 source.n143 185
R131 source.n165 source.n164 185
R132 source.n167 source.n166 185
R133 source.n27 source.n26 185
R134 source.n25 source.n24 185
R135 source.n4 source.n3 185
R136 source.n19 source.n18 185
R137 source.n17 source.n16 185
R138 source.n8 source.n7 185
R139 source.n11 source.n10 185
R140 source.n65 source.n64 185
R141 source.n63 source.n62 185
R142 source.n42 source.n41 185
R143 source.n57 source.n56 185
R144 source.n55 source.n54 185
R145 source.n46 source.n45 185
R146 source.n49 source.n48 185
R147 source.n97 source.n96 185
R148 source.n95 source.n94 185
R149 source.n74 source.n73 185
R150 source.n89 source.n88 185
R151 source.n87 source.n86 185
R152 source.n78 source.n77 185
R153 source.n81 source.n80 185
R154 source.n135 source.n134 185
R155 source.n133 source.n132 185
R156 source.n112 source.n111 185
R157 source.n127 source.n126 185
R158 source.n125 source.n124 185
R159 source.n116 source.n115 185
R160 source.n119 source.n118 185
R161 source.t17 source.n257 147.661
R162 source.t22 source.n219 147.661
R163 source.t8 source.n187 147.661
R164 source.t14 source.n149 147.661
R165 source.t2 source.n9 147.661
R166 source.t0 source.n47 147.661
R167 source.t25 source.n79 147.661
R168 source.t20 source.n117 147.661
R169 source.n258 source.n255 104.615
R170 source.n265 source.n255 104.615
R171 source.n266 source.n265 104.615
R172 source.n266 source.n251 104.615
R173 source.n273 source.n251 104.615
R174 source.n274 source.n273 104.615
R175 source.n220 source.n217 104.615
R176 source.n227 source.n217 104.615
R177 source.n228 source.n227 104.615
R178 source.n228 source.n213 104.615
R179 source.n235 source.n213 104.615
R180 source.n236 source.n235 104.615
R181 source.n188 source.n185 104.615
R182 source.n195 source.n185 104.615
R183 source.n196 source.n195 104.615
R184 source.n196 source.n181 104.615
R185 source.n203 source.n181 104.615
R186 source.n204 source.n203 104.615
R187 source.n150 source.n147 104.615
R188 source.n157 source.n147 104.615
R189 source.n158 source.n157 104.615
R190 source.n158 source.n143 104.615
R191 source.n165 source.n143 104.615
R192 source.n166 source.n165 104.615
R193 source.n26 source.n25 104.615
R194 source.n25 source.n3 104.615
R195 source.n18 source.n3 104.615
R196 source.n18 source.n17 104.615
R197 source.n17 source.n7 104.615
R198 source.n10 source.n7 104.615
R199 source.n64 source.n63 104.615
R200 source.n63 source.n41 104.615
R201 source.n56 source.n41 104.615
R202 source.n56 source.n55 104.615
R203 source.n55 source.n45 104.615
R204 source.n48 source.n45 104.615
R205 source.n96 source.n95 104.615
R206 source.n95 source.n73 104.615
R207 source.n88 source.n73 104.615
R208 source.n88 source.n87 104.615
R209 source.n87 source.n77 104.615
R210 source.n80 source.n77 104.615
R211 source.n134 source.n133 104.615
R212 source.n133 source.n111 104.615
R213 source.n126 source.n111 104.615
R214 source.n126 source.n125 104.615
R215 source.n125 source.n115 104.615
R216 source.n118 source.n115 104.615
R217 source.n258 source.t17 52.3082
R218 source.n220 source.t22 52.3082
R219 source.n188 source.t8 52.3082
R220 source.n150 source.t14 52.3082
R221 source.n10 source.t2 52.3082
R222 source.n48 source.t0 52.3082
R223 source.n80 source.t25 52.3082
R224 source.n118 source.t20 52.3082
R225 source.n33 source.n32 50.512
R226 source.n35 source.n34 50.512
R227 source.n37 source.n36 50.512
R228 source.n103 source.n102 50.512
R229 source.n105 source.n104 50.512
R230 source.n107 source.n106 50.512
R231 source.n247 source.n246 50.5119
R232 source.n245 source.n244 50.5119
R233 source.n243 source.n242 50.5119
R234 source.n177 source.n176 50.5119
R235 source.n175 source.n174 50.5119
R236 source.n173 source.n172 50.5119
R237 source.n279 source.n278 32.1853
R238 source.n241 source.n240 32.1853
R239 source.n209 source.n208 32.1853
R240 source.n171 source.n170 32.1853
R241 source.n31 source.n30 32.1853
R242 source.n69 source.n68 32.1853
R243 source.n101 source.n100 32.1853
R244 source.n139 source.n138 32.1853
R245 source.n171 source.n139 17.1992
R246 source.n259 source.n257 15.6674
R247 source.n221 source.n219 15.6674
R248 source.n189 source.n187 15.6674
R249 source.n151 source.n149 15.6674
R250 source.n11 source.n9 15.6674
R251 source.n49 source.n47 15.6674
R252 source.n81 source.n79 15.6674
R253 source.n119 source.n117 15.6674
R254 source.n260 source.n256 12.8005
R255 source.n222 source.n218 12.8005
R256 source.n190 source.n186 12.8005
R257 source.n152 source.n148 12.8005
R258 source.n12 source.n8 12.8005
R259 source.n50 source.n46 12.8005
R260 source.n82 source.n78 12.8005
R261 source.n120 source.n116 12.8005
R262 source.n264 source.n263 12.0247
R263 source.n226 source.n225 12.0247
R264 source.n194 source.n193 12.0247
R265 source.n156 source.n155 12.0247
R266 source.n16 source.n15 12.0247
R267 source.n54 source.n53 12.0247
R268 source.n86 source.n85 12.0247
R269 source.n124 source.n123 12.0247
R270 source.n280 source.n31 11.7078
R271 source.n267 source.n254 11.249
R272 source.n229 source.n216 11.249
R273 source.n197 source.n184 11.249
R274 source.n159 source.n146 11.249
R275 source.n19 source.n6 11.249
R276 source.n57 source.n44 11.249
R277 source.n89 source.n76 11.249
R278 source.n127 source.n114 11.249
R279 source.n268 source.n252 10.4732
R280 source.n230 source.n214 10.4732
R281 source.n198 source.n182 10.4732
R282 source.n160 source.n144 10.4732
R283 source.n20 source.n4 10.4732
R284 source.n58 source.n42 10.4732
R285 source.n90 source.n74 10.4732
R286 source.n128 source.n112 10.4732
R287 source.n272 source.n271 9.69747
R288 source.n234 source.n233 9.69747
R289 source.n202 source.n201 9.69747
R290 source.n164 source.n163 9.69747
R291 source.n24 source.n23 9.69747
R292 source.n62 source.n61 9.69747
R293 source.n94 source.n93 9.69747
R294 source.n132 source.n131 9.69747
R295 source.n278 source.n277 9.45567
R296 source.n240 source.n239 9.45567
R297 source.n208 source.n207 9.45567
R298 source.n170 source.n169 9.45567
R299 source.n30 source.n29 9.45567
R300 source.n68 source.n67 9.45567
R301 source.n100 source.n99 9.45567
R302 source.n138 source.n137 9.45567
R303 source.n277 source.n276 9.3005
R304 source.n250 source.n249 9.3005
R305 source.n271 source.n270 9.3005
R306 source.n269 source.n268 9.3005
R307 source.n254 source.n253 9.3005
R308 source.n263 source.n262 9.3005
R309 source.n261 source.n260 9.3005
R310 source.n239 source.n238 9.3005
R311 source.n212 source.n211 9.3005
R312 source.n233 source.n232 9.3005
R313 source.n231 source.n230 9.3005
R314 source.n216 source.n215 9.3005
R315 source.n225 source.n224 9.3005
R316 source.n223 source.n222 9.3005
R317 source.n207 source.n206 9.3005
R318 source.n180 source.n179 9.3005
R319 source.n201 source.n200 9.3005
R320 source.n199 source.n198 9.3005
R321 source.n184 source.n183 9.3005
R322 source.n193 source.n192 9.3005
R323 source.n191 source.n190 9.3005
R324 source.n169 source.n168 9.3005
R325 source.n142 source.n141 9.3005
R326 source.n163 source.n162 9.3005
R327 source.n161 source.n160 9.3005
R328 source.n146 source.n145 9.3005
R329 source.n155 source.n154 9.3005
R330 source.n153 source.n152 9.3005
R331 source.n29 source.n28 9.3005
R332 source.n2 source.n1 9.3005
R333 source.n23 source.n22 9.3005
R334 source.n21 source.n20 9.3005
R335 source.n6 source.n5 9.3005
R336 source.n15 source.n14 9.3005
R337 source.n13 source.n12 9.3005
R338 source.n67 source.n66 9.3005
R339 source.n40 source.n39 9.3005
R340 source.n61 source.n60 9.3005
R341 source.n59 source.n58 9.3005
R342 source.n44 source.n43 9.3005
R343 source.n53 source.n52 9.3005
R344 source.n51 source.n50 9.3005
R345 source.n99 source.n98 9.3005
R346 source.n72 source.n71 9.3005
R347 source.n93 source.n92 9.3005
R348 source.n91 source.n90 9.3005
R349 source.n76 source.n75 9.3005
R350 source.n85 source.n84 9.3005
R351 source.n83 source.n82 9.3005
R352 source.n137 source.n136 9.3005
R353 source.n110 source.n109 9.3005
R354 source.n131 source.n130 9.3005
R355 source.n129 source.n128 9.3005
R356 source.n114 source.n113 9.3005
R357 source.n123 source.n122 9.3005
R358 source.n121 source.n120 9.3005
R359 source.n275 source.n250 8.92171
R360 source.n237 source.n212 8.92171
R361 source.n205 source.n180 8.92171
R362 source.n167 source.n142 8.92171
R363 source.n27 source.n2 8.92171
R364 source.n65 source.n40 8.92171
R365 source.n97 source.n72 8.92171
R366 source.n135 source.n110 8.92171
R367 source.n276 source.n248 8.14595
R368 source.n238 source.n210 8.14595
R369 source.n206 source.n178 8.14595
R370 source.n168 source.n140 8.14595
R371 source.n28 source.n0 8.14595
R372 source.n66 source.n38 8.14595
R373 source.n98 source.n70 8.14595
R374 source.n136 source.n108 8.14595
R375 source.n278 source.n248 5.81868
R376 source.n240 source.n210 5.81868
R377 source.n208 source.n178 5.81868
R378 source.n170 source.n140 5.81868
R379 source.n30 source.n0 5.81868
R380 source.n68 source.n38 5.81868
R381 source.n100 source.n70 5.81868
R382 source.n138 source.n108 5.81868
R383 source.n280 source.n279 5.49188
R384 source.n276 source.n275 5.04292
R385 source.n238 source.n237 5.04292
R386 source.n206 source.n205 5.04292
R387 source.n168 source.n167 5.04292
R388 source.n28 source.n27 5.04292
R389 source.n66 source.n65 5.04292
R390 source.n98 source.n97 5.04292
R391 source.n136 source.n135 5.04292
R392 source.n261 source.n257 4.38594
R393 source.n223 source.n219 4.38594
R394 source.n191 source.n187 4.38594
R395 source.n153 source.n149 4.38594
R396 source.n13 source.n9 4.38594
R397 source.n51 source.n47 4.38594
R398 source.n83 source.n79 4.38594
R399 source.n121 source.n117 4.38594
R400 source.n272 source.n250 4.26717
R401 source.n234 source.n212 4.26717
R402 source.n202 source.n180 4.26717
R403 source.n164 source.n142 4.26717
R404 source.n24 source.n2 4.26717
R405 source.n62 source.n40 4.26717
R406 source.n94 source.n72 4.26717
R407 source.n132 source.n110 4.26717
R408 source.n271 source.n252 3.49141
R409 source.n233 source.n214 3.49141
R410 source.n201 source.n182 3.49141
R411 source.n163 source.n144 3.49141
R412 source.n23 source.n4 3.49141
R413 source.n61 source.n42 3.49141
R414 source.n93 source.n74 3.49141
R415 source.n131 source.n112 3.49141
R416 source.n246 source.t16 3.3005
R417 source.n246 source.t31 3.3005
R418 source.n244 source.t19 3.3005
R419 source.n244 source.t28 3.3005
R420 source.n242 source.t18 3.3005
R421 source.n242 source.t23 3.3005
R422 source.n176 source.t13 3.3005
R423 source.n176 source.t11 3.3005
R424 source.n174 source.t1 3.3005
R425 source.n174 source.t5 3.3005
R426 source.n172 source.t7 3.3005
R427 source.n172 source.t6 3.3005
R428 source.n32 source.t12 3.3005
R429 source.n32 source.t4 3.3005
R430 source.n34 source.t9 3.3005
R431 source.n34 source.t3 3.3005
R432 source.n36 source.t15 3.3005
R433 source.n36 source.t10 3.3005
R434 source.n102 source.t30 3.3005
R435 source.n102 source.t26 3.3005
R436 source.n104 source.t24 3.3005
R437 source.n104 source.t21 3.3005
R438 source.n106 source.t29 3.3005
R439 source.n106 source.t27 3.3005
R440 source.n268 source.n267 2.71565
R441 source.n230 source.n229 2.71565
R442 source.n198 source.n197 2.71565
R443 source.n160 source.n159 2.71565
R444 source.n20 source.n19 2.71565
R445 source.n58 source.n57 2.71565
R446 source.n90 source.n89 2.71565
R447 source.n128 source.n127 2.71565
R448 source.n264 source.n254 1.93989
R449 source.n226 source.n216 1.93989
R450 source.n194 source.n184 1.93989
R451 source.n156 source.n146 1.93989
R452 source.n16 source.n6 1.93989
R453 source.n54 source.n44 1.93989
R454 source.n86 source.n76 1.93989
R455 source.n124 source.n114 1.93989
R456 source.n263 source.n256 1.16414
R457 source.n225 source.n218 1.16414
R458 source.n193 source.n186 1.16414
R459 source.n155 source.n148 1.16414
R460 source.n15 source.n8 1.16414
R461 source.n53 source.n46 1.16414
R462 source.n85 source.n78 1.16414
R463 source.n123 source.n116 1.16414
R464 source.n101 source.n69 0.470328
R465 source.n241 source.n209 0.470328
R466 source.n139 source.n107 0.457397
R467 source.n107 source.n105 0.457397
R468 source.n105 source.n103 0.457397
R469 source.n103 source.n101 0.457397
R470 source.n69 source.n37 0.457397
R471 source.n37 source.n35 0.457397
R472 source.n35 source.n33 0.457397
R473 source.n33 source.n31 0.457397
R474 source.n173 source.n171 0.457397
R475 source.n175 source.n173 0.457397
R476 source.n177 source.n175 0.457397
R477 source.n209 source.n177 0.457397
R478 source.n243 source.n241 0.457397
R479 source.n245 source.n243 0.457397
R480 source.n247 source.n245 0.457397
R481 source.n279 source.n247 0.457397
R482 source.n260 source.n259 0.388379
R483 source.n222 source.n221 0.388379
R484 source.n190 source.n189 0.388379
R485 source.n152 source.n151 0.388379
R486 source.n12 source.n11 0.388379
R487 source.n50 source.n49 0.388379
R488 source.n82 source.n81 0.388379
R489 source.n120 source.n119 0.388379
R490 source source.n280 0.188
R491 source.n262 source.n261 0.155672
R492 source.n262 source.n253 0.155672
R493 source.n269 source.n253 0.155672
R494 source.n270 source.n269 0.155672
R495 source.n270 source.n249 0.155672
R496 source.n277 source.n249 0.155672
R497 source.n224 source.n223 0.155672
R498 source.n224 source.n215 0.155672
R499 source.n231 source.n215 0.155672
R500 source.n232 source.n231 0.155672
R501 source.n232 source.n211 0.155672
R502 source.n239 source.n211 0.155672
R503 source.n192 source.n191 0.155672
R504 source.n192 source.n183 0.155672
R505 source.n199 source.n183 0.155672
R506 source.n200 source.n199 0.155672
R507 source.n200 source.n179 0.155672
R508 source.n207 source.n179 0.155672
R509 source.n154 source.n153 0.155672
R510 source.n154 source.n145 0.155672
R511 source.n161 source.n145 0.155672
R512 source.n162 source.n161 0.155672
R513 source.n162 source.n141 0.155672
R514 source.n169 source.n141 0.155672
R515 source.n29 source.n1 0.155672
R516 source.n22 source.n1 0.155672
R517 source.n22 source.n21 0.155672
R518 source.n21 source.n5 0.155672
R519 source.n14 source.n5 0.155672
R520 source.n14 source.n13 0.155672
R521 source.n67 source.n39 0.155672
R522 source.n60 source.n39 0.155672
R523 source.n60 source.n59 0.155672
R524 source.n59 source.n43 0.155672
R525 source.n52 source.n43 0.155672
R526 source.n52 source.n51 0.155672
R527 source.n99 source.n71 0.155672
R528 source.n92 source.n71 0.155672
R529 source.n92 source.n91 0.155672
R530 source.n91 source.n75 0.155672
R531 source.n84 source.n75 0.155672
R532 source.n84 source.n83 0.155672
R533 source.n137 source.n109 0.155672
R534 source.n130 source.n109 0.155672
R535 source.n130 source.n129 0.155672
R536 source.n129 source.n113 0.155672
R537 source.n122 source.n113 0.155672
R538 source.n122 source.n121 0.155672
R539 plus.n4 plus.t7 931.503
R540 plus.n17 plus.t14 931.503
R541 plus.n23 plus.t10 931.503
R542 plus.n36 plus.t2 931.503
R543 plus.n3 plus.t1 879.65
R544 plus.n7 plus.t15 879.65
R545 plus.n9 plus.t13 879.65
R546 plus.n1 plus.t12 879.65
R547 plus.n14 plus.t6 879.65
R548 plus.n16 plus.t0 879.65
R549 plus.n22 plus.t11 879.65
R550 plus.n26 plus.t8 879.65
R551 plus.n28 plus.t4 879.65
R552 plus.n20 plus.t9 879.65
R553 plus.n33 plus.t3 879.65
R554 plus.n35 plus.t5 879.65
R555 plus.n5 plus.n4 161.489
R556 plus.n24 plus.n23 161.489
R557 plus.n6 plus.n5 161.3
R558 plus.n8 plus.n2 161.3
R559 plus.n11 plus.n10 161.3
R560 plus.n13 plus.n12 161.3
R561 plus.n15 plus.n0 161.3
R562 plus.n18 plus.n17 161.3
R563 plus.n25 plus.n24 161.3
R564 plus.n27 plus.n21 161.3
R565 plus.n30 plus.n29 161.3
R566 plus.n32 plus.n31 161.3
R567 plus.n34 plus.n19 161.3
R568 plus.n37 plus.n36 161.3
R569 plus.n6 plus.n3 47.4702
R570 plus.n16 plus.n15 47.4702
R571 plus.n35 plus.n34 47.4702
R572 plus.n25 plus.n22 47.4702
R573 plus.n8 plus.n7 43.0884
R574 plus.n14 plus.n13 43.0884
R575 plus.n33 plus.n32 43.0884
R576 plus.n27 plus.n26 43.0884
R577 plus.n10 plus.n9 38.7066
R578 plus.n10 plus.n1 38.7066
R579 plus.n29 plus.n20 38.7066
R580 plus.n29 plus.n28 38.7066
R581 plus.n9 plus.n8 34.3247
R582 plus.n13 plus.n1 34.3247
R583 plus.n32 plus.n20 34.3247
R584 plus.n28 plus.n27 34.3247
R585 plus.n7 plus.n6 29.9429
R586 plus.n15 plus.n14 29.9429
R587 plus.n34 plus.n33 29.9429
R588 plus.n26 plus.n25 29.9429
R589 plus plus.n37 27.0217
R590 plus.n4 plus.n3 25.5611
R591 plus.n17 plus.n16 25.5611
R592 plus.n36 plus.n35 25.5611
R593 plus.n23 plus.n22 25.5611
R594 plus plus.n18 9.83762
R595 plus.n5 plus.n2 0.189894
R596 plus.n11 plus.n2 0.189894
R597 plus.n12 plus.n11 0.189894
R598 plus.n12 plus.n0 0.189894
R599 plus.n18 plus.n0 0.189894
R600 plus.n37 plus.n19 0.189894
R601 plus.n31 plus.n19 0.189894
R602 plus.n31 plus.n30 0.189894
R603 plus.n30 plus.n21 0.189894
R604 plus.n24 plus.n21 0.189894
R605 drain_left.n9 drain_left.n7 67.6477
R606 drain_left.n5 drain_left.n3 67.6476
R607 drain_left.n2 drain_left.n0 67.6476
R608 drain_left.n11 drain_left.n10 67.1908
R609 drain_left.n9 drain_left.n8 67.1908
R610 drain_left.n13 drain_left.n12 67.1907
R611 drain_left.n5 drain_left.n4 67.1907
R612 drain_left.n2 drain_left.n1 67.1907
R613 drain_left drain_left.n6 25.7914
R614 drain_left drain_left.n13 6.11011
R615 drain_left.n3 drain_left.t4 3.3005
R616 drain_left.n3 drain_left.t5 3.3005
R617 drain_left.n4 drain_left.t11 3.3005
R618 drain_left.n4 drain_left.t7 3.3005
R619 drain_left.n1 drain_left.t12 3.3005
R620 drain_left.n1 drain_left.t6 3.3005
R621 drain_left.n0 drain_left.t13 3.3005
R622 drain_left.n0 drain_left.t10 3.3005
R623 drain_left.n12 drain_left.t15 3.3005
R624 drain_left.n12 drain_left.t1 3.3005
R625 drain_left.n10 drain_left.t3 3.3005
R626 drain_left.n10 drain_left.t9 3.3005
R627 drain_left.n8 drain_left.t0 3.3005
R628 drain_left.n8 drain_left.t2 3.3005
R629 drain_left.n7 drain_left.t8 3.3005
R630 drain_left.n7 drain_left.t14 3.3005
R631 drain_left.n11 drain_left.n9 0.457397
R632 drain_left.n13 drain_left.n11 0.457397
R633 drain_left.n6 drain_left.n5 0.173602
R634 drain_left.n6 drain_left.n2 0.173602
C0 drain_left source 19.7024f
C1 source plus 2.37886f
C2 drain_left minus 0.170856f
C3 plus minus 4.12612f
C4 drain_right source 19.702f
C5 drain_left plus 2.62482f
C6 drain_right minus 2.46385f
C7 drain_right drain_left 0.846053f
C8 drain_right plus 0.314737f
C9 source minus 2.36484f
C10 drain_right a_n1670_n2088# 5.28617f
C11 drain_left a_n1670_n2088# 5.55084f
C12 source a_n1670_n2088# 5.233456f
C13 minus a_n1670_n2088# 6.006576f
C14 plus a_n1670_n2088# 7.63938f
C15 drain_left.t13 a_n1670_n2088# 0.177955f
C16 drain_left.t10 a_n1670_n2088# 0.177955f
C17 drain_left.n0 a_n1670_n2088# 1.48706f
C18 drain_left.t12 a_n1670_n2088# 0.177955f
C19 drain_left.t6 a_n1670_n2088# 0.177955f
C20 drain_left.n1 a_n1670_n2088# 1.48415f
C21 drain_left.n2 a_n1670_n2088# 0.813193f
C22 drain_left.t4 a_n1670_n2088# 0.177955f
C23 drain_left.t5 a_n1670_n2088# 0.177955f
C24 drain_left.n3 a_n1670_n2088# 1.48706f
C25 drain_left.t11 a_n1670_n2088# 0.177955f
C26 drain_left.t7 a_n1670_n2088# 0.177955f
C27 drain_left.n4 a_n1670_n2088# 1.48415f
C28 drain_left.n5 a_n1670_n2088# 0.813193f
C29 drain_left.n6 a_n1670_n2088# 1.27169f
C30 drain_left.t8 a_n1670_n2088# 0.177955f
C31 drain_left.t14 a_n1670_n2088# 0.177955f
C32 drain_left.n7 a_n1670_n2088# 1.48706f
C33 drain_left.t0 a_n1670_n2088# 0.177955f
C34 drain_left.t2 a_n1670_n2088# 0.177955f
C35 drain_left.n8 a_n1670_n2088# 1.48416f
C36 drain_left.n9 a_n1670_n2088# 0.842474f
C37 drain_left.t3 a_n1670_n2088# 0.177955f
C38 drain_left.t9 a_n1670_n2088# 0.177955f
C39 drain_left.n10 a_n1670_n2088# 1.48416f
C40 drain_left.n11 a_n1670_n2088# 0.415131f
C41 drain_left.t15 a_n1670_n2088# 0.177955f
C42 drain_left.t1 a_n1670_n2088# 0.177955f
C43 drain_left.n12 a_n1670_n2088# 1.48415f
C44 drain_left.n13 a_n1670_n2088# 0.722305f
C45 plus.n0 a_n1670_n2088# 0.055152f
C46 plus.t0 a_n1670_n2088# 0.188565f
C47 plus.t6 a_n1670_n2088# 0.188565f
C48 plus.t12 a_n1670_n2088# 0.188565f
C49 plus.n1 a_n1670_n2088# 0.092222f
C50 plus.n2 a_n1670_n2088# 0.055152f
C51 plus.t13 a_n1670_n2088# 0.188565f
C52 plus.t15 a_n1670_n2088# 0.188565f
C53 plus.t1 a_n1670_n2088# 0.188565f
C54 plus.n3 a_n1670_n2088# 0.092222f
C55 plus.t7 a_n1670_n2088# 0.193803f
C56 plus.n4 a_n1670_n2088# 0.108251f
C57 plus.n5 a_n1670_n2088# 0.124164f
C58 plus.n6 a_n1670_n2088# 0.019316f
C59 plus.n7 a_n1670_n2088# 0.092222f
C60 plus.n8 a_n1670_n2088# 0.019316f
C61 plus.n9 a_n1670_n2088# 0.092222f
C62 plus.n10 a_n1670_n2088# 0.019316f
C63 plus.n11 a_n1670_n2088# 0.055152f
C64 plus.n12 a_n1670_n2088# 0.055152f
C65 plus.n13 a_n1670_n2088# 0.019316f
C66 plus.n14 a_n1670_n2088# 0.092222f
C67 plus.n15 a_n1670_n2088# 0.019316f
C68 plus.n16 a_n1670_n2088# 0.092222f
C69 plus.t14 a_n1670_n2088# 0.193803f
C70 plus.n17 a_n1670_n2088# 0.10817f
C71 plus.n18 a_n1670_n2088# 0.468037f
C72 plus.n19 a_n1670_n2088# 0.055152f
C73 plus.t2 a_n1670_n2088# 0.193803f
C74 plus.t5 a_n1670_n2088# 0.188565f
C75 plus.t3 a_n1670_n2088# 0.188565f
C76 plus.t9 a_n1670_n2088# 0.188565f
C77 plus.n20 a_n1670_n2088# 0.092222f
C78 plus.n21 a_n1670_n2088# 0.055152f
C79 plus.t4 a_n1670_n2088# 0.188565f
C80 plus.t8 a_n1670_n2088# 0.188565f
C81 plus.t11 a_n1670_n2088# 0.188565f
C82 plus.n22 a_n1670_n2088# 0.092222f
C83 plus.t10 a_n1670_n2088# 0.193803f
C84 plus.n23 a_n1670_n2088# 0.108251f
C85 plus.n24 a_n1670_n2088# 0.124164f
C86 plus.n25 a_n1670_n2088# 0.019316f
C87 plus.n26 a_n1670_n2088# 0.092222f
C88 plus.n27 a_n1670_n2088# 0.019316f
C89 plus.n28 a_n1670_n2088# 0.092222f
C90 plus.n29 a_n1670_n2088# 0.019316f
C91 plus.n30 a_n1670_n2088# 0.055152f
C92 plus.n31 a_n1670_n2088# 0.055152f
C93 plus.n32 a_n1670_n2088# 0.019316f
C94 plus.n33 a_n1670_n2088# 0.092222f
C95 plus.n34 a_n1670_n2088# 0.019316f
C96 plus.n35 a_n1670_n2088# 0.092222f
C97 plus.n36 a_n1670_n2088# 0.10817f
C98 plus.n37 a_n1670_n2088# 1.35855f
C99 source.n0 a_n1670_n2088# 0.046514f
C100 source.n1 a_n1670_n2088# 0.033092f
C101 source.n2 a_n1670_n2088# 0.017782f
C102 source.n3 a_n1670_n2088# 0.042031f
C103 source.n4 a_n1670_n2088# 0.018828f
C104 source.n5 a_n1670_n2088# 0.033092f
C105 source.n6 a_n1670_n2088# 0.017782f
C106 source.n7 a_n1670_n2088# 0.042031f
C107 source.n8 a_n1670_n2088# 0.018828f
C108 source.n9 a_n1670_n2088# 0.141611f
C109 source.t2 a_n1670_n2088# 0.068505f
C110 source.n10 a_n1670_n2088# 0.031523f
C111 source.n11 a_n1670_n2088# 0.024827f
C112 source.n12 a_n1670_n2088# 0.017782f
C113 source.n13 a_n1670_n2088# 0.787395f
C114 source.n14 a_n1670_n2088# 0.033092f
C115 source.n15 a_n1670_n2088# 0.017782f
C116 source.n16 a_n1670_n2088# 0.018828f
C117 source.n17 a_n1670_n2088# 0.042031f
C118 source.n18 a_n1670_n2088# 0.042031f
C119 source.n19 a_n1670_n2088# 0.018828f
C120 source.n20 a_n1670_n2088# 0.017782f
C121 source.n21 a_n1670_n2088# 0.033092f
C122 source.n22 a_n1670_n2088# 0.033092f
C123 source.n23 a_n1670_n2088# 0.017782f
C124 source.n24 a_n1670_n2088# 0.018828f
C125 source.n25 a_n1670_n2088# 0.042031f
C126 source.n26 a_n1670_n2088# 0.09099f
C127 source.n27 a_n1670_n2088# 0.018828f
C128 source.n28 a_n1670_n2088# 0.017782f
C129 source.n29 a_n1670_n2088# 0.076491f
C130 source.n30 a_n1670_n2088# 0.050912f
C131 source.n31 a_n1670_n2088# 0.78579f
C132 source.t12 a_n1670_n2088# 0.156902f
C133 source.t4 a_n1670_n2088# 0.156902f
C134 source.n32 a_n1670_n2088# 1.22197f
C135 source.n33 a_n1670_n2088# 0.407645f
C136 source.t9 a_n1670_n2088# 0.156902f
C137 source.t3 a_n1670_n2088# 0.156902f
C138 source.n34 a_n1670_n2088# 1.22197f
C139 source.n35 a_n1670_n2088# 0.407645f
C140 source.t15 a_n1670_n2088# 0.156902f
C141 source.t10 a_n1670_n2088# 0.156902f
C142 source.n36 a_n1670_n2088# 1.22197f
C143 source.n37 a_n1670_n2088# 0.407645f
C144 source.n38 a_n1670_n2088# 0.046514f
C145 source.n39 a_n1670_n2088# 0.033092f
C146 source.n40 a_n1670_n2088# 0.017782f
C147 source.n41 a_n1670_n2088# 0.042031f
C148 source.n42 a_n1670_n2088# 0.018828f
C149 source.n43 a_n1670_n2088# 0.033092f
C150 source.n44 a_n1670_n2088# 0.017782f
C151 source.n45 a_n1670_n2088# 0.042031f
C152 source.n46 a_n1670_n2088# 0.018828f
C153 source.n47 a_n1670_n2088# 0.141611f
C154 source.t0 a_n1670_n2088# 0.068505f
C155 source.n48 a_n1670_n2088# 0.031523f
C156 source.n49 a_n1670_n2088# 0.024827f
C157 source.n50 a_n1670_n2088# 0.017782f
C158 source.n51 a_n1670_n2088# 0.787395f
C159 source.n52 a_n1670_n2088# 0.033092f
C160 source.n53 a_n1670_n2088# 0.017782f
C161 source.n54 a_n1670_n2088# 0.018828f
C162 source.n55 a_n1670_n2088# 0.042031f
C163 source.n56 a_n1670_n2088# 0.042031f
C164 source.n57 a_n1670_n2088# 0.018828f
C165 source.n58 a_n1670_n2088# 0.017782f
C166 source.n59 a_n1670_n2088# 0.033092f
C167 source.n60 a_n1670_n2088# 0.033092f
C168 source.n61 a_n1670_n2088# 0.017782f
C169 source.n62 a_n1670_n2088# 0.018828f
C170 source.n63 a_n1670_n2088# 0.042031f
C171 source.n64 a_n1670_n2088# 0.09099f
C172 source.n65 a_n1670_n2088# 0.018828f
C173 source.n66 a_n1670_n2088# 0.017782f
C174 source.n67 a_n1670_n2088# 0.076491f
C175 source.n68 a_n1670_n2088# 0.050912f
C176 source.n69 a_n1670_n2088# 0.12708f
C177 source.n70 a_n1670_n2088# 0.046514f
C178 source.n71 a_n1670_n2088# 0.033092f
C179 source.n72 a_n1670_n2088# 0.017782f
C180 source.n73 a_n1670_n2088# 0.042031f
C181 source.n74 a_n1670_n2088# 0.018828f
C182 source.n75 a_n1670_n2088# 0.033092f
C183 source.n76 a_n1670_n2088# 0.017782f
C184 source.n77 a_n1670_n2088# 0.042031f
C185 source.n78 a_n1670_n2088# 0.018828f
C186 source.n79 a_n1670_n2088# 0.141611f
C187 source.t25 a_n1670_n2088# 0.068505f
C188 source.n80 a_n1670_n2088# 0.031523f
C189 source.n81 a_n1670_n2088# 0.024827f
C190 source.n82 a_n1670_n2088# 0.017782f
C191 source.n83 a_n1670_n2088# 0.787395f
C192 source.n84 a_n1670_n2088# 0.033092f
C193 source.n85 a_n1670_n2088# 0.017782f
C194 source.n86 a_n1670_n2088# 0.018828f
C195 source.n87 a_n1670_n2088# 0.042031f
C196 source.n88 a_n1670_n2088# 0.042031f
C197 source.n89 a_n1670_n2088# 0.018828f
C198 source.n90 a_n1670_n2088# 0.017782f
C199 source.n91 a_n1670_n2088# 0.033092f
C200 source.n92 a_n1670_n2088# 0.033092f
C201 source.n93 a_n1670_n2088# 0.017782f
C202 source.n94 a_n1670_n2088# 0.018828f
C203 source.n95 a_n1670_n2088# 0.042031f
C204 source.n96 a_n1670_n2088# 0.09099f
C205 source.n97 a_n1670_n2088# 0.018828f
C206 source.n98 a_n1670_n2088# 0.017782f
C207 source.n99 a_n1670_n2088# 0.076491f
C208 source.n100 a_n1670_n2088# 0.050912f
C209 source.n101 a_n1670_n2088# 0.12708f
C210 source.t30 a_n1670_n2088# 0.156902f
C211 source.t26 a_n1670_n2088# 0.156902f
C212 source.n102 a_n1670_n2088# 1.22197f
C213 source.n103 a_n1670_n2088# 0.407645f
C214 source.t24 a_n1670_n2088# 0.156902f
C215 source.t21 a_n1670_n2088# 0.156902f
C216 source.n104 a_n1670_n2088# 1.22197f
C217 source.n105 a_n1670_n2088# 0.407645f
C218 source.t29 a_n1670_n2088# 0.156902f
C219 source.t27 a_n1670_n2088# 0.156902f
C220 source.n106 a_n1670_n2088# 1.22197f
C221 source.n107 a_n1670_n2088# 0.407645f
C222 source.n108 a_n1670_n2088# 0.046514f
C223 source.n109 a_n1670_n2088# 0.033092f
C224 source.n110 a_n1670_n2088# 0.017782f
C225 source.n111 a_n1670_n2088# 0.042031f
C226 source.n112 a_n1670_n2088# 0.018828f
C227 source.n113 a_n1670_n2088# 0.033092f
C228 source.n114 a_n1670_n2088# 0.017782f
C229 source.n115 a_n1670_n2088# 0.042031f
C230 source.n116 a_n1670_n2088# 0.018828f
C231 source.n117 a_n1670_n2088# 0.141611f
C232 source.t20 a_n1670_n2088# 0.068505f
C233 source.n118 a_n1670_n2088# 0.031523f
C234 source.n119 a_n1670_n2088# 0.024827f
C235 source.n120 a_n1670_n2088# 0.017782f
C236 source.n121 a_n1670_n2088# 0.787395f
C237 source.n122 a_n1670_n2088# 0.033092f
C238 source.n123 a_n1670_n2088# 0.017782f
C239 source.n124 a_n1670_n2088# 0.018828f
C240 source.n125 a_n1670_n2088# 0.042031f
C241 source.n126 a_n1670_n2088# 0.042031f
C242 source.n127 a_n1670_n2088# 0.018828f
C243 source.n128 a_n1670_n2088# 0.017782f
C244 source.n129 a_n1670_n2088# 0.033092f
C245 source.n130 a_n1670_n2088# 0.033092f
C246 source.n131 a_n1670_n2088# 0.017782f
C247 source.n132 a_n1670_n2088# 0.018828f
C248 source.n133 a_n1670_n2088# 0.042031f
C249 source.n134 a_n1670_n2088# 0.09099f
C250 source.n135 a_n1670_n2088# 0.018828f
C251 source.n136 a_n1670_n2088# 0.017782f
C252 source.n137 a_n1670_n2088# 0.076491f
C253 source.n138 a_n1670_n2088# 0.050912f
C254 source.n139 a_n1670_n2088# 1.2092f
C255 source.n140 a_n1670_n2088# 0.046514f
C256 source.n141 a_n1670_n2088# 0.033092f
C257 source.n142 a_n1670_n2088# 0.017782f
C258 source.n143 a_n1670_n2088# 0.042031f
C259 source.n144 a_n1670_n2088# 0.018828f
C260 source.n145 a_n1670_n2088# 0.033092f
C261 source.n146 a_n1670_n2088# 0.017782f
C262 source.n147 a_n1670_n2088# 0.042031f
C263 source.n148 a_n1670_n2088# 0.018828f
C264 source.n149 a_n1670_n2088# 0.141611f
C265 source.t14 a_n1670_n2088# 0.068505f
C266 source.n150 a_n1670_n2088# 0.031523f
C267 source.n151 a_n1670_n2088# 0.024827f
C268 source.n152 a_n1670_n2088# 0.017782f
C269 source.n153 a_n1670_n2088# 0.787395f
C270 source.n154 a_n1670_n2088# 0.033092f
C271 source.n155 a_n1670_n2088# 0.017782f
C272 source.n156 a_n1670_n2088# 0.018828f
C273 source.n157 a_n1670_n2088# 0.042031f
C274 source.n158 a_n1670_n2088# 0.042031f
C275 source.n159 a_n1670_n2088# 0.018828f
C276 source.n160 a_n1670_n2088# 0.017782f
C277 source.n161 a_n1670_n2088# 0.033092f
C278 source.n162 a_n1670_n2088# 0.033092f
C279 source.n163 a_n1670_n2088# 0.017782f
C280 source.n164 a_n1670_n2088# 0.018828f
C281 source.n165 a_n1670_n2088# 0.042031f
C282 source.n166 a_n1670_n2088# 0.09099f
C283 source.n167 a_n1670_n2088# 0.018828f
C284 source.n168 a_n1670_n2088# 0.017782f
C285 source.n169 a_n1670_n2088# 0.076491f
C286 source.n170 a_n1670_n2088# 0.050912f
C287 source.n171 a_n1670_n2088# 1.2092f
C288 source.t7 a_n1670_n2088# 0.156902f
C289 source.t6 a_n1670_n2088# 0.156902f
C290 source.n172 a_n1670_n2088# 1.22196f
C291 source.n173 a_n1670_n2088# 0.407653f
C292 source.t1 a_n1670_n2088# 0.156902f
C293 source.t5 a_n1670_n2088# 0.156902f
C294 source.n174 a_n1670_n2088# 1.22196f
C295 source.n175 a_n1670_n2088# 0.407653f
C296 source.t13 a_n1670_n2088# 0.156902f
C297 source.t11 a_n1670_n2088# 0.156902f
C298 source.n176 a_n1670_n2088# 1.22196f
C299 source.n177 a_n1670_n2088# 0.407653f
C300 source.n178 a_n1670_n2088# 0.046514f
C301 source.n179 a_n1670_n2088# 0.033092f
C302 source.n180 a_n1670_n2088# 0.017782f
C303 source.n181 a_n1670_n2088# 0.042031f
C304 source.n182 a_n1670_n2088# 0.018828f
C305 source.n183 a_n1670_n2088# 0.033092f
C306 source.n184 a_n1670_n2088# 0.017782f
C307 source.n185 a_n1670_n2088# 0.042031f
C308 source.n186 a_n1670_n2088# 0.018828f
C309 source.n187 a_n1670_n2088# 0.141611f
C310 source.t8 a_n1670_n2088# 0.068505f
C311 source.n188 a_n1670_n2088# 0.031523f
C312 source.n189 a_n1670_n2088# 0.024827f
C313 source.n190 a_n1670_n2088# 0.017782f
C314 source.n191 a_n1670_n2088# 0.787395f
C315 source.n192 a_n1670_n2088# 0.033092f
C316 source.n193 a_n1670_n2088# 0.017782f
C317 source.n194 a_n1670_n2088# 0.018828f
C318 source.n195 a_n1670_n2088# 0.042031f
C319 source.n196 a_n1670_n2088# 0.042031f
C320 source.n197 a_n1670_n2088# 0.018828f
C321 source.n198 a_n1670_n2088# 0.017782f
C322 source.n199 a_n1670_n2088# 0.033092f
C323 source.n200 a_n1670_n2088# 0.033092f
C324 source.n201 a_n1670_n2088# 0.017782f
C325 source.n202 a_n1670_n2088# 0.018828f
C326 source.n203 a_n1670_n2088# 0.042031f
C327 source.n204 a_n1670_n2088# 0.09099f
C328 source.n205 a_n1670_n2088# 0.018828f
C329 source.n206 a_n1670_n2088# 0.017782f
C330 source.n207 a_n1670_n2088# 0.076491f
C331 source.n208 a_n1670_n2088# 0.050912f
C332 source.n209 a_n1670_n2088# 0.12708f
C333 source.n210 a_n1670_n2088# 0.046514f
C334 source.n211 a_n1670_n2088# 0.033092f
C335 source.n212 a_n1670_n2088# 0.017782f
C336 source.n213 a_n1670_n2088# 0.042031f
C337 source.n214 a_n1670_n2088# 0.018828f
C338 source.n215 a_n1670_n2088# 0.033092f
C339 source.n216 a_n1670_n2088# 0.017782f
C340 source.n217 a_n1670_n2088# 0.042031f
C341 source.n218 a_n1670_n2088# 0.018828f
C342 source.n219 a_n1670_n2088# 0.141611f
C343 source.t22 a_n1670_n2088# 0.068505f
C344 source.n220 a_n1670_n2088# 0.031523f
C345 source.n221 a_n1670_n2088# 0.024827f
C346 source.n222 a_n1670_n2088# 0.017782f
C347 source.n223 a_n1670_n2088# 0.787395f
C348 source.n224 a_n1670_n2088# 0.033092f
C349 source.n225 a_n1670_n2088# 0.017782f
C350 source.n226 a_n1670_n2088# 0.018828f
C351 source.n227 a_n1670_n2088# 0.042031f
C352 source.n228 a_n1670_n2088# 0.042031f
C353 source.n229 a_n1670_n2088# 0.018828f
C354 source.n230 a_n1670_n2088# 0.017782f
C355 source.n231 a_n1670_n2088# 0.033092f
C356 source.n232 a_n1670_n2088# 0.033092f
C357 source.n233 a_n1670_n2088# 0.017782f
C358 source.n234 a_n1670_n2088# 0.018828f
C359 source.n235 a_n1670_n2088# 0.042031f
C360 source.n236 a_n1670_n2088# 0.09099f
C361 source.n237 a_n1670_n2088# 0.018828f
C362 source.n238 a_n1670_n2088# 0.017782f
C363 source.n239 a_n1670_n2088# 0.076491f
C364 source.n240 a_n1670_n2088# 0.050912f
C365 source.n241 a_n1670_n2088# 0.12708f
C366 source.t18 a_n1670_n2088# 0.156902f
C367 source.t23 a_n1670_n2088# 0.156902f
C368 source.n242 a_n1670_n2088# 1.22196f
C369 source.n243 a_n1670_n2088# 0.407653f
C370 source.t19 a_n1670_n2088# 0.156902f
C371 source.t28 a_n1670_n2088# 0.156902f
C372 source.n244 a_n1670_n2088# 1.22196f
C373 source.n245 a_n1670_n2088# 0.407653f
C374 source.t16 a_n1670_n2088# 0.156902f
C375 source.t31 a_n1670_n2088# 0.156902f
C376 source.n246 a_n1670_n2088# 1.22196f
C377 source.n247 a_n1670_n2088# 0.407653f
C378 source.n248 a_n1670_n2088# 0.046514f
C379 source.n249 a_n1670_n2088# 0.033092f
C380 source.n250 a_n1670_n2088# 0.017782f
C381 source.n251 a_n1670_n2088# 0.042031f
C382 source.n252 a_n1670_n2088# 0.018828f
C383 source.n253 a_n1670_n2088# 0.033092f
C384 source.n254 a_n1670_n2088# 0.017782f
C385 source.n255 a_n1670_n2088# 0.042031f
C386 source.n256 a_n1670_n2088# 0.018828f
C387 source.n257 a_n1670_n2088# 0.141611f
C388 source.t17 a_n1670_n2088# 0.068505f
C389 source.n258 a_n1670_n2088# 0.031523f
C390 source.n259 a_n1670_n2088# 0.024827f
C391 source.n260 a_n1670_n2088# 0.017782f
C392 source.n261 a_n1670_n2088# 0.787395f
C393 source.n262 a_n1670_n2088# 0.033092f
C394 source.n263 a_n1670_n2088# 0.017782f
C395 source.n264 a_n1670_n2088# 0.018828f
C396 source.n265 a_n1670_n2088# 0.042031f
C397 source.n266 a_n1670_n2088# 0.042031f
C398 source.n267 a_n1670_n2088# 0.018828f
C399 source.n268 a_n1670_n2088# 0.017782f
C400 source.n269 a_n1670_n2088# 0.033092f
C401 source.n270 a_n1670_n2088# 0.033092f
C402 source.n271 a_n1670_n2088# 0.017782f
C403 source.n272 a_n1670_n2088# 0.018828f
C404 source.n273 a_n1670_n2088# 0.042031f
C405 source.n274 a_n1670_n2088# 0.09099f
C406 source.n275 a_n1670_n2088# 0.018828f
C407 source.n276 a_n1670_n2088# 0.017782f
C408 source.n277 a_n1670_n2088# 0.076491f
C409 source.n278 a_n1670_n2088# 0.050912f
C410 source.n279 a_n1670_n2088# 0.306516f
C411 source.n280 a_n1670_n2088# 1.34963f
C412 drain_right.t13 a_n1670_n2088# 0.178331f
C413 drain_right.t11 a_n1670_n2088# 0.178331f
C414 drain_right.n0 a_n1670_n2088# 1.4902f
C415 drain_right.t14 a_n1670_n2088# 0.178331f
C416 drain_right.t15 a_n1670_n2088# 0.178331f
C417 drain_right.n1 a_n1670_n2088# 1.48729f
C418 drain_right.n2 a_n1670_n2088# 0.814911f
C419 drain_right.t1 a_n1670_n2088# 0.178331f
C420 drain_right.t9 a_n1670_n2088# 0.178331f
C421 drain_right.n3 a_n1670_n2088# 1.4902f
C422 drain_right.t7 a_n1670_n2088# 0.178331f
C423 drain_right.t4 a_n1670_n2088# 0.178331f
C424 drain_right.n4 a_n1670_n2088# 1.48729f
C425 drain_right.n5 a_n1670_n2088# 0.814911f
C426 drain_right.n6 a_n1670_n2088# 1.19782f
C427 drain_right.t2 a_n1670_n2088# 0.178331f
C428 drain_right.t0 a_n1670_n2088# 0.178331f
C429 drain_right.n7 a_n1670_n2088# 1.4902f
C430 drain_right.t12 a_n1670_n2088# 0.178331f
C431 drain_right.t10 a_n1670_n2088# 0.178331f
C432 drain_right.n8 a_n1670_n2088# 1.48729f
C433 drain_right.n9 a_n1670_n2088# 0.844261f
C434 drain_right.t3 a_n1670_n2088# 0.178331f
C435 drain_right.t6 a_n1670_n2088# 0.178331f
C436 drain_right.n10 a_n1670_n2088# 1.48729f
C437 drain_right.n11 a_n1670_n2088# 0.416009f
C438 drain_right.t5 a_n1670_n2088# 0.178331f
C439 drain_right.t8 a_n1670_n2088# 0.178331f
C440 drain_right.n12 a_n1670_n2088# 1.48729f
C441 drain_right.n13 a_n1670_n2088# 0.723825f
C442 minus.n0 a_n1670_n2088# 0.053886f
C443 minus.t11 a_n1670_n2088# 0.189353f
C444 minus.t2 a_n1670_n2088# 0.184235f
C445 minus.t4 a_n1670_n2088# 0.184235f
C446 minus.t7 a_n1670_n2088# 0.184235f
C447 minus.n1 a_n1670_n2088# 0.090104f
C448 minus.n2 a_n1670_n2088# 0.053886f
C449 minus.t10 a_n1670_n2088# 0.184235f
C450 minus.t1 a_n1670_n2088# 0.184235f
C451 minus.t5 a_n1670_n2088# 0.184235f
C452 minus.n3 a_n1670_n2088# 0.090104f
C453 minus.t6 a_n1670_n2088# 0.189353f
C454 minus.n4 a_n1670_n2088# 0.105766f
C455 minus.n5 a_n1670_n2088# 0.121313f
C456 minus.n6 a_n1670_n2088# 0.018872f
C457 minus.n7 a_n1670_n2088# 0.090104f
C458 minus.n8 a_n1670_n2088# 0.018872f
C459 minus.n9 a_n1670_n2088# 0.090104f
C460 minus.n10 a_n1670_n2088# 0.018872f
C461 minus.n11 a_n1670_n2088# 0.053886f
C462 minus.n12 a_n1670_n2088# 0.053886f
C463 minus.n13 a_n1670_n2088# 0.018872f
C464 minus.n14 a_n1670_n2088# 0.090104f
C465 minus.n15 a_n1670_n2088# 0.018872f
C466 minus.n16 a_n1670_n2088# 0.090104f
C467 minus.n17 a_n1670_n2088# 0.105686f
C468 minus.n18 a_n1670_n2088# 1.4696f
C469 minus.n19 a_n1670_n2088# 0.053886f
C470 minus.t0 a_n1670_n2088# 0.184235f
C471 minus.t15 a_n1670_n2088# 0.184235f
C472 minus.t3 a_n1670_n2088# 0.184235f
C473 minus.n20 a_n1670_n2088# 0.090104f
C474 minus.n21 a_n1670_n2088# 0.053886f
C475 minus.t12 a_n1670_n2088# 0.184235f
C476 minus.t8 a_n1670_n2088# 0.184235f
C477 minus.t13 a_n1670_n2088# 0.184235f
C478 minus.n22 a_n1670_n2088# 0.090104f
C479 minus.t9 a_n1670_n2088# 0.189353f
C480 minus.n23 a_n1670_n2088# 0.105766f
C481 minus.n24 a_n1670_n2088# 0.121313f
C482 minus.n25 a_n1670_n2088# 0.018872f
C483 minus.n26 a_n1670_n2088# 0.090104f
C484 minus.n27 a_n1670_n2088# 0.018872f
C485 minus.n28 a_n1670_n2088# 0.090104f
C486 minus.n29 a_n1670_n2088# 0.018872f
C487 minus.n30 a_n1670_n2088# 0.053886f
C488 minus.n31 a_n1670_n2088# 0.053886f
C489 minus.n32 a_n1670_n2088# 0.018872f
C490 minus.n33 a_n1670_n2088# 0.090104f
C491 minus.n34 a_n1670_n2088# 0.018872f
C492 minus.n35 a_n1670_n2088# 0.090104f
C493 minus.t14 a_n1670_n2088# 0.189353f
C494 minus.n36 a_n1670_n2088# 0.105686f
C495 minus.n37 a_n1670_n2088# 0.348019f
C496 minus.n38 a_n1670_n2088# 1.81218f
.ends

