* NGSPICE file created from diffpair646.ext - technology: sky130A

.subckt diffpair646 minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t9 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 drain_right.t8 minus.t1 source.t26 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X2 source.t0 plus.t0 drain_left.t13 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X3 a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X4 a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X5 drain_left.t12 plus.t1 source.t1 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X6 a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X7 drain_left.t11 plus.t2 source.t3 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X8 a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X9 source.t25 minus.t2 drain_right.t13 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X10 source.t6 plus.t3 drain_left.t10 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X11 drain_right.t12 minus.t3 source.t24 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X12 drain_right.t11 minus.t4 source.t23 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X13 drain_right.t10 minus.t5 source.t22 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X14 drain_left.t9 plus.t4 source.t8 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X15 source.t21 minus.t6 drain_right.t1 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X16 drain_left.t8 plus.t5 source.t7 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 drain_left.t7 plus.t6 source.t13 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X18 drain_right.t0 minus.t7 source.t20 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 drain_right.t7 minus.t8 source.t19 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X20 source.t18 minus.t9 drain_right.t6 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X21 source.t5 plus.t7 drain_left.t6 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 source.t17 minus.t10 drain_right.t3 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X23 source.t16 minus.t11 drain_right.t2 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X24 source.t9 plus.t8 drain_left.t5 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X25 drain_left.t4 plus.t9 source.t11 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X26 drain_left.t3 plus.t10 source.t2 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X27 source.t10 plus.t11 drain_left.t2 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X28 source.t4 plus.t12 drain_left.t1 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X29 drain_right.t5 minus.t12 source.t15 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X30 drain_left.t0 plus.t13 source.t12 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X31 drain_right.t4 minus.t13 source.t14 a_n1756_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
R0 minus.n15 minus.t8 4291.26
R1 minus.n3 minus.t3 4291.26
R2 minus.n32 minus.t13 4291.26
R3 minus.n20 minus.t1 4291.26
R4 minus.n1 minus.t6 4225.53
R5 minus.n14 minus.t10 4225.53
R6 minus.n12 minus.t4 4225.53
R7 minus.n6 minus.t7 4225.53
R8 minus.n4 minus.t2 4225.53
R9 minus.n18 minus.t0 4225.53
R10 minus.n31 minus.t11 4225.53
R11 minus.n29 minus.t5 4225.53
R12 minus.n23 minus.t12 4225.53
R13 minus.n21 minus.t9 4225.53
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 51.1217
R33 minus.n6 minus.n5 51.1217
R34 minus.n23 minus.n22 51.1217
R35 minus.n30 minus.n29 51.1217
R36 minus.n34 minus.n16 45.6918
R37 minus.n14 minus.n13 43.8187
R38 minus.n5 minus.n4 43.8187
R39 minus.n22 minus.n21 43.8187
R40 minus.n31 minus.n30 43.8187
R41 minus.n15 minus.n14 29.2126
R42 minus.n4 minus.n3 29.2126
R43 minus.n21 minus.n20 29.2126
R44 minus.n32 minus.n31 29.2126
R45 minus.n12 minus.n11 21.9096
R46 minus.n7 minus.n6 21.9096
R47 minus.n24 minus.n23 21.9096
R48 minus.n29 minus.n28 21.9096
R49 minus.n34 minus.n33 6.57058
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n1 drain_right.t8 60.4756
R62 drain_right.n11 drain_right.t7 59.9154
R63 drain_right.n4 drain_right.n2 59.2758
R64 drain_right.n8 drain_right.n6 59.2756
R65 drain_right.n4 drain_right.n3 58.7154
R66 drain_right.n1 drain_right.n0 58.7154
R67 drain_right.n8 drain_right.n7 58.7154
R68 drain_right.n10 drain_right.n9 58.7154
R69 drain_right drain_right.n5 39.8843
R70 drain_right drain_right.n11 5.93339
R71 drain_right.n2 drain_right.t2 1.2005
R72 drain_right.n2 drain_right.t4 1.2005
R73 drain_right.n3 drain_right.t9 1.2005
R74 drain_right.n3 drain_right.t10 1.2005
R75 drain_right.n0 drain_right.t6 1.2005
R76 drain_right.n0 drain_right.t5 1.2005
R77 drain_right.n6 drain_right.t13 1.2005
R78 drain_right.n6 drain_right.t12 1.2005
R79 drain_right.n7 drain_right.t1 1.2005
R80 drain_right.n7 drain_right.t0 1.2005
R81 drain_right.n9 drain_right.t3 1.2005
R82 drain_right.n9 drain_right.t11 1.2005
R83 drain_right.n11 drain_right.n10 0.560845
R84 drain_right.n10 drain_right.n8 0.560845
R85 drain_right.n5 drain_right.n1 0.365413
R86 drain_right.n5 drain_right.n4 0.0852402
R87 source.n7 source.t24 43.2366
R88 source.n27 source.t14 43.2365
R89 source.n20 source.t8 43.2365
R90 source.n0 source.t11 43.2365
R91 source.n26 source.n25 42.0366
R92 source.n24 source.n23 42.0366
R93 source.n22 source.n21 42.0366
R94 source.n19 source.n18 42.0366
R95 source.n17 source.n16 42.0366
R96 source.n15 source.n14 42.0366
R97 source.n2 source.n1 42.0366
R98 source.n4 source.n3 42.0366
R99 source.n6 source.n5 42.0366
R100 source.n9 source.n8 42.0366
R101 source.n11 source.n10 42.0366
R102 source.n13 source.n12 42.0366
R103 source.n15 source.n13 32.2569
R104 source.n28 source.n0 26.1535
R105 source.n28 source.n27 5.5436
R106 source.n25 source.t22 1.2005
R107 source.n25 source.t16 1.2005
R108 source.n23 source.t15 1.2005
R109 source.n23 source.t27 1.2005
R110 source.n21 source.t26 1.2005
R111 source.n21 source.t18 1.2005
R112 source.n18 source.t1 1.2005
R113 source.n18 source.t9 1.2005
R114 source.n16 source.t7 1.2005
R115 source.n16 source.t6 1.2005
R116 source.n14 source.t3 1.2005
R117 source.n14 source.t0 1.2005
R118 source.n1 source.t12 1.2005
R119 source.n1 source.t10 1.2005
R120 source.n3 source.t2 1.2005
R121 source.n3 source.t5 1.2005
R122 source.n5 source.t13 1.2005
R123 source.n5 source.t4 1.2005
R124 source.n8 source.t20 1.2005
R125 source.n8 source.t25 1.2005
R126 source.n10 source.t23 1.2005
R127 source.n10 source.t21 1.2005
R128 source.n12 source.t19 1.2005
R129 source.n12 source.t17 1.2005
R130 source.n7 source.n6 0.7505
R131 source.n22 source.n20 0.7505
R132 source.n13 source.n11 0.560845
R133 source.n11 source.n9 0.560845
R134 source.n9 source.n7 0.560845
R135 source.n6 source.n4 0.560845
R136 source.n4 source.n2 0.560845
R137 source.n2 source.n0 0.560845
R138 source.n17 source.n15 0.560845
R139 source.n19 source.n17 0.560845
R140 source.n20 source.n19 0.560845
R141 source.n24 source.n22 0.560845
R142 source.n26 source.n24 0.560845
R143 source.n27 source.n26 0.560845
R144 source source.n28 0.188
R145 plus.n3 plus.t6 4291.26
R146 plus.n15 plus.t9 4291.26
R147 plus.n20 plus.t4 4291.26
R148 plus.n32 plus.t2 4291.26
R149 plus.n1 plus.t7 4225.53
R150 plus.n4 plus.t12 4225.53
R151 plus.n6 plus.t10 4225.53
R152 plus.n12 plus.t13 4225.53
R153 plus.n14 plus.t11 4225.53
R154 plus.n18 plus.t3 4225.53
R155 plus.n21 plus.t8 4225.53
R156 plus.n23 plus.t1 4225.53
R157 plus.n29 plus.t5 4225.53
R158 plus.n31 plus.t0 4225.53
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 51.1217
R178 plus.n13 plus.n12 51.1217
R179 plus.n30 plus.n29 51.1217
R180 plus.n23 plus.n22 51.1217
R181 plus.n5 plus.n4 43.8187
R182 plus.n14 plus.n13 43.8187
R183 plus.n31 plus.n30 43.8187
R184 plus.n22 plus.n21 43.8187
R185 plus plus.n33 34.6486
R186 plus.n4 plus.n3 29.2126
R187 plus.n15 plus.n14 29.2126
R188 plus.n32 plus.n31 29.2126
R189 plus.n21 plus.n20 29.2126
R190 plus.n7 plus.n6 21.9096
R191 plus.n12 plus.n11 21.9096
R192 plus.n29 plus.n28 21.9096
R193 plus.n24 plus.n23 21.9096
R194 plus plus.n16 17.1388
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t7 60.4758
R206 drain_left.n1 drain_left.t11 60.4756
R207 drain_left.n4 drain_left.n2 59.2758
R208 drain_left.n4 drain_left.n3 58.7154
R209 drain_left.n1 drain_left.n0 58.7154
R210 drain_left.n9 drain_left.n8 58.7154
R211 drain_left.n7 drain_left.n6 58.7154
R212 drain_left.n11 drain_left.n10 58.7153
R213 drain_left drain_left.n5 40.4375
R214 drain_left drain_left.n11 6.21356
R215 drain_left.n2 drain_left.t5 1.2005
R216 drain_left.n2 drain_left.t9 1.2005
R217 drain_left.n3 drain_left.t10 1.2005
R218 drain_left.n3 drain_left.t12 1.2005
R219 drain_left.n0 drain_left.t13 1.2005
R220 drain_left.n0 drain_left.t8 1.2005
R221 drain_left.n10 drain_left.t2 1.2005
R222 drain_left.n10 drain_left.t4 1.2005
R223 drain_left.n8 drain_left.t6 1.2005
R224 drain_left.n8 drain_left.t0 1.2005
R225 drain_left.n6 drain_left.t1 1.2005
R226 drain_left.n6 drain_left.t3 1.2005
R227 drain_left.n9 drain_left.n7 0.560845
R228 drain_left.n11 drain_left.n9 0.560845
R229 drain_left.n5 drain_left.n1 0.365413
R230 drain_left.n5 drain_left.n4 0.0852402
C0 source drain_left 56.6125f
C1 plus minus 7.73138f
C2 drain_right minus 6.14735f
C3 plus drain_right 0.328442f
C4 source minus 5.02453f
C5 plus source 5.03991f
C6 source drain_right 56.591896f
C7 drain_left minus 0.171187f
C8 plus drain_left 6.3116f
C9 drain_left drain_right 0.906572f
C10 drain_right a_n1756_n5888# 10.57128f
C11 drain_left a_n1756_n5888# 10.84485f
C12 source a_n1756_n5888# 10.757905f
C13 minus a_n1756_n5888# 7.336607f
C14 plus a_n1756_n5888# 10.4395f
C15 drain_left.t11 a_n1756_n5888# 6.56173f
C16 drain_left.t13 a_n1756_n5888# 0.779689f
C17 drain_left.t8 a_n1756_n5888# 0.779689f
C18 drain_left.n0 a_n1756_n5888# 5.27273f
C19 drain_left.n1 a_n1756_n5888# 0.691636f
C20 drain_left.t5 a_n1756_n5888# 0.779689f
C21 drain_left.t9 a_n1756_n5888# 0.779689f
C22 drain_left.n2 a_n1756_n5888# 5.2758f
C23 drain_left.t10 a_n1756_n5888# 0.779689f
C24 drain_left.t12 a_n1756_n5888# 0.779689f
C25 drain_left.n3 a_n1756_n5888# 5.27273f
C26 drain_left.n4 a_n1756_n5888# 0.603113f
C27 drain_left.n5 a_n1756_n5888# 2.10338f
C28 drain_left.t7 a_n1756_n5888# 6.56174f
C29 drain_left.t1 a_n1756_n5888# 0.779689f
C30 drain_left.t3 a_n1756_n5888# 0.779689f
C31 drain_left.n6 a_n1756_n5888# 5.27273f
C32 drain_left.n7 a_n1756_n5888# 0.706371f
C33 drain_left.t6 a_n1756_n5888# 0.779689f
C34 drain_left.t0 a_n1756_n5888# 0.779689f
C35 drain_left.n8 a_n1756_n5888# 5.27273f
C36 drain_left.n9 a_n1756_n5888# 0.31424f
C37 drain_left.t2 a_n1756_n5888# 0.779689f
C38 drain_left.t4 a_n1756_n5888# 0.779689f
C39 drain_left.n10 a_n1756_n5888# 5.27272f
C40 drain_left.n11 a_n1756_n5888# 0.531779f
C41 plus.n0 a_n1756_n5888# 0.056397f
C42 plus.t11 a_n1756_n5888# 0.59506f
C43 plus.t13 a_n1756_n5888# 0.59506f
C44 plus.t7 a_n1756_n5888# 0.59506f
C45 plus.n1 a_n1756_n5888# 0.243931f
C46 plus.n2 a_n1756_n5888# 0.131829f
C47 plus.t10 a_n1756_n5888# 0.59506f
C48 plus.t12 a_n1756_n5888# 0.59506f
C49 plus.t6 a_n1756_n5888# 0.598563f
C50 plus.n3 a_n1756_n5888# 0.249209f
C51 plus.n4 a_n1756_n5888# 0.225222f
C52 plus.n5 a_n1756_n5888# 0.023924f
C53 plus.n6 a_n1756_n5888# 0.225222f
C54 plus.n7 a_n1756_n5888# 0.023924f
C55 plus.n8 a_n1756_n5888# 0.056397f
C56 plus.n9 a_n1756_n5888# 0.056397f
C57 plus.n10 a_n1756_n5888# 0.056397f
C58 plus.n11 a_n1756_n5888# 0.023924f
C59 plus.n12 a_n1756_n5888# 0.225222f
C60 plus.n13 a_n1756_n5888# 0.023924f
C61 plus.n14 a_n1756_n5888# 0.225222f
C62 plus.t9 a_n1756_n5888# 0.598563f
C63 plus.n15 a_n1756_n5888# 0.249121f
C64 plus.n16 a_n1756_n5888# 1.01566f
C65 plus.n17 a_n1756_n5888# 0.056397f
C66 plus.t2 a_n1756_n5888# 0.598563f
C67 plus.t0 a_n1756_n5888# 0.59506f
C68 plus.t5 a_n1756_n5888# 0.59506f
C69 plus.t3 a_n1756_n5888# 0.59506f
C70 plus.n18 a_n1756_n5888# 0.243931f
C71 plus.n19 a_n1756_n5888# 0.131829f
C72 plus.t1 a_n1756_n5888# 0.59506f
C73 plus.t8 a_n1756_n5888# 0.59506f
C74 plus.t4 a_n1756_n5888# 0.598563f
C75 plus.n20 a_n1756_n5888# 0.249209f
C76 plus.n21 a_n1756_n5888# 0.225222f
C77 plus.n22 a_n1756_n5888# 0.023924f
C78 plus.n23 a_n1756_n5888# 0.225222f
C79 plus.n24 a_n1756_n5888# 0.023924f
C80 plus.n25 a_n1756_n5888# 0.056397f
C81 plus.n26 a_n1756_n5888# 0.056397f
C82 plus.n27 a_n1756_n5888# 0.056397f
C83 plus.n28 a_n1756_n5888# 0.023924f
C84 plus.n29 a_n1756_n5888# 0.225222f
C85 plus.n30 a_n1756_n5888# 0.023924f
C86 plus.n31 a_n1756_n5888# 0.225222f
C87 plus.n32 a_n1756_n5888# 0.249121f
C88 plus.n33 a_n1756_n5888# 2.15981f
C89 source.t11 a_n1756_n5888# 6.437819f
C90 source.n0 a_n1756_n5888# 2.46341f
C91 source.t12 a_n1756_n5888# 0.7807f
C92 source.t10 a_n1756_n5888# 0.7807f
C93 source.n1 a_n1756_n5888# 5.19407f
C94 source.n2 a_n1756_n5888# 0.364702f
C95 source.t2 a_n1756_n5888# 0.7807f
C96 source.t5 a_n1756_n5888# 0.7807f
C97 source.n3 a_n1756_n5888# 5.19407f
C98 source.n4 a_n1756_n5888# 0.364702f
C99 source.t13 a_n1756_n5888# 0.7807f
C100 source.t4 a_n1756_n5888# 0.7807f
C101 source.n5 a_n1756_n5888# 5.19407f
C102 source.n6 a_n1756_n5888# 0.38064f
C103 source.t24 a_n1756_n5888# 6.43784f
C104 source.n7 a_n1756_n5888# 0.542134f
C105 source.t20 a_n1756_n5888# 0.7807f
C106 source.t25 a_n1756_n5888# 0.7807f
C107 source.n8 a_n1756_n5888# 5.19407f
C108 source.n9 a_n1756_n5888# 0.364702f
C109 source.t23 a_n1756_n5888# 0.7807f
C110 source.t21 a_n1756_n5888# 0.7807f
C111 source.n10 a_n1756_n5888# 5.19407f
C112 source.n11 a_n1756_n5888# 0.364702f
C113 source.t19 a_n1756_n5888# 0.7807f
C114 source.t17 a_n1756_n5888# 0.7807f
C115 source.n12 a_n1756_n5888# 5.19407f
C116 source.n13 a_n1756_n5888# 2.83215f
C117 source.t3 a_n1756_n5888# 0.7807f
C118 source.t0 a_n1756_n5888# 0.7807f
C119 source.n14 a_n1756_n5888# 5.19407f
C120 source.n15 a_n1756_n5888# 2.83215f
C121 source.t7 a_n1756_n5888# 0.7807f
C122 source.t6 a_n1756_n5888# 0.7807f
C123 source.n16 a_n1756_n5888# 5.19407f
C124 source.n17 a_n1756_n5888# 0.364703f
C125 source.t1 a_n1756_n5888# 0.7807f
C126 source.t9 a_n1756_n5888# 0.7807f
C127 source.n18 a_n1756_n5888# 5.19407f
C128 source.n19 a_n1756_n5888# 0.364703f
C129 source.t8 a_n1756_n5888# 6.437819f
C130 source.n20 a_n1756_n5888# 0.542151f
C131 source.t26 a_n1756_n5888# 0.7807f
C132 source.t18 a_n1756_n5888# 0.7807f
C133 source.n21 a_n1756_n5888# 5.19407f
C134 source.n22 a_n1756_n5888# 0.380642f
C135 source.t15 a_n1756_n5888# 0.7807f
C136 source.t27 a_n1756_n5888# 0.7807f
C137 source.n23 a_n1756_n5888# 5.19407f
C138 source.n24 a_n1756_n5888# 0.364703f
C139 source.t22 a_n1756_n5888# 0.7807f
C140 source.t16 a_n1756_n5888# 0.7807f
C141 source.n25 a_n1756_n5888# 5.19407f
C142 source.n26 a_n1756_n5888# 0.364703f
C143 source.t14 a_n1756_n5888# 6.437819f
C144 source.n27 a_n1756_n5888# 0.666993f
C145 source.n28 a_n1756_n5888# 2.78128f
C146 drain_right.t8 a_n1756_n5888# 6.55148f
C147 drain_right.t6 a_n1756_n5888# 0.778471f
C148 drain_right.t5 a_n1756_n5888# 0.778471f
C149 drain_right.n0 a_n1756_n5888# 5.2645f
C150 drain_right.n1 a_n1756_n5888# 0.690555f
C151 drain_right.t2 a_n1756_n5888# 0.778471f
C152 drain_right.t4 a_n1756_n5888# 0.778471f
C153 drain_right.n2 a_n1756_n5888# 5.26756f
C154 drain_right.t9 a_n1756_n5888# 0.778471f
C155 drain_right.t10 a_n1756_n5888# 0.778471f
C156 drain_right.n3 a_n1756_n5888# 5.2645f
C157 drain_right.n4 a_n1756_n5888# 0.60217f
C158 drain_right.n5 a_n1756_n5888# 2.04611f
C159 drain_right.t13 a_n1756_n5888# 0.778471f
C160 drain_right.t12 a_n1756_n5888# 0.778471f
C161 drain_right.n6 a_n1756_n5888# 5.26755f
C162 drain_right.t1 a_n1756_n5888# 0.778471f
C163 drain_right.t0 a_n1756_n5888# 0.778471f
C164 drain_right.n7 a_n1756_n5888# 5.2645f
C165 drain_right.n8 a_n1756_n5888# 0.63492f
C166 drain_right.t3 a_n1756_n5888# 0.778471f
C167 drain_right.t11 a_n1756_n5888# 0.778471f
C168 drain_right.n9 a_n1756_n5888# 5.2645f
C169 drain_right.n10 a_n1756_n5888# 0.313749f
C170 drain_right.t7 a_n1756_n5888# 6.54783f
C171 drain_right.n11 a_n1756_n5888# 0.613257f
C172 minus.n0 a_n1756_n5888# 0.05547f
C173 minus.t8 a_n1756_n5888# 0.588729f
C174 minus.t10 a_n1756_n5888# 0.585284f
C175 minus.t4 a_n1756_n5888# 0.585284f
C176 minus.t6 a_n1756_n5888# 0.585284f
C177 minus.n1 a_n1756_n5888# 0.239923f
C178 minus.n2 a_n1756_n5888# 0.129663f
C179 minus.t7 a_n1756_n5888# 0.585284f
C180 minus.t2 a_n1756_n5888# 0.585284f
C181 minus.t3 a_n1756_n5888# 0.588729f
C182 minus.n3 a_n1756_n5888# 0.245115f
C183 minus.n4 a_n1756_n5888# 0.221522f
C184 minus.n5 a_n1756_n5888# 0.023531f
C185 minus.n6 a_n1756_n5888# 0.221522f
C186 minus.n7 a_n1756_n5888# 0.023531f
C187 minus.n8 a_n1756_n5888# 0.05547f
C188 minus.n9 a_n1756_n5888# 0.05547f
C189 minus.n10 a_n1756_n5888# 0.05547f
C190 minus.n11 a_n1756_n5888# 0.023531f
C191 minus.n12 a_n1756_n5888# 0.221522f
C192 minus.n13 a_n1756_n5888# 0.023531f
C193 minus.n14 a_n1756_n5888# 0.221522f
C194 minus.n15 a_n1756_n5888# 0.245028f
C195 minus.n16 a_n1756_n5888# 2.77818f
C196 minus.n17 a_n1756_n5888# 0.05547f
C197 minus.t11 a_n1756_n5888# 0.585284f
C198 minus.t5 a_n1756_n5888# 0.585284f
C199 minus.t0 a_n1756_n5888# 0.585284f
C200 minus.n18 a_n1756_n5888# 0.239923f
C201 minus.n19 a_n1756_n5888# 0.129663f
C202 minus.t12 a_n1756_n5888# 0.585284f
C203 minus.t9 a_n1756_n5888# 0.585284f
C204 minus.t1 a_n1756_n5888# 0.588729f
C205 minus.n20 a_n1756_n5888# 0.245115f
C206 minus.n21 a_n1756_n5888# 0.221522f
C207 minus.n22 a_n1756_n5888# 0.023531f
C208 minus.n23 a_n1756_n5888# 0.221522f
C209 minus.n24 a_n1756_n5888# 0.023531f
C210 minus.n25 a_n1756_n5888# 0.05547f
C211 minus.n26 a_n1756_n5888# 0.05547f
C212 minus.n27 a_n1756_n5888# 0.05547f
C213 minus.n28 a_n1756_n5888# 0.023531f
C214 minus.n29 a_n1756_n5888# 0.221522f
C215 minus.n30 a_n1756_n5888# 0.023531f
C216 minus.n31 a_n1756_n5888# 0.221522f
C217 minus.t13 a_n1756_n5888# 0.588729f
C218 minus.n32 a_n1756_n5888# 0.245028f
C219 minus.n33 a_n1756_n5888# 0.371843f
C220 minus.n34 a_n1756_n5888# 3.28216f
.ends

