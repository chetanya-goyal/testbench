* NGSPICE file created from diffpair175.ext - technology: sky130A

.subckt diffpair175 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t15 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X1 drain_right.t11 minus.t0 source.t1 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X2 drain_right.t10 minus.t1 source.t7 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X3 source.t13 plus.t1 drain_left.t10 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X4 drain_left.t9 plus.t2 source.t18 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X5 source.t9 minus.t2 drain_right.t9 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X6 drain_left.t8 plus.t3 source.t23 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X7 source.t5 minus.t3 drain_right.t8 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X8 source.t6 minus.t4 drain_right.t7 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X9 source.t10 minus.t5 drain_right.t6 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X10 drain_left.t7 plus.t4 source.t22 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X11 source.t17 plus.t5 drain_left.t6 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X12 drain_right.t5 minus.t6 source.t4 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X13 source.t21 plus.t6 drain_left.t5 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X14 source.t16 plus.t7 drain_left.t4 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X15 a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X16 drain_right.t4 minus.t7 source.t8 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X17 drain_right.t3 minus.t8 source.t11 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X18 a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X19 drain_left.t3 plus.t8 source.t14 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X20 a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X21 source.t12 plus.t9 drain_left.t2 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X22 drain_left.t1 plus.t10 source.t20 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X23 a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X24 source.t0 minus.t9 drain_right.t2 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X25 drain_right.t1 minus.t10 source.t2 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X26 source.t19 plus.t11 drain_left.t0 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X27 source.t3 minus.t11 drain_right.t0 a_n1458_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n2 plus.t5 565.62
R1 plus.n11 plus.t4 565.62
R2 plus.n15 plus.t3 565.62
R3 plus.n24 plus.t1 565.62
R4 plus.n3 plus.t2 518.15
R5 plus.n1 plus.t11 518.15
R6 plus.n8 plus.t10 518.15
R7 plus.n10 plus.t9 518.15
R8 plus.n16 plus.t7 518.15
R9 plus.n14 plus.t0 518.15
R10 plus.n21 plus.t6 518.15
R11 plus.n23 plus.t8 518.15
R12 plus.n5 plus.n2 161.489
R13 plus.n18 plus.n15 161.489
R14 plus.n5 plus.n4 161.3
R15 plus.n7 plus.n6 161.3
R16 plus.n9 plus.n0 161.3
R17 plus.n12 plus.n11 161.3
R18 plus.n18 plus.n17 161.3
R19 plus.n20 plus.n19 161.3
R20 plus.n22 plus.n13 161.3
R21 plus.n25 plus.n24 161.3
R22 plus.n4 plus.n3 43.0884
R23 plus.n10 plus.n9 43.0884
R24 plus.n23 plus.n22 43.0884
R25 plus.n17 plus.n16 43.0884
R26 plus.n7 plus.n1 38.7066
R27 plus.n8 plus.n7 38.7066
R28 plus.n21 plus.n20 38.7066
R29 plus.n20 plus.n14 38.7066
R30 plus.n4 plus.n1 34.3247
R31 plus.n9 plus.n8 34.3247
R32 plus.n22 plus.n21 34.3247
R33 plus.n17 plus.n14 34.3247
R34 plus.n3 plus.n2 29.9429
R35 plus.n11 plus.n10 29.9429
R36 plus.n24 plus.n23 29.9429
R37 plus.n16 plus.n15 29.9429
R38 plus plus.n25 25.071
R39 plus plus.n12 8.68989
R40 plus.n6 plus.n5 0.189894
R41 plus.n6 plus.n0 0.189894
R42 plus.n12 plus.n0 0.189894
R43 plus.n25 plus.n13 0.189894
R44 plus.n19 plus.n13 0.189894
R45 plus.n19 plus.n18 0.189894
R46 source.n0 source.t22 69.6943
R47 source.n5 source.t17 69.6943
R48 source.n6 source.t8 69.6943
R49 source.n11 source.t5 69.6943
R50 source.n23 source.t2 69.6942
R51 source.n18 source.t9 69.6942
R52 source.n17 source.t23 69.6942
R53 source.n12 source.t13 69.6942
R54 source.n2 source.n1 63.0943
R55 source.n4 source.n3 63.0943
R56 source.n8 source.n7 63.0943
R57 source.n10 source.n9 63.0943
R58 source.n22 source.n21 63.0942
R59 source.n20 source.n19 63.0942
R60 source.n16 source.n15 63.0942
R61 source.n14 source.n13 63.0942
R62 source.n12 source.n11 14.9264
R63 source.n24 source.n0 9.43506
R64 source.n21 source.t7 6.6005
R65 source.n21 source.t10 6.6005
R66 source.n19 source.t4 6.6005
R67 source.n19 source.t3 6.6005
R68 source.n15 source.t15 6.6005
R69 source.n15 source.t16 6.6005
R70 source.n13 source.t14 6.6005
R71 source.n13 source.t21 6.6005
R72 source.n1 source.t20 6.6005
R73 source.n1 source.t12 6.6005
R74 source.n3 source.t18 6.6005
R75 source.n3 source.t19 6.6005
R76 source.n7 source.t1 6.6005
R77 source.n7 source.t6 6.6005
R78 source.n9 source.t11 6.6005
R79 source.n9 source.t0 6.6005
R80 source.n24 source.n23 5.49188
R81 source.n6 source.n5 0.470328
R82 source.n18 source.n17 0.470328
R83 source.n11 source.n10 0.457397
R84 source.n10 source.n8 0.457397
R85 source.n8 source.n6 0.457397
R86 source.n5 source.n4 0.457397
R87 source.n4 source.n2 0.457397
R88 source.n2 source.n0 0.457397
R89 source.n14 source.n12 0.457397
R90 source.n16 source.n14 0.457397
R91 source.n17 source.n16 0.457397
R92 source.n20 source.n18 0.457397
R93 source.n22 source.n20 0.457397
R94 source.n23 source.n22 0.457397
R95 source source.n24 0.188
R96 drain_left.n6 drain_left.n4 80.23
R97 drain_left.n3 drain_left.n2 80.1746
R98 drain_left.n3 drain_left.n0 80.1746
R99 drain_left.n8 drain_left.n7 79.7731
R100 drain_left.n6 drain_left.n5 79.7731
R101 drain_left.n3 drain_left.n1 79.773
R102 drain_left drain_left.n3 22.8334
R103 drain_left.n1 drain_left.t5 6.6005
R104 drain_left.n1 drain_left.t11 6.6005
R105 drain_left.n2 drain_left.t4 6.6005
R106 drain_left.n2 drain_left.t8 6.6005
R107 drain_left.n0 drain_left.t10 6.6005
R108 drain_left.n0 drain_left.t3 6.6005
R109 drain_left.n7 drain_left.t2 6.6005
R110 drain_left.n7 drain_left.t7 6.6005
R111 drain_left.n5 drain_left.t0 6.6005
R112 drain_left.n5 drain_left.t1 6.6005
R113 drain_left.n4 drain_left.t6 6.6005
R114 drain_left.n4 drain_left.t9 6.6005
R115 drain_left drain_left.n8 6.11011
R116 drain_left.n8 drain_left.n6 0.457397
R117 minus.n11 minus.t3 565.62
R118 minus.n2 minus.t7 565.62
R119 minus.n24 minus.t10 565.62
R120 minus.n15 minus.t2 565.62
R121 minus.n10 minus.t8 518.15
R122 minus.n8 minus.t9 518.15
R123 minus.n1 minus.t0 518.15
R124 minus.n3 minus.t4 518.15
R125 minus.n23 minus.t5 518.15
R126 minus.n21 minus.t1 518.15
R127 minus.n14 minus.t11 518.15
R128 minus.n16 minus.t6 518.15
R129 minus.n5 minus.n2 161.489
R130 minus.n18 minus.n15 161.489
R131 minus.n12 minus.n11 161.3
R132 minus.n9 minus.n0 161.3
R133 minus.n7 minus.n6 161.3
R134 minus.n5 minus.n4 161.3
R135 minus.n25 minus.n24 161.3
R136 minus.n22 minus.n13 161.3
R137 minus.n20 minus.n19 161.3
R138 minus.n18 minus.n17 161.3
R139 minus.n10 minus.n9 43.0884
R140 minus.n4 minus.n3 43.0884
R141 minus.n17 minus.n16 43.0884
R142 minus.n23 minus.n22 43.0884
R143 minus.n8 minus.n7 38.7066
R144 minus.n7 minus.n1 38.7066
R145 minus.n20 minus.n14 38.7066
R146 minus.n21 minus.n20 38.7066
R147 minus.n9 minus.n8 34.3247
R148 minus.n4 minus.n1 34.3247
R149 minus.n17 minus.n14 34.3247
R150 minus.n22 minus.n21 34.3247
R151 minus.n11 minus.n10 29.9429
R152 minus.n3 minus.n2 29.9429
R153 minus.n16 minus.n15 29.9429
R154 minus.n24 minus.n23 29.9429
R155 minus.n26 minus.n12 27.7808
R156 minus.n26 minus.n25 6.45505
R157 minus.n12 minus.n0 0.189894
R158 minus.n6 minus.n0 0.189894
R159 minus.n6 minus.n5 0.189894
R160 minus.n19 minus.n18 0.189894
R161 minus.n19 minus.n13 0.189894
R162 minus.n25 minus.n13 0.189894
R163 minus minus.n26 0.188
R164 drain_right.n6 drain_right.n4 80.23
R165 drain_right.n3 drain_right.n2 80.1746
R166 drain_right.n3 drain_right.n0 80.1746
R167 drain_right.n6 drain_right.n5 79.7731
R168 drain_right.n8 drain_right.n7 79.7731
R169 drain_right.n3 drain_right.n1 79.773
R170 drain_right drain_right.n3 22.2801
R171 drain_right.n1 drain_right.t0 6.6005
R172 drain_right.n1 drain_right.t10 6.6005
R173 drain_right.n2 drain_right.t6 6.6005
R174 drain_right.n2 drain_right.t1 6.6005
R175 drain_right.n0 drain_right.t9 6.6005
R176 drain_right.n0 drain_right.t5 6.6005
R177 drain_right.n4 drain_right.t7 6.6005
R178 drain_right.n4 drain_right.t4 6.6005
R179 drain_right.n5 drain_right.t2 6.6005
R180 drain_right.n5 drain_right.t11 6.6005
R181 drain_right.n7 drain_right.t8 6.6005
R182 drain_right.n7 drain_right.t3 6.6005
R183 drain_right drain_right.n8 6.11011
R184 drain_right.n8 drain_right.n6 0.457397
C0 plus drain_right 0.297597f
C1 drain_right minus 1.20122f
C2 drain_left drain_right 0.711854f
C3 plus source 1.22401f
C4 source minus 1.21001f
C5 source drain_left 8.71548f
C6 plus minus 3.3127f
C7 plus drain_left 1.34012f
C8 drain_left minus 0.175432f
C9 source drain_right 8.71461f
C10 drain_right a_n1458_n1488# 3.82233f
C11 drain_left a_n1458_n1488# 4.0319f
C12 source a_n1458_n1488# 3.492841f
C13 minus a_n1458_n1488# 4.920253f
C14 plus a_n1458_n1488# 5.623342f
C15 drain_right.t9 a_n1458_n1488# 0.072907f
C16 drain_right.t5 a_n1458_n1488# 0.072907f
C17 drain_right.n0 a_n1458_n1488# 0.527531f
C18 drain_right.t0 a_n1458_n1488# 0.072907f
C19 drain_right.t10 a_n1458_n1488# 0.072907f
C20 drain_right.n1 a_n1458_n1488# 0.525801f
C21 drain_right.t6 a_n1458_n1488# 0.072907f
C22 drain_right.t1 a_n1458_n1488# 0.072907f
C23 drain_right.n2 a_n1458_n1488# 0.527531f
C24 drain_right.n3 a_n1458_n1488# 1.72636f
C25 drain_right.t7 a_n1458_n1488# 0.072907f
C26 drain_right.t4 a_n1458_n1488# 0.072907f
C27 drain_right.n4 a_n1458_n1488# 0.527792f
C28 drain_right.t2 a_n1458_n1488# 0.072907f
C29 drain_right.t11 a_n1458_n1488# 0.072907f
C30 drain_right.n5 a_n1458_n1488# 0.525804f
C31 drain_right.n6 a_n1458_n1488# 0.683856f
C32 drain_right.t8 a_n1458_n1488# 0.072907f
C33 drain_right.t3 a_n1458_n1488# 0.072907f
C34 drain_right.n7 a_n1458_n1488# 0.525804f
C35 drain_right.n8 a_n1458_n1488# 0.588418f
C36 minus.n0 a_n1458_n1488# 0.031695f
C37 minus.t3 a_n1458_n1488# 0.058069f
C38 minus.t8 a_n1458_n1488# 0.055071f
C39 minus.t9 a_n1458_n1488# 0.055071f
C40 minus.t0 a_n1458_n1488# 0.055071f
C41 minus.n1 a_n1458_n1488# 0.035234f
C42 minus.t7 a_n1458_n1488# 0.058069f
C43 minus.n2 a_n1458_n1488# 0.04387f
C44 minus.t4 a_n1458_n1488# 0.055071f
C45 minus.n3 a_n1458_n1488# 0.035234f
C46 minus.n4 a_n1458_n1488# 0.011101f
C47 minus.n5 a_n1458_n1488# 0.070185f
C48 minus.n6 a_n1458_n1488# 0.031695f
C49 minus.n7 a_n1458_n1488# 0.011101f
C50 minus.n8 a_n1458_n1488# 0.035234f
C51 minus.n9 a_n1458_n1488# 0.011101f
C52 minus.n10 a_n1458_n1488# 0.035234f
C53 minus.n11 a_n1458_n1488# 0.043825f
C54 minus.n12 a_n1458_n1488# 0.71977f
C55 minus.n13 a_n1458_n1488# 0.031695f
C56 minus.t5 a_n1458_n1488# 0.055071f
C57 minus.t1 a_n1458_n1488# 0.055071f
C58 minus.t11 a_n1458_n1488# 0.055071f
C59 minus.n14 a_n1458_n1488# 0.035234f
C60 minus.t2 a_n1458_n1488# 0.058069f
C61 minus.n15 a_n1458_n1488# 0.04387f
C62 minus.t6 a_n1458_n1488# 0.055071f
C63 minus.n16 a_n1458_n1488# 0.035234f
C64 minus.n17 a_n1458_n1488# 0.011101f
C65 minus.n18 a_n1458_n1488# 0.070185f
C66 minus.n19 a_n1458_n1488# 0.031695f
C67 minus.n20 a_n1458_n1488# 0.011101f
C68 minus.n21 a_n1458_n1488# 0.035234f
C69 minus.n22 a_n1458_n1488# 0.011101f
C70 minus.n23 a_n1458_n1488# 0.035234f
C71 minus.t10 a_n1458_n1488# 0.058069f
C72 minus.n24 a_n1458_n1488# 0.043825f
C73 minus.n25 a_n1458_n1488# 0.203851f
C74 minus.n26 a_n1458_n1488# 0.891706f
C75 drain_left.t10 a_n1458_n1488# 0.071913f
C76 drain_left.t3 a_n1458_n1488# 0.071913f
C77 drain_left.n0 a_n1458_n1488# 0.520336f
C78 drain_left.t5 a_n1458_n1488# 0.071913f
C79 drain_left.t11 a_n1458_n1488# 0.071913f
C80 drain_left.n1 a_n1458_n1488# 0.51863f
C81 drain_left.t4 a_n1458_n1488# 0.071913f
C82 drain_left.t8 a_n1458_n1488# 0.071913f
C83 drain_left.n2 a_n1458_n1488# 0.520336f
C84 drain_left.n3 a_n1458_n1488# 1.7632f
C85 drain_left.t6 a_n1458_n1488# 0.071913f
C86 drain_left.t9 a_n1458_n1488# 0.071913f
C87 drain_left.n4 a_n1458_n1488# 0.520593f
C88 drain_left.t0 a_n1458_n1488# 0.071913f
C89 drain_left.t1 a_n1458_n1488# 0.071913f
C90 drain_left.n5 a_n1458_n1488# 0.518632f
C91 drain_left.n6 a_n1458_n1488# 0.674529f
C92 drain_left.t2 a_n1458_n1488# 0.071913f
C93 drain_left.t7 a_n1458_n1488# 0.071913f
C94 drain_left.n7 a_n1458_n1488# 0.518632f
C95 drain_left.n8 a_n1458_n1488# 0.580393f
C96 source.t22 a_n1458_n1488# 0.559466f
C97 source.n0 a_n1458_n1488# 0.749386f
C98 source.t20 a_n1458_n1488# 0.067374f
C99 source.t12 a_n1458_n1488# 0.067374f
C100 source.n1 a_n1458_n1488# 0.427193f
C101 source.n2 a_n1458_n1488# 0.331253f
C102 source.t18 a_n1458_n1488# 0.067374f
C103 source.t19 a_n1458_n1488# 0.067374f
C104 source.n3 a_n1458_n1488# 0.427193f
C105 source.n4 a_n1458_n1488# 0.331253f
C106 source.t17 a_n1458_n1488# 0.559466f
C107 source.n5 a_n1458_n1488# 0.383913f
C108 source.t8 a_n1458_n1488# 0.559466f
C109 source.n6 a_n1458_n1488# 0.383913f
C110 source.t1 a_n1458_n1488# 0.067374f
C111 source.t6 a_n1458_n1488# 0.067374f
C112 source.n7 a_n1458_n1488# 0.427193f
C113 source.n8 a_n1458_n1488# 0.331253f
C114 source.t11 a_n1458_n1488# 0.067374f
C115 source.t0 a_n1458_n1488# 0.067374f
C116 source.n9 a_n1458_n1488# 0.427193f
C117 source.n10 a_n1458_n1488# 0.331253f
C118 source.t5 a_n1458_n1488# 0.559466f
C119 source.n11 a_n1458_n1488# 1.04375f
C120 source.t13 a_n1458_n1488# 0.559463f
C121 source.n12 a_n1458_n1488# 1.04375f
C122 source.t14 a_n1458_n1488# 0.067374f
C123 source.t21 a_n1458_n1488# 0.067374f
C124 source.n13 a_n1458_n1488# 0.42719f
C125 source.n14 a_n1458_n1488# 0.331257f
C126 source.t15 a_n1458_n1488# 0.067374f
C127 source.t16 a_n1458_n1488# 0.067374f
C128 source.n15 a_n1458_n1488# 0.42719f
C129 source.n16 a_n1458_n1488# 0.331257f
C130 source.t23 a_n1458_n1488# 0.559463f
C131 source.n17 a_n1458_n1488# 0.383916f
C132 source.t9 a_n1458_n1488# 0.559463f
C133 source.n18 a_n1458_n1488# 0.383916f
C134 source.t4 a_n1458_n1488# 0.067374f
C135 source.t3 a_n1458_n1488# 0.067374f
C136 source.n19 a_n1458_n1488# 0.42719f
C137 source.n20 a_n1458_n1488# 0.331257f
C138 source.t7 a_n1458_n1488# 0.067374f
C139 source.t10 a_n1458_n1488# 0.067374f
C140 source.n21 a_n1458_n1488# 0.42719f
C141 source.n22 a_n1458_n1488# 0.331257f
C142 source.t2 a_n1458_n1488# 0.559463f
C143 source.n23 a_n1458_n1488# 0.538017f
C144 source.n24 a_n1458_n1488# 0.820311f
C145 plus.n0 a_n1458_n1488# 0.032323f
C146 plus.t9 a_n1458_n1488# 0.056162f
C147 plus.t10 a_n1458_n1488# 0.056162f
C148 plus.t11 a_n1458_n1488# 0.056162f
C149 plus.n1 a_n1458_n1488# 0.035932f
C150 plus.t5 a_n1458_n1488# 0.05922f
C151 plus.n2 a_n1458_n1488# 0.044739f
C152 plus.t2 a_n1458_n1488# 0.056162f
C153 plus.n3 a_n1458_n1488# 0.035932f
C154 plus.n4 a_n1458_n1488# 0.01132f
C155 plus.n5 a_n1458_n1488# 0.071575f
C156 plus.n6 a_n1458_n1488# 0.032323f
C157 plus.n7 a_n1458_n1488# 0.01132f
C158 plus.n8 a_n1458_n1488# 0.035932f
C159 plus.n9 a_n1458_n1488# 0.01132f
C160 plus.n10 a_n1458_n1488# 0.035932f
C161 plus.t4 a_n1458_n1488# 0.05922f
C162 plus.n11 a_n1458_n1488# 0.044693f
C163 plus.n12 a_n1458_n1488# 0.23784f
C164 plus.n13 a_n1458_n1488# 0.032323f
C165 plus.t1 a_n1458_n1488# 0.05922f
C166 plus.t8 a_n1458_n1488# 0.056162f
C167 plus.t6 a_n1458_n1488# 0.056162f
C168 plus.t0 a_n1458_n1488# 0.056162f
C169 plus.n14 a_n1458_n1488# 0.035932f
C170 plus.t3 a_n1458_n1488# 0.05922f
C171 plus.n15 a_n1458_n1488# 0.044739f
C172 plus.t7 a_n1458_n1488# 0.056162f
C173 plus.n16 a_n1458_n1488# 0.035932f
C174 plus.n17 a_n1458_n1488# 0.01132f
C175 plus.n18 a_n1458_n1488# 0.071575f
C176 plus.n19 a_n1458_n1488# 0.032323f
C177 plus.n20 a_n1458_n1488# 0.01132f
C178 plus.n21 a_n1458_n1488# 0.035932f
C179 plus.n22 a_n1458_n1488# 0.01132f
C180 plus.n23 a_n1458_n1488# 0.035932f
C181 plus.n24 a_n1458_n1488# 0.044693f
C182 plus.n25 a_n1458_n1488# 0.692522f
.ends

