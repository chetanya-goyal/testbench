* NGSPICE file created from diffpair265.ext - technology: sky130A

.subckt diffpair265 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t13 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_left.t10 plus.t1 source.t19 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t9 plus.t2 source.t16 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X4 source.t5 minus.t0 drain_right.t11 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X5 source.t8 minus.t1 drain_right.t10 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X6 a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X7 source.t11 plus.t3 drain_left.t8 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X8 drain_right.t9 minus.t2 source.t3 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X9 source.t7 minus.t3 drain_right.t8 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X10 source.t17 plus.t4 drain_left.t7 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X11 source.t9 minus.t4 drain_right.t7 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X12 source.t14 plus.t5 drain_left.t6 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X13 source.t18 plus.t6 drain_left.t5 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X14 source.t20 plus.t7 drain_left.t4 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X16 drain_left.t3 plus.t8 source.t15 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X17 drain_right.t6 minus.t5 source.t0 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X18 drain_right.t5 minus.t6 source.t1 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 source.t2 minus.t7 drain_right.t4 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X20 drain_right.t3 minus.t8 source.t6 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X21 a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X22 source.t12 plus.t9 drain_left.t2 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X23 drain_right.t2 minus.t9 source.t10 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X24 drain_left.t1 plus.t10 source.t22 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X25 drain_right.t1 minus.t10 source.t23 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X26 source.t4 minus.t11 drain_right.t0 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X27 drain_left.t0 plus.t11 source.t21 a_n1528_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
R0 plus.n2 plus.t3 732.933
R1 plus.n13 plus.t11 732.933
R2 plus.n17 plus.t8 732.933
R3 plus.n28 plus.t5 732.933
R4 plus.n3 plus.t1 703.721
R5 plus.n4 plus.t7 703.721
R6 plus.n10 plus.t0 703.721
R7 plus.n12 plus.t6 703.721
R8 plus.n19 plus.t4 703.721
R9 plus.n18 plus.t2 703.721
R10 plus.n25 plus.t9 703.721
R11 plus.n27 plus.t10 703.721
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 26.4536
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 9.80732
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n266 source.n240 289.615
R53 source.n230 source.n204 289.615
R54 source.n198 source.n172 289.615
R55 source.n162 source.n136 289.615
R56 source.n26 source.n0 289.615
R57 source.n62 source.n36 289.615
R58 source.n94 source.n68 289.615
R59 source.n130 source.n104 289.615
R60 source.n251 source.n250 185
R61 source.n248 source.n247 185
R62 source.n257 source.n256 185
R63 source.n259 source.n258 185
R64 source.n244 source.n243 185
R65 source.n265 source.n264 185
R66 source.n267 source.n266 185
R67 source.n215 source.n214 185
R68 source.n212 source.n211 185
R69 source.n221 source.n220 185
R70 source.n223 source.n222 185
R71 source.n208 source.n207 185
R72 source.n229 source.n228 185
R73 source.n231 source.n230 185
R74 source.n183 source.n182 185
R75 source.n180 source.n179 185
R76 source.n189 source.n188 185
R77 source.n191 source.n190 185
R78 source.n176 source.n175 185
R79 source.n197 source.n196 185
R80 source.n199 source.n198 185
R81 source.n147 source.n146 185
R82 source.n144 source.n143 185
R83 source.n153 source.n152 185
R84 source.n155 source.n154 185
R85 source.n140 source.n139 185
R86 source.n161 source.n160 185
R87 source.n163 source.n162 185
R88 source.n27 source.n26 185
R89 source.n25 source.n24 185
R90 source.n4 source.n3 185
R91 source.n19 source.n18 185
R92 source.n17 source.n16 185
R93 source.n8 source.n7 185
R94 source.n11 source.n10 185
R95 source.n63 source.n62 185
R96 source.n61 source.n60 185
R97 source.n40 source.n39 185
R98 source.n55 source.n54 185
R99 source.n53 source.n52 185
R100 source.n44 source.n43 185
R101 source.n47 source.n46 185
R102 source.n95 source.n94 185
R103 source.n93 source.n92 185
R104 source.n72 source.n71 185
R105 source.n87 source.n86 185
R106 source.n85 source.n84 185
R107 source.n76 source.n75 185
R108 source.n79 source.n78 185
R109 source.n131 source.n130 185
R110 source.n129 source.n128 185
R111 source.n108 source.n107 185
R112 source.n123 source.n122 185
R113 source.n121 source.n120 185
R114 source.n112 source.n111 185
R115 source.n115 source.n114 185
R116 source.t0 source.n249 147.661
R117 source.t2 source.n213 147.661
R118 source.t15 source.n181 147.661
R119 source.t14 source.n145 147.661
R120 source.t21 source.n9 147.661
R121 source.t11 source.n45 147.661
R122 source.t6 source.n77 147.661
R123 source.t7 source.n113 147.661
R124 source.n250 source.n247 104.615
R125 source.n257 source.n247 104.615
R126 source.n258 source.n257 104.615
R127 source.n258 source.n243 104.615
R128 source.n265 source.n243 104.615
R129 source.n266 source.n265 104.615
R130 source.n214 source.n211 104.615
R131 source.n221 source.n211 104.615
R132 source.n222 source.n221 104.615
R133 source.n222 source.n207 104.615
R134 source.n229 source.n207 104.615
R135 source.n230 source.n229 104.615
R136 source.n182 source.n179 104.615
R137 source.n189 source.n179 104.615
R138 source.n190 source.n189 104.615
R139 source.n190 source.n175 104.615
R140 source.n197 source.n175 104.615
R141 source.n198 source.n197 104.615
R142 source.n146 source.n143 104.615
R143 source.n153 source.n143 104.615
R144 source.n154 source.n153 104.615
R145 source.n154 source.n139 104.615
R146 source.n161 source.n139 104.615
R147 source.n162 source.n161 104.615
R148 source.n26 source.n25 104.615
R149 source.n25 source.n3 104.615
R150 source.n18 source.n3 104.615
R151 source.n18 source.n17 104.615
R152 source.n17 source.n7 104.615
R153 source.n10 source.n7 104.615
R154 source.n62 source.n61 104.615
R155 source.n61 source.n39 104.615
R156 source.n54 source.n39 104.615
R157 source.n54 source.n53 104.615
R158 source.n53 source.n43 104.615
R159 source.n46 source.n43 104.615
R160 source.n94 source.n93 104.615
R161 source.n93 source.n71 104.615
R162 source.n86 source.n71 104.615
R163 source.n86 source.n85 104.615
R164 source.n85 source.n75 104.615
R165 source.n78 source.n75 104.615
R166 source.n130 source.n129 104.615
R167 source.n129 source.n107 104.615
R168 source.n122 source.n107 104.615
R169 source.n122 source.n121 104.615
R170 source.n121 source.n111 104.615
R171 source.n114 source.n111 104.615
R172 source.n250 source.t0 52.3082
R173 source.n214 source.t2 52.3082
R174 source.n182 source.t15 52.3082
R175 source.n146 source.t14 52.3082
R176 source.n10 source.t21 52.3082
R177 source.n46 source.t11 52.3082
R178 source.n78 source.t6 52.3082
R179 source.n114 source.t7 52.3082
R180 source.n33 source.n32 50.512
R181 source.n35 source.n34 50.512
R182 source.n101 source.n100 50.512
R183 source.n103 source.n102 50.512
R184 source.n239 source.n238 50.5119
R185 source.n237 source.n236 50.5119
R186 source.n171 source.n170 50.5119
R187 source.n169 source.n168 50.5119
R188 source.n271 source.n270 32.1853
R189 source.n235 source.n234 32.1853
R190 source.n203 source.n202 32.1853
R191 source.n167 source.n166 32.1853
R192 source.n31 source.n30 32.1853
R193 source.n67 source.n66 32.1853
R194 source.n99 source.n98 32.1853
R195 source.n135 source.n134 32.1853
R196 source.n167 source.n135 17.2423
R197 source.n251 source.n249 15.6674
R198 source.n215 source.n213 15.6674
R199 source.n183 source.n181 15.6674
R200 source.n147 source.n145 15.6674
R201 source.n11 source.n9 15.6674
R202 source.n47 source.n45 15.6674
R203 source.n79 source.n77 15.6674
R204 source.n115 source.n113 15.6674
R205 source.n252 source.n248 12.8005
R206 source.n216 source.n212 12.8005
R207 source.n184 source.n180 12.8005
R208 source.n148 source.n144 12.8005
R209 source.n12 source.n8 12.8005
R210 source.n48 source.n44 12.8005
R211 source.n80 source.n76 12.8005
R212 source.n116 source.n112 12.8005
R213 source.n256 source.n255 12.0247
R214 source.n220 source.n219 12.0247
R215 source.n188 source.n187 12.0247
R216 source.n152 source.n151 12.0247
R217 source.n16 source.n15 12.0247
R218 source.n52 source.n51 12.0247
R219 source.n84 source.n83 12.0247
R220 source.n120 source.n119 12.0247
R221 source.n272 source.n31 11.7293
R222 source.n259 source.n246 11.249
R223 source.n223 source.n210 11.249
R224 source.n191 source.n178 11.249
R225 source.n155 source.n142 11.249
R226 source.n19 source.n6 11.249
R227 source.n55 source.n42 11.249
R228 source.n87 source.n74 11.249
R229 source.n123 source.n110 11.249
R230 source.n260 source.n244 10.4732
R231 source.n224 source.n208 10.4732
R232 source.n192 source.n176 10.4732
R233 source.n156 source.n140 10.4732
R234 source.n20 source.n4 10.4732
R235 source.n56 source.n40 10.4732
R236 source.n88 source.n72 10.4732
R237 source.n124 source.n108 10.4732
R238 source.n264 source.n263 9.69747
R239 source.n228 source.n227 9.69747
R240 source.n196 source.n195 9.69747
R241 source.n160 source.n159 9.69747
R242 source.n24 source.n23 9.69747
R243 source.n60 source.n59 9.69747
R244 source.n92 source.n91 9.69747
R245 source.n128 source.n127 9.69747
R246 source.n270 source.n269 9.45567
R247 source.n234 source.n233 9.45567
R248 source.n202 source.n201 9.45567
R249 source.n166 source.n165 9.45567
R250 source.n30 source.n29 9.45567
R251 source.n66 source.n65 9.45567
R252 source.n98 source.n97 9.45567
R253 source.n134 source.n133 9.45567
R254 source.n269 source.n268 9.3005
R255 source.n242 source.n241 9.3005
R256 source.n263 source.n262 9.3005
R257 source.n261 source.n260 9.3005
R258 source.n246 source.n245 9.3005
R259 source.n255 source.n254 9.3005
R260 source.n253 source.n252 9.3005
R261 source.n233 source.n232 9.3005
R262 source.n206 source.n205 9.3005
R263 source.n227 source.n226 9.3005
R264 source.n225 source.n224 9.3005
R265 source.n210 source.n209 9.3005
R266 source.n219 source.n218 9.3005
R267 source.n217 source.n216 9.3005
R268 source.n201 source.n200 9.3005
R269 source.n174 source.n173 9.3005
R270 source.n195 source.n194 9.3005
R271 source.n193 source.n192 9.3005
R272 source.n178 source.n177 9.3005
R273 source.n187 source.n186 9.3005
R274 source.n185 source.n184 9.3005
R275 source.n165 source.n164 9.3005
R276 source.n138 source.n137 9.3005
R277 source.n159 source.n158 9.3005
R278 source.n157 source.n156 9.3005
R279 source.n142 source.n141 9.3005
R280 source.n151 source.n150 9.3005
R281 source.n149 source.n148 9.3005
R282 source.n29 source.n28 9.3005
R283 source.n2 source.n1 9.3005
R284 source.n23 source.n22 9.3005
R285 source.n21 source.n20 9.3005
R286 source.n6 source.n5 9.3005
R287 source.n15 source.n14 9.3005
R288 source.n13 source.n12 9.3005
R289 source.n65 source.n64 9.3005
R290 source.n38 source.n37 9.3005
R291 source.n59 source.n58 9.3005
R292 source.n57 source.n56 9.3005
R293 source.n42 source.n41 9.3005
R294 source.n51 source.n50 9.3005
R295 source.n49 source.n48 9.3005
R296 source.n97 source.n96 9.3005
R297 source.n70 source.n69 9.3005
R298 source.n91 source.n90 9.3005
R299 source.n89 source.n88 9.3005
R300 source.n74 source.n73 9.3005
R301 source.n83 source.n82 9.3005
R302 source.n81 source.n80 9.3005
R303 source.n133 source.n132 9.3005
R304 source.n106 source.n105 9.3005
R305 source.n127 source.n126 9.3005
R306 source.n125 source.n124 9.3005
R307 source.n110 source.n109 9.3005
R308 source.n119 source.n118 9.3005
R309 source.n117 source.n116 9.3005
R310 source.n267 source.n242 8.92171
R311 source.n231 source.n206 8.92171
R312 source.n199 source.n174 8.92171
R313 source.n163 source.n138 8.92171
R314 source.n27 source.n2 8.92171
R315 source.n63 source.n38 8.92171
R316 source.n95 source.n70 8.92171
R317 source.n131 source.n106 8.92171
R318 source.n268 source.n240 8.14595
R319 source.n232 source.n204 8.14595
R320 source.n200 source.n172 8.14595
R321 source.n164 source.n136 8.14595
R322 source.n28 source.n0 8.14595
R323 source.n64 source.n36 8.14595
R324 source.n96 source.n68 8.14595
R325 source.n132 source.n104 8.14595
R326 source.n270 source.n240 5.81868
R327 source.n234 source.n204 5.81868
R328 source.n202 source.n172 5.81868
R329 source.n166 source.n136 5.81868
R330 source.n30 source.n0 5.81868
R331 source.n66 source.n36 5.81868
R332 source.n98 source.n68 5.81868
R333 source.n134 source.n104 5.81868
R334 source.n272 source.n271 5.51343
R335 source.n268 source.n267 5.04292
R336 source.n232 source.n231 5.04292
R337 source.n200 source.n199 5.04292
R338 source.n164 source.n163 5.04292
R339 source.n28 source.n27 5.04292
R340 source.n64 source.n63 5.04292
R341 source.n96 source.n95 5.04292
R342 source.n132 source.n131 5.04292
R343 source.n253 source.n249 4.38594
R344 source.n217 source.n213 4.38594
R345 source.n185 source.n181 4.38594
R346 source.n149 source.n145 4.38594
R347 source.n13 source.n9 4.38594
R348 source.n49 source.n45 4.38594
R349 source.n81 source.n77 4.38594
R350 source.n117 source.n113 4.38594
R351 source.n264 source.n242 4.26717
R352 source.n228 source.n206 4.26717
R353 source.n196 source.n174 4.26717
R354 source.n160 source.n138 4.26717
R355 source.n24 source.n2 4.26717
R356 source.n60 source.n38 4.26717
R357 source.n92 source.n70 4.26717
R358 source.n128 source.n106 4.26717
R359 source.n263 source.n244 3.49141
R360 source.n227 source.n208 3.49141
R361 source.n195 source.n176 3.49141
R362 source.n159 source.n140 3.49141
R363 source.n23 source.n4 3.49141
R364 source.n59 source.n40 3.49141
R365 source.n91 source.n72 3.49141
R366 source.n127 source.n108 3.49141
R367 source.n238 source.t3 3.3005
R368 source.n238 source.t4 3.3005
R369 source.n236 source.t10 3.3005
R370 source.n236 source.t9 3.3005
R371 source.n170 source.t16 3.3005
R372 source.n170 source.t17 3.3005
R373 source.n168 source.t22 3.3005
R374 source.n168 source.t12 3.3005
R375 source.n32 source.t13 3.3005
R376 source.n32 source.t18 3.3005
R377 source.n34 source.t19 3.3005
R378 source.n34 source.t20 3.3005
R379 source.n100 source.t1 3.3005
R380 source.n100 source.t8 3.3005
R381 source.n102 source.t23 3.3005
R382 source.n102 source.t5 3.3005
R383 source.n260 source.n259 2.71565
R384 source.n224 source.n223 2.71565
R385 source.n192 source.n191 2.71565
R386 source.n156 source.n155 2.71565
R387 source.n20 source.n19 2.71565
R388 source.n56 source.n55 2.71565
R389 source.n88 source.n87 2.71565
R390 source.n124 source.n123 2.71565
R391 source.n256 source.n246 1.93989
R392 source.n220 source.n210 1.93989
R393 source.n188 source.n178 1.93989
R394 source.n152 source.n142 1.93989
R395 source.n16 source.n6 1.93989
R396 source.n52 source.n42 1.93989
R397 source.n84 source.n74 1.93989
R398 source.n120 source.n110 1.93989
R399 source.n255 source.n248 1.16414
R400 source.n219 source.n212 1.16414
R401 source.n187 source.n180 1.16414
R402 source.n151 source.n144 1.16414
R403 source.n15 source.n8 1.16414
R404 source.n51 source.n44 1.16414
R405 source.n83 source.n76 1.16414
R406 source.n119 source.n112 1.16414
R407 source.n135 source.n103 0.5005
R408 source.n103 source.n101 0.5005
R409 source.n101 source.n99 0.5005
R410 source.n67 source.n35 0.5005
R411 source.n35 source.n33 0.5005
R412 source.n33 source.n31 0.5005
R413 source.n169 source.n167 0.5005
R414 source.n171 source.n169 0.5005
R415 source.n203 source.n171 0.5005
R416 source.n237 source.n235 0.5005
R417 source.n239 source.n237 0.5005
R418 source.n271 source.n239 0.5005
R419 source.n99 source.n67 0.470328
R420 source.n235 source.n203 0.470328
R421 source.n252 source.n251 0.388379
R422 source.n216 source.n215 0.388379
R423 source.n184 source.n183 0.388379
R424 source.n148 source.n147 0.388379
R425 source.n12 source.n11 0.388379
R426 source.n48 source.n47 0.388379
R427 source.n80 source.n79 0.388379
R428 source.n116 source.n115 0.388379
R429 source source.n272 0.188
R430 source.n254 source.n253 0.155672
R431 source.n254 source.n245 0.155672
R432 source.n261 source.n245 0.155672
R433 source.n262 source.n261 0.155672
R434 source.n262 source.n241 0.155672
R435 source.n269 source.n241 0.155672
R436 source.n218 source.n217 0.155672
R437 source.n218 source.n209 0.155672
R438 source.n225 source.n209 0.155672
R439 source.n226 source.n225 0.155672
R440 source.n226 source.n205 0.155672
R441 source.n233 source.n205 0.155672
R442 source.n186 source.n185 0.155672
R443 source.n186 source.n177 0.155672
R444 source.n193 source.n177 0.155672
R445 source.n194 source.n193 0.155672
R446 source.n194 source.n173 0.155672
R447 source.n201 source.n173 0.155672
R448 source.n150 source.n149 0.155672
R449 source.n150 source.n141 0.155672
R450 source.n157 source.n141 0.155672
R451 source.n158 source.n157 0.155672
R452 source.n158 source.n137 0.155672
R453 source.n165 source.n137 0.155672
R454 source.n29 source.n1 0.155672
R455 source.n22 source.n1 0.155672
R456 source.n22 source.n21 0.155672
R457 source.n21 source.n5 0.155672
R458 source.n14 source.n5 0.155672
R459 source.n14 source.n13 0.155672
R460 source.n65 source.n37 0.155672
R461 source.n58 source.n37 0.155672
R462 source.n58 source.n57 0.155672
R463 source.n57 source.n41 0.155672
R464 source.n50 source.n41 0.155672
R465 source.n50 source.n49 0.155672
R466 source.n97 source.n69 0.155672
R467 source.n90 source.n69 0.155672
R468 source.n90 source.n89 0.155672
R469 source.n89 source.n73 0.155672
R470 source.n82 source.n73 0.155672
R471 source.n82 source.n81 0.155672
R472 source.n133 source.n105 0.155672
R473 source.n126 source.n105 0.155672
R474 source.n126 source.n125 0.155672
R475 source.n125 source.n109 0.155672
R476 source.n118 source.n109 0.155672
R477 source.n118 source.n117 0.155672
R478 drain_left.n6 drain_left.n4 67.6908
R479 drain_left.n3 drain_left.n2 67.6353
R480 drain_left.n3 drain_left.n0 67.6353
R481 drain_left.n6 drain_left.n5 67.1908
R482 drain_left.n8 drain_left.n7 67.1907
R483 drain_left.n3 drain_left.n1 67.1907
R484 drain_left drain_left.n3 25.3216
R485 drain_left drain_left.n8 6.15322
R486 drain_left.n1 drain_left.t2 3.3005
R487 drain_left.n1 drain_left.t9 3.3005
R488 drain_left.n2 drain_left.t7 3.3005
R489 drain_left.n2 drain_left.t3 3.3005
R490 drain_left.n0 drain_left.t6 3.3005
R491 drain_left.n0 drain_left.t1 3.3005
R492 drain_left.n7 drain_left.t5 3.3005
R493 drain_left.n7 drain_left.t0 3.3005
R494 drain_left.n5 drain_left.t4 3.3005
R495 drain_left.n5 drain_left.t11 3.3005
R496 drain_left.n4 drain_left.t8 3.3005
R497 drain_left.n4 drain_left.t10 3.3005
R498 drain_left.n8 drain_left.n6 0.5005
R499 minus.n13 minus.t3 732.933
R500 minus.n2 minus.t8 732.933
R501 minus.n28 minus.t5 732.933
R502 minus.n17 minus.t7 732.933
R503 minus.n12 minus.t10 703.721
R504 minus.n10 minus.t0 703.721
R505 minus.n3 minus.t6 703.721
R506 minus.n4 minus.t1 703.721
R507 minus.n27 minus.t11 703.721
R508 minus.n25 minus.t2 703.721
R509 minus.n19 minus.t4 703.721
R510 minus.n18 minus.t9 703.721
R511 minus.n6 minus.n2 161.489
R512 minus.n21 minus.n17 161.489
R513 minus.n14 minus.n13 161.3
R514 minus.n11 minus.n0 161.3
R515 minus.n9 minus.n8 161.3
R516 minus.n7 minus.n1 161.3
R517 minus.n6 minus.n5 161.3
R518 minus.n29 minus.n28 161.3
R519 minus.n26 minus.n15 161.3
R520 minus.n24 minus.n23 161.3
R521 minus.n22 minus.n16 161.3
R522 minus.n21 minus.n20 161.3
R523 minus.n9 minus.n1 73.0308
R524 minus.n24 minus.n16 73.0308
R525 minus.n11 minus.n10 67.1884
R526 minus.n5 minus.n3 67.1884
R527 minus.n20 minus.n19 67.1884
R528 minus.n26 minus.n25 67.1884
R529 minus.n13 minus.n12 55.5035
R530 minus.n4 minus.n2 55.5035
R531 minus.n18 minus.n17 55.5035
R532 minus.n28 minus.n27 55.5035
R533 minus.n30 minus.n14 30.2997
R534 minus.n12 minus.n11 17.5278
R535 minus.n5 minus.n4 17.5278
R536 minus.n20 minus.n18 17.5278
R537 minus.n27 minus.n26 17.5278
R538 minus.n30 minus.n29 6.43611
R539 minus.n10 minus.n9 5.84292
R540 minus.n3 minus.n1 5.84292
R541 minus.n19 minus.n16 5.84292
R542 minus.n25 minus.n24 5.84292
R543 minus.n14 minus.n0 0.189894
R544 minus.n8 minus.n0 0.189894
R545 minus.n8 minus.n7 0.189894
R546 minus.n7 minus.n6 0.189894
R547 minus.n22 minus.n21 0.189894
R548 minus.n23 minus.n22 0.189894
R549 minus.n23 minus.n15 0.189894
R550 minus.n29 minus.n15 0.189894
R551 minus minus.n30 0.188
R552 drain_right.n6 drain_right.n4 67.6907
R553 drain_right.n3 drain_right.n2 67.6353
R554 drain_right.n3 drain_right.n0 67.6353
R555 drain_right.n6 drain_right.n5 67.1908
R556 drain_right.n8 drain_right.n7 67.1908
R557 drain_right.n3 drain_right.n1 67.1907
R558 drain_right drain_right.n3 24.7684
R559 drain_right drain_right.n8 6.15322
R560 drain_right.n1 drain_right.t7 3.3005
R561 drain_right.n1 drain_right.t9 3.3005
R562 drain_right.n2 drain_right.t0 3.3005
R563 drain_right.n2 drain_right.t6 3.3005
R564 drain_right.n0 drain_right.t4 3.3005
R565 drain_right.n0 drain_right.t2 3.3005
R566 drain_right.n4 drain_right.t10 3.3005
R567 drain_right.n4 drain_right.t3 3.3005
R568 drain_right.n5 drain_right.t11 3.3005
R569 drain_right.n5 drain_right.t5 3.3005
R570 drain_right.n7 drain_right.t8 3.3005
R571 drain_right.n7 drain_right.t1 3.3005
R572 drain_right.n8 drain_right.n6 0.5005
C0 plus source 2.16251f
C1 plus drain_right 0.300071f
C2 plus drain_left 2.40371f
C3 plus minus 3.95112f
C4 drain_right source 13.9247f
C5 drain_left source 13.9253f
C6 drain_right drain_left 0.751086f
C7 minus source 2.14849f
C8 minus drain_right 2.25754f
C9 minus drain_left 0.171004f
C10 drain_right a_n1528_n2088# 4.82884f
C11 drain_left a_n1528_n2088# 5.06928f
C12 source a_n1528_n2088# 5.204087f
C13 minus a_n1528_n2088# 5.459149f
C14 plus a_n1528_n2088# 7.05838f
C15 drain_right.t4 a_n1528_n2088# 0.163829f
C16 drain_right.t2 a_n1528_n2088# 0.163829f
C17 drain_right.n0 a_n1528_n2088# 1.36897f
C18 drain_right.t7 a_n1528_n2088# 0.163829f
C19 drain_right.t9 a_n1528_n2088# 0.163829f
C20 drain_right.n1 a_n1528_n2088# 1.36633f
C21 drain_right.t0 a_n1528_n2088# 0.163829f
C22 drain_right.t6 a_n1528_n2088# 0.163829f
C23 drain_right.n2 a_n1528_n2088# 1.36897f
C24 drain_right.n3 a_n1528_n2088# 2.19311f
C25 drain_right.t10 a_n1528_n2088# 0.163829f
C26 drain_right.t3 a_n1528_n2088# 0.163829f
C27 drain_right.n4 a_n1528_n2088# 1.36933f
C28 drain_right.t11 a_n1528_n2088# 0.163829f
C29 drain_right.t5 a_n1528_n2088# 0.163829f
C30 drain_right.n5 a_n1528_n2088# 1.36634f
C31 drain_right.n6 a_n1528_n2088# 0.794476f
C32 drain_right.t8 a_n1528_n2088# 0.163829f
C33 drain_right.t1 a_n1528_n2088# 0.163829f
C34 drain_right.n7 a_n1528_n2088# 1.36634f
C35 drain_right.n8 a_n1528_n2088# 0.676985f
C36 minus.n0 a_n1528_n2088# 0.05383f
C37 minus.t3 a_n1528_n2088# 0.234308f
C38 minus.t10 a_n1528_n2088# 0.230055f
C39 minus.t0 a_n1528_n2088# 0.230055f
C40 minus.n1 a_n1528_n2088# 0.019185f
C41 minus.t8 a_n1528_n2088# 0.234308f
C42 minus.n2 a_n1528_n2088# 0.123034f
C43 minus.t6 a_n1528_n2088# 0.230055f
C44 minus.n3 a_n1528_n2088# 0.108365f
C45 minus.t1 a_n1528_n2088# 0.230055f
C46 minus.n4 a_n1528_n2088# 0.108365f
C47 minus.n5 a_n1528_n2088# 0.020512f
C48 minus.n6 a_n1528_n2088# 0.112569f
C49 minus.n7 a_n1528_n2088# 0.05383f
C50 minus.n8 a_n1528_n2088# 0.05383f
C51 minus.n9 a_n1528_n2088# 0.019185f
C52 minus.n10 a_n1528_n2088# 0.108365f
C53 minus.n11 a_n1528_n2088# 0.020512f
C54 minus.n12 a_n1528_n2088# 0.108365f
C55 minus.n13 a_n1528_n2088# 0.122965f
C56 minus.n14 a_n1528_n2088# 1.42108f
C57 minus.n15 a_n1528_n2088# 0.05383f
C58 minus.t11 a_n1528_n2088# 0.230055f
C59 minus.t2 a_n1528_n2088# 0.230055f
C60 minus.n16 a_n1528_n2088# 0.019185f
C61 minus.t7 a_n1528_n2088# 0.234308f
C62 minus.n17 a_n1528_n2088# 0.123034f
C63 minus.t9 a_n1528_n2088# 0.230055f
C64 minus.n18 a_n1528_n2088# 0.108365f
C65 minus.t4 a_n1528_n2088# 0.230055f
C66 minus.n19 a_n1528_n2088# 0.108365f
C67 minus.n20 a_n1528_n2088# 0.020512f
C68 minus.n21 a_n1528_n2088# 0.112569f
C69 minus.n22 a_n1528_n2088# 0.05383f
C70 minus.n23 a_n1528_n2088# 0.05383f
C71 minus.n24 a_n1528_n2088# 0.019185f
C72 minus.n25 a_n1528_n2088# 0.108365f
C73 minus.n26 a_n1528_n2088# 0.020512f
C74 minus.n27 a_n1528_n2088# 0.108365f
C75 minus.t5 a_n1528_n2088# 0.234308f
C76 minus.n28 a_n1528_n2088# 0.122965f
C77 minus.n29 a_n1528_n2088# 0.343797f
C78 minus.n30 a_n1528_n2088# 1.75628f
C79 drain_left.t6 a_n1528_n2088# 0.163476f
C80 drain_left.t1 a_n1528_n2088# 0.163476f
C81 drain_left.n0 a_n1528_n2088# 1.36602f
C82 drain_left.t2 a_n1528_n2088# 0.163476f
C83 drain_left.t9 a_n1528_n2088# 0.163476f
C84 drain_left.n1 a_n1528_n2088# 1.36339f
C85 drain_left.t7 a_n1528_n2088# 0.163476f
C86 drain_left.t3 a_n1528_n2088# 0.163476f
C87 drain_left.n2 a_n1528_n2088# 1.36602f
C88 drain_left.n3 a_n1528_n2088# 2.25874f
C89 drain_left.t8 a_n1528_n2088# 0.163476f
C90 drain_left.t10 a_n1528_n2088# 0.163476f
C91 drain_left.n4 a_n1528_n2088# 1.36639f
C92 drain_left.t4 a_n1528_n2088# 0.163476f
C93 drain_left.t11 a_n1528_n2088# 0.163476f
C94 drain_left.n5 a_n1528_n2088# 1.3634f
C95 drain_left.n6 a_n1528_n2088# 0.792759f
C96 drain_left.t5 a_n1528_n2088# 0.163476f
C97 drain_left.t0 a_n1528_n2088# 0.163476f
C98 drain_left.n7 a_n1528_n2088# 1.36339f
C99 drain_left.n8 a_n1528_n2088# 0.675534f
C100 source.n0 a_n1528_n2088# 0.040845f
C101 source.n1 a_n1528_n2088# 0.029059f
C102 source.n2 a_n1528_n2088# 0.015615f
C103 source.n3 a_n1528_n2088# 0.036908f
C104 source.n4 a_n1528_n2088# 0.016534f
C105 source.n5 a_n1528_n2088# 0.029059f
C106 source.n6 a_n1528_n2088# 0.015615f
C107 source.n7 a_n1528_n2088# 0.036908f
C108 source.n8 a_n1528_n2088# 0.016534f
C109 source.n9 a_n1528_n2088# 0.124353f
C110 source.t21 a_n1528_n2088# 0.060156f
C111 source.n10 a_n1528_n2088# 0.027681f
C112 source.n11 a_n1528_n2088# 0.021801f
C113 source.n12 a_n1528_n2088# 0.015615f
C114 source.n13 a_n1528_n2088# 0.691434f
C115 source.n14 a_n1528_n2088# 0.029059f
C116 source.n15 a_n1528_n2088# 0.015615f
C117 source.n16 a_n1528_n2088# 0.016534f
C118 source.n17 a_n1528_n2088# 0.036908f
C119 source.n18 a_n1528_n2088# 0.036908f
C120 source.n19 a_n1528_n2088# 0.016534f
C121 source.n20 a_n1528_n2088# 0.015615f
C122 source.n21 a_n1528_n2088# 0.029059f
C123 source.n22 a_n1528_n2088# 0.029059f
C124 source.n23 a_n1528_n2088# 0.015615f
C125 source.n24 a_n1528_n2088# 0.016534f
C126 source.n25 a_n1528_n2088# 0.036908f
C127 source.n26 a_n1528_n2088# 0.079901f
C128 source.n27 a_n1528_n2088# 0.016534f
C129 source.n28 a_n1528_n2088# 0.015615f
C130 source.n29 a_n1528_n2088# 0.067169f
C131 source.n30 a_n1528_n2088# 0.044707f
C132 source.n31 a_n1528_n2088# 0.696949f
C133 source.t13 a_n1528_n2088# 0.13778f
C134 source.t18 a_n1528_n2088# 0.13778f
C135 source.n32 a_n1528_n2088# 1.07305f
C136 source.n33 a_n1528_n2088# 0.366037f
C137 source.t19 a_n1528_n2088# 0.13778f
C138 source.t20 a_n1528_n2088# 0.13778f
C139 source.n34 a_n1528_n2088# 1.07305f
C140 source.n35 a_n1528_n2088# 0.366037f
C141 source.n36 a_n1528_n2088# 0.040845f
C142 source.n37 a_n1528_n2088# 0.029059f
C143 source.n38 a_n1528_n2088# 0.015615f
C144 source.n39 a_n1528_n2088# 0.036908f
C145 source.n40 a_n1528_n2088# 0.016534f
C146 source.n41 a_n1528_n2088# 0.029059f
C147 source.n42 a_n1528_n2088# 0.015615f
C148 source.n43 a_n1528_n2088# 0.036908f
C149 source.n44 a_n1528_n2088# 0.016534f
C150 source.n45 a_n1528_n2088# 0.124353f
C151 source.t11 a_n1528_n2088# 0.060156f
C152 source.n46 a_n1528_n2088# 0.027681f
C153 source.n47 a_n1528_n2088# 0.021801f
C154 source.n48 a_n1528_n2088# 0.015615f
C155 source.n49 a_n1528_n2088# 0.691434f
C156 source.n50 a_n1528_n2088# 0.029059f
C157 source.n51 a_n1528_n2088# 0.015615f
C158 source.n52 a_n1528_n2088# 0.016534f
C159 source.n53 a_n1528_n2088# 0.036908f
C160 source.n54 a_n1528_n2088# 0.036908f
C161 source.n55 a_n1528_n2088# 0.016534f
C162 source.n56 a_n1528_n2088# 0.015615f
C163 source.n57 a_n1528_n2088# 0.029059f
C164 source.n58 a_n1528_n2088# 0.029059f
C165 source.n59 a_n1528_n2088# 0.015615f
C166 source.n60 a_n1528_n2088# 0.016534f
C167 source.n61 a_n1528_n2088# 0.036908f
C168 source.n62 a_n1528_n2088# 0.079901f
C169 source.n63 a_n1528_n2088# 0.016534f
C170 source.n64 a_n1528_n2088# 0.015615f
C171 source.n65 a_n1528_n2088# 0.067169f
C172 source.n66 a_n1528_n2088# 0.044707f
C173 source.n67 a_n1528_n2088# 0.115628f
C174 source.n68 a_n1528_n2088# 0.040845f
C175 source.n69 a_n1528_n2088# 0.029059f
C176 source.n70 a_n1528_n2088# 0.015615f
C177 source.n71 a_n1528_n2088# 0.036908f
C178 source.n72 a_n1528_n2088# 0.016534f
C179 source.n73 a_n1528_n2088# 0.029059f
C180 source.n74 a_n1528_n2088# 0.015615f
C181 source.n75 a_n1528_n2088# 0.036908f
C182 source.n76 a_n1528_n2088# 0.016534f
C183 source.n77 a_n1528_n2088# 0.124353f
C184 source.t6 a_n1528_n2088# 0.060156f
C185 source.n78 a_n1528_n2088# 0.027681f
C186 source.n79 a_n1528_n2088# 0.021801f
C187 source.n80 a_n1528_n2088# 0.015615f
C188 source.n81 a_n1528_n2088# 0.691434f
C189 source.n82 a_n1528_n2088# 0.029059f
C190 source.n83 a_n1528_n2088# 0.015615f
C191 source.n84 a_n1528_n2088# 0.016534f
C192 source.n85 a_n1528_n2088# 0.036908f
C193 source.n86 a_n1528_n2088# 0.036908f
C194 source.n87 a_n1528_n2088# 0.016534f
C195 source.n88 a_n1528_n2088# 0.015615f
C196 source.n89 a_n1528_n2088# 0.029059f
C197 source.n90 a_n1528_n2088# 0.029059f
C198 source.n91 a_n1528_n2088# 0.015615f
C199 source.n92 a_n1528_n2088# 0.016534f
C200 source.n93 a_n1528_n2088# 0.036908f
C201 source.n94 a_n1528_n2088# 0.079901f
C202 source.n95 a_n1528_n2088# 0.016534f
C203 source.n96 a_n1528_n2088# 0.015615f
C204 source.n97 a_n1528_n2088# 0.067169f
C205 source.n98 a_n1528_n2088# 0.044707f
C206 source.n99 a_n1528_n2088# 0.115628f
C207 source.t1 a_n1528_n2088# 0.13778f
C208 source.t8 a_n1528_n2088# 0.13778f
C209 source.n100 a_n1528_n2088# 1.07305f
C210 source.n101 a_n1528_n2088# 0.366037f
C211 source.t23 a_n1528_n2088# 0.13778f
C212 source.t5 a_n1528_n2088# 0.13778f
C213 source.n102 a_n1528_n2088# 1.07305f
C214 source.n103 a_n1528_n2088# 0.366037f
C215 source.n104 a_n1528_n2088# 0.040845f
C216 source.n105 a_n1528_n2088# 0.029059f
C217 source.n106 a_n1528_n2088# 0.015615f
C218 source.n107 a_n1528_n2088# 0.036908f
C219 source.n108 a_n1528_n2088# 0.016534f
C220 source.n109 a_n1528_n2088# 0.029059f
C221 source.n110 a_n1528_n2088# 0.015615f
C222 source.n111 a_n1528_n2088# 0.036908f
C223 source.n112 a_n1528_n2088# 0.016534f
C224 source.n113 a_n1528_n2088# 0.124353f
C225 source.t7 a_n1528_n2088# 0.060156f
C226 source.n114 a_n1528_n2088# 0.027681f
C227 source.n115 a_n1528_n2088# 0.021801f
C228 source.n116 a_n1528_n2088# 0.015615f
C229 source.n117 a_n1528_n2088# 0.691434f
C230 source.n118 a_n1528_n2088# 0.029059f
C231 source.n119 a_n1528_n2088# 0.015615f
C232 source.n120 a_n1528_n2088# 0.016534f
C233 source.n121 a_n1528_n2088# 0.036908f
C234 source.n122 a_n1528_n2088# 0.036908f
C235 source.n123 a_n1528_n2088# 0.016534f
C236 source.n124 a_n1528_n2088# 0.015615f
C237 source.n125 a_n1528_n2088# 0.029059f
C238 source.n126 a_n1528_n2088# 0.029059f
C239 source.n127 a_n1528_n2088# 0.015615f
C240 source.n128 a_n1528_n2088# 0.016534f
C241 source.n129 a_n1528_n2088# 0.036908f
C242 source.n130 a_n1528_n2088# 0.079901f
C243 source.n131 a_n1528_n2088# 0.016534f
C244 source.n132 a_n1528_n2088# 0.015615f
C245 source.n133 a_n1528_n2088# 0.067169f
C246 source.n134 a_n1528_n2088# 0.044707f
C247 source.n135 a_n1528_n2088# 1.0699f
C248 source.n136 a_n1528_n2088# 0.040845f
C249 source.n137 a_n1528_n2088# 0.029059f
C250 source.n138 a_n1528_n2088# 0.015615f
C251 source.n139 a_n1528_n2088# 0.036908f
C252 source.n140 a_n1528_n2088# 0.016534f
C253 source.n141 a_n1528_n2088# 0.029059f
C254 source.n142 a_n1528_n2088# 0.015615f
C255 source.n143 a_n1528_n2088# 0.036908f
C256 source.n144 a_n1528_n2088# 0.016534f
C257 source.n145 a_n1528_n2088# 0.124353f
C258 source.t14 a_n1528_n2088# 0.060156f
C259 source.n146 a_n1528_n2088# 0.027681f
C260 source.n147 a_n1528_n2088# 0.021801f
C261 source.n148 a_n1528_n2088# 0.015615f
C262 source.n149 a_n1528_n2088# 0.691434f
C263 source.n150 a_n1528_n2088# 0.029059f
C264 source.n151 a_n1528_n2088# 0.015615f
C265 source.n152 a_n1528_n2088# 0.016534f
C266 source.n153 a_n1528_n2088# 0.036908f
C267 source.n154 a_n1528_n2088# 0.036908f
C268 source.n155 a_n1528_n2088# 0.016534f
C269 source.n156 a_n1528_n2088# 0.015615f
C270 source.n157 a_n1528_n2088# 0.029059f
C271 source.n158 a_n1528_n2088# 0.029059f
C272 source.n159 a_n1528_n2088# 0.015615f
C273 source.n160 a_n1528_n2088# 0.016534f
C274 source.n161 a_n1528_n2088# 0.036908f
C275 source.n162 a_n1528_n2088# 0.079901f
C276 source.n163 a_n1528_n2088# 0.016534f
C277 source.n164 a_n1528_n2088# 0.015615f
C278 source.n165 a_n1528_n2088# 0.067169f
C279 source.n166 a_n1528_n2088# 0.044707f
C280 source.n167 a_n1528_n2088# 1.0699f
C281 source.t22 a_n1528_n2088# 0.13778f
C282 source.t12 a_n1528_n2088# 0.13778f
C283 source.n168 a_n1528_n2088# 1.07304f
C284 source.n169 a_n1528_n2088# 0.366044f
C285 source.t16 a_n1528_n2088# 0.13778f
C286 source.t17 a_n1528_n2088# 0.13778f
C287 source.n170 a_n1528_n2088# 1.07304f
C288 source.n171 a_n1528_n2088# 0.366044f
C289 source.n172 a_n1528_n2088# 0.040845f
C290 source.n173 a_n1528_n2088# 0.029059f
C291 source.n174 a_n1528_n2088# 0.015615f
C292 source.n175 a_n1528_n2088# 0.036908f
C293 source.n176 a_n1528_n2088# 0.016534f
C294 source.n177 a_n1528_n2088# 0.029059f
C295 source.n178 a_n1528_n2088# 0.015615f
C296 source.n179 a_n1528_n2088# 0.036908f
C297 source.n180 a_n1528_n2088# 0.016534f
C298 source.n181 a_n1528_n2088# 0.124353f
C299 source.t15 a_n1528_n2088# 0.060156f
C300 source.n182 a_n1528_n2088# 0.027681f
C301 source.n183 a_n1528_n2088# 0.021801f
C302 source.n184 a_n1528_n2088# 0.015615f
C303 source.n185 a_n1528_n2088# 0.691434f
C304 source.n186 a_n1528_n2088# 0.029059f
C305 source.n187 a_n1528_n2088# 0.015615f
C306 source.n188 a_n1528_n2088# 0.016534f
C307 source.n189 a_n1528_n2088# 0.036908f
C308 source.n190 a_n1528_n2088# 0.036908f
C309 source.n191 a_n1528_n2088# 0.016534f
C310 source.n192 a_n1528_n2088# 0.015615f
C311 source.n193 a_n1528_n2088# 0.029059f
C312 source.n194 a_n1528_n2088# 0.029059f
C313 source.n195 a_n1528_n2088# 0.015615f
C314 source.n196 a_n1528_n2088# 0.016534f
C315 source.n197 a_n1528_n2088# 0.036908f
C316 source.n198 a_n1528_n2088# 0.079901f
C317 source.n199 a_n1528_n2088# 0.016534f
C318 source.n200 a_n1528_n2088# 0.015615f
C319 source.n201 a_n1528_n2088# 0.067169f
C320 source.n202 a_n1528_n2088# 0.044707f
C321 source.n203 a_n1528_n2088# 0.115628f
C322 source.n204 a_n1528_n2088# 0.040845f
C323 source.n205 a_n1528_n2088# 0.029059f
C324 source.n206 a_n1528_n2088# 0.015615f
C325 source.n207 a_n1528_n2088# 0.036908f
C326 source.n208 a_n1528_n2088# 0.016534f
C327 source.n209 a_n1528_n2088# 0.029059f
C328 source.n210 a_n1528_n2088# 0.015615f
C329 source.n211 a_n1528_n2088# 0.036908f
C330 source.n212 a_n1528_n2088# 0.016534f
C331 source.n213 a_n1528_n2088# 0.124353f
C332 source.t2 a_n1528_n2088# 0.060156f
C333 source.n214 a_n1528_n2088# 0.027681f
C334 source.n215 a_n1528_n2088# 0.021801f
C335 source.n216 a_n1528_n2088# 0.015615f
C336 source.n217 a_n1528_n2088# 0.691434f
C337 source.n218 a_n1528_n2088# 0.029059f
C338 source.n219 a_n1528_n2088# 0.015615f
C339 source.n220 a_n1528_n2088# 0.016534f
C340 source.n221 a_n1528_n2088# 0.036908f
C341 source.n222 a_n1528_n2088# 0.036908f
C342 source.n223 a_n1528_n2088# 0.016534f
C343 source.n224 a_n1528_n2088# 0.015615f
C344 source.n225 a_n1528_n2088# 0.029059f
C345 source.n226 a_n1528_n2088# 0.029059f
C346 source.n227 a_n1528_n2088# 0.015615f
C347 source.n228 a_n1528_n2088# 0.016534f
C348 source.n229 a_n1528_n2088# 0.036908f
C349 source.n230 a_n1528_n2088# 0.079901f
C350 source.n231 a_n1528_n2088# 0.016534f
C351 source.n232 a_n1528_n2088# 0.015615f
C352 source.n233 a_n1528_n2088# 0.067169f
C353 source.n234 a_n1528_n2088# 0.044707f
C354 source.n235 a_n1528_n2088# 0.115628f
C355 source.t10 a_n1528_n2088# 0.13778f
C356 source.t9 a_n1528_n2088# 0.13778f
C357 source.n236 a_n1528_n2088# 1.07304f
C358 source.n237 a_n1528_n2088# 0.366044f
C359 source.t3 a_n1528_n2088# 0.13778f
C360 source.t4 a_n1528_n2088# 0.13778f
C361 source.n238 a_n1528_n2088# 1.07304f
C362 source.n239 a_n1528_n2088# 0.366044f
C363 source.n240 a_n1528_n2088# 0.040845f
C364 source.n241 a_n1528_n2088# 0.029059f
C365 source.n242 a_n1528_n2088# 0.015615f
C366 source.n243 a_n1528_n2088# 0.036908f
C367 source.n244 a_n1528_n2088# 0.016534f
C368 source.n245 a_n1528_n2088# 0.029059f
C369 source.n246 a_n1528_n2088# 0.015615f
C370 source.n247 a_n1528_n2088# 0.036908f
C371 source.n248 a_n1528_n2088# 0.016534f
C372 source.n249 a_n1528_n2088# 0.124353f
C373 source.t0 a_n1528_n2088# 0.060156f
C374 source.n250 a_n1528_n2088# 0.027681f
C375 source.n251 a_n1528_n2088# 0.021801f
C376 source.n252 a_n1528_n2088# 0.015615f
C377 source.n253 a_n1528_n2088# 0.691434f
C378 source.n254 a_n1528_n2088# 0.029059f
C379 source.n255 a_n1528_n2088# 0.015615f
C380 source.n256 a_n1528_n2088# 0.016534f
C381 source.n257 a_n1528_n2088# 0.036908f
C382 source.n258 a_n1528_n2088# 0.036908f
C383 source.n259 a_n1528_n2088# 0.016534f
C384 source.n260 a_n1528_n2088# 0.015615f
C385 source.n261 a_n1528_n2088# 0.029059f
C386 source.n262 a_n1528_n2088# 0.029059f
C387 source.n263 a_n1528_n2088# 0.015615f
C388 source.n264 a_n1528_n2088# 0.016534f
C389 source.n265 a_n1528_n2088# 0.036908f
C390 source.n266 a_n1528_n2088# 0.079901f
C391 source.n267 a_n1528_n2088# 0.016534f
C392 source.n268 a_n1528_n2088# 0.015615f
C393 source.n269 a_n1528_n2088# 0.067169f
C394 source.n270 a_n1528_n2088# 0.044707f
C395 source.n271 a_n1528_n2088# 0.276436f
C396 source.n272 a_n1528_n2088# 1.18709f
C397 plus.n0 a_n1528_n2088# 0.055835f
C398 plus.t6 a_n1528_n2088# 0.238625f
C399 plus.t0 a_n1528_n2088# 0.238625f
C400 plus.n1 a_n1528_n2088# 0.019899f
C401 plus.t3 a_n1528_n2088# 0.243037f
C402 plus.n2 a_n1528_n2088# 0.127617f
C403 plus.t1 a_n1528_n2088# 0.238625f
C404 plus.n3 a_n1528_n2088# 0.112402f
C405 plus.t7 a_n1528_n2088# 0.238625f
C406 plus.n4 a_n1528_n2088# 0.112402f
C407 plus.n5 a_n1528_n2088# 0.021276f
C408 plus.n6 a_n1528_n2088# 0.116762f
C409 plus.n7 a_n1528_n2088# 0.055835f
C410 plus.n8 a_n1528_n2088# 0.055835f
C411 plus.n9 a_n1528_n2088# 0.019899f
C412 plus.n10 a_n1528_n2088# 0.112402f
C413 plus.n11 a_n1528_n2088# 0.021276f
C414 plus.n12 a_n1528_n2088# 0.112402f
C415 plus.t11 a_n1528_n2088# 0.243037f
C416 plus.n13 a_n1528_n2088# 0.127545f
C417 plus.n14 a_n1528_n2088# 0.46966f
C418 plus.n15 a_n1528_n2088# 0.055835f
C419 plus.t5 a_n1528_n2088# 0.243037f
C420 plus.t10 a_n1528_n2088# 0.238625f
C421 plus.t9 a_n1528_n2088# 0.238625f
C422 plus.n16 a_n1528_n2088# 0.019899f
C423 plus.t8 a_n1528_n2088# 0.243037f
C424 plus.n17 a_n1528_n2088# 0.127617f
C425 plus.t2 a_n1528_n2088# 0.238625f
C426 plus.n18 a_n1528_n2088# 0.112402f
C427 plus.t4 a_n1528_n2088# 0.238625f
C428 plus.n19 a_n1528_n2088# 0.112402f
C429 plus.n20 a_n1528_n2088# 0.021276f
C430 plus.n21 a_n1528_n2088# 0.116762f
C431 plus.n22 a_n1528_n2088# 0.055835f
C432 plus.n23 a_n1528_n2088# 0.055835f
C433 plus.n24 a_n1528_n2088# 0.019899f
C434 plus.n25 a_n1528_n2088# 0.112402f
C435 plus.n26 a_n1528_n2088# 0.021276f
C436 plus.n27 a_n1528_n2088# 0.112402f
C437 plus.n28 a_n1528_n2088# 0.127545f
C438 plus.n29 a_n1528_n2088# 1.33139f
.ends

