* NGSPICE file created from diffpair206.ext - technology: sky130A

.subckt diffpair206 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t25 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X1 a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X2 drain_right.t12 minus.t1 source.t20 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X3 source.t23 minus.t2 drain_right.t11 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X4 drain_left.t13 plus.t0 source.t8 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X5 drain_left.t12 plus.t1 source.t4 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X6 drain_right.t10 minus.t3 source.t24 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 drain_right.t9 minus.t4 source.t15 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X8 source.t16 minus.t5 drain_right.t8 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X9 drain_left.t11 plus.t2 source.t6 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X10 drain_right.t7 minus.t6 source.t17 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X11 source.t10 plus.t3 drain_left.t10 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X12 source.t18 minus.t7 drain_right.t6 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X13 a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X14 source.t22 minus.t8 drain_right.t5 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X15 source.t0 plus.t4 drain_left.t9 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X16 drain_left.t8 plus.t5 source.t11 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X17 source.t14 minus.t9 drain_right.t4 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X18 a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X19 source.t1 plus.t6 drain_left.t7 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X20 a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X21 drain_right.t3 minus.t10 source.t26 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X22 source.t5 plus.t7 drain_left.t6 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X23 drain_left.t5 plus.t8 source.t9 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X24 drain_right.t2 minus.t11 source.t19 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X25 source.t2 plus.t9 drain_left.t4 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X26 drain_right.t1 minus.t12 source.t27 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X27 source.t21 minus.t13 drain_right.t0 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X28 drain_left.t3 plus.t10 source.t13 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X29 drain_left.t2 plus.t11 source.t12 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X30 drain_left.t1 plus.t12 source.t3 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X31 source.t7 plus.t13 drain_left.t0 a_n2044_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
R0 minus.n4 minus.t11 244.149
R1 minus.n20 minus.t3 244.149
R2 minus.n3 minus.t2 223.167
R3 minus.n7 minus.t6 223.167
R4 minus.n8 minus.t13 223.167
R5 minus.n1 minus.t4 223.167
R6 minus.n13 minus.t9 223.167
R7 minus.n14 minus.t0 223.167
R8 minus.n19 minus.t7 223.167
R9 minus.n23 minus.t1 223.167
R10 minus.n24 minus.t5 223.167
R11 minus.n17 minus.t12 223.167
R12 minus.n29 minus.t8 223.167
R13 minus.n30 minus.t10 223.167
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n0 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n1 161.3
R18 minus.n7 minus.n2 161.3
R19 minus.n6 minus.n5 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n16 161.3
R22 minus.n28 minus.n27 161.3
R23 minus.n26 minus.n17 161.3
R24 minus.n23 minus.n18 161.3
R25 minus.n22 minus.n21 161.3
R26 minus.n9 minus.n8 80.6037
R27 minus.n25 minus.n24 80.6037
R28 minus.n5 minus.n4 70.4033
R29 minus.n21 minus.n20 70.4033
R30 minus.n8 minus.n7 48.2005
R31 minus.n8 minus.n1 48.2005
R32 minus.n14 minus.n13 48.2005
R33 minus.n24 minus.n23 48.2005
R34 minus.n24 minus.n17 48.2005
R35 minus.n30 minus.n29 48.2005
R36 minus.n32 minus.n15 30.1388
R37 minus.n7 minus.n6 24.8308
R38 minus.n12 minus.n1 24.8308
R39 minus.n23 minus.n22 24.8308
R40 minus.n28 minus.n17 24.8308
R41 minus.n6 minus.n3 23.3702
R42 minus.n13 minus.n12 23.3702
R43 minus.n22 minus.n19 23.3702
R44 minus.n29 minus.n28 23.3702
R45 minus.n4 minus.n3 20.9576
R46 minus.n20 minus.n19 20.9576
R47 minus.n32 minus.n31 6.5933
R48 minus.n10 minus.n9 0.285035
R49 minus.n9 minus.n2 0.285035
R50 minus.n25 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n5 minus.n2 0.189894
R56 minus.n21 minus.n18 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n16 0.189894
R59 minus.n31 minus.n16 0.189894
R60 minus minus.n32 0.188
R61 source.n0 source.t11 69.6943
R62 source.n7 source.t19 69.6943
R63 source.n27 source.t26 69.6942
R64 source.n20 source.t6 69.6942
R65 source.n2 source.n1 63.0943
R66 source.n4 source.n3 63.0943
R67 source.n6 source.n5 63.0943
R68 source.n9 source.n8 63.0943
R69 source.n11 source.n10 63.0943
R70 source.n13 source.n12 63.0943
R71 source.n26 source.n25 63.0942
R72 source.n24 source.n23 63.0942
R73 source.n22 source.n21 63.0942
R74 source.n19 source.n18 63.0942
R75 source.n17 source.n16 63.0942
R76 source.n15 source.n14 63.0942
R77 source.n15 source.n13 15.9006
R78 source.n28 source.n0 9.56437
R79 source.n25 source.t27 6.6005
R80 source.n25 source.t22 6.6005
R81 source.n23 source.t20 6.6005
R82 source.n23 source.t16 6.6005
R83 source.n21 source.t24 6.6005
R84 source.n21 source.t18 6.6005
R85 source.n18 source.t8 6.6005
R86 source.n18 source.t1 6.6005
R87 source.n16 source.t13 6.6005
R88 source.n16 source.t5 6.6005
R89 source.n14 source.t9 6.6005
R90 source.n14 source.t0 6.6005
R91 source.n1 source.t12 6.6005
R92 source.n1 source.t7 6.6005
R93 source.n3 source.t3 6.6005
R94 source.n3 source.t10 6.6005
R95 source.n5 source.t4 6.6005
R96 source.n5 source.t2 6.6005
R97 source.n8 source.t17 6.6005
R98 source.n8 source.t23 6.6005
R99 source.n10 source.t15 6.6005
R100 source.n10 source.t21 6.6005
R101 source.n12 source.t25 6.6005
R102 source.n12 source.t14 6.6005
R103 source.n28 source.n27 5.62119
R104 source.n7 source.n6 0.828086
R105 source.n22 source.n20 0.828086
R106 source.n13 source.n11 0.716017
R107 source.n11 source.n9 0.716017
R108 source.n9 source.n7 0.716017
R109 source.n6 source.n4 0.716017
R110 source.n4 source.n2 0.716017
R111 source.n2 source.n0 0.716017
R112 source.n17 source.n15 0.716017
R113 source.n19 source.n17 0.716017
R114 source.n20 source.n19 0.716017
R115 source.n24 source.n22 0.716017
R116 source.n26 source.n24 0.716017
R117 source.n27 source.n26 0.716017
R118 source source.n28 0.188
R119 drain_right.n1 drain_right.t10 87.0885
R120 drain_right.n11 drain_right.t13 86.3731
R121 drain_right.n8 drain_right.n6 80.4886
R122 drain_right.n4 drain_right.n2 80.4885
R123 drain_right.n8 drain_right.n7 79.7731
R124 drain_right.n10 drain_right.n9 79.7731
R125 drain_right.n4 drain_right.n3 79.773
R126 drain_right.n1 drain_right.n0 79.773
R127 drain_right drain_right.n5 24.1099
R128 drain_right.n2 drain_right.t5 6.6005
R129 drain_right.n2 drain_right.t3 6.6005
R130 drain_right.n3 drain_right.t8 6.6005
R131 drain_right.n3 drain_right.t1 6.6005
R132 drain_right.n0 drain_right.t6 6.6005
R133 drain_right.n0 drain_right.t12 6.6005
R134 drain_right.n6 drain_right.t11 6.6005
R135 drain_right.n6 drain_right.t2 6.6005
R136 drain_right.n7 drain_right.t0 6.6005
R137 drain_right.n7 drain_right.t7 6.6005
R138 drain_right.n9 drain_right.t4 6.6005
R139 drain_right.n9 drain_right.t9 6.6005
R140 drain_right drain_right.n11 6.01097
R141 drain_right.n11 drain_right.n10 0.716017
R142 drain_right.n10 drain_right.n8 0.716017
R143 drain_right.n5 drain_right.n1 0.481792
R144 drain_right.n5 drain_right.n4 0.124033
R145 plus.n4 plus.t1 244.149
R146 plus.n20 plus.t2 244.149
R147 plus.n14 plus.t5 223.167
R148 plus.n13 plus.t13 223.167
R149 plus.n1 plus.t11 223.167
R150 plus.n8 plus.t3 223.167
R151 plus.n7 plus.t12 223.167
R152 plus.n3 plus.t9 223.167
R153 plus.n30 plus.t8 223.167
R154 plus.n29 plus.t4 223.167
R155 plus.n17 plus.t10 223.167
R156 plus.n24 plus.t7 223.167
R157 plus.n23 plus.t0 223.167
R158 plus.n19 plus.t6 223.167
R159 plus.n6 plus.n5 161.3
R160 plus.n7 plus.n2 161.3
R161 plus.n10 plus.n1 161.3
R162 plus.n12 plus.n11 161.3
R163 plus.n13 plus.n0 161.3
R164 plus.n15 plus.n14 161.3
R165 plus.n22 plus.n21 161.3
R166 plus.n23 plus.n18 161.3
R167 plus.n26 plus.n17 161.3
R168 plus.n28 plus.n27 161.3
R169 plus.n29 plus.n16 161.3
R170 plus.n31 plus.n30 161.3
R171 plus.n9 plus.n8 80.6037
R172 plus.n25 plus.n24 80.6037
R173 plus.n5 plus.n4 70.4033
R174 plus.n21 plus.n20 70.4033
R175 plus.n14 plus.n13 48.2005
R176 plus.n8 plus.n1 48.2005
R177 plus.n8 plus.n7 48.2005
R178 plus.n30 plus.n29 48.2005
R179 plus.n24 plus.n17 48.2005
R180 plus.n24 plus.n23 48.2005
R181 plus plus.n31 27.4289
R182 plus.n12 plus.n1 24.8308
R183 plus.n7 plus.n6 24.8308
R184 plus.n28 plus.n17 24.8308
R185 plus.n23 plus.n22 24.8308
R186 plus.n13 plus.n12 23.3702
R187 plus.n6 plus.n3 23.3702
R188 plus.n29 plus.n28 23.3702
R189 plus.n22 plus.n19 23.3702
R190 plus.n4 plus.n3 20.9576
R191 plus.n20 plus.n19 20.9576
R192 plus plus.n15 8.82815
R193 plus.n9 plus.n2 0.285035
R194 plus.n10 plus.n9 0.285035
R195 plus.n26 plus.n25 0.285035
R196 plus.n25 plus.n18 0.285035
R197 plus.n5 plus.n2 0.189894
R198 plus.n11 plus.n10 0.189894
R199 plus.n11 plus.n0 0.189894
R200 plus.n15 plus.n0 0.189894
R201 plus.n31 plus.n16 0.189894
R202 plus.n27 plus.n16 0.189894
R203 plus.n27 plus.n26 0.189894
R204 plus.n21 plus.n18 0.189894
R205 drain_left.n7 drain_left.t12 87.0886
R206 drain_left.n1 drain_left.t5 87.0885
R207 drain_left.n4 drain_left.n2 80.4885
R208 drain_left.n11 drain_left.n10 79.7731
R209 drain_left.n9 drain_left.n8 79.7731
R210 drain_left.n7 drain_left.n6 79.7731
R211 drain_left.n4 drain_left.n3 79.773
R212 drain_left.n1 drain_left.n0 79.773
R213 drain_left drain_left.n5 24.6631
R214 drain_left.n2 drain_left.t7 6.6005
R215 drain_left.n2 drain_left.t11 6.6005
R216 drain_left.n3 drain_left.t6 6.6005
R217 drain_left.n3 drain_left.t13 6.6005
R218 drain_left.n0 drain_left.t9 6.6005
R219 drain_left.n0 drain_left.t3 6.6005
R220 drain_left.n10 drain_left.t0 6.6005
R221 drain_left.n10 drain_left.t8 6.6005
R222 drain_left.n8 drain_left.t10 6.6005
R223 drain_left.n8 drain_left.t2 6.6005
R224 drain_left.n6 drain_left.t4 6.6005
R225 drain_left.n6 drain_left.t1 6.6005
R226 drain_left drain_left.n11 6.36873
R227 drain_left.n9 drain_left.n7 0.716017
R228 drain_left.n11 drain_left.n9 0.716017
R229 drain_left.n5 drain_left.n1 0.481792
R230 drain_left.n5 drain_left.n4 0.124033
C0 drain_left plus 2.43735f
C1 plus minus 4.03581f
C2 plus source 2.5421f
C3 drain_right drain_left 1.05608f
C4 drain_right minus 2.23818f
C5 drain_left minus 0.177607f
C6 drain_right source 7.66105f
C7 drain_left source 7.662951f
C8 source minus 2.52796f
C9 drain_right plus 0.361665f
C10 drain_right a_n2044_n1488# 4.71377f
C11 drain_left a_n2044_n1488# 5.037f
C12 source a_n2044_n1488# 3.048583f
C13 minus a_n2044_n1488# 7.314109f
C14 plus a_n2044_n1488# 8.628071f
C15 drain_left.t5 a_n2044_n1488# 0.590311f
C16 drain_left.t9 a_n2044_n1488# 0.063482f
C17 drain_left.t3 a_n2044_n1488# 0.063482f
C18 drain_left.n0 a_n2044_n1488# 0.457827f
C19 drain_left.n1 a_n2044_n1488# 0.646436f
C20 drain_left.t7 a_n2044_n1488# 0.063482f
C21 drain_left.t11 a_n2044_n1488# 0.063482f
C22 drain_left.n2 a_n2044_n1488# 0.460927f
C23 drain_left.t6 a_n2044_n1488# 0.063482f
C24 drain_left.t13 a_n2044_n1488# 0.063482f
C25 drain_left.n3 a_n2044_n1488# 0.457827f
C26 drain_left.n4 a_n2044_n1488# 0.637292f
C27 drain_left.n5 a_n2044_n1488# 0.873823f
C28 drain_left.t12 a_n2044_n1488# 0.590313f
C29 drain_left.t4 a_n2044_n1488# 0.063482f
C30 drain_left.t1 a_n2044_n1488# 0.063482f
C31 drain_left.n6 a_n2044_n1488# 0.45783f
C32 drain_left.n7 a_n2044_n1488# 0.665352f
C33 drain_left.t10 a_n2044_n1488# 0.063482f
C34 drain_left.t2 a_n2044_n1488# 0.063482f
C35 drain_left.n8 a_n2044_n1488# 0.45783f
C36 drain_left.n9 a_n2044_n1488# 0.337827f
C37 drain_left.t0 a_n2044_n1488# 0.063482f
C38 drain_left.t8 a_n2044_n1488# 0.063482f
C39 drain_left.n10 a_n2044_n1488# 0.45783f
C40 drain_left.n11 a_n2044_n1488# 0.567887f
C41 plus.n0 a_n2044_n1488# 0.047967f
C42 plus.t5 a_n2044_n1488# 0.215756f
C43 plus.t13 a_n2044_n1488# 0.215756f
C44 plus.t11 a_n2044_n1488# 0.215756f
C45 plus.n1 a_n2044_n1488# 0.134432f
C46 plus.n2 a_n2044_n1488# 0.064007f
C47 plus.t3 a_n2044_n1488# 0.215756f
C48 plus.t12 a_n2044_n1488# 0.215756f
C49 plus.t9 a_n2044_n1488# 0.215756f
C50 plus.n3 a_n2044_n1488# 0.134137f
C51 plus.t1 a_n2044_n1488# 0.226883f
C52 plus.n4 a_n2044_n1488# 0.118647f
C53 plus.n5 a_n2044_n1488# 0.157729f
C54 plus.n6 a_n2044_n1488# 0.010885f
C55 plus.n7 a_n2044_n1488# 0.134432f
C56 plus.n8 a_n2044_n1488# 0.14029f
C57 plus.n9 a_n2044_n1488# 0.063857f
C58 plus.n10 a_n2044_n1488# 0.064007f
C59 plus.n11 a_n2044_n1488# 0.047967f
C60 plus.n12 a_n2044_n1488# 0.010885f
C61 plus.n13 a_n2044_n1488# 0.134137f
C62 plus.n14 a_n2044_n1488# 0.129405f
C63 plus.n15 a_n2044_n1488# 0.369367f
C64 plus.n16 a_n2044_n1488# 0.047967f
C65 plus.t8 a_n2044_n1488# 0.215756f
C66 plus.t4 a_n2044_n1488# 0.215756f
C67 plus.t10 a_n2044_n1488# 0.215756f
C68 plus.n17 a_n2044_n1488# 0.134432f
C69 plus.n18 a_n2044_n1488# 0.064007f
C70 plus.t7 a_n2044_n1488# 0.215756f
C71 plus.t0 a_n2044_n1488# 0.215756f
C72 plus.t6 a_n2044_n1488# 0.215756f
C73 plus.n19 a_n2044_n1488# 0.134137f
C74 plus.t2 a_n2044_n1488# 0.226883f
C75 plus.n20 a_n2044_n1488# 0.118647f
C76 plus.n21 a_n2044_n1488# 0.157729f
C77 plus.n22 a_n2044_n1488# 0.010885f
C78 plus.n23 a_n2044_n1488# 0.134432f
C79 plus.n24 a_n2044_n1488# 0.14029f
C80 plus.n25 a_n2044_n1488# 0.063857f
C81 plus.n26 a_n2044_n1488# 0.064007f
C82 plus.n27 a_n2044_n1488# 0.047967f
C83 plus.n28 a_n2044_n1488# 0.010885f
C84 plus.n29 a_n2044_n1488# 0.134137f
C85 plus.n30 a_n2044_n1488# 0.129405f
C86 plus.n31 a_n2044_n1488# 1.18621f
C87 drain_right.t10 a_n2044_n1488# 0.584686f
C88 drain_right.t6 a_n2044_n1488# 0.062877f
C89 drain_right.t12 a_n2044_n1488# 0.062877f
C90 drain_right.n0 a_n2044_n1488# 0.453465f
C91 drain_right.n1 a_n2044_n1488# 0.640276f
C92 drain_right.t5 a_n2044_n1488# 0.062877f
C93 drain_right.t3 a_n2044_n1488# 0.062877f
C94 drain_right.n2 a_n2044_n1488# 0.456534f
C95 drain_right.t8 a_n2044_n1488# 0.062877f
C96 drain_right.t1 a_n2044_n1488# 0.062877f
C97 drain_right.n3 a_n2044_n1488# 0.453465f
C98 drain_right.n4 a_n2044_n1488# 0.631219f
C99 drain_right.n5 a_n2044_n1488# 0.81307f
C100 drain_right.t11 a_n2044_n1488# 0.062877f
C101 drain_right.t2 a_n2044_n1488# 0.062877f
C102 drain_right.n6 a_n2044_n1488# 0.456536f
C103 drain_right.t0 a_n2044_n1488# 0.062877f
C104 drain_right.t7 a_n2044_n1488# 0.062877f
C105 drain_right.n7 a_n2044_n1488# 0.453467f
C106 drain_right.n8 a_n2044_n1488# 0.676829f
C107 drain_right.t4 a_n2044_n1488# 0.062877f
C108 drain_right.t9 a_n2044_n1488# 0.062877f
C109 drain_right.n9 a_n2044_n1488# 0.453467f
C110 drain_right.n10 a_n2044_n1488# 0.334608f
C111 drain_right.t13 a_n2044_n1488# 0.582001f
C112 drain_right.n11 a_n2044_n1488# 0.559659f
C113 source.t11 a_n2044_n1488# 0.629542f
C114 source.n0 a_n2044_n1488# 0.890155f
C115 source.t12 a_n2044_n1488# 0.075814f
C116 source.t7 a_n2044_n1488# 0.075814f
C117 source.n1 a_n2044_n1488# 0.480701f
C118 source.n2 a_n2044_n1488# 0.426044f
C119 source.t3 a_n2044_n1488# 0.075814f
C120 source.t10 a_n2044_n1488# 0.075814f
C121 source.n3 a_n2044_n1488# 0.480701f
C122 source.n4 a_n2044_n1488# 0.426044f
C123 source.t4 a_n2044_n1488# 0.075814f
C124 source.t2 a_n2044_n1488# 0.075814f
C125 source.n5 a_n2044_n1488# 0.480701f
C126 source.n6 a_n2044_n1488# 0.437592f
C127 source.t19 a_n2044_n1488# 0.629542f
C128 source.n7 a_n2044_n1488# 0.495515f
C129 source.t17 a_n2044_n1488# 0.075814f
C130 source.t23 a_n2044_n1488# 0.075814f
C131 source.n8 a_n2044_n1488# 0.480701f
C132 source.n9 a_n2044_n1488# 0.426044f
C133 source.t15 a_n2044_n1488# 0.075814f
C134 source.t21 a_n2044_n1488# 0.075814f
C135 source.n10 a_n2044_n1488# 0.480701f
C136 source.n11 a_n2044_n1488# 0.426044f
C137 source.t25 a_n2044_n1488# 0.075814f
C138 source.t14 a_n2044_n1488# 0.075814f
C139 source.n12 a_n2044_n1488# 0.480701f
C140 source.n13 a_n2044_n1488# 1.24359f
C141 source.t9 a_n2044_n1488# 0.075814f
C142 source.t0 a_n2044_n1488# 0.075814f
C143 source.n14 a_n2044_n1488# 0.480698f
C144 source.n15 a_n2044_n1488# 1.24359f
C145 source.t13 a_n2044_n1488# 0.075814f
C146 source.t5 a_n2044_n1488# 0.075814f
C147 source.n16 a_n2044_n1488# 0.480698f
C148 source.n17 a_n2044_n1488# 0.426047f
C149 source.t8 a_n2044_n1488# 0.075814f
C150 source.t1 a_n2044_n1488# 0.075814f
C151 source.n18 a_n2044_n1488# 0.480698f
C152 source.n19 a_n2044_n1488# 0.426047f
C153 source.t6 a_n2044_n1488# 0.629539f
C154 source.n20 a_n2044_n1488# 0.495519f
C155 source.t24 a_n2044_n1488# 0.075814f
C156 source.t18 a_n2044_n1488# 0.075814f
C157 source.n21 a_n2044_n1488# 0.480698f
C158 source.n22 a_n2044_n1488# 0.437595f
C159 source.t20 a_n2044_n1488# 0.075814f
C160 source.t16 a_n2044_n1488# 0.075814f
C161 source.n23 a_n2044_n1488# 0.480698f
C162 source.n24 a_n2044_n1488# 0.426047f
C163 source.t27 a_n2044_n1488# 0.075814f
C164 source.t22 a_n2044_n1488# 0.075814f
C165 source.n25 a_n2044_n1488# 0.480698f
C166 source.n26 a_n2044_n1488# 0.426047f
C167 source.t26 a_n2044_n1488# 0.629539f
C168 source.n27 a_n2044_n1488# 0.653296f
C169 source.n28 a_n2044_n1488# 0.934863f
C170 minus.n0 a_n2044_n1488# 0.046384f
C171 minus.t4 a_n2044_n1488# 0.208633f
C172 minus.n1 a_n2044_n1488# 0.129995f
C173 minus.n2 a_n2044_n1488# 0.061894f
C174 minus.t2 a_n2044_n1488# 0.208633f
C175 minus.n3 a_n2044_n1488# 0.129709f
C176 minus.t11 a_n2044_n1488# 0.219393f
C177 minus.n4 a_n2044_n1488# 0.11473f
C178 minus.n5 a_n2044_n1488# 0.152522f
C179 minus.n6 a_n2044_n1488# 0.010526f
C180 minus.t6 a_n2044_n1488# 0.208633f
C181 minus.n7 a_n2044_n1488# 0.129995f
C182 minus.t13 a_n2044_n1488# 0.208633f
C183 minus.n8 a_n2044_n1488# 0.135659f
C184 minus.n9 a_n2044_n1488# 0.061749f
C185 minus.n10 a_n2044_n1488# 0.061894f
C186 minus.n11 a_n2044_n1488# 0.046384f
C187 minus.n12 a_n2044_n1488# 0.010526f
C188 minus.t9 a_n2044_n1488# 0.208633f
C189 minus.n13 a_n2044_n1488# 0.129709f
C190 minus.t0 a_n2044_n1488# 0.208633f
C191 minus.n14 a_n2044_n1488# 0.125133f
C192 minus.n15 a_n2044_n1488# 1.22019f
C193 minus.n16 a_n2044_n1488# 0.046384f
C194 minus.t12 a_n2044_n1488# 0.208633f
C195 minus.n17 a_n2044_n1488# 0.129995f
C196 minus.n18 a_n2044_n1488# 0.061894f
C197 minus.t7 a_n2044_n1488# 0.208633f
C198 minus.n19 a_n2044_n1488# 0.129709f
C199 minus.t3 a_n2044_n1488# 0.219393f
C200 minus.n20 a_n2044_n1488# 0.11473f
C201 minus.n21 a_n2044_n1488# 0.152522f
C202 minus.n22 a_n2044_n1488# 0.010526f
C203 minus.t1 a_n2044_n1488# 0.208633f
C204 minus.n23 a_n2044_n1488# 0.129995f
C205 minus.t5 a_n2044_n1488# 0.208633f
C206 minus.n24 a_n2044_n1488# 0.135659f
C207 minus.n25 a_n2044_n1488# 0.061749f
C208 minus.n26 a_n2044_n1488# 0.061894f
C209 minus.n27 a_n2044_n1488# 0.046384f
C210 minus.n28 a_n2044_n1488# 0.010526f
C211 minus.t8 a_n2044_n1488# 0.208633f
C212 minus.n29 a_n2044_n1488# 0.129709f
C213 minus.t10 a_n2044_n1488# 0.208633f
C214 minus.n30 a_n2044_n1488# 0.125133f
C215 minus.n31 a_n2044_n1488# 0.313398f
C216 minus.n32 a_n2044_n1488# 1.49996f
.ends

