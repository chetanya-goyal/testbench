* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X1 drain_right.t9 minus.t0 source.t18 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X2 source.t13 minus.t1 drain_right.t8 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t5 plus.t0 drain_left.t9 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 drain_right.t7 minus.t2 source.t14 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 source.t2 plus.t1 drain_left.t8 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X6 a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X7 source.t9 plus.t2 drain_left.t7 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X8 drain_left.t6 plus.t3 source.t8 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X9 source.t15 minus.t3 drain_right.t6 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X10 drain_left.t5 plus.t4 source.t3 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X11 drain_right.t5 minus.t4 source.t17 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 drain_left.t4 plus.t5 source.t4 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X13 drain_right.t4 minus.t5 source.t19 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X14 drain_right.t3 minus.t6 source.t16 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X15 a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X16 drain_left.t3 plus.t6 source.t6 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X17 source.t0 plus.t7 drain_left.t2 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X18 source.t10 minus.t7 drain_right.t2 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X19 source.t11 minus.t8 drain_right.t1 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X20 a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X21 drain_right.t0 minus.t9 source.t12 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X22 drain_left.t1 plus.t8 source.t1 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X23 drain_left.t0 plus.t9 source.t7 a_n1352_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 minus.n8 minus.t6 442.93
R1 minus.n2 minus.t5 442.93
R2 minus.n18 minus.t0 442.93
R3 minus.n12 minus.t9 442.93
R4 minus.n7 minus.t8 397.651
R5 minus.n5 minus.t2 397.651
R6 minus.n1 minus.t3 397.651
R7 minus.n17 minus.t7 397.651
R8 minus.n15 minus.t4 397.651
R9 minus.n11 minus.t1 397.651
R10 minus.n3 minus.n2 161.489
R11 minus.n13 minus.n12 161.489
R12 minus.n9 minus.n8 161.3
R13 minus.n6 minus.n0 161.3
R14 minus.n4 minus.n3 161.3
R15 minus.n19 minus.n18 161.3
R16 minus.n16 minus.n10 161.3
R17 minus.n14 minus.n13 161.3
R18 minus.n7 minus.n6 40.8975
R19 minus.n4 minus.n1 40.8975
R20 minus.n14 minus.n11 40.8975
R21 minus.n17 minus.n16 40.8975
R22 minus.n6 minus.n5 36.5157
R23 minus.n5 minus.n4 36.5157
R24 minus.n15 minus.n14 36.5157
R25 minus.n16 minus.n15 36.5157
R26 minus.n8 minus.n7 32.1338
R27 minus.n2 minus.n1 32.1338
R28 minus.n12 minus.n11 32.1338
R29 minus.n18 minus.n17 32.1338
R30 minus.n20 minus.n9 26.616
R31 minus.n20 minus.n19 6.44936
R32 minus.n9 minus.n0 0.189894
R33 minus.n3 minus.n0 0.189894
R34 minus.n13 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n42 source.n40 289.615
R38 source.n30 source.n28 289.615
R39 source.n2 source.n0 289.615
R40 source.n14 source.n12 289.615
R41 source.n43 source.n42 185
R42 source.n31 source.n30 185
R43 source.n3 source.n2 185
R44 source.n15 source.n14 185
R45 source.t18 source.n41 167.117
R46 source.t1 source.n29 167.117
R47 source.t6 source.n1 167.117
R48 source.t19 source.n13 167.117
R49 source.n9 source.n8 84.1169
R50 source.n11 source.n10 84.1169
R51 source.n21 source.n20 84.1169
R52 source.n23 source.n22 84.1169
R53 source.n39 source.n38 84.1168
R54 source.n37 source.n36 84.1168
R55 source.n27 source.n26 84.1168
R56 source.n25 source.n24 84.1168
R57 source.n42 source.t18 52.3082
R58 source.n30 source.t1 52.3082
R59 source.n2 source.t6 52.3082
R60 source.n14 source.t19 52.3082
R61 source.n47 source.n46 31.4096
R62 source.n35 source.n34 31.4096
R63 source.n7 source.n6 31.4096
R64 source.n19 source.n18 31.4096
R65 source.n25 source.n23 14.6258
R66 source.n38 source.t17 9.9005
R67 source.n38 source.t10 9.9005
R68 source.n36 source.t12 9.9005
R69 source.n36 source.t13 9.9005
R70 source.n26 source.t4 9.9005
R71 source.n26 source.t2 9.9005
R72 source.n24 source.t8 9.9005
R73 source.n24 source.t5 9.9005
R74 source.n8 source.t7 9.9005
R75 source.n8 source.t0 9.9005
R76 source.n10 source.t3 9.9005
R77 source.n10 source.t9 9.9005
R78 source.n20 source.t14 9.9005
R79 source.n20 source.t15 9.9005
R80 source.n22 source.t16 9.9005
R81 source.n22 source.t11 9.9005
R82 source.n43 source.n41 9.71174
R83 source.n31 source.n29 9.71174
R84 source.n3 source.n1 9.71174
R85 source.n15 source.n13 9.71174
R86 source.n46 source.n45 9.45567
R87 source.n34 source.n33 9.45567
R88 source.n6 source.n5 9.45567
R89 source.n18 source.n17 9.45567
R90 source.n45 source.n44 9.3005
R91 source.n33 source.n32 9.3005
R92 source.n5 source.n4 9.3005
R93 source.n17 source.n16 9.3005
R94 source.n48 source.n7 8.67749
R95 source.n46 source.n40 8.14595
R96 source.n34 source.n28 8.14595
R97 source.n6 source.n0 8.14595
R98 source.n18 source.n12 8.14595
R99 source.n44 source.n43 7.3702
R100 source.n32 source.n31 7.3702
R101 source.n4 source.n3 7.3702
R102 source.n16 source.n15 7.3702
R103 source.n44 source.n40 5.81868
R104 source.n32 source.n28 5.81868
R105 source.n4 source.n0 5.81868
R106 source.n16 source.n12 5.81868
R107 source.n48 source.n47 5.49188
R108 source.n45 source.n41 3.44771
R109 source.n33 source.n29 3.44771
R110 source.n5 source.n1 3.44771
R111 source.n17 source.n13 3.44771
R112 source.n19 source.n11 0.698776
R113 source.n37 source.n35 0.698776
R114 source.n23 source.n21 0.457397
R115 source.n21 source.n19 0.457397
R116 source.n11 source.n9 0.457397
R117 source.n9 source.n7 0.457397
R118 source.n27 source.n25 0.457397
R119 source.n35 source.n27 0.457397
R120 source.n39 source.n37 0.457397
R121 source.n47 source.n39 0.457397
R122 source source.n48 0.188
R123 drain_right.n2 drain_right.n0 289.615
R124 drain_right.n16 drain_right.n14 289.615
R125 drain_right.n3 drain_right.n2 185
R126 drain_right.n17 drain_right.n16 185
R127 drain_right.t0 drain_right.n1 167.117
R128 drain_right.t3 drain_right.n15 167.117
R129 drain_right.n13 drain_right.n11 101.252
R130 drain_right.n10 drain_right.n9 101.082
R131 drain_right.n13 drain_right.n12 100.796
R132 drain_right.n8 drain_right.n7 100.796
R133 drain_right.n2 drain_right.t0 52.3082
R134 drain_right.n16 drain_right.t3 52.3082
R135 drain_right.n8 drain_right.n6 48.5453
R136 drain_right.n21 drain_right.n20 48.0884
R137 drain_right drain_right.n10 21.1799
R138 drain_right.n9 drain_right.t2 9.9005
R139 drain_right.n9 drain_right.t9 9.9005
R140 drain_right.n7 drain_right.t8 9.9005
R141 drain_right.n7 drain_right.t5 9.9005
R142 drain_right.n11 drain_right.t6 9.9005
R143 drain_right.n11 drain_right.t4 9.9005
R144 drain_right.n12 drain_right.t1 9.9005
R145 drain_right.n12 drain_right.t7 9.9005
R146 drain_right.n3 drain_right.n1 9.71174
R147 drain_right.n17 drain_right.n15 9.71174
R148 drain_right.n6 drain_right.n5 9.45567
R149 drain_right.n20 drain_right.n19 9.45567
R150 drain_right.n5 drain_right.n4 9.3005
R151 drain_right.n19 drain_right.n18 9.3005
R152 drain_right.n6 drain_right.n0 8.14595
R153 drain_right.n20 drain_right.n14 8.14595
R154 drain_right.n4 drain_right.n3 7.3702
R155 drain_right.n18 drain_right.n17 7.3702
R156 drain_right drain_right.n21 5.88166
R157 drain_right.n4 drain_right.n0 5.81868
R158 drain_right.n18 drain_right.n14 5.81868
R159 drain_right.n5 drain_right.n1 3.44771
R160 drain_right.n19 drain_right.n15 3.44771
R161 drain_right.n21 drain_right.n13 0.457397
R162 drain_right.n10 drain_right.n8 0.0593781
R163 plus.n2 plus.t4 442.93
R164 plus.n8 plus.t6 442.93
R165 plus.n12 plus.t8 442.93
R166 plus.n18 plus.t3 442.93
R167 plus.n1 plus.t2 397.651
R168 plus.n5 plus.t9 397.651
R169 plus.n7 plus.t7 397.651
R170 plus.n11 plus.t1 397.651
R171 plus.n15 plus.t5 397.651
R172 plus.n17 plus.t0 397.651
R173 plus.n3 plus.n2 161.489
R174 plus.n13 plus.n12 161.489
R175 plus.n4 plus.n3 161.3
R176 plus.n6 plus.n0 161.3
R177 plus.n9 plus.n8 161.3
R178 plus.n14 plus.n13 161.3
R179 plus.n16 plus.n10 161.3
R180 plus.n19 plus.n18 161.3
R181 plus.n4 plus.n1 40.8975
R182 plus.n7 plus.n6 40.8975
R183 plus.n17 plus.n16 40.8975
R184 plus.n14 plus.n11 40.8975
R185 plus.n5 plus.n4 36.5157
R186 plus.n6 plus.n5 36.5157
R187 plus.n16 plus.n15 36.5157
R188 plus.n15 plus.n14 36.5157
R189 plus.n2 plus.n1 32.1338
R190 plus.n8 plus.n7 32.1338
R191 plus.n18 plus.n17 32.1338
R192 plus.n12 plus.n11 32.1338
R193 plus plus.n19 24.285
R194 plus plus.n9 8.30542
R195 plus.n3 plus.n0 0.189894
R196 plus.n9 plus.n0 0.189894
R197 plus.n19 plus.n10 0.189894
R198 plus.n13 plus.n10 0.189894
R199 drain_left.n2 drain_left.n0 289.615
R200 drain_left.n13 drain_left.n11 289.615
R201 drain_left.n3 drain_left.n2 185
R202 drain_left.n14 drain_left.n13 185
R203 drain_left.t6 drain_left.n1 167.117
R204 drain_left.t5 drain_left.n12 167.117
R205 drain_left.n10 drain_left.n9 101.082
R206 drain_left.n21 drain_left.n20 100.796
R207 drain_left.n19 drain_left.n18 100.796
R208 drain_left.n8 drain_left.n7 100.796
R209 drain_left.n2 drain_left.t6 52.3082
R210 drain_left.n13 drain_left.t5 52.3082
R211 drain_left.n8 drain_left.n6 48.5453
R212 drain_left.n19 drain_left.n17 48.5453
R213 drain_left drain_left.n10 21.7331
R214 drain_left.n9 drain_left.t8 9.9005
R215 drain_left.n9 drain_left.t1 9.9005
R216 drain_left.n7 drain_left.t9 9.9005
R217 drain_left.n7 drain_left.t4 9.9005
R218 drain_left.n20 drain_left.t2 9.9005
R219 drain_left.n20 drain_left.t3 9.9005
R220 drain_left.n18 drain_left.t7 9.9005
R221 drain_left.n18 drain_left.t0 9.9005
R222 drain_left.n3 drain_left.n1 9.71174
R223 drain_left.n14 drain_left.n12 9.71174
R224 drain_left.n6 drain_left.n5 9.45567
R225 drain_left.n17 drain_left.n16 9.45567
R226 drain_left.n5 drain_left.n4 9.3005
R227 drain_left.n16 drain_left.n15 9.3005
R228 drain_left.n6 drain_left.n0 8.14595
R229 drain_left.n17 drain_left.n11 8.14595
R230 drain_left.n4 drain_left.n3 7.3702
R231 drain_left.n15 drain_left.n14 7.3702
R232 drain_left drain_left.n21 6.11011
R233 drain_left.n4 drain_left.n0 5.81868
R234 drain_left.n15 drain_left.n11 5.81868
R235 drain_left.n5 drain_left.n1 3.44771
R236 drain_left.n16 drain_left.n12 3.44771
R237 drain_left.n21 drain_left.n19 0.457397
R238 drain_left.n10 drain_left.n8 0.0593781
C0 drain_right minus 0.830732f
C1 source drain_left 5.88398f
C2 plus drain_right 0.28857f
C3 minus drain_left 0.17691f
C4 minus source 0.892382f
C5 plus drain_left 0.958152f
C6 plus source 0.906462f
C7 drain_right drain_left 0.658684f
C8 drain_right source 5.88024f
C9 plus minus 2.99637f
C10 drain_right a_n1352_n1288# 3.52233f
C11 drain_left a_n1352_n1288# 3.7062f
C12 source a_n1352_n1288# 2.374134f
C13 minus a_n1352_n1288# 4.420642f
C14 plus a_n1352_n1288# 5.14544f
C15 drain_left.n0 a_n1352_n1288# 0.038611f
C16 drain_left.n1 a_n1352_n1288# 0.085431f
C17 drain_left.t6 a_n1352_n1288# 0.064112f
C18 drain_left.n2 a_n1352_n1288# 0.066862f
C19 drain_left.n3 a_n1352_n1288# 0.021554f
C20 drain_left.n4 a_n1352_n1288# 0.014215f
C21 drain_left.n5 a_n1352_n1288# 0.188311f
C22 drain_left.n6 a_n1352_n1288# 0.061442f
C23 drain_left.t9 a_n1352_n1288# 0.041809f
C24 drain_left.t4 a_n1352_n1288# 0.041809f
C25 drain_left.n7 a_n1352_n1288# 0.262657f
C26 drain_left.n8 a_n1352_n1288# 0.345074f
C27 drain_left.t8 a_n1352_n1288# 0.041809f
C28 drain_left.t1 a_n1352_n1288# 0.041809f
C29 drain_left.n9 a_n1352_n1288# 0.263449f
C30 drain_left.n10 a_n1352_n1288# 0.892273f
C31 drain_left.n11 a_n1352_n1288# 0.038611f
C32 drain_left.n12 a_n1352_n1288# 0.085431f
C33 drain_left.t5 a_n1352_n1288# 0.064112f
C34 drain_left.n13 a_n1352_n1288# 0.066862f
C35 drain_left.n14 a_n1352_n1288# 0.021554f
C36 drain_left.n15 a_n1352_n1288# 0.014215f
C37 drain_left.n16 a_n1352_n1288# 0.188311f
C38 drain_left.n17 a_n1352_n1288# 0.061442f
C39 drain_left.t7 a_n1352_n1288# 0.041809f
C40 drain_left.t0 a_n1352_n1288# 0.041809f
C41 drain_left.n18 a_n1352_n1288# 0.262658f
C42 drain_left.n19 a_n1352_n1288# 0.368584f
C43 drain_left.t2 a_n1352_n1288# 0.041809f
C44 drain_left.t3 a_n1352_n1288# 0.041809f
C45 drain_left.n20 a_n1352_n1288# 0.262658f
C46 drain_left.n21 a_n1352_n1288# 0.496863f
C47 plus.n0 a_n1352_n1288# 0.036435f
C48 plus.t7 a_n1352_n1288# 0.042885f
C49 plus.t9 a_n1352_n1288# 0.042885f
C50 plus.t2 a_n1352_n1288# 0.042885f
C51 plus.n1 a_n1352_n1288# 0.033696f
C52 plus.t4 a_n1352_n1288# 0.046353f
C53 plus.n2 a_n1352_n1288# 0.043265f
C54 plus.n3 a_n1352_n1288# 0.080007f
C55 plus.n4 a_n1352_n1288# 0.012761f
C56 plus.n5 a_n1352_n1288# 0.033696f
C57 plus.n6 a_n1352_n1288# 0.012761f
C58 plus.n7 a_n1352_n1288# 0.033696f
C59 plus.t6 a_n1352_n1288# 0.046353f
C60 plus.n8 a_n1352_n1288# 0.043213f
C61 plus.n9 a_n1352_n1288# 0.255881f
C62 plus.n10 a_n1352_n1288# 0.036435f
C63 plus.t3 a_n1352_n1288# 0.046353f
C64 plus.t0 a_n1352_n1288# 0.042885f
C65 plus.t5 a_n1352_n1288# 0.042885f
C66 plus.t1 a_n1352_n1288# 0.042885f
C67 plus.n11 a_n1352_n1288# 0.033696f
C68 plus.t8 a_n1352_n1288# 0.046353f
C69 plus.n12 a_n1352_n1288# 0.043265f
C70 plus.n13 a_n1352_n1288# 0.080007f
C71 plus.n14 a_n1352_n1288# 0.012761f
C72 plus.n15 a_n1352_n1288# 0.033696f
C73 plus.n16 a_n1352_n1288# 0.012761f
C74 plus.n17 a_n1352_n1288# 0.033696f
C75 plus.n18 a_n1352_n1288# 0.043213f
C76 plus.n19 a_n1352_n1288# 0.73509f
C77 drain_right.n0 a_n1352_n1288# 0.0393f
C78 drain_right.n1 a_n1352_n1288# 0.086956f
C79 drain_right.t0 a_n1352_n1288# 0.065256f
C80 drain_right.n2 a_n1352_n1288# 0.068055f
C81 drain_right.n3 a_n1352_n1288# 0.021939f
C82 drain_right.n4 a_n1352_n1288# 0.014469f
C83 drain_right.n5 a_n1352_n1288# 0.191673f
C84 drain_right.n6 a_n1352_n1288# 0.062539f
C85 drain_right.t8 a_n1352_n1288# 0.042555f
C86 drain_right.t5 a_n1352_n1288# 0.042555f
C87 drain_right.n7 a_n1352_n1288# 0.267346f
C88 drain_right.n8 a_n1352_n1288# 0.351234f
C89 drain_right.t2 a_n1352_n1288# 0.042555f
C90 drain_right.t9 a_n1352_n1288# 0.042555f
C91 drain_right.n9 a_n1352_n1288# 0.268153f
C92 drain_right.n10 a_n1352_n1288# 0.855192f
C93 drain_right.t6 a_n1352_n1288# 0.042555f
C94 drain_right.t4 a_n1352_n1288# 0.042555f
C95 drain_right.n11 a_n1352_n1288# 0.268684f
C96 drain_right.t1 a_n1352_n1288# 0.042555f
C97 drain_right.t7 a_n1352_n1288# 0.042555f
C98 drain_right.n12 a_n1352_n1288# 0.267348f
C99 drain_right.n13 a_n1352_n1288# 0.580249f
C100 drain_right.n14 a_n1352_n1288# 0.0393f
C101 drain_right.n15 a_n1352_n1288# 0.086956f
C102 drain_right.t3 a_n1352_n1288# 0.065256f
C103 drain_right.n16 a_n1352_n1288# 0.068055f
C104 drain_right.n17 a_n1352_n1288# 0.021939f
C105 drain_right.n18 a_n1352_n1288# 0.014469f
C106 drain_right.n19 a_n1352_n1288# 0.191673f
C107 drain_right.n20 a_n1352_n1288# 0.061686f
C108 drain_right.n21 a_n1352_n1288# 0.309495f
C109 source.n0 a_n1352_n1288# 0.047657f
C110 source.n1 a_n1352_n1288# 0.105448f
C111 source.t6 a_n1352_n1288# 0.079133f
C112 source.n2 a_n1352_n1288# 0.082528f
C113 source.n3 a_n1352_n1288# 0.026604f
C114 source.n4 a_n1352_n1288# 0.017546f
C115 source.n5 a_n1352_n1288# 0.232433f
C116 source.n6 a_n1352_n1288# 0.052244f
C117 source.n7 a_n1352_n1288# 0.476859f
C118 source.t7 a_n1352_n1288# 0.051605f
C119 source.t0 a_n1352_n1288# 0.051605f
C120 source.n8 a_n1352_n1288# 0.275879f
C121 source.n9 a_n1352_n1288# 0.349995f
C122 source.t3 a_n1352_n1288# 0.051605f
C123 source.t9 a_n1352_n1288# 0.051605f
C124 source.n10 a_n1352_n1288# 0.275879f
C125 source.n11 a_n1352_n1288# 0.37539f
C126 source.n12 a_n1352_n1288# 0.047657f
C127 source.n13 a_n1352_n1288# 0.105448f
C128 source.t19 a_n1352_n1288# 0.079133f
C129 source.n14 a_n1352_n1288# 0.082528f
C130 source.n15 a_n1352_n1288# 0.026604f
C131 source.n16 a_n1352_n1288# 0.017546f
C132 source.n17 a_n1352_n1288# 0.232433f
C133 source.n18 a_n1352_n1288# 0.052244f
C134 source.n19 a_n1352_n1288# 0.148418f
C135 source.t14 a_n1352_n1288# 0.051605f
C136 source.t15 a_n1352_n1288# 0.051605f
C137 source.n20 a_n1352_n1288# 0.275879f
C138 source.n21 a_n1352_n1288# 0.349995f
C139 source.t16 a_n1352_n1288# 0.051605f
C140 source.t11 a_n1352_n1288# 0.051605f
C141 source.n22 a_n1352_n1288# 0.275879f
C142 source.n23 a_n1352_n1288# 1.05431f
C143 source.t8 a_n1352_n1288# 0.051605f
C144 source.t5 a_n1352_n1288# 0.051605f
C145 source.n24 a_n1352_n1288# 0.275877f
C146 source.n25 a_n1352_n1288# 1.05431f
C147 source.t4 a_n1352_n1288# 0.051605f
C148 source.t2 a_n1352_n1288# 0.051605f
C149 source.n26 a_n1352_n1288# 0.275877f
C150 source.n27 a_n1352_n1288# 0.349996f
C151 source.n28 a_n1352_n1288# 0.047657f
C152 source.n29 a_n1352_n1288# 0.105448f
C153 source.t1 a_n1352_n1288# 0.079133f
C154 source.n30 a_n1352_n1288# 0.082528f
C155 source.n31 a_n1352_n1288# 0.026604f
C156 source.n32 a_n1352_n1288# 0.017546f
C157 source.n33 a_n1352_n1288# 0.232433f
C158 source.n34 a_n1352_n1288# 0.052244f
C159 source.n35 a_n1352_n1288# 0.148418f
C160 source.t12 a_n1352_n1288# 0.051605f
C161 source.t13 a_n1352_n1288# 0.051605f
C162 source.n36 a_n1352_n1288# 0.275877f
C163 source.n37 a_n1352_n1288# 0.375392f
C164 source.t17 a_n1352_n1288# 0.051605f
C165 source.t10 a_n1352_n1288# 0.051605f
C166 source.n38 a_n1352_n1288# 0.275877f
C167 source.n39 a_n1352_n1288# 0.349996f
C168 source.n40 a_n1352_n1288# 0.047657f
C169 source.n41 a_n1352_n1288# 0.105448f
C170 source.t18 a_n1352_n1288# 0.079133f
C171 source.n42 a_n1352_n1288# 0.082528f
C172 source.n43 a_n1352_n1288# 0.026604f
C173 source.n44 a_n1352_n1288# 0.017546f
C174 source.n45 a_n1352_n1288# 0.232433f
C175 source.n46 a_n1352_n1288# 0.052244f
C176 source.n47 a_n1352_n1288# 0.301431f
C177 source.n48 a_n1352_n1288# 0.803463f
C178 minus.n0 a_n1352_n1288# 0.035562f
C179 minus.t6 a_n1352_n1288# 0.045242f
C180 minus.t8 a_n1352_n1288# 0.041857f
C181 minus.t2 a_n1352_n1288# 0.041857f
C182 minus.t3 a_n1352_n1288# 0.041857f
C183 minus.n1 a_n1352_n1288# 0.032888f
C184 minus.t5 a_n1352_n1288# 0.045242f
C185 minus.n2 a_n1352_n1288# 0.042227f
C186 minus.n3 a_n1352_n1288# 0.078089f
C187 minus.n4 a_n1352_n1288# 0.012455f
C188 minus.n5 a_n1352_n1288# 0.032888f
C189 minus.n6 a_n1352_n1288# 0.012455f
C190 minus.n7 a_n1352_n1288# 0.032888f
C191 minus.n8 a_n1352_n1288# 0.042178f
C192 minus.n9 a_n1352_n1288# 0.747282f
C193 minus.n10 a_n1352_n1288# 0.035562f
C194 minus.t7 a_n1352_n1288# 0.041857f
C195 minus.t4 a_n1352_n1288# 0.041857f
C196 minus.t1 a_n1352_n1288# 0.041857f
C197 minus.n11 a_n1352_n1288# 0.032888f
C198 minus.t9 a_n1352_n1288# 0.045242f
C199 minus.n12 a_n1352_n1288# 0.042227f
C200 minus.n13 a_n1352_n1288# 0.078089f
C201 minus.n14 a_n1352_n1288# 0.012455f
C202 minus.n15 a_n1352_n1288# 0.032888f
C203 minus.n16 a_n1352_n1288# 0.012455f
C204 minus.n17 a_n1352_n1288# 0.032888f
C205 minus.t0 a_n1352_n1288# 0.045242f
C206 minus.n18 a_n1352_n1288# 0.042178f
C207 minus.n19 a_n1352_n1288# 0.22824f
C208 minus.n20 a_n1352_n1288# 0.925757f
.ends

