* NGSPICE file created from diffpair281.ext - technology: sky130A

.subckt diffpair281 minus drain_right drain_left source plus
X0 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X1 source.t6 minus.t0 drain_right.t2 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X2 source.t1 plus.t0 drain_left.t3 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X3 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X4 drain_left.t2 plus.t1 source.t0 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X5 source.t7 plus.t2 drain_left.t1 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X6 drain_right.t0 minus.t1 source.t5 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X7 drain_left.t0 plus.t3 source.t2 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X8 drain_right.t3 minus.t2 source.t4 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X9 source.t3 minus.t3 drain_right.t1 a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X10 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X11 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
R0 minus.n0 minus.t1 388.748
R1 minus.n1 minus.t3 388.748
R2 minus.n0 minus.t0 388.724
R3 minus.n1 minus.t2 388.724
R4 minus.n2 minus.n0 99.4525
R5 minus.n2 minus.n1 76.7783
R6 minus minus.n2 0.188
R7 drain_right drain_right.n0 90.8896
R8 drain_right drain_right.n1 73.5589
R9 drain_right.n0 drain_right.t1 3.3005
R10 drain_right.n0 drain_right.t3 3.3005
R11 drain_right.n1 drain_right.t2 3.3005
R12 drain_right.n1 drain_right.t0 3.3005
R13 source.n250 source.n224 289.615
R14 source.n218 source.n192 289.615
R15 source.n186 source.n160 289.615
R16 source.n154 source.n128 289.615
R17 source.n26 source.n0 289.615
R18 source.n58 source.n32 289.615
R19 source.n90 source.n64 289.615
R20 source.n122 source.n96 289.615
R21 source.n235 source.n234 185
R22 source.n232 source.n231 185
R23 source.n241 source.n240 185
R24 source.n243 source.n242 185
R25 source.n228 source.n227 185
R26 source.n249 source.n248 185
R27 source.n251 source.n250 185
R28 source.n203 source.n202 185
R29 source.n200 source.n199 185
R30 source.n209 source.n208 185
R31 source.n211 source.n210 185
R32 source.n196 source.n195 185
R33 source.n217 source.n216 185
R34 source.n219 source.n218 185
R35 source.n171 source.n170 185
R36 source.n168 source.n167 185
R37 source.n177 source.n176 185
R38 source.n179 source.n178 185
R39 source.n164 source.n163 185
R40 source.n185 source.n184 185
R41 source.n187 source.n186 185
R42 source.n139 source.n138 185
R43 source.n136 source.n135 185
R44 source.n145 source.n144 185
R45 source.n147 source.n146 185
R46 source.n132 source.n131 185
R47 source.n153 source.n152 185
R48 source.n155 source.n154 185
R49 source.n27 source.n26 185
R50 source.n25 source.n24 185
R51 source.n4 source.n3 185
R52 source.n19 source.n18 185
R53 source.n17 source.n16 185
R54 source.n8 source.n7 185
R55 source.n11 source.n10 185
R56 source.n59 source.n58 185
R57 source.n57 source.n56 185
R58 source.n36 source.n35 185
R59 source.n51 source.n50 185
R60 source.n49 source.n48 185
R61 source.n40 source.n39 185
R62 source.n43 source.n42 185
R63 source.n91 source.n90 185
R64 source.n89 source.n88 185
R65 source.n68 source.n67 185
R66 source.n83 source.n82 185
R67 source.n81 source.n80 185
R68 source.n72 source.n71 185
R69 source.n75 source.n74 185
R70 source.n123 source.n122 185
R71 source.n121 source.n120 185
R72 source.n100 source.n99 185
R73 source.n115 source.n114 185
R74 source.n113 source.n112 185
R75 source.n104 source.n103 185
R76 source.n107 source.n106 185
R77 source.t4 source.n233 147.661
R78 source.t3 source.n201 147.661
R79 source.t0 source.n169 147.661
R80 source.t7 source.n137 147.661
R81 source.t2 source.n9 147.661
R82 source.t1 source.n41 147.661
R83 source.t5 source.n73 147.661
R84 source.t6 source.n105 147.661
R85 source.n234 source.n231 104.615
R86 source.n241 source.n231 104.615
R87 source.n242 source.n241 104.615
R88 source.n242 source.n227 104.615
R89 source.n249 source.n227 104.615
R90 source.n250 source.n249 104.615
R91 source.n202 source.n199 104.615
R92 source.n209 source.n199 104.615
R93 source.n210 source.n209 104.615
R94 source.n210 source.n195 104.615
R95 source.n217 source.n195 104.615
R96 source.n218 source.n217 104.615
R97 source.n170 source.n167 104.615
R98 source.n177 source.n167 104.615
R99 source.n178 source.n177 104.615
R100 source.n178 source.n163 104.615
R101 source.n185 source.n163 104.615
R102 source.n186 source.n185 104.615
R103 source.n138 source.n135 104.615
R104 source.n145 source.n135 104.615
R105 source.n146 source.n145 104.615
R106 source.n146 source.n131 104.615
R107 source.n153 source.n131 104.615
R108 source.n154 source.n153 104.615
R109 source.n26 source.n25 104.615
R110 source.n25 source.n3 104.615
R111 source.n18 source.n3 104.615
R112 source.n18 source.n17 104.615
R113 source.n17 source.n7 104.615
R114 source.n10 source.n7 104.615
R115 source.n58 source.n57 104.615
R116 source.n57 source.n35 104.615
R117 source.n50 source.n35 104.615
R118 source.n50 source.n49 104.615
R119 source.n49 source.n39 104.615
R120 source.n42 source.n39 104.615
R121 source.n90 source.n89 104.615
R122 source.n89 source.n67 104.615
R123 source.n82 source.n67 104.615
R124 source.n82 source.n81 104.615
R125 source.n81 source.n71 104.615
R126 source.n74 source.n71 104.615
R127 source.n122 source.n121 104.615
R128 source.n121 source.n99 104.615
R129 source.n114 source.n99 104.615
R130 source.n114 source.n113 104.615
R131 source.n113 source.n103 104.615
R132 source.n106 source.n103 104.615
R133 source.n234 source.t4 52.3082
R134 source.n202 source.t3 52.3082
R135 source.n170 source.t0 52.3082
R136 source.n138 source.t7 52.3082
R137 source.n10 source.t2 52.3082
R138 source.n42 source.t1 52.3082
R139 source.n74 source.t5 52.3082
R140 source.n106 source.t6 52.3082
R141 source.n255 source.n254 32.1853
R142 source.n223 source.n222 32.1853
R143 source.n191 source.n190 32.1853
R144 source.n159 source.n158 32.1853
R145 source.n31 source.n30 32.1853
R146 source.n63 source.n62 32.1853
R147 source.n95 source.n94 32.1853
R148 source.n127 source.n126 32.1853
R149 source.n159 source.n127 17.4578
R150 source.n235 source.n233 15.6674
R151 source.n203 source.n201 15.6674
R152 source.n171 source.n169 15.6674
R153 source.n139 source.n137 15.6674
R154 source.n11 source.n9 15.6674
R155 source.n43 source.n41 15.6674
R156 source.n75 source.n73 15.6674
R157 source.n107 source.n105 15.6674
R158 source.n236 source.n232 12.8005
R159 source.n204 source.n200 12.8005
R160 source.n172 source.n168 12.8005
R161 source.n140 source.n136 12.8005
R162 source.n12 source.n8 12.8005
R163 source.n44 source.n40 12.8005
R164 source.n76 source.n72 12.8005
R165 source.n108 source.n104 12.8005
R166 source.n240 source.n239 12.0247
R167 source.n208 source.n207 12.0247
R168 source.n176 source.n175 12.0247
R169 source.n144 source.n143 12.0247
R170 source.n16 source.n15 12.0247
R171 source.n48 source.n47 12.0247
R172 source.n80 source.n79 12.0247
R173 source.n112 source.n111 12.0247
R174 source.n256 source.n31 11.8371
R175 source.n243 source.n230 11.249
R176 source.n211 source.n198 11.249
R177 source.n179 source.n166 11.249
R178 source.n147 source.n134 11.249
R179 source.n19 source.n6 11.249
R180 source.n51 source.n38 11.249
R181 source.n83 source.n70 11.249
R182 source.n115 source.n102 11.249
R183 source.n244 source.n228 10.4732
R184 source.n212 source.n196 10.4732
R185 source.n180 source.n164 10.4732
R186 source.n148 source.n132 10.4732
R187 source.n20 source.n4 10.4732
R188 source.n52 source.n36 10.4732
R189 source.n84 source.n68 10.4732
R190 source.n116 source.n100 10.4732
R191 source.n248 source.n247 9.69747
R192 source.n216 source.n215 9.69747
R193 source.n184 source.n183 9.69747
R194 source.n152 source.n151 9.69747
R195 source.n24 source.n23 9.69747
R196 source.n56 source.n55 9.69747
R197 source.n88 source.n87 9.69747
R198 source.n120 source.n119 9.69747
R199 source.n254 source.n253 9.45567
R200 source.n222 source.n221 9.45567
R201 source.n190 source.n189 9.45567
R202 source.n158 source.n157 9.45567
R203 source.n30 source.n29 9.45567
R204 source.n62 source.n61 9.45567
R205 source.n94 source.n93 9.45567
R206 source.n126 source.n125 9.45567
R207 source.n253 source.n252 9.3005
R208 source.n226 source.n225 9.3005
R209 source.n247 source.n246 9.3005
R210 source.n245 source.n244 9.3005
R211 source.n230 source.n229 9.3005
R212 source.n239 source.n238 9.3005
R213 source.n237 source.n236 9.3005
R214 source.n221 source.n220 9.3005
R215 source.n194 source.n193 9.3005
R216 source.n215 source.n214 9.3005
R217 source.n213 source.n212 9.3005
R218 source.n198 source.n197 9.3005
R219 source.n207 source.n206 9.3005
R220 source.n205 source.n204 9.3005
R221 source.n189 source.n188 9.3005
R222 source.n162 source.n161 9.3005
R223 source.n183 source.n182 9.3005
R224 source.n181 source.n180 9.3005
R225 source.n166 source.n165 9.3005
R226 source.n175 source.n174 9.3005
R227 source.n173 source.n172 9.3005
R228 source.n157 source.n156 9.3005
R229 source.n130 source.n129 9.3005
R230 source.n151 source.n150 9.3005
R231 source.n149 source.n148 9.3005
R232 source.n134 source.n133 9.3005
R233 source.n143 source.n142 9.3005
R234 source.n141 source.n140 9.3005
R235 source.n29 source.n28 9.3005
R236 source.n2 source.n1 9.3005
R237 source.n23 source.n22 9.3005
R238 source.n21 source.n20 9.3005
R239 source.n6 source.n5 9.3005
R240 source.n15 source.n14 9.3005
R241 source.n13 source.n12 9.3005
R242 source.n61 source.n60 9.3005
R243 source.n34 source.n33 9.3005
R244 source.n55 source.n54 9.3005
R245 source.n53 source.n52 9.3005
R246 source.n38 source.n37 9.3005
R247 source.n47 source.n46 9.3005
R248 source.n45 source.n44 9.3005
R249 source.n93 source.n92 9.3005
R250 source.n66 source.n65 9.3005
R251 source.n87 source.n86 9.3005
R252 source.n85 source.n84 9.3005
R253 source.n70 source.n69 9.3005
R254 source.n79 source.n78 9.3005
R255 source.n77 source.n76 9.3005
R256 source.n125 source.n124 9.3005
R257 source.n98 source.n97 9.3005
R258 source.n119 source.n118 9.3005
R259 source.n117 source.n116 9.3005
R260 source.n102 source.n101 9.3005
R261 source.n111 source.n110 9.3005
R262 source.n109 source.n108 9.3005
R263 source.n251 source.n226 8.92171
R264 source.n219 source.n194 8.92171
R265 source.n187 source.n162 8.92171
R266 source.n155 source.n130 8.92171
R267 source.n27 source.n2 8.92171
R268 source.n59 source.n34 8.92171
R269 source.n91 source.n66 8.92171
R270 source.n123 source.n98 8.92171
R271 source.n252 source.n224 8.14595
R272 source.n220 source.n192 8.14595
R273 source.n188 source.n160 8.14595
R274 source.n156 source.n128 8.14595
R275 source.n28 source.n0 8.14595
R276 source.n60 source.n32 8.14595
R277 source.n92 source.n64 8.14595
R278 source.n124 source.n96 8.14595
R279 source.n254 source.n224 5.81868
R280 source.n222 source.n192 5.81868
R281 source.n190 source.n160 5.81868
R282 source.n158 source.n128 5.81868
R283 source.n30 source.n0 5.81868
R284 source.n62 source.n32 5.81868
R285 source.n94 source.n64 5.81868
R286 source.n126 source.n96 5.81868
R287 source.n256 source.n255 5.62119
R288 source.n252 source.n251 5.04292
R289 source.n220 source.n219 5.04292
R290 source.n188 source.n187 5.04292
R291 source.n156 source.n155 5.04292
R292 source.n28 source.n27 5.04292
R293 source.n60 source.n59 5.04292
R294 source.n92 source.n91 5.04292
R295 source.n124 source.n123 5.04292
R296 source.n237 source.n233 4.38594
R297 source.n205 source.n201 4.38594
R298 source.n173 source.n169 4.38594
R299 source.n141 source.n137 4.38594
R300 source.n13 source.n9 4.38594
R301 source.n45 source.n41 4.38594
R302 source.n77 source.n73 4.38594
R303 source.n109 source.n105 4.38594
R304 source.n248 source.n226 4.26717
R305 source.n216 source.n194 4.26717
R306 source.n184 source.n162 4.26717
R307 source.n152 source.n130 4.26717
R308 source.n24 source.n2 4.26717
R309 source.n56 source.n34 4.26717
R310 source.n88 source.n66 4.26717
R311 source.n120 source.n98 4.26717
R312 source.n247 source.n228 3.49141
R313 source.n215 source.n196 3.49141
R314 source.n183 source.n164 3.49141
R315 source.n151 source.n132 3.49141
R316 source.n23 source.n4 3.49141
R317 source.n55 source.n36 3.49141
R318 source.n87 source.n68 3.49141
R319 source.n119 source.n100 3.49141
R320 source.n244 source.n243 2.71565
R321 source.n212 source.n211 2.71565
R322 source.n180 source.n179 2.71565
R323 source.n148 source.n147 2.71565
R324 source.n20 source.n19 2.71565
R325 source.n52 source.n51 2.71565
R326 source.n84 source.n83 2.71565
R327 source.n116 source.n115 2.71565
R328 source.n240 source.n230 1.93989
R329 source.n208 source.n198 1.93989
R330 source.n176 source.n166 1.93989
R331 source.n144 source.n134 1.93989
R332 source.n16 source.n6 1.93989
R333 source.n48 source.n38 1.93989
R334 source.n80 source.n70 1.93989
R335 source.n112 source.n102 1.93989
R336 source.n239 source.n232 1.16414
R337 source.n207 source.n200 1.16414
R338 source.n175 source.n168 1.16414
R339 source.n143 source.n136 1.16414
R340 source.n15 source.n8 1.16414
R341 source.n47 source.n40 1.16414
R342 source.n79 source.n72 1.16414
R343 source.n111 source.n104 1.16414
R344 source.n127 source.n95 0.716017
R345 source.n63 source.n31 0.716017
R346 source.n191 source.n159 0.716017
R347 source.n255 source.n223 0.716017
R348 source.n95 source.n63 0.470328
R349 source.n223 source.n191 0.470328
R350 source.n236 source.n235 0.388379
R351 source.n204 source.n203 0.388379
R352 source.n172 source.n171 0.388379
R353 source.n140 source.n139 0.388379
R354 source.n12 source.n11 0.388379
R355 source.n44 source.n43 0.388379
R356 source.n76 source.n75 0.388379
R357 source.n108 source.n107 0.388379
R358 source source.n256 0.188
R359 source.n238 source.n237 0.155672
R360 source.n238 source.n229 0.155672
R361 source.n245 source.n229 0.155672
R362 source.n246 source.n245 0.155672
R363 source.n246 source.n225 0.155672
R364 source.n253 source.n225 0.155672
R365 source.n206 source.n205 0.155672
R366 source.n206 source.n197 0.155672
R367 source.n213 source.n197 0.155672
R368 source.n214 source.n213 0.155672
R369 source.n214 source.n193 0.155672
R370 source.n221 source.n193 0.155672
R371 source.n174 source.n173 0.155672
R372 source.n174 source.n165 0.155672
R373 source.n181 source.n165 0.155672
R374 source.n182 source.n181 0.155672
R375 source.n182 source.n161 0.155672
R376 source.n189 source.n161 0.155672
R377 source.n142 source.n141 0.155672
R378 source.n142 source.n133 0.155672
R379 source.n149 source.n133 0.155672
R380 source.n150 source.n149 0.155672
R381 source.n150 source.n129 0.155672
R382 source.n157 source.n129 0.155672
R383 source.n29 source.n1 0.155672
R384 source.n22 source.n1 0.155672
R385 source.n22 source.n21 0.155672
R386 source.n21 source.n5 0.155672
R387 source.n14 source.n5 0.155672
R388 source.n14 source.n13 0.155672
R389 source.n61 source.n33 0.155672
R390 source.n54 source.n33 0.155672
R391 source.n54 source.n53 0.155672
R392 source.n53 source.n37 0.155672
R393 source.n46 source.n37 0.155672
R394 source.n46 source.n45 0.155672
R395 source.n93 source.n65 0.155672
R396 source.n86 source.n65 0.155672
R397 source.n86 source.n85 0.155672
R398 source.n85 source.n69 0.155672
R399 source.n78 source.n69 0.155672
R400 source.n78 source.n77 0.155672
R401 source.n125 source.n97 0.155672
R402 source.n118 source.n97 0.155672
R403 source.n118 source.n117 0.155672
R404 source.n117 source.n101 0.155672
R405 source.n110 source.n101 0.155672
R406 source.n110 source.n109 0.155672
R407 plus.n0 plus.t0 388.748
R408 plus.n1 plus.t1 388.748
R409 plus.n0 plus.t3 388.724
R410 plus.n1 plus.t2 388.724
R411 plus plus.n1 95.6064
R412 plus plus.n0 80.1495
R413 drain_left drain_left.n0 91.4428
R414 drain_left drain_left.n1 73.5589
R415 drain_left.n0 drain_left.t1 3.3005
R416 drain_left.n0 drain_left.t2 3.3005
R417 drain_left.n1 drain_left.t3 3.3005
R418 drain_left.n1 drain_left.t0 3.3005
C0 drain_right minus 1.49211f
C1 source minus 1.33827f
C2 drain_left plus 1.60556f
C3 drain_right drain_left 0.522435f
C4 source drain_left 4.63548f
C5 drain_right plus 0.266739f
C6 source plus 1.35229f
C7 drain_left minus 0.170454f
C8 plus minus 3.54726f
C9 drain_right source 4.63523f
C10 drain_right a_n1214_n2088# 4.34672f
C11 drain_left a_n1214_n2088# 4.49327f
C12 source a_n1214_n2088# 5.186623f
C13 minus a_n1214_n2088# 4.108154f
C14 plus a_n1214_n2088# 5.664f
C15 drain_left.t1 a_n1214_n2088# 0.099391f
C16 drain_left.t2 a_n1214_n2088# 0.099391f
C17 drain_left.n0 a_n1214_n2088# 1.01002f
C18 drain_left.t3 a_n1214_n2088# 0.099391f
C19 drain_left.t0 a_n1214_n2088# 0.099391f
C20 drain_left.n1 a_n1214_n2088# 0.868347f
C21 plus.t3 a_n1214_n2088# 0.272451f
C22 plus.t0 a_n1214_n2088# 0.272461f
C23 plus.n0 a_n1214_n2088# 0.274449f
C24 plus.t2 a_n1214_n2088# 0.272451f
C25 plus.t1 a_n1214_n2088# 0.272461f
C26 plus.n1 a_n1214_n2088# 0.429854f
C27 source.n0 a_n1214_n2088# 0.020176f
C28 source.n1 a_n1214_n2088# 0.014354f
C29 source.n2 a_n1214_n2088# 0.007713f
C30 source.n3 a_n1214_n2088# 0.018231f
C31 source.n4 a_n1214_n2088# 0.008167f
C32 source.n5 a_n1214_n2088# 0.014354f
C33 source.n6 a_n1214_n2088# 0.007713f
C34 source.n7 a_n1214_n2088# 0.018231f
C35 source.n8 a_n1214_n2088# 0.008167f
C36 source.n9 a_n1214_n2088# 0.061425f
C37 source.t2 a_n1214_n2088# 0.029715f
C38 source.n10 a_n1214_n2088# 0.013674f
C39 source.n11 a_n1214_n2088# 0.010769f
C40 source.n12 a_n1214_n2088# 0.007713f
C41 source.n13 a_n1214_n2088# 0.34154f
C42 source.n14 a_n1214_n2088# 0.014354f
C43 source.n15 a_n1214_n2088# 0.007713f
C44 source.n16 a_n1214_n2088# 0.008167f
C45 source.n17 a_n1214_n2088# 0.018231f
C46 source.n18 a_n1214_n2088# 0.018231f
C47 source.n19 a_n1214_n2088# 0.008167f
C48 source.n20 a_n1214_n2088# 0.007713f
C49 source.n21 a_n1214_n2088# 0.014354f
C50 source.n22 a_n1214_n2088# 0.014354f
C51 source.n23 a_n1214_n2088# 0.007713f
C52 source.n24 a_n1214_n2088# 0.008167f
C53 source.n25 a_n1214_n2088# 0.018231f
C54 source.n26 a_n1214_n2088# 0.039468f
C55 source.n27 a_n1214_n2088# 0.008167f
C56 source.n28 a_n1214_n2088# 0.007713f
C57 source.n29 a_n1214_n2088# 0.033179f
C58 source.n30 a_n1214_n2088# 0.022084f
C59 source.n31 a_n1214_n2088# 0.361343f
C60 source.n32 a_n1214_n2088# 0.020176f
C61 source.n33 a_n1214_n2088# 0.014354f
C62 source.n34 a_n1214_n2088# 0.007713f
C63 source.n35 a_n1214_n2088# 0.018231f
C64 source.n36 a_n1214_n2088# 0.008167f
C65 source.n37 a_n1214_n2088# 0.014354f
C66 source.n38 a_n1214_n2088# 0.007713f
C67 source.n39 a_n1214_n2088# 0.018231f
C68 source.n40 a_n1214_n2088# 0.008167f
C69 source.n41 a_n1214_n2088# 0.061425f
C70 source.t1 a_n1214_n2088# 0.029715f
C71 source.n42 a_n1214_n2088# 0.013674f
C72 source.n43 a_n1214_n2088# 0.010769f
C73 source.n44 a_n1214_n2088# 0.007713f
C74 source.n45 a_n1214_n2088# 0.34154f
C75 source.n46 a_n1214_n2088# 0.014354f
C76 source.n47 a_n1214_n2088# 0.007713f
C77 source.n48 a_n1214_n2088# 0.008167f
C78 source.n49 a_n1214_n2088# 0.018231f
C79 source.n50 a_n1214_n2088# 0.018231f
C80 source.n51 a_n1214_n2088# 0.008167f
C81 source.n52 a_n1214_n2088# 0.007713f
C82 source.n53 a_n1214_n2088# 0.014354f
C83 source.n54 a_n1214_n2088# 0.014354f
C84 source.n55 a_n1214_n2088# 0.007713f
C85 source.n56 a_n1214_n2088# 0.008167f
C86 source.n57 a_n1214_n2088# 0.018231f
C87 source.n58 a_n1214_n2088# 0.039468f
C88 source.n59 a_n1214_n2088# 0.008167f
C89 source.n60 a_n1214_n2088# 0.007713f
C90 source.n61 a_n1214_n2088# 0.033179f
C91 source.n62 a_n1214_n2088# 0.022084f
C92 source.n63 a_n1214_n2088# 0.067084f
C93 source.n64 a_n1214_n2088# 0.020176f
C94 source.n65 a_n1214_n2088# 0.014354f
C95 source.n66 a_n1214_n2088# 0.007713f
C96 source.n67 a_n1214_n2088# 0.018231f
C97 source.n68 a_n1214_n2088# 0.008167f
C98 source.n69 a_n1214_n2088# 0.014354f
C99 source.n70 a_n1214_n2088# 0.007713f
C100 source.n71 a_n1214_n2088# 0.018231f
C101 source.n72 a_n1214_n2088# 0.008167f
C102 source.n73 a_n1214_n2088# 0.061425f
C103 source.t5 a_n1214_n2088# 0.029715f
C104 source.n74 a_n1214_n2088# 0.013674f
C105 source.n75 a_n1214_n2088# 0.010769f
C106 source.n76 a_n1214_n2088# 0.007713f
C107 source.n77 a_n1214_n2088# 0.34154f
C108 source.n78 a_n1214_n2088# 0.014354f
C109 source.n79 a_n1214_n2088# 0.007713f
C110 source.n80 a_n1214_n2088# 0.008167f
C111 source.n81 a_n1214_n2088# 0.018231f
C112 source.n82 a_n1214_n2088# 0.018231f
C113 source.n83 a_n1214_n2088# 0.008167f
C114 source.n84 a_n1214_n2088# 0.007713f
C115 source.n85 a_n1214_n2088# 0.014354f
C116 source.n86 a_n1214_n2088# 0.014354f
C117 source.n87 a_n1214_n2088# 0.007713f
C118 source.n88 a_n1214_n2088# 0.008167f
C119 source.n89 a_n1214_n2088# 0.018231f
C120 source.n90 a_n1214_n2088# 0.039468f
C121 source.n91 a_n1214_n2088# 0.008167f
C122 source.n92 a_n1214_n2088# 0.007713f
C123 source.n93 a_n1214_n2088# 0.033179f
C124 source.n94 a_n1214_n2088# 0.022084f
C125 source.n95 a_n1214_n2088# 0.067084f
C126 source.n96 a_n1214_n2088# 0.020176f
C127 source.n97 a_n1214_n2088# 0.014354f
C128 source.n98 a_n1214_n2088# 0.007713f
C129 source.n99 a_n1214_n2088# 0.018231f
C130 source.n100 a_n1214_n2088# 0.008167f
C131 source.n101 a_n1214_n2088# 0.014354f
C132 source.n102 a_n1214_n2088# 0.007713f
C133 source.n103 a_n1214_n2088# 0.018231f
C134 source.n104 a_n1214_n2088# 0.008167f
C135 source.n105 a_n1214_n2088# 0.061425f
C136 source.t6 a_n1214_n2088# 0.029715f
C137 source.n106 a_n1214_n2088# 0.013674f
C138 source.n107 a_n1214_n2088# 0.010769f
C139 source.n108 a_n1214_n2088# 0.007713f
C140 source.n109 a_n1214_n2088# 0.34154f
C141 source.n110 a_n1214_n2088# 0.014354f
C142 source.n111 a_n1214_n2088# 0.007713f
C143 source.n112 a_n1214_n2088# 0.008167f
C144 source.n113 a_n1214_n2088# 0.018231f
C145 source.n114 a_n1214_n2088# 0.018231f
C146 source.n115 a_n1214_n2088# 0.008167f
C147 source.n116 a_n1214_n2088# 0.007713f
C148 source.n117 a_n1214_n2088# 0.014354f
C149 source.n118 a_n1214_n2088# 0.014354f
C150 source.n119 a_n1214_n2088# 0.007713f
C151 source.n120 a_n1214_n2088# 0.008167f
C152 source.n121 a_n1214_n2088# 0.018231f
C153 source.n122 a_n1214_n2088# 0.039468f
C154 source.n123 a_n1214_n2088# 0.008167f
C155 source.n124 a_n1214_n2088# 0.007713f
C156 source.n125 a_n1214_n2088# 0.033179f
C157 source.n126 a_n1214_n2088# 0.022084f
C158 source.n127 a_n1214_n2088# 0.548425f
C159 source.n128 a_n1214_n2088# 0.020176f
C160 source.n129 a_n1214_n2088# 0.014354f
C161 source.n130 a_n1214_n2088# 0.007713f
C162 source.n131 a_n1214_n2088# 0.018231f
C163 source.n132 a_n1214_n2088# 0.008167f
C164 source.n133 a_n1214_n2088# 0.014354f
C165 source.n134 a_n1214_n2088# 0.007713f
C166 source.n135 a_n1214_n2088# 0.018231f
C167 source.n136 a_n1214_n2088# 0.008167f
C168 source.n137 a_n1214_n2088# 0.061425f
C169 source.t7 a_n1214_n2088# 0.029715f
C170 source.n138 a_n1214_n2088# 0.013674f
C171 source.n139 a_n1214_n2088# 0.010769f
C172 source.n140 a_n1214_n2088# 0.007713f
C173 source.n141 a_n1214_n2088# 0.34154f
C174 source.n142 a_n1214_n2088# 0.014354f
C175 source.n143 a_n1214_n2088# 0.007713f
C176 source.n144 a_n1214_n2088# 0.008167f
C177 source.n145 a_n1214_n2088# 0.018231f
C178 source.n146 a_n1214_n2088# 0.018231f
C179 source.n147 a_n1214_n2088# 0.008167f
C180 source.n148 a_n1214_n2088# 0.007713f
C181 source.n149 a_n1214_n2088# 0.014354f
C182 source.n150 a_n1214_n2088# 0.014354f
C183 source.n151 a_n1214_n2088# 0.007713f
C184 source.n152 a_n1214_n2088# 0.008167f
C185 source.n153 a_n1214_n2088# 0.018231f
C186 source.n154 a_n1214_n2088# 0.039468f
C187 source.n155 a_n1214_n2088# 0.008167f
C188 source.n156 a_n1214_n2088# 0.007713f
C189 source.n157 a_n1214_n2088# 0.033179f
C190 source.n158 a_n1214_n2088# 0.022084f
C191 source.n159 a_n1214_n2088# 0.548425f
C192 source.n160 a_n1214_n2088# 0.020176f
C193 source.n161 a_n1214_n2088# 0.014354f
C194 source.n162 a_n1214_n2088# 0.007713f
C195 source.n163 a_n1214_n2088# 0.018231f
C196 source.n164 a_n1214_n2088# 0.008167f
C197 source.n165 a_n1214_n2088# 0.014354f
C198 source.n166 a_n1214_n2088# 0.007713f
C199 source.n167 a_n1214_n2088# 0.018231f
C200 source.n168 a_n1214_n2088# 0.008167f
C201 source.n169 a_n1214_n2088# 0.061425f
C202 source.t0 a_n1214_n2088# 0.029715f
C203 source.n170 a_n1214_n2088# 0.013674f
C204 source.n171 a_n1214_n2088# 0.010769f
C205 source.n172 a_n1214_n2088# 0.007713f
C206 source.n173 a_n1214_n2088# 0.34154f
C207 source.n174 a_n1214_n2088# 0.014354f
C208 source.n175 a_n1214_n2088# 0.007713f
C209 source.n176 a_n1214_n2088# 0.008167f
C210 source.n177 a_n1214_n2088# 0.018231f
C211 source.n178 a_n1214_n2088# 0.018231f
C212 source.n179 a_n1214_n2088# 0.008167f
C213 source.n180 a_n1214_n2088# 0.007713f
C214 source.n181 a_n1214_n2088# 0.014354f
C215 source.n182 a_n1214_n2088# 0.014354f
C216 source.n183 a_n1214_n2088# 0.007713f
C217 source.n184 a_n1214_n2088# 0.008167f
C218 source.n185 a_n1214_n2088# 0.018231f
C219 source.n186 a_n1214_n2088# 0.039468f
C220 source.n187 a_n1214_n2088# 0.008167f
C221 source.n188 a_n1214_n2088# 0.007713f
C222 source.n189 a_n1214_n2088# 0.033179f
C223 source.n190 a_n1214_n2088# 0.022084f
C224 source.n191 a_n1214_n2088# 0.067084f
C225 source.n192 a_n1214_n2088# 0.020176f
C226 source.n193 a_n1214_n2088# 0.014354f
C227 source.n194 a_n1214_n2088# 0.007713f
C228 source.n195 a_n1214_n2088# 0.018231f
C229 source.n196 a_n1214_n2088# 0.008167f
C230 source.n197 a_n1214_n2088# 0.014354f
C231 source.n198 a_n1214_n2088# 0.007713f
C232 source.n199 a_n1214_n2088# 0.018231f
C233 source.n200 a_n1214_n2088# 0.008167f
C234 source.n201 a_n1214_n2088# 0.061425f
C235 source.t3 a_n1214_n2088# 0.029715f
C236 source.n202 a_n1214_n2088# 0.013674f
C237 source.n203 a_n1214_n2088# 0.010769f
C238 source.n204 a_n1214_n2088# 0.007713f
C239 source.n205 a_n1214_n2088# 0.34154f
C240 source.n206 a_n1214_n2088# 0.014354f
C241 source.n207 a_n1214_n2088# 0.007713f
C242 source.n208 a_n1214_n2088# 0.008167f
C243 source.n209 a_n1214_n2088# 0.018231f
C244 source.n210 a_n1214_n2088# 0.018231f
C245 source.n211 a_n1214_n2088# 0.008167f
C246 source.n212 a_n1214_n2088# 0.007713f
C247 source.n213 a_n1214_n2088# 0.014354f
C248 source.n214 a_n1214_n2088# 0.014354f
C249 source.n215 a_n1214_n2088# 0.007713f
C250 source.n216 a_n1214_n2088# 0.008167f
C251 source.n217 a_n1214_n2088# 0.018231f
C252 source.n218 a_n1214_n2088# 0.039468f
C253 source.n219 a_n1214_n2088# 0.008167f
C254 source.n220 a_n1214_n2088# 0.007713f
C255 source.n221 a_n1214_n2088# 0.033179f
C256 source.n222 a_n1214_n2088# 0.022084f
C257 source.n223 a_n1214_n2088# 0.067084f
C258 source.n224 a_n1214_n2088# 0.020176f
C259 source.n225 a_n1214_n2088# 0.014354f
C260 source.n226 a_n1214_n2088# 0.007713f
C261 source.n227 a_n1214_n2088# 0.018231f
C262 source.n228 a_n1214_n2088# 0.008167f
C263 source.n229 a_n1214_n2088# 0.014354f
C264 source.n230 a_n1214_n2088# 0.007713f
C265 source.n231 a_n1214_n2088# 0.018231f
C266 source.n232 a_n1214_n2088# 0.008167f
C267 source.n233 a_n1214_n2088# 0.061425f
C268 source.t4 a_n1214_n2088# 0.029715f
C269 source.n234 a_n1214_n2088# 0.013674f
C270 source.n235 a_n1214_n2088# 0.010769f
C271 source.n236 a_n1214_n2088# 0.007713f
C272 source.n237 a_n1214_n2088# 0.34154f
C273 source.n238 a_n1214_n2088# 0.014354f
C274 source.n239 a_n1214_n2088# 0.007713f
C275 source.n240 a_n1214_n2088# 0.008167f
C276 source.n241 a_n1214_n2088# 0.018231f
C277 source.n242 a_n1214_n2088# 0.018231f
C278 source.n243 a_n1214_n2088# 0.008167f
C279 source.n244 a_n1214_n2088# 0.007713f
C280 source.n245 a_n1214_n2088# 0.014354f
C281 source.n246 a_n1214_n2088# 0.014354f
C282 source.n247 a_n1214_n2088# 0.007713f
C283 source.n248 a_n1214_n2088# 0.008167f
C284 source.n249 a_n1214_n2088# 0.018231f
C285 source.n250 a_n1214_n2088# 0.039468f
C286 source.n251 a_n1214_n2088# 0.008167f
C287 source.n252 a_n1214_n2088# 0.007713f
C288 source.n253 a_n1214_n2088# 0.033179f
C289 source.n254 a_n1214_n2088# 0.022084f
C290 source.n255 a_n1214_n2088# 0.154449f
C291 source.n256 a_n1214_n2088# 0.591268f
C292 drain_right.t1 a_n1214_n2088# 0.101196f
C293 drain_right.t3 a_n1214_n2088# 0.101196f
C294 drain_right.n0 a_n1214_n2088# 1.01382f
C295 drain_right.t2 a_n1214_n2088# 0.101196f
C296 drain_right.t0 a_n1214_n2088# 0.101196f
C297 drain_right.n1 a_n1214_n2088# 0.884107f
C298 minus.t1 a_n1214_n2088# 0.267737f
C299 minus.t0 a_n1214_n2088# 0.267727f
C300 minus.n0 a_n1214_n2088# 0.463477f
C301 minus.t3 a_n1214_n2088# 0.267737f
C302 minus.t2 a_n1214_n2088# 0.267727f
C303 minus.n1 a_n1214_n2088# 0.253002f
C304 minus.n2 a_n1214_n2088# 1.69289f
.ends

