* NGSPICE file created from diffpair439.ext - technology: sky130A

.subckt diffpair439 minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t1 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X1 source.t9 minus.t0 drain_right.t23 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X2 source.t4 minus.t1 drain_right.t22 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X3 drain_left.t0 plus.t1 source.t46 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X4 source.t10 minus.t2 drain_right.t21 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X5 drain_right.t20 minus.t3 source.t14 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X6 drain_right.t19 minus.t4 source.t6 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X7 drain_right.t18 minus.t5 source.t19 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X8 drain_right.t17 minus.t6 source.t23 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X9 source.t13 minus.t7 drain_right.t16 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X10 drain_left.t7 plus.t2 source.t45 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X11 source.t44 plus.t3 drain_left.t6 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X12 drain_left.t3 plus.t4 source.t43 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X13 source.t42 plus.t5 drain_left.t2 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X14 drain_left.t9 plus.t6 source.t41 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X15 drain_left.t8 plus.t7 source.t40 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X16 a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.3
X17 drain_right.t15 minus.t8 source.t0 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X18 source.t20 minus.t9 drain_right.t14 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X19 source.t12 minus.t10 drain_right.t13 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X20 source.t16 minus.t11 drain_right.t12 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X21 a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X22 source.t39 plus.t8 drain_left.t11 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X23 source.t21 minus.t12 drain_right.t11 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X24 drain_left.t10 plus.t9 source.t38 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X25 source.t37 plus.t10 drain_left.t15 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X26 drain_left.t14 plus.t11 source.t36 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X27 source.t1 minus.t13 drain_right.t10 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X28 source.t35 plus.t12 drain_left.t19 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X29 source.t34 plus.t13 drain_left.t18 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X30 source.t33 plus.t14 drain_left.t13 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X31 drain_right.t9 minus.t14 source.t8 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X32 drain_left.t12 plus.t15 source.t32 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X33 drain_right.t8 minus.t15 source.t11 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X34 drain_right.t7 minus.t16 source.t15 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X35 source.t5 minus.t17 drain_right.t6 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X36 source.t31 plus.t16 drain_left.t17 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X37 a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X38 drain_right.t5 minus.t18 source.t3 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X39 source.t30 plus.t17 drain_left.t16 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X40 drain_right.t4 minus.t19 source.t18 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X41 source.t29 plus.t18 drain_left.t5 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X42 drain_left.t4 plus.t19 source.t28 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X43 drain_right.t3 minus.t20 source.t17 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X44 drain_right.t2 minus.t21 source.t22 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X45 a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X46 drain_left.t23 plus.t20 source.t27 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X47 drain_left.t22 plus.t21 source.t26 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X48 source.t2 minus.t22 drain_right.t1 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X49 source.t7 minus.t23 drain_right.t0 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X50 source.t25 plus.t22 drain_left.t21 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X51 drain_left.t20 plus.t23 source.t24 a_n2354_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
R0 plus.n9 plus.t5 1099.84
R1 plus.n35 plus.t7 1099.84
R2 plus.n46 plus.t20 1099.84
R3 plus.n72 plus.t3 1099.84
R4 plus.n8 plus.t11 1068.43
R5 plus.n13 plus.t16 1068.43
R6 plus.n15 plus.t23 1068.43
R7 plus.n5 plus.t8 1068.43
R8 plus.n20 plus.t15 1068.43
R9 plus.n3 plus.t22 1068.43
R10 plus.n26 plus.t1 1068.43
R11 plus.n28 plus.t14 1068.43
R12 plus.n1 plus.t19 1068.43
R13 plus.n34 plus.t0 1068.43
R14 plus.n45 plus.t10 1068.43
R15 plus.n50 plus.t21 1068.43
R16 plus.n52 plus.t12 1068.43
R17 plus.n42 plus.t4 1068.43
R18 plus.n57 plus.t13 1068.43
R19 plus.n40 plus.t6 1068.43
R20 plus.n63 plus.t17 1068.43
R21 plus.n65 plus.t2 1068.43
R22 plus.n38 plus.t18 1068.43
R23 plus.n71 plus.t9 1068.43
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 31.8892
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus.n8 plus.n7 12.4157
R88 plus.n34 plus.n33 12.4157
R89 plus.n71 plus.n70 12.4157
R90 plus.n45 plus.n44 12.4157
R91 plus plus.n36 12.1141
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 drain_left.n13 drain_left.n11 60.0958
R125 drain_left.n7 drain_left.n5 60.0956
R126 drain_left.n2 drain_left.n0 60.0956
R127 drain_left.n19 drain_left.n18 59.5527
R128 drain_left.n17 drain_left.n16 59.5527
R129 drain_left.n15 drain_left.n14 59.5527
R130 drain_left.n13 drain_left.n12 59.5527
R131 drain_left.n7 drain_left.n6 59.5525
R132 drain_left.n9 drain_left.n8 59.5525
R133 drain_left.n4 drain_left.n3 59.5525
R134 drain_left.n2 drain_left.n1 59.5525
R135 drain_left.n21 drain_left.n20 59.5525
R136 drain_left drain_left.n10 32.5266
R137 drain_left drain_left.n21 6.19632
R138 drain_left.n5 drain_left.t15 1.6505
R139 drain_left.n5 drain_left.t23 1.6505
R140 drain_left.n6 drain_left.t19 1.6505
R141 drain_left.n6 drain_left.t22 1.6505
R142 drain_left.n8 drain_left.t18 1.6505
R143 drain_left.n8 drain_left.t3 1.6505
R144 drain_left.n3 drain_left.t16 1.6505
R145 drain_left.n3 drain_left.t9 1.6505
R146 drain_left.n1 drain_left.t5 1.6505
R147 drain_left.n1 drain_left.t7 1.6505
R148 drain_left.n0 drain_left.t6 1.6505
R149 drain_left.n0 drain_left.t10 1.6505
R150 drain_left.n20 drain_left.t1 1.6505
R151 drain_left.n20 drain_left.t8 1.6505
R152 drain_left.n18 drain_left.t13 1.6505
R153 drain_left.n18 drain_left.t4 1.6505
R154 drain_left.n16 drain_left.t21 1.6505
R155 drain_left.n16 drain_left.t0 1.6505
R156 drain_left.n14 drain_left.t11 1.6505
R157 drain_left.n14 drain_left.t12 1.6505
R158 drain_left.n12 drain_left.t17 1.6505
R159 drain_left.n12 drain_left.t20 1.6505
R160 drain_left.n11 drain_left.t2 1.6505
R161 drain_left.n11 drain_left.t14 1.6505
R162 drain_left.n9 drain_left.n7 0.543603
R163 drain_left.n4 drain_left.n2 0.543603
R164 drain_left.n15 drain_left.n13 0.543603
R165 drain_left.n17 drain_left.n15 0.543603
R166 drain_left.n19 drain_left.n17 0.543603
R167 drain_left.n21 drain_left.n19 0.543603
R168 drain_left.n10 drain_left.n9 0.216706
R169 drain_left.n10 drain_left.n4 0.216706
R170 source.n562 source.n502 289.615
R171 source.n486 source.n426 289.615
R172 source.n420 source.n360 289.615
R173 source.n344 source.n284 289.615
R174 source.n60 source.n0 289.615
R175 source.n136 source.n76 289.615
R176 source.n202 source.n142 289.615
R177 source.n278 source.n218 289.615
R178 source.n522 source.n521 185
R179 source.n527 source.n526 185
R180 source.n529 source.n528 185
R181 source.n518 source.n517 185
R182 source.n535 source.n534 185
R183 source.n537 source.n536 185
R184 source.n514 source.n513 185
R185 source.n544 source.n543 185
R186 source.n545 source.n512 185
R187 source.n547 source.n546 185
R188 source.n510 source.n509 185
R189 source.n553 source.n552 185
R190 source.n555 source.n554 185
R191 source.n506 source.n505 185
R192 source.n561 source.n560 185
R193 source.n563 source.n562 185
R194 source.n446 source.n445 185
R195 source.n451 source.n450 185
R196 source.n453 source.n452 185
R197 source.n442 source.n441 185
R198 source.n459 source.n458 185
R199 source.n461 source.n460 185
R200 source.n438 source.n437 185
R201 source.n468 source.n467 185
R202 source.n469 source.n436 185
R203 source.n471 source.n470 185
R204 source.n434 source.n433 185
R205 source.n477 source.n476 185
R206 source.n479 source.n478 185
R207 source.n430 source.n429 185
R208 source.n485 source.n484 185
R209 source.n487 source.n486 185
R210 source.n380 source.n379 185
R211 source.n385 source.n384 185
R212 source.n387 source.n386 185
R213 source.n376 source.n375 185
R214 source.n393 source.n392 185
R215 source.n395 source.n394 185
R216 source.n372 source.n371 185
R217 source.n402 source.n401 185
R218 source.n403 source.n370 185
R219 source.n405 source.n404 185
R220 source.n368 source.n367 185
R221 source.n411 source.n410 185
R222 source.n413 source.n412 185
R223 source.n364 source.n363 185
R224 source.n419 source.n418 185
R225 source.n421 source.n420 185
R226 source.n304 source.n303 185
R227 source.n309 source.n308 185
R228 source.n311 source.n310 185
R229 source.n300 source.n299 185
R230 source.n317 source.n316 185
R231 source.n319 source.n318 185
R232 source.n296 source.n295 185
R233 source.n326 source.n325 185
R234 source.n327 source.n294 185
R235 source.n329 source.n328 185
R236 source.n292 source.n291 185
R237 source.n335 source.n334 185
R238 source.n337 source.n336 185
R239 source.n288 source.n287 185
R240 source.n343 source.n342 185
R241 source.n345 source.n344 185
R242 source.n61 source.n60 185
R243 source.n59 source.n58 185
R244 source.n4 source.n3 185
R245 source.n53 source.n52 185
R246 source.n51 source.n50 185
R247 source.n8 source.n7 185
R248 source.n45 source.n44 185
R249 source.n43 source.n10 185
R250 source.n42 source.n41 185
R251 source.n13 source.n11 185
R252 source.n36 source.n35 185
R253 source.n34 source.n33 185
R254 source.n17 source.n16 185
R255 source.n28 source.n27 185
R256 source.n26 source.n25 185
R257 source.n21 source.n20 185
R258 source.n137 source.n136 185
R259 source.n135 source.n134 185
R260 source.n80 source.n79 185
R261 source.n129 source.n128 185
R262 source.n127 source.n126 185
R263 source.n84 source.n83 185
R264 source.n121 source.n120 185
R265 source.n119 source.n86 185
R266 source.n118 source.n117 185
R267 source.n89 source.n87 185
R268 source.n112 source.n111 185
R269 source.n110 source.n109 185
R270 source.n93 source.n92 185
R271 source.n104 source.n103 185
R272 source.n102 source.n101 185
R273 source.n97 source.n96 185
R274 source.n203 source.n202 185
R275 source.n201 source.n200 185
R276 source.n146 source.n145 185
R277 source.n195 source.n194 185
R278 source.n193 source.n192 185
R279 source.n150 source.n149 185
R280 source.n187 source.n186 185
R281 source.n185 source.n152 185
R282 source.n184 source.n183 185
R283 source.n155 source.n153 185
R284 source.n178 source.n177 185
R285 source.n176 source.n175 185
R286 source.n159 source.n158 185
R287 source.n170 source.n169 185
R288 source.n168 source.n167 185
R289 source.n163 source.n162 185
R290 source.n279 source.n278 185
R291 source.n277 source.n276 185
R292 source.n222 source.n221 185
R293 source.n271 source.n270 185
R294 source.n269 source.n268 185
R295 source.n226 source.n225 185
R296 source.n263 source.n262 185
R297 source.n261 source.n228 185
R298 source.n260 source.n259 185
R299 source.n231 source.n229 185
R300 source.n254 source.n253 185
R301 source.n252 source.n251 185
R302 source.n235 source.n234 185
R303 source.n246 source.n245 185
R304 source.n244 source.n243 185
R305 source.n239 source.n238 185
R306 source.n523 source.t14 149.524
R307 source.n447 source.t4 149.524
R308 source.n381 source.t27 149.524
R309 source.n305 source.t44 149.524
R310 source.n22 source.t40 149.524
R311 source.n98 source.t42 149.524
R312 source.n164 source.t8 149.524
R313 source.n240 source.t13 149.524
R314 source.n527 source.n521 104.615
R315 source.n528 source.n527 104.615
R316 source.n528 source.n517 104.615
R317 source.n535 source.n517 104.615
R318 source.n536 source.n535 104.615
R319 source.n536 source.n513 104.615
R320 source.n544 source.n513 104.615
R321 source.n545 source.n544 104.615
R322 source.n546 source.n545 104.615
R323 source.n546 source.n509 104.615
R324 source.n553 source.n509 104.615
R325 source.n554 source.n553 104.615
R326 source.n554 source.n505 104.615
R327 source.n561 source.n505 104.615
R328 source.n562 source.n561 104.615
R329 source.n451 source.n445 104.615
R330 source.n452 source.n451 104.615
R331 source.n452 source.n441 104.615
R332 source.n459 source.n441 104.615
R333 source.n460 source.n459 104.615
R334 source.n460 source.n437 104.615
R335 source.n468 source.n437 104.615
R336 source.n469 source.n468 104.615
R337 source.n470 source.n469 104.615
R338 source.n470 source.n433 104.615
R339 source.n477 source.n433 104.615
R340 source.n478 source.n477 104.615
R341 source.n478 source.n429 104.615
R342 source.n485 source.n429 104.615
R343 source.n486 source.n485 104.615
R344 source.n385 source.n379 104.615
R345 source.n386 source.n385 104.615
R346 source.n386 source.n375 104.615
R347 source.n393 source.n375 104.615
R348 source.n394 source.n393 104.615
R349 source.n394 source.n371 104.615
R350 source.n402 source.n371 104.615
R351 source.n403 source.n402 104.615
R352 source.n404 source.n403 104.615
R353 source.n404 source.n367 104.615
R354 source.n411 source.n367 104.615
R355 source.n412 source.n411 104.615
R356 source.n412 source.n363 104.615
R357 source.n419 source.n363 104.615
R358 source.n420 source.n419 104.615
R359 source.n309 source.n303 104.615
R360 source.n310 source.n309 104.615
R361 source.n310 source.n299 104.615
R362 source.n317 source.n299 104.615
R363 source.n318 source.n317 104.615
R364 source.n318 source.n295 104.615
R365 source.n326 source.n295 104.615
R366 source.n327 source.n326 104.615
R367 source.n328 source.n327 104.615
R368 source.n328 source.n291 104.615
R369 source.n335 source.n291 104.615
R370 source.n336 source.n335 104.615
R371 source.n336 source.n287 104.615
R372 source.n343 source.n287 104.615
R373 source.n344 source.n343 104.615
R374 source.n60 source.n59 104.615
R375 source.n59 source.n3 104.615
R376 source.n52 source.n3 104.615
R377 source.n52 source.n51 104.615
R378 source.n51 source.n7 104.615
R379 source.n44 source.n7 104.615
R380 source.n44 source.n43 104.615
R381 source.n43 source.n42 104.615
R382 source.n42 source.n11 104.615
R383 source.n35 source.n11 104.615
R384 source.n35 source.n34 104.615
R385 source.n34 source.n16 104.615
R386 source.n27 source.n16 104.615
R387 source.n27 source.n26 104.615
R388 source.n26 source.n20 104.615
R389 source.n136 source.n135 104.615
R390 source.n135 source.n79 104.615
R391 source.n128 source.n79 104.615
R392 source.n128 source.n127 104.615
R393 source.n127 source.n83 104.615
R394 source.n120 source.n83 104.615
R395 source.n120 source.n119 104.615
R396 source.n119 source.n118 104.615
R397 source.n118 source.n87 104.615
R398 source.n111 source.n87 104.615
R399 source.n111 source.n110 104.615
R400 source.n110 source.n92 104.615
R401 source.n103 source.n92 104.615
R402 source.n103 source.n102 104.615
R403 source.n102 source.n96 104.615
R404 source.n202 source.n201 104.615
R405 source.n201 source.n145 104.615
R406 source.n194 source.n145 104.615
R407 source.n194 source.n193 104.615
R408 source.n193 source.n149 104.615
R409 source.n186 source.n149 104.615
R410 source.n186 source.n185 104.615
R411 source.n185 source.n184 104.615
R412 source.n184 source.n153 104.615
R413 source.n177 source.n153 104.615
R414 source.n177 source.n176 104.615
R415 source.n176 source.n158 104.615
R416 source.n169 source.n158 104.615
R417 source.n169 source.n168 104.615
R418 source.n168 source.n162 104.615
R419 source.n278 source.n277 104.615
R420 source.n277 source.n221 104.615
R421 source.n270 source.n221 104.615
R422 source.n270 source.n269 104.615
R423 source.n269 source.n225 104.615
R424 source.n262 source.n225 104.615
R425 source.n262 source.n261 104.615
R426 source.n261 source.n260 104.615
R427 source.n260 source.n229 104.615
R428 source.n253 source.n229 104.615
R429 source.n253 source.n252 104.615
R430 source.n252 source.n234 104.615
R431 source.n245 source.n234 104.615
R432 source.n245 source.n244 104.615
R433 source.n244 source.n238 104.615
R434 source.t14 source.n521 52.3082
R435 source.t4 source.n445 52.3082
R436 source.t27 source.n379 52.3082
R437 source.t44 source.n303 52.3082
R438 source.t40 source.n20 52.3082
R439 source.t42 source.n96 52.3082
R440 source.t8 source.n162 52.3082
R441 source.t13 source.n238 52.3082
R442 source.n67 source.n66 42.8739
R443 source.n69 source.n68 42.8739
R444 source.n71 source.n70 42.8739
R445 source.n73 source.n72 42.8739
R446 source.n75 source.n74 42.8739
R447 source.n209 source.n208 42.8739
R448 source.n211 source.n210 42.8739
R449 source.n213 source.n212 42.8739
R450 source.n215 source.n214 42.8739
R451 source.n217 source.n216 42.8739
R452 source.n501 source.n500 42.8737
R453 source.n499 source.n498 42.8737
R454 source.n497 source.n496 42.8737
R455 source.n495 source.n494 42.8737
R456 source.n493 source.n492 42.8737
R457 source.n359 source.n358 42.8737
R458 source.n357 source.n356 42.8737
R459 source.n355 source.n354 42.8737
R460 source.n353 source.n352 42.8737
R461 source.n351 source.n350 42.8737
R462 source.n567 source.n566 29.8581
R463 source.n491 source.n490 29.8581
R464 source.n425 source.n424 29.8581
R465 source.n349 source.n348 29.8581
R466 source.n65 source.n64 29.8581
R467 source.n141 source.n140 29.8581
R468 source.n207 source.n206 29.8581
R469 source.n283 source.n282 29.8581
R470 source.n349 source.n283 21.8308
R471 source.n568 source.n65 16.2963
R472 source.n547 source.n512 13.1884
R473 source.n471 source.n436 13.1884
R474 source.n405 source.n370 13.1884
R475 source.n329 source.n294 13.1884
R476 source.n45 source.n10 13.1884
R477 source.n121 source.n86 13.1884
R478 source.n187 source.n152 13.1884
R479 source.n263 source.n228 13.1884
R480 source.n543 source.n542 12.8005
R481 source.n548 source.n510 12.8005
R482 source.n467 source.n466 12.8005
R483 source.n472 source.n434 12.8005
R484 source.n401 source.n400 12.8005
R485 source.n406 source.n368 12.8005
R486 source.n325 source.n324 12.8005
R487 source.n330 source.n292 12.8005
R488 source.n46 source.n8 12.8005
R489 source.n41 source.n12 12.8005
R490 source.n122 source.n84 12.8005
R491 source.n117 source.n88 12.8005
R492 source.n188 source.n150 12.8005
R493 source.n183 source.n154 12.8005
R494 source.n264 source.n226 12.8005
R495 source.n259 source.n230 12.8005
R496 source.n541 source.n514 12.0247
R497 source.n552 source.n551 12.0247
R498 source.n465 source.n438 12.0247
R499 source.n476 source.n475 12.0247
R500 source.n399 source.n372 12.0247
R501 source.n410 source.n409 12.0247
R502 source.n323 source.n296 12.0247
R503 source.n334 source.n333 12.0247
R504 source.n50 source.n49 12.0247
R505 source.n40 source.n13 12.0247
R506 source.n126 source.n125 12.0247
R507 source.n116 source.n89 12.0247
R508 source.n192 source.n191 12.0247
R509 source.n182 source.n155 12.0247
R510 source.n268 source.n267 12.0247
R511 source.n258 source.n231 12.0247
R512 source.n538 source.n537 11.249
R513 source.n555 source.n508 11.249
R514 source.n462 source.n461 11.249
R515 source.n479 source.n432 11.249
R516 source.n396 source.n395 11.249
R517 source.n413 source.n366 11.249
R518 source.n320 source.n319 11.249
R519 source.n337 source.n290 11.249
R520 source.n53 source.n6 11.249
R521 source.n37 source.n36 11.249
R522 source.n129 source.n82 11.249
R523 source.n113 source.n112 11.249
R524 source.n195 source.n148 11.249
R525 source.n179 source.n178 11.249
R526 source.n271 source.n224 11.249
R527 source.n255 source.n254 11.249
R528 source.n534 source.n516 10.4732
R529 source.n556 source.n506 10.4732
R530 source.n458 source.n440 10.4732
R531 source.n480 source.n430 10.4732
R532 source.n392 source.n374 10.4732
R533 source.n414 source.n364 10.4732
R534 source.n316 source.n298 10.4732
R535 source.n338 source.n288 10.4732
R536 source.n54 source.n4 10.4732
R537 source.n33 source.n15 10.4732
R538 source.n130 source.n80 10.4732
R539 source.n109 source.n91 10.4732
R540 source.n196 source.n146 10.4732
R541 source.n175 source.n157 10.4732
R542 source.n272 source.n222 10.4732
R543 source.n251 source.n233 10.4732
R544 source.n523 source.n522 10.2747
R545 source.n447 source.n446 10.2747
R546 source.n381 source.n380 10.2747
R547 source.n305 source.n304 10.2747
R548 source.n22 source.n21 10.2747
R549 source.n98 source.n97 10.2747
R550 source.n164 source.n163 10.2747
R551 source.n240 source.n239 10.2747
R552 source.n533 source.n518 9.69747
R553 source.n560 source.n559 9.69747
R554 source.n457 source.n442 9.69747
R555 source.n484 source.n483 9.69747
R556 source.n391 source.n376 9.69747
R557 source.n418 source.n417 9.69747
R558 source.n315 source.n300 9.69747
R559 source.n342 source.n341 9.69747
R560 source.n58 source.n57 9.69747
R561 source.n32 source.n17 9.69747
R562 source.n134 source.n133 9.69747
R563 source.n108 source.n93 9.69747
R564 source.n200 source.n199 9.69747
R565 source.n174 source.n159 9.69747
R566 source.n276 source.n275 9.69747
R567 source.n250 source.n235 9.69747
R568 source.n566 source.n565 9.45567
R569 source.n490 source.n489 9.45567
R570 source.n424 source.n423 9.45567
R571 source.n348 source.n347 9.45567
R572 source.n64 source.n63 9.45567
R573 source.n140 source.n139 9.45567
R574 source.n206 source.n205 9.45567
R575 source.n282 source.n281 9.45567
R576 source.n565 source.n564 9.3005
R577 source.n504 source.n503 9.3005
R578 source.n559 source.n558 9.3005
R579 source.n557 source.n556 9.3005
R580 source.n508 source.n507 9.3005
R581 source.n551 source.n550 9.3005
R582 source.n549 source.n548 9.3005
R583 source.n525 source.n524 9.3005
R584 source.n520 source.n519 9.3005
R585 source.n531 source.n530 9.3005
R586 source.n533 source.n532 9.3005
R587 source.n516 source.n515 9.3005
R588 source.n539 source.n538 9.3005
R589 source.n541 source.n540 9.3005
R590 source.n542 source.n511 9.3005
R591 source.n489 source.n488 9.3005
R592 source.n428 source.n427 9.3005
R593 source.n483 source.n482 9.3005
R594 source.n481 source.n480 9.3005
R595 source.n432 source.n431 9.3005
R596 source.n475 source.n474 9.3005
R597 source.n473 source.n472 9.3005
R598 source.n449 source.n448 9.3005
R599 source.n444 source.n443 9.3005
R600 source.n455 source.n454 9.3005
R601 source.n457 source.n456 9.3005
R602 source.n440 source.n439 9.3005
R603 source.n463 source.n462 9.3005
R604 source.n465 source.n464 9.3005
R605 source.n466 source.n435 9.3005
R606 source.n423 source.n422 9.3005
R607 source.n362 source.n361 9.3005
R608 source.n417 source.n416 9.3005
R609 source.n415 source.n414 9.3005
R610 source.n366 source.n365 9.3005
R611 source.n409 source.n408 9.3005
R612 source.n407 source.n406 9.3005
R613 source.n383 source.n382 9.3005
R614 source.n378 source.n377 9.3005
R615 source.n389 source.n388 9.3005
R616 source.n391 source.n390 9.3005
R617 source.n374 source.n373 9.3005
R618 source.n397 source.n396 9.3005
R619 source.n399 source.n398 9.3005
R620 source.n400 source.n369 9.3005
R621 source.n347 source.n346 9.3005
R622 source.n286 source.n285 9.3005
R623 source.n341 source.n340 9.3005
R624 source.n339 source.n338 9.3005
R625 source.n290 source.n289 9.3005
R626 source.n333 source.n332 9.3005
R627 source.n331 source.n330 9.3005
R628 source.n307 source.n306 9.3005
R629 source.n302 source.n301 9.3005
R630 source.n313 source.n312 9.3005
R631 source.n315 source.n314 9.3005
R632 source.n298 source.n297 9.3005
R633 source.n321 source.n320 9.3005
R634 source.n323 source.n322 9.3005
R635 source.n324 source.n293 9.3005
R636 source.n24 source.n23 9.3005
R637 source.n19 source.n18 9.3005
R638 source.n30 source.n29 9.3005
R639 source.n32 source.n31 9.3005
R640 source.n15 source.n14 9.3005
R641 source.n38 source.n37 9.3005
R642 source.n40 source.n39 9.3005
R643 source.n12 source.n9 9.3005
R644 source.n63 source.n62 9.3005
R645 source.n2 source.n1 9.3005
R646 source.n57 source.n56 9.3005
R647 source.n55 source.n54 9.3005
R648 source.n6 source.n5 9.3005
R649 source.n49 source.n48 9.3005
R650 source.n47 source.n46 9.3005
R651 source.n100 source.n99 9.3005
R652 source.n95 source.n94 9.3005
R653 source.n106 source.n105 9.3005
R654 source.n108 source.n107 9.3005
R655 source.n91 source.n90 9.3005
R656 source.n114 source.n113 9.3005
R657 source.n116 source.n115 9.3005
R658 source.n88 source.n85 9.3005
R659 source.n139 source.n138 9.3005
R660 source.n78 source.n77 9.3005
R661 source.n133 source.n132 9.3005
R662 source.n131 source.n130 9.3005
R663 source.n82 source.n81 9.3005
R664 source.n125 source.n124 9.3005
R665 source.n123 source.n122 9.3005
R666 source.n166 source.n165 9.3005
R667 source.n161 source.n160 9.3005
R668 source.n172 source.n171 9.3005
R669 source.n174 source.n173 9.3005
R670 source.n157 source.n156 9.3005
R671 source.n180 source.n179 9.3005
R672 source.n182 source.n181 9.3005
R673 source.n154 source.n151 9.3005
R674 source.n205 source.n204 9.3005
R675 source.n144 source.n143 9.3005
R676 source.n199 source.n198 9.3005
R677 source.n197 source.n196 9.3005
R678 source.n148 source.n147 9.3005
R679 source.n191 source.n190 9.3005
R680 source.n189 source.n188 9.3005
R681 source.n242 source.n241 9.3005
R682 source.n237 source.n236 9.3005
R683 source.n248 source.n247 9.3005
R684 source.n250 source.n249 9.3005
R685 source.n233 source.n232 9.3005
R686 source.n256 source.n255 9.3005
R687 source.n258 source.n257 9.3005
R688 source.n230 source.n227 9.3005
R689 source.n281 source.n280 9.3005
R690 source.n220 source.n219 9.3005
R691 source.n275 source.n274 9.3005
R692 source.n273 source.n272 9.3005
R693 source.n224 source.n223 9.3005
R694 source.n267 source.n266 9.3005
R695 source.n265 source.n264 9.3005
R696 source.n530 source.n529 8.92171
R697 source.n563 source.n504 8.92171
R698 source.n454 source.n453 8.92171
R699 source.n487 source.n428 8.92171
R700 source.n388 source.n387 8.92171
R701 source.n421 source.n362 8.92171
R702 source.n312 source.n311 8.92171
R703 source.n345 source.n286 8.92171
R704 source.n61 source.n2 8.92171
R705 source.n29 source.n28 8.92171
R706 source.n137 source.n78 8.92171
R707 source.n105 source.n104 8.92171
R708 source.n203 source.n144 8.92171
R709 source.n171 source.n170 8.92171
R710 source.n279 source.n220 8.92171
R711 source.n247 source.n246 8.92171
R712 source.n526 source.n520 8.14595
R713 source.n564 source.n502 8.14595
R714 source.n450 source.n444 8.14595
R715 source.n488 source.n426 8.14595
R716 source.n384 source.n378 8.14595
R717 source.n422 source.n360 8.14595
R718 source.n308 source.n302 8.14595
R719 source.n346 source.n284 8.14595
R720 source.n62 source.n0 8.14595
R721 source.n25 source.n19 8.14595
R722 source.n138 source.n76 8.14595
R723 source.n101 source.n95 8.14595
R724 source.n204 source.n142 8.14595
R725 source.n167 source.n161 8.14595
R726 source.n280 source.n218 8.14595
R727 source.n243 source.n237 8.14595
R728 source.n525 source.n522 7.3702
R729 source.n449 source.n446 7.3702
R730 source.n383 source.n380 7.3702
R731 source.n307 source.n304 7.3702
R732 source.n24 source.n21 7.3702
R733 source.n100 source.n97 7.3702
R734 source.n166 source.n163 7.3702
R735 source.n242 source.n239 7.3702
R736 source.n526 source.n525 5.81868
R737 source.n566 source.n502 5.81868
R738 source.n450 source.n449 5.81868
R739 source.n490 source.n426 5.81868
R740 source.n384 source.n383 5.81868
R741 source.n424 source.n360 5.81868
R742 source.n308 source.n307 5.81868
R743 source.n348 source.n284 5.81868
R744 source.n64 source.n0 5.81868
R745 source.n25 source.n24 5.81868
R746 source.n140 source.n76 5.81868
R747 source.n101 source.n100 5.81868
R748 source.n206 source.n142 5.81868
R749 source.n167 source.n166 5.81868
R750 source.n282 source.n218 5.81868
R751 source.n243 source.n242 5.81868
R752 source.n568 source.n567 5.53498
R753 source.n529 source.n520 5.04292
R754 source.n564 source.n563 5.04292
R755 source.n453 source.n444 5.04292
R756 source.n488 source.n487 5.04292
R757 source.n387 source.n378 5.04292
R758 source.n422 source.n421 5.04292
R759 source.n311 source.n302 5.04292
R760 source.n346 source.n345 5.04292
R761 source.n62 source.n61 5.04292
R762 source.n28 source.n19 5.04292
R763 source.n138 source.n137 5.04292
R764 source.n104 source.n95 5.04292
R765 source.n204 source.n203 5.04292
R766 source.n170 source.n161 5.04292
R767 source.n280 source.n279 5.04292
R768 source.n246 source.n237 5.04292
R769 source.n530 source.n518 4.26717
R770 source.n560 source.n504 4.26717
R771 source.n454 source.n442 4.26717
R772 source.n484 source.n428 4.26717
R773 source.n388 source.n376 4.26717
R774 source.n418 source.n362 4.26717
R775 source.n312 source.n300 4.26717
R776 source.n342 source.n286 4.26717
R777 source.n58 source.n2 4.26717
R778 source.n29 source.n17 4.26717
R779 source.n134 source.n78 4.26717
R780 source.n105 source.n93 4.26717
R781 source.n200 source.n144 4.26717
R782 source.n171 source.n159 4.26717
R783 source.n276 source.n220 4.26717
R784 source.n247 source.n235 4.26717
R785 source.n534 source.n533 3.49141
R786 source.n559 source.n506 3.49141
R787 source.n458 source.n457 3.49141
R788 source.n483 source.n430 3.49141
R789 source.n392 source.n391 3.49141
R790 source.n417 source.n364 3.49141
R791 source.n316 source.n315 3.49141
R792 source.n341 source.n288 3.49141
R793 source.n57 source.n4 3.49141
R794 source.n33 source.n32 3.49141
R795 source.n133 source.n80 3.49141
R796 source.n109 source.n108 3.49141
R797 source.n199 source.n146 3.49141
R798 source.n175 source.n174 3.49141
R799 source.n275 source.n222 3.49141
R800 source.n251 source.n250 3.49141
R801 source.n524 source.n523 2.84303
R802 source.n448 source.n447 2.84303
R803 source.n382 source.n381 2.84303
R804 source.n306 source.n305 2.84303
R805 source.n23 source.n22 2.84303
R806 source.n99 source.n98 2.84303
R807 source.n165 source.n164 2.84303
R808 source.n241 source.n240 2.84303
R809 source.n537 source.n516 2.71565
R810 source.n556 source.n555 2.71565
R811 source.n461 source.n440 2.71565
R812 source.n480 source.n479 2.71565
R813 source.n395 source.n374 2.71565
R814 source.n414 source.n413 2.71565
R815 source.n319 source.n298 2.71565
R816 source.n338 source.n337 2.71565
R817 source.n54 source.n53 2.71565
R818 source.n36 source.n15 2.71565
R819 source.n130 source.n129 2.71565
R820 source.n112 source.n91 2.71565
R821 source.n196 source.n195 2.71565
R822 source.n178 source.n157 2.71565
R823 source.n272 source.n271 2.71565
R824 source.n254 source.n233 2.71565
R825 source.n538 source.n514 1.93989
R826 source.n552 source.n508 1.93989
R827 source.n462 source.n438 1.93989
R828 source.n476 source.n432 1.93989
R829 source.n396 source.n372 1.93989
R830 source.n410 source.n366 1.93989
R831 source.n320 source.n296 1.93989
R832 source.n334 source.n290 1.93989
R833 source.n50 source.n6 1.93989
R834 source.n37 source.n13 1.93989
R835 source.n126 source.n82 1.93989
R836 source.n113 source.n89 1.93989
R837 source.n192 source.n148 1.93989
R838 source.n179 source.n155 1.93989
R839 source.n268 source.n224 1.93989
R840 source.n255 source.n231 1.93989
R841 source.n500 source.t6 1.6505
R842 source.n500 source.t21 1.6505
R843 source.n498 source.t3 1.6505
R844 source.n498 source.t5 1.6505
R845 source.n496 source.t18 1.6505
R846 source.n496 source.t12 1.6505
R847 source.n494 source.t11 1.6505
R848 source.n494 source.t16 1.6505
R849 source.n492 source.t15 1.6505
R850 source.n492 source.t9 1.6505
R851 source.n358 source.t26 1.6505
R852 source.n358 source.t37 1.6505
R853 source.n356 source.t43 1.6505
R854 source.n356 source.t35 1.6505
R855 source.n354 source.t41 1.6505
R856 source.n354 source.t34 1.6505
R857 source.n352 source.t45 1.6505
R858 source.n352 source.t30 1.6505
R859 source.n350 source.t38 1.6505
R860 source.n350 source.t29 1.6505
R861 source.n66 source.t28 1.6505
R862 source.n66 source.t47 1.6505
R863 source.n68 source.t46 1.6505
R864 source.n68 source.t33 1.6505
R865 source.n70 source.t32 1.6505
R866 source.n70 source.t25 1.6505
R867 source.n72 source.t24 1.6505
R868 source.n72 source.t39 1.6505
R869 source.n74 source.t36 1.6505
R870 source.n74 source.t31 1.6505
R871 source.n208 source.t19 1.6505
R872 source.n208 source.t2 1.6505
R873 source.n210 source.t17 1.6505
R874 source.n210 source.t1 1.6505
R875 source.n212 source.t0 1.6505
R876 source.n212 source.t10 1.6505
R877 source.n214 source.t23 1.6505
R878 source.n214 source.t7 1.6505
R879 source.n216 source.t22 1.6505
R880 source.n216 source.t20 1.6505
R881 source.n543 source.n541 1.16414
R882 source.n551 source.n510 1.16414
R883 source.n467 source.n465 1.16414
R884 source.n475 source.n434 1.16414
R885 source.n401 source.n399 1.16414
R886 source.n409 source.n368 1.16414
R887 source.n325 source.n323 1.16414
R888 source.n333 source.n292 1.16414
R889 source.n49 source.n8 1.16414
R890 source.n41 source.n40 1.16414
R891 source.n125 source.n84 1.16414
R892 source.n117 source.n116 1.16414
R893 source.n191 source.n150 1.16414
R894 source.n183 source.n182 1.16414
R895 source.n267 source.n226 1.16414
R896 source.n259 source.n258 1.16414
R897 source.n283 source.n217 0.543603
R898 source.n217 source.n215 0.543603
R899 source.n215 source.n213 0.543603
R900 source.n213 source.n211 0.543603
R901 source.n211 source.n209 0.543603
R902 source.n209 source.n207 0.543603
R903 source.n141 source.n75 0.543603
R904 source.n75 source.n73 0.543603
R905 source.n73 source.n71 0.543603
R906 source.n71 source.n69 0.543603
R907 source.n69 source.n67 0.543603
R908 source.n67 source.n65 0.543603
R909 source.n351 source.n349 0.543603
R910 source.n353 source.n351 0.543603
R911 source.n355 source.n353 0.543603
R912 source.n357 source.n355 0.543603
R913 source.n359 source.n357 0.543603
R914 source.n425 source.n359 0.543603
R915 source.n493 source.n491 0.543603
R916 source.n495 source.n493 0.543603
R917 source.n497 source.n495 0.543603
R918 source.n499 source.n497 0.543603
R919 source.n501 source.n499 0.543603
R920 source.n567 source.n501 0.543603
R921 source.n207 source.n141 0.470328
R922 source.n491 source.n425 0.470328
R923 source.n542 source.n512 0.388379
R924 source.n548 source.n547 0.388379
R925 source.n466 source.n436 0.388379
R926 source.n472 source.n471 0.388379
R927 source.n400 source.n370 0.388379
R928 source.n406 source.n405 0.388379
R929 source.n324 source.n294 0.388379
R930 source.n330 source.n329 0.388379
R931 source.n46 source.n45 0.388379
R932 source.n12 source.n10 0.388379
R933 source.n122 source.n121 0.388379
R934 source.n88 source.n86 0.388379
R935 source.n188 source.n187 0.388379
R936 source.n154 source.n152 0.388379
R937 source.n264 source.n263 0.388379
R938 source.n230 source.n228 0.388379
R939 source source.n568 0.188
R940 source.n524 source.n519 0.155672
R941 source.n531 source.n519 0.155672
R942 source.n532 source.n531 0.155672
R943 source.n532 source.n515 0.155672
R944 source.n539 source.n515 0.155672
R945 source.n540 source.n539 0.155672
R946 source.n540 source.n511 0.155672
R947 source.n549 source.n511 0.155672
R948 source.n550 source.n549 0.155672
R949 source.n550 source.n507 0.155672
R950 source.n557 source.n507 0.155672
R951 source.n558 source.n557 0.155672
R952 source.n558 source.n503 0.155672
R953 source.n565 source.n503 0.155672
R954 source.n448 source.n443 0.155672
R955 source.n455 source.n443 0.155672
R956 source.n456 source.n455 0.155672
R957 source.n456 source.n439 0.155672
R958 source.n463 source.n439 0.155672
R959 source.n464 source.n463 0.155672
R960 source.n464 source.n435 0.155672
R961 source.n473 source.n435 0.155672
R962 source.n474 source.n473 0.155672
R963 source.n474 source.n431 0.155672
R964 source.n481 source.n431 0.155672
R965 source.n482 source.n481 0.155672
R966 source.n482 source.n427 0.155672
R967 source.n489 source.n427 0.155672
R968 source.n382 source.n377 0.155672
R969 source.n389 source.n377 0.155672
R970 source.n390 source.n389 0.155672
R971 source.n390 source.n373 0.155672
R972 source.n397 source.n373 0.155672
R973 source.n398 source.n397 0.155672
R974 source.n398 source.n369 0.155672
R975 source.n407 source.n369 0.155672
R976 source.n408 source.n407 0.155672
R977 source.n408 source.n365 0.155672
R978 source.n415 source.n365 0.155672
R979 source.n416 source.n415 0.155672
R980 source.n416 source.n361 0.155672
R981 source.n423 source.n361 0.155672
R982 source.n306 source.n301 0.155672
R983 source.n313 source.n301 0.155672
R984 source.n314 source.n313 0.155672
R985 source.n314 source.n297 0.155672
R986 source.n321 source.n297 0.155672
R987 source.n322 source.n321 0.155672
R988 source.n322 source.n293 0.155672
R989 source.n331 source.n293 0.155672
R990 source.n332 source.n331 0.155672
R991 source.n332 source.n289 0.155672
R992 source.n339 source.n289 0.155672
R993 source.n340 source.n339 0.155672
R994 source.n340 source.n285 0.155672
R995 source.n347 source.n285 0.155672
R996 source.n63 source.n1 0.155672
R997 source.n56 source.n1 0.155672
R998 source.n56 source.n55 0.155672
R999 source.n55 source.n5 0.155672
R1000 source.n48 source.n5 0.155672
R1001 source.n48 source.n47 0.155672
R1002 source.n47 source.n9 0.155672
R1003 source.n39 source.n9 0.155672
R1004 source.n39 source.n38 0.155672
R1005 source.n38 source.n14 0.155672
R1006 source.n31 source.n14 0.155672
R1007 source.n31 source.n30 0.155672
R1008 source.n30 source.n18 0.155672
R1009 source.n23 source.n18 0.155672
R1010 source.n139 source.n77 0.155672
R1011 source.n132 source.n77 0.155672
R1012 source.n132 source.n131 0.155672
R1013 source.n131 source.n81 0.155672
R1014 source.n124 source.n81 0.155672
R1015 source.n124 source.n123 0.155672
R1016 source.n123 source.n85 0.155672
R1017 source.n115 source.n85 0.155672
R1018 source.n115 source.n114 0.155672
R1019 source.n114 source.n90 0.155672
R1020 source.n107 source.n90 0.155672
R1021 source.n107 source.n106 0.155672
R1022 source.n106 source.n94 0.155672
R1023 source.n99 source.n94 0.155672
R1024 source.n205 source.n143 0.155672
R1025 source.n198 source.n143 0.155672
R1026 source.n198 source.n197 0.155672
R1027 source.n197 source.n147 0.155672
R1028 source.n190 source.n147 0.155672
R1029 source.n190 source.n189 0.155672
R1030 source.n189 source.n151 0.155672
R1031 source.n181 source.n151 0.155672
R1032 source.n181 source.n180 0.155672
R1033 source.n180 source.n156 0.155672
R1034 source.n173 source.n156 0.155672
R1035 source.n173 source.n172 0.155672
R1036 source.n172 source.n160 0.155672
R1037 source.n165 source.n160 0.155672
R1038 source.n281 source.n219 0.155672
R1039 source.n274 source.n219 0.155672
R1040 source.n274 source.n273 0.155672
R1041 source.n273 source.n223 0.155672
R1042 source.n266 source.n223 0.155672
R1043 source.n266 source.n265 0.155672
R1044 source.n265 source.n227 0.155672
R1045 source.n257 source.n227 0.155672
R1046 source.n257 source.n256 0.155672
R1047 source.n256 source.n232 0.155672
R1048 source.n249 source.n232 0.155672
R1049 source.n249 source.n248 0.155672
R1050 source.n248 source.n236 0.155672
R1051 source.n241 source.n236 0.155672
R1052 minus.n35 minus.t7 1099.84
R1053 minus.n9 minus.t14 1099.84
R1054 minus.n72 minus.t3 1099.84
R1055 minus.n46 minus.t1 1099.84
R1056 minus.n34 minus.t21 1068.43
R1057 minus.n1 minus.t9 1068.43
R1058 minus.n28 minus.t6 1068.43
R1059 minus.n26 minus.t23 1068.43
R1060 minus.n3 minus.t8 1068.43
R1061 minus.n20 minus.t2 1068.43
R1062 minus.n5 minus.t20 1068.43
R1063 minus.n15 minus.t13 1068.43
R1064 minus.n13 minus.t5 1068.43
R1065 minus.n8 minus.t22 1068.43
R1066 minus.n71 minus.t12 1068.43
R1067 minus.n38 minus.t4 1068.43
R1068 minus.n65 minus.t17 1068.43
R1069 minus.n63 minus.t18 1068.43
R1070 minus.n40 minus.t10 1068.43
R1071 minus.n57 minus.t19 1068.43
R1072 minus.n42 minus.t11 1068.43
R1073 minus.n52 minus.t15 1068.43
R1074 minus.n50 minus.t0 1068.43
R1075 minus.n45 minus.t16 1068.43
R1076 minus.n10 minus.n9 161.489
R1077 minus.n47 minus.n46 161.489
R1078 minus.n36 minus.n35 161.3
R1079 minus.n33 minus.n0 161.3
R1080 minus.n32 minus.n31 161.3
R1081 minus.n30 minus.n29 161.3
R1082 minus.n27 minus.n2 161.3
R1083 minus.n25 minus.n24 161.3
R1084 minus.n23 minus.n22 161.3
R1085 minus.n21 minus.n4 161.3
R1086 minus.n19 minus.n18 161.3
R1087 minus.n17 minus.n16 161.3
R1088 minus.n14 minus.n6 161.3
R1089 minus.n12 minus.n11 161.3
R1090 minus.n10 minus.n7 161.3
R1091 minus.n73 minus.n72 161.3
R1092 minus.n70 minus.n37 161.3
R1093 minus.n69 minus.n68 161.3
R1094 minus.n67 minus.n66 161.3
R1095 minus.n64 minus.n39 161.3
R1096 minus.n62 minus.n61 161.3
R1097 minus.n60 minus.n59 161.3
R1098 minus.n58 minus.n41 161.3
R1099 minus.n56 minus.n55 161.3
R1100 minus.n54 minus.n53 161.3
R1101 minus.n51 minus.n43 161.3
R1102 minus.n49 minus.n48 161.3
R1103 minus.n47 minus.n44 161.3
R1104 minus.n33 minus.n32 73.0308
R1105 minus.n22 minus.n21 73.0308
R1106 minus.n12 minus.n7 73.0308
R1107 minus.n49 minus.n44 73.0308
R1108 minus.n59 minus.n58 73.0308
R1109 minus.n70 minus.n69 73.0308
R1110 minus.n29 minus.n1 66.4581
R1111 minus.n14 minus.n13 66.4581
R1112 minus.n51 minus.n50 66.4581
R1113 minus.n66 minus.n38 66.4581
R1114 minus.n25 minus.n3 63.5369
R1115 minus.n20 minus.n19 63.5369
R1116 minus.n57 minus.n56 63.5369
R1117 minus.n62 minus.n40 63.5369
R1118 minus.n35 minus.n34 60.6157
R1119 minus.n9 minus.n8 60.6157
R1120 minus.n46 minus.n45 60.6157
R1121 minus.n72 minus.n71 60.6157
R1122 minus.n28 minus.n27 47.4702
R1123 minus.n16 minus.n15 47.4702
R1124 minus.n53 minus.n52 47.4702
R1125 minus.n65 minus.n64 47.4702
R1126 minus.n27 minus.n26 44.549
R1127 minus.n16 minus.n5 44.549
R1128 minus.n53 minus.n42 44.549
R1129 minus.n64 minus.n63 44.549
R1130 minus.n74 minus.n36 38.0081
R1131 minus.n26 minus.n25 28.4823
R1132 minus.n19 minus.n5 28.4823
R1133 minus.n56 minus.n42 28.4823
R1134 minus.n63 minus.n62 28.4823
R1135 minus.n29 minus.n28 25.5611
R1136 minus.n15 minus.n14 25.5611
R1137 minus.n52 minus.n51 25.5611
R1138 minus.n66 minus.n65 25.5611
R1139 minus.n34 minus.n33 12.4157
R1140 minus.n8 minus.n7 12.4157
R1141 minus.n45 minus.n44 12.4157
R1142 minus.n71 minus.n70 12.4157
R1143 minus.n22 minus.n3 9.49444
R1144 minus.n21 minus.n20 9.49444
R1145 minus.n58 minus.n57 9.49444
R1146 minus.n59 minus.n40 9.49444
R1147 minus.n32 minus.n1 6.57323
R1148 minus.n13 minus.n12 6.57323
R1149 minus.n50 minus.n49 6.57323
R1150 minus.n69 minus.n38 6.57323
R1151 minus.n74 minus.n73 6.4702
R1152 minus.n36 minus.n0 0.189894
R1153 minus.n31 minus.n0 0.189894
R1154 minus.n31 minus.n30 0.189894
R1155 minus.n30 minus.n2 0.189894
R1156 minus.n24 minus.n2 0.189894
R1157 minus.n24 minus.n23 0.189894
R1158 minus.n23 minus.n4 0.189894
R1159 minus.n18 minus.n4 0.189894
R1160 minus.n18 minus.n17 0.189894
R1161 minus.n17 minus.n6 0.189894
R1162 minus.n11 minus.n6 0.189894
R1163 minus.n11 minus.n10 0.189894
R1164 minus.n48 minus.n47 0.189894
R1165 minus.n48 minus.n43 0.189894
R1166 minus.n54 minus.n43 0.189894
R1167 minus.n55 minus.n54 0.189894
R1168 minus.n55 minus.n41 0.189894
R1169 minus.n60 minus.n41 0.189894
R1170 minus.n61 minus.n60 0.189894
R1171 minus.n61 minus.n39 0.189894
R1172 minus.n67 minus.n39 0.189894
R1173 minus.n68 minus.n67 0.189894
R1174 minus.n68 minus.n37 0.189894
R1175 minus.n73 minus.n37 0.189894
R1176 minus minus.n74 0.188
R1177 drain_right.n7 drain_right.n5 60.0956
R1178 drain_right.n2 drain_right.n0 60.0956
R1179 drain_right.n13 drain_right.n11 60.0956
R1180 drain_right.n13 drain_right.n12 59.5527
R1181 drain_right.n15 drain_right.n14 59.5527
R1182 drain_right.n17 drain_right.n16 59.5527
R1183 drain_right.n19 drain_right.n18 59.5527
R1184 drain_right.n21 drain_right.n20 59.5527
R1185 drain_right.n7 drain_right.n6 59.5525
R1186 drain_right.n9 drain_right.n8 59.5525
R1187 drain_right.n4 drain_right.n3 59.5525
R1188 drain_right.n2 drain_right.n1 59.5525
R1189 drain_right drain_right.n10 31.9733
R1190 drain_right drain_right.n21 6.19632
R1191 drain_right.n5 drain_right.t11 1.6505
R1192 drain_right.n5 drain_right.t20 1.6505
R1193 drain_right.n6 drain_right.t6 1.6505
R1194 drain_right.n6 drain_right.t19 1.6505
R1195 drain_right.n8 drain_right.t13 1.6505
R1196 drain_right.n8 drain_right.t5 1.6505
R1197 drain_right.n3 drain_right.t12 1.6505
R1198 drain_right.n3 drain_right.t4 1.6505
R1199 drain_right.n1 drain_right.t23 1.6505
R1200 drain_right.n1 drain_right.t8 1.6505
R1201 drain_right.n0 drain_right.t22 1.6505
R1202 drain_right.n0 drain_right.t7 1.6505
R1203 drain_right.n11 drain_right.t1 1.6505
R1204 drain_right.n11 drain_right.t9 1.6505
R1205 drain_right.n12 drain_right.t10 1.6505
R1206 drain_right.n12 drain_right.t18 1.6505
R1207 drain_right.n14 drain_right.t21 1.6505
R1208 drain_right.n14 drain_right.t3 1.6505
R1209 drain_right.n16 drain_right.t0 1.6505
R1210 drain_right.n16 drain_right.t15 1.6505
R1211 drain_right.n18 drain_right.t14 1.6505
R1212 drain_right.n18 drain_right.t17 1.6505
R1213 drain_right.n20 drain_right.t16 1.6505
R1214 drain_right.n20 drain_right.t2 1.6505
R1215 drain_right.n9 drain_right.n7 0.543603
R1216 drain_right.n4 drain_right.n2 0.543603
R1217 drain_right.n21 drain_right.n19 0.543603
R1218 drain_right.n19 drain_right.n17 0.543603
R1219 drain_right.n17 drain_right.n15 0.543603
R1220 drain_right.n15 drain_right.n13 0.543603
R1221 drain_right.n10 drain_right.n9 0.216706
R1222 drain_right.n10 drain_right.n4 0.216706
C0 drain_right plus 0.387992f
C1 plus minus 6.09401f
C2 drain_right minus 8.43656f
C3 source plus 8.26809f
C4 drain_left plus 8.668759f
C5 source drain_right 44.431396f
C6 source minus 8.254049f
C7 drain_left drain_right 1.26597f
C8 drain_left minus 0.172624f
C9 drain_left source 44.4307f
C10 drain_right a_n2354_n3288# 7.35467f
C11 drain_left a_n2354_n3288# 7.71183f
C12 source a_n2354_n3288# 8.916337f
C13 minus a_n2354_n3288# 9.27826f
C14 plus a_n2354_n3288# 11.341109f
C15 drain_right.t22 a_n2354_n3288# 0.324124f
C16 drain_right.t7 a_n2354_n3288# 0.324124f
C17 drain_right.n0 a_n2354_n3288# 2.888f
C18 drain_right.t23 a_n2354_n3288# 0.324124f
C19 drain_right.t8 a_n2354_n3288# 0.324124f
C20 drain_right.n1 a_n2354_n3288# 2.8842f
C21 drain_right.n2 a_n2354_n3288# 0.822952f
C22 drain_right.t12 a_n2354_n3288# 0.324124f
C23 drain_right.t4 a_n2354_n3288# 0.324124f
C24 drain_right.n3 a_n2354_n3288# 2.8842f
C25 drain_right.n4 a_n2354_n3288# 0.374153f
C26 drain_right.t11 a_n2354_n3288# 0.324124f
C27 drain_right.t20 a_n2354_n3288# 0.324124f
C28 drain_right.n5 a_n2354_n3288# 2.888f
C29 drain_right.t6 a_n2354_n3288# 0.324124f
C30 drain_right.t19 a_n2354_n3288# 0.324124f
C31 drain_right.n6 a_n2354_n3288# 2.8842f
C32 drain_right.n7 a_n2354_n3288# 0.822952f
C33 drain_right.t13 a_n2354_n3288# 0.324124f
C34 drain_right.t5 a_n2354_n3288# 0.324124f
C35 drain_right.n8 a_n2354_n3288# 2.8842f
C36 drain_right.n9 a_n2354_n3288# 0.374153f
C37 drain_right.n10 a_n2354_n3288# 1.78411f
C38 drain_right.t1 a_n2354_n3288# 0.324124f
C39 drain_right.t9 a_n2354_n3288# 0.324124f
C40 drain_right.n11 a_n2354_n3288# 2.888f
C41 drain_right.t10 a_n2354_n3288# 0.324124f
C42 drain_right.t18 a_n2354_n3288# 0.324124f
C43 drain_right.n12 a_n2354_n3288# 2.88421f
C44 drain_right.n13 a_n2354_n3288# 0.82294f
C45 drain_right.t21 a_n2354_n3288# 0.324124f
C46 drain_right.t3 a_n2354_n3288# 0.324124f
C47 drain_right.n14 a_n2354_n3288# 2.88421f
C48 drain_right.n15 a_n2354_n3288# 0.40648f
C49 drain_right.t0 a_n2354_n3288# 0.324124f
C50 drain_right.t15 a_n2354_n3288# 0.324124f
C51 drain_right.n16 a_n2354_n3288# 2.88421f
C52 drain_right.n17 a_n2354_n3288# 0.40648f
C53 drain_right.t14 a_n2354_n3288# 0.324124f
C54 drain_right.t17 a_n2354_n3288# 0.324124f
C55 drain_right.n18 a_n2354_n3288# 2.88421f
C56 drain_right.n19 a_n2354_n3288# 0.40648f
C57 drain_right.t16 a_n2354_n3288# 0.324124f
C58 drain_right.t2 a_n2354_n3288# 0.324124f
C59 drain_right.n20 a_n2354_n3288# 2.88421f
C60 drain_right.n21 a_n2354_n3288# 0.690984f
C61 minus.n0 a_n2354_n3288# 0.048547f
C62 minus.t7 a_n2354_n3288# 0.49947f
C63 minus.t21 a_n2354_n3288# 0.493864f
C64 minus.t9 a_n2354_n3288# 0.493864f
C65 minus.n1 a_n2354_n3288# 0.195913f
C66 minus.n2 a_n2354_n3288# 0.048547f
C67 minus.t6 a_n2354_n3288# 0.493864f
C68 minus.t23 a_n2354_n3288# 0.493864f
C69 minus.t8 a_n2354_n3288# 0.493864f
C70 minus.n3 a_n2354_n3288# 0.195913f
C71 minus.n4 a_n2354_n3288# 0.048547f
C72 minus.t2 a_n2354_n3288# 0.493864f
C73 minus.t20 a_n2354_n3288# 0.493864f
C74 minus.n5 a_n2354_n3288# 0.195913f
C75 minus.n6 a_n2354_n3288# 0.048547f
C76 minus.t13 a_n2354_n3288# 0.493864f
C77 minus.t5 a_n2354_n3288# 0.493864f
C78 minus.n7 a_n2354_n3288# 0.018649f
C79 minus.t22 a_n2354_n3288# 0.493864f
C80 minus.n8 a_n2354_n3288# 0.195913f
C81 minus.t14 a_n2354_n3288# 0.49947f
C82 minus.n9 a_n2354_n3288# 0.210816f
C83 minus.n10 a_n2354_n3288# 0.103913f
C84 minus.n11 a_n2354_n3288# 0.048547f
C85 minus.n12 a_n2354_n3288# 0.017451f
C86 minus.n13 a_n2354_n3288# 0.195913f
C87 minus.n14 a_n2354_n3288# 0.019996f
C88 minus.n15 a_n2354_n3288# 0.195913f
C89 minus.n16 a_n2354_n3288# 0.019996f
C90 minus.n17 a_n2354_n3288# 0.048547f
C91 minus.n18 a_n2354_n3288# 0.048547f
C92 minus.n19 a_n2354_n3288# 0.019996f
C93 minus.n20 a_n2354_n3288# 0.195913f
C94 minus.n21 a_n2354_n3288# 0.01805f
C95 minus.n22 a_n2354_n3288# 0.01805f
C96 minus.n23 a_n2354_n3288# 0.048547f
C97 minus.n24 a_n2354_n3288# 0.048547f
C98 minus.n25 a_n2354_n3288# 0.019996f
C99 minus.n26 a_n2354_n3288# 0.195913f
C100 minus.n27 a_n2354_n3288# 0.019996f
C101 minus.n28 a_n2354_n3288# 0.195913f
C102 minus.n29 a_n2354_n3288# 0.019996f
C103 minus.n30 a_n2354_n3288# 0.048547f
C104 minus.n31 a_n2354_n3288# 0.048547f
C105 minus.n32 a_n2354_n3288# 0.017451f
C106 minus.n33 a_n2354_n3288# 0.018649f
C107 minus.n34 a_n2354_n3288# 0.195913f
C108 minus.n35 a_n2354_n3288# 0.210751f
C109 minus.n36 a_n2354_n3288# 1.84952f
C110 minus.n37 a_n2354_n3288# 0.048547f
C111 minus.t12 a_n2354_n3288# 0.493864f
C112 minus.t4 a_n2354_n3288# 0.493864f
C113 minus.n38 a_n2354_n3288# 0.195913f
C114 minus.n39 a_n2354_n3288# 0.048547f
C115 minus.t17 a_n2354_n3288# 0.493864f
C116 minus.t18 a_n2354_n3288# 0.493864f
C117 minus.t10 a_n2354_n3288# 0.493864f
C118 minus.n40 a_n2354_n3288# 0.195913f
C119 minus.n41 a_n2354_n3288# 0.048547f
C120 minus.t19 a_n2354_n3288# 0.493864f
C121 minus.t11 a_n2354_n3288# 0.493864f
C122 minus.n42 a_n2354_n3288# 0.195913f
C123 minus.n43 a_n2354_n3288# 0.048547f
C124 minus.t15 a_n2354_n3288# 0.493864f
C125 minus.t0 a_n2354_n3288# 0.493864f
C126 minus.n44 a_n2354_n3288# 0.018649f
C127 minus.t1 a_n2354_n3288# 0.49947f
C128 minus.t16 a_n2354_n3288# 0.493864f
C129 minus.n45 a_n2354_n3288# 0.195913f
C130 minus.n46 a_n2354_n3288# 0.210816f
C131 minus.n47 a_n2354_n3288# 0.103913f
C132 minus.n48 a_n2354_n3288# 0.048547f
C133 minus.n49 a_n2354_n3288# 0.017451f
C134 minus.n50 a_n2354_n3288# 0.195913f
C135 minus.n51 a_n2354_n3288# 0.019996f
C136 minus.n52 a_n2354_n3288# 0.195913f
C137 minus.n53 a_n2354_n3288# 0.019996f
C138 minus.n54 a_n2354_n3288# 0.048547f
C139 minus.n55 a_n2354_n3288# 0.048547f
C140 minus.n56 a_n2354_n3288# 0.019996f
C141 minus.n57 a_n2354_n3288# 0.195913f
C142 minus.n58 a_n2354_n3288# 0.01805f
C143 minus.n59 a_n2354_n3288# 0.01805f
C144 minus.n60 a_n2354_n3288# 0.048547f
C145 minus.n61 a_n2354_n3288# 0.048547f
C146 minus.n62 a_n2354_n3288# 0.019996f
C147 minus.n63 a_n2354_n3288# 0.195913f
C148 minus.n64 a_n2354_n3288# 0.019996f
C149 minus.n65 a_n2354_n3288# 0.195913f
C150 minus.n66 a_n2354_n3288# 0.019996f
C151 minus.n67 a_n2354_n3288# 0.048547f
C152 minus.n68 a_n2354_n3288# 0.048547f
C153 minus.n69 a_n2354_n3288# 0.017451f
C154 minus.n70 a_n2354_n3288# 0.018649f
C155 minus.n71 a_n2354_n3288# 0.195913f
C156 minus.t3 a_n2354_n3288# 0.49947f
C157 minus.n72 a_n2354_n3288# 0.210751f
C158 minus.n73 a_n2354_n3288# 0.313973f
C159 minus.n74 a_n2354_n3288# 2.23567f
C160 source.n0 a_n2354_n3288# 0.040444f
C161 source.n1 a_n2354_n3288# 0.030532f
C162 source.n2 a_n2354_n3288# 0.016407f
C163 source.n3 a_n2354_n3288# 0.038779f
C164 source.n4 a_n2354_n3288# 0.017372f
C165 source.n5 a_n2354_n3288# 0.030532f
C166 source.n6 a_n2354_n3288# 0.016407f
C167 source.n7 a_n2354_n3288# 0.038779f
C168 source.n8 a_n2354_n3288# 0.017372f
C169 source.n9 a_n2354_n3288# 0.030532f
C170 source.n10 a_n2354_n3288# 0.016889f
C171 source.n11 a_n2354_n3288# 0.038779f
C172 source.n12 a_n2354_n3288# 0.016407f
C173 source.n13 a_n2354_n3288# 0.017372f
C174 source.n14 a_n2354_n3288# 0.030532f
C175 source.n15 a_n2354_n3288# 0.016407f
C176 source.n16 a_n2354_n3288# 0.038779f
C177 source.n17 a_n2354_n3288# 0.017372f
C178 source.n18 a_n2354_n3288# 0.030532f
C179 source.n19 a_n2354_n3288# 0.016407f
C180 source.n20 a_n2354_n3288# 0.029084f
C181 source.n21 a_n2354_n3288# 0.027414f
C182 source.t40 a_n2354_n3288# 0.065495f
C183 source.n22 a_n2354_n3288# 0.220132f
C184 source.n23 a_n2354_n3288# 1.54029f
C185 source.n24 a_n2354_n3288# 0.016407f
C186 source.n25 a_n2354_n3288# 0.017372f
C187 source.n26 a_n2354_n3288# 0.038779f
C188 source.n27 a_n2354_n3288# 0.038779f
C189 source.n28 a_n2354_n3288# 0.017372f
C190 source.n29 a_n2354_n3288# 0.016407f
C191 source.n30 a_n2354_n3288# 0.030532f
C192 source.n31 a_n2354_n3288# 0.030532f
C193 source.n32 a_n2354_n3288# 0.016407f
C194 source.n33 a_n2354_n3288# 0.017372f
C195 source.n34 a_n2354_n3288# 0.038779f
C196 source.n35 a_n2354_n3288# 0.038779f
C197 source.n36 a_n2354_n3288# 0.017372f
C198 source.n37 a_n2354_n3288# 0.016407f
C199 source.n38 a_n2354_n3288# 0.030532f
C200 source.n39 a_n2354_n3288# 0.030532f
C201 source.n40 a_n2354_n3288# 0.016407f
C202 source.n41 a_n2354_n3288# 0.017372f
C203 source.n42 a_n2354_n3288# 0.038779f
C204 source.n43 a_n2354_n3288# 0.038779f
C205 source.n44 a_n2354_n3288# 0.038779f
C206 source.n45 a_n2354_n3288# 0.016889f
C207 source.n46 a_n2354_n3288# 0.016407f
C208 source.n47 a_n2354_n3288# 0.030532f
C209 source.n48 a_n2354_n3288# 0.030532f
C210 source.n49 a_n2354_n3288# 0.016407f
C211 source.n50 a_n2354_n3288# 0.017372f
C212 source.n51 a_n2354_n3288# 0.038779f
C213 source.n52 a_n2354_n3288# 0.038779f
C214 source.n53 a_n2354_n3288# 0.017372f
C215 source.n54 a_n2354_n3288# 0.016407f
C216 source.n55 a_n2354_n3288# 0.030532f
C217 source.n56 a_n2354_n3288# 0.030532f
C218 source.n57 a_n2354_n3288# 0.016407f
C219 source.n58 a_n2354_n3288# 0.017372f
C220 source.n59 a_n2354_n3288# 0.038779f
C221 source.n60 a_n2354_n3288# 0.079579f
C222 source.n61 a_n2354_n3288# 0.017372f
C223 source.n62 a_n2354_n3288# 0.016407f
C224 source.n63 a_n2354_n3288# 0.065568f
C225 source.n64 a_n2354_n3288# 0.043919f
C226 source.n65 a_n2354_n3288# 1.22876f
C227 source.t28 a_n2354_n3288# 0.289528f
C228 source.t47 a_n2354_n3288# 0.289528f
C229 source.n66 a_n2354_n3288# 2.47894f
C230 source.n67 a_n2354_n3288# 0.419013f
C231 source.t46 a_n2354_n3288# 0.289528f
C232 source.t33 a_n2354_n3288# 0.289528f
C233 source.n68 a_n2354_n3288# 2.47894f
C234 source.n69 a_n2354_n3288# 0.419013f
C235 source.t32 a_n2354_n3288# 0.289528f
C236 source.t25 a_n2354_n3288# 0.289528f
C237 source.n70 a_n2354_n3288# 2.47894f
C238 source.n71 a_n2354_n3288# 0.419013f
C239 source.t24 a_n2354_n3288# 0.289528f
C240 source.t39 a_n2354_n3288# 0.289528f
C241 source.n72 a_n2354_n3288# 2.47894f
C242 source.n73 a_n2354_n3288# 0.419013f
C243 source.t36 a_n2354_n3288# 0.289528f
C244 source.t31 a_n2354_n3288# 0.289528f
C245 source.n74 a_n2354_n3288# 2.47894f
C246 source.n75 a_n2354_n3288# 0.419013f
C247 source.n76 a_n2354_n3288# 0.040444f
C248 source.n77 a_n2354_n3288# 0.030532f
C249 source.n78 a_n2354_n3288# 0.016407f
C250 source.n79 a_n2354_n3288# 0.038779f
C251 source.n80 a_n2354_n3288# 0.017372f
C252 source.n81 a_n2354_n3288# 0.030532f
C253 source.n82 a_n2354_n3288# 0.016407f
C254 source.n83 a_n2354_n3288# 0.038779f
C255 source.n84 a_n2354_n3288# 0.017372f
C256 source.n85 a_n2354_n3288# 0.030532f
C257 source.n86 a_n2354_n3288# 0.016889f
C258 source.n87 a_n2354_n3288# 0.038779f
C259 source.n88 a_n2354_n3288# 0.016407f
C260 source.n89 a_n2354_n3288# 0.017372f
C261 source.n90 a_n2354_n3288# 0.030532f
C262 source.n91 a_n2354_n3288# 0.016407f
C263 source.n92 a_n2354_n3288# 0.038779f
C264 source.n93 a_n2354_n3288# 0.017372f
C265 source.n94 a_n2354_n3288# 0.030532f
C266 source.n95 a_n2354_n3288# 0.016407f
C267 source.n96 a_n2354_n3288# 0.029084f
C268 source.n97 a_n2354_n3288# 0.027414f
C269 source.t42 a_n2354_n3288# 0.065495f
C270 source.n98 a_n2354_n3288# 0.220132f
C271 source.n99 a_n2354_n3288# 1.54029f
C272 source.n100 a_n2354_n3288# 0.016407f
C273 source.n101 a_n2354_n3288# 0.017372f
C274 source.n102 a_n2354_n3288# 0.038779f
C275 source.n103 a_n2354_n3288# 0.038779f
C276 source.n104 a_n2354_n3288# 0.017372f
C277 source.n105 a_n2354_n3288# 0.016407f
C278 source.n106 a_n2354_n3288# 0.030532f
C279 source.n107 a_n2354_n3288# 0.030532f
C280 source.n108 a_n2354_n3288# 0.016407f
C281 source.n109 a_n2354_n3288# 0.017372f
C282 source.n110 a_n2354_n3288# 0.038779f
C283 source.n111 a_n2354_n3288# 0.038779f
C284 source.n112 a_n2354_n3288# 0.017372f
C285 source.n113 a_n2354_n3288# 0.016407f
C286 source.n114 a_n2354_n3288# 0.030532f
C287 source.n115 a_n2354_n3288# 0.030532f
C288 source.n116 a_n2354_n3288# 0.016407f
C289 source.n117 a_n2354_n3288# 0.017372f
C290 source.n118 a_n2354_n3288# 0.038779f
C291 source.n119 a_n2354_n3288# 0.038779f
C292 source.n120 a_n2354_n3288# 0.038779f
C293 source.n121 a_n2354_n3288# 0.016889f
C294 source.n122 a_n2354_n3288# 0.016407f
C295 source.n123 a_n2354_n3288# 0.030532f
C296 source.n124 a_n2354_n3288# 0.030532f
C297 source.n125 a_n2354_n3288# 0.016407f
C298 source.n126 a_n2354_n3288# 0.017372f
C299 source.n127 a_n2354_n3288# 0.038779f
C300 source.n128 a_n2354_n3288# 0.038779f
C301 source.n129 a_n2354_n3288# 0.017372f
C302 source.n130 a_n2354_n3288# 0.016407f
C303 source.n131 a_n2354_n3288# 0.030532f
C304 source.n132 a_n2354_n3288# 0.030532f
C305 source.n133 a_n2354_n3288# 0.016407f
C306 source.n134 a_n2354_n3288# 0.017372f
C307 source.n135 a_n2354_n3288# 0.038779f
C308 source.n136 a_n2354_n3288# 0.079579f
C309 source.n137 a_n2354_n3288# 0.017372f
C310 source.n138 a_n2354_n3288# 0.016407f
C311 source.n139 a_n2354_n3288# 0.065568f
C312 source.n140 a_n2354_n3288# 0.043919f
C313 source.n141 a_n2354_n3288# 0.12291f
C314 source.n142 a_n2354_n3288# 0.040444f
C315 source.n143 a_n2354_n3288# 0.030532f
C316 source.n144 a_n2354_n3288# 0.016407f
C317 source.n145 a_n2354_n3288# 0.038779f
C318 source.n146 a_n2354_n3288# 0.017372f
C319 source.n147 a_n2354_n3288# 0.030532f
C320 source.n148 a_n2354_n3288# 0.016407f
C321 source.n149 a_n2354_n3288# 0.038779f
C322 source.n150 a_n2354_n3288# 0.017372f
C323 source.n151 a_n2354_n3288# 0.030532f
C324 source.n152 a_n2354_n3288# 0.016889f
C325 source.n153 a_n2354_n3288# 0.038779f
C326 source.n154 a_n2354_n3288# 0.016407f
C327 source.n155 a_n2354_n3288# 0.017372f
C328 source.n156 a_n2354_n3288# 0.030532f
C329 source.n157 a_n2354_n3288# 0.016407f
C330 source.n158 a_n2354_n3288# 0.038779f
C331 source.n159 a_n2354_n3288# 0.017372f
C332 source.n160 a_n2354_n3288# 0.030532f
C333 source.n161 a_n2354_n3288# 0.016407f
C334 source.n162 a_n2354_n3288# 0.029084f
C335 source.n163 a_n2354_n3288# 0.027414f
C336 source.t8 a_n2354_n3288# 0.065495f
C337 source.n164 a_n2354_n3288# 0.220132f
C338 source.n165 a_n2354_n3288# 1.54029f
C339 source.n166 a_n2354_n3288# 0.016407f
C340 source.n167 a_n2354_n3288# 0.017372f
C341 source.n168 a_n2354_n3288# 0.038779f
C342 source.n169 a_n2354_n3288# 0.038779f
C343 source.n170 a_n2354_n3288# 0.017372f
C344 source.n171 a_n2354_n3288# 0.016407f
C345 source.n172 a_n2354_n3288# 0.030532f
C346 source.n173 a_n2354_n3288# 0.030532f
C347 source.n174 a_n2354_n3288# 0.016407f
C348 source.n175 a_n2354_n3288# 0.017372f
C349 source.n176 a_n2354_n3288# 0.038779f
C350 source.n177 a_n2354_n3288# 0.038779f
C351 source.n178 a_n2354_n3288# 0.017372f
C352 source.n179 a_n2354_n3288# 0.016407f
C353 source.n180 a_n2354_n3288# 0.030532f
C354 source.n181 a_n2354_n3288# 0.030532f
C355 source.n182 a_n2354_n3288# 0.016407f
C356 source.n183 a_n2354_n3288# 0.017372f
C357 source.n184 a_n2354_n3288# 0.038779f
C358 source.n185 a_n2354_n3288# 0.038779f
C359 source.n186 a_n2354_n3288# 0.038779f
C360 source.n187 a_n2354_n3288# 0.016889f
C361 source.n188 a_n2354_n3288# 0.016407f
C362 source.n189 a_n2354_n3288# 0.030532f
C363 source.n190 a_n2354_n3288# 0.030532f
C364 source.n191 a_n2354_n3288# 0.016407f
C365 source.n192 a_n2354_n3288# 0.017372f
C366 source.n193 a_n2354_n3288# 0.038779f
C367 source.n194 a_n2354_n3288# 0.038779f
C368 source.n195 a_n2354_n3288# 0.017372f
C369 source.n196 a_n2354_n3288# 0.016407f
C370 source.n197 a_n2354_n3288# 0.030532f
C371 source.n198 a_n2354_n3288# 0.030532f
C372 source.n199 a_n2354_n3288# 0.016407f
C373 source.n200 a_n2354_n3288# 0.017372f
C374 source.n201 a_n2354_n3288# 0.038779f
C375 source.n202 a_n2354_n3288# 0.079579f
C376 source.n203 a_n2354_n3288# 0.017372f
C377 source.n204 a_n2354_n3288# 0.016407f
C378 source.n205 a_n2354_n3288# 0.065568f
C379 source.n206 a_n2354_n3288# 0.043919f
C380 source.n207 a_n2354_n3288# 0.12291f
C381 source.t19 a_n2354_n3288# 0.289528f
C382 source.t2 a_n2354_n3288# 0.289528f
C383 source.n208 a_n2354_n3288# 2.47894f
C384 source.n209 a_n2354_n3288# 0.419013f
C385 source.t17 a_n2354_n3288# 0.289528f
C386 source.t1 a_n2354_n3288# 0.289528f
C387 source.n210 a_n2354_n3288# 2.47894f
C388 source.n211 a_n2354_n3288# 0.419013f
C389 source.t0 a_n2354_n3288# 0.289528f
C390 source.t10 a_n2354_n3288# 0.289528f
C391 source.n212 a_n2354_n3288# 2.47894f
C392 source.n213 a_n2354_n3288# 0.419013f
C393 source.t23 a_n2354_n3288# 0.289528f
C394 source.t7 a_n2354_n3288# 0.289528f
C395 source.n214 a_n2354_n3288# 2.47894f
C396 source.n215 a_n2354_n3288# 0.419013f
C397 source.t22 a_n2354_n3288# 0.289528f
C398 source.t20 a_n2354_n3288# 0.289528f
C399 source.n216 a_n2354_n3288# 2.47894f
C400 source.n217 a_n2354_n3288# 0.419013f
C401 source.n218 a_n2354_n3288# 0.040444f
C402 source.n219 a_n2354_n3288# 0.030532f
C403 source.n220 a_n2354_n3288# 0.016407f
C404 source.n221 a_n2354_n3288# 0.038779f
C405 source.n222 a_n2354_n3288# 0.017372f
C406 source.n223 a_n2354_n3288# 0.030532f
C407 source.n224 a_n2354_n3288# 0.016407f
C408 source.n225 a_n2354_n3288# 0.038779f
C409 source.n226 a_n2354_n3288# 0.017372f
C410 source.n227 a_n2354_n3288# 0.030532f
C411 source.n228 a_n2354_n3288# 0.016889f
C412 source.n229 a_n2354_n3288# 0.038779f
C413 source.n230 a_n2354_n3288# 0.016407f
C414 source.n231 a_n2354_n3288# 0.017372f
C415 source.n232 a_n2354_n3288# 0.030532f
C416 source.n233 a_n2354_n3288# 0.016407f
C417 source.n234 a_n2354_n3288# 0.038779f
C418 source.n235 a_n2354_n3288# 0.017372f
C419 source.n236 a_n2354_n3288# 0.030532f
C420 source.n237 a_n2354_n3288# 0.016407f
C421 source.n238 a_n2354_n3288# 0.029084f
C422 source.n239 a_n2354_n3288# 0.027414f
C423 source.t13 a_n2354_n3288# 0.065495f
C424 source.n240 a_n2354_n3288# 0.220132f
C425 source.n241 a_n2354_n3288# 1.54029f
C426 source.n242 a_n2354_n3288# 0.016407f
C427 source.n243 a_n2354_n3288# 0.017372f
C428 source.n244 a_n2354_n3288# 0.038779f
C429 source.n245 a_n2354_n3288# 0.038779f
C430 source.n246 a_n2354_n3288# 0.017372f
C431 source.n247 a_n2354_n3288# 0.016407f
C432 source.n248 a_n2354_n3288# 0.030532f
C433 source.n249 a_n2354_n3288# 0.030532f
C434 source.n250 a_n2354_n3288# 0.016407f
C435 source.n251 a_n2354_n3288# 0.017372f
C436 source.n252 a_n2354_n3288# 0.038779f
C437 source.n253 a_n2354_n3288# 0.038779f
C438 source.n254 a_n2354_n3288# 0.017372f
C439 source.n255 a_n2354_n3288# 0.016407f
C440 source.n256 a_n2354_n3288# 0.030532f
C441 source.n257 a_n2354_n3288# 0.030532f
C442 source.n258 a_n2354_n3288# 0.016407f
C443 source.n259 a_n2354_n3288# 0.017372f
C444 source.n260 a_n2354_n3288# 0.038779f
C445 source.n261 a_n2354_n3288# 0.038779f
C446 source.n262 a_n2354_n3288# 0.038779f
C447 source.n263 a_n2354_n3288# 0.016889f
C448 source.n264 a_n2354_n3288# 0.016407f
C449 source.n265 a_n2354_n3288# 0.030532f
C450 source.n266 a_n2354_n3288# 0.030532f
C451 source.n267 a_n2354_n3288# 0.016407f
C452 source.n268 a_n2354_n3288# 0.017372f
C453 source.n269 a_n2354_n3288# 0.038779f
C454 source.n270 a_n2354_n3288# 0.038779f
C455 source.n271 a_n2354_n3288# 0.017372f
C456 source.n272 a_n2354_n3288# 0.016407f
C457 source.n273 a_n2354_n3288# 0.030532f
C458 source.n274 a_n2354_n3288# 0.030532f
C459 source.n275 a_n2354_n3288# 0.016407f
C460 source.n276 a_n2354_n3288# 0.017372f
C461 source.n277 a_n2354_n3288# 0.038779f
C462 source.n278 a_n2354_n3288# 0.079579f
C463 source.n279 a_n2354_n3288# 0.017372f
C464 source.n280 a_n2354_n3288# 0.016407f
C465 source.n281 a_n2354_n3288# 0.065568f
C466 source.n282 a_n2354_n3288# 0.043919f
C467 source.n283 a_n2354_n3288# 1.70885f
C468 source.n284 a_n2354_n3288# 0.040444f
C469 source.n285 a_n2354_n3288# 0.030532f
C470 source.n286 a_n2354_n3288# 0.016407f
C471 source.n287 a_n2354_n3288# 0.038779f
C472 source.n288 a_n2354_n3288# 0.017372f
C473 source.n289 a_n2354_n3288# 0.030532f
C474 source.n290 a_n2354_n3288# 0.016407f
C475 source.n291 a_n2354_n3288# 0.038779f
C476 source.n292 a_n2354_n3288# 0.017372f
C477 source.n293 a_n2354_n3288# 0.030532f
C478 source.n294 a_n2354_n3288# 0.016889f
C479 source.n295 a_n2354_n3288# 0.038779f
C480 source.n296 a_n2354_n3288# 0.017372f
C481 source.n297 a_n2354_n3288# 0.030532f
C482 source.n298 a_n2354_n3288# 0.016407f
C483 source.n299 a_n2354_n3288# 0.038779f
C484 source.n300 a_n2354_n3288# 0.017372f
C485 source.n301 a_n2354_n3288# 0.030532f
C486 source.n302 a_n2354_n3288# 0.016407f
C487 source.n303 a_n2354_n3288# 0.029084f
C488 source.n304 a_n2354_n3288# 0.027414f
C489 source.t44 a_n2354_n3288# 0.065495f
C490 source.n305 a_n2354_n3288# 0.220132f
C491 source.n306 a_n2354_n3288# 1.54029f
C492 source.n307 a_n2354_n3288# 0.016407f
C493 source.n308 a_n2354_n3288# 0.017372f
C494 source.n309 a_n2354_n3288# 0.038779f
C495 source.n310 a_n2354_n3288# 0.038779f
C496 source.n311 a_n2354_n3288# 0.017372f
C497 source.n312 a_n2354_n3288# 0.016407f
C498 source.n313 a_n2354_n3288# 0.030532f
C499 source.n314 a_n2354_n3288# 0.030532f
C500 source.n315 a_n2354_n3288# 0.016407f
C501 source.n316 a_n2354_n3288# 0.017372f
C502 source.n317 a_n2354_n3288# 0.038779f
C503 source.n318 a_n2354_n3288# 0.038779f
C504 source.n319 a_n2354_n3288# 0.017372f
C505 source.n320 a_n2354_n3288# 0.016407f
C506 source.n321 a_n2354_n3288# 0.030532f
C507 source.n322 a_n2354_n3288# 0.030532f
C508 source.n323 a_n2354_n3288# 0.016407f
C509 source.n324 a_n2354_n3288# 0.016407f
C510 source.n325 a_n2354_n3288# 0.017372f
C511 source.n326 a_n2354_n3288# 0.038779f
C512 source.n327 a_n2354_n3288# 0.038779f
C513 source.n328 a_n2354_n3288# 0.038779f
C514 source.n329 a_n2354_n3288# 0.016889f
C515 source.n330 a_n2354_n3288# 0.016407f
C516 source.n331 a_n2354_n3288# 0.030532f
C517 source.n332 a_n2354_n3288# 0.030532f
C518 source.n333 a_n2354_n3288# 0.016407f
C519 source.n334 a_n2354_n3288# 0.017372f
C520 source.n335 a_n2354_n3288# 0.038779f
C521 source.n336 a_n2354_n3288# 0.038779f
C522 source.n337 a_n2354_n3288# 0.017372f
C523 source.n338 a_n2354_n3288# 0.016407f
C524 source.n339 a_n2354_n3288# 0.030532f
C525 source.n340 a_n2354_n3288# 0.030532f
C526 source.n341 a_n2354_n3288# 0.016407f
C527 source.n342 a_n2354_n3288# 0.017372f
C528 source.n343 a_n2354_n3288# 0.038779f
C529 source.n344 a_n2354_n3288# 0.079579f
C530 source.n345 a_n2354_n3288# 0.017372f
C531 source.n346 a_n2354_n3288# 0.016407f
C532 source.n347 a_n2354_n3288# 0.065568f
C533 source.n348 a_n2354_n3288# 0.043919f
C534 source.n349 a_n2354_n3288# 1.70885f
C535 source.t38 a_n2354_n3288# 0.289528f
C536 source.t29 a_n2354_n3288# 0.289528f
C537 source.n350 a_n2354_n3288# 2.47893f
C538 source.n351 a_n2354_n3288# 0.419028f
C539 source.t45 a_n2354_n3288# 0.289528f
C540 source.t30 a_n2354_n3288# 0.289528f
C541 source.n352 a_n2354_n3288# 2.47893f
C542 source.n353 a_n2354_n3288# 0.419028f
C543 source.t41 a_n2354_n3288# 0.289528f
C544 source.t34 a_n2354_n3288# 0.289528f
C545 source.n354 a_n2354_n3288# 2.47893f
C546 source.n355 a_n2354_n3288# 0.419028f
C547 source.t43 a_n2354_n3288# 0.289528f
C548 source.t35 a_n2354_n3288# 0.289528f
C549 source.n356 a_n2354_n3288# 2.47893f
C550 source.n357 a_n2354_n3288# 0.419028f
C551 source.t26 a_n2354_n3288# 0.289528f
C552 source.t37 a_n2354_n3288# 0.289528f
C553 source.n358 a_n2354_n3288# 2.47893f
C554 source.n359 a_n2354_n3288# 0.419028f
C555 source.n360 a_n2354_n3288# 0.040444f
C556 source.n361 a_n2354_n3288# 0.030532f
C557 source.n362 a_n2354_n3288# 0.016407f
C558 source.n363 a_n2354_n3288# 0.038779f
C559 source.n364 a_n2354_n3288# 0.017372f
C560 source.n365 a_n2354_n3288# 0.030532f
C561 source.n366 a_n2354_n3288# 0.016407f
C562 source.n367 a_n2354_n3288# 0.038779f
C563 source.n368 a_n2354_n3288# 0.017372f
C564 source.n369 a_n2354_n3288# 0.030532f
C565 source.n370 a_n2354_n3288# 0.016889f
C566 source.n371 a_n2354_n3288# 0.038779f
C567 source.n372 a_n2354_n3288# 0.017372f
C568 source.n373 a_n2354_n3288# 0.030532f
C569 source.n374 a_n2354_n3288# 0.016407f
C570 source.n375 a_n2354_n3288# 0.038779f
C571 source.n376 a_n2354_n3288# 0.017372f
C572 source.n377 a_n2354_n3288# 0.030532f
C573 source.n378 a_n2354_n3288# 0.016407f
C574 source.n379 a_n2354_n3288# 0.029084f
C575 source.n380 a_n2354_n3288# 0.027414f
C576 source.t27 a_n2354_n3288# 0.065495f
C577 source.n381 a_n2354_n3288# 0.220132f
C578 source.n382 a_n2354_n3288# 1.54029f
C579 source.n383 a_n2354_n3288# 0.016407f
C580 source.n384 a_n2354_n3288# 0.017372f
C581 source.n385 a_n2354_n3288# 0.038779f
C582 source.n386 a_n2354_n3288# 0.038779f
C583 source.n387 a_n2354_n3288# 0.017372f
C584 source.n388 a_n2354_n3288# 0.016407f
C585 source.n389 a_n2354_n3288# 0.030532f
C586 source.n390 a_n2354_n3288# 0.030532f
C587 source.n391 a_n2354_n3288# 0.016407f
C588 source.n392 a_n2354_n3288# 0.017372f
C589 source.n393 a_n2354_n3288# 0.038779f
C590 source.n394 a_n2354_n3288# 0.038779f
C591 source.n395 a_n2354_n3288# 0.017372f
C592 source.n396 a_n2354_n3288# 0.016407f
C593 source.n397 a_n2354_n3288# 0.030532f
C594 source.n398 a_n2354_n3288# 0.030532f
C595 source.n399 a_n2354_n3288# 0.016407f
C596 source.n400 a_n2354_n3288# 0.016407f
C597 source.n401 a_n2354_n3288# 0.017372f
C598 source.n402 a_n2354_n3288# 0.038779f
C599 source.n403 a_n2354_n3288# 0.038779f
C600 source.n404 a_n2354_n3288# 0.038779f
C601 source.n405 a_n2354_n3288# 0.016889f
C602 source.n406 a_n2354_n3288# 0.016407f
C603 source.n407 a_n2354_n3288# 0.030532f
C604 source.n408 a_n2354_n3288# 0.030532f
C605 source.n409 a_n2354_n3288# 0.016407f
C606 source.n410 a_n2354_n3288# 0.017372f
C607 source.n411 a_n2354_n3288# 0.038779f
C608 source.n412 a_n2354_n3288# 0.038779f
C609 source.n413 a_n2354_n3288# 0.017372f
C610 source.n414 a_n2354_n3288# 0.016407f
C611 source.n415 a_n2354_n3288# 0.030532f
C612 source.n416 a_n2354_n3288# 0.030532f
C613 source.n417 a_n2354_n3288# 0.016407f
C614 source.n418 a_n2354_n3288# 0.017372f
C615 source.n419 a_n2354_n3288# 0.038779f
C616 source.n420 a_n2354_n3288# 0.079579f
C617 source.n421 a_n2354_n3288# 0.017372f
C618 source.n422 a_n2354_n3288# 0.016407f
C619 source.n423 a_n2354_n3288# 0.065568f
C620 source.n424 a_n2354_n3288# 0.043919f
C621 source.n425 a_n2354_n3288# 0.12291f
C622 source.n426 a_n2354_n3288# 0.040444f
C623 source.n427 a_n2354_n3288# 0.030532f
C624 source.n428 a_n2354_n3288# 0.016407f
C625 source.n429 a_n2354_n3288# 0.038779f
C626 source.n430 a_n2354_n3288# 0.017372f
C627 source.n431 a_n2354_n3288# 0.030532f
C628 source.n432 a_n2354_n3288# 0.016407f
C629 source.n433 a_n2354_n3288# 0.038779f
C630 source.n434 a_n2354_n3288# 0.017372f
C631 source.n435 a_n2354_n3288# 0.030532f
C632 source.n436 a_n2354_n3288# 0.016889f
C633 source.n437 a_n2354_n3288# 0.038779f
C634 source.n438 a_n2354_n3288# 0.017372f
C635 source.n439 a_n2354_n3288# 0.030532f
C636 source.n440 a_n2354_n3288# 0.016407f
C637 source.n441 a_n2354_n3288# 0.038779f
C638 source.n442 a_n2354_n3288# 0.017372f
C639 source.n443 a_n2354_n3288# 0.030532f
C640 source.n444 a_n2354_n3288# 0.016407f
C641 source.n445 a_n2354_n3288# 0.029084f
C642 source.n446 a_n2354_n3288# 0.027414f
C643 source.t4 a_n2354_n3288# 0.065495f
C644 source.n447 a_n2354_n3288# 0.220132f
C645 source.n448 a_n2354_n3288# 1.54029f
C646 source.n449 a_n2354_n3288# 0.016407f
C647 source.n450 a_n2354_n3288# 0.017372f
C648 source.n451 a_n2354_n3288# 0.038779f
C649 source.n452 a_n2354_n3288# 0.038779f
C650 source.n453 a_n2354_n3288# 0.017372f
C651 source.n454 a_n2354_n3288# 0.016407f
C652 source.n455 a_n2354_n3288# 0.030532f
C653 source.n456 a_n2354_n3288# 0.030532f
C654 source.n457 a_n2354_n3288# 0.016407f
C655 source.n458 a_n2354_n3288# 0.017372f
C656 source.n459 a_n2354_n3288# 0.038779f
C657 source.n460 a_n2354_n3288# 0.038779f
C658 source.n461 a_n2354_n3288# 0.017372f
C659 source.n462 a_n2354_n3288# 0.016407f
C660 source.n463 a_n2354_n3288# 0.030532f
C661 source.n464 a_n2354_n3288# 0.030532f
C662 source.n465 a_n2354_n3288# 0.016407f
C663 source.n466 a_n2354_n3288# 0.016407f
C664 source.n467 a_n2354_n3288# 0.017372f
C665 source.n468 a_n2354_n3288# 0.038779f
C666 source.n469 a_n2354_n3288# 0.038779f
C667 source.n470 a_n2354_n3288# 0.038779f
C668 source.n471 a_n2354_n3288# 0.016889f
C669 source.n472 a_n2354_n3288# 0.016407f
C670 source.n473 a_n2354_n3288# 0.030532f
C671 source.n474 a_n2354_n3288# 0.030532f
C672 source.n475 a_n2354_n3288# 0.016407f
C673 source.n476 a_n2354_n3288# 0.017372f
C674 source.n477 a_n2354_n3288# 0.038779f
C675 source.n478 a_n2354_n3288# 0.038779f
C676 source.n479 a_n2354_n3288# 0.017372f
C677 source.n480 a_n2354_n3288# 0.016407f
C678 source.n481 a_n2354_n3288# 0.030532f
C679 source.n482 a_n2354_n3288# 0.030532f
C680 source.n483 a_n2354_n3288# 0.016407f
C681 source.n484 a_n2354_n3288# 0.017372f
C682 source.n485 a_n2354_n3288# 0.038779f
C683 source.n486 a_n2354_n3288# 0.079579f
C684 source.n487 a_n2354_n3288# 0.017372f
C685 source.n488 a_n2354_n3288# 0.016407f
C686 source.n489 a_n2354_n3288# 0.065568f
C687 source.n490 a_n2354_n3288# 0.043919f
C688 source.n491 a_n2354_n3288# 0.12291f
C689 source.t15 a_n2354_n3288# 0.289528f
C690 source.t9 a_n2354_n3288# 0.289528f
C691 source.n492 a_n2354_n3288# 2.47893f
C692 source.n493 a_n2354_n3288# 0.419028f
C693 source.t11 a_n2354_n3288# 0.289528f
C694 source.t16 a_n2354_n3288# 0.289528f
C695 source.n494 a_n2354_n3288# 2.47893f
C696 source.n495 a_n2354_n3288# 0.419028f
C697 source.t18 a_n2354_n3288# 0.289528f
C698 source.t12 a_n2354_n3288# 0.289528f
C699 source.n496 a_n2354_n3288# 2.47893f
C700 source.n497 a_n2354_n3288# 0.419028f
C701 source.t3 a_n2354_n3288# 0.289528f
C702 source.t5 a_n2354_n3288# 0.289528f
C703 source.n498 a_n2354_n3288# 2.47893f
C704 source.n499 a_n2354_n3288# 0.419028f
C705 source.t6 a_n2354_n3288# 0.289528f
C706 source.t21 a_n2354_n3288# 0.289528f
C707 source.n500 a_n2354_n3288# 2.47893f
C708 source.n501 a_n2354_n3288# 0.419028f
C709 source.n502 a_n2354_n3288# 0.040444f
C710 source.n503 a_n2354_n3288# 0.030532f
C711 source.n504 a_n2354_n3288# 0.016407f
C712 source.n505 a_n2354_n3288# 0.038779f
C713 source.n506 a_n2354_n3288# 0.017372f
C714 source.n507 a_n2354_n3288# 0.030532f
C715 source.n508 a_n2354_n3288# 0.016407f
C716 source.n509 a_n2354_n3288# 0.038779f
C717 source.n510 a_n2354_n3288# 0.017372f
C718 source.n511 a_n2354_n3288# 0.030532f
C719 source.n512 a_n2354_n3288# 0.016889f
C720 source.n513 a_n2354_n3288# 0.038779f
C721 source.n514 a_n2354_n3288# 0.017372f
C722 source.n515 a_n2354_n3288# 0.030532f
C723 source.n516 a_n2354_n3288# 0.016407f
C724 source.n517 a_n2354_n3288# 0.038779f
C725 source.n518 a_n2354_n3288# 0.017372f
C726 source.n519 a_n2354_n3288# 0.030532f
C727 source.n520 a_n2354_n3288# 0.016407f
C728 source.n521 a_n2354_n3288# 0.029084f
C729 source.n522 a_n2354_n3288# 0.027414f
C730 source.t14 a_n2354_n3288# 0.065495f
C731 source.n523 a_n2354_n3288# 0.220132f
C732 source.n524 a_n2354_n3288# 1.54029f
C733 source.n525 a_n2354_n3288# 0.016407f
C734 source.n526 a_n2354_n3288# 0.017372f
C735 source.n527 a_n2354_n3288# 0.038779f
C736 source.n528 a_n2354_n3288# 0.038779f
C737 source.n529 a_n2354_n3288# 0.017372f
C738 source.n530 a_n2354_n3288# 0.016407f
C739 source.n531 a_n2354_n3288# 0.030532f
C740 source.n532 a_n2354_n3288# 0.030532f
C741 source.n533 a_n2354_n3288# 0.016407f
C742 source.n534 a_n2354_n3288# 0.017372f
C743 source.n535 a_n2354_n3288# 0.038779f
C744 source.n536 a_n2354_n3288# 0.038779f
C745 source.n537 a_n2354_n3288# 0.017372f
C746 source.n538 a_n2354_n3288# 0.016407f
C747 source.n539 a_n2354_n3288# 0.030532f
C748 source.n540 a_n2354_n3288# 0.030532f
C749 source.n541 a_n2354_n3288# 0.016407f
C750 source.n542 a_n2354_n3288# 0.016407f
C751 source.n543 a_n2354_n3288# 0.017372f
C752 source.n544 a_n2354_n3288# 0.038779f
C753 source.n545 a_n2354_n3288# 0.038779f
C754 source.n546 a_n2354_n3288# 0.038779f
C755 source.n547 a_n2354_n3288# 0.016889f
C756 source.n548 a_n2354_n3288# 0.016407f
C757 source.n549 a_n2354_n3288# 0.030532f
C758 source.n550 a_n2354_n3288# 0.030532f
C759 source.n551 a_n2354_n3288# 0.016407f
C760 source.n552 a_n2354_n3288# 0.017372f
C761 source.n553 a_n2354_n3288# 0.038779f
C762 source.n554 a_n2354_n3288# 0.038779f
C763 source.n555 a_n2354_n3288# 0.017372f
C764 source.n556 a_n2354_n3288# 0.016407f
C765 source.n557 a_n2354_n3288# 0.030532f
C766 source.n558 a_n2354_n3288# 0.030532f
C767 source.n559 a_n2354_n3288# 0.016407f
C768 source.n560 a_n2354_n3288# 0.017372f
C769 source.n561 a_n2354_n3288# 0.038779f
C770 source.n562 a_n2354_n3288# 0.079579f
C771 source.n563 a_n2354_n3288# 0.017372f
C772 source.n564 a_n2354_n3288# 0.016407f
C773 source.n565 a_n2354_n3288# 0.065568f
C774 source.n566 a_n2354_n3288# 0.043919f
C775 source.n567 a_n2354_n3288# 0.295263f
C776 source.n568 a_n2354_n3288# 1.91539f
C777 drain_left.t6 a_n2354_n3288# 0.325142f
C778 drain_left.t10 a_n2354_n3288# 0.325142f
C779 drain_left.n0 a_n2354_n3288# 2.89707f
C780 drain_left.t5 a_n2354_n3288# 0.325142f
C781 drain_left.t7 a_n2354_n3288# 0.325142f
C782 drain_left.n1 a_n2354_n3288# 2.89326f
C783 drain_left.n2 a_n2354_n3288# 0.825538f
C784 drain_left.t16 a_n2354_n3288# 0.325142f
C785 drain_left.t9 a_n2354_n3288# 0.325142f
C786 drain_left.n3 a_n2354_n3288# 2.89326f
C787 drain_left.n4 a_n2354_n3288# 0.375329f
C788 drain_left.t15 a_n2354_n3288# 0.325142f
C789 drain_left.t23 a_n2354_n3288# 0.325142f
C790 drain_left.n5 a_n2354_n3288# 2.89707f
C791 drain_left.t19 a_n2354_n3288# 0.325142f
C792 drain_left.t22 a_n2354_n3288# 0.325142f
C793 drain_left.n6 a_n2354_n3288# 2.89326f
C794 drain_left.n7 a_n2354_n3288# 0.825538f
C795 drain_left.t18 a_n2354_n3288# 0.325142f
C796 drain_left.t3 a_n2354_n3288# 0.325142f
C797 drain_left.n8 a_n2354_n3288# 2.89326f
C798 drain_left.n9 a_n2354_n3288# 0.375329f
C799 drain_left.n10 a_n2354_n3288# 1.8602f
C800 drain_left.t2 a_n2354_n3288# 0.325142f
C801 drain_left.t14 a_n2354_n3288# 0.325142f
C802 drain_left.n11 a_n2354_n3288# 2.89709f
C803 drain_left.t17 a_n2354_n3288# 0.325142f
C804 drain_left.t20 a_n2354_n3288# 0.325142f
C805 drain_left.n12 a_n2354_n3288# 2.89328f
C806 drain_left.n13 a_n2354_n3288# 0.825514f
C807 drain_left.t11 a_n2354_n3288# 0.325142f
C808 drain_left.t12 a_n2354_n3288# 0.325142f
C809 drain_left.n14 a_n2354_n3288# 2.89328f
C810 drain_left.n15 a_n2354_n3288# 0.407757f
C811 drain_left.t21 a_n2354_n3288# 0.325142f
C812 drain_left.t0 a_n2354_n3288# 0.325142f
C813 drain_left.n16 a_n2354_n3288# 2.89328f
C814 drain_left.n17 a_n2354_n3288# 0.407757f
C815 drain_left.t13 a_n2354_n3288# 0.325142f
C816 drain_left.t4 a_n2354_n3288# 0.325142f
C817 drain_left.n18 a_n2354_n3288# 2.89328f
C818 drain_left.n19 a_n2354_n3288# 0.407757f
C819 drain_left.t1 a_n2354_n3288# 0.325142f
C820 drain_left.t8 a_n2354_n3288# 0.325142f
C821 drain_left.n20 a_n2354_n3288# 2.89326f
C822 drain_left.n21 a_n2354_n3288# 0.693166f
C823 plus.n0 a_n2354_n3288# 0.049398f
C824 plus.t0 a_n2354_n3288# 0.502526f
C825 plus.t19 a_n2354_n3288# 0.502526f
C826 plus.n1 a_n2354_n3288# 0.199349f
C827 plus.n2 a_n2354_n3288# 0.049398f
C828 plus.t14 a_n2354_n3288# 0.502526f
C829 plus.t1 a_n2354_n3288# 0.502526f
C830 plus.t22 a_n2354_n3288# 0.502526f
C831 plus.n3 a_n2354_n3288# 0.199349f
C832 plus.n4 a_n2354_n3288# 0.049398f
C833 plus.t15 a_n2354_n3288# 0.502526f
C834 plus.t8 a_n2354_n3288# 0.502526f
C835 plus.n5 a_n2354_n3288# 0.199349f
C836 plus.n6 a_n2354_n3288# 0.049398f
C837 plus.t23 a_n2354_n3288# 0.502526f
C838 plus.t16 a_n2354_n3288# 0.502526f
C839 plus.n7 a_n2354_n3288# 0.018976f
C840 plus.t5 a_n2354_n3288# 0.508231f
C841 plus.t11 a_n2354_n3288# 0.502526f
C842 plus.n8 a_n2354_n3288# 0.199349f
C843 plus.n9 a_n2354_n3288# 0.214513f
C844 plus.n10 a_n2354_n3288# 0.105735f
C845 plus.n11 a_n2354_n3288# 0.049398f
C846 plus.n12 a_n2354_n3288# 0.017757f
C847 plus.n13 a_n2354_n3288# 0.199349f
C848 plus.n14 a_n2354_n3288# 0.020346f
C849 plus.n15 a_n2354_n3288# 0.199349f
C850 plus.n16 a_n2354_n3288# 0.020346f
C851 plus.n17 a_n2354_n3288# 0.049398f
C852 plus.n18 a_n2354_n3288# 0.049398f
C853 plus.n19 a_n2354_n3288# 0.020346f
C854 plus.n20 a_n2354_n3288# 0.199349f
C855 plus.n21 a_n2354_n3288# 0.018367f
C856 plus.n22 a_n2354_n3288# 0.018367f
C857 plus.n23 a_n2354_n3288# 0.049398f
C858 plus.n24 a_n2354_n3288# 0.049398f
C859 plus.n25 a_n2354_n3288# 0.020346f
C860 plus.n26 a_n2354_n3288# 0.199349f
C861 plus.n27 a_n2354_n3288# 0.020346f
C862 plus.n28 a_n2354_n3288# 0.199349f
C863 plus.n29 a_n2354_n3288# 0.020346f
C864 plus.n30 a_n2354_n3288# 0.049398f
C865 plus.n31 a_n2354_n3288# 0.049398f
C866 plus.n32 a_n2354_n3288# 0.017757f
C867 plus.n33 a_n2354_n3288# 0.018976f
C868 plus.n34 a_n2354_n3288# 0.199349f
C869 plus.t7 a_n2354_n3288# 0.508231f
C870 plus.n35 a_n2354_n3288# 0.214447f
C871 plus.n36 a_n2354_n3288# 0.549168f
C872 plus.n37 a_n2354_n3288# 0.049398f
C873 plus.t3 a_n2354_n3288# 0.508231f
C874 plus.t9 a_n2354_n3288# 0.502526f
C875 plus.t18 a_n2354_n3288# 0.502526f
C876 plus.n38 a_n2354_n3288# 0.199349f
C877 plus.n39 a_n2354_n3288# 0.049398f
C878 plus.t2 a_n2354_n3288# 0.502526f
C879 plus.t17 a_n2354_n3288# 0.502526f
C880 plus.t6 a_n2354_n3288# 0.502526f
C881 plus.n40 a_n2354_n3288# 0.199349f
C882 plus.n41 a_n2354_n3288# 0.049398f
C883 plus.t13 a_n2354_n3288# 0.502526f
C884 plus.t4 a_n2354_n3288# 0.502526f
C885 plus.n42 a_n2354_n3288# 0.199349f
C886 plus.n43 a_n2354_n3288# 0.049398f
C887 plus.t12 a_n2354_n3288# 0.502526f
C888 plus.t21 a_n2354_n3288# 0.502526f
C889 plus.n44 a_n2354_n3288# 0.018976f
C890 plus.t10 a_n2354_n3288# 0.502526f
C891 plus.n45 a_n2354_n3288# 0.199349f
C892 plus.t20 a_n2354_n3288# 0.508231f
C893 plus.n46 a_n2354_n3288# 0.214513f
C894 plus.n47 a_n2354_n3288# 0.105735f
C895 plus.n48 a_n2354_n3288# 0.049398f
C896 plus.n49 a_n2354_n3288# 0.017757f
C897 plus.n50 a_n2354_n3288# 0.199349f
C898 plus.n51 a_n2354_n3288# 0.020346f
C899 plus.n52 a_n2354_n3288# 0.199349f
C900 plus.n53 a_n2354_n3288# 0.020346f
C901 plus.n54 a_n2354_n3288# 0.049398f
C902 plus.n55 a_n2354_n3288# 0.049398f
C903 plus.n56 a_n2354_n3288# 0.020346f
C904 plus.n57 a_n2354_n3288# 0.199349f
C905 plus.n58 a_n2354_n3288# 0.018367f
C906 plus.n59 a_n2354_n3288# 0.018367f
C907 plus.n60 a_n2354_n3288# 0.049398f
C908 plus.n61 a_n2354_n3288# 0.049398f
C909 plus.n62 a_n2354_n3288# 0.020346f
C910 plus.n63 a_n2354_n3288# 0.199349f
C911 plus.n64 a_n2354_n3288# 0.020346f
C912 plus.n65 a_n2354_n3288# 0.199349f
C913 plus.n66 a_n2354_n3288# 0.020346f
C914 plus.n67 a_n2354_n3288# 0.049398f
C915 plus.n68 a_n2354_n3288# 0.049398f
C916 plus.n69 a_n2354_n3288# 0.017757f
C917 plus.n70 a_n2354_n3288# 0.018976f
C918 plus.n71 a_n2354_n3288# 0.199349f
C919 plus.n72 a_n2354_n3288# 0.214447f
C920 plus.n73 a_n2354_n3288# 1.5981f
.ends

