* NGSPICE file created from diffpair611.ext - technology: sky130A

.subckt diffpair611 minus drain_right drain_left source plus
X0 drain_left plus source a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X1 a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X2 a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X3 drain_right minus source a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X4 a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X5 source plus drain_left a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X6 source minus drain_right a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X7 drain_right minus source a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X8 drain_left plus source a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X9 source plus drain_left a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X10 source minus drain_right a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X11 a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# a_n1274_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
.ends

