* NGSPICE file created from diffpair507.ext - technology: sky130A

.subckt diffpair507 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t24 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X1 drain_left.t14 plus.t1 source.t17 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X2 source.t21 plus.t2 drain_left.t13 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X3 drain_right.t15 minus.t0 source.t15 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X4 drain_left.t12 plus.t3 source.t27 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X5 source.t6 minus.t1 drain_right.t14 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X6 a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X7 drain_left.t11 plus.t4 source.t28 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X8 source.t14 minus.t2 drain_right.t13 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X9 source.t2 minus.t3 drain_right.t12 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X10 a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X11 source.t22 plus.t5 drain_left.t10 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X12 source.t31 plus.t6 drain_left.t9 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X13 source.t9 minus.t4 drain_right.t11 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X14 source.t12 minus.t5 drain_right.t10 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X15 drain_right.t9 minus.t6 source.t7 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X16 drain_left.t8 plus.t7 source.t25 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X17 source.t8 minus.t7 drain_right.t8 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X18 source.t18 plus.t8 drain_left.t7 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X19 source.t19 plus.t9 drain_left.t6 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X20 source.t23 plus.t10 drain_left.t5 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X21 a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X22 source.t20 plus.t11 drain_left.t4 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X23 drain_left.t3 plus.t12 source.t30 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X24 drain_right.t7 minus.t8 source.t11 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X25 drain_right.t6 minus.t9 source.t0 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X26 a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X27 drain_right.t5 minus.t10 source.t13 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X28 drain_right.t4 minus.t11 source.t4 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X29 drain_right.t3 minus.t12 source.t1 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X30 drain_right.t2 minus.t13 source.t3 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X31 drain_left.t2 plus.t13 source.t29 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X32 source.t16 plus.t14 drain_left.t1 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X33 drain_left.t0 plus.t15 source.t26 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X34 source.t5 minus.t14 drain_right.t1 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X35 source.t10 minus.t15 drain_right.t0 a_n1760_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
R0 plus.n4 plus.t6 1612.22
R1 plus.n19 plus.t4 1612.22
R2 plus.n25 plus.t3 1612.22
R3 plus.n40 plus.t11 1612.22
R4 plus.n5 plus.t1 1571.32
R5 plus.n3 plus.t10 1571.32
R6 plus.n10 plus.t0 1571.32
R7 plus.n1 plus.t9 1571.32
R8 plus.n16 plus.t15 1571.32
R9 plus.n18 plus.t8 1571.32
R10 plus.n26 plus.t14 1571.32
R11 plus.n24 plus.t12 1571.32
R12 plus.n31 plus.t5 1571.32
R13 plus.n22 plus.t7 1571.32
R14 plus.n37 plus.t2 1571.32
R15 plus.n39 plus.t13 1571.32
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus plus.n41 30.7717
R47 plus.n6 plus.n5 29.2126
R48 plus.n18 plus.n17 29.2126
R49 plus.n39 plus.n38 29.2126
R50 plus.n27 plus.n26 29.2126
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 13.2467
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n7 source.t31 45.521
R73 source.n8 source.t0 45.521
R74 source.n15 source.t9 45.521
R75 source.n31 source.t3 45.5208
R76 source.n24 source.t2 45.5208
R77 source.n23 source.t27 45.5208
R78 source.n16 source.t20 45.5208
R79 source.n0 source.t28 45.5208
R80 source.n2 source.n1 44.201
R81 source.n4 source.n3 44.201
R82 source.n6 source.n5 44.201
R83 source.n10 source.n9 44.201
R84 source.n12 source.n11 44.201
R85 source.n14 source.n13 44.201
R86 source.n30 source.n29 44.2008
R87 source.n28 source.n27 44.2008
R88 source.n26 source.n25 44.2008
R89 source.n22 source.n21 44.2008
R90 source.n20 source.n19 44.2008
R91 source.n18 source.n17 44.2008
R92 source.n16 source.n15 24.0605
R93 source.n32 source.n0 18.5475
R94 source.n32 source.n31 5.51343
R95 source.n29 source.t15 1.3205
R96 source.n29 source.t5 1.3205
R97 source.n27 source.t13 1.3205
R98 source.n27 source.t8 1.3205
R99 source.n25 source.t7 1.3205
R100 source.n25 source.t10 1.3205
R101 source.n21 source.t30 1.3205
R102 source.n21 source.t16 1.3205
R103 source.n19 source.t25 1.3205
R104 source.n19 source.t22 1.3205
R105 source.n17 source.t29 1.3205
R106 source.n17 source.t21 1.3205
R107 source.n1 source.t26 1.3205
R108 source.n1 source.t18 1.3205
R109 source.n3 source.t24 1.3205
R110 source.n3 source.t19 1.3205
R111 source.n5 source.t17 1.3205
R112 source.n5 source.t23 1.3205
R113 source.n9 source.t11 1.3205
R114 source.n9 source.t14 1.3205
R115 source.n11 source.t4 1.3205
R116 source.n11 source.t6 1.3205
R117 source.n13 source.t1 1.3205
R118 source.n13 source.t12 1.3205
R119 source.n15 source.n14 0.5005
R120 source.n14 source.n12 0.5005
R121 source.n12 source.n10 0.5005
R122 source.n10 source.n8 0.5005
R123 source.n7 source.n6 0.5005
R124 source.n6 source.n4 0.5005
R125 source.n4 source.n2 0.5005
R126 source.n2 source.n0 0.5005
R127 source.n18 source.n16 0.5005
R128 source.n20 source.n18 0.5005
R129 source.n22 source.n20 0.5005
R130 source.n23 source.n22 0.5005
R131 source.n26 source.n24 0.5005
R132 source.n28 source.n26 0.5005
R133 source.n30 source.n28 0.5005
R134 source.n31 source.n30 0.5005
R135 source.n8 source.n7 0.470328
R136 source.n24 source.n23 0.470328
R137 source source.n32 0.188
R138 drain_left.n9 drain_left.n7 61.3798
R139 drain_left.n5 drain_left.n3 61.3796
R140 drain_left.n2 drain_left.n0 61.3796
R141 drain_left.n11 drain_left.n10 60.8798
R142 drain_left.n9 drain_left.n8 60.8798
R143 drain_left.n13 drain_left.n12 60.8796
R144 drain_left.n5 drain_left.n4 60.8796
R145 drain_left.n2 drain_left.n1 60.8796
R146 drain_left drain_left.n6 32.8898
R147 drain_left drain_left.n13 6.15322
R148 drain_left.n3 drain_left.t1 1.3205
R149 drain_left.n3 drain_left.t12 1.3205
R150 drain_left.n4 drain_left.t10 1.3205
R151 drain_left.n4 drain_left.t3 1.3205
R152 drain_left.n1 drain_left.t13 1.3205
R153 drain_left.n1 drain_left.t8 1.3205
R154 drain_left.n0 drain_left.t4 1.3205
R155 drain_left.n0 drain_left.t2 1.3205
R156 drain_left.n12 drain_left.t7 1.3205
R157 drain_left.n12 drain_left.t11 1.3205
R158 drain_left.n10 drain_left.t6 1.3205
R159 drain_left.n10 drain_left.t0 1.3205
R160 drain_left.n8 drain_left.t5 1.3205
R161 drain_left.n8 drain_left.t15 1.3205
R162 drain_left.n7 drain_left.t9 1.3205
R163 drain_left.n7 drain_left.t14 1.3205
R164 drain_left.n11 drain_left.n9 0.5005
R165 drain_left.n13 drain_left.n11 0.5005
R166 drain_left.n6 drain_left.n5 0.195154
R167 drain_left.n6 drain_left.n2 0.195154
R168 minus.n19 minus.t4 1612.22
R169 minus.n4 minus.t9 1612.22
R170 minus.n40 minus.t13 1612.22
R171 minus.n25 minus.t3 1612.22
R172 minus.n18 minus.t12 1571.32
R173 minus.n16 minus.t5 1571.32
R174 minus.n1 minus.t11 1571.32
R175 minus.n10 minus.t1 1571.32
R176 minus.n3 minus.t8 1571.32
R177 minus.n5 minus.t2 1571.32
R178 minus.n39 minus.t14 1571.32
R179 minus.n37 minus.t0 1571.32
R180 minus.n22 minus.t7 1571.32
R181 minus.n31 minus.t10 1571.32
R182 minus.n24 minus.t15 1571.32
R183 minus.n26 minus.t6 1571.32
R184 minus.n7 minus.n4 161.489
R185 minus.n28 minus.n25 161.489
R186 minus.n20 minus.n19 161.3
R187 minus.n17 minus.n0 161.3
R188 minus.n15 minus.n14 161.3
R189 minus.n13 minus.n12 161.3
R190 minus.n11 minus.n2 161.3
R191 minus.n9 minus.n8 161.3
R192 minus.n7 minus.n6 161.3
R193 minus.n41 minus.n40 161.3
R194 minus.n38 minus.n21 161.3
R195 minus.n36 minus.n35 161.3
R196 minus.n34 minus.n33 161.3
R197 minus.n32 minus.n23 161.3
R198 minus.n30 minus.n29 161.3
R199 minus.n28 minus.n27 161.3
R200 minus.n12 minus.n11 73.0308
R201 minus.n33 minus.n32 73.0308
R202 minus.n15 minus.n1 67.1884
R203 minus.n10 minus.n9 67.1884
R204 minus.n31 minus.n30 67.1884
R205 minus.n36 minus.n22 67.1884
R206 minus.n17 minus.n16 55.5035
R207 minus.n6 minus.n3 55.5035
R208 minus.n27 minus.n24 55.5035
R209 minus.n38 minus.n37 55.5035
R210 minus.n19 minus.n18 43.8187
R211 minus.n5 minus.n4 43.8187
R212 minus.n26 minus.n25 43.8187
R213 minus.n40 minus.n39 43.8187
R214 minus.n42 minus.n20 38.027
R215 minus.n18 minus.n17 29.2126
R216 minus.n6 minus.n5 29.2126
R217 minus.n27 minus.n26 29.2126
R218 minus.n39 minus.n38 29.2126
R219 minus.n16 minus.n15 17.5278
R220 minus.n9 minus.n3 17.5278
R221 minus.n30 minus.n24 17.5278
R222 minus.n37 minus.n36 17.5278
R223 minus.n42 minus.n41 6.46641
R224 minus.n12 minus.n1 5.84292
R225 minus.n11 minus.n10 5.84292
R226 minus.n32 minus.n31 5.84292
R227 minus.n33 minus.n22 5.84292
R228 minus.n20 minus.n0 0.189894
R229 minus.n14 minus.n0 0.189894
R230 minus.n14 minus.n13 0.189894
R231 minus.n13 minus.n2 0.189894
R232 minus.n8 minus.n2 0.189894
R233 minus.n8 minus.n7 0.189894
R234 minus.n29 minus.n28 0.189894
R235 minus.n29 minus.n23 0.189894
R236 minus.n34 minus.n23 0.189894
R237 minus.n35 minus.n34 0.189894
R238 minus.n35 minus.n21 0.189894
R239 minus.n41 minus.n21 0.189894
R240 minus minus.n42 0.188
R241 drain_right.n9 drain_right.n7 61.3796
R242 drain_right.n5 drain_right.n3 61.3796
R243 drain_right.n2 drain_right.n0 61.3796
R244 drain_right.n9 drain_right.n8 60.8798
R245 drain_right.n11 drain_right.n10 60.8798
R246 drain_right.n13 drain_right.n12 60.8798
R247 drain_right.n5 drain_right.n4 60.8796
R248 drain_right.n2 drain_right.n1 60.8796
R249 drain_right drain_right.n6 32.3366
R250 drain_right drain_right.n13 6.15322
R251 drain_right.n3 drain_right.t1 1.3205
R252 drain_right.n3 drain_right.t2 1.3205
R253 drain_right.n4 drain_right.t8 1.3205
R254 drain_right.n4 drain_right.t15 1.3205
R255 drain_right.n1 drain_right.t0 1.3205
R256 drain_right.n1 drain_right.t5 1.3205
R257 drain_right.n0 drain_right.t12 1.3205
R258 drain_right.n0 drain_right.t9 1.3205
R259 drain_right.n7 drain_right.t13 1.3205
R260 drain_right.n7 drain_right.t6 1.3205
R261 drain_right.n8 drain_right.t14 1.3205
R262 drain_right.n8 drain_right.t7 1.3205
R263 drain_right.n10 drain_right.t10 1.3205
R264 drain_right.n10 drain_right.t4 1.3205
R265 drain_right.n12 drain_right.t11 1.3205
R266 drain_right.n12 drain_right.t3 1.3205
R267 drain_right.n13 drain_right.n11 0.5005
R268 drain_right.n11 drain_right.n9 0.5005
R269 drain_right.n6 drain_right.n5 0.195154
R270 drain_right.n6 drain_right.n2 0.195154
C0 drain_left minus 0.171252f
C1 drain_right plus 0.324551f
C2 minus plus 5.90572f
C3 drain_left plus 6.52242f
C4 drain_right source 40.862f
C5 source minus 5.86201f
C6 source drain_left 40.862103f
C7 drain_right minus 6.35208f
C8 source plus 5.87605f
C9 drain_right drain_left 0.897273f
C10 drain_right a_n1760_n3888# 7.33627f
C11 drain_left a_n1760_n3888# 7.60889f
C12 source a_n1760_n3888# 10.253778f
C13 minus a_n1760_n3888# 7.052824f
C14 plus a_n1760_n3888# 9.28068f
C15 drain_right.t12 a_n1760_n3888# 0.429145f
C16 drain_right.t9 a_n1760_n3888# 0.429145f
C17 drain_right.n0 a_n1760_n3888# 3.88245f
C18 drain_right.t0 a_n1760_n3888# 0.429145f
C19 drain_right.t5 a_n1760_n3888# 0.429145f
C20 drain_right.n1 a_n1760_n3888# 3.87897f
C21 drain_right.n2 a_n1760_n3888# 0.806174f
C22 drain_right.t1 a_n1760_n3888# 0.429145f
C23 drain_right.t2 a_n1760_n3888# 0.429145f
C24 drain_right.n3 a_n1760_n3888# 3.88245f
C25 drain_right.t8 a_n1760_n3888# 0.429145f
C26 drain_right.t15 a_n1760_n3888# 0.429145f
C27 drain_right.n4 a_n1760_n3888# 3.87897f
C28 drain_right.n5 a_n1760_n3888# 0.806174f
C29 drain_right.n6 a_n1760_n3888# 1.91864f
C30 drain_right.t13 a_n1760_n3888# 0.429145f
C31 drain_right.t6 a_n1760_n3888# 0.429145f
C32 drain_right.n7 a_n1760_n3888# 3.88244f
C33 drain_right.t14 a_n1760_n3888# 0.429145f
C34 drain_right.t7 a_n1760_n3888# 0.429145f
C35 drain_right.n8 a_n1760_n3888# 3.87897f
C36 drain_right.n9 a_n1760_n3888# 0.83749f
C37 drain_right.t10 a_n1760_n3888# 0.429145f
C38 drain_right.t4 a_n1760_n3888# 0.429145f
C39 drain_right.n10 a_n1760_n3888# 3.87897f
C40 drain_right.n11 a_n1760_n3888# 0.413189f
C41 drain_right.t11 a_n1760_n3888# 0.429145f
C42 drain_right.t3 a_n1760_n3888# 0.429145f
C43 drain_right.n12 a_n1760_n3888# 3.87897f
C44 drain_right.n13 a_n1760_n3888# 0.712031f
C45 minus.n0 a_n1760_n3888# 0.052467f
C46 minus.t4 a_n1760_n3888# 0.560564f
C47 minus.t12 a_n1760_n3888# 0.555063f
C48 minus.t5 a_n1760_n3888# 0.555063f
C49 minus.t11 a_n1760_n3888# 0.555063f
C50 minus.n1 a_n1760_n3888# 0.215899f
C51 minus.n2 a_n1760_n3888# 0.052467f
C52 minus.t1 a_n1760_n3888# 0.555063f
C53 minus.t8 a_n1760_n3888# 0.555063f
C54 minus.n3 a_n1760_n3888# 0.215899f
C55 minus.t9 a_n1760_n3888# 0.560564f
C56 minus.n4 a_n1760_n3888# 0.231434f
C57 minus.t2 a_n1760_n3888# 0.555063f
C58 minus.n5 a_n1760_n3888# 0.215899f
C59 minus.n6 a_n1760_n3888# 0.019993f
C60 minus.n7 a_n1760_n3888# 0.114888f
C61 minus.n8 a_n1760_n3888# 0.052467f
C62 minus.n9 a_n1760_n3888# 0.019993f
C63 minus.n10 a_n1760_n3888# 0.215899f
C64 minus.n11 a_n1760_n3888# 0.018699f
C65 minus.n12 a_n1760_n3888# 0.018699f
C66 minus.n13 a_n1760_n3888# 0.052467f
C67 minus.n14 a_n1760_n3888# 0.052467f
C68 minus.n15 a_n1760_n3888# 0.019993f
C69 minus.n16 a_n1760_n3888# 0.215899f
C70 minus.n17 a_n1760_n3888# 0.019993f
C71 minus.n18 a_n1760_n3888# 0.215899f
C72 minus.n19 a_n1760_n3888# 0.231361f
C73 minus.n20 a_n1760_n3888# 2.00025f
C74 minus.n21 a_n1760_n3888# 0.052467f
C75 minus.t14 a_n1760_n3888# 0.555063f
C76 minus.t0 a_n1760_n3888# 0.555063f
C77 minus.t7 a_n1760_n3888# 0.555063f
C78 minus.n22 a_n1760_n3888# 0.215899f
C79 minus.n23 a_n1760_n3888# 0.052467f
C80 minus.t10 a_n1760_n3888# 0.555063f
C81 minus.t15 a_n1760_n3888# 0.555063f
C82 minus.n24 a_n1760_n3888# 0.215899f
C83 minus.t3 a_n1760_n3888# 0.560564f
C84 minus.n25 a_n1760_n3888# 0.231434f
C85 minus.t6 a_n1760_n3888# 0.555063f
C86 minus.n26 a_n1760_n3888# 0.215899f
C87 minus.n27 a_n1760_n3888# 0.019993f
C88 minus.n28 a_n1760_n3888# 0.114888f
C89 minus.n29 a_n1760_n3888# 0.052467f
C90 minus.n30 a_n1760_n3888# 0.019993f
C91 minus.n31 a_n1760_n3888# 0.215899f
C92 minus.n32 a_n1760_n3888# 0.018699f
C93 minus.n33 a_n1760_n3888# 0.018699f
C94 minus.n34 a_n1760_n3888# 0.052467f
C95 minus.n35 a_n1760_n3888# 0.052467f
C96 minus.n36 a_n1760_n3888# 0.019993f
C97 minus.n37 a_n1760_n3888# 0.215899f
C98 minus.n38 a_n1760_n3888# 0.019993f
C99 minus.n39 a_n1760_n3888# 0.215899f
C100 minus.t13 a_n1760_n3888# 0.560564f
C101 minus.n40 a_n1760_n3888# 0.231361f
C102 minus.n41 a_n1760_n3888# 0.338856f
C103 minus.n42 a_n1760_n3888# 2.41788f
C104 drain_left.t4 a_n1760_n3888# 0.428768f
C105 drain_left.t2 a_n1760_n3888# 0.428768f
C106 drain_left.n0 a_n1760_n3888# 3.87905f
C107 drain_left.t13 a_n1760_n3888# 0.428768f
C108 drain_left.t8 a_n1760_n3888# 0.428768f
C109 drain_left.n1 a_n1760_n3888# 3.87556f
C110 drain_left.n2 a_n1760_n3888# 0.805466f
C111 drain_left.t1 a_n1760_n3888# 0.428768f
C112 drain_left.t12 a_n1760_n3888# 0.428768f
C113 drain_left.n3 a_n1760_n3888# 3.87905f
C114 drain_left.t10 a_n1760_n3888# 0.428768f
C115 drain_left.t3 a_n1760_n3888# 0.428768f
C116 drain_left.n4 a_n1760_n3888# 3.87556f
C117 drain_left.n5 a_n1760_n3888# 0.805466f
C118 drain_left.n6 a_n1760_n3888# 1.99234f
C119 drain_left.t9 a_n1760_n3888# 0.428768f
C120 drain_left.t14 a_n1760_n3888# 0.428768f
C121 drain_left.n7 a_n1760_n3888# 3.87905f
C122 drain_left.t5 a_n1760_n3888# 0.428768f
C123 drain_left.t15 a_n1760_n3888# 0.428768f
C124 drain_left.n8 a_n1760_n3888# 3.87557f
C125 drain_left.n9 a_n1760_n3888# 0.836742f
C126 drain_left.t6 a_n1760_n3888# 0.428768f
C127 drain_left.t0 a_n1760_n3888# 0.428768f
C128 drain_left.n10 a_n1760_n3888# 3.87557f
C129 drain_left.n11 a_n1760_n3888# 0.412827f
C130 drain_left.t7 a_n1760_n3888# 0.428768f
C131 drain_left.t11 a_n1760_n3888# 0.428768f
C132 drain_left.n12 a_n1760_n3888# 3.87555f
C133 drain_left.n13 a_n1760_n3888# 0.711419f
C134 source.t28 a_n1760_n3888# 3.9676f
C135 source.n0 a_n1760_n3888# 1.83102f
C136 source.t26 a_n1760_n3888# 0.354041f
C137 source.t18 a_n1760_n3888# 0.354041f
C138 source.n1 a_n1760_n3888# 3.10995f
C139 source.n2 a_n1760_n3888# 0.390447f
C140 source.t24 a_n1760_n3888# 0.354041f
C141 source.t19 a_n1760_n3888# 0.354041f
C142 source.n3 a_n1760_n3888# 3.10995f
C143 source.n4 a_n1760_n3888# 0.390447f
C144 source.t17 a_n1760_n3888# 0.354041f
C145 source.t23 a_n1760_n3888# 0.354041f
C146 source.n5 a_n1760_n3888# 3.10995f
C147 source.n6 a_n1760_n3888# 0.390447f
C148 source.t31 a_n1760_n3888# 3.9676f
C149 source.n7 a_n1760_n3888# 0.495458f
C150 source.t0 a_n1760_n3888# 3.9676f
C151 source.n8 a_n1760_n3888# 0.495458f
C152 source.t11 a_n1760_n3888# 0.354041f
C153 source.t14 a_n1760_n3888# 0.354041f
C154 source.n9 a_n1760_n3888# 3.10995f
C155 source.n10 a_n1760_n3888# 0.390447f
C156 source.t4 a_n1760_n3888# 0.354041f
C157 source.t6 a_n1760_n3888# 0.354041f
C158 source.n11 a_n1760_n3888# 3.10995f
C159 source.n12 a_n1760_n3888# 0.390447f
C160 source.t1 a_n1760_n3888# 0.354041f
C161 source.t12 a_n1760_n3888# 0.354041f
C162 source.n13 a_n1760_n3888# 3.10995f
C163 source.n14 a_n1760_n3888# 0.390447f
C164 source.t9 a_n1760_n3888# 3.9676f
C165 source.n15 a_n1760_n3888# 2.326f
C166 source.t20 a_n1760_n3888# 3.9676f
C167 source.n16 a_n1760_n3888# 2.32601f
C168 source.t29 a_n1760_n3888# 0.354041f
C169 source.t21 a_n1760_n3888# 0.354041f
C170 source.n17 a_n1760_n3888# 3.10995f
C171 source.n18 a_n1760_n3888# 0.390451f
C172 source.t25 a_n1760_n3888# 0.354041f
C173 source.t22 a_n1760_n3888# 0.354041f
C174 source.n19 a_n1760_n3888# 3.10995f
C175 source.n20 a_n1760_n3888# 0.390451f
C176 source.t30 a_n1760_n3888# 0.354041f
C177 source.t16 a_n1760_n3888# 0.354041f
C178 source.n21 a_n1760_n3888# 3.10995f
C179 source.n22 a_n1760_n3888# 0.390451f
C180 source.t27 a_n1760_n3888# 3.9676f
C181 source.n23 a_n1760_n3888# 0.495463f
C182 source.t2 a_n1760_n3888# 3.9676f
C183 source.n24 a_n1760_n3888# 0.495463f
C184 source.t7 a_n1760_n3888# 0.354041f
C185 source.t10 a_n1760_n3888# 0.354041f
C186 source.n25 a_n1760_n3888# 3.10995f
C187 source.n26 a_n1760_n3888# 0.390451f
C188 source.t13 a_n1760_n3888# 0.354041f
C189 source.t8 a_n1760_n3888# 0.354041f
C190 source.n27 a_n1760_n3888# 3.10995f
C191 source.n28 a_n1760_n3888# 0.390451f
C192 source.t15 a_n1760_n3888# 0.354041f
C193 source.t5 a_n1760_n3888# 0.354041f
C194 source.n29 a_n1760_n3888# 3.10995f
C195 source.n30 a_n1760_n3888# 0.390451f
C196 source.t3 a_n1760_n3888# 3.9676f
C197 source.n31 a_n1760_n3888# 0.660748f
C198 source.n32 a_n1760_n3888# 2.18148f
C199 plus.n0 a_n1760_n3888# 0.053064f
C200 plus.t8 a_n1760_n3888# 0.561385f
C201 plus.t15 a_n1760_n3888# 0.561385f
C202 plus.t9 a_n1760_n3888# 0.561385f
C203 plus.n1 a_n1760_n3888# 0.218358f
C204 plus.n2 a_n1760_n3888# 0.053064f
C205 plus.t0 a_n1760_n3888# 0.561385f
C206 plus.t10 a_n1760_n3888# 0.561385f
C207 plus.n3 a_n1760_n3888# 0.218358f
C208 plus.t6 a_n1760_n3888# 0.566949f
C209 plus.n4 a_n1760_n3888# 0.23407f
C210 plus.t1 a_n1760_n3888# 0.561385f
C211 plus.n5 a_n1760_n3888# 0.218358f
C212 plus.n6 a_n1760_n3888# 0.020221f
C213 plus.n7 a_n1760_n3888# 0.116197f
C214 plus.n8 a_n1760_n3888# 0.053064f
C215 plus.n9 a_n1760_n3888# 0.020221f
C216 plus.n10 a_n1760_n3888# 0.218358f
C217 plus.n11 a_n1760_n3888# 0.018912f
C218 plus.n12 a_n1760_n3888# 0.018912f
C219 plus.n13 a_n1760_n3888# 0.053064f
C220 plus.n14 a_n1760_n3888# 0.053064f
C221 plus.n15 a_n1760_n3888# 0.020221f
C222 plus.n16 a_n1760_n3888# 0.218358f
C223 plus.n17 a_n1760_n3888# 0.020221f
C224 plus.n18 a_n1760_n3888# 0.218358f
C225 plus.t4 a_n1760_n3888# 0.566949f
C226 plus.n19 a_n1760_n3888# 0.233996f
C227 plus.n20 a_n1760_n3888# 0.666364f
C228 plus.n21 a_n1760_n3888# 0.053064f
C229 plus.t11 a_n1760_n3888# 0.566949f
C230 plus.t13 a_n1760_n3888# 0.561385f
C231 plus.t2 a_n1760_n3888# 0.561385f
C232 plus.t7 a_n1760_n3888# 0.561385f
C233 plus.n22 a_n1760_n3888# 0.218358f
C234 plus.n23 a_n1760_n3888# 0.053064f
C235 plus.t5 a_n1760_n3888# 0.561385f
C236 plus.t12 a_n1760_n3888# 0.561385f
C237 plus.n24 a_n1760_n3888# 0.218358f
C238 plus.t3 a_n1760_n3888# 0.566949f
C239 plus.n25 a_n1760_n3888# 0.23407f
C240 plus.t14 a_n1760_n3888# 0.561385f
C241 plus.n26 a_n1760_n3888# 0.218358f
C242 plus.n27 a_n1760_n3888# 0.020221f
C243 plus.n28 a_n1760_n3888# 0.116197f
C244 plus.n29 a_n1760_n3888# 0.053064f
C245 plus.n30 a_n1760_n3888# 0.020221f
C246 plus.n31 a_n1760_n3888# 0.218358f
C247 plus.n32 a_n1760_n3888# 0.018912f
C248 plus.n33 a_n1760_n3888# 0.018912f
C249 plus.n34 a_n1760_n3888# 0.053064f
C250 plus.n35 a_n1760_n3888# 0.053064f
C251 plus.n36 a_n1760_n3888# 0.020221f
C252 plus.n37 a_n1760_n3888# 0.218358f
C253 plus.n38 a_n1760_n3888# 0.020221f
C254 plus.n39 a_n1760_n3888# 0.218358f
C255 plus.n40 a_n1760_n3888# 0.233996f
C256 plus.n41 a_n1760_n3888# 1.66215f
.ends

