* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t37 plus.t0 drain_left.t9 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 drain_right.t19 minus.t0 source.t2 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 drain_right.t18 minus.t1 source.t9 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X3 source.t36 plus.t1 drain_left.t19 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X4 source.t1 minus.t2 drain_right.t17 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X5 source.t35 plus.t2 drain_left.t14 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X6 drain_left.t2 plus.t3 source.t34 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X7 drain_right.t16 minus.t3 source.t5 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X8 a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X9 drain_left.t3 plus.t4 source.t33 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 source.t12 minus.t4 drain_right.t15 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X11 a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X12 source.t16 minus.t5 drain_right.t14 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X13 drain_right.t13 minus.t6 source.t11 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X14 source.t10 minus.t7 drain_right.t12 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X15 a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X16 source.t32 plus.t5 drain_left.t10 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 drain_left.t6 plus.t6 source.t31 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X19 drain_right.t11 minus.t8 source.t38 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X20 drain_right.t10 minus.t9 source.t39 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X21 source.t4 minus.t10 drain_right.t9 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X22 source.t0 minus.t11 drain_right.t8 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 drain_left.t0 plus.t7 source.t30 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X24 drain_right.t7 minus.t12 source.t3 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X25 source.t29 plus.t8 drain_left.t7 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X26 drain_left.t4 plus.t9 source.t28 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X27 source.t27 plus.t10 drain_left.t8 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X28 drain_right.t6 minus.t13 source.t17 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X29 drain_right.t5 minus.t14 source.t15 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X30 source.t7 minus.t15 drain_right.t4 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X31 drain_left.t11 plus.t11 source.t26 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X32 source.t13 minus.t16 drain_right.t3 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X33 drain_right.t2 minus.t17 source.t14 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X34 drain_left.t5 plus.t12 source.t25 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X35 source.t24 plus.t13 drain_left.t1 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X36 source.t23 plus.t14 drain_left.t13 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X37 drain_left.t12 plus.t15 source.t22 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X38 source.t6 minus.t18 drain_right.t1 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X39 source.t21 plus.t16 drain_left.t15 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X40 drain_left.t16 plus.t17 source.t20 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X41 drain_left.t17 plus.t18 source.t19 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X42 source.t8 minus.t19 drain_right.t0 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X43 source.t18 plus.t19 drain_left.t18 a_n2146_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
R0 plus.n6 plus.t10 752.942
R1 plus.n27 plus.t12 752.942
R2 plus.n36 plus.t3 752.942
R3 plus.n56 plus.t2 752.942
R4 plus.n5 plus.t18 690.867
R5 plus.n9 plus.t14 690.867
R6 plus.n3 plus.t11 690.867
R7 plus.n15 plus.t19 690.867
R8 plus.n17 plus.t17 690.867
R9 plus.n18 plus.t13 690.867
R10 plus.n24 plus.t9 690.867
R11 plus.n26 plus.t16 690.867
R12 plus.n35 plus.t1 690.867
R13 plus.n39 plus.t7 690.867
R14 plus.n33 plus.t5 690.867
R15 plus.n45 plus.t4 690.867
R16 plus.n47 plus.t0 690.867
R17 plus.n32 plus.t15 690.867
R18 plus.n53 plus.t8 690.867
R19 plus.n55 plus.t6 690.867
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 69.3793
R47 plus.n19 plus.n18 69.3793
R48 plus.n48 plus.n32 69.3793
R49 plus.n44 plus.n33 69.3793
R50 plus.n9 plus.n8 54.7732
R51 plus.n25 plus.n24 54.7732
R52 plus.n54 plus.n53 54.7732
R53 plus.n39 plus.n38 54.7732
R54 plus.n16 plus.n15 47.4702
R55 plus.n17 plus.n16 47.4702
R56 plus.n47 plus.n46 47.4702
R57 plus.n46 plus.n45 47.4702
R58 plus.n8 plus.n5 40.1672
R59 plus.n26 plus.n25 40.1672
R60 plus.n55 plus.n54 40.1672
R61 plus.n38 plus.n35 40.1672
R62 plus.n6 plus.n5 32.8641
R63 plus.n27 plus.n26 32.8641
R64 plus.n56 plus.n55 32.8641
R65 plus.n36 plus.n35 32.8641
R66 plus plus.n57 27.7831
R67 plus.n15 plus.n14 25.5611
R68 plus.n19 plus.n17 25.5611
R69 plus.n48 plus.n47 25.5611
R70 plus.n45 plus.n44 25.5611
R71 plus.n10 plus.n9 18.2581
R72 plus.n24 plus.n23 18.2581
R73 plus.n53 plus.n52 18.2581
R74 plus.n40 plus.n39 18.2581
R75 plus plus.n28 8.79595
R76 plus.n11 plus.n3 3.65202
R77 plus.n18 plus.n1 3.65202
R78 plus.n32 plus.n30 3.65202
R79 plus.n41 plus.n33 3.65202
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 drain_left.n10 drain_left.n8 80.3335
R99 drain_left.n6 drain_left.n4 80.3334
R100 drain_left.n2 drain_left.n0 80.3334
R101 drain_left.n16 drain_left.n15 79.7731
R102 drain_left.n14 drain_left.n13 79.7731
R103 drain_left.n12 drain_left.n11 79.7731
R104 drain_left.n10 drain_left.n9 79.7731
R105 drain_left.n7 drain_left.n3 79.773
R106 drain_left.n6 drain_left.n5 79.773
R107 drain_left.n2 drain_left.n1 79.773
R108 drain_left drain_left.n7 25.0317
R109 drain_left.n3 drain_left.t9 10.0005
R110 drain_left.n3 drain_left.t3 10.0005
R111 drain_left.n4 drain_left.t19 10.0005
R112 drain_left.n4 drain_left.t2 10.0005
R113 drain_left.n5 drain_left.t10 10.0005
R114 drain_left.n5 drain_left.t0 10.0005
R115 drain_left.n1 drain_left.t7 10.0005
R116 drain_left.n1 drain_left.t12 10.0005
R117 drain_left.n0 drain_left.t14 10.0005
R118 drain_left.n0 drain_left.t6 10.0005
R119 drain_left.n15 drain_left.t15 10.0005
R120 drain_left.n15 drain_left.t5 10.0005
R121 drain_left.n13 drain_left.t1 10.0005
R122 drain_left.n13 drain_left.t4 10.0005
R123 drain_left.n11 drain_left.t18 10.0005
R124 drain_left.n11 drain_left.t16 10.0005
R125 drain_left.n9 drain_left.t13 10.0005
R126 drain_left.n9 drain_left.t11 10.0005
R127 drain_left.n8 drain_left.t8 10.0005
R128 drain_left.n8 drain_left.t17 10.0005
R129 drain_left drain_left.n16 6.21356
R130 drain_left.n12 drain_left.n10 0.560845
R131 drain_left.n14 drain_left.n12 0.560845
R132 drain_left.n16 drain_left.n14 0.560845
R133 drain_left.n7 drain_left.n6 0.505499
R134 drain_left.n7 drain_left.n2 0.505499
R135 source.n0 source.t25 73.0943
R136 source.n9 source.t27 73.0943
R137 source.n10 source.t38 73.0943
R138 source.n19 source.t6 73.0943
R139 source.n39 source.t11 73.0942
R140 source.n30 source.t16 73.0942
R141 source.n29 source.t34 73.0942
R142 source.n20 source.t35 73.0942
R143 source.n2 source.n1 63.0943
R144 source.n4 source.n3 63.0943
R145 source.n6 source.n5 63.0943
R146 source.n8 source.n7 63.0943
R147 source.n12 source.n11 63.0943
R148 source.n14 source.n13 63.0943
R149 source.n16 source.n15 63.0943
R150 source.n18 source.n17 63.0943
R151 source.n38 source.n37 63.0942
R152 source.n36 source.n35 63.0942
R153 source.n34 source.n33 63.0942
R154 source.n32 source.n31 63.0942
R155 source.n28 source.n27 63.0942
R156 source.n26 source.n25 63.0942
R157 source.n24 source.n23 63.0942
R158 source.n22 source.n21 63.0942
R159 source.n20 source.n19 15.0299
R160 source.n37 source.t2 10.0005
R161 source.n37 source.t0 10.0005
R162 source.n35 source.t5 10.0005
R163 source.n35 source.t1 10.0005
R164 source.n33 source.t14 10.0005
R165 source.n33 source.t12 10.0005
R166 source.n31 source.t9 10.0005
R167 source.n31 source.t8 10.0005
R168 source.n27 source.t30 10.0005
R169 source.n27 source.t36 10.0005
R170 source.n25 source.t33 10.0005
R171 source.n25 source.t32 10.0005
R172 source.n23 source.t22 10.0005
R173 source.n23 source.t37 10.0005
R174 source.n21 source.t31 10.0005
R175 source.n21 source.t29 10.0005
R176 source.n1 source.t28 10.0005
R177 source.n1 source.t21 10.0005
R178 source.n3 source.t20 10.0005
R179 source.n3 source.t24 10.0005
R180 source.n5 source.t26 10.0005
R181 source.n5 source.t18 10.0005
R182 source.n7 source.t19 10.0005
R183 source.n7 source.t23 10.0005
R184 source.n11 source.t17 10.0005
R185 source.n11 source.t10 10.0005
R186 source.n13 source.t39 10.0005
R187 source.n13 source.t4 10.0005
R188 source.n15 source.t15 10.0005
R189 source.n15 source.t13 10.0005
R190 source.n17 source.t3 10.0005
R191 source.n17 source.t7 10.0005
R192 source.n40 source.n0 9.48679
R193 source.n40 source.n39 5.5436
R194 source.n19 source.n18 0.560845
R195 source.n18 source.n16 0.560845
R196 source.n16 source.n14 0.560845
R197 source.n14 source.n12 0.560845
R198 source.n12 source.n10 0.560845
R199 source.n9 source.n8 0.560845
R200 source.n8 source.n6 0.560845
R201 source.n6 source.n4 0.560845
R202 source.n4 source.n2 0.560845
R203 source.n2 source.n0 0.560845
R204 source.n22 source.n20 0.560845
R205 source.n24 source.n22 0.560845
R206 source.n26 source.n24 0.560845
R207 source.n28 source.n26 0.560845
R208 source.n29 source.n28 0.560845
R209 source.n32 source.n30 0.560845
R210 source.n34 source.n32 0.560845
R211 source.n36 source.n34 0.560845
R212 source.n38 source.n36 0.560845
R213 source.n39 source.n38 0.560845
R214 source.n10 source.n9 0.470328
R215 source.n30 source.n29 0.470328
R216 source source.n40 0.188
R217 minus.n27 minus.t18 752.942
R218 minus.n7 minus.t8 752.942
R219 minus.n56 minus.t6 752.942
R220 minus.n35 minus.t5 752.942
R221 minus.n26 minus.t12 690.867
R222 minus.n24 minus.t15 690.867
R223 minus.n3 minus.t14 690.867
R224 minus.n18 minus.t16 690.867
R225 minus.n16 minus.t9 690.867
R226 minus.n4 minus.t10 690.867
R227 minus.n10 minus.t13 690.867
R228 minus.n6 minus.t7 690.867
R229 minus.n55 minus.t11 690.867
R230 minus.n53 minus.t0 690.867
R231 minus.n47 minus.t2 690.867
R232 minus.n46 minus.t3 690.867
R233 minus.n44 minus.t4 690.867
R234 minus.n32 minus.t17 690.867
R235 minus.n38 minus.t19 690.867
R236 minus.n34 minus.t1 690.867
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 69.3793
R264 minus.n15 minus.n4 69.3793
R265 minus.n43 minus.n32 69.3793
R266 minus.n48 minus.n47 69.3793
R267 minus.n25 minus.n24 54.7732
R268 minus.n10 minus.n9 54.7732
R269 minus.n38 minus.n37 54.7732
R270 minus.n54 minus.n53 54.7732
R271 minus.n18 minus.n17 47.4702
R272 minus.n17 minus.n16 47.4702
R273 minus.n45 minus.n44 47.4702
R274 minus.n46 minus.n45 47.4702
R275 minus.n26 minus.n25 40.1672
R276 minus.n9 minus.n6 40.1672
R277 minus.n37 minus.n34 40.1672
R278 minus.n55 minus.n54 40.1672
R279 minus.n27 minus.n26 32.8641
R280 minus.n7 minus.n6 32.8641
R281 minus.n35 minus.n34 32.8641
R282 minus.n56 minus.n55 32.8641
R283 minus.n58 minus.n28 30.4929
R284 minus.n19 minus.n18 25.5611
R285 minus.n16 minus.n15 25.5611
R286 minus.n44 minus.n43 25.5611
R287 minus.n48 minus.n46 25.5611
R288 minus.n24 minus.n23 18.2581
R289 minus.n11 minus.n10 18.2581
R290 minus.n39 minus.n38 18.2581
R291 minus.n53 minus.n52 18.2581
R292 minus.n58 minus.n57 6.56111
R293 minus.n3 minus.n1 3.65202
R294 minus.n12 minus.n4 3.65202
R295 minus.n40 minus.n32 3.65202
R296 minus.n47 minus.n30 3.65202
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 80.3335
R317 drain_right.n6 drain_right.n4 80.3334
R318 drain_right.n2 drain_right.n0 80.3334
R319 drain_right.n10 drain_right.n9 79.7731
R320 drain_right.n12 drain_right.n11 79.7731
R321 drain_right.n14 drain_right.n13 79.7731
R322 drain_right.n16 drain_right.n15 79.7731
R323 drain_right.n7 drain_right.n3 79.773
R324 drain_right.n6 drain_right.n5 79.773
R325 drain_right.n2 drain_right.n1 79.773
R326 drain_right drain_right.n7 24.4784
R327 drain_right.n3 drain_right.t15 10.0005
R328 drain_right.n3 drain_right.t16 10.0005
R329 drain_right.n4 drain_right.t8 10.0005
R330 drain_right.n4 drain_right.t13 10.0005
R331 drain_right.n5 drain_right.t17 10.0005
R332 drain_right.n5 drain_right.t19 10.0005
R333 drain_right.n1 drain_right.t0 10.0005
R334 drain_right.n1 drain_right.t2 10.0005
R335 drain_right.n0 drain_right.t14 10.0005
R336 drain_right.n0 drain_right.t18 10.0005
R337 drain_right.n8 drain_right.t12 10.0005
R338 drain_right.n8 drain_right.t11 10.0005
R339 drain_right.n9 drain_right.t9 10.0005
R340 drain_right.n9 drain_right.t6 10.0005
R341 drain_right.n11 drain_right.t3 10.0005
R342 drain_right.n11 drain_right.t10 10.0005
R343 drain_right.n13 drain_right.t4 10.0005
R344 drain_right.n13 drain_right.t5 10.0005
R345 drain_right.n15 drain_right.t1 10.0005
R346 drain_right.n15 drain_right.t7 10.0005
R347 drain_right drain_right.n16 6.21356
R348 drain_right.n16 drain_right.n14 0.560845
R349 drain_right.n14 drain_right.n12 0.560845
R350 drain_right.n12 drain_right.n10 0.560845
R351 drain_right.n7 drain_right.n6 0.505499
R352 drain_right.n7 drain_right.n2 0.505499
C0 drain_right source 12.1051f
C1 drain_left plus 1.71372f
C2 drain_left minus 0.176528f
C3 plus minus 4.15326f
C4 drain_left source 12.1046f
C5 plus source 1.58957f
C6 minus source 1.57557f
C7 drain_left drain_right 1.13565f
C8 drain_right plus 0.370515f
C9 drain_right minus 1.50305f
C10 drain_right a_n2146_n1488# 4.48305f
C11 drain_left a_n2146_n1488# 4.77538f
C12 source a_n2146_n1488# 3.899197f
C13 minus a_n2146_n1488# 7.197741f
C14 plus a_n2146_n1488# 7.97783f
C15 drain_right.t14 a_n2146_n1488# 0.089787f
C16 drain_right.t18 a_n2146_n1488# 0.089787f
C17 drain_right.n0 a_n2146_n1488# 0.490526f
C18 drain_right.t0 a_n2146_n1488# 0.089787f
C19 drain_right.t2 a_n2146_n1488# 0.089787f
C20 drain_right.n1 a_n2146_n1488# 0.488431f
C21 drain_right.n2 a_n2146_n1488# 0.585386f
C22 drain_right.t15 a_n2146_n1488# 0.089787f
C23 drain_right.t16 a_n2146_n1488# 0.089787f
C24 drain_right.n3 a_n2146_n1488# 0.488431f
C25 drain_right.t8 a_n2146_n1488# 0.089787f
C26 drain_right.t13 a_n2146_n1488# 0.089787f
C27 drain_right.n4 a_n2146_n1488# 0.490526f
C28 drain_right.t17 a_n2146_n1488# 0.089787f
C29 drain_right.t19 a_n2146_n1488# 0.089787f
C30 drain_right.n5 a_n2146_n1488# 0.488431f
C31 drain_right.n6 a_n2146_n1488# 0.585386f
C32 drain_right.n7 a_n2146_n1488# 1.03111f
C33 drain_right.t12 a_n2146_n1488# 0.089787f
C34 drain_right.t11 a_n2146_n1488# 0.089787f
C35 drain_right.n8 a_n2146_n1488# 0.490528f
C36 drain_right.t9 a_n2146_n1488# 0.089787f
C37 drain_right.t6 a_n2146_n1488# 0.089787f
C38 drain_right.n9 a_n2146_n1488# 0.488433f
C39 drain_right.n10 a_n2146_n1488# 0.588693f
C40 drain_right.t3 a_n2146_n1488# 0.089787f
C41 drain_right.t10 a_n2146_n1488# 0.089787f
C42 drain_right.n11 a_n2146_n1488# 0.488433f
C43 drain_right.n12 a_n2146_n1488# 0.29036f
C44 drain_right.t4 a_n2146_n1488# 0.089787f
C45 drain_right.t5 a_n2146_n1488# 0.089787f
C46 drain_right.n13 a_n2146_n1488# 0.488433f
C47 drain_right.n14 a_n2146_n1488# 0.29036f
C48 drain_right.t1 a_n2146_n1488# 0.089787f
C49 drain_right.t7 a_n2146_n1488# 0.089787f
C50 drain_right.n15 a_n2146_n1488# 0.488433f
C51 drain_right.n16 a_n2146_n1488# 0.49911f
C52 minus.n0 a_n2146_n1488# 0.029756f
C53 minus.t18 a_n2146_n1488# 0.041124f
C54 minus.t12 a_n2146_n1488# 0.038776f
C55 minus.t15 a_n2146_n1488# 0.038776f
C56 minus.n1 a_n2146_n1488# 0.01033f
C57 minus.n2 a_n2146_n1488# 0.029756f
C58 minus.t14 a_n2146_n1488# 0.038776f
C59 minus.n3 a_n2146_n1488# 0.027102f
C60 minus.t16 a_n2146_n1488# 0.038776f
C61 minus.t9 a_n2146_n1488# 0.038776f
C62 minus.t10 a_n2146_n1488# 0.038776f
C63 minus.n4 a_n2146_n1488# 0.027102f
C64 minus.n5 a_n2146_n1488# 0.029756f
C65 minus.t13 a_n2146_n1488# 0.038776f
C66 minus.t7 a_n2146_n1488# 0.038776f
C67 minus.n6 a_n2146_n1488# 0.027102f
C68 minus.t8 a_n2146_n1488# 0.041124f
C69 minus.n7 a_n2146_n1488# 0.038798f
C70 minus.n8 a_n2146_n1488# 0.068639f
C71 minus.n9 a_n2146_n1488# 0.012623f
C72 minus.n10 a_n2146_n1488# 0.027102f
C73 minus.n11 a_n2146_n1488# 0.012164f
C74 minus.n12 a_n2146_n1488# 0.01033f
C75 minus.n13 a_n2146_n1488# 0.029756f
C76 minus.n14 a_n2146_n1488# 0.029756f
C77 minus.n15 a_n2146_n1488# 0.012623f
C78 minus.n16 a_n2146_n1488# 0.027102f
C79 minus.n17 a_n2146_n1488# 0.012623f
C80 minus.n18 a_n2146_n1488# 0.027102f
C81 minus.n19 a_n2146_n1488# 0.012623f
C82 minus.n20 a_n2146_n1488# 0.029756f
C83 minus.n21 a_n2146_n1488# 0.029756f
C84 minus.n22 a_n2146_n1488# 0.029756f
C85 minus.n23 a_n2146_n1488# 0.012164f
C86 minus.n24 a_n2146_n1488# 0.027102f
C87 minus.n25 a_n2146_n1488# 0.012623f
C88 minus.n26 a_n2146_n1488# 0.027102f
C89 minus.n27 a_n2146_n1488# 0.038753f
C90 minus.n28 a_n2146_n1488# 0.797492f
C91 minus.n29 a_n2146_n1488# 0.029756f
C92 minus.t11 a_n2146_n1488# 0.038776f
C93 minus.t0 a_n2146_n1488# 0.038776f
C94 minus.n30 a_n2146_n1488# 0.01033f
C95 minus.n31 a_n2146_n1488# 0.029756f
C96 minus.t3 a_n2146_n1488# 0.038776f
C97 minus.t4 a_n2146_n1488# 0.038776f
C98 minus.t17 a_n2146_n1488# 0.038776f
C99 minus.n32 a_n2146_n1488# 0.027102f
C100 minus.n33 a_n2146_n1488# 0.029756f
C101 minus.t19 a_n2146_n1488# 0.038776f
C102 minus.t1 a_n2146_n1488# 0.038776f
C103 minus.n34 a_n2146_n1488# 0.027102f
C104 minus.t5 a_n2146_n1488# 0.041124f
C105 minus.n35 a_n2146_n1488# 0.038798f
C106 minus.n36 a_n2146_n1488# 0.068639f
C107 minus.n37 a_n2146_n1488# 0.012623f
C108 minus.n38 a_n2146_n1488# 0.027102f
C109 minus.n39 a_n2146_n1488# 0.012164f
C110 minus.n40 a_n2146_n1488# 0.01033f
C111 minus.n41 a_n2146_n1488# 0.029756f
C112 minus.n42 a_n2146_n1488# 0.029756f
C113 minus.n43 a_n2146_n1488# 0.012623f
C114 minus.n44 a_n2146_n1488# 0.027102f
C115 minus.n45 a_n2146_n1488# 0.012623f
C116 minus.n46 a_n2146_n1488# 0.027102f
C117 minus.t2 a_n2146_n1488# 0.038776f
C118 minus.n47 a_n2146_n1488# 0.027102f
C119 minus.n48 a_n2146_n1488# 0.012623f
C120 minus.n49 a_n2146_n1488# 0.029756f
C121 minus.n50 a_n2146_n1488# 0.029756f
C122 minus.n51 a_n2146_n1488# 0.029756f
C123 minus.n52 a_n2146_n1488# 0.012164f
C124 minus.n53 a_n2146_n1488# 0.027102f
C125 minus.n54 a_n2146_n1488# 0.012623f
C126 minus.n55 a_n2146_n1488# 0.027102f
C127 minus.t6 a_n2146_n1488# 0.041124f
C128 minus.n56 a_n2146_n1488# 0.038753f
C129 minus.n57 a_n2146_n1488# 0.198807f
C130 minus.n58 a_n2146_n1488# 0.98094f
C131 source.t25 a_n2146_n1488# 0.524536f
C132 source.n0 a_n2146_n1488# 0.692453f
C133 source.t28 a_n2146_n1488# 0.089059f
C134 source.t21 a_n2146_n1488# 0.089059f
C135 source.n1 a_n2146_n1488# 0.43325f
C136 source.n2 a_n2146_n1488# 0.30552f
C137 source.t20 a_n2146_n1488# 0.089059f
C138 source.t24 a_n2146_n1488# 0.089059f
C139 source.n3 a_n2146_n1488# 0.43325f
C140 source.n4 a_n2146_n1488# 0.30552f
C141 source.t26 a_n2146_n1488# 0.089059f
C142 source.t18 a_n2146_n1488# 0.089059f
C143 source.n5 a_n2146_n1488# 0.43325f
C144 source.n6 a_n2146_n1488# 0.30552f
C145 source.t19 a_n2146_n1488# 0.089059f
C146 source.t23 a_n2146_n1488# 0.089059f
C147 source.n7 a_n2146_n1488# 0.43325f
C148 source.n8 a_n2146_n1488# 0.30552f
C149 source.t27 a_n2146_n1488# 0.524535f
C150 source.n9 a_n2146_n1488# 0.367309f
C151 source.t38 a_n2146_n1488# 0.524535f
C152 source.n10 a_n2146_n1488# 0.367309f
C153 source.t17 a_n2146_n1488# 0.089059f
C154 source.t10 a_n2146_n1488# 0.089059f
C155 source.n11 a_n2146_n1488# 0.43325f
C156 source.n12 a_n2146_n1488# 0.30552f
C157 source.t39 a_n2146_n1488# 0.089059f
C158 source.t4 a_n2146_n1488# 0.089059f
C159 source.n13 a_n2146_n1488# 0.43325f
C160 source.n14 a_n2146_n1488# 0.30552f
C161 source.t15 a_n2146_n1488# 0.089059f
C162 source.t13 a_n2146_n1488# 0.089059f
C163 source.n15 a_n2146_n1488# 0.43325f
C164 source.n16 a_n2146_n1488# 0.30552f
C165 source.t3 a_n2146_n1488# 0.089059f
C166 source.t7 a_n2146_n1488# 0.089059f
C167 source.n17 a_n2146_n1488# 0.43325f
C168 source.n18 a_n2146_n1488# 0.30552f
C169 source.t6 a_n2146_n1488# 0.524535f
C170 source.n19 a_n2146_n1488# 0.951225f
C171 source.t35 a_n2146_n1488# 0.524533f
C172 source.n20 a_n2146_n1488# 0.951227f
C173 source.t31 a_n2146_n1488# 0.089059f
C174 source.t29 a_n2146_n1488# 0.089059f
C175 source.n21 a_n2146_n1488# 0.433248f
C176 source.n22 a_n2146_n1488# 0.305523f
C177 source.t22 a_n2146_n1488# 0.089059f
C178 source.t37 a_n2146_n1488# 0.089059f
C179 source.n23 a_n2146_n1488# 0.433248f
C180 source.n24 a_n2146_n1488# 0.305523f
C181 source.t33 a_n2146_n1488# 0.089059f
C182 source.t32 a_n2146_n1488# 0.089059f
C183 source.n25 a_n2146_n1488# 0.433248f
C184 source.n26 a_n2146_n1488# 0.305523f
C185 source.t30 a_n2146_n1488# 0.089059f
C186 source.t36 a_n2146_n1488# 0.089059f
C187 source.n27 a_n2146_n1488# 0.433248f
C188 source.n28 a_n2146_n1488# 0.305523f
C189 source.t34 a_n2146_n1488# 0.524533f
C190 source.n29 a_n2146_n1488# 0.367312f
C191 source.t16 a_n2146_n1488# 0.524533f
C192 source.n30 a_n2146_n1488# 0.367312f
C193 source.t9 a_n2146_n1488# 0.089059f
C194 source.t8 a_n2146_n1488# 0.089059f
C195 source.n31 a_n2146_n1488# 0.433248f
C196 source.n32 a_n2146_n1488# 0.305523f
C197 source.t14 a_n2146_n1488# 0.089059f
C198 source.t12 a_n2146_n1488# 0.089059f
C199 source.n33 a_n2146_n1488# 0.433248f
C200 source.n34 a_n2146_n1488# 0.305523f
C201 source.t5 a_n2146_n1488# 0.089059f
C202 source.t1 a_n2146_n1488# 0.089059f
C203 source.n35 a_n2146_n1488# 0.433248f
C204 source.n36 a_n2146_n1488# 0.305523f
C205 source.t2 a_n2146_n1488# 0.089059f
C206 source.t0 a_n2146_n1488# 0.089059f
C207 source.n37 a_n2146_n1488# 0.433248f
C208 source.n38 a_n2146_n1488# 0.305523f
C209 source.t11 a_n2146_n1488# 0.524533f
C210 source.n39 a_n2146_n1488# 0.508374f
C211 source.n40 a_n2146_n1488# 0.719262f
C212 drain_left.t14 a_n2146_n1488# 0.089068f
C213 drain_left.t6 a_n2146_n1488# 0.089068f
C214 drain_left.n0 a_n2146_n1488# 0.486594f
C215 drain_left.t7 a_n2146_n1488# 0.089068f
C216 drain_left.t12 a_n2146_n1488# 0.089068f
C217 drain_left.n1 a_n2146_n1488# 0.484515f
C218 drain_left.n2 a_n2146_n1488# 0.580693f
C219 drain_left.t9 a_n2146_n1488# 0.089068f
C220 drain_left.t3 a_n2146_n1488# 0.089068f
C221 drain_left.n3 a_n2146_n1488# 0.484515f
C222 drain_left.t19 a_n2146_n1488# 0.089068f
C223 drain_left.t2 a_n2146_n1488# 0.089068f
C224 drain_left.n4 a_n2146_n1488# 0.486594f
C225 drain_left.t10 a_n2146_n1488# 0.089068f
C226 drain_left.t0 a_n2146_n1488# 0.089068f
C227 drain_left.n5 a_n2146_n1488# 0.484515f
C228 drain_left.n6 a_n2146_n1488# 0.580694f
C229 drain_left.n7 a_n2146_n1488# 1.07179f
C230 drain_left.t8 a_n2146_n1488# 0.089068f
C231 drain_left.t17 a_n2146_n1488# 0.089068f
C232 drain_left.n8 a_n2146_n1488# 0.486596f
C233 drain_left.t13 a_n2146_n1488# 0.089068f
C234 drain_left.t11 a_n2146_n1488# 0.089068f
C235 drain_left.n9 a_n2146_n1488# 0.484517f
C236 drain_left.n10 a_n2146_n1488# 0.583973f
C237 drain_left.t18 a_n2146_n1488# 0.089068f
C238 drain_left.t16 a_n2146_n1488# 0.089068f
C239 drain_left.n11 a_n2146_n1488# 0.484517f
C240 drain_left.n12 a_n2146_n1488# 0.288032f
C241 drain_left.t1 a_n2146_n1488# 0.089068f
C242 drain_left.t4 a_n2146_n1488# 0.089068f
C243 drain_left.n13 a_n2146_n1488# 0.484517f
C244 drain_left.n14 a_n2146_n1488# 0.288032f
C245 drain_left.t15 a_n2146_n1488# 0.089068f
C246 drain_left.t5 a_n2146_n1488# 0.089068f
C247 drain_left.n15 a_n2146_n1488# 0.484517f
C248 drain_left.n16 a_n2146_n1488# 0.495109f
C249 plus.n0 a_n2146_n1488# 0.030188f
C250 plus.t16 a_n2146_n1488# 0.03934f
C251 plus.t9 a_n2146_n1488# 0.03934f
C252 plus.n1 a_n2146_n1488# 0.01048f
C253 plus.n2 a_n2146_n1488# 0.030188f
C254 plus.t17 a_n2146_n1488# 0.03934f
C255 plus.t19 a_n2146_n1488# 0.03934f
C256 plus.t11 a_n2146_n1488# 0.03934f
C257 plus.n3 a_n2146_n1488# 0.027496f
C258 plus.n4 a_n2146_n1488# 0.030188f
C259 plus.t14 a_n2146_n1488# 0.03934f
C260 plus.t18 a_n2146_n1488# 0.03934f
C261 plus.n5 a_n2146_n1488# 0.027496f
C262 plus.t10 a_n2146_n1488# 0.041722f
C263 plus.n6 a_n2146_n1488# 0.039362f
C264 plus.n7 a_n2146_n1488# 0.069637f
C265 plus.n8 a_n2146_n1488# 0.012806f
C266 plus.n9 a_n2146_n1488# 0.027496f
C267 plus.n10 a_n2146_n1488# 0.012341f
C268 plus.n11 a_n2146_n1488# 0.01048f
C269 plus.n12 a_n2146_n1488# 0.030188f
C270 plus.n13 a_n2146_n1488# 0.030188f
C271 plus.n14 a_n2146_n1488# 0.012806f
C272 plus.n15 a_n2146_n1488# 0.027496f
C273 plus.n16 a_n2146_n1488# 0.012806f
C274 plus.n17 a_n2146_n1488# 0.027496f
C275 plus.t13 a_n2146_n1488# 0.03934f
C276 plus.n18 a_n2146_n1488# 0.027496f
C277 plus.n19 a_n2146_n1488# 0.012806f
C278 plus.n20 a_n2146_n1488# 0.030188f
C279 plus.n21 a_n2146_n1488# 0.030188f
C280 plus.n22 a_n2146_n1488# 0.030188f
C281 plus.n23 a_n2146_n1488# 0.012341f
C282 plus.n24 a_n2146_n1488# 0.027496f
C283 plus.n25 a_n2146_n1488# 0.012806f
C284 plus.n26 a_n2146_n1488# 0.027496f
C285 plus.t12 a_n2146_n1488# 0.041722f
C286 plus.n27 a_n2146_n1488# 0.039316f
C287 plus.n28 a_n2146_n1488# 0.230066f
C288 plus.n29 a_n2146_n1488# 0.030188f
C289 plus.t2 a_n2146_n1488# 0.041722f
C290 plus.t6 a_n2146_n1488# 0.03934f
C291 plus.t8 a_n2146_n1488# 0.03934f
C292 plus.n30 a_n2146_n1488# 0.01048f
C293 plus.n31 a_n2146_n1488# 0.030188f
C294 plus.t15 a_n2146_n1488# 0.03934f
C295 plus.n32 a_n2146_n1488# 0.027496f
C296 plus.t0 a_n2146_n1488# 0.03934f
C297 plus.t4 a_n2146_n1488# 0.03934f
C298 plus.t5 a_n2146_n1488# 0.03934f
C299 plus.n33 a_n2146_n1488# 0.027496f
C300 plus.n34 a_n2146_n1488# 0.030188f
C301 plus.t7 a_n2146_n1488# 0.03934f
C302 plus.t1 a_n2146_n1488# 0.03934f
C303 plus.n35 a_n2146_n1488# 0.027496f
C304 plus.t3 a_n2146_n1488# 0.041722f
C305 plus.n36 a_n2146_n1488# 0.039362f
C306 plus.n37 a_n2146_n1488# 0.069637f
C307 plus.n38 a_n2146_n1488# 0.012806f
C308 plus.n39 a_n2146_n1488# 0.027496f
C309 plus.n40 a_n2146_n1488# 0.012341f
C310 plus.n41 a_n2146_n1488# 0.01048f
C311 plus.n42 a_n2146_n1488# 0.030188f
C312 plus.n43 a_n2146_n1488# 0.030188f
C313 plus.n44 a_n2146_n1488# 0.012806f
C314 plus.n45 a_n2146_n1488# 0.027496f
C315 plus.n46 a_n2146_n1488# 0.012806f
C316 plus.n47 a_n2146_n1488# 0.027496f
C317 plus.n48 a_n2146_n1488# 0.012806f
C318 plus.n49 a_n2146_n1488# 0.030188f
C319 plus.n50 a_n2146_n1488# 0.030188f
C320 plus.n51 a_n2146_n1488# 0.030188f
C321 plus.n52 a_n2146_n1488# 0.012341f
C322 plus.n53 a_n2146_n1488# 0.027496f
C323 plus.n54 a_n2146_n1488# 0.012806f
C324 plus.n55 a_n2146_n1488# 0.027496f
C325 plus.n56 a_n2146_n1488# 0.039316f
C326 plus.n57 a_n2146_n1488# 0.760157f
.ends

