* NGSPICE file created from diffpair221.ext - technology: sky130A

.subckt diffpair221 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t3 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X1 source.t2 minus.t1 drain_right.t2 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X3 source.t4 minus.t2 drain_right.t1 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X4 source.t5 plus.t0 drain_left.t3 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X5 drain_left.t2 plus.t1 source.t6 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X6 source.t7 plus.t2 drain_left.t1 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X7 a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X8 drain_right.t0 minus.t3 source.t1 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X9 drain_left.t0 plus.t3 source.t0 a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X10 a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X11 a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# a_n1334_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
R0 minus.n0 minus.t3 180.4
R1 minus.n1 minus.t1 180.4
R2 minus.n0 minus.t2 180.351
R3 minus.n1 minus.t0 180.351
R4 minus.n2 minus.n0 72.1394
R5 minus.n2 minus.n1 51.2833
R6 minus minus.n2 0.188
R7 source.n0 source.t0 69.6943
R8 source.n1 source.t5 69.6943
R9 source.n2 source.t1 69.6943
R10 source.n3 source.t4 69.6943
R11 source.n7 source.t3 69.6942
R12 source.n6 source.t2 69.6942
R13 source.n5 source.t6 69.6942
R14 source.n4 source.t7 69.6942
R15 source.n4 source.n3 15.3575
R16 source.n8 source.n0 9.65058
R17 source.n8 source.n7 5.7074
R18 source.n3 source.n2 0.888431
R19 source.n1 source.n0 0.888431
R20 source.n5 source.n4 0.888431
R21 source.n7 source.n6 0.888431
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 101.544
R26 drain_right drain_right.n1 86.3138
R27 drain_right.n0 drain_right.t2 6.6005
R28 drain_right.n0 drain_right.t3 6.6005
R29 drain_right.n1 drain_right.t1 6.6005
R30 drain_right.n1 drain_right.t0 6.6005
R31 plus.n0 plus.t0 180.4
R32 plus.n1 plus.t1 180.4
R33 plus.n0 plus.t3 180.351
R34 plus.n1 plus.t2 180.351
R35 plus plus.n1 69.4295
R36 plus plus.n0 53.5181
R37 drain_left drain_left.n0 102.097
R38 drain_left drain_left.n1 86.3138
R39 drain_left.n0 drain_left.t1 6.6005
R40 drain_left.n0 drain_left.t2 6.6005
R41 drain_left.n1 drain_left.t3 6.6005
R42 drain_left.n1 drain_left.t0 6.6005
C0 drain_left minus 0.175207f
C1 source drain_right 2.87532f
C2 minus drain_right 1.01615f
C3 source minus 1.06179f
C4 plus drain_left 1.14209f
C5 plus drain_right 0.284499f
C6 plus source 1.07579f
C7 plus minus 3.14373f
C8 drain_left drain_right 0.565395f
C9 drain_left source 2.87434f
C10 drain_right a_n1334_n1488# 3.784f
C11 drain_left a_n1334_n1488# 3.93163f
C12 source a_n1334_n1488# 3.520694f
C13 minus a_n1334_n1488# 4.298367f
C14 plus a_n1334_n1488# 5.67655f
C15 drain_left.t1 a_n1334_n1488# 0.046249f
C16 drain_left.t2 a_n1334_n1488# 0.046249f
C17 drain_left.n0 a_n1334_n1488# 0.448272f
C18 drain_left.t3 a_n1334_n1488# 0.046249f
C19 drain_left.t0 a_n1334_n1488# 0.046249f
C20 drain_left.n1 a_n1334_n1488# 0.367505f
C21 plus.t3 a_n1334_n1488# 0.208943f
C22 plus.t0 a_n1334_n1488# 0.208985f
C23 plus.n0 a_n1334_n1488# 0.254607f
C24 plus.t1 a_n1334_n1488# 0.208985f
C25 plus.t2 a_n1334_n1488# 0.208943f
C26 plus.n1 a_n1334_n1488# 0.462586f
C27 drain_right.t2 a_n1334_n1488# 0.047499f
C28 drain_right.t3 a_n1334_n1488# 0.047499f
C29 drain_right.n0 a_n1334_n1488# 0.449522f
C30 drain_right.t1 a_n1334_n1488# 0.047499f
C31 drain_right.t0 a_n1334_n1488# 0.047499f
C32 drain_right.n1 a_n1334_n1488# 0.377438f
C33 source.t0 a_n1334_n1488# 0.302468f
C34 source.n0 a_n1334_n1488# 0.442655f
C35 source.t5 a_n1334_n1488# 0.302468f
C36 source.n1 a_n1334_n1488# 0.228898f
C37 source.t1 a_n1334_n1488# 0.302468f
C38 source.n2 a_n1334_n1488# 0.228898f
C39 source.t4 a_n1334_n1488# 0.302468f
C40 source.n3 a_n1334_n1488# 0.606968f
C41 source.t7 a_n1334_n1488# 0.302466f
C42 source.n4 a_n1334_n1488# 0.60697f
C43 source.t6 a_n1334_n1488# 0.302466f
C44 source.n5 a_n1334_n1488# 0.228899f
C45 source.t2 a_n1334_n1488# 0.302466f
C46 source.n6 a_n1334_n1488# 0.228899f
C47 source.t3 a_n1334_n1488# 0.302466f
C48 source.n7 a_n1334_n1488# 0.329124f
C49 source.n8 a_n1334_n1488# 0.453088f
C50 minus.t3 a_n1334_n1488# 0.204832f
C51 minus.t2 a_n1334_n1488# 0.204791f
C52 minus.n0 a_n1334_n1488# 0.484759f
C53 minus.t1 a_n1334_n1488# 0.204832f
C54 minus.t0 a_n1334_n1488# 0.204791f
C55 minus.n1 a_n1334_n1488# 0.234845f
C56 minus.n2 a_n1334_n1488# 1.54115f
.ends

