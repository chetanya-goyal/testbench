* NGSPICE file created from diffpair527.ext - technology: sky130A

.subckt diffpair527 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t20 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X1 source.t6 plus.t0 drain_left.t15 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X2 drain_left.t14 plus.t1 source.t2 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X3 a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X4 source.t24 minus.t1 drain_right.t14 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X5 source.t14 plus.t2 drain_left.t13 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X6 source.t15 plus.t3 drain_left.t12 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X7 source.t3 plus.t4 drain_left.t11 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X8 drain_left.t10 plus.t5 source.t9 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X9 drain_right.t13 minus.t2 source.t25 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X10 a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X11 drain_right.t12 minus.t3 source.t21 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X12 source.t31 minus.t4 drain_right.t11 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X13 drain_right.t10 minus.t5 source.t23 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X14 drain_left.t9 plus.t6 source.t12 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 source.t16 minus.t6 drain_right.t9 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X16 drain_left.t8 plus.t7 source.t1 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X17 drain_left.t7 plus.t8 source.t11 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X18 source.t4 plus.t9 drain_left.t6 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 source.t17 minus.t7 drain_right.t8 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X20 source.t22 minus.t8 drain_right.t7 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X21 drain_right.t6 minus.t9 source.t18 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X22 source.t13 plus.t10 drain_left.t5 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X23 drain_right.t5 minus.t10 source.t30 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X24 drain_right.t4 minus.t11 source.t26 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X25 source.t28 minus.t12 drain_right.t3 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X26 a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X27 drain_left.t4 plus.t11 source.t0 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X28 a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X29 source.t27 minus.t13 drain_right.t2 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X30 source.t29 minus.t14 drain_right.t1 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X31 drain_right.t0 minus.t15 source.t19 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X32 source.t8 plus.t12 drain_left.t3 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X33 drain_left.t2 plus.t13 source.t10 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X34 source.t5 plus.t14 drain_left.t1 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X35 drain_left.t0 plus.t15 source.t7 a_n2210_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
R0 minus.n5 minus.t10 822.548
R1 minus.n27 minus.t4 822.548
R2 minus.n6 minus.t1 801.567
R3 minus.n8 minus.t5 801.567
R4 minus.n12 minus.t13 801.567
R5 minus.n13 minus.t2 801.567
R6 minus.n1 minus.t7 801.567
R7 minus.n19 minus.t0 801.567
R8 minus.n20 minus.t8 801.567
R9 minus.n28 minus.t3 801.567
R10 minus.n30 minus.t12 801.567
R11 minus.n34 minus.t11 801.567
R12 minus.n35 minus.t6 801.567
R13 minus.n23 minus.t15 801.567
R14 minus.n41 minus.t14 801.567
R15 minus.n42 minus.t9 801.567
R16 minus.n21 minus.n20 161.3
R17 minus.n19 minus.n0 161.3
R18 minus.n18 minus.n17 161.3
R19 minus.n16 minus.n1 161.3
R20 minus.n15 minus.n14 161.3
R21 minus.n13 minus.n2 161.3
R22 minus.n12 minus.n11 161.3
R23 minus.n10 minus.n3 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n43 minus.n42 161.3
R27 minus.n41 minus.n22 161.3
R28 minus.n40 minus.n39 161.3
R29 minus.n38 minus.n23 161.3
R30 minus.n37 minus.n36 161.3
R31 minus.n35 minus.n24 161.3
R32 minus.n34 minus.n33 161.3
R33 minus.n32 minus.n25 161.3
R34 minus.n31 minus.n30 161.3
R35 minus.n29 minus.n26 161.3
R36 minus.n5 minus.n4 70.4033
R37 minus.n27 minus.n26 70.4033
R38 minus.n13 minus.n12 48.2005
R39 minus.n20 minus.n19 48.2005
R40 minus.n35 minus.n34 48.2005
R41 minus.n42 minus.n41 48.2005
R42 minus.n44 minus.n21 39.8263
R43 minus.n8 minus.n7 37.246
R44 minus.n18 minus.n1 37.246
R45 minus.n30 minus.n29 37.246
R46 minus.n40 minus.n23 37.246
R47 minus.n8 minus.n3 35.7853
R48 minus.n14 minus.n1 35.7853
R49 minus.n30 minus.n25 35.7853
R50 minus.n36 minus.n23 35.7853
R51 minus.n6 minus.n5 20.9576
R52 minus.n28 minus.n27 20.9576
R53 minus.n12 minus.n3 12.4157
R54 minus.n14 minus.n13 12.4157
R55 minus.n34 minus.n25 12.4157
R56 minus.n36 minus.n35 12.4157
R57 minus.n7 minus.n6 10.955
R58 minus.n19 minus.n18 10.955
R59 minus.n29 minus.n28 10.955
R60 minus.n41 minus.n40 10.955
R61 minus.n44 minus.n43 6.56111
R62 minus.n21 minus.n0 0.189894
R63 minus.n17 minus.n0 0.189894
R64 minus.n17 minus.n16 0.189894
R65 minus.n16 minus.n15 0.189894
R66 minus.n15 minus.n2 0.189894
R67 minus.n11 minus.n2 0.189894
R68 minus.n11 minus.n10 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n31 minus.n26 0.189894
R72 minus.n32 minus.n31 0.189894
R73 minus.n33 minus.n32 0.189894
R74 minus.n33 minus.n24 0.189894
R75 minus.n37 minus.n24 0.189894
R76 minus.n38 minus.n37 0.189894
R77 minus.n39 minus.n38 0.189894
R78 minus.n39 minus.n22 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 source.n7 source.t15 45.521
R82 source.n8 source.t30 45.521
R83 source.n15 source.t22 45.521
R84 source.n31 source.t18 45.5208
R85 source.n24 source.t31 45.5208
R86 source.n23 source.t2 45.5208
R87 source.n16 source.t14 45.5208
R88 source.n0 source.t10 45.5208
R89 source.n2 source.n1 44.201
R90 source.n4 source.n3 44.201
R91 source.n6 source.n5 44.201
R92 source.n10 source.n9 44.201
R93 source.n12 source.n11 44.201
R94 source.n14 source.n13 44.201
R95 source.n30 source.n29 44.2008
R96 source.n28 source.n27 44.2008
R97 source.n26 source.n25 44.2008
R98 source.n22 source.n21 44.2008
R99 source.n20 source.n19 44.2008
R100 source.n18 source.n17 44.2008
R101 source.n16 source.n15 24.276
R102 source.n32 source.n0 18.6553
R103 source.n32 source.n31 5.62119
R104 source.n29 source.t19 1.3205
R105 source.n29 source.t29 1.3205
R106 source.n27 source.t26 1.3205
R107 source.n27 source.t16 1.3205
R108 source.n25 source.t21 1.3205
R109 source.n25 source.t28 1.3205
R110 source.n21 source.t11 1.3205
R111 source.n21 source.t6 1.3205
R112 source.n19 source.t9 1.3205
R113 source.n19 source.t3 1.3205
R114 source.n17 source.t1 1.3205
R115 source.n17 source.t13 1.3205
R116 source.n1 source.t7 1.3205
R117 source.n1 source.t4 1.3205
R118 source.n3 source.t12 1.3205
R119 source.n3 source.t8 1.3205
R120 source.n5 source.t0 1.3205
R121 source.n5 source.t5 1.3205
R122 source.n9 source.t23 1.3205
R123 source.n9 source.t24 1.3205
R124 source.n11 source.t25 1.3205
R125 source.n11 source.t27 1.3205
R126 source.n13 source.t20 1.3205
R127 source.n13 source.t17 1.3205
R128 source.n15 source.n14 0.716017
R129 source.n14 source.n12 0.716017
R130 source.n12 source.n10 0.716017
R131 source.n10 source.n8 0.716017
R132 source.n7 source.n6 0.716017
R133 source.n6 source.n4 0.716017
R134 source.n4 source.n2 0.716017
R135 source.n2 source.n0 0.716017
R136 source.n18 source.n16 0.716017
R137 source.n20 source.n18 0.716017
R138 source.n22 source.n20 0.716017
R139 source.n23 source.n22 0.716017
R140 source.n26 source.n24 0.716017
R141 source.n28 source.n26 0.716017
R142 source.n30 source.n28 0.716017
R143 source.n31 source.n30 0.716017
R144 source.n8 source.n7 0.470328
R145 source.n24 source.n23 0.470328
R146 source source.n32 0.188
R147 drain_right.n9 drain_right.n7 61.5952
R148 drain_right.n5 drain_right.n3 61.5951
R149 drain_right.n2 drain_right.n0 61.5951
R150 drain_right.n9 drain_right.n8 60.8798
R151 drain_right.n11 drain_right.n10 60.8798
R152 drain_right.n13 drain_right.n12 60.8798
R153 drain_right.n5 drain_right.n4 60.8796
R154 drain_right.n2 drain_right.n1 60.8796
R155 drain_right drain_right.n6 33.7374
R156 drain_right drain_right.n13 6.36873
R157 drain_right.n3 drain_right.t1 1.3205
R158 drain_right.n3 drain_right.t6 1.3205
R159 drain_right.n4 drain_right.t9 1.3205
R160 drain_right.n4 drain_right.t0 1.3205
R161 drain_right.n1 drain_right.t3 1.3205
R162 drain_right.n1 drain_right.t4 1.3205
R163 drain_right.n0 drain_right.t11 1.3205
R164 drain_right.n0 drain_right.t12 1.3205
R165 drain_right.n7 drain_right.t14 1.3205
R166 drain_right.n7 drain_right.t5 1.3205
R167 drain_right.n8 drain_right.t2 1.3205
R168 drain_right.n8 drain_right.t10 1.3205
R169 drain_right.n10 drain_right.t8 1.3205
R170 drain_right.n10 drain_right.t13 1.3205
R171 drain_right.n12 drain_right.t7 1.3205
R172 drain_right.n12 drain_right.t15 1.3205
R173 drain_right.n13 drain_right.n11 0.716017
R174 drain_right.n11 drain_right.n9 0.716017
R175 drain_right.n6 drain_right.n5 0.302913
R176 drain_right.n6 drain_right.n2 0.302913
R177 plus.n5 plus.t3 822.548
R178 plus.n27 plus.t1 822.548
R179 plus.n20 plus.t13 801.567
R180 plus.n19 plus.t9 801.567
R181 plus.n1 plus.t15 801.567
R182 plus.n13 plus.t12 801.567
R183 plus.n12 plus.t6 801.567
R184 plus.n4 plus.t14 801.567
R185 plus.n6 plus.t11 801.567
R186 plus.n42 plus.t2 801.567
R187 plus.n41 plus.t7 801.567
R188 plus.n23 plus.t10 801.567
R189 plus.n35 plus.t5 801.567
R190 plus.n34 plus.t4 801.567
R191 plus.n26 plus.t8 801.567
R192 plus.n28 plus.t0 801.567
R193 plus.n8 plus.n7 161.3
R194 plus.n9 plus.n4 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n12 plus.n3 161.3
R197 plus.n13 plus.n2 161.3
R198 plus.n15 plus.n14 161.3
R199 plus.n16 plus.n1 161.3
R200 plus.n18 plus.n17 161.3
R201 plus.n19 plus.n0 161.3
R202 plus.n21 plus.n20 161.3
R203 plus.n30 plus.n29 161.3
R204 plus.n31 plus.n26 161.3
R205 plus.n33 plus.n32 161.3
R206 plus.n34 plus.n25 161.3
R207 plus.n35 plus.n24 161.3
R208 plus.n37 plus.n36 161.3
R209 plus.n38 plus.n23 161.3
R210 plus.n40 plus.n39 161.3
R211 plus.n41 plus.n22 161.3
R212 plus.n43 plus.n42 161.3
R213 plus.n8 plus.n5 70.4033
R214 plus.n30 plus.n27 70.4033
R215 plus.n20 plus.n19 48.2005
R216 plus.n13 plus.n12 48.2005
R217 plus.n42 plus.n41 48.2005
R218 plus.n35 plus.n34 48.2005
R219 plus.n18 plus.n1 37.246
R220 plus.n7 plus.n4 37.246
R221 plus.n40 plus.n23 37.246
R222 plus.n29 plus.n26 37.246
R223 plus.n14 plus.n1 35.7853
R224 plus.n11 plus.n4 35.7853
R225 plus.n36 plus.n23 35.7853
R226 plus.n33 plus.n26 35.7853
R227 plus plus.n43 32.571
R228 plus.n6 plus.n5 20.9576
R229 plus.n28 plus.n27 20.9576
R230 plus plus.n21 13.3414
R231 plus.n14 plus.n13 12.4157
R232 plus.n12 plus.n11 12.4157
R233 plus.n36 plus.n35 12.4157
R234 plus.n34 plus.n33 12.4157
R235 plus.n19 plus.n18 10.955
R236 plus.n7 plus.n6 10.955
R237 plus.n41 plus.n40 10.955
R238 plus.n29 plus.n28 10.955
R239 plus.n9 plus.n8 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n3 0.189894
R242 plus.n3 plus.n2 0.189894
R243 plus.n15 plus.n2 0.189894
R244 plus.n16 plus.n15 0.189894
R245 plus.n17 plus.n16 0.189894
R246 plus.n17 plus.n0 0.189894
R247 plus.n21 plus.n0 0.189894
R248 plus.n43 plus.n22 0.189894
R249 plus.n39 plus.n22 0.189894
R250 plus.n39 plus.n38 0.189894
R251 plus.n38 plus.n37 0.189894
R252 plus.n37 plus.n24 0.189894
R253 plus.n25 plus.n24 0.189894
R254 plus.n32 plus.n25 0.189894
R255 plus.n32 plus.n31 0.189894
R256 plus.n31 plus.n30 0.189894
R257 drain_left.n9 drain_left.n7 61.5953
R258 drain_left.n5 drain_left.n3 61.5951
R259 drain_left.n2 drain_left.n0 61.5951
R260 drain_left.n11 drain_left.n10 60.8798
R261 drain_left.n9 drain_left.n8 60.8798
R262 drain_left.n13 drain_left.n12 60.8796
R263 drain_left.n5 drain_left.n4 60.8796
R264 drain_left.n2 drain_left.n1 60.8796
R265 drain_left drain_left.n6 34.2907
R266 drain_left drain_left.n13 6.36873
R267 drain_left.n3 drain_left.t15 1.3205
R268 drain_left.n3 drain_left.t14 1.3205
R269 drain_left.n4 drain_left.t11 1.3205
R270 drain_left.n4 drain_left.t7 1.3205
R271 drain_left.n1 drain_left.t5 1.3205
R272 drain_left.n1 drain_left.t10 1.3205
R273 drain_left.n0 drain_left.t13 1.3205
R274 drain_left.n0 drain_left.t8 1.3205
R275 drain_left.n12 drain_left.t6 1.3205
R276 drain_left.n12 drain_left.t2 1.3205
R277 drain_left.n10 drain_left.t3 1.3205
R278 drain_left.n10 drain_left.t0 1.3205
R279 drain_left.n8 drain_left.t1 1.3205
R280 drain_left.n8 drain_left.t9 1.3205
R281 drain_left.n7 drain_left.t12 1.3205
R282 drain_left.n7 drain_left.t4 1.3205
R283 drain_left.n11 drain_left.n9 0.716017
R284 drain_left.n13 drain_left.n11 0.716017
R285 drain_left.n6 drain_left.n5 0.302913
R286 drain_left.n6 drain_left.n2 0.302913
C0 source drain_left 28.632801f
C1 drain_right plus 0.372806f
C2 minus plus 6.46219f
C3 drain_right minus 10.3135f
C4 plus drain_left 10.5307f
C5 plus source 10.087f
C6 drain_right drain_left 1.15071f
C7 drain_right source 28.633999f
C8 minus drain_left 0.172419f
C9 minus source 10.073f
C10 drain_right a_n2210_n3888# 7.15129f
C11 drain_left a_n2210_n3888# 7.47272f
C12 source a_n2210_n3888# 10.651047f
C13 minus a_n2210_n3888# 8.94237f
C14 plus a_n2210_n3888# 10.97665f
C15 drain_left.t13 a_n2210_n3888# 0.348154f
C16 drain_left.t8 a_n2210_n3888# 0.348154f
C17 drain_left.n0 a_n2210_n3888# 3.15141f
C18 drain_left.t5 a_n2210_n3888# 0.348154f
C19 drain_left.t10 a_n2210_n3888# 0.348154f
C20 drain_left.n1 a_n2210_n3888# 3.1469f
C21 drain_left.n2 a_n2210_n3888# 0.722491f
C22 drain_left.t15 a_n2210_n3888# 0.348154f
C23 drain_left.t14 a_n2210_n3888# 0.348154f
C24 drain_left.n3 a_n2210_n3888# 3.15141f
C25 drain_left.t11 a_n2210_n3888# 0.348154f
C26 drain_left.t7 a_n2210_n3888# 0.348154f
C27 drain_left.n4 a_n2210_n3888# 3.1469f
C28 drain_left.n5 a_n2210_n3888# 0.722491f
C29 drain_left.n6 a_n2210_n3888# 1.77314f
C30 drain_left.t12 a_n2210_n3888# 0.348154f
C31 drain_left.t4 a_n2210_n3888# 0.348154f
C32 drain_left.n7 a_n2210_n3888# 3.15141f
C33 drain_left.t1 a_n2210_n3888# 0.348154f
C34 drain_left.t9 a_n2210_n3888# 0.348154f
C35 drain_left.n8 a_n2210_n3888# 3.1469f
C36 drain_left.n9 a_n2210_n3888# 0.759331f
C37 drain_left.t3 a_n2210_n3888# 0.348154f
C38 drain_left.t0 a_n2210_n3888# 0.348154f
C39 drain_left.n10 a_n2210_n3888# 3.1469f
C40 drain_left.n11 a_n2210_n3888# 0.376003f
C41 drain_left.t6 a_n2210_n3888# 0.348154f
C42 drain_left.t2 a_n2210_n3888# 0.348154f
C43 drain_left.n12 a_n2210_n3888# 3.14689f
C44 drain_left.n13 a_n2210_n3888# 0.628356f
C45 plus.n0 a_n2210_n3888# 0.045598f
C46 plus.t13 a_n2210_n3888# 0.971818f
C47 plus.t9 a_n2210_n3888# 0.971818f
C48 plus.t15 a_n2210_n3888# 0.971818f
C49 plus.n1 a_n2210_n3888# 0.383365f
C50 plus.n2 a_n2210_n3888# 0.045598f
C51 plus.t12 a_n2210_n3888# 0.971818f
C52 plus.t6 a_n2210_n3888# 0.971818f
C53 plus.n3 a_n2210_n3888# 0.045598f
C54 plus.t14 a_n2210_n3888# 0.971818f
C55 plus.n4 a_n2210_n3888# 0.383365f
C56 plus.t3 a_n2210_n3888# 0.981477f
C57 plus.n5 a_n2210_n3888# 0.36926f
C58 plus.t11 a_n2210_n3888# 0.971818f
C59 plus.n6 a_n2210_n3888# 0.380694f
C60 plus.n7 a_n2210_n3888# 0.010347f
C61 plus.n8 a_n2210_n3888# 0.145177f
C62 plus.n9 a_n2210_n3888# 0.045598f
C63 plus.n10 a_n2210_n3888# 0.045598f
C64 plus.n11 a_n2210_n3888# 0.010347f
C65 plus.n12 a_n2210_n3888# 0.380975f
C66 plus.n13 a_n2210_n3888# 0.380975f
C67 plus.n14 a_n2210_n3888# 0.010347f
C68 plus.n15 a_n2210_n3888# 0.045598f
C69 plus.n16 a_n2210_n3888# 0.045598f
C70 plus.n17 a_n2210_n3888# 0.045598f
C71 plus.n18 a_n2210_n3888# 0.010347f
C72 plus.n19 a_n2210_n3888# 0.380694f
C73 plus.n20 a_n2210_n3888# 0.378586f
C74 plus.n21 a_n2210_n3888# 0.582768f
C75 plus.n22 a_n2210_n3888# 0.045598f
C76 plus.t2 a_n2210_n3888# 0.971818f
C77 plus.t7 a_n2210_n3888# 0.971818f
C78 plus.t10 a_n2210_n3888# 0.971818f
C79 plus.n23 a_n2210_n3888# 0.383365f
C80 plus.n24 a_n2210_n3888# 0.045598f
C81 plus.t5 a_n2210_n3888# 0.971818f
C82 plus.n25 a_n2210_n3888# 0.045598f
C83 plus.t4 a_n2210_n3888# 0.971818f
C84 plus.t8 a_n2210_n3888# 0.971818f
C85 plus.n26 a_n2210_n3888# 0.383365f
C86 plus.t1 a_n2210_n3888# 0.981477f
C87 plus.n27 a_n2210_n3888# 0.36926f
C88 plus.t0 a_n2210_n3888# 0.971818f
C89 plus.n28 a_n2210_n3888# 0.380694f
C90 plus.n29 a_n2210_n3888# 0.010347f
C91 plus.n30 a_n2210_n3888# 0.145177f
C92 plus.n31 a_n2210_n3888# 0.045598f
C93 plus.n32 a_n2210_n3888# 0.045598f
C94 plus.n33 a_n2210_n3888# 0.010347f
C95 plus.n34 a_n2210_n3888# 0.380975f
C96 plus.n35 a_n2210_n3888# 0.380975f
C97 plus.n36 a_n2210_n3888# 0.010347f
C98 plus.n37 a_n2210_n3888# 0.045598f
C99 plus.n38 a_n2210_n3888# 0.045598f
C100 plus.n39 a_n2210_n3888# 0.045598f
C101 plus.n40 a_n2210_n3888# 0.010347f
C102 plus.n41 a_n2210_n3888# 0.380694f
C103 plus.n42 a_n2210_n3888# 0.378586f
C104 plus.n43 a_n2210_n3888# 1.5442f
C105 drain_right.t11 a_n2210_n3888# 0.347394f
C106 drain_right.t12 a_n2210_n3888# 0.347394f
C107 drain_right.n0 a_n2210_n3888# 3.14453f
C108 drain_right.t3 a_n2210_n3888# 0.347394f
C109 drain_right.t4 a_n2210_n3888# 0.347394f
C110 drain_right.n1 a_n2210_n3888# 3.14003f
C111 drain_right.n2 a_n2210_n3888# 0.720914f
C112 drain_right.t1 a_n2210_n3888# 0.347394f
C113 drain_right.t6 a_n2210_n3888# 0.347394f
C114 drain_right.n3 a_n2210_n3888# 3.14453f
C115 drain_right.t9 a_n2210_n3888# 0.347394f
C116 drain_right.t0 a_n2210_n3888# 0.347394f
C117 drain_right.n4 a_n2210_n3888# 3.14003f
C118 drain_right.n5 a_n2210_n3888# 0.720914f
C119 drain_right.n6 a_n2210_n3888# 1.70863f
C120 drain_right.t14 a_n2210_n3888# 0.347394f
C121 drain_right.t5 a_n2210_n3888# 0.347394f
C122 drain_right.n7 a_n2210_n3888# 3.14452f
C123 drain_right.t2 a_n2210_n3888# 0.347394f
C124 drain_right.t10 a_n2210_n3888# 0.347394f
C125 drain_right.n8 a_n2210_n3888# 3.14003f
C126 drain_right.n9 a_n2210_n3888# 0.757684f
C127 drain_right.t8 a_n2210_n3888# 0.347394f
C128 drain_right.t13 a_n2210_n3888# 0.347394f
C129 drain_right.n10 a_n2210_n3888# 3.14003f
C130 drain_right.n11 a_n2210_n3888# 0.375182f
C131 drain_right.t7 a_n2210_n3888# 0.347394f
C132 drain_right.t15 a_n2210_n3888# 0.347394f
C133 drain_right.n12 a_n2210_n3888# 3.14003f
C134 drain_right.n13 a_n2210_n3888# 0.626973f
C135 source.t10 a_n2210_n3888# 3.25493f
C136 source.n0 a_n2210_n3888# 1.52957f
C137 source.t7 a_n2210_n3888# 0.290448f
C138 source.t4 a_n2210_n3888# 0.290448f
C139 source.n1 a_n2210_n3888# 2.55134f
C140 source.n2 a_n2210_n3888# 0.354347f
C141 source.t12 a_n2210_n3888# 0.290448f
C142 source.t8 a_n2210_n3888# 0.290448f
C143 source.n3 a_n2210_n3888# 2.55134f
C144 source.n4 a_n2210_n3888# 0.354347f
C145 source.t0 a_n2210_n3888# 0.290448f
C146 source.t5 a_n2210_n3888# 0.290448f
C147 source.n5 a_n2210_n3888# 2.55134f
C148 source.n6 a_n2210_n3888# 0.354347f
C149 source.t15 a_n2210_n3888# 3.25494f
C150 source.n7 a_n2210_n3888# 0.423479f
C151 source.t30 a_n2210_n3888# 3.25494f
C152 source.n8 a_n2210_n3888# 0.423479f
C153 source.t23 a_n2210_n3888# 0.290448f
C154 source.t24 a_n2210_n3888# 0.290448f
C155 source.n9 a_n2210_n3888# 2.55134f
C156 source.n10 a_n2210_n3888# 0.354347f
C157 source.t25 a_n2210_n3888# 0.290448f
C158 source.t27 a_n2210_n3888# 0.290448f
C159 source.n11 a_n2210_n3888# 2.55134f
C160 source.n12 a_n2210_n3888# 0.354347f
C161 source.t20 a_n2210_n3888# 0.290448f
C162 source.t17 a_n2210_n3888# 0.290448f
C163 source.n13 a_n2210_n3888# 2.55134f
C164 source.n14 a_n2210_n3888# 0.354347f
C165 source.t22 a_n2210_n3888# 3.25494f
C166 source.n15 a_n2210_n3888# 1.94223f
C167 source.t14 a_n2210_n3888# 3.25493f
C168 source.n16 a_n2210_n3888# 1.94224f
C169 source.t1 a_n2210_n3888# 0.290448f
C170 source.t13 a_n2210_n3888# 0.290448f
C171 source.n17 a_n2210_n3888# 2.55134f
C172 source.n18 a_n2210_n3888# 0.35435f
C173 source.t9 a_n2210_n3888# 0.290448f
C174 source.t3 a_n2210_n3888# 0.290448f
C175 source.n19 a_n2210_n3888# 2.55134f
C176 source.n20 a_n2210_n3888# 0.35435f
C177 source.t11 a_n2210_n3888# 0.290448f
C178 source.t6 a_n2210_n3888# 0.290448f
C179 source.n21 a_n2210_n3888# 2.55134f
C180 source.n22 a_n2210_n3888# 0.35435f
C181 source.t2 a_n2210_n3888# 3.25493f
C182 source.n23 a_n2210_n3888# 0.423483f
C183 source.t31 a_n2210_n3888# 3.25493f
C184 source.n24 a_n2210_n3888# 0.423483f
C185 source.t21 a_n2210_n3888# 0.290448f
C186 source.t28 a_n2210_n3888# 0.290448f
C187 source.n25 a_n2210_n3888# 2.55134f
C188 source.n26 a_n2210_n3888# 0.35435f
C189 source.t26 a_n2210_n3888# 0.290448f
C190 source.t16 a_n2210_n3888# 0.290448f
C191 source.n27 a_n2210_n3888# 2.55134f
C192 source.n28 a_n2210_n3888# 0.35435f
C193 source.t19 a_n2210_n3888# 0.290448f
C194 source.t29 a_n2210_n3888# 0.290448f
C195 source.n29 a_n2210_n3888# 2.55134f
C196 source.n30 a_n2210_n3888# 0.35435f
C197 source.t18 a_n2210_n3888# 3.25493f
C198 source.n31 a_n2210_n3888# 0.572622f
C199 source.n32 a_n2210_n3888# 1.79971f
C200 minus.n0 a_n2210_n3888# 0.045108f
C201 minus.t7 a_n2210_n3888# 0.961375f
C202 minus.n1 a_n2210_n3888# 0.379245f
C203 minus.n2 a_n2210_n3888# 0.045108f
C204 minus.n3 a_n2210_n3888# 0.010236f
C205 minus.t13 a_n2210_n3888# 0.961375f
C206 minus.n4 a_n2210_n3888# 0.143616f
C207 minus.t1 a_n2210_n3888# 0.961375f
C208 minus.t10 a_n2210_n3888# 0.97093f
C209 minus.n5 a_n2210_n3888# 0.365291f
C210 minus.n6 a_n2210_n3888# 0.376603f
C211 minus.n7 a_n2210_n3888# 0.010236f
C212 minus.t5 a_n2210_n3888# 0.961375f
C213 minus.n8 a_n2210_n3888# 0.379245f
C214 minus.n9 a_n2210_n3888# 0.045108f
C215 minus.n10 a_n2210_n3888# 0.045108f
C216 minus.n11 a_n2210_n3888# 0.045108f
C217 minus.n12 a_n2210_n3888# 0.376882f
C218 minus.t2 a_n2210_n3888# 0.961375f
C219 minus.n13 a_n2210_n3888# 0.376882f
C220 minus.n14 a_n2210_n3888# 0.010236f
C221 minus.n15 a_n2210_n3888# 0.045108f
C222 minus.n16 a_n2210_n3888# 0.045108f
C223 minus.n17 a_n2210_n3888# 0.045108f
C224 minus.n18 a_n2210_n3888# 0.010236f
C225 minus.t0 a_n2210_n3888# 0.961375f
C226 minus.n19 a_n2210_n3888# 0.376603f
C227 minus.t8 a_n2210_n3888# 0.961375f
C228 minus.n20 a_n2210_n3888# 0.374518f
C229 minus.n21 a_n2210_n3888# 1.84776f
C230 minus.n22 a_n2210_n3888# 0.045108f
C231 minus.t15 a_n2210_n3888# 0.961375f
C232 minus.n23 a_n2210_n3888# 0.379245f
C233 minus.n24 a_n2210_n3888# 0.045108f
C234 minus.n25 a_n2210_n3888# 0.010236f
C235 minus.n26 a_n2210_n3888# 0.143616f
C236 minus.t4 a_n2210_n3888# 0.97093f
C237 minus.n27 a_n2210_n3888# 0.365291f
C238 minus.t3 a_n2210_n3888# 0.961375f
C239 minus.n28 a_n2210_n3888# 0.376603f
C240 minus.n29 a_n2210_n3888# 0.010236f
C241 minus.t12 a_n2210_n3888# 0.961375f
C242 minus.n30 a_n2210_n3888# 0.379245f
C243 minus.n31 a_n2210_n3888# 0.045108f
C244 minus.n32 a_n2210_n3888# 0.045108f
C245 minus.n33 a_n2210_n3888# 0.045108f
C246 minus.t11 a_n2210_n3888# 0.961375f
C247 minus.n34 a_n2210_n3888# 0.376882f
C248 minus.t6 a_n2210_n3888# 0.961375f
C249 minus.n35 a_n2210_n3888# 0.376882f
C250 minus.n36 a_n2210_n3888# 0.010236f
C251 minus.n37 a_n2210_n3888# 0.045108f
C252 minus.n38 a_n2210_n3888# 0.045108f
C253 minus.n39 a_n2210_n3888# 0.045108f
C254 minus.n40 a_n2210_n3888# 0.010236f
C255 minus.t14 a_n2210_n3888# 0.961375f
C256 minus.n41 a_n2210_n3888# 0.376603f
C257 minus.t9 a_n2210_n3888# 0.961375f
C258 minus.n42 a_n2210_n3888# 0.374518f
C259 minus.n43 a_n2210_n3888# 0.301379f
C260 minus.n44 a_n2210_n3888# 2.21875f
.ends

