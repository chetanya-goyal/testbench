* NGSPICE file created from diffpair377.ext - technology: sky130A

.subckt diffpair377 minus drain_right drain_left source plus
X0 a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X1 drain_left.t15 plus.t0 source.t22 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X2 source.t15 plus.t1 drain_left.t14 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X3 drain_left.t13 plus.t2 source.t21 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 source.t1 minus.t0 drain_right.t15 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X6 source.t13 minus.t1 drain_right.t14 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X7 drain_right.t13 minus.t2 source.t2 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X8 drain_right.t12 minus.t3 source.t7 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X9 source.t30 plus.t3 drain_left.t12 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 source.t10 minus.t4 drain_right.t11 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 source.t3 minus.t5 drain_right.t10 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X12 source.t12 minus.t6 drain_right.t9 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X13 source.t29 plus.t4 drain_left.t11 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X14 drain_left.t10 plus.t5 source.t16 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X15 drain_left.t9 plus.t6 source.t17 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X16 source.t6 minus.t7 drain_right.t8 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X17 drain_right.t7 minus.t8 source.t8 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X18 a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X19 drain_left.t8 plus.t7 source.t26 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X20 source.t11 minus.t9 drain_right.t6 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X21 source.t23 plus.t8 drain_left.t7 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X22 drain_right.t5 minus.t10 source.t5 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X23 drain_right.t4 minus.t11 source.t14 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X24 drain_left.t6 plus.t9 source.t28 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X25 source.t25 plus.t10 drain_left.t5 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X26 a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X27 drain_right.t3 minus.t12 source.t31 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X28 drain_left.t4 plus.t11 source.t18 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X29 source.t27 plus.t12 drain_left.t3 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X30 source.t19 plus.t13 drain_left.t2 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X31 drain_right.t2 minus.t13 source.t9 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X32 drain_left.t1 plus.t14 source.t24 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X33 source.t0 minus.t14 drain_right.t1 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X34 drain_right.t0 minus.t15 source.t4 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X35 source.t20 plus.t15 drain_left.t0 a_n2390_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
R0 plus.n6 plus.t10 447.954
R1 plus.n30 plus.t11 447.954
R2 plus.n22 plus.t0 426.973
R3 plus.n21 plus.t1 426.973
R4 plus.n1 plus.t2 426.973
R5 plus.n15 plus.t4 426.973
R6 plus.n3 plus.t7 426.973
R7 plus.n9 plus.t8 426.973
R8 plus.n5 plus.t9 426.973
R9 plus.n46 plus.t13 426.973
R10 plus.n45 plus.t6 426.973
R11 plus.n25 plus.t15 426.973
R12 plus.n39 plus.t14 426.973
R13 plus.n27 plus.t12 426.973
R14 plus.n33 plus.t5 426.973
R15 plus.n29 plus.t3 426.973
R16 plus.n8 plus.n7 161.3
R17 plus.n9 plus.n4 161.3
R18 plus.n11 plus.n10 161.3
R19 plus.n12 plus.n3 161.3
R20 plus.n14 plus.n13 161.3
R21 plus.n15 plus.n2 161.3
R22 plus.n17 plus.n16 161.3
R23 plus.n18 plus.n1 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n21 plus.n0 161.3
R26 plus.n23 plus.n22 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n33 plus.n28 161.3
R29 plus.n35 plus.n34 161.3
R30 plus.n36 plus.n27 161.3
R31 plus.n38 plus.n37 161.3
R32 plus.n39 plus.n26 161.3
R33 plus.n41 plus.n40 161.3
R34 plus.n42 plus.n25 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n45 plus.n24 161.3
R37 plus.n47 plus.n46 161.3
R38 plus.n7 plus.n6 70.4033
R39 plus.n31 plus.n30 70.4033
R40 plus.n22 plus.n21 48.2005
R41 plus.n46 plus.n45 48.2005
R42 plus.n20 plus.n1 44.549
R43 plus.n9 plus.n8 44.549
R44 plus.n44 plus.n25 44.549
R45 plus.n33 plus.n32 44.549
R46 plus.n16 plus.n15 34.3247
R47 plus.n10 plus.n3 34.3247
R48 plus.n40 plus.n39 34.3247
R49 plus.n34 plus.n27 34.3247
R50 plus plus.n47 31.0748
R51 plus.n14 plus.n3 24.1005
R52 plus.n15 plus.n14 24.1005
R53 plus.n39 plus.n38 24.1005
R54 plus.n38 plus.n27 24.1005
R55 plus.n6 plus.n5 20.9576
R56 plus.n30 plus.n29 20.9576
R57 plus.n16 plus.n1 13.8763
R58 plus.n10 plus.n9 13.8763
R59 plus.n40 plus.n25 13.8763
R60 plus.n34 plus.n33 13.8763
R61 plus plus.n23 11.1634
R62 plus.n21 plus.n20 3.65202
R63 plus.n8 plus.n5 3.65202
R64 plus.n45 plus.n44 3.65202
R65 plus.n32 plus.n29 3.65202
R66 plus.n7 plus.n4 0.189894
R67 plus.n11 plus.n4 0.189894
R68 plus.n12 plus.n11 0.189894
R69 plus.n13 plus.n12 0.189894
R70 plus.n13 plus.n2 0.189894
R71 plus.n17 plus.n2 0.189894
R72 plus.n18 plus.n17 0.189894
R73 plus.n19 plus.n18 0.189894
R74 plus.n19 plus.n0 0.189894
R75 plus.n23 plus.n0 0.189894
R76 plus.n47 plus.n24 0.189894
R77 plus.n43 plus.n24 0.189894
R78 plus.n43 plus.n42 0.189894
R79 plus.n42 plus.n41 0.189894
R80 plus.n41 plus.n26 0.189894
R81 plus.n37 plus.n26 0.189894
R82 plus.n37 plus.n36 0.189894
R83 plus.n36 plus.n35 0.189894
R84 plus.n35 plus.n28 0.189894
R85 plus.n31 plus.n28 0.189894
R86 source.n7 source.t25 51.0588
R87 source.n8 source.t5 51.0588
R88 source.n15 source.t1 51.0588
R89 source.n31 source.t14 51.0586
R90 source.n24 source.t12 51.0586
R91 source.n23 source.t18 51.0586
R92 source.n16 source.t19 51.0586
R93 source.n0 source.t22 51.0586
R94 source.n2 source.n1 48.8588
R95 source.n4 source.n3 48.8588
R96 source.n6 source.n5 48.8588
R97 source.n10 source.n9 48.8588
R98 source.n12 source.n11 48.8588
R99 source.n14 source.n13 48.8588
R100 source.n30 source.n29 48.8586
R101 source.n28 source.n27 48.8586
R102 source.n26 source.n25 48.8586
R103 source.n22 source.n21 48.8586
R104 source.n20 source.n19 48.8586
R105 source.n18 source.n17 48.8586
R106 source.n16 source.n15 19.8167
R107 source.n32 source.n0 14.1529
R108 source.n32 source.n31 5.66429
R109 source.n29 source.t9 2.2005
R110 source.n29 source.t3 2.2005
R111 source.n27 source.t31 2.2005
R112 source.n27 source.t0 2.2005
R113 source.n25 source.t4 2.2005
R114 source.n25 source.t13 2.2005
R115 source.n21 source.t16 2.2005
R116 source.n21 source.t30 2.2005
R117 source.n19 source.t24 2.2005
R118 source.n19 source.t27 2.2005
R119 source.n17 source.t17 2.2005
R120 source.n17 source.t20 2.2005
R121 source.n1 source.t21 2.2005
R122 source.n1 source.t15 2.2005
R123 source.n3 source.t26 2.2005
R124 source.n3 source.t29 2.2005
R125 source.n5 source.t28 2.2005
R126 source.n5 source.t23 2.2005
R127 source.n9 source.t8 2.2005
R128 source.n9 source.t11 2.2005
R129 source.n11 source.t2 2.2005
R130 source.n11 source.t6 2.2005
R131 source.n13 source.t7 2.2005
R132 source.n13 source.t10 2.2005
R133 source.n15 source.n14 0.802224
R134 source.n14 source.n12 0.802224
R135 source.n12 source.n10 0.802224
R136 source.n10 source.n8 0.802224
R137 source.n7 source.n6 0.802224
R138 source.n6 source.n4 0.802224
R139 source.n4 source.n2 0.802224
R140 source.n2 source.n0 0.802224
R141 source.n18 source.n16 0.802224
R142 source.n20 source.n18 0.802224
R143 source.n22 source.n20 0.802224
R144 source.n23 source.n22 0.802224
R145 source.n26 source.n24 0.802224
R146 source.n28 source.n26 0.802224
R147 source.n30 source.n28 0.802224
R148 source.n31 source.n30 0.802224
R149 source.n8 source.n7 0.470328
R150 source.n24 source.n23 0.470328
R151 source source.n32 0.188
R152 drain_left.n9 drain_left.n7 66.3393
R153 drain_left.n5 drain_left.n3 66.3391
R154 drain_left.n2 drain_left.n0 66.3391
R155 drain_left.n11 drain_left.n10 65.5376
R156 drain_left.n9 drain_left.n8 65.5376
R157 drain_left.n13 drain_left.n12 65.5374
R158 drain_left.n5 drain_left.n4 65.5373
R159 drain_left.n2 drain_left.n1 65.5373
R160 drain_left drain_left.n6 30.3056
R161 drain_left drain_left.n13 6.45494
R162 drain_left.n3 drain_left.t12 2.2005
R163 drain_left.n3 drain_left.t4 2.2005
R164 drain_left.n4 drain_left.t3 2.2005
R165 drain_left.n4 drain_left.t10 2.2005
R166 drain_left.n1 drain_left.t0 2.2005
R167 drain_left.n1 drain_left.t1 2.2005
R168 drain_left.n0 drain_left.t2 2.2005
R169 drain_left.n0 drain_left.t9 2.2005
R170 drain_left.n12 drain_left.t14 2.2005
R171 drain_left.n12 drain_left.t15 2.2005
R172 drain_left.n10 drain_left.t11 2.2005
R173 drain_left.n10 drain_left.t13 2.2005
R174 drain_left.n8 drain_left.t7 2.2005
R175 drain_left.n8 drain_left.t8 2.2005
R176 drain_left.n7 drain_left.t5 2.2005
R177 drain_left.n7 drain_left.t6 2.2005
R178 drain_left.n11 drain_left.n9 0.802224
R179 drain_left.n13 drain_left.n11 0.802224
R180 drain_left.n6 drain_left.n5 0.346016
R181 drain_left.n6 drain_left.n2 0.346016
R182 minus.n6 minus.t10 447.954
R183 minus.n30 minus.t6 447.954
R184 minus.n5 minus.t9 426.973
R185 minus.n9 minus.t8 426.973
R186 minus.n3 minus.t7 426.973
R187 minus.n15 minus.t2 426.973
R188 minus.n1 minus.t4 426.973
R189 minus.n21 minus.t3 426.973
R190 minus.n22 minus.t0 426.973
R191 minus.n29 minus.t15 426.973
R192 minus.n33 minus.t1 426.973
R193 minus.n27 minus.t12 426.973
R194 minus.n39 minus.t14 426.973
R195 minus.n25 minus.t13 426.973
R196 minus.n45 minus.t5 426.973
R197 minus.n46 minus.t11 426.973
R198 minus.n23 minus.n22 161.3
R199 minus.n21 minus.n0 161.3
R200 minus.n20 minus.n19 161.3
R201 minus.n18 minus.n1 161.3
R202 minus.n17 minus.n16 161.3
R203 minus.n15 minus.n2 161.3
R204 minus.n14 minus.n13 161.3
R205 minus.n12 minus.n3 161.3
R206 minus.n11 minus.n10 161.3
R207 minus.n9 minus.n4 161.3
R208 minus.n8 minus.n7 161.3
R209 minus.n47 minus.n46 161.3
R210 minus.n45 minus.n24 161.3
R211 minus.n44 minus.n43 161.3
R212 minus.n42 minus.n25 161.3
R213 minus.n41 minus.n40 161.3
R214 minus.n39 minus.n26 161.3
R215 minus.n38 minus.n37 161.3
R216 minus.n36 minus.n27 161.3
R217 minus.n35 minus.n34 161.3
R218 minus.n33 minus.n28 161.3
R219 minus.n32 minus.n31 161.3
R220 minus.n7 minus.n6 70.4033
R221 minus.n31 minus.n30 70.4033
R222 minus.n22 minus.n21 48.2005
R223 minus.n46 minus.n45 48.2005
R224 minus.n9 minus.n8 44.549
R225 minus.n20 minus.n1 44.549
R226 minus.n33 minus.n32 44.549
R227 minus.n44 minus.n25 44.549
R228 minus.n48 minus.n23 36.0573
R229 minus.n10 minus.n3 34.3247
R230 minus.n16 minus.n15 34.3247
R231 minus.n34 minus.n27 34.3247
R232 minus.n40 minus.n39 34.3247
R233 minus.n15 minus.n14 24.1005
R234 minus.n14 minus.n3 24.1005
R235 minus.n38 minus.n27 24.1005
R236 minus.n39 minus.n38 24.1005
R237 minus.n6 minus.n5 20.9576
R238 minus.n30 minus.n29 20.9576
R239 minus.n10 minus.n9 13.8763
R240 minus.n16 minus.n1 13.8763
R241 minus.n34 minus.n33 13.8763
R242 minus.n40 minus.n25 13.8763
R243 minus.n48 minus.n47 6.6558
R244 minus.n8 minus.n5 3.65202
R245 minus.n21 minus.n20 3.65202
R246 minus.n32 minus.n29 3.65202
R247 minus.n45 minus.n44 3.65202
R248 minus.n23 minus.n0 0.189894
R249 minus.n19 minus.n0 0.189894
R250 minus.n19 minus.n18 0.189894
R251 minus.n18 minus.n17 0.189894
R252 minus.n17 minus.n2 0.189894
R253 minus.n13 minus.n2 0.189894
R254 minus.n13 minus.n12 0.189894
R255 minus.n12 minus.n11 0.189894
R256 minus.n11 minus.n4 0.189894
R257 minus.n7 minus.n4 0.189894
R258 minus.n31 minus.n28 0.189894
R259 minus.n35 minus.n28 0.189894
R260 minus.n36 minus.n35 0.189894
R261 minus.n37 minus.n36 0.189894
R262 minus.n37 minus.n26 0.189894
R263 minus.n41 minus.n26 0.189894
R264 minus.n42 minus.n41 0.189894
R265 minus.n43 minus.n42 0.189894
R266 minus.n43 minus.n24 0.189894
R267 minus.n47 minus.n24 0.189894
R268 minus minus.n48 0.188
R269 drain_right.n9 drain_right.n7 66.3391
R270 drain_right.n5 drain_right.n3 66.3391
R271 drain_right.n2 drain_right.n0 66.3391
R272 drain_right.n9 drain_right.n8 65.5376
R273 drain_right.n11 drain_right.n10 65.5376
R274 drain_right.n13 drain_right.n12 65.5376
R275 drain_right.n5 drain_right.n4 65.5373
R276 drain_right.n2 drain_right.n1 65.5373
R277 drain_right drain_right.n6 29.7523
R278 drain_right drain_right.n13 6.45494
R279 drain_right.n3 drain_right.t10 2.2005
R280 drain_right.n3 drain_right.t4 2.2005
R281 drain_right.n4 drain_right.t1 2.2005
R282 drain_right.n4 drain_right.t2 2.2005
R283 drain_right.n1 drain_right.t14 2.2005
R284 drain_right.n1 drain_right.t3 2.2005
R285 drain_right.n0 drain_right.t9 2.2005
R286 drain_right.n0 drain_right.t0 2.2005
R287 drain_right.n7 drain_right.t6 2.2005
R288 drain_right.n7 drain_right.t5 2.2005
R289 drain_right.n8 drain_right.t8 2.2005
R290 drain_right.n8 drain_right.t7 2.2005
R291 drain_right.n10 drain_right.t11 2.2005
R292 drain_right.n10 drain_right.t13 2.2005
R293 drain_right.n12 drain_right.t15 2.2005
R294 drain_right.n12 drain_right.t12 2.2005
R295 drain_right.n13 drain_right.n11 0.802224
R296 drain_right.n11 drain_right.n9 0.802224
R297 drain_right.n6 drain_right.n5 0.346016
R298 drain_right.n6 drain_right.n2 0.346016
C0 source minus 7.23524f
C1 drain_right minus 7.16065f
C2 source plus 7.24928f
C3 drain_right plus 0.391974f
C4 drain_left source 16.8791f
C5 drain_left drain_right 1.24373f
C6 plus minus 5.56869f
C7 source drain_right 16.8808f
C8 drain_left minus 0.172752f
C9 drain_left plus 7.39655f
C10 drain_right a_n2390_n2688# 6.0974f
C11 drain_left a_n2390_n2688# 6.4397f
C12 source a_n2390_n2688# 7.476986f
C13 minus a_n2390_n2688# 9.281727f
C14 plus a_n2390_n2688# 10.93406f
C15 drain_right.t9 a_n2390_n2688# 0.199088f
C16 drain_right.t0 a_n2390_n2688# 0.199088f
C17 drain_right.n0 a_n2390_n2688# 1.74595f
C18 drain_right.t14 a_n2390_n2688# 0.199088f
C19 drain_right.t3 a_n2390_n2688# 0.199088f
C20 drain_right.n1 a_n2390_n2688# 1.74135f
C21 drain_right.n2 a_n2390_n2688# 0.705123f
C22 drain_right.t10 a_n2390_n2688# 0.199088f
C23 drain_right.t4 a_n2390_n2688# 0.199088f
C24 drain_right.n3 a_n2390_n2688# 1.74595f
C25 drain_right.t1 a_n2390_n2688# 0.199088f
C26 drain_right.t2 a_n2390_n2688# 0.199088f
C27 drain_right.n4 a_n2390_n2688# 1.74135f
C28 drain_right.n5 a_n2390_n2688# 0.705123f
C29 drain_right.n6 a_n2390_n2688# 1.30185f
C30 drain_right.t6 a_n2390_n2688# 0.199088f
C31 drain_right.t5 a_n2390_n2688# 0.199088f
C32 drain_right.n7 a_n2390_n2688# 1.74594f
C33 drain_right.t8 a_n2390_n2688# 0.199088f
C34 drain_right.t7 a_n2390_n2688# 0.199088f
C35 drain_right.n8 a_n2390_n2688# 1.74136f
C36 drain_right.n9 a_n2390_n2688# 0.744395f
C37 drain_right.t11 a_n2390_n2688# 0.199088f
C38 drain_right.t13 a_n2390_n2688# 0.199088f
C39 drain_right.n10 a_n2390_n2688# 1.74136f
C40 drain_right.n11 a_n2390_n2688# 0.368853f
C41 drain_right.t15 a_n2390_n2688# 0.199088f
C42 drain_right.t12 a_n2390_n2688# 0.199088f
C43 drain_right.n12 a_n2390_n2688# 1.74136f
C44 drain_right.n13 a_n2390_n2688# 0.612949f
C45 minus.n0 a_n2390_n2688# 0.042954f
C46 minus.t4 a_n2390_n2688# 0.6652f
C47 minus.n1 a_n2390_n2688# 0.283411f
C48 minus.n2 a_n2390_n2688# 0.042954f
C49 minus.t7 a_n2390_n2688# 0.6652f
C50 minus.n3 a_n2390_n2688# 0.283411f
C51 minus.n4 a_n2390_n2688# 0.042954f
C52 minus.t9 a_n2390_n2688# 0.6652f
C53 minus.n5 a_n2390_n2688# 0.282219f
C54 minus.t10 a_n2390_n2688# 0.678391f
C55 minus.n6 a_n2390_n2688# 0.26871f
C56 minus.n7 a_n2390_n2688# 0.144672f
C57 minus.n8 a_n2390_n2688# 0.009747f
C58 minus.t8 a_n2390_n2688# 0.6652f
C59 minus.n9 a_n2390_n2688# 0.283411f
C60 minus.n10 a_n2390_n2688# 0.009747f
C61 minus.n11 a_n2390_n2688# 0.042954f
C62 minus.n12 a_n2390_n2688# 0.042954f
C63 minus.n13 a_n2390_n2688# 0.042954f
C64 minus.n14 a_n2390_n2688# 0.009747f
C65 minus.t2 a_n2390_n2688# 0.6652f
C66 minus.n15 a_n2390_n2688# 0.283411f
C67 minus.n16 a_n2390_n2688# 0.009747f
C68 minus.n17 a_n2390_n2688# 0.042954f
C69 minus.n18 a_n2390_n2688# 0.042954f
C70 minus.n19 a_n2390_n2688# 0.042954f
C71 minus.n20 a_n2390_n2688# 0.009747f
C72 minus.t3 a_n2390_n2688# 0.6652f
C73 minus.n21 a_n2390_n2688# 0.282219f
C74 minus.t0 a_n2390_n2688# 0.6652f
C75 minus.n22 a_n2390_n2688# 0.281557f
C76 minus.n23 a_n2390_n2688# 1.51427f
C77 minus.n24 a_n2390_n2688# 0.042954f
C78 minus.t13 a_n2390_n2688# 0.6652f
C79 minus.n25 a_n2390_n2688# 0.283411f
C80 minus.n26 a_n2390_n2688# 0.042954f
C81 minus.t12 a_n2390_n2688# 0.6652f
C82 minus.n27 a_n2390_n2688# 0.283411f
C83 minus.n28 a_n2390_n2688# 0.042954f
C84 minus.t15 a_n2390_n2688# 0.6652f
C85 minus.n29 a_n2390_n2688# 0.282219f
C86 minus.t6 a_n2390_n2688# 0.678391f
C87 minus.n30 a_n2390_n2688# 0.26871f
C88 minus.n31 a_n2390_n2688# 0.144672f
C89 minus.n32 a_n2390_n2688# 0.009747f
C90 minus.t1 a_n2390_n2688# 0.6652f
C91 minus.n33 a_n2390_n2688# 0.283411f
C92 minus.n34 a_n2390_n2688# 0.009747f
C93 minus.n35 a_n2390_n2688# 0.042954f
C94 minus.n36 a_n2390_n2688# 0.042954f
C95 minus.n37 a_n2390_n2688# 0.042954f
C96 minus.n38 a_n2390_n2688# 0.009747f
C97 minus.t14 a_n2390_n2688# 0.6652f
C98 minus.n39 a_n2390_n2688# 0.283411f
C99 minus.n40 a_n2390_n2688# 0.009747f
C100 minus.n41 a_n2390_n2688# 0.042954f
C101 minus.n42 a_n2390_n2688# 0.042954f
C102 minus.n43 a_n2390_n2688# 0.042954f
C103 minus.n44 a_n2390_n2688# 0.009747f
C104 minus.t5 a_n2390_n2688# 0.6652f
C105 minus.n45 a_n2390_n2688# 0.282219f
C106 minus.t11 a_n2390_n2688# 0.6652f
C107 minus.n46 a_n2390_n2688# 0.281557f
C108 minus.n47 a_n2390_n2688# 0.296473f
C109 minus.n48 a_n2390_n2688# 1.83479f
C110 drain_left.t2 a_n2390_n2688# 0.199832f
C111 drain_left.t9 a_n2390_n2688# 0.199832f
C112 drain_left.n0 a_n2390_n2688# 1.75247f
C113 drain_left.t0 a_n2390_n2688# 0.199832f
C114 drain_left.t1 a_n2390_n2688# 0.199832f
C115 drain_left.n1 a_n2390_n2688# 1.74786f
C116 drain_left.n2 a_n2390_n2688# 0.707759f
C117 drain_left.t12 a_n2390_n2688# 0.199832f
C118 drain_left.t4 a_n2390_n2688# 0.199832f
C119 drain_left.n3 a_n2390_n2688# 1.75247f
C120 drain_left.t3 a_n2390_n2688# 0.199832f
C121 drain_left.t10 a_n2390_n2688# 0.199832f
C122 drain_left.n4 a_n2390_n2688# 1.74786f
C123 drain_left.n5 a_n2390_n2688# 0.707759f
C124 drain_left.n6 a_n2390_n2688# 1.36402f
C125 drain_left.t5 a_n2390_n2688# 0.199832f
C126 drain_left.t6 a_n2390_n2688# 0.199832f
C127 drain_left.n7 a_n2390_n2688# 1.75248f
C128 drain_left.t7 a_n2390_n2688# 0.199832f
C129 drain_left.t8 a_n2390_n2688# 0.199832f
C130 drain_left.n8 a_n2390_n2688# 1.74787f
C131 drain_left.n9 a_n2390_n2688# 0.74717f
C132 drain_left.t11 a_n2390_n2688# 0.199832f
C133 drain_left.t13 a_n2390_n2688# 0.199832f
C134 drain_left.n10 a_n2390_n2688# 1.74787f
C135 drain_left.n11 a_n2390_n2688# 0.370232f
C136 drain_left.t14 a_n2390_n2688# 0.199832f
C137 drain_left.t15 a_n2390_n2688# 0.199832f
C138 drain_left.n12 a_n2390_n2688# 1.74786f
C139 drain_left.n13 a_n2390_n2688# 0.615248f
C140 source.t22 a_n2390_n2688# 1.8524f
C141 source.n0 a_n2390_n2688# 1.09922f
C142 source.t21 a_n2390_n2688# 0.173714f
C143 source.t15 a_n2390_n2688# 0.173714f
C144 source.n1 a_n2390_n2688# 1.45422f
C145 source.n2 a_n2390_n2688# 0.353845f
C146 source.t26 a_n2390_n2688# 0.173714f
C147 source.t29 a_n2390_n2688# 0.173714f
C148 source.n3 a_n2390_n2688# 1.45422f
C149 source.n4 a_n2390_n2688# 0.353845f
C150 source.t28 a_n2390_n2688# 0.173714f
C151 source.t23 a_n2390_n2688# 0.173714f
C152 source.n5 a_n2390_n2688# 1.45422f
C153 source.n6 a_n2390_n2688# 0.353845f
C154 source.t25 a_n2390_n2688# 1.8524f
C155 source.n7 a_n2390_n2688# 0.403311f
C156 source.t5 a_n2390_n2688# 1.8524f
C157 source.n8 a_n2390_n2688# 0.403311f
C158 source.t8 a_n2390_n2688# 0.173714f
C159 source.t11 a_n2390_n2688# 0.173714f
C160 source.n9 a_n2390_n2688# 1.45422f
C161 source.n10 a_n2390_n2688# 0.353845f
C162 source.t2 a_n2390_n2688# 0.173714f
C163 source.t6 a_n2390_n2688# 0.173714f
C164 source.n11 a_n2390_n2688# 1.45422f
C165 source.n12 a_n2390_n2688# 0.353845f
C166 source.t7 a_n2390_n2688# 0.173714f
C167 source.t10 a_n2390_n2688# 0.173714f
C168 source.n13 a_n2390_n2688# 1.45422f
C169 source.n14 a_n2390_n2688# 0.353845f
C170 source.t1 a_n2390_n2688# 1.8524f
C171 source.n15 a_n2390_n2688# 1.46078f
C172 source.t19 a_n2390_n2688# 1.8524f
C173 source.n16 a_n2390_n2688# 1.46079f
C174 source.t17 a_n2390_n2688# 0.173714f
C175 source.t20 a_n2390_n2688# 0.173714f
C176 source.n17 a_n2390_n2688# 1.45422f
C177 source.n18 a_n2390_n2688# 0.353849f
C178 source.t24 a_n2390_n2688# 0.173714f
C179 source.t27 a_n2390_n2688# 0.173714f
C180 source.n19 a_n2390_n2688# 1.45422f
C181 source.n20 a_n2390_n2688# 0.353849f
C182 source.t16 a_n2390_n2688# 0.173714f
C183 source.t30 a_n2390_n2688# 0.173714f
C184 source.n21 a_n2390_n2688# 1.45422f
C185 source.n22 a_n2390_n2688# 0.353849f
C186 source.t18 a_n2390_n2688# 1.8524f
C187 source.n23 a_n2390_n2688# 0.403316f
C188 source.t12 a_n2390_n2688# 1.8524f
C189 source.n24 a_n2390_n2688# 0.403316f
C190 source.t4 a_n2390_n2688# 0.173714f
C191 source.t13 a_n2390_n2688# 0.173714f
C192 source.n25 a_n2390_n2688# 1.45422f
C193 source.n26 a_n2390_n2688# 0.353849f
C194 source.t31 a_n2390_n2688# 0.173714f
C195 source.t0 a_n2390_n2688# 0.173714f
C196 source.n27 a_n2390_n2688# 1.45422f
C197 source.n28 a_n2390_n2688# 0.353849f
C198 source.t9 a_n2390_n2688# 0.173714f
C199 source.t3 a_n2390_n2688# 0.173714f
C200 source.n29 a_n2390_n2688# 1.45422f
C201 source.n30 a_n2390_n2688# 0.353849f
C202 source.t14 a_n2390_n2688# 1.8524f
C203 source.n31 a_n2390_n2688# 0.557326f
C204 source.n32 a_n2390_n2688# 1.2824f
C205 plus.n0 a_n2390_n2688# 0.043573f
C206 plus.t0 a_n2390_n2688# 0.674783f
C207 plus.t1 a_n2390_n2688# 0.674783f
C208 plus.t2 a_n2390_n2688# 0.674783f
C209 plus.n1 a_n2390_n2688# 0.287494f
C210 plus.n2 a_n2390_n2688# 0.043573f
C211 plus.t4 a_n2390_n2688# 0.674783f
C212 plus.t7 a_n2390_n2688# 0.674783f
C213 plus.n3 a_n2390_n2688# 0.287494f
C214 plus.n4 a_n2390_n2688# 0.043573f
C215 plus.t8 a_n2390_n2688# 0.674783f
C216 plus.t9 a_n2390_n2688# 0.674783f
C217 plus.n5 a_n2390_n2688# 0.286285f
C218 plus.t10 a_n2390_n2688# 0.688164f
C219 plus.n6 a_n2390_n2688# 0.272581f
C220 plus.n7 a_n2390_n2688# 0.146756f
C221 plus.n8 a_n2390_n2688# 0.009887f
C222 plus.n9 a_n2390_n2688# 0.287494f
C223 plus.n10 a_n2390_n2688# 0.009887f
C224 plus.n11 a_n2390_n2688# 0.043573f
C225 plus.n12 a_n2390_n2688# 0.043573f
C226 plus.n13 a_n2390_n2688# 0.043573f
C227 plus.n14 a_n2390_n2688# 0.009887f
C228 plus.n15 a_n2390_n2688# 0.287494f
C229 plus.n16 a_n2390_n2688# 0.009887f
C230 plus.n17 a_n2390_n2688# 0.043573f
C231 plus.n18 a_n2390_n2688# 0.043573f
C232 plus.n19 a_n2390_n2688# 0.043573f
C233 plus.n20 a_n2390_n2688# 0.009887f
C234 plus.n21 a_n2390_n2688# 0.286285f
C235 plus.n22 a_n2390_n2688# 0.285613f
C236 plus.n23 a_n2390_n2688# 0.444404f
C237 plus.n24 a_n2390_n2688# 0.043573f
C238 plus.t13 a_n2390_n2688# 0.674783f
C239 plus.t6 a_n2390_n2688# 0.674783f
C240 plus.t15 a_n2390_n2688# 0.674783f
C241 plus.n25 a_n2390_n2688# 0.287494f
C242 plus.n26 a_n2390_n2688# 0.043573f
C243 plus.t14 a_n2390_n2688# 0.674783f
C244 plus.t12 a_n2390_n2688# 0.674783f
C245 plus.n27 a_n2390_n2688# 0.287494f
C246 plus.n28 a_n2390_n2688# 0.043573f
C247 plus.t5 a_n2390_n2688# 0.674783f
C248 plus.t3 a_n2390_n2688# 0.674783f
C249 plus.n29 a_n2390_n2688# 0.286285f
C250 plus.t11 a_n2390_n2688# 0.688164f
C251 plus.n30 a_n2390_n2688# 0.272581f
C252 plus.n31 a_n2390_n2688# 0.146756f
C253 plus.n32 a_n2390_n2688# 0.009887f
C254 plus.n33 a_n2390_n2688# 0.287494f
C255 plus.n34 a_n2390_n2688# 0.009887f
C256 plus.n35 a_n2390_n2688# 0.043573f
C257 plus.n36 a_n2390_n2688# 0.043573f
C258 plus.n37 a_n2390_n2688# 0.043573f
C259 plus.n38 a_n2390_n2688# 0.009887f
C260 plus.n39 a_n2390_n2688# 0.287494f
C261 plus.n40 a_n2390_n2688# 0.009887f
C262 plus.n41 a_n2390_n2688# 0.043573f
C263 plus.n42 a_n2390_n2688# 0.043573f
C264 plus.n43 a_n2390_n2688# 0.043573f
C265 plus.n44 a_n2390_n2688# 0.009887f
C266 plus.n45 a_n2390_n2688# 0.286285f
C267 plus.n46 a_n2390_n2688# 0.285613f
C268 plus.n47 a_n2390_n2688# 1.34566f
.ends

