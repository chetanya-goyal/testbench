* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X1 drain_left.t5 plus.t0 source.t4 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X2 source.t1 minus.t0 drain_right.t5 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 drain_left.t4 plus.t1 source.t9 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X4 drain_left.t3 plus.t2 source.t8 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X5 a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X6 drain_right.t4 minus.t1 source.t2 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X7 a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X8 a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X9 source.t3 minus.t2 drain_right.t3 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X10 drain_right.t2 minus.t3 source.t0 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X11 drain_right.t1 minus.t4 source.t10 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X12 source.t7 plus.t3 drain_left.t2 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 drain_right.t0 minus.t5 source.t11 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X14 source.t6 plus.t4 drain_left.t1 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X15 drain_left.t0 plus.t5 source.t5 a_n1540_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
R0 plus.n3 plus.n0 161.3
R1 plus.n5 plus.n4 161.3
R2 plus.n9 plus.n6 161.3
R3 plus.n11 plus.n10 161.3
R4 plus.n1 plus.t2 146.571
R5 plus.n7 plus.t5 146.571
R6 plus.n4 plus.t0 124.977
R7 plus.n2 plus.t3 124.977
R8 plus.n10 plus.t1 124.977
R9 plus.n8 plus.t4 124.977
R10 plus.n1 plus.n0 44.8545
R11 plus.n7 plus.n6 44.8545
R12 plus.n4 plus.n3 26.2914
R13 plus.n10 plus.n9 26.2914
R14 plus plus.n11 25.1752
R15 plus.n3 plus.n2 21.9096
R16 plus.n9 plus.n8 21.9096
R17 plus.n2 plus.n1 20.3348
R18 plus.n8 plus.n7 20.3348
R19 plus plus.n5 8.48345
R20 plus.n5 plus.n0 0.189894
R21 plus.n11 plus.n6 0.189894
R22 source.n34 source.n32 289.615
R23 source.n24 source.n22 289.615
R24 source.n2 source.n0 289.615
R25 source.n12 source.n10 289.615
R26 source.n35 source.n34 185
R27 source.n25 source.n24 185
R28 source.n3 source.n2 185
R29 source.n13 source.n12 185
R30 source.t11 source.n33 167.117
R31 source.t5 source.n23 167.117
R32 source.t4 source.n1 167.117
R33 source.t0 source.n11 167.117
R34 source.n9 source.n8 84.1169
R35 source.n19 source.n18 84.1169
R36 source.n31 source.n30 84.1168
R37 source.n21 source.n20 84.1168
R38 source.n34 source.t11 52.3082
R39 source.n24 source.t5 52.3082
R40 source.n2 source.t4 52.3082
R41 source.n12 source.t0 52.3082
R42 source.n39 source.n38 31.4096
R43 source.n29 source.n28 31.4096
R44 source.n7 source.n6 31.4096
R45 source.n17 source.n16 31.4096
R46 source.n21 source.n19 15.4878
R47 source.n30 source.t10 9.9005
R48 source.n30 source.t3 9.9005
R49 source.n20 source.t9 9.9005
R50 source.n20 source.t6 9.9005
R51 source.n8 source.t8 9.9005
R52 source.n8 source.t7 9.9005
R53 source.n18 source.t2 9.9005
R54 source.n18 source.t1 9.9005
R55 source.n35 source.n33 9.71174
R56 source.n25 source.n23 9.71174
R57 source.n3 source.n1 9.71174
R58 source.n13 source.n11 9.71174
R59 source.n38 source.n37 9.45567
R60 source.n28 source.n27 9.45567
R61 source.n6 source.n5 9.45567
R62 source.n16 source.n15 9.45567
R63 source.n37 source.n36 9.3005
R64 source.n27 source.n26 9.3005
R65 source.n5 source.n4 9.3005
R66 source.n15 source.n14 9.3005
R67 source.n40 source.n7 8.893
R68 source.n38 source.n32 8.14595
R69 source.n28 source.n22 8.14595
R70 source.n6 source.n0 8.14595
R71 source.n16 source.n10 8.14595
R72 source.n36 source.n35 7.3702
R73 source.n26 source.n25 7.3702
R74 source.n4 source.n3 7.3702
R75 source.n14 source.n13 7.3702
R76 source.n36 source.n32 5.81868
R77 source.n26 source.n22 5.81868
R78 source.n4 source.n0 5.81868
R79 source.n14 source.n10 5.81868
R80 source.n40 source.n39 5.7074
R81 source.n37 source.n33 3.44771
R82 source.n27 source.n23 3.44771
R83 source.n5 source.n1 3.44771
R84 source.n15 source.n11 3.44771
R85 source.n17 source.n9 0.914293
R86 source.n31 source.n29 0.914293
R87 source.n19 source.n17 0.888431
R88 source.n9 source.n7 0.888431
R89 source.n29 source.n21 0.888431
R90 source.n39 source.n31 0.888431
R91 source source.n40 0.188
R92 drain_left.n2 drain_left.n0 289.615
R93 drain_left.n11 drain_left.n9 289.615
R94 drain_left.n3 drain_left.n2 185
R95 drain_left.n12 drain_left.n11 185
R96 drain_left.t4 drain_left.n1 167.117
R97 drain_left.t3 drain_left.n10 167.117
R98 drain_left.n8 drain_left.n7 100.963
R99 drain_left.n17 drain_left.n16 100.796
R100 drain_left.n2 drain_left.t4 52.3082
R101 drain_left.n11 drain_left.t3 52.3082
R102 drain_left.n17 drain_left.n15 48.9763
R103 drain_left.n8 drain_left.n6 48.699
R104 drain_left drain_left.n8 22.2331
R105 drain_left.n7 drain_left.t1 9.9005
R106 drain_left.n7 drain_left.t0 9.9005
R107 drain_left.n16 drain_left.t2 9.9005
R108 drain_left.n16 drain_left.t5 9.9005
R109 drain_left.n3 drain_left.n1 9.71174
R110 drain_left.n12 drain_left.n10 9.71174
R111 drain_left.n6 drain_left.n5 9.45567
R112 drain_left.n15 drain_left.n14 9.45567
R113 drain_left.n5 drain_left.n4 9.3005
R114 drain_left.n14 drain_left.n13 9.3005
R115 drain_left.n6 drain_left.n0 8.14595
R116 drain_left.n15 drain_left.n9 8.14595
R117 drain_left.n4 drain_left.n3 7.3702
R118 drain_left.n13 drain_left.n12 7.3702
R119 drain_left drain_left.n17 6.54115
R120 drain_left.n4 drain_left.n0 5.81868
R121 drain_left.n13 drain_left.n9 5.81868
R122 drain_left.n5 drain_left.n1 3.44771
R123 drain_left.n14 drain_left.n10 3.44771
R124 minus.n5 minus.n4 161.3
R125 minus.n3 minus.n0 161.3
R126 minus.n11 minus.n10 161.3
R127 minus.n9 minus.n6 161.3
R128 minus.n1 minus.t3 146.571
R129 minus.n7 minus.t4 146.571
R130 minus.n2 minus.t0 124.977
R131 minus.n4 minus.t1 124.977
R132 minus.n8 minus.t2 124.977
R133 minus.n10 minus.t5 124.977
R134 minus.n1 minus.n0 44.8545
R135 minus.n7 minus.n6 44.8545
R136 minus.n12 minus.n5 27.5062
R137 minus.n4 minus.n3 26.2914
R138 minus.n10 minus.n9 26.2914
R139 minus.n3 minus.n2 21.9096
R140 minus.n9 minus.n8 21.9096
R141 minus.n2 minus.n1 20.3348
R142 minus.n8 minus.n7 20.3348
R143 minus.n12 minus.n11 6.62739
R144 minus.n5 minus.n0 0.189894
R145 minus.n11 minus.n6 0.189894
R146 minus minus.n12 0.188
R147 drain_right.n2 drain_right.n0 289.615
R148 drain_right.n12 drain_right.n10 289.615
R149 drain_right.n3 drain_right.n2 185
R150 drain_right.n13 drain_right.n12 185
R151 drain_right.t1 drain_right.n1 167.117
R152 drain_right.t4 drain_right.n11 167.117
R153 drain_right.n17 drain_right.n9 101.683
R154 drain_right.n8 drain_right.n7 100.963
R155 drain_right.n2 drain_right.t1 52.3082
R156 drain_right.n12 drain_right.t4 52.3082
R157 drain_right.n8 drain_right.n6 48.699
R158 drain_right.n17 drain_right.n16 48.0884
R159 drain_right drain_right.n8 21.6799
R160 drain_right.n7 drain_right.t3 9.9005
R161 drain_right.n7 drain_right.t0 9.9005
R162 drain_right.n9 drain_right.t5 9.9005
R163 drain_right.n9 drain_right.t2 9.9005
R164 drain_right.n3 drain_right.n1 9.71174
R165 drain_right.n13 drain_right.n11 9.71174
R166 drain_right.n6 drain_right.n5 9.45567
R167 drain_right.n16 drain_right.n15 9.45567
R168 drain_right.n5 drain_right.n4 9.3005
R169 drain_right.n15 drain_right.n14 9.3005
R170 drain_right.n6 drain_right.n0 8.14595
R171 drain_right.n16 drain_right.n10 8.14595
R172 drain_right.n4 drain_right.n3 7.3702
R173 drain_right.n14 drain_right.n13 7.3702
R174 drain_right drain_right.n17 6.09718
R175 drain_right.n4 drain_right.n0 5.81868
R176 drain_right.n14 drain_right.n10 5.81868
R177 drain_right.n5 drain_right.n1 3.44771
R178 drain_right.n15 drain_right.n11 3.44771
C0 source drain_right 3.2832f
C1 drain_left drain_right 0.705446f
C2 source plus 1.22652f
C3 drain_left plus 1.15941f
C4 source minus 1.21248f
C5 drain_left minus 0.17749f
C6 drain_right plus 0.308856f
C7 drain_right minus 1.01246f
C8 source drain_left 3.28387f
C9 plus minus 3.21739f
C10 drain_right a_n1540_n1288# 3.227851f
C11 drain_left a_n1540_n1288# 3.430266f
C12 source a_n1540_n1288# 2.480082f
C13 minus a_n1540_n1288# 5.080446f
C14 plus a_n1540_n1288# 5.679356f
C15 drain_right.n0 a_n1540_n1288# 0.02608f
C16 drain_right.n1 a_n1540_n1288# 0.057704f
C17 drain_right.t1 a_n1540_n1288# 0.043304f
C18 drain_right.n2 a_n1540_n1288# 0.045162f
C19 drain_right.n3 a_n1540_n1288# 0.014558f
C20 drain_right.n4 a_n1540_n1288# 0.009602f
C21 drain_right.n5 a_n1540_n1288# 0.127194f
C22 drain_right.n6 a_n1540_n1288# 0.041808f
C23 drain_right.t3 a_n1540_n1288# 0.02824f
C24 drain_right.t0 a_n1540_n1288# 0.02824f
C25 drain_right.n7 a_n1540_n1288# 0.177753f
C26 drain_right.n8 a_n1540_n1288# 0.712567f
C27 drain_right.t5 a_n1540_n1288# 0.02824f
C28 drain_right.t2 a_n1540_n1288# 0.02824f
C29 drain_right.n9 a_n1540_n1288# 0.179561f
C30 drain_right.n10 a_n1540_n1288# 0.02608f
C31 drain_right.n11 a_n1540_n1288# 0.057704f
C32 drain_right.t4 a_n1540_n1288# 0.043304f
C33 drain_right.n12 a_n1540_n1288# 0.045162f
C34 drain_right.n13 a_n1540_n1288# 0.014558f
C35 drain_right.n14 a_n1540_n1288# 0.009602f
C36 drain_right.n15 a_n1540_n1288# 0.127194f
C37 drain_right.n16 a_n1540_n1288# 0.040935f
C38 drain_right.n17 a_n1540_n1288# 0.493239f
C39 minus.n0 a_n1540_n1288# 0.11976f
C40 minus.t3 a_n1540_n1288# 0.138224f
C41 minus.n1 a_n1540_n1288# 0.077025f
C42 minus.t0 a_n1540_n1288# 0.125408f
C43 minus.n2 a_n1540_n1288# 0.089517f
C44 minus.n3 a_n1540_n1288# 0.006564f
C45 minus.t1 a_n1540_n1288# 0.125408f
C46 minus.n4 a_n1540_n1288# 0.085035f
C47 minus.n5 a_n1540_n1288# 0.650387f
C48 minus.n6 a_n1540_n1288# 0.11976f
C49 minus.t4 a_n1540_n1288# 0.138224f
C50 minus.n7 a_n1540_n1288# 0.077025f
C51 minus.t2 a_n1540_n1288# 0.125408f
C52 minus.n8 a_n1540_n1288# 0.089517f
C53 minus.n9 a_n1540_n1288# 0.006564f
C54 minus.t5 a_n1540_n1288# 0.125408f
C55 minus.n10 a_n1540_n1288# 0.085035f
C56 minus.n11 a_n1540_n1288# 0.197744f
C57 minus.n12 a_n1540_n1288# 0.79899f
C58 drain_left.n0 a_n1540_n1288# 0.025539f
C59 drain_left.n1 a_n1540_n1288# 0.056507f
C60 drain_left.t4 a_n1540_n1288# 0.042406f
C61 drain_left.n2 a_n1540_n1288# 0.044225f
C62 drain_left.n3 a_n1540_n1288# 0.014256f
C63 drain_left.n4 a_n1540_n1288# 0.009402f
C64 drain_left.n5 a_n1540_n1288# 0.124556f
C65 drain_left.n6 a_n1540_n1288# 0.040941f
C66 drain_left.t1 a_n1540_n1288# 0.027654f
C67 drain_left.t0 a_n1540_n1288# 0.027654f
C68 drain_left.n7 a_n1540_n1288# 0.174066f
C69 drain_left.n8 a_n1540_n1288# 0.732181f
C70 drain_left.n9 a_n1540_n1288# 0.025539f
C71 drain_left.n10 a_n1540_n1288# 0.056507f
C72 drain_left.t3 a_n1540_n1288# 0.042406f
C73 drain_left.n11 a_n1540_n1288# 0.044225f
C74 drain_left.n12 a_n1540_n1288# 0.014256f
C75 drain_left.n13 a_n1540_n1288# 0.009402f
C76 drain_left.n14 a_n1540_n1288# 0.124556f
C77 drain_left.n15 a_n1540_n1288# 0.041594f
C78 drain_left.t2 a_n1540_n1288# 0.027654f
C79 drain_left.t5 a_n1540_n1288# 0.027654f
C80 drain_left.n16 a_n1540_n1288# 0.173732f
C81 drain_left.n17 a_n1540_n1288# 0.470512f
C82 source.n0 a_n1540_n1288# 0.032733f
C83 source.n1 a_n1540_n1288# 0.072425f
C84 source.t4 a_n1540_n1288# 0.054352f
C85 source.n2 a_n1540_n1288# 0.056683f
C86 source.n3 a_n1540_n1288# 0.018272f
C87 source.n4 a_n1540_n1288# 0.012051f
C88 source.n5 a_n1540_n1288# 0.159643f
C89 source.n6 a_n1540_n1288# 0.035883f
C90 source.n7 a_n1540_n1288# 0.382753f
C91 source.t8 a_n1540_n1288# 0.035444f
C92 source.t7 a_n1540_n1288# 0.035444f
C93 source.n8 a_n1540_n1288# 0.189484f
C94 source.n9 a_n1540_n1288# 0.304554f
C95 source.n10 a_n1540_n1288# 0.032733f
C96 source.n11 a_n1540_n1288# 0.072425f
C97 source.t0 a_n1540_n1288# 0.054352f
C98 source.n12 a_n1540_n1288# 0.056683f
C99 source.n13 a_n1540_n1288# 0.018272f
C100 source.n14 a_n1540_n1288# 0.012051f
C101 source.n15 a_n1540_n1288# 0.159643f
C102 source.n16 a_n1540_n1288# 0.035883f
C103 source.n17 a_n1540_n1288# 0.148661f
C104 source.t2 a_n1540_n1288# 0.035444f
C105 source.t1 a_n1540_n1288# 0.035444f
C106 source.n18 a_n1540_n1288# 0.189484f
C107 source.n19 a_n1540_n1288# 0.817581f
C108 source.t9 a_n1540_n1288# 0.035444f
C109 source.t6 a_n1540_n1288# 0.035444f
C110 source.n20 a_n1540_n1288# 0.189482f
C111 source.n21 a_n1540_n1288# 0.817582f
C112 source.n22 a_n1540_n1288# 0.032733f
C113 source.n23 a_n1540_n1288# 0.072425f
C114 source.t5 a_n1540_n1288# 0.054352f
C115 source.n24 a_n1540_n1288# 0.056683f
C116 source.n25 a_n1540_n1288# 0.018272f
C117 source.n26 a_n1540_n1288# 0.012051f
C118 source.n27 a_n1540_n1288# 0.159643f
C119 source.n28 a_n1540_n1288# 0.035883f
C120 source.n29 a_n1540_n1288# 0.148661f
C121 source.t10 a_n1540_n1288# 0.035444f
C122 source.t3 a_n1540_n1288# 0.035444f
C123 source.n30 a_n1540_n1288# 0.189482f
C124 source.n31 a_n1540_n1288# 0.304555f
C125 source.n32 a_n1540_n1288# 0.032733f
C126 source.n33 a_n1540_n1288# 0.072425f
C127 source.t11 a_n1540_n1288# 0.054352f
C128 source.n34 a_n1540_n1288# 0.056683f
C129 source.n35 a_n1540_n1288# 0.018272f
C130 source.n36 a_n1540_n1288# 0.012051f
C131 source.n37 a_n1540_n1288# 0.159643f
C132 source.n38 a_n1540_n1288# 0.035883f
C133 source.n39 a_n1540_n1288# 0.262867f
C134 source.n40 a_n1540_n1288# 0.565378f
C135 plus.n0 a_n1540_n1288# 0.12199f
C136 plus.t0 a_n1540_n1288# 0.127743f
C137 plus.t3 a_n1540_n1288# 0.127743f
C138 plus.t2 a_n1540_n1288# 0.140798f
C139 plus.n1 a_n1540_n1288# 0.078459f
C140 plus.n2 a_n1540_n1288# 0.091184f
C141 plus.n3 a_n1540_n1288# 0.006686f
C142 plus.n4 a_n1540_n1288# 0.086619f
C143 plus.n5 a_n1540_n1288# 0.219914f
C144 plus.n6 a_n1540_n1288# 0.12199f
C145 plus.t1 a_n1540_n1288# 0.127743f
C146 plus.t5 a_n1540_n1288# 0.140798f
C147 plus.n7 a_n1540_n1288# 0.078459f
C148 plus.t4 a_n1540_n1288# 0.127743f
C149 plus.n8 a_n1540_n1288# 0.091184f
C150 plus.n9 a_n1540_n1288# 0.006686f
C151 plus.n10 a_n1540_n1288# 0.086619f
C152 plus.n11 a_n1540_n1288# 0.634775f
.ends

