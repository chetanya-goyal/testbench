* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t11 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X1 a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X2 a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X3 drain_right.t9 minus.t0 source.t1 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X4 source.t0 minus.t1 drain_right.t8 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X5 source.t16 plus.t1 drain_left.t8 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X6 drain_right.t7 minus.t2 source.t3 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X7 drain_left.t7 plus.t2 source.t17 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X8 source.t6 minus.t3 drain_right.t6 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X9 drain_right.t5 minus.t4 source.t8 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X10 drain_left.t6 plus.t3 source.t13 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X11 source.t7 minus.t5 drain_right.t4 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X12 source.t12 plus.t4 drain_left.t5 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X13 source.t14 plus.t5 drain_left.t4 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X14 a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X15 drain_right.t3 minus.t6 source.t2 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X16 drain_right.t2 minus.t7 source.t4 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X17 drain_left.t3 plus.t6 source.t10 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X18 drain_left.t2 plus.t7 source.t18 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X19 source.t19 plus.t8 drain_left.t1 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X20 source.t5 minus.t8 drain_right.t1 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X21 a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X22 drain_left.t0 plus.t9 source.t15 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X23 drain_right.t0 minus.t9 source.t9 a_n1352_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n2 plus.t3 563.429
R1 plus.n8 plus.t7 563.429
R2 plus.n12 plus.t2 563.429
R3 plus.n18 plus.t6 563.429
R4 plus.n1 plus.t1 518.15
R5 plus.n5 plus.t9 518.15
R6 plus.n7 plus.t8 518.15
R7 plus.n11 plus.t5 518.15
R8 plus.n15 plus.t0 518.15
R9 plus.n17 plus.t4 518.15
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 40.8975
R19 plus.n7 plus.n6 40.8975
R20 plus.n17 plus.n16 40.8975
R21 plus.n14 plus.n11 40.8975
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus.n2 plus.n1 32.1338
R27 plus.n8 plus.n7 32.1338
R28 plus.n18 plus.n17 32.1338
R29 plus.n12 plus.n11 32.1338
R30 plus plus.n19 24.6638
R31 plus plus.n9 8.68421
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 source.n0 source.t18 69.6943
R37 source.n5 source.t2 69.6943
R38 source.n19 source.t8 69.6942
R39 source.n14 source.t17 69.6942
R40 source.n2 source.n1 63.0943
R41 source.n4 source.n3 63.0943
R42 source.n7 source.n6 63.0943
R43 source.n9 source.n8 63.0943
R44 source.n18 source.n17 63.0942
R45 source.n16 source.n15 63.0942
R46 source.n13 source.n12 63.0942
R47 source.n11 source.n10 63.0942
R48 source.n11 source.n9 15.3833
R49 source.n20 source.n0 9.43506
R50 source.n17 source.t9 6.6005
R51 source.n17 source.t0 6.6005
R52 source.n15 source.t3 6.6005
R53 source.n15 source.t7 6.6005
R54 source.n12 source.t11 6.6005
R55 source.n12 source.t14 6.6005
R56 source.n10 source.t10 6.6005
R57 source.n10 source.t12 6.6005
R58 source.n1 source.t15 6.6005
R59 source.n1 source.t19 6.6005
R60 source.n3 source.t13 6.6005
R61 source.n3 source.t16 6.6005
R62 source.n6 source.t1 6.6005
R63 source.n6 source.t6 6.6005
R64 source.n8 source.t4 6.6005
R65 source.n8 source.t5 6.6005
R66 source.n20 source.n19 5.49188
R67 source.n5 source.n4 0.698776
R68 source.n16 source.n14 0.698776
R69 source.n9 source.n7 0.457397
R70 source.n7 source.n5 0.457397
R71 source.n4 source.n2 0.457397
R72 source.n2 source.n0 0.457397
R73 source.n13 source.n11 0.457397
R74 source.n14 source.n13 0.457397
R75 source.n18 source.n16 0.457397
R76 source.n19 source.n18 0.457397
R77 source source.n20 0.188
R78 drain_left.n5 drain_left.t6 86.83
R79 drain_left.n1 drain_left.t3 86.8299
R80 drain_left.n3 drain_left.n2 80.0603
R81 drain_left.n7 drain_left.n6 79.7731
R82 drain_left.n5 drain_left.n4 79.7731
R83 drain_left.n1 drain_left.n0 79.773
R84 drain_left drain_left.n3 22.4907
R85 drain_left.n2 drain_left.t4 6.6005
R86 drain_left.n2 drain_left.t7 6.6005
R87 drain_left.n0 drain_left.t5 6.6005
R88 drain_left.n0 drain_left.t9 6.6005
R89 drain_left.n6 drain_left.t1 6.6005
R90 drain_left.n6 drain_left.t2 6.6005
R91 drain_left.n4 drain_left.t8 6.6005
R92 drain_left.n4 drain_left.t0 6.6005
R93 drain_left drain_left.n7 6.11011
R94 drain_left.n7 drain_left.n5 0.457397
R95 drain_left.n3 drain_left.n1 0.0593781
R96 minus.n8 minus.t7 563.429
R97 minus.n2 minus.t6 563.429
R98 minus.n18 minus.t4 563.429
R99 minus.n12 minus.t2 563.429
R100 minus.n7 minus.t8 518.15
R101 minus.n5 minus.t0 518.15
R102 minus.n1 minus.t3 518.15
R103 minus.n17 minus.t1 518.15
R104 minus.n15 minus.t9 518.15
R105 minus.n11 minus.t5 518.15
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 40.8975
R115 minus.n4 minus.n1 40.8975
R116 minus.n14 minus.n11 40.8975
R117 minus.n17 minus.n16 40.8975
R118 minus.n6 minus.n5 36.5157
R119 minus.n5 minus.n4 36.5157
R120 minus.n15 minus.n14 36.5157
R121 minus.n16 minus.n15 36.5157
R122 minus.n8 minus.n7 32.1338
R123 minus.n2 minus.n1 32.1338
R124 minus.n12 minus.n11 32.1338
R125 minus.n18 minus.n17 32.1338
R126 minus.n20 minus.n9 27.3736
R127 minus.n20 minus.n19 6.44936
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t7 86.8299
R134 drain_right.n7 drain_right.t2 86.3731
R135 drain_right.n6 drain_right.n4 80.23
R136 drain_right.n3 drain_right.n2 80.0603
R137 drain_right.n6 drain_right.n5 79.7731
R138 drain_right.n1 drain_right.n0 79.773
R139 drain_right drain_right.n3 21.9375
R140 drain_right.n2 drain_right.t8 6.6005
R141 drain_right.n2 drain_right.t5 6.6005
R142 drain_right.n0 drain_right.t4 6.6005
R143 drain_right.n0 drain_right.t0 6.6005
R144 drain_right.n4 drain_right.t6 6.6005
R145 drain_right.n4 drain_right.t3 6.6005
R146 drain_right.n5 drain_right.t1 6.6005
R147 drain_right.n5 drain_right.t9 6.6005
R148 drain_right drain_right.n7 5.88166
R149 drain_right.n7 drain_right.n6 0.457397
R150 drain_right.n3 drain_right.n1 0.0593781
C0 plus minus 3.18042f
C1 plus source 1.06826f
C2 drain_left minus 0.175826f
C3 drain_right minus 1.05528f
C4 drain_left source 7.78861f
C5 drain_right source 7.78401f
C6 drain_left plus 1.18246f
C7 drain_right plus 0.287486f
C8 drain_left drain_right 0.659063f
C9 minus source 1.05409f
C10 drain_right a_n1352_n1488# 3.87348f
C11 drain_left a_n1352_n1488# 4.061181f
C12 source a_n1352_n1488# 2.741466f
C13 minus a_n1352_n1488# 4.503664f
C14 plus a_n1352_n1488# 5.2451f
C15 drain_right.t7 a_n1352_n1488# 0.610374f
C16 drain_right.t4 a_n1352_n1488# 0.065762f
C17 drain_right.t0 a_n1352_n1488# 0.065762f
C18 drain_right.n0 a_n1352_n1488# 0.474266f
C19 drain_right.n1 a_n1352_n1488# 0.596376f
C20 drain_right.t8 a_n1352_n1488# 0.065762f
C21 drain_right.t5 a_n1352_n1488# 0.065762f
C22 drain_right.n2 a_n1352_n1488# 0.475349f
C23 drain_right.n3 a_n1352_n1488# 0.936072f
C24 drain_right.t6 a_n1352_n1488# 0.065762f
C25 drain_right.t3 a_n1352_n1488# 0.065762f
C26 drain_right.n4 a_n1352_n1488# 0.476061f
C27 drain_right.t1 a_n1352_n1488# 0.065762f
C28 drain_right.t9 a_n1352_n1488# 0.065762f
C29 drain_right.n5 a_n1352_n1488# 0.474268f
C30 drain_right.n6 a_n1352_n1488# 0.616829f
C31 drain_right.t2 a_n1352_n1488# 0.608698f
C32 drain_right.n7 a_n1352_n1488# 0.544438f
C33 minus.n0 a_n1352_n1488# 0.033934f
C34 minus.t7 a_n1352_n1488# 0.06201f
C35 minus.t8 a_n1352_n1488# 0.058962f
C36 minus.t0 a_n1352_n1488# 0.058962f
C37 minus.t3 a_n1352_n1488# 0.058962f
C38 minus.n1 a_n1352_n1488# 0.037723f
C39 minus.t6 a_n1352_n1488# 0.06201f
C40 minus.n2 a_n1352_n1488# 0.046816f
C41 minus.n3 a_n1352_n1488# 0.074516f
C42 minus.n4 a_n1352_n1488# 0.011885f
C43 minus.n5 a_n1352_n1488# 0.037723f
C44 minus.n6 a_n1352_n1488# 0.011885f
C45 minus.n7 a_n1352_n1488# 0.037723f
C46 minus.n8 a_n1352_n1488# 0.046769f
C47 minus.n9 a_n1352_n1488# 0.750311f
C48 minus.n10 a_n1352_n1488# 0.033934f
C49 minus.t1 a_n1352_n1488# 0.058962f
C50 minus.t9 a_n1352_n1488# 0.058962f
C51 minus.t5 a_n1352_n1488# 0.058962f
C52 minus.n11 a_n1352_n1488# 0.037723f
C53 minus.t2 a_n1352_n1488# 0.06201f
C54 minus.n12 a_n1352_n1488# 0.046816f
C55 minus.n13 a_n1352_n1488# 0.074516f
C56 minus.n14 a_n1352_n1488# 0.011885f
C57 minus.n15 a_n1352_n1488# 0.037723f
C58 minus.n16 a_n1352_n1488# 0.011885f
C59 minus.n17 a_n1352_n1488# 0.037723f
C60 minus.t4 a_n1352_n1488# 0.06201f
C61 minus.n18 a_n1352_n1488# 0.046769f
C62 minus.n19 a_n1352_n1488# 0.217795f
C63 minus.n20 a_n1352_n1488# 0.929854f
C64 drain_left.t3 a_n1352_n1488# 0.601999f
C65 drain_left.t5 a_n1352_n1488# 0.064859f
C66 drain_left.t9 a_n1352_n1488# 0.064859f
C67 drain_left.n0 a_n1352_n1488# 0.467758f
C68 drain_left.n1 a_n1352_n1488# 0.588193f
C69 drain_left.t4 a_n1352_n1488# 0.064859f
C70 drain_left.t7 a_n1352_n1488# 0.064859f
C71 drain_left.n2 a_n1352_n1488# 0.468827f
C72 drain_left.n3 a_n1352_n1488# 0.977777f
C73 drain_left.t6 a_n1352_n1488# 0.602001f
C74 drain_left.t8 a_n1352_n1488# 0.064859f
C75 drain_left.t0 a_n1352_n1488# 0.064859f
C76 drain_left.n4 a_n1352_n1488# 0.467761f
C77 drain_left.n5 a_n1352_n1488# 0.612504f
C78 drain_left.t1 a_n1352_n1488# 0.064859f
C79 drain_left.t2 a_n1352_n1488# 0.064859f
C80 drain_left.n6 a_n1352_n1488# 0.467761f
C81 drain_left.n7 a_n1352_n1488# 0.523463f
C82 source.t18 a_n1352_n1488# 0.632505f
C83 source.n0 a_n1352_n1488# 0.84722f
C84 source.t15 a_n1352_n1488# 0.07617f
C85 source.t19 a_n1352_n1488# 0.07617f
C86 source.n1 a_n1352_n1488# 0.482964f
C87 source.n2 a_n1352_n1488# 0.374499f
C88 source.t13 a_n1352_n1488# 0.07617f
C89 source.t16 a_n1352_n1488# 0.07617f
C90 source.n3 a_n1352_n1488# 0.482964f
C91 source.n4 a_n1352_n1488# 0.399489f
C92 source.t2 a_n1352_n1488# 0.632505f
C93 source.n5 a_n1352_n1488# 0.457685f
C94 source.t1 a_n1352_n1488# 0.07617f
C95 source.t6 a_n1352_n1488# 0.07617f
C96 source.n6 a_n1352_n1488# 0.482964f
C97 source.n7 a_n1352_n1488# 0.374499f
C98 source.t4 a_n1352_n1488# 0.07617f
C99 source.t5 a_n1352_n1488# 0.07617f
C100 source.n8 a_n1352_n1488# 0.482964f
C101 source.n9 a_n1352_n1488# 1.16912f
C102 source.t10 a_n1352_n1488# 0.07617f
C103 source.t12 a_n1352_n1488# 0.07617f
C104 source.n10 a_n1352_n1488# 0.48296f
C105 source.n11 a_n1352_n1488# 1.16912f
C106 source.t11 a_n1352_n1488# 0.07617f
C107 source.t14 a_n1352_n1488# 0.07617f
C108 source.n12 a_n1352_n1488# 0.48296f
C109 source.n13 a_n1352_n1488# 0.374503f
C110 source.t17 a_n1352_n1488# 0.632502f
C111 source.n14 a_n1352_n1488# 0.457688f
C112 source.t3 a_n1352_n1488# 0.07617f
C113 source.t7 a_n1352_n1488# 0.07617f
C114 source.n15 a_n1352_n1488# 0.48296f
C115 source.n16 a_n1352_n1488# 0.399493f
C116 source.t9 a_n1352_n1488# 0.07617f
C117 source.t0 a_n1352_n1488# 0.07617f
C118 source.n17 a_n1352_n1488# 0.48296f
C119 source.n18 a_n1352_n1488# 0.374503f
C120 source.t8 a_n1352_n1488# 0.632502f
C121 source.n19 a_n1352_n1488# 0.608256f
C122 source.n20 a_n1352_n1488# 0.927403f
C123 plus.n0 a_n1352_n1488# 0.034678f
C124 plus.t8 a_n1352_n1488# 0.060254f
C125 plus.t9 a_n1352_n1488# 0.060254f
C126 plus.t1 a_n1352_n1488# 0.060254f
C127 plus.n1 a_n1352_n1488# 0.038549f
C128 plus.t3 a_n1352_n1488# 0.063369f
C129 plus.n2 a_n1352_n1488# 0.047842f
C130 plus.n3 a_n1352_n1488# 0.076149f
C131 plus.n4 a_n1352_n1488# 0.012145f
C132 plus.n5 a_n1352_n1488# 0.038549f
C133 plus.n6 a_n1352_n1488# 0.012145f
C134 plus.n7 a_n1352_n1488# 0.038549f
C135 plus.t7 a_n1352_n1488# 0.063369f
C136 plus.n8 a_n1352_n1488# 0.047793f
C137 plus.n9 a_n1352_n1488# 0.254678f
C138 plus.n10 a_n1352_n1488# 0.034678f
C139 plus.t6 a_n1352_n1488# 0.063369f
C140 plus.t4 a_n1352_n1488# 0.060254f
C141 plus.t0 a_n1352_n1488# 0.060254f
C142 plus.t5 a_n1352_n1488# 0.060254f
C143 plus.n11 a_n1352_n1488# 0.038549f
C144 plus.t2 a_n1352_n1488# 0.063369f
C145 plus.n12 a_n1352_n1488# 0.047842f
C146 plus.n13 a_n1352_n1488# 0.076149f
C147 plus.n14 a_n1352_n1488# 0.012145f
C148 plus.n15 a_n1352_n1488# 0.038549f
C149 plus.n16 a_n1352_n1488# 0.012145f
C150 plus.n17 a_n1352_n1488# 0.038549f
C151 plus.n18 a_n1352_n1488# 0.047793f
C152 plus.n19 a_n1352_n1488# 0.724261f
.ends

