* NGSPICE file created from diffpair151.ext - technology: sky130A

.subckt diffpair151 minus drain_right drain_left source plus
X0 a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X1 drain_right minus source a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X2 a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X3 a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X4 source plus drain_left a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X5 a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X6 source minus drain_right a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X7 drain_right minus source a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X8 source minus drain_right a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X9 drain_left plus source a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X10 drain_left plus source a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X11 source plus drain_left a_n1394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
.ends

