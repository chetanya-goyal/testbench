* NGSPICE file created from diffpair678.ext - technology: sky130A

.subckt diffpair678 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t31 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X1 source.t8 minus.t0 drain_right.t19 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X2 drain_right.t18 minus.t1 source.t1 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X3 drain_right.t17 minus.t2 source.t4 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X4 source.t11 minus.t3 drain_right.t16 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X5 source.t13 minus.t4 drain_right.t15 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X6 drain_right.t14 minus.t5 source.t14 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X7 source.t23 plus.t1 drain_left.t18 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X8 drain_left.t17 plus.t2 source.t30 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X9 drain_right.t13 minus.t6 source.t9 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X10 drain_left.t16 plus.t3 source.t22 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X11 source.t38 minus.t7 drain_right.t12 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X12 drain_left.t15 plus.t4 source.t21 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X13 a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X14 source.t20 plus.t5 drain_left.t14 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X15 drain_left.t13 plus.t6 source.t28 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X16 source.t39 minus.t8 drain_right.t11 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X17 source.t3 minus.t9 drain_right.t10 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X18 a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X19 source.t0 minus.t10 drain_right.t9 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X20 a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X21 source.t19 plus.t7 drain_left.t12 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X22 source.t24 plus.t8 drain_left.t11 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X23 drain_right.t8 minus.t11 source.t2 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X24 drain_left.t10 plus.t9 source.t18 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X25 source.t27 plus.t10 drain_left.t9 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X26 source.t32 plus.t11 drain_left.t8 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X27 source.t25 plus.t12 drain_left.t7 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X28 a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X29 drain_right.t7 minus.t12 source.t16 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X30 drain_right.t6 minus.t13 source.t10 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X31 drain_left.t6 plus.t13 source.t37 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X32 source.t6 minus.t14 drain_right.t5 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X33 drain_right.t4 minus.t15 source.t12 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X34 drain_right.t3 minus.t16 source.t15 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X35 source.t29 plus.t14 drain_left.t5 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X36 source.t5 minus.t17 drain_right.t2 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X37 source.t7 minus.t18 drain_right.t1 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X38 drain_right.t0 minus.t19 source.t17 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X39 source.t26 plus.t15 drain_left.t4 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X40 source.t33 plus.t16 drain_left.t3 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X41 drain_left.t2 plus.t17 source.t34 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X42 drain_left.t1 plus.t18 source.t35 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X43 drain_left.t0 plus.t19 source.t36 a_n2102_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
R0 plus.n6 plus.t1 2161.7
R1 plus.n27 plus.t13 2161.7
R2 plus.n36 plus.t18 2161.7
R3 plus.n56 plus.t15 2161.7
R4 plus.n5 plus.t6 2112.77
R5 plus.n9 plus.t11 2112.77
R6 plus.n3 plus.t17 2112.77
R7 plus.n15 plus.t5 2112.77
R8 plus.n17 plus.t9 2112.77
R9 plus.n18 plus.t16 2112.77
R10 plus.n24 plus.t0 2112.77
R11 plus.n26 plus.t7 2112.77
R12 plus.n35 plus.t8 2112.77
R13 plus.n39 plus.t19 2112.77
R14 plus.n33 plus.t10 2112.77
R15 plus.n45 plus.t3 2112.77
R16 plus.n47 plus.t12 2112.77
R17 plus.n32 plus.t4 2112.77
R18 plus.n53 plus.t14 2112.77
R19 plus.n55 plus.t2 2112.77
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 64.9975
R47 plus.n19 plus.n18 64.9975
R48 plus.n48 plus.n32 64.9975
R49 plus.n44 plus.n33 64.9975
R50 plus.n9 plus.n8 62.0763
R51 plus.n25 plus.n24 62.0763
R52 plus.n54 plus.n53 62.0763
R53 plus.n39 plus.n38 62.0763
R54 plus.n16 plus.n15 46.0096
R55 plus.n17 plus.n16 46.0096
R56 plus.n47 plus.n46 46.0096
R57 plus.n46 plus.n45 46.0096
R58 plus.n6 plus.n5 43.0884
R59 plus.n27 plus.n26 43.0884
R60 plus.n56 plus.n55 43.0884
R61 plus.n36 plus.n35 43.0884
R62 plus plus.n57 35.9043
R63 plus.n8 plus.n5 29.9429
R64 plus.n26 plus.n25 29.9429
R65 plus.n55 plus.n54 29.9429
R66 plus.n38 plus.n35 29.9429
R67 plus.n15 plus.n14 27.0217
R68 plus.n19 plus.n17 27.0217
R69 plus.n48 plus.n47 27.0217
R70 plus.n45 plus.n44 27.0217
R71 plus plus.n28 17.0838
R72 plus.n10 plus.n9 10.955
R73 plus.n24 plus.n23 10.955
R74 plus.n53 plus.n52 10.955
R75 plus.n40 plus.n39 10.955
R76 plus.n11 plus.n3 8.03383
R77 plus.n18 plus.n1 8.03383
R78 plus.n32 plus.n30 8.03383
R79 plus.n41 plus.n33 8.03383
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n1146 source.n1012 289.615
R99 source.n998 source.n864 289.615
R100 source.n858 source.n724 289.615
R101 source.n710 source.n576 289.615
R102 source.n134 source.n0 289.615
R103 source.n282 source.n148 289.615
R104 source.n422 source.n288 289.615
R105 source.n570 source.n436 289.615
R106 source.n1056 source.n1055 185
R107 source.n1061 source.n1060 185
R108 source.n1063 source.n1062 185
R109 source.n1052 source.n1051 185
R110 source.n1069 source.n1068 185
R111 source.n1071 source.n1070 185
R112 source.n1048 source.n1047 185
R113 source.n1078 source.n1077 185
R114 source.n1079 source.n1046 185
R115 source.n1081 source.n1080 185
R116 source.n1044 source.n1043 185
R117 source.n1087 source.n1086 185
R118 source.n1089 source.n1088 185
R119 source.n1040 source.n1039 185
R120 source.n1095 source.n1094 185
R121 source.n1097 source.n1096 185
R122 source.n1036 source.n1035 185
R123 source.n1103 source.n1102 185
R124 source.n1105 source.n1104 185
R125 source.n1032 source.n1031 185
R126 source.n1111 source.n1110 185
R127 source.n1113 source.n1112 185
R128 source.n1028 source.n1027 185
R129 source.n1119 source.n1118 185
R130 source.n1122 source.n1121 185
R131 source.n1120 source.n1024 185
R132 source.n1127 source.n1023 185
R133 source.n1129 source.n1128 185
R134 source.n1131 source.n1130 185
R135 source.n1020 source.n1019 185
R136 source.n1137 source.n1136 185
R137 source.n1139 source.n1138 185
R138 source.n1016 source.n1015 185
R139 source.n1145 source.n1144 185
R140 source.n1147 source.n1146 185
R141 source.n908 source.n907 185
R142 source.n913 source.n912 185
R143 source.n915 source.n914 185
R144 source.n904 source.n903 185
R145 source.n921 source.n920 185
R146 source.n923 source.n922 185
R147 source.n900 source.n899 185
R148 source.n930 source.n929 185
R149 source.n931 source.n898 185
R150 source.n933 source.n932 185
R151 source.n896 source.n895 185
R152 source.n939 source.n938 185
R153 source.n941 source.n940 185
R154 source.n892 source.n891 185
R155 source.n947 source.n946 185
R156 source.n949 source.n948 185
R157 source.n888 source.n887 185
R158 source.n955 source.n954 185
R159 source.n957 source.n956 185
R160 source.n884 source.n883 185
R161 source.n963 source.n962 185
R162 source.n965 source.n964 185
R163 source.n880 source.n879 185
R164 source.n971 source.n970 185
R165 source.n974 source.n973 185
R166 source.n972 source.n876 185
R167 source.n979 source.n875 185
R168 source.n981 source.n980 185
R169 source.n983 source.n982 185
R170 source.n872 source.n871 185
R171 source.n989 source.n988 185
R172 source.n991 source.n990 185
R173 source.n868 source.n867 185
R174 source.n997 source.n996 185
R175 source.n999 source.n998 185
R176 source.n768 source.n767 185
R177 source.n773 source.n772 185
R178 source.n775 source.n774 185
R179 source.n764 source.n763 185
R180 source.n781 source.n780 185
R181 source.n783 source.n782 185
R182 source.n760 source.n759 185
R183 source.n790 source.n789 185
R184 source.n791 source.n758 185
R185 source.n793 source.n792 185
R186 source.n756 source.n755 185
R187 source.n799 source.n798 185
R188 source.n801 source.n800 185
R189 source.n752 source.n751 185
R190 source.n807 source.n806 185
R191 source.n809 source.n808 185
R192 source.n748 source.n747 185
R193 source.n815 source.n814 185
R194 source.n817 source.n816 185
R195 source.n744 source.n743 185
R196 source.n823 source.n822 185
R197 source.n825 source.n824 185
R198 source.n740 source.n739 185
R199 source.n831 source.n830 185
R200 source.n834 source.n833 185
R201 source.n832 source.n736 185
R202 source.n839 source.n735 185
R203 source.n841 source.n840 185
R204 source.n843 source.n842 185
R205 source.n732 source.n731 185
R206 source.n849 source.n848 185
R207 source.n851 source.n850 185
R208 source.n728 source.n727 185
R209 source.n857 source.n856 185
R210 source.n859 source.n858 185
R211 source.n620 source.n619 185
R212 source.n625 source.n624 185
R213 source.n627 source.n626 185
R214 source.n616 source.n615 185
R215 source.n633 source.n632 185
R216 source.n635 source.n634 185
R217 source.n612 source.n611 185
R218 source.n642 source.n641 185
R219 source.n643 source.n610 185
R220 source.n645 source.n644 185
R221 source.n608 source.n607 185
R222 source.n651 source.n650 185
R223 source.n653 source.n652 185
R224 source.n604 source.n603 185
R225 source.n659 source.n658 185
R226 source.n661 source.n660 185
R227 source.n600 source.n599 185
R228 source.n667 source.n666 185
R229 source.n669 source.n668 185
R230 source.n596 source.n595 185
R231 source.n675 source.n674 185
R232 source.n677 source.n676 185
R233 source.n592 source.n591 185
R234 source.n683 source.n682 185
R235 source.n686 source.n685 185
R236 source.n684 source.n588 185
R237 source.n691 source.n587 185
R238 source.n693 source.n692 185
R239 source.n695 source.n694 185
R240 source.n584 source.n583 185
R241 source.n701 source.n700 185
R242 source.n703 source.n702 185
R243 source.n580 source.n579 185
R244 source.n709 source.n708 185
R245 source.n711 source.n710 185
R246 source.n135 source.n134 185
R247 source.n133 source.n132 185
R248 source.n4 source.n3 185
R249 source.n127 source.n126 185
R250 source.n125 source.n124 185
R251 source.n8 source.n7 185
R252 source.n119 source.n118 185
R253 source.n117 source.n116 185
R254 source.n115 source.n11 185
R255 source.n15 source.n12 185
R256 source.n110 source.n109 185
R257 source.n108 source.n107 185
R258 source.n17 source.n16 185
R259 source.n102 source.n101 185
R260 source.n100 source.n99 185
R261 source.n21 source.n20 185
R262 source.n94 source.n93 185
R263 source.n92 source.n91 185
R264 source.n25 source.n24 185
R265 source.n86 source.n85 185
R266 source.n84 source.n83 185
R267 source.n29 source.n28 185
R268 source.n78 source.n77 185
R269 source.n76 source.n75 185
R270 source.n33 source.n32 185
R271 source.n70 source.n69 185
R272 source.n68 source.n35 185
R273 source.n67 source.n66 185
R274 source.n38 source.n36 185
R275 source.n61 source.n60 185
R276 source.n59 source.n58 185
R277 source.n42 source.n41 185
R278 source.n53 source.n52 185
R279 source.n51 source.n50 185
R280 source.n46 source.n45 185
R281 source.n283 source.n282 185
R282 source.n281 source.n280 185
R283 source.n152 source.n151 185
R284 source.n275 source.n274 185
R285 source.n273 source.n272 185
R286 source.n156 source.n155 185
R287 source.n267 source.n266 185
R288 source.n265 source.n264 185
R289 source.n263 source.n159 185
R290 source.n163 source.n160 185
R291 source.n258 source.n257 185
R292 source.n256 source.n255 185
R293 source.n165 source.n164 185
R294 source.n250 source.n249 185
R295 source.n248 source.n247 185
R296 source.n169 source.n168 185
R297 source.n242 source.n241 185
R298 source.n240 source.n239 185
R299 source.n173 source.n172 185
R300 source.n234 source.n233 185
R301 source.n232 source.n231 185
R302 source.n177 source.n176 185
R303 source.n226 source.n225 185
R304 source.n224 source.n223 185
R305 source.n181 source.n180 185
R306 source.n218 source.n217 185
R307 source.n216 source.n183 185
R308 source.n215 source.n214 185
R309 source.n186 source.n184 185
R310 source.n209 source.n208 185
R311 source.n207 source.n206 185
R312 source.n190 source.n189 185
R313 source.n201 source.n200 185
R314 source.n199 source.n198 185
R315 source.n194 source.n193 185
R316 source.n423 source.n422 185
R317 source.n421 source.n420 185
R318 source.n292 source.n291 185
R319 source.n415 source.n414 185
R320 source.n413 source.n412 185
R321 source.n296 source.n295 185
R322 source.n407 source.n406 185
R323 source.n405 source.n404 185
R324 source.n403 source.n299 185
R325 source.n303 source.n300 185
R326 source.n398 source.n397 185
R327 source.n396 source.n395 185
R328 source.n305 source.n304 185
R329 source.n390 source.n389 185
R330 source.n388 source.n387 185
R331 source.n309 source.n308 185
R332 source.n382 source.n381 185
R333 source.n380 source.n379 185
R334 source.n313 source.n312 185
R335 source.n374 source.n373 185
R336 source.n372 source.n371 185
R337 source.n317 source.n316 185
R338 source.n366 source.n365 185
R339 source.n364 source.n363 185
R340 source.n321 source.n320 185
R341 source.n358 source.n357 185
R342 source.n356 source.n323 185
R343 source.n355 source.n354 185
R344 source.n326 source.n324 185
R345 source.n349 source.n348 185
R346 source.n347 source.n346 185
R347 source.n330 source.n329 185
R348 source.n341 source.n340 185
R349 source.n339 source.n338 185
R350 source.n334 source.n333 185
R351 source.n571 source.n570 185
R352 source.n569 source.n568 185
R353 source.n440 source.n439 185
R354 source.n563 source.n562 185
R355 source.n561 source.n560 185
R356 source.n444 source.n443 185
R357 source.n555 source.n554 185
R358 source.n553 source.n552 185
R359 source.n551 source.n447 185
R360 source.n451 source.n448 185
R361 source.n546 source.n545 185
R362 source.n544 source.n543 185
R363 source.n453 source.n452 185
R364 source.n538 source.n537 185
R365 source.n536 source.n535 185
R366 source.n457 source.n456 185
R367 source.n530 source.n529 185
R368 source.n528 source.n527 185
R369 source.n461 source.n460 185
R370 source.n522 source.n521 185
R371 source.n520 source.n519 185
R372 source.n465 source.n464 185
R373 source.n514 source.n513 185
R374 source.n512 source.n511 185
R375 source.n469 source.n468 185
R376 source.n506 source.n505 185
R377 source.n504 source.n471 185
R378 source.n503 source.n502 185
R379 source.n474 source.n472 185
R380 source.n497 source.n496 185
R381 source.n495 source.n494 185
R382 source.n478 source.n477 185
R383 source.n489 source.n488 185
R384 source.n487 source.n486 185
R385 source.n482 source.n481 185
R386 source.n1057 source.t14 149.524
R387 source.n909 source.t13 149.524
R388 source.n769 source.t35 149.524
R389 source.n621 source.t26 149.524
R390 source.n47 source.t37 149.524
R391 source.n195 source.t23 149.524
R392 source.n335 source.t2 149.524
R393 source.n483 source.t38 149.524
R394 source.n1061 source.n1055 104.615
R395 source.n1062 source.n1061 104.615
R396 source.n1062 source.n1051 104.615
R397 source.n1069 source.n1051 104.615
R398 source.n1070 source.n1069 104.615
R399 source.n1070 source.n1047 104.615
R400 source.n1078 source.n1047 104.615
R401 source.n1079 source.n1078 104.615
R402 source.n1080 source.n1079 104.615
R403 source.n1080 source.n1043 104.615
R404 source.n1087 source.n1043 104.615
R405 source.n1088 source.n1087 104.615
R406 source.n1088 source.n1039 104.615
R407 source.n1095 source.n1039 104.615
R408 source.n1096 source.n1095 104.615
R409 source.n1096 source.n1035 104.615
R410 source.n1103 source.n1035 104.615
R411 source.n1104 source.n1103 104.615
R412 source.n1104 source.n1031 104.615
R413 source.n1111 source.n1031 104.615
R414 source.n1112 source.n1111 104.615
R415 source.n1112 source.n1027 104.615
R416 source.n1119 source.n1027 104.615
R417 source.n1121 source.n1119 104.615
R418 source.n1121 source.n1120 104.615
R419 source.n1120 source.n1023 104.615
R420 source.n1129 source.n1023 104.615
R421 source.n1130 source.n1129 104.615
R422 source.n1130 source.n1019 104.615
R423 source.n1137 source.n1019 104.615
R424 source.n1138 source.n1137 104.615
R425 source.n1138 source.n1015 104.615
R426 source.n1145 source.n1015 104.615
R427 source.n1146 source.n1145 104.615
R428 source.n913 source.n907 104.615
R429 source.n914 source.n913 104.615
R430 source.n914 source.n903 104.615
R431 source.n921 source.n903 104.615
R432 source.n922 source.n921 104.615
R433 source.n922 source.n899 104.615
R434 source.n930 source.n899 104.615
R435 source.n931 source.n930 104.615
R436 source.n932 source.n931 104.615
R437 source.n932 source.n895 104.615
R438 source.n939 source.n895 104.615
R439 source.n940 source.n939 104.615
R440 source.n940 source.n891 104.615
R441 source.n947 source.n891 104.615
R442 source.n948 source.n947 104.615
R443 source.n948 source.n887 104.615
R444 source.n955 source.n887 104.615
R445 source.n956 source.n955 104.615
R446 source.n956 source.n883 104.615
R447 source.n963 source.n883 104.615
R448 source.n964 source.n963 104.615
R449 source.n964 source.n879 104.615
R450 source.n971 source.n879 104.615
R451 source.n973 source.n971 104.615
R452 source.n973 source.n972 104.615
R453 source.n972 source.n875 104.615
R454 source.n981 source.n875 104.615
R455 source.n982 source.n981 104.615
R456 source.n982 source.n871 104.615
R457 source.n989 source.n871 104.615
R458 source.n990 source.n989 104.615
R459 source.n990 source.n867 104.615
R460 source.n997 source.n867 104.615
R461 source.n998 source.n997 104.615
R462 source.n773 source.n767 104.615
R463 source.n774 source.n773 104.615
R464 source.n774 source.n763 104.615
R465 source.n781 source.n763 104.615
R466 source.n782 source.n781 104.615
R467 source.n782 source.n759 104.615
R468 source.n790 source.n759 104.615
R469 source.n791 source.n790 104.615
R470 source.n792 source.n791 104.615
R471 source.n792 source.n755 104.615
R472 source.n799 source.n755 104.615
R473 source.n800 source.n799 104.615
R474 source.n800 source.n751 104.615
R475 source.n807 source.n751 104.615
R476 source.n808 source.n807 104.615
R477 source.n808 source.n747 104.615
R478 source.n815 source.n747 104.615
R479 source.n816 source.n815 104.615
R480 source.n816 source.n743 104.615
R481 source.n823 source.n743 104.615
R482 source.n824 source.n823 104.615
R483 source.n824 source.n739 104.615
R484 source.n831 source.n739 104.615
R485 source.n833 source.n831 104.615
R486 source.n833 source.n832 104.615
R487 source.n832 source.n735 104.615
R488 source.n841 source.n735 104.615
R489 source.n842 source.n841 104.615
R490 source.n842 source.n731 104.615
R491 source.n849 source.n731 104.615
R492 source.n850 source.n849 104.615
R493 source.n850 source.n727 104.615
R494 source.n857 source.n727 104.615
R495 source.n858 source.n857 104.615
R496 source.n625 source.n619 104.615
R497 source.n626 source.n625 104.615
R498 source.n626 source.n615 104.615
R499 source.n633 source.n615 104.615
R500 source.n634 source.n633 104.615
R501 source.n634 source.n611 104.615
R502 source.n642 source.n611 104.615
R503 source.n643 source.n642 104.615
R504 source.n644 source.n643 104.615
R505 source.n644 source.n607 104.615
R506 source.n651 source.n607 104.615
R507 source.n652 source.n651 104.615
R508 source.n652 source.n603 104.615
R509 source.n659 source.n603 104.615
R510 source.n660 source.n659 104.615
R511 source.n660 source.n599 104.615
R512 source.n667 source.n599 104.615
R513 source.n668 source.n667 104.615
R514 source.n668 source.n595 104.615
R515 source.n675 source.n595 104.615
R516 source.n676 source.n675 104.615
R517 source.n676 source.n591 104.615
R518 source.n683 source.n591 104.615
R519 source.n685 source.n683 104.615
R520 source.n685 source.n684 104.615
R521 source.n684 source.n587 104.615
R522 source.n693 source.n587 104.615
R523 source.n694 source.n693 104.615
R524 source.n694 source.n583 104.615
R525 source.n701 source.n583 104.615
R526 source.n702 source.n701 104.615
R527 source.n702 source.n579 104.615
R528 source.n709 source.n579 104.615
R529 source.n710 source.n709 104.615
R530 source.n134 source.n133 104.615
R531 source.n133 source.n3 104.615
R532 source.n126 source.n3 104.615
R533 source.n126 source.n125 104.615
R534 source.n125 source.n7 104.615
R535 source.n118 source.n7 104.615
R536 source.n118 source.n117 104.615
R537 source.n117 source.n11 104.615
R538 source.n15 source.n11 104.615
R539 source.n109 source.n15 104.615
R540 source.n109 source.n108 104.615
R541 source.n108 source.n16 104.615
R542 source.n101 source.n16 104.615
R543 source.n101 source.n100 104.615
R544 source.n100 source.n20 104.615
R545 source.n93 source.n20 104.615
R546 source.n93 source.n92 104.615
R547 source.n92 source.n24 104.615
R548 source.n85 source.n24 104.615
R549 source.n85 source.n84 104.615
R550 source.n84 source.n28 104.615
R551 source.n77 source.n28 104.615
R552 source.n77 source.n76 104.615
R553 source.n76 source.n32 104.615
R554 source.n69 source.n32 104.615
R555 source.n69 source.n68 104.615
R556 source.n68 source.n67 104.615
R557 source.n67 source.n36 104.615
R558 source.n60 source.n36 104.615
R559 source.n60 source.n59 104.615
R560 source.n59 source.n41 104.615
R561 source.n52 source.n41 104.615
R562 source.n52 source.n51 104.615
R563 source.n51 source.n45 104.615
R564 source.n282 source.n281 104.615
R565 source.n281 source.n151 104.615
R566 source.n274 source.n151 104.615
R567 source.n274 source.n273 104.615
R568 source.n273 source.n155 104.615
R569 source.n266 source.n155 104.615
R570 source.n266 source.n265 104.615
R571 source.n265 source.n159 104.615
R572 source.n163 source.n159 104.615
R573 source.n257 source.n163 104.615
R574 source.n257 source.n256 104.615
R575 source.n256 source.n164 104.615
R576 source.n249 source.n164 104.615
R577 source.n249 source.n248 104.615
R578 source.n248 source.n168 104.615
R579 source.n241 source.n168 104.615
R580 source.n241 source.n240 104.615
R581 source.n240 source.n172 104.615
R582 source.n233 source.n172 104.615
R583 source.n233 source.n232 104.615
R584 source.n232 source.n176 104.615
R585 source.n225 source.n176 104.615
R586 source.n225 source.n224 104.615
R587 source.n224 source.n180 104.615
R588 source.n217 source.n180 104.615
R589 source.n217 source.n216 104.615
R590 source.n216 source.n215 104.615
R591 source.n215 source.n184 104.615
R592 source.n208 source.n184 104.615
R593 source.n208 source.n207 104.615
R594 source.n207 source.n189 104.615
R595 source.n200 source.n189 104.615
R596 source.n200 source.n199 104.615
R597 source.n199 source.n193 104.615
R598 source.n422 source.n421 104.615
R599 source.n421 source.n291 104.615
R600 source.n414 source.n291 104.615
R601 source.n414 source.n413 104.615
R602 source.n413 source.n295 104.615
R603 source.n406 source.n295 104.615
R604 source.n406 source.n405 104.615
R605 source.n405 source.n299 104.615
R606 source.n303 source.n299 104.615
R607 source.n397 source.n303 104.615
R608 source.n397 source.n396 104.615
R609 source.n396 source.n304 104.615
R610 source.n389 source.n304 104.615
R611 source.n389 source.n388 104.615
R612 source.n388 source.n308 104.615
R613 source.n381 source.n308 104.615
R614 source.n381 source.n380 104.615
R615 source.n380 source.n312 104.615
R616 source.n373 source.n312 104.615
R617 source.n373 source.n372 104.615
R618 source.n372 source.n316 104.615
R619 source.n365 source.n316 104.615
R620 source.n365 source.n364 104.615
R621 source.n364 source.n320 104.615
R622 source.n357 source.n320 104.615
R623 source.n357 source.n356 104.615
R624 source.n356 source.n355 104.615
R625 source.n355 source.n324 104.615
R626 source.n348 source.n324 104.615
R627 source.n348 source.n347 104.615
R628 source.n347 source.n329 104.615
R629 source.n340 source.n329 104.615
R630 source.n340 source.n339 104.615
R631 source.n339 source.n333 104.615
R632 source.n570 source.n569 104.615
R633 source.n569 source.n439 104.615
R634 source.n562 source.n439 104.615
R635 source.n562 source.n561 104.615
R636 source.n561 source.n443 104.615
R637 source.n554 source.n443 104.615
R638 source.n554 source.n553 104.615
R639 source.n553 source.n447 104.615
R640 source.n451 source.n447 104.615
R641 source.n545 source.n451 104.615
R642 source.n545 source.n544 104.615
R643 source.n544 source.n452 104.615
R644 source.n537 source.n452 104.615
R645 source.n537 source.n536 104.615
R646 source.n536 source.n456 104.615
R647 source.n529 source.n456 104.615
R648 source.n529 source.n528 104.615
R649 source.n528 source.n460 104.615
R650 source.n521 source.n460 104.615
R651 source.n521 source.n520 104.615
R652 source.n520 source.n464 104.615
R653 source.n513 source.n464 104.615
R654 source.n513 source.n512 104.615
R655 source.n512 source.n468 104.615
R656 source.n505 source.n468 104.615
R657 source.n505 source.n504 104.615
R658 source.n504 source.n503 104.615
R659 source.n503 source.n472 104.615
R660 source.n496 source.n472 104.615
R661 source.n496 source.n495 104.615
R662 source.n495 source.n477 104.615
R663 source.n488 source.n477 104.615
R664 source.n488 source.n487 104.615
R665 source.n487 source.n481 104.615
R666 source.t14 source.n1055 52.3082
R667 source.t13 source.n907 52.3082
R668 source.t35 source.n767 52.3082
R669 source.t26 source.n619 52.3082
R670 source.t37 source.n45 52.3082
R671 source.t23 source.n193 52.3082
R672 source.t2 source.n333 52.3082
R673 source.t38 source.n481 52.3082
R674 source.n1011 source.n1010 42.0366
R675 source.n1009 source.n1008 42.0366
R676 source.n1007 source.n1006 42.0366
R677 source.n1005 source.n1004 42.0366
R678 source.n723 source.n722 42.0366
R679 source.n721 source.n720 42.0366
R680 source.n719 source.n718 42.0366
R681 source.n717 source.n716 42.0366
R682 source.n141 source.n140 42.0366
R683 source.n143 source.n142 42.0366
R684 source.n145 source.n144 42.0366
R685 source.n147 source.n146 42.0366
R686 source.n429 source.n428 42.0366
R687 source.n431 source.n430 42.0366
R688 source.n433 source.n432 42.0366
R689 source.n435 source.n434 42.0366
R690 source.n715 source.n575 31.6793
R691 source.n1151 source.n1150 30.6338
R692 source.n1003 source.n1002 30.6338
R693 source.n863 source.n862 30.6338
R694 source.n715 source.n714 30.6338
R695 source.n139 source.n138 30.6338
R696 source.n287 source.n286 30.6338
R697 source.n427 source.n426 30.6338
R698 source.n575 source.n574 30.6338
R699 source.n1152 source.n139 26.1448
R700 source.n1081 source.n1046 13.1884
R701 source.n1128 source.n1127 13.1884
R702 source.n933 source.n898 13.1884
R703 source.n980 source.n979 13.1884
R704 source.n793 source.n758 13.1884
R705 source.n840 source.n839 13.1884
R706 source.n645 source.n610 13.1884
R707 source.n692 source.n691 13.1884
R708 source.n116 source.n115 13.1884
R709 source.n70 source.n35 13.1884
R710 source.n264 source.n263 13.1884
R711 source.n218 source.n183 13.1884
R712 source.n404 source.n403 13.1884
R713 source.n358 source.n323 13.1884
R714 source.n552 source.n551 13.1884
R715 source.n506 source.n471 13.1884
R716 source.n1077 source.n1076 12.8005
R717 source.n1082 source.n1044 12.8005
R718 source.n1126 source.n1024 12.8005
R719 source.n1131 source.n1022 12.8005
R720 source.n929 source.n928 12.8005
R721 source.n934 source.n896 12.8005
R722 source.n978 source.n876 12.8005
R723 source.n983 source.n874 12.8005
R724 source.n789 source.n788 12.8005
R725 source.n794 source.n756 12.8005
R726 source.n838 source.n736 12.8005
R727 source.n843 source.n734 12.8005
R728 source.n641 source.n640 12.8005
R729 source.n646 source.n608 12.8005
R730 source.n690 source.n588 12.8005
R731 source.n695 source.n586 12.8005
R732 source.n119 source.n10 12.8005
R733 source.n114 source.n12 12.8005
R734 source.n71 source.n33 12.8005
R735 source.n66 source.n37 12.8005
R736 source.n267 source.n158 12.8005
R737 source.n262 source.n160 12.8005
R738 source.n219 source.n181 12.8005
R739 source.n214 source.n185 12.8005
R740 source.n407 source.n298 12.8005
R741 source.n402 source.n300 12.8005
R742 source.n359 source.n321 12.8005
R743 source.n354 source.n325 12.8005
R744 source.n555 source.n446 12.8005
R745 source.n550 source.n448 12.8005
R746 source.n507 source.n469 12.8005
R747 source.n502 source.n473 12.8005
R748 source.n1075 source.n1048 12.0247
R749 source.n1086 source.n1085 12.0247
R750 source.n1123 source.n1122 12.0247
R751 source.n1132 source.n1020 12.0247
R752 source.n927 source.n900 12.0247
R753 source.n938 source.n937 12.0247
R754 source.n975 source.n974 12.0247
R755 source.n984 source.n872 12.0247
R756 source.n787 source.n760 12.0247
R757 source.n798 source.n797 12.0247
R758 source.n835 source.n834 12.0247
R759 source.n844 source.n732 12.0247
R760 source.n639 source.n612 12.0247
R761 source.n650 source.n649 12.0247
R762 source.n687 source.n686 12.0247
R763 source.n696 source.n584 12.0247
R764 source.n120 source.n8 12.0247
R765 source.n111 source.n110 12.0247
R766 source.n75 source.n74 12.0247
R767 source.n65 source.n38 12.0247
R768 source.n268 source.n156 12.0247
R769 source.n259 source.n258 12.0247
R770 source.n223 source.n222 12.0247
R771 source.n213 source.n186 12.0247
R772 source.n408 source.n296 12.0247
R773 source.n399 source.n398 12.0247
R774 source.n363 source.n362 12.0247
R775 source.n353 source.n326 12.0247
R776 source.n556 source.n444 12.0247
R777 source.n547 source.n546 12.0247
R778 source.n511 source.n510 12.0247
R779 source.n501 source.n474 12.0247
R780 source.n1072 source.n1071 11.249
R781 source.n1089 source.n1042 11.249
R782 source.n1118 source.n1026 11.249
R783 source.n1136 source.n1135 11.249
R784 source.n924 source.n923 11.249
R785 source.n941 source.n894 11.249
R786 source.n970 source.n878 11.249
R787 source.n988 source.n987 11.249
R788 source.n784 source.n783 11.249
R789 source.n801 source.n754 11.249
R790 source.n830 source.n738 11.249
R791 source.n848 source.n847 11.249
R792 source.n636 source.n635 11.249
R793 source.n653 source.n606 11.249
R794 source.n682 source.n590 11.249
R795 source.n700 source.n699 11.249
R796 source.n124 source.n123 11.249
R797 source.n107 source.n14 11.249
R798 source.n78 source.n31 11.249
R799 source.n62 source.n61 11.249
R800 source.n272 source.n271 11.249
R801 source.n255 source.n162 11.249
R802 source.n226 source.n179 11.249
R803 source.n210 source.n209 11.249
R804 source.n412 source.n411 11.249
R805 source.n395 source.n302 11.249
R806 source.n366 source.n319 11.249
R807 source.n350 source.n349 11.249
R808 source.n560 source.n559 11.249
R809 source.n543 source.n450 11.249
R810 source.n514 source.n467 11.249
R811 source.n498 source.n497 11.249
R812 source.n1068 source.n1050 10.4732
R813 source.n1090 source.n1040 10.4732
R814 source.n1117 source.n1028 10.4732
R815 source.n1139 source.n1018 10.4732
R816 source.n920 source.n902 10.4732
R817 source.n942 source.n892 10.4732
R818 source.n969 source.n880 10.4732
R819 source.n991 source.n870 10.4732
R820 source.n780 source.n762 10.4732
R821 source.n802 source.n752 10.4732
R822 source.n829 source.n740 10.4732
R823 source.n851 source.n730 10.4732
R824 source.n632 source.n614 10.4732
R825 source.n654 source.n604 10.4732
R826 source.n681 source.n592 10.4732
R827 source.n703 source.n582 10.4732
R828 source.n127 source.n6 10.4732
R829 source.n106 source.n17 10.4732
R830 source.n79 source.n29 10.4732
R831 source.n58 source.n40 10.4732
R832 source.n275 source.n154 10.4732
R833 source.n254 source.n165 10.4732
R834 source.n227 source.n177 10.4732
R835 source.n206 source.n188 10.4732
R836 source.n415 source.n294 10.4732
R837 source.n394 source.n305 10.4732
R838 source.n367 source.n317 10.4732
R839 source.n346 source.n328 10.4732
R840 source.n563 source.n442 10.4732
R841 source.n542 source.n453 10.4732
R842 source.n515 source.n465 10.4732
R843 source.n494 source.n476 10.4732
R844 source.n1057 source.n1056 10.2747
R845 source.n909 source.n908 10.2747
R846 source.n769 source.n768 10.2747
R847 source.n621 source.n620 10.2747
R848 source.n47 source.n46 10.2747
R849 source.n195 source.n194 10.2747
R850 source.n335 source.n334 10.2747
R851 source.n483 source.n482 10.2747
R852 source.n1067 source.n1052 9.69747
R853 source.n1094 source.n1093 9.69747
R854 source.n1114 source.n1113 9.69747
R855 source.n1140 source.n1016 9.69747
R856 source.n919 source.n904 9.69747
R857 source.n946 source.n945 9.69747
R858 source.n966 source.n965 9.69747
R859 source.n992 source.n868 9.69747
R860 source.n779 source.n764 9.69747
R861 source.n806 source.n805 9.69747
R862 source.n826 source.n825 9.69747
R863 source.n852 source.n728 9.69747
R864 source.n631 source.n616 9.69747
R865 source.n658 source.n657 9.69747
R866 source.n678 source.n677 9.69747
R867 source.n704 source.n580 9.69747
R868 source.n128 source.n4 9.69747
R869 source.n103 source.n102 9.69747
R870 source.n83 source.n82 9.69747
R871 source.n57 source.n42 9.69747
R872 source.n276 source.n152 9.69747
R873 source.n251 source.n250 9.69747
R874 source.n231 source.n230 9.69747
R875 source.n205 source.n190 9.69747
R876 source.n416 source.n292 9.69747
R877 source.n391 source.n390 9.69747
R878 source.n371 source.n370 9.69747
R879 source.n345 source.n330 9.69747
R880 source.n564 source.n440 9.69747
R881 source.n539 source.n538 9.69747
R882 source.n519 source.n518 9.69747
R883 source.n493 source.n478 9.69747
R884 source.n1150 source.n1149 9.45567
R885 source.n1002 source.n1001 9.45567
R886 source.n862 source.n861 9.45567
R887 source.n714 source.n713 9.45567
R888 source.n138 source.n137 9.45567
R889 source.n286 source.n285 9.45567
R890 source.n426 source.n425 9.45567
R891 source.n574 source.n573 9.45567
R892 source.n1014 source.n1013 9.3005
R893 source.n1143 source.n1142 9.3005
R894 source.n1141 source.n1140 9.3005
R895 source.n1018 source.n1017 9.3005
R896 source.n1135 source.n1134 9.3005
R897 source.n1133 source.n1132 9.3005
R898 source.n1022 source.n1021 9.3005
R899 source.n1101 source.n1100 9.3005
R900 source.n1099 source.n1098 9.3005
R901 source.n1038 source.n1037 9.3005
R902 source.n1093 source.n1092 9.3005
R903 source.n1091 source.n1090 9.3005
R904 source.n1042 source.n1041 9.3005
R905 source.n1085 source.n1084 9.3005
R906 source.n1083 source.n1082 9.3005
R907 source.n1059 source.n1058 9.3005
R908 source.n1054 source.n1053 9.3005
R909 source.n1065 source.n1064 9.3005
R910 source.n1067 source.n1066 9.3005
R911 source.n1050 source.n1049 9.3005
R912 source.n1073 source.n1072 9.3005
R913 source.n1075 source.n1074 9.3005
R914 source.n1076 source.n1045 9.3005
R915 source.n1034 source.n1033 9.3005
R916 source.n1107 source.n1106 9.3005
R917 source.n1109 source.n1108 9.3005
R918 source.n1030 source.n1029 9.3005
R919 source.n1115 source.n1114 9.3005
R920 source.n1117 source.n1116 9.3005
R921 source.n1026 source.n1025 9.3005
R922 source.n1124 source.n1123 9.3005
R923 source.n1126 source.n1125 9.3005
R924 source.n1149 source.n1148 9.3005
R925 source.n866 source.n865 9.3005
R926 source.n995 source.n994 9.3005
R927 source.n993 source.n992 9.3005
R928 source.n870 source.n869 9.3005
R929 source.n987 source.n986 9.3005
R930 source.n985 source.n984 9.3005
R931 source.n874 source.n873 9.3005
R932 source.n953 source.n952 9.3005
R933 source.n951 source.n950 9.3005
R934 source.n890 source.n889 9.3005
R935 source.n945 source.n944 9.3005
R936 source.n943 source.n942 9.3005
R937 source.n894 source.n893 9.3005
R938 source.n937 source.n936 9.3005
R939 source.n935 source.n934 9.3005
R940 source.n911 source.n910 9.3005
R941 source.n906 source.n905 9.3005
R942 source.n917 source.n916 9.3005
R943 source.n919 source.n918 9.3005
R944 source.n902 source.n901 9.3005
R945 source.n925 source.n924 9.3005
R946 source.n927 source.n926 9.3005
R947 source.n928 source.n897 9.3005
R948 source.n886 source.n885 9.3005
R949 source.n959 source.n958 9.3005
R950 source.n961 source.n960 9.3005
R951 source.n882 source.n881 9.3005
R952 source.n967 source.n966 9.3005
R953 source.n969 source.n968 9.3005
R954 source.n878 source.n877 9.3005
R955 source.n976 source.n975 9.3005
R956 source.n978 source.n977 9.3005
R957 source.n1001 source.n1000 9.3005
R958 source.n726 source.n725 9.3005
R959 source.n855 source.n854 9.3005
R960 source.n853 source.n852 9.3005
R961 source.n730 source.n729 9.3005
R962 source.n847 source.n846 9.3005
R963 source.n845 source.n844 9.3005
R964 source.n734 source.n733 9.3005
R965 source.n813 source.n812 9.3005
R966 source.n811 source.n810 9.3005
R967 source.n750 source.n749 9.3005
R968 source.n805 source.n804 9.3005
R969 source.n803 source.n802 9.3005
R970 source.n754 source.n753 9.3005
R971 source.n797 source.n796 9.3005
R972 source.n795 source.n794 9.3005
R973 source.n771 source.n770 9.3005
R974 source.n766 source.n765 9.3005
R975 source.n777 source.n776 9.3005
R976 source.n779 source.n778 9.3005
R977 source.n762 source.n761 9.3005
R978 source.n785 source.n784 9.3005
R979 source.n787 source.n786 9.3005
R980 source.n788 source.n757 9.3005
R981 source.n746 source.n745 9.3005
R982 source.n819 source.n818 9.3005
R983 source.n821 source.n820 9.3005
R984 source.n742 source.n741 9.3005
R985 source.n827 source.n826 9.3005
R986 source.n829 source.n828 9.3005
R987 source.n738 source.n737 9.3005
R988 source.n836 source.n835 9.3005
R989 source.n838 source.n837 9.3005
R990 source.n861 source.n860 9.3005
R991 source.n578 source.n577 9.3005
R992 source.n707 source.n706 9.3005
R993 source.n705 source.n704 9.3005
R994 source.n582 source.n581 9.3005
R995 source.n699 source.n698 9.3005
R996 source.n697 source.n696 9.3005
R997 source.n586 source.n585 9.3005
R998 source.n665 source.n664 9.3005
R999 source.n663 source.n662 9.3005
R1000 source.n602 source.n601 9.3005
R1001 source.n657 source.n656 9.3005
R1002 source.n655 source.n654 9.3005
R1003 source.n606 source.n605 9.3005
R1004 source.n649 source.n648 9.3005
R1005 source.n647 source.n646 9.3005
R1006 source.n623 source.n622 9.3005
R1007 source.n618 source.n617 9.3005
R1008 source.n629 source.n628 9.3005
R1009 source.n631 source.n630 9.3005
R1010 source.n614 source.n613 9.3005
R1011 source.n637 source.n636 9.3005
R1012 source.n639 source.n638 9.3005
R1013 source.n640 source.n609 9.3005
R1014 source.n598 source.n597 9.3005
R1015 source.n671 source.n670 9.3005
R1016 source.n673 source.n672 9.3005
R1017 source.n594 source.n593 9.3005
R1018 source.n679 source.n678 9.3005
R1019 source.n681 source.n680 9.3005
R1020 source.n590 source.n589 9.3005
R1021 source.n688 source.n687 9.3005
R1022 source.n690 source.n689 9.3005
R1023 source.n713 source.n712 9.3005
R1024 source.n49 source.n48 9.3005
R1025 source.n44 source.n43 9.3005
R1026 source.n55 source.n54 9.3005
R1027 source.n57 source.n56 9.3005
R1028 source.n40 source.n39 9.3005
R1029 source.n63 source.n62 9.3005
R1030 source.n65 source.n64 9.3005
R1031 source.n37 source.n34 9.3005
R1032 source.n96 source.n95 9.3005
R1033 source.n98 source.n97 9.3005
R1034 source.n19 source.n18 9.3005
R1035 source.n104 source.n103 9.3005
R1036 source.n106 source.n105 9.3005
R1037 source.n14 source.n13 9.3005
R1038 source.n112 source.n111 9.3005
R1039 source.n114 source.n113 9.3005
R1040 source.n137 source.n136 9.3005
R1041 source.n2 source.n1 9.3005
R1042 source.n131 source.n130 9.3005
R1043 source.n129 source.n128 9.3005
R1044 source.n6 source.n5 9.3005
R1045 source.n123 source.n122 9.3005
R1046 source.n121 source.n120 9.3005
R1047 source.n10 source.n9 9.3005
R1048 source.n23 source.n22 9.3005
R1049 source.n90 source.n89 9.3005
R1050 source.n88 source.n87 9.3005
R1051 source.n27 source.n26 9.3005
R1052 source.n82 source.n81 9.3005
R1053 source.n80 source.n79 9.3005
R1054 source.n31 source.n30 9.3005
R1055 source.n74 source.n73 9.3005
R1056 source.n72 source.n71 9.3005
R1057 source.n197 source.n196 9.3005
R1058 source.n192 source.n191 9.3005
R1059 source.n203 source.n202 9.3005
R1060 source.n205 source.n204 9.3005
R1061 source.n188 source.n187 9.3005
R1062 source.n211 source.n210 9.3005
R1063 source.n213 source.n212 9.3005
R1064 source.n185 source.n182 9.3005
R1065 source.n244 source.n243 9.3005
R1066 source.n246 source.n245 9.3005
R1067 source.n167 source.n166 9.3005
R1068 source.n252 source.n251 9.3005
R1069 source.n254 source.n253 9.3005
R1070 source.n162 source.n161 9.3005
R1071 source.n260 source.n259 9.3005
R1072 source.n262 source.n261 9.3005
R1073 source.n285 source.n284 9.3005
R1074 source.n150 source.n149 9.3005
R1075 source.n279 source.n278 9.3005
R1076 source.n277 source.n276 9.3005
R1077 source.n154 source.n153 9.3005
R1078 source.n271 source.n270 9.3005
R1079 source.n269 source.n268 9.3005
R1080 source.n158 source.n157 9.3005
R1081 source.n171 source.n170 9.3005
R1082 source.n238 source.n237 9.3005
R1083 source.n236 source.n235 9.3005
R1084 source.n175 source.n174 9.3005
R1085 source.n230 source.n229 9.3005
R1086 source.n228 source.n227 9.3005
R1087 source.n179 source.n178 9.3005
R1088 source.n222 source.n221 9.3005
R1089 source.n220 source.n219 9.3005
R1090 source.n337 source.n336 9.3005
R1091 source.n332 source.n331 9.3005
R1092 source.n343 source.n342 9.3005
R1093 source.n345 source.n344 9.3005
R1094 source.n328 source.n327 9.3005
R1095 source.n351 source.n350 9.3005
R1096 source.n353 source.n352 9.3005
R1097 source.n325 source.n322 9.3005
R1098 source.n384 source.n383 9.3005
R1099 source.n386 source.n385 9.3005
R1100 source.n307 source.n306 9.3005
R1101 source.n392 source.n391 9.3005
R1102 source.n394 source.n393 9.3005
R1103 source.n302 source.n301 9.3005
R1104 source.n400 source.n399 9.3005
R1105 source.n402 source.n401 9.3005
R1106 source.n425 source.n424 9.3005
R1107 source.n290 source.n289 9.3005
R1108 source.n419 source.n418 9.3005
R1109 source.n417 source.n416 9.3005
R1110 source.n294 source.n293 9.3005
R1111 source.n411 source.n410 9.3005
R1112 source.n409 source.n408 9.3005
R1113 source.n298 source.n297 9.3005
R1114 source.n311 source.n310 9.3005
R1115 source.n378 source.n377 9.3005
R1116 source.n376 source.n375 9.3005
R1117 source.n315 source.n314 9.3005
R1118 source.n370 source.n369 9.3005
R1119 source.n368 source.n367 9.3005
R1120 source.n319 source.n318 9.3005
R1121 source.n362 source.n361 9.3005
R1122 source.n360 source.n359 9.3005
R1123 source.n485 source.n484 9.3005
R1124 source.n480 source.n479 9.3005
R1125 source.n491 source.n490 9.3005
R1126 source.n493 source.n492 9.3005
R1127 source.n476 source.n475 9.3005
R1128 source.n499 source.n498 9.3005
R1129 source.n501 source.n500 9.3005
R1130 source.n473 source.n470 9.3005
R1131 source.n532 source.n531 9.3005
R1132 source.n534 source.n533 9.3005
R1133 source.n455 source.n454 9.3005
R1134 source.n540 source.n539 9.3005
R1135 source.n542 source.n541 9.3005
R1136 source.n450 source.n449 9.3005
R1137 source.n548 source.n547 9.3005
R1138 source.n550 source.n549 9.3005
R1139 source.n573 source.n572 9.3005
R1140 source.n438 source.n437 9.3005
R1141 source.n567 source.n566 9.3005
R1142 source.n565 source.n564 9.3005
R1143 source.n442 source.n441 9.3005
R1144 source.n559 source.n558 9.3005
R1145 source.n557 source.n556 9.3005
R1146 source.n446 source.n445 9.3005
R1147 source.n459 source.n458 9.3005
R1148 source.n526 source.n525 9.3005
R1149 source.n524 source.n523 9.3005
R1150 source.n463 source.n462 9.3005
R1151 source.n518 source.n517 9.3005
R1152 source.n516 source.n515 9.3005
R1153 source.n467 source.n466 9.3005
R1154 source.n510 source.n509 9.3005
R1155 source.n508 source.n507 9.3005
R1156 source.n1064 source.n1063 8.92171
R1157 source.n1097 source.n1038 8.92171
R1158 source.n1110 source.n1030 8.92171
R1159 source.n1144 source.n1143 8.92171
R1160 source.n916 source.n915 8.92171
R1161 source.n949 source.n890 8.92171
R1162 source.n962 source.n882 8.92171
R1163 source.n996 source.n995 8.92171
R1164 source.n776 source.n775 8.92171
R1165 source.n809 source.n750 8.92171
R1166 source.n822 source.n742 8.92171
R1167 source.n856 source.n855 8.92171
R1168 source.n628 source.n627 8.92171
R1169 source.n661 source.n602 8.92171
R1170 source.n674 source.n594 8.92171
R1171 source.n708 source.n707 8.92171
R1172 source.n132 source.n131 8.92171
R1173 source.n99 source.n19 8.92171
R1174 source.n86 source.n27 8.92171
R1175 source.n54 source.n53 8.92171
R1176 source.n280 source.n279 8.92171
R1177 source.n247 source.n167 8.92171
R1178 source.n234 source.n175 8.92171
R1179 source.n202 source.n201 8.92171
R1180 source.n420 source.n419 8.92171
R1181 source.n387 source.n307 8.92171
R1182 source.n374 source.n315 8.92171
R1183 source.n342 source.n341 8.92171
R1184 source.n568 source.n567 8.92171
R1185 source.n535 source.n455 8.92171
R1186 source.n522 source.n463 8.92171
R1187 source.n490 source.n489 8.92171
R1188 source.n1060 source.n1054 8.14595
R1189 source.n1098 source.n1036 8.14595
R1190 source.n1109 source.n1032 8.14595
R1191 source.n1147 source.n1014 8.14595
R1192 source.n912 source.n906 8.14595
R1193 source.n950 source.n888 8.14595
R1194 source.n961 source.n884 8.14595
R1195 source.n999 source.n866 8.14595
R1196 source.n772 source.n766 8.14595
R1197 source.n810 source.n748 8.14595
R1198 source.n821 source.n744 8.14595
R1199 source.n859 source.n726 8.14595
R1200 source.n624 source.n618 8.14595
R1201 source.n662 source.n600 8.14595
R1202 source.n673 source.n596 8.14595
R1203 source.n711 source.n578 8.14595
R1204 source.n135 source.n2 8.14595
R1205 source.n98 source.n21 8.14595
R1206 source.n87 source.n25 8.14595
R1207 source.n50 source.n44 8.14595
R1208 source.n283 source.n150 8.14595
R1209 source.n246 source.n169 8.14595
R1210 source.n235 source.n173 8.14595
R1211 source.n198 source.n192 8.14595
R1212 source.n423 source.n290 8.14595
R1213 source.n386 source.n309 8.14595
R1214 source.n375 source.n313 8.14595
R1215 source.n338 source.n332 8.14595
R1216 source.n571 source.n438 8.14595
R1217 source.n534 source.n457 8.14595
R1218 source.n523 source.n461 8.14595
R1219 source.n486 source.n480 8.14595
R1220 source.n1059 source.n1056 7.3702
R1221 source.n1102 source.n1101 7.3702
R1222 source.n1106 source.n1105 7.3702
R1223 source.n1148 source.n1012 7.3702
R1224 source.n911 source.n908 7.3702
R1225 source.n954 source.n953 7.3702
R1226 source.n958 source.n957 7.3702
R1227 source.n1000 source.n864 7.3702
R1228 source.n771 source.n768 7.3702
R1229 source.n814 source.n813 7.3702
R1230 source.n818 source.n817 7.3702
R1231 source.n860 source.n724 7.3702
R1232 source.n623 source.n620 7.3702
R1233 source.n666 source.n665 7.3702
R1234 source.n670 source.n669 7.3702
R1235 source.n712 source.n576 7.3702
R1236 source.n136 source.n0 7.3702
R1237 source.n95 source.n94 7.3702
R1238 source.n91 source.n90 7.3702
R1239 source.n49 source.n46 7.3702
R1240 source.n284 source.n148 7.3702
R1241 source.n243 source.n242 7.3702
R1242 source.n239 source.n238 7.3702
R1243 source.n197 source.n194 7.3702
R1244 source.n424 source.n288 7.3702
R1245 source.n383 source.n382 7.3702
R1246 source.n379 source.n378 7.3702
R1247 source.n337 source.n334 7.3702
R1248 source.n572 source.n436 7.3702
R1249 source.n531 source.n530 7.3702
R1250 source.n527 source.n526 7.3702
R1251 source.n485 source.n482 7.3702
R1252 source.n1102 source.n1034 6.59444
R1253 source.n1105 source.n1034 6.59444
R1254 source.n1150 source.n1012 6.59444
R1255 source.n954 source.n886 6.59444
R1256 source.n957 source.n886 6.59444
R1257 source.n1002 source.n864 6.59444
R1258 source.n814 source.n746 6.59444
R1259 source.n817 source.n746 6.59444
R1260 source.n862 source.n724 6.59444
R1261 source.n666 source.n598 6.59444
R1262 source.n669 source.n598 6.59444
R1263 source.n714 source.n576 6.59444
R1264 source.n138 source.n0 6.59444
R1265 source.n94 source.n23 6.59444
R1266 source.n91 source.n23 6.59444
R1267 source.n286 source.n148 6.59444
R1268 source.n242 source.n171 6.59444
R1269 source.n239 source.n171 6.59444
R1270 source.n426 source.n288 6.59444
R1271 source.n382 source.n311 6.59444
R1272 source.n379 source.n311 6.59444
R1273 source.n574 source.n436 6.59444
R1274 source.n530 source.n459 6.59444
R1275 source.n527 source.n459 6.59444
R1276 source.n1060 source.n1059 5.81868
R1277 source.n1101 source.n1036 5.81868
R1278 source.n1106 source.n1032 5.81868
R1279 source.n1148 source.n1147 5.81868
R1280 source.n912 source.n911 5.81868
R1281 source.n953 source.n888 5.81868
R1282 source.n958 source.n884 5.81868
R1283 source.n1000 source.n999 5.81868
R1284 source.n772 source.n771 5.81868
R1285 source.n813 source.n748 5.81868
R1286 source.n818 source.n744 5.81868
R1287 source.n860 source.n859 5.81868
R1288 source.n624 source.n623 5.81868
R1289 source.n665 source.n600 5.81868
R1290 source.n670 source.n596 5.81868
R1291 source.n712 source.n711 5.81868
R1292 source.n136 source.n135 5.81868
R1293 source.n95 source.n21 5.81868
R1294 source.n90 source.n25 5.81868
R1295 source.n50 source.n49 5.81868
R1296 source.n284 source.n283 5.81868
R1297 source.n243 source.n169 5.81868
R1298 source.n238 source.n173 5.81868
R1299 source.n198 source.n197 5.81868
R1300 source.n424 source.n423 5.81868
R1301 source.n383 source.n309 5.81868
R1302 source.n378 source.n313 5.81868
R1303 source.n338 source.n337 5.81868
R1304 source.n572 source.n571 5.81868
R1305 source.n531 source.n457 5.81868
R1306 source.n526 source.n461 5.81868
R1307 source.n486 source.n485 5.81868
R1308 source.n1152 source.n1151 5.53498
R1309 source.n1063 source.n1054 5.04292
R1310 source.n1098 source.n1097 5.04292
R1311 source.n1110 source.n1109 5.04292
R1312 source.n1144 source.n1014 5.04292
R1313 source.n915 source.n906 5.04292
R1314 source.n950 source.n949 5.04292
R1315 source.n962 source.n961 5.04292
R1316 source.n996 source.n866 5.04292
R1317 source.n775 source.n766 5.04292
R1318 source.n810 source.n809 5.04292
R1319 source.n822 source.n821 5.04292
R1320 source.n856 source.n726 5.04292
R1321 source.n627 source.n618 5.04292
R1322 source.n662 source.n661 5.04292
R1323 source.n674 source.n673 5.04292
R1324 source.n708 source.n578 5.04292
R1325 source.n132 source.n2 5.04292
R1326 source.n99 source.n98 5.04292
R1327 source.n87 source.n86 5.04292
R1328 source.n53 source.n44 5.04292
R1329 source.n280 source.n150 5.04292
R1330 source.n247 source.n246 5.04292
R1331 source.n235 source.n234 5.04292
R1332 source.n201 source.n192 5.04292
R1333 source.n420 source.n290 5.04292
R1334 source.n387 source.n386 5.04292
R1335 source.n375 source.n374 5.04292
R1336 source.n341 source.n332 5.04292
R1337 source.n568 source.n438 5.04292
R1338 source.n535 source.n534 5.04292
R1339 source.n523 source.n522 5.04292
R1340 source.n489 source.n480 5.04292
R1341 source.n1064 source.n1052 4.26717
R1342 source.n1094 source.n1038 4.26717
R1343 source.n1113 source.n1030 4.26717
R1344 source.n1143 source.n1016 4.26717
R1345 source.n916 source.n904 4.26717
R1346 source.n946 source.n890 4.26717
R1347 source.n965 source.n882 4.26717
R1348 source.n995 source.n868 4.26717
R1349 source.n776 source.n764 4.26717
R1350 source.n806 source.n750 4.26717
R1351 source.n825 source.n742 4.26717
R1352 source.n855 source.n728 4.26717
R1353 source.n628 source.n616 4.26717
R1354 source.n658 source.n602 4.26717
R1355 source.n677 source.n594 4.26717
R1356 source.n707 source.n580 4.26717
R1357 source.n131 source.n4 4.26717
R1358 source.n102 source.n19 4.26717
R1359 source.n83 source.n27 4.26717
R1360 source.n54 source.n42 4.26717
R1361 source.n279 source.n152 4.26717
R1362 source.n250 source.n167 4.26717
R1363 source.n231 source.n175 4.26717
R1364 source.n202 source.n190 4.26717
R1365 source.n419 source.n292 4.26717
R1366 source.n390 source.n307 4.26717
R1367 source.n371 source.n315 4.26717
R1368 source.n342 source.n330 4.26717
R1369 source.n567 source.n440 4.26717
R1370 source.n538 source.n455 4.26717
R1371 source.n519 source.n463 4.26717
R1372 source.n490 source.n478 4.26717
R1373 source.n1068 source.n1067 3.49141
R1374 source.n1093 source.n1040 3.49141
R1375 source.n1114 source.n1028 3.49141
R1376 source.n1140 source.n1139 3.49141
R1377 source.n920 source.n919 3.49141
R1378 source.n945 source.n892 3.49141
R1379 source.n966 source.n880 3.49141
R1380 source.n992 source.n991 3.49141
R1381 source.n780 source.n779 3.49141
R1382 source.n805 source.n752 3.49141
R1383 source.n826 source.n740 3.49141
R1384 source.n852 source.n851 3.49141
R1385 source.n632 source.n631 3.49141
R1386 source.n657 source.n604 3.49141
R1387 source.n678 source.n592 3.49141
R1388 source.n704 source.n703 3.49141
R1389 source.n128 source.n127 3.49141
R1390 source.n103 source.n17 3.49141
R1391 source.n82 source.n29 3.49141
R1392 source.n58 source.n57 3.49141
R1393 source.n276 source.n275 3.49141
R1394 source.n251 source.n165 3.49141
R1395 source.n230 source.n177 3.49141
R1396 source.n206 source.n205 3.49141
R1397 source.n416 source.n415 3.49141
R1398 source.n391 source.n305 3.49141
R1399 source.n370 source.n317 3.49141
R1400 source.n346 source.n345 3.49141
R1401 source.n564 source.n563 3.49141
R1402 source.n539 source.n453 3.49141
R1403 source.n518 source.n465 3.49141
R1404 source.n494 source.n493 3.49141
R1405 source.n48 source.n47 2.84303
R1406 source.n196 source.n195 2.84303
R1407 source.n336 source.n335 2.84303
R1408 source.n484 source.n483 2.84303
R1409 source.n1058 source.n1057 2.84303
R1410 source.n910 source.n909 2.84303
R1411 source.n770 source.n769 2.84303
R1412 source.n622 source.n621 2.84303
R1413 source.n1071 source.n1050 2.71565
R1414 source.n1090 source.n1089 2.71565
R1415 source.n1118 source.n1117 2.71565
R1416 source.n1136 source.n1018 2.71565
R1417 source.n923 source.n902 2.71565
R1418 source.n942 source.n941 2.71565
R1419 source.n970 source.n969 2.71565
R1420 source.n988 source.n870 2.71565
R1421 source.n783 source.n762 2.71565
R1422 source.n802 source.n801 2.71565
R1423 source.n830 source.n829 2.71565
R1424 source.n848 source.n730 2.71565
R1425 source.n635 source.n614 2.71565
R1426 source.n654 source.n653 2.71565
R1427 source.n682 source.n681 2.71565
R1428 source.n700 source.n582 2.71565
R1429 source.n124 source.n6 2.71565
R1430 source.n107 source.n106 2.71565
R1431 source.n79 source.n78 2.71565
R1432 source.n61 source.n40 2.71565
R1433 source.n272 source.n154 2.71565
R1434 source.n255 source.n254 2.71565
R1435 source.n227 source.n226 2.71565
R1436 source.n209 source.n188 2.71565
R1437 source.n412 source.n294 2.71565
R1438 source.n395 source.n394 2.71565
R1439 source.n367 source.n366 2.71565
R1440 source.n349 source.n328 2.71565
R1441 source.n560 source.n442 2.71565
R1442 source.n543 source.n542 2.71565
R1443 source.n515 source.n514 2.71565
R1444 source.n497 source.n476 2.71565
R1445 source.n1072 source.n1048 1.93989
R1446 source.n1086 source.n1042 1.93989
R1447 source.n1122 source.n1026 1.93989
R1448 source.n1135 source.n1020 1.93989
R1449 source.n924 source.n900 1.93989
R1450 source.n938 source.n894 1.93989
R1451 source.n974 source.n878 1.93989
R1452 source.n987 source.n872 1.93989
R1453 source.n784 source.n760 1.93989
R1454 source.n798 source.n754 1.93989
R1455 source.n834 source.n738 1.93989
R1456 source.n847 source.n732 1.93989
R1457 source.n636 source.n612 1.93989
R1458 source.n650 source.n606 1.93989
R1459 source.n686 source.n590 1.93989
R1460 source.n699 source.n584 1.93989
R1461 source.n123 source.n8 1.93989
R1462 source.n110 source.n14 1.93989
R1463 source.n75 source.n31 1.93989
R1464 source.n62 source.n38 1.93989
R1465 source.n271 source.n156 1.93989
R1466 source.n258 source.n162 1.93989
R1467 source.n223 source.n179 1.93989
R1468 source.n210 source.n186 1.93989
R1469 source.n411 source.n296 1.93989
R1470 source.n398 source.n302 1.93989
R1471 source.n363 source.n319 1.93989
R1472 source.n350 source.n326 1.93989
R1473 source.n559 source.n444 1.93989
R1474 source.n546 source.n450 1.93989
R1475 source.n511 source.n467 1.93989
R1476 source.n498 source.n474 1.93989
R1477 source.n1077 source.n1075 1.16414
R1478 source.n1085 source.n1044 1.16414
R1479 source.n1123 source.n1024 1.16414
R1480 source.n1132 source.n1131 1.16414
R1481 source.n929 source.n927 1.16414
R1482 source.n937 source.n896 1.16414
R1483 source.n975 source.n876 1.16414
R1484 source.n984 source.n983 1.16414
R1485 source.n789 source.n787 1.16414
R1486 source.n797 source.n756 1.16414
R1487 source.n835 source.n736 1.16414
R1488 source.n844 source.n843 1.16414
R1489 source.n641 source.n639 1.16414
R1490 source.n649 source.n608 1.16414
R1491 source.n687 source.n588 1.16414
R1492 source.n696 source.n695 1.16414
R1493 source.n120 source.n119 1.16414
R1494 source.n111 source.n12 1.16414
R1495 source.n74 source.n33 1.16414
R1496 source.n66 source.n65 1.16414
R1497 source.n268 source.n267 1.16414
R1498 source.n259 source.n160 1.16414
R1499 source.n222 source.n181 1.16414
R1500 source.n214 source.n213 1.16414
R1501 source.n408 source.n407 1.16414
R1502 source.n399 source.n300 1.16414
R1503 source.n362 source.n321 1.16414
R1504 source.n354 source.n353 1.16414
R1505 source.n556 source.n555 1.16414
R1506 source.n547 source.n448 1.16414
R1507 source.n510 source.n469 1.16414
R1508 source.n502 source.n501 1.16414
R1509 source.n1010 source.t15 0.7925
R1510 source.n1010 source.t6 0.7925
R1511 source.n1008 source.t17 0.7925
R1512 source.n1008 source.t39 0.7925
R1513 source.n1006 source.t16 0.7925
R1514 source.n1006 source.t3 0.7925
R1515 source.n1004 source.t10 0.7925
R1516 source.n1004 source.t11 0.7925
R1517 source.n722 source.t36 0.7925
R1518 source.n722 source.t24 0.7925
R1519 source.n720 source.t22 0.7925
R1520 source.n720 source.t27 0.7925
R1521 source.n718 source.t21 0.7925
R1522 source.n718 source.t25 0.7925
R1523 source.n716 source.t30 0.7925
R1524 source.n716 source.t29 0.7925
R1525 source.n140 source.t31 0.7925
R1526 source.n140 source.t19 0.7925
R1527 source.n142 source.t18 0.7925
R1528 source.n142 source.t33 0.7925
R1529 source.n144 source.t34 0.7925
R1530 source.n144 source.t20 0.7925
R1531 source.n146 source.t28 0.7925
R1532 source.n146 source.t32 0.7925
R1533 source.n428 source.t1 0.7925
R1534 source.n428 source.t5 0.7925
R1535 source.n430 source.t12 0.7925
R1536 source.n430 source.t0 0.7925
R1537 source.n432 source.t9 0.7925
R1538 source.n432 source.t8 0.7925
R1539 source.n434 source.t4 0.7925
R1540 source.n434 source.t7 0.7925
R1541 source.n575 source.n435 0.543603
R1542 source.n435 source.n433 0.543603
R1543 source.n433 source.n431 0.543603
R1544 source.n431 source.n429 0.543603
R1545 source.n429 source.n427 0.543603
R1546 source.n287 source.n147 0.543603
R1547 source.n147 source.n145 0.543603
R1548 source.n145 source.n143 0.543603
R1549 source.n143 source.n141 0.543603
R1550 source.n141 source.n139 0.543603
R1551 source.n717 source.n715 0.543603
R1552 source.n719 source.n717 0.543603
R1553 source.n721 source.n719 0.543603
R1554 source.n723 source.n721 0.543603
R1555 source.n863 source.n723 0.543603
R1556 source.n1005 source.n1003 0.543603
R1557 source.n1007 source.n1005 0.543603
R1558 source.n1009 source.n1007 0.543603
R1559 source.n1011 source.n1009 0.543603
R1560 source.n1151 source.n1011 0.543603
R1561 source.n427 source.n287 0.470328
R1562 source.n1003 source.n863 0.470328
R1563 source.n1076 source.n1046 0.388379
R1564 source.n1082 source.n1081 0.388379
R1565 source.n1127 source.n1126 0.388379
R1566 source.n1128 source.n1022 0.388379
R1567 source.n928 source.n898 0.388379
R1568 source.n934 source.n933 0.388379
R1569 source.n979 source.n978 0.388379
R1570 source.n980 source.n874 0.388379
R1571 source.n788 source.n758 0.388379
R1572 source.n794 source.n793 0.388379
R1573 source.n839 source.n838 0.388379
R1574 source.n840 source.n734 0.388379
R1575 source.n640 source.n610 0.388379
R1576 source.n646 source.n645 0.388379
R1577 source.n691 source.n690 0.388379
R1578 source.n692 source.n586 0.388379
R1579 source.n116 source.n10 0.388379
R1580 source.n115 source.n114 0.388379
R1581 source.n71 source.n70 0.388379
R1582 source.n37 source.n35 0.388379
R1583 source.n264 source.n158 0.388379
R1584 source.n263 source.n262 0.388379
R1585 source.n219 source.n218 0.388379
R1586 source.n185 source.n183 0.388379
R1587 source.n404 source.n298 0.388379
R1588 source.n403 source.n402 0.388379
R1589 source.n359 source.n358 0.388379
R1590 source.n325 source.n323 0.388379
R1591 source.n552 source.n446 0.388379
R1592 source.n551 source.n550 0.388379
R1593 source.n507 source.n506 0.388379
R1594 source.n473 source.n471 0.388379
R1595 source source.n1152 0.188
R1596 source.n1058 source.n1053 0.155672
R1597 source.n1065 source.n1053 0.155672
R1598 source.n1066 source.n1065 0.155672
R1599 source.n1066 source.n1049 0.155672
R1600 source.n1073 source.n1049 0.155672
R1601 source.n1074 source.n1073 0.155672
R1602 source.n1074 source.n1045 0.155672
R1603 source.n1083 source.n1045 0.155672
R1604 source.n1084 source.n1083 0.155672
R1605 source.n1084 source.n1041 0.155672
R1606 source.n1091 source.n1041 0.155672
R1607 source.n1092 source.n1091 0.155672
R1608 source.n1092 source.n1037 0.155672
R1609 source.n1099 source.n1037 0.155672
R1610 source.n1100 source.n1099 0.155672
R1611 source.n1100 source.n1033 0.155672
R1612 source.n1107 source.n1033 0.155672
R1613 source.n1108 source.n1107 0.155672
R1614 source.n1108 source.n1029 0.155672
R1615 source.n1115 source.n1029 0.155672
R1616 source.n1116 source.n1115 0.155672
R1617 source.n1116 source.n1025 0.155672
R1618 source.n1124 source.n1025 0.155672
R1619 source.n1125 source.n1124 0.155672
R1620 source.n1125 source.n1021 0.155672
R1621 source.n1133 source.n1021 0.155672
R1622 source.n1134 source.n1133 0.155672
R1623 source.n1134 source.n1017 0.155672
R1624 source.n1141 source.n1017 0.155672
R1625 source.n1142 source.n1141 0.155672
R1626 source.n1142 source.n1013 0.155672
R1627 source.n1149 source.n1013 0.155672
R1628 source.n910 source.n905 0.155672
R1629 source.n917 source.n905 0.155672
R1630 source.n918 source.n917 0.155672
R1631 source.n918 source.n901 0.155672
R1632 source.n925 source.n901 0.155672
R1633 source.n926 source.n925 0.155672
R1634 source.n926 source.n897 0.155672
R1635 source.n935 source.n897 0.155672
R1636 source.n936 source.n935 0.155672
R1637 source.n936 source.n893 0.155672
R1638 source.n943 source.n893 0.155672
R1639 source.n944 source.n943 0.155672
R1640 source.n944 source.n889 0.155672
R1641 source.n951 source.n889 0.155672
R1642 source.n952 source.n951 0.155672
R1643 source.n952 source.n885 0.155672
R1644 source.n959 source.n885 0.155672
R1645 source.n960 source.n959 0.155672
R1646 source.n960 source.n881 0.155672
R1647 source.n967 source.n881 0.155672
R1648 source.n968 source.n967 0.155672
R1649 source.n968 source.n877 0.155672
R1650 source.n976 source.n877 0.155672
R1651 source.n977 source.n976 0.155672
R1652 source.n977 source.n873 0.155672
R1653 source.n985 source.n873 0.155672
R1654 source.n986 source.n985 0.155672
R1655 source.n986 source.n869 0.155672
R1656 source.n993 source.n869 0.155672
R1657 source.n994 source.n993 0.155672
R1658 source.n994 source.n865 0.155672
R1659 source.n1001 source.n865 0.155672
R1660 source.n770 source.n765 0.155672
R1661 source.n777 source.n765 0.155672
R1662 source.n778 source.n777 0.155672
R1663 source.n778 source.n761 0.155672
R1664 source.n785 source.n761 0.155672
R1665 source.n786 source.n785 0.155672
R1666 source.n786 source.n757 0.155672
R1667 source.n795 source.n757 0.155672
R1668 source.n796 source.n795 0.155672
R1669 source.n796 source.n753 0.155672
R1670 source.n803 source.n753 0.155672
R1671 source.n804 source.n803 0.155672
R1672 source.n804 source.n749 0.155672
R1673 source.n811 source.n749 0.155672
R1674 source.n812 source.n811 0.155672
R1675 source.n812 source.n745 0.155672
R1676 source.n819 source.n745 0.155672
R1677 source.n820 source.n819 0.155672
R1678 source.n820 source.n741 0.155672
R1679 source.n827 source.n741 0.155672
R1680 source.n828 source.n827 0.155672
R1681 source.n828 source.n737 0.155672
R1682 source.n836 source.n737 0.155672
R1683 source.n837 source.n836 0.155672
R1684 source.n837 source.n733 0.155672
R1685 source.n845 source.n733 0.155672
R1686 source.n846 source.n845 0.155672
R1687 source.n846 source.n729 0.155672
R1688 source.n853 source.n729 0.155672
R1689 source.n854 source.n853 0.155672
R1690 source.n854 source.n725 0.155672
R1691 source.n861 source.n725 0.155672
R1692 source.n622 source.n617 0.155672
R1693 source.n629 source.n617 0.155672
R1694 source.n630 source.n629 0.155672
R1695 source.n630 source.n613 0.155672
R1696 source.n637 source.n613 0.155672
R1697 source.n638 source.n637 0.155672
R1698 source.n638 source.n609 0.155672
R1699 source.n647 source.n609 0.155672
R1700 source.n648 source.n647 0.155672
R1701 source.n648 source.n605 0.155672
R1702 source.n655 source.n605 0.155672
R1703 source.n656 source.n655 0.155672
R1704 source.n656 source.n601 0.155672
R1705 source.n663 source.n601 0.155672
R1706 source.n664 source.n663 0.155672
R1707 source.n664 source.n597 0.155672
R1708 source.n671 source.n597 0.155672
R1709 source.n672 source.n671 0.155672
R1710 source.n672 source.n593 0.155672
R1711 source.n679 source.n593 0.155672
R1712 source.n680 source.n679 0.155672
R1713 source.n680 source.n589 0.155672
R1714 source.n688 source.n589 0.155672
R1715 source.n689 source.n688 0.155672
R1716 source.n689 source.n585 0.155672
R1717 source.n697 source.n585 0.155672
R1718 source.n698 source.n697 0.155672
R1719 source.n698 source.n581 0.155672
R1720 source.n705 source.n581 0.155672
R1721 source.n706 source.n705 0.155672
R1722 source.n706 source.n577 0.155672
R1723 source.n713 source.n577 0.155672
R1724 source.n137 source.n1 0.155672
R1725 source.n130 source.n1 0.155672
R1726 source.n130 source.n129 0.155672
R1727 source.n129 source.n5 0.155672
R1728 source.n122 source.n5 0.155672
R1729 source.n122 source.n121 0.155672
R1730 source.n121 source.n9 0.155672
R1731 source.n113 source.n9 0.155672
R1732 source.n113 source.n112 0.155672
R1733 source.n112 source.n13 0.155672
R1734 source.n105 source.n13 0.155672
R1735 source.n105 source.n104 0.155672
R1736 source.n104 source.n18 0.155672
R1737 source.n97 source.n18 0.155672
R1738 source.n97 source.n96 0.155672
R1739 source.n96 source.n22 0.155672
R1740 source.n89 source.n22 0.155672
R1741 source.n89 source.n88 0.155672
R1742 source.n88 source.n26 0.155672
R1743 source.n81 source.n26 0.155672
R1744 source.n81 source.n80 0.155672
R1745 source.n80 source.n30 0.155672
R1746 source.n73 source.n30 0.155672
R1747 source.n73 source.n72 0.155672
R1748 source.n72 source.n34 0.155672
R1749 source.n64 source.n34 0.155672
R1750 source.n64 source.n63 0.155672
R1751 source.n63 source.n39 0.155672
R1752 source.n56 source.n39 0.155672
R1753 source.n56 source.n55 0.155672
R1754 source.n55 source.n43 0.155672
R1755 source.n48 source.n43 0.155672
R1756 source.n285 source.n149 0.155672
R1757 source.n278 source.n149 0.155672
R1758 source.n278 source.n277 0.155672
R1759 source.n277 source.n153 0.155672
R1760 source.n270 source.n153 0.155672
R1761 source.n270 source.n269 0.155672
R1762 source.n269 source.n157 0.155672
R1763 source.n261 source.n157 0.155672
R1764 source.n261 source.n260 0.155672
R1765 source.n260 source.n161 0.155672
R1766 source.n253 source.n161 0.155672
R1767 source.n253 source.n252 0.155672
R1768 source.n252 source.n166 0.155672
R1769 source.n245 source.n166 0.155672
R1770 source.n245 source.n244 0.155672
R1771 source.n244 source.n170 0.155672
R1772 source.n237 source.n170 0.155672
R1773 source.n237 source.n236 0.155672
R1774 source.n236 source.n174 0.155672
R1775 source.n229 source.n174 0.155672
R1776 source.n229 source.n228 0.155672
R1777 source.n228 source.n178 0.155672
R1778 source.n221 source.n178 0.155672
R1779 source.n221 source.n220 0.155672
R1780 source.n220 source.n182 0.155672
R1781 source.n212 source.n182 0.155672
R1782 source.n212 source.n211 0.155672
R1783 source.n211 source.n187 0.155672
R1784 source.n204 source.n187 0.155672
R1785 source.n204 source.n203 0.155672
R1786 source.n203 source.n191 0.155672
R1787 source.n196 source.n191 0.155672
R1788 source.n425 source.n289 0.155672
R1789 source.n418 source.n289 0.155672
R1790 source.n418 source.n417 0.155672
R1791 source.n417 source.n293 0.155672
R1792 source.n410 source.n293 0.155672
R1793 source.n410 source.n409 0.155672
R1794 source.n409 source.n297 0.155672
R1795 source.n401 source.n297 0.155672
R1796 source.n401 source.n400 0.155672
R1797 source.n400 source.n301 0.155672
R1798 source.n393 source.n301 0.155672
R1799 source.n393 source.n392 0.155672
R1800 source.n392 source.n306 0.155672
R1801 source.n385 source.n306 0.155672
R1802 source.n385 source.n384 0.155672
R1803 source.n384 source.n310 0.155672
R1804 source.n377 source.n310 0.155672
R1805 source.n377 source.n376 0.155672
R1806 source.n376 source.n314 0.155672
R1807 source.n369 source.n314 0.155672
R1808 source.n369 source.n368 0.155672
R1809 source.n368 source.n318 0.155672
R1810 source.n361 source.n318 0.155672
R1811 source.n361 source.n360 0.155672
R1812 source.n360 source.n322 0.155672
R1813 source.n352 source.n322 0.155672
R1814 source.n352 source.n351 0.155672
R1815 source.n351 source.n327 0.155672
R1816 source.n344 source.n327 0.155672
R1817 source.n344 source.n343 0.155672
R1818 source.n343 source.n331 0.155672
R1819 source.n336 source.n331 0.155672
R1820 source.n573 source.n437 0.155672
R1821 source.n566 source.n437 0.155672
R1822 source.n566 source.n565 0.155672
R1823 source.n565 source.n441 0.155672
R1824 source.n558 source.n441 0.155672
R1825 source.n558 source.n557 0.155672
R1826 source.n557 source.n445 0.155672
R1827 source.n549 source.n445 0.155672
R1828 source.n549 source.n548 0.155672
R1829 source.n548 source.n449 0.155672
R1830 source.n541 source.n449 0.155672
R1831 source.n541 source.n540 0.155672
R1832 source.n540 source.n454 0.155672
R1833 source.n533 source.n454 0.155672
R1834 source.n533 source.n532 0.155672
R1835 source.n532 source.n458 0.155672
R1836 source.n525 source.n458 0.155672
R1837 source.n525 source.n524 0.155672
R1838 source.n524 source.n462 0.155672
R1839 source.n517 source.n462 0.155672
R1840 source.n517 source.n516 0.155672
R1841 source.n516 source.n466 0.155672
R1842 source.n509 source.n466 0.155672
R1843 source.n509 source.n508 0.155672
R1844 source.n508 source.n470 0.155672
R1845 source.n500 source.n470 0.155672
R1846 source.n500 source.n499 0.155672
R1847 source.n499 source.n475 0.155672
R1848 source.n492 source.n475 0.155672
R1849 source.n492 source.n491 0.155672
R1850 source.n491 source.n479 0.155672
R1851 source.n484 source.n479 0.155672
R1852 drain_left.n6 drain_left.n4 59.2585
R1853 drain_left.n2 drain_left.n0 59.2585
R1854 drain_left.n10 drain_left.n8 59.2585
R1855 drain_left.n7 drain_left.n3 58.7154
R1856 drain_left.n6 drain_left.n5 58.7154
R1857 drain_left.n2 drain_left.n1 58.7154
R1858 drain_left.n14 drain_left.n13 58.7154
R1859 drain_left.n12 drain_left.n11 58.7154
R1860 drain_left.n10 drain_left.n9 58.7154
R1861 drain_left.n16 drain_left.n15 58.7153
R1862 drain_left drain_left.n7 41.5604
R1863 drain_left drain_left.n16 6.19632
R1864 drain_left.n3 drain_left.t7 0.7925
R1865 drain_left.n3 drain_left.t16 0.7925
R1866 drain_left.n4 drain_left.t11 0.7925
R1867 drain_left.n4 drain_left.t1 0.7925
R1868 drain_left.n5 drain_left.t9 0.7925
R1869 drain_left.n5 drain_left.t0 0.7925
R1870 drain_left.n1 drain_left.t5 0.7925
R1871 drain_left.n1 drain_left.t15 0.7925
R1872 drain_left.n0 drain_left.t4 0.7925
R1873 drain_left.n0 drain_left.t17 0.7925
R1874 drain_left.n15 drain_left.t12 0.7925
R1875 drain_left.n15 drain_left.t6 0.7925
R1876 drain_left.n13 drain_left.t3 0.7925
R1877 drain_left.n13 drain_left.t19 0.7925
R1878 drain_left.n11 drain_left.t14 0.7925
R1879 drain_left.n11 drain_left.t10 0.7925
R1880 drain_left.n9 drain_left.t8 0.7925
R1881 drain_left.n9 drain_left.t2 0.7925
R1882 drain_left.n8 drain_left.t18 0.7925
R1883 drain_left.n8 drain_left.t13 0.7925
R1884 drain_left.n12 drain_left.n10 0.543603
R1885 drain_left.n14 drain_left.n12 0.543603
R1886 drain_left.n16 drain_left.n14 0.543603
R1887 drain_left.n7 drain_left.n6 0.488257
R1888 drain_left.n7 drain_left.n2 0.488257
R1889 minus.n27 minus.t7 2161.7
R1890 minus.n7 minus.t11 2161.7
R1891 minus.n56 minus.t5 2161.7
R1892 minus.n35 minus.t4 2161.7
R1893 minus.n26 minus.t2 2112.77
R1894 minus.n24 minus.t18 2112.77
R1895 minus.n3 minus.t6 2112.77
R1896 minus.n18 minus.t0 2112.77
R1897 minus.n16 minus.t15 2112.77
R1898 minus.n4 minus.t10 2112.77
R1899 minus.n10 minus.t1 2112.77
R1900 minus.n6 minus.t17 2112.77
R1901 minus.n55 minus.t14 2112.77
R1902 minus.n53 minus.t16 2112.77
R1903 minus.n47 minus.t8 2112.77
R1904 minus.n46 minus.t19 2112.77
R1905 minus.n44 minus.t9 2112.77
R1906 minus.n32 minus.t12 2112.77
R1907 minus.n38 minus.t3 2112.77
R1908 minus.n34 minus.t13 2112.77
R1909 minus.n8 minus.n7 161.489
R1910 minus.n36 minus.n35 161.489
R1911 minus.n28 minus.n27 161.3
R1912 minus.n25 minus.n0 161.3
R1913 minus.n23 minus.n22 161.3
R1914 minus.n21 minus.n1 161.3
R1915 minus.n20 minus.n19 161.3
R1916 minus.n17 minus.n2 161.3
R1917 minus.n15 minus.n14 161.3
R1918 minus.n13 minus.n12 161.3
R1919 minus.n11 minus.n5 161.3
R1920 minus.n9 minus.n8 161.3
R1921 minus.n57 minus.n56 161.3
R1922 minus.n54 minus.n29 161.3
R1923 minus.n52 minus.n51 161.3
R1924 minus.n50 minus.n30 161.3
R1925 minus.n49 minus.n48 161.3
R1926 minus.n45 minus.n31 161.3
R1927 minus.n43 minus.n42 161.3
R1928 minus.n41 minus.n40 161.3
R1929 minus.n39 minus.n33 161.3
R1930 minus.n37 minus.n36 161.3
R1931 minus.n23 minus.n1 73.0308
R1932 minus.n12 minus.n11 73.0308
R1933 minus.n40 minus.n39 73.0308
R1934 minus.n52 minus.n30 73.0308
R1935 minus.n19 minus.n3 64.9975
R1936 minus.n15 minus.n4 64.9975
R1937 minus.n43 minus.n32 64.9975
R1938 minus.n48 minus.n47 64.9975
R1939 minus.n25 minus.n24 62.0763
R1940 minus.n10 minus.n9 62.0763
R1941 minus.n38 minus.n37 62.0763
R1942 minus.n54 minus.n53 62.0763
R1943 minus.n58 minus.n28 46.9475
R1944 minus.n18 minus.n17 46.0096
R1945 minus.n17 minus.n16 46.0096
R1946 minus.n45 minus.n44 46.0096
R1947 minus.n46 minus.n45 46.0096
R1948 minus.n27 minus.n26 43.0884
R1949 minus.n7 minus.n6 43.0884
R1950 minus.n35 minus.n34 43.0884
R1951 minus.n56 minus.n55 43.0884
R1952 minus.n26 minus.n25 29.9429
R1953 minus.n9 minus.n6 29.9429
R1954 minus.n37 minus.n34 29.9429
R1955 minus.n55 minus.n54 29.9429
R1956 minus.n19 minus.n18 27.0217
R1957 minus.n16 minus.n15 27.0217
R1958 minus.n44 minus.n43 27.0217
R1959 minus.n48 minus.n46 27.0217
R1960 minus.n24 minus.n23 10.955
R1961 minus.n11 minus.n10 10.955
R1962 minus.n39 minus.n38 10.955
R1963 minus.n53 minus.n52 10.955
R1964 minus.n3 minus.n1 8.03383
R1965 minus.n12 minus.n4 8.03383
R1966 minus.n40 minus.n32 8.03383
R1967 minus.n47 minus.n30 8.03383
R1968 minus.n58 minus.n57 6.51565
R1969 minus.n28 minus.n0 0.189894
R1970 minus.n22 minus.n0 0.189894
R1971 minus.n22 minus.n21 0.189894
R1972 minus.n21 minus.n20 0.189894
R1973 minus.n20 minus.n2 0.189894
R1974 minus.n14 minus.n2 0.189894
R1975 minus.n14 minus.n13 0.189894
R1976 minus.n13 minus.n5 0.189894
R1977 minus.n8 minus.n5 0.189894
R1978 minus.n36 minus.n33 0.189894
R1979 minus.n41 minus.n33 0.189894
R1980 minus.n42 minus.n41 0.189894
R1981 minus.n42 minus.n31 0.189894
R1982 minus.n49 minus.n31 0.189894
R1983 minus.n50 minus.n49 0.189894
R1984 minus.n51 minus.n50 0.189894
R1985 minus.n51 minus.n29 0.189894
R1986 minus.n57 minus.n29 0.189894
R1987 minus minus.n58 0.188
R1988 drain_right.n6 drain_right.n4 59.2585
R1989 drain_right.n2 drain_right.n0 59.2585
R1990 drain_right.n10 drain_right.n8 59.2584
R1991 drain_right.n7 drain_right.n3 58.7154
R1992 drain_right.n6 drain_right.n5 58.7154
R1993 drain_right.n2 drain_right.n1 58.7154
R1994 drain_right.n10 drain_right.n9 58.7154
R1995 drain_right.n12 drain_right.n11 58.7154
R1996 drain_right.n14 drain_right.n13 58.7154
R1997 drain_right.n16 drain_right.n15 58.7154
R1998 drain_right drain_right.n7 41.0072
R1999 drain_right drain_right.n16 6.19632
R2000 drain_right.n3 drain_right.t10 0.7925
R2001 drain_right.n3 drain_right.t0 0.7925
R2002 drain_right.n4 drain_right.t5 0.7925
R2003 drain_right.n4 drain_right.t14 0.7925
R2004 drain_right.n5 drain_right.t11 0.7925
R2005 drain_right.n5 drain_right.t3 0.7925
R2006 drain_right.n1 drain_right.t16 0.7925
R2007 drain_right.n1 drain_right.t7 0.7925
R2008 drain_right.n0 drain_right.t15 0.7925
R2009 drain_right.n0 drain_right.t6 0.7925
R2010 drain_right.n8 drain_right.t2 0.7925
R2011 drain_right.n8 drain_right.t8 0.7925
R2012 drain_right.n9 drain_right.t9 0.7925
R2013 drain_right.n9 drain_right.t18 0.7925
R2014 drain_right.n11 drain_right.t19 0.7925
R2015 drain_right.n11 drain_right.t4 0.7925
R2016 drain_right.n13 drain_right.t1 0.7925
R2017 drain_right.n13 drain_right.t13 0.7925
R2018 drain_right.n15 drain_right.t12 0.7925
R2019 drain_right.n15 drain_right.t17 0.7925
R2020 drain_right.n16 drain_right.n14 0.543603
R2021 drain_right.n14 drain_right.n12 0.543603
R2022 drain_right.n12 drain_right.n10 0.543603
R2023 drain_right.n7 drain_right.n6 0.488257
R2024 drain_right.n7 drain_right.n2 0.488257
C0 drain_left minus 0.171748f
C1 plus minus 8.18185f
C2 plus drain_left 14.509f
C3 drain_right minus 14.3031f
C4 source minus 13.519199f
C5 drain_right drain_left 1.10832f
C6 drain_right plus 0.36079f
C7 source drain_left 74.4487f
C8 source plus 13.533299f
C9 source drain_right 74.4491f
C10 drain_right a_n2102_n5888# 9.66289f
C11 drain_left a_n2102_n5888# 9.98152f
C12 source a_n2102_n5888# 15.784036f
C13 minus a_n2102_n5888# 9.121881f
C14 plus a_n2102_n5888# 11.96322f
C15 drain_right.t15 a_n2102_n5888# 0.680743f
C16 drain_right.t6 a_n2102_n5888# 0.680743f
C17 drain_right.n0 a_n2102_n5888# 6.27768f
C18 drain_right.t16 a_n2102_n5888# 0.680743f
C19 drain_right.t7 a_n2102_n5888# 0.680743f
C20 drain_right.n1 a_n2102_n5888# 6.27378f
C21 drain_right.n2 a_n2102_n5888# 0.829215f
C22 drain_right.t10 a_n2102_n5888# 0.680743f
C23 drain_right.t0 a_n2102_n5888# 0.680743f
C24 drain_right.n3 a_n2102_n5888# 6.27378f
C25 drain_right.t5 a_n2102_n5888# 0.680743f
C26 drain_right.t14 a_n2102_n5888# 0.680743f
C27 drain_right.n4 a_n2102_n5888# 6.27768f
C28 drain_right.t11 a_n2102_n5888# 0.680743f
C29 drain_right.t3 a_n2102_n5888# 0.680743f
C30 drain_right.n5 a_n2102_n5888# 6.27378f
C31 drain_right.n6 a_n2102_n5888# 0.829215f
C32 drain_right.n7 a_n2102_n5888# 3.19274f
C33 drain_right.t2 a_n2102_n5888# 0.680743f
C34 drain_right.t8 a_n2102_n5888# 0.680743f
C35 drain_right.n8 a_n2102_n5888# 6.27767f
C36 drain_right.t9 a_n2102_n5888# 0.680743f
C37 drain_right.t18 a_n2102_n5888# 0.680743f
C38 drain_right.n9 a_n2102_n5888# 6.27378f
C39 drain_right.n10 a_n2102_n5888# 0.833734f
C40 drain_right.t19 a_n2102_n5888# 0.680743f
C41 drain_right.t4 a_n2102_n5888# 0.680743f
C42 drain_right.n11 a_n2102_n5888# 6.27378f
C43 drain_right.n12 a_n2102_n5888# 0.411871f
C44 drain_right.t1 a_n2102_n5888# 0.680743f
C45 drain_right.t13 a_n2102_n5888# 0.680743f
C46 drain_right.n13 a_n2102_n5888# 6.27378f
C47 drain_right.n14 a_n2102_n5888# 0.411871f
C48 drain_right.t12 a_n2102_n5888# 0.680743f
C49 drain_right.t17 a_n2102_n5888# 0.680743f
C50 drain_right.n15 a_n2102_n5888# 6.27378f
C51 drain_right.n16 a_n2102_n5888# 0.698685f
C52 minus.n0 a_n2102_n5888# 0.0496f
C53 minus.t7 a_n2102_n5888# 1.05541f
C54 minus.t2 a_n2102_n5888# 1.04669f
C55 minus.t18 a_n2102_n5888# 1.04669f
C56 minus.n1 a_n2102_n5888# 0.018136f
C57 minus.n2 a_n2102_n5888# 0.0496f
C58 minus.t6 a_n2102_n5888# 1.04669f
C59 minus.n3 a_n2102_n5888# 0.380868f
C60 minus.t0 a_n2102_n5888# 1.04669f
C61 minus.t15 a_n2102_n5888# 1.04669f
C62 minus.t10 a_n2102_n5888# 1.04669f
C63 minus.n4 a_n2102_n5888# 0.380868f
C64 minus.n5 a_n2102_n5888# 0.0496f
C65 minus.t1 a_n2102_n5888# 1.04669f
C66 minus.t17 a_n2102_n5888# 1.04669f
C67 minus.n6 a_n2102_n5888# 0.380868f
C68 minus.t11 a_n2102_n5888# 1.05541f
C69 minus.n7 a_n2102_n5888# 0.396787f
C70 minus.n8 a_n2102_n5888# 0.113498f
C71 minus.n9 a_n2102_n5888# 0.020429f
C72 minus.n10 a_n2102_n5888# 0.380868f
C73 minus.n11 a_n2102_n5888# 0.018748f
C74 minus.n12 a_n2102_n5888# 0.018136f
C75 minus.n13 a_n2102_n5888# 0.0496f
C76 minus.n14 a_n2102_n5888# 0.0496f
C77 minus.n15 a_n2102_n5888# 0.020429f
C78 minus.n16 a_n2102_n5888# 0.380868f
C79 minus.n17 a_n2102_n5888# 0.020429f
C80 minus.n18 a_n2102_n5888# 0.380868f
C81 minus.n19 a_n2102_n5888# 0.020429f
C82 minus.n20 a_n2102_n5888# 0.0496f
C83 minus.n21 a_n2102_n5888# 0.0496f
C84 minus.n22 a_n2102_n5888# 0.0496f
C85 minus.n23 a_n2102_n5888# 0.018748f
C86 minus.n24 a_n2102_n5888# 0.380868f
C87 minus.n25 a_n2102_n5888# 0.020429f
C88 minus.n26 a_n2102_n5888# 0.380868f
C89 minus.n27 a_n2102_n5888# 0.396712f
C90 minus.n28 a_n2102_n5888# 2.58004f
C91 minus.n29 a_n2102_n5888# 0.0496f
C92 minus.t14 a_n2102_n5888# 1.04669f
C93 minus.t16 a_n2102_n5888# 1.04669f
C94 minus.n30 a_n2102_n5888# 0.018136f
C95 minus.n31 a_n2102_n5888# 0.0496f
C96 minus.t19 a_n2102_n5888# 1.04669f
C97 minus.t9 a_n2102_n5888# 1.04669f
C98 minus.t12 a_n2102_n5888# 1.04669f
C99 minus.n32 a_n2102_n5888# 0.380868f
C100 minus.n33 a_n2102_n5888# 0.0496f
C101 minus.t3 a_n2102_n5888# 1.04669f
C102 minus.t13 a_n2102_n5888# 1.04669f
C103 minus.n34 a_n2102_n5888# 0.380868f
C104 minus.t4 a_n2102_n5888# 1.05541f
C105 minus.n35 a_n2102_n5888# 0.396787f
C106 minus.n36 a_n2102_n5888# 0.113498f
C107 minus.n37 a_n2102_n5888# 0.020429f
C108 minus.n38 a_n2102_n5888# 0.380868f
C109 minus.n39 a_n2102_n5888# 0.018748f
C110 minus.n40 a_n2102_n5888# 0.018136f
C111 minus.n41 a_n2102_n5888# 0.0496f
C112 minus.n42 a_n2102_n5888# 0.0496f
C113 minus.n43 a_n2102_n5888# 0.020429f
C114 minus.n44 a_n2102_n5888# 0.380868f
C115 minus.n45 a_n2102_n5888# 0.020429f
C116 minus.n46 a_n2102_n5888# 0.380868f
C117 minus.t8 a_n2102_n5888# 1.04669f
C118 minus.n47 a_n2102_n5888# 0.380868f
C119 minus.n48 a_n2102_n5888# 0.020429f
C120 minus.n49 a_n2102_n5888# 0.0496f
C121 minus.n50 a_n2102_n5888# 0.0496f
C122 minus.n51 a_n2102_n5888# 0.0496f
C123 minus.n52 a_n2102_n5888# 0.018748f
C124 minus.n53 a_n2102_n5888# 0.380868f
C125 minus.n54 a_n2102_n5888# 0.020429f
C126 minus.n55 a_n2102_n5888# 0.380868f
C127 minus.t5 a_n2102_n5888# 1.05541f
C128 minus.n56 a_n2102_n5888# 0.396712f
C129 minus.n57 a_n2102_n5888# 0.326101f
C130 minus.n58 a_n2102_n5888# 3.03924f
C131 drain_left.t4 a_n2102_n5888# 0.681242f
C132 drain_left.t17 a_n2102_n5888# 0.681242f
C133 drain_left.n0 a_n2102_n5888# 6.28229f
C134 drain_left.t5 a_n2102_n5888# 0.681242f
C135 drain_left.t15 a_n2102_n5888# 0.681242f
C136 drain_left.n1 a_n2102_n5888# 6.27838f
C137 drain_left.n2 a_n2102_n5888# 0.829823f
C138 drain_left.t7 a_n2102_n5888# 0.681242f
C139 drain_left.t16 a_n2102_n5888# 0.681242f
C140 drain_left.n3 a_n2102_n5888# 6.27838f
C141 drain_left.t11 a_n2102_n5888# 0.681242f
C142 drain_left.t1 a_n2102_n5888# 0.681242f
C143 drain_left.n4 a_n2102_n5888# 6.28229f
C144 drain_left.t9 a_n2102_n5888# 0.681242f
C145 drain_left.t0 a_n2102_n5888# 0.681242f
C146 drain_left.n5 a_n2102_n5888# 6.27838f
C147 drain_left.n6 a_n2102_n5888# 0.829823f
C148 drain_left.n7 a_n2102_n5888# 3.26633f
C149 drain_left.t18 a_n2102_n5888# 0.681242f
C150 drain_left.t13 a_n2102_n5888# 0.681242f
C151 drain_left.n8 a_n2102_n5888# 6.28229f
C152 drain_left.t8 a_n2102_n5888# 0.681242f
C153 drain_left.t2 a_n2102_n5888# 0.681242f
C154 drain_left.n9 a_n2102_n5888# 6.27839f
C155 drain_left.n10 a_n2102_n5888# 0.834331f
C156 drain_left.t14 a_n2102_n5888# 0.681242f
C157 drain_left.t10 a_n2102_n5888# 0.681242f
C158 drain_left.n11 a_n2102_n5888# 6.27839f
C159 drain_left.n12 a_n2102_n5888# 0.412173f
C160 drain_left.t3 a_n2102_n5888# 0.681242f
C161 drain_left.t19 a_n2102_n5888# 0.681242f
C162 drain_left.n13 a_n2102_n5888# 6.27839f
C163 drain_left.n14 a_n2102_n5888# 0.412173f
C164 drain_left.t12 a_n2102_n5888# 0.681242f
C165 drain_left.t6 a_n2102_n5888# 0.681242f
C166 drain_left.n15 a_n2102_n5888# 6.27837f
C167 drain_left.n16 a_n2102_n5888# 0.699214f
C168 source.n0 a_n2102_n5888# 0.039994f
C169 source.n1 a_n2102_n5888# 0.029011f
C170 source.n2 a_n2102_n5888# 0.015589f
C171 source.n3 a_n2102_n5888# 0.036847f
C172 source.n4 a_n2102_n5888# 0.016506f
C173 source.n5 a_n2102_n5888# 0.029011f
C174 source.n6 a_n2102_n5888# 0.015589f
C175 source.n7 a_n2102_n5888# 0.036847f
C176 source.n8 a_n2102_n5888# 0.016506f
C177 source.n9 a_n2102_n5888# 0.029011f
C178 source.n10 a_n2102_n5888# 0.015589f
C179 source.n11 a_n2102_n5888# 0.036847f
C180 source.n12 a_n2102_n5888# 0.016506f
C181 source.n13 a_n2102_n5888# 0.029011f
C182 source.n14 a_n2102_n5888# 0.015589f
C183 source.n15 a_n2102_n5888# 0.036847f
C184 source.n16 a_n2102_n5888# 0.036847f
C185 source.n17 a_n2102_n5888# 0.016506f
C186 source.n18 a_n2102_n5888# 0.029011f
C187 source.n19 a_n2102_n5888# 0.015589f
C188 source.n20 a_n2102_n5888# 0.036847f
C189 source.n21 a_n2102_n5888# 0.016506f
C190 source.n22 a_n2102_n5888# 0.029011f
C191 source.n23 a_n2102_n5888# 0.015589f
C192 source.n24 a_n2102_n5888# 0.036847f
C193 source.n25 a_n2102_n5888# 0.016506f
C194 source.n26 a_n2102_n5888# 0.029011f
C195 source.n27 a_n2102_n5888# 0.015589f
C196 source.n28 a_n2102_n5888# 0.036847f
C197 source.n29 a_n2102_n5888# 0.016506f
C198 source.n30 a_n2102_n5888# 0.029011f
C199 source.n31 a_n2102_n5888# 0.015589f
C200 source.n32 a_n2102_n5888# 0.036847f
C201 source.n33 a_n2102_n5888# 0.016506f
C202 source.n34 a_n2102_n5888# 0.029011f
C203 source.n35 a_n2102_n5888# 0.016048f
C204 source.n36 a_n2102_n5888# 0.036847f
C205 source.n37 a_n2102_n5888# 0.015589f
C206 source.n38 a_n2102_n5888# 0.016506f
C207 source.n39 a_n2102_n5888# 0.029011f
C208 source.n40 a_n2102_n5888# 0.015589f
C209 source.n41 a_n2102_n5888# 0.036847f
C210 source.n42 a_n2102_n5888# 0.016506f
C211 source.n43 a_n2102_n5888# 0.029011f
C212 source.n44 a_n2102_n5888# 0.015589f
C213 source.n45 a_n2102_n5888# 0.027635f
C214 source.n46 a_n2102_n5888# 0.026048f
C215 source.t37 a_n2102_n5888# 0.064263f
C216 source.n47 a_n2102_n5888# 0.353956f
C217 source.n48 a_n2102_n5888# 3.14101f
C218 source.n49 a_n2102_n5888# 0.015589f
C219 source.n50 a_n2102_n5888# 0.016506f
C220 source.n51 a_n2102_n5888# 0.036847f
C221 source.n52 a_n2102_n5888# 0.036847f
C222 source.n53 a_n2102_n5888# 0.016506f
C223 source.n54 a_n2102_n5888# 0.015589f
C224 source.n55 a_n2102_n5888# 0.029011f
C225 source.n56 a_n2102_n5888# 0.029011f
C226 source.n57 a_n2102_n5888# 0.015589f
C227 source.n58 a_n2102_n5888# 0.016506f
C228 source.n59 a_n2102_n5888# 0.036847f
C229 source.n60 a_n2102_n5888# 0.036847f
C230 source.n61 a_n2102_n5888# 0.016506f
C231 source.n62 a_n2102_n5888# 0.015589f
C232 source.n63 a_n2102_n5888# 0.029011f
C233 source.n64 a_n2102_n5888# 0.029011f
C234 source.n65 a_n2102_n5888# 0.015589f
C235 source.n66 a_n2102_n5888# 0.016506f
C236 source.n67 a_n2102_n5888# 0.036847f
C237 source.n68 a_n2102_n5888# 0.036847f
C238 source.n69 a_n2102_n5888# 0.036847f
C239 source.n70 a_n2102_n5888# 0.016048f
C240 source.n71 a_n2102_n5888# 0.015589f
C241 source.n72 a_n2102_n5888# 0.029011f
C242 source.n73 a_n2102_n5888# 0.029011f
C243 source.n74 a_n2102_n5888# 0.015589f
C244 source.n75 a_n2102_n5888# 0.016506f
C245 source.n76 a_n2102_n5888# 0.036847f
C246 source.n77 a_n2102_n5888# 0.036847f
C247 source.n78 a_n2102_n5888# 0.016506f
C248 source.n79 a_n2102_n5888# 0.015589f
C249 source.n80 a_n2102_n5888# 0.029011f
C250 source.n81 a_n2102_n5888# 0.029011f
C251 source.n82 a_n2102_n5888# 0.015589f
C252 source.n83 a_n2102_n5888# 0.016506f
C253 source.n84 a_n2102_n5888# 0.036847f
C254 source.n85 a_n2102_n5888# 0.036847f
C255 source.n86 a_n2102_n5888# 0.016506f
C256 source.n87 a_n2102_n5888# 0.015589f
C257 source.n88 a_n2102_n5888# 0.029011f
C258 source.n89 a_n2102_n5888# 0.029011f
C259 source.n90 a_n2102_n5888# 0.015589f
C260 source.n91 a_n2102_n5888# 0.016506f
C261 source.n92 a_n2102_n5888# 0.036847f
C262 source.n93 a_n2102_n5888# 0.036847f
C263 source.n94 a_n2102_n5888# 0.016506f
C264 source.n95 a_n2102_n5888# 0.015589f
C265 source.n96 a_n2102_n5888# 0.029011f
C266 source.n97 a_n2102_n5888# 0.029011f
C267 source.n98 a_n2102_n5888# 0.015589f
C268 source.n99 a_n2102_n5888# 0.016506f
C269 source.n100 a_n2102_n5888# 0.036847f
C270 source.n101 a_n2102_n5888# 0.036847f
C271 source.n102 a_n2102_n5888# 0.016506f
C272 source.n103 a_n2102_n5888# 0.015589f
C273 source.n104 a_n2102_n5888# 0.029011f
C274 source.n105 a_n2102_n5888# 0.029011f
C275 source.n106 a_n2102_n5888# 0.015589f
C276 source.n107 a_n2102_n5888# 0.016506f
C277 source.n108 a_n2102_n5888# 0.036847f
C278 source.n109 a_n2102_n5888# 0.036847f
C279 source.n110 a_n2102_n5888# 0.016506f
C280 source.n111 a_n2102_n5888# 0.015589f
C281 source.n112 a_n2102_n5888# 0.029011f
C282 source.n113 a_n2102_n5888# 0.029011f
C283 source.n114 a_n2102_n5888# 0.015589f
C284 source.n115 a_n2102_n5888# 0.016048f
C285 source.n116 a_n2102_n5888# 0.016048f
C286 source.n117 a_n2102_n5888# 0.036847f
C287 source.n118 a_n2102_n5888# 0.036847f
C288 source.n119 a_n2102_n5888# 0.016506f
C289 source.n120 a_n2102_n5888# 0.015589f
C290 source.n121 a_n2102_n5888# 0.029011f
C291 source.n122 a_n2102_n5888# 0.029011f
C292 source.n123 a_n2102_n5888# 0.015589f
C293 source.n124 a_n2102_n5888# 0.016506f
C294 source.n125 a_n2102_n5888# 0.036847f
C295 source.n126 a_n2102_n5888# 0.036847f
C296 source.n127 a_n2102_n5888# 0.016506f
C297 source.n128 a_n2102_n5888# 0.015589f
C298 source.n129 a_n2102_n5888# 0.029011f
C299 source.n130 a_n2102_n5888# 0.029011f
C300 source.n131 a_n2102_n5888# 0.015589f
C301 source.n132 a_n2102_n5888# 0.016506f
C302 source.n133 a_n2102_n5888# 0.036847f
C303 source.n134 a_n2102_n5888# 0.078383f
C304 source.n135 a_n2102_n5888# 0.016506f
C305 source.n136 a_n2102_n5888# 0.015589f
C306 source.n137 a_n2102_n5888# 0.063887f
C307 source.n138 a_n2102_n5888# 0.043617f
C308 source.n139 a_n2102_n5888# 2.28002f
C309 source.t31 a_n2102_n5888# 0.57313f
C310 source.t19 a_n2102_n5888# 0.57313f
C311 source.n140 a_n2102_n5888# 5.18691f
C312 source.n141 a_n2102_n5888# 0.402437f
C313 source.t18 a_n2102_n5888# 0.57313f
C314 source.t33 a_n2102_n5888# 0.57313f
C315 source.n142 a_n2102_n5888# 5.18691f
C316 source.n143 a_n2102_n5888# 0.402437f
C317 source.t34 a_n2102_n5888# 0.57313f
C318 source.t20 a_n2102_n5888# 0.57313f
C319 source.n144 a_n2102_n5888# 5.18691f
C320 source.n145 a_n2102_n5888# 0.402437f
C321 source.t28 a_n2102_n5888# 0.57313f
C322 source.t32 a_n2102_n5888# 0.57313f
C323 source.n146 a_n2102_n5888# 5.18691f
C324 source.n147 a_n2102_n5888# 0.402437f
C325 source.n148 a_n2102_n5888# 0.039994f
C326 source.n149 a_n2102_n5888# 0.029011f
C327 source.n150 a_n2102_n5888# 0.015589f
C328 source.n151 a_n2102_n5888# 0.036847f
C329 source.n152 a_n2102_n5888# 0.016506f
C330 source.n153 a_n2102_n5888# 0.029011f
C331 source.n154 a_n2102_n5888# 0.015589f
C332 source.n155 a_n2102_n5888# 0.036847f
C333 source.n156 a_n2102_n5888# 0.016506f
C334 source.n157 a_n2102_n5888# 0.029011f
C335 source.n158 a_n2102_n5888# 0.015589f
C336 source.n159 a_n2102_n5888# 0.036847f
C337 source.n160 a_n2102_n5888# 0.016506f
C338 source.n161 a_n2102_n5888# 0.029011f
C339 source.n162 a_n2102_n5888# 0.015589f
C340 source.n163 a_n2102_n5888# 0.036847f
C341 source.n164 a_n2102_n5888# 0.036847f
C342 source.n165 a_n2102_n5888# 0.016506f
C343 source.n166 a_n2102_n5888# 0.029011f
C344 source.n167 a_n2102_n5888# 0.015589f
C345 source.n168 a_n2102_n5888# 0.036847f
C346 source.n169 a_n2102_n5888# 0.016506f
C347 source.n170 a_n2102_n5888# 0.029011f
C348 source.n171 a_n2102_n5888# 0.015589f
C349 source.n172 a_n2102_n5888# 0.036847f
C350 source.n173 a_n2102_n5888# 0.016506f
C351 source.n174 a_n2102_n5888# 0.029011f
C352 source.n175 a_n2102_n5888# 0.015589f
C353 source.n176 a_n2102_n5888# 0.036847f
C354 source.n177 a_n2102_n5888# 0.016506f
C355 source.n178 a_n2102_n5888# 0.029011f
C356 source.n179 a_n2102_n5888# 0.015589f
C357 source.n180 a_n2102_n5888# 0.036847f
C358 source.n181 a_n2102_n5888# 0.016506f
C359 source.n182 a_n2102_n5888# 0.029011f
C360 source.n183 a_n2102_n5888# 0.016048f
C361 source.n184 a_n2102_n5888# 0.036847f
C362 source.n185 a_n2102_n5888# 0.015589f
C363 source.n186 a_n2102_n5888# 0.016506f
C364 source.n187 a_n2102_n5888# 0.029011f
C365 source.n188 a_n2102_n5888# 0.015589f
C366 source.n189 a_n2102_n5888# 0.036847f
C367 source.n190 a_n2102_n5888# 0.016506f
C368 source.n191 a_n2102_n5888# 0.029011f
C369 source.n192 a_n2102_n5888# 0.015589f
C370 source.n193 a_n2102_n5888# 0.027635f
C371 source.n194 a_n2102_n5888# 0.026048f
C372 source.t23 a_n2102_n5888# 0.064263f
C373 source.n195 a_n2102_n5888# 0.353956f
C374 source.n196 a_n2102_n5888# 3.14101f
C375 source.n197 a_n2102_n5888# 0.015589f
C376 source.n198 a_n2102_n5888# 0.016506f
C377 source.n199 a_n2102_n5888# 0.036847f
C378 source.n200 a_n2102_n5888# 0.036847f
C379 source.n201 a_n2102_n5888# 0.016506f
C380 source.n202 a_n2102_n5888# 0.015589f
C381 source.n203 a_n2102_n5888# 0.029011f
C382 source.n204 a_n2102_n5888# 0.029011f
C383 source.n205 a_n2102_n5888# 0.015589f
C384 source.n206 a_n2102_n5888# 0.016506f
C385 source.n207 a_n2102_n5888# 0.036847f
C386 source.n208 a_n2102_n5888# 0.036847f
C387 source.n209 a_n2102_n5888# 0.016506f
C388 source.n210 a_n2102_n5888# 0.015589f
C389 source.n211 a_n2102_n5888# 0.029011f
C390 source.n212 a_n2102_n5888# 0.029011f
C391 source.n213 a_n2102_n5888# 0.015589f
C392 source.n214 a_n2102_n5888# 0.016506f
C393 source.n215 a_n2102_n5888# 0.036847f
C394 source.n216 a_n2102_n5888# 0.036847f
C395 source.n217 a_n2102_n5888# 0.036847f
C396 source.n218 a_n2102_n5888# 0.016048f
C397 source.n219 a_n2102_n5888# 0.015589f
C398 source.n220 a_n2102_n5888# 0.029011f
C399 source.n221 a_n2102_n5888# 0.029011f
C400 source.n222 a_n2102_n5888# 0.015589f
C401 source.n223 a_n2102_n5888# 0.016506f
C402 source.n224 a_n2102_n5888# 0.036847f
C403 source.n225 a_n2102_n5888# 0.036847f
C404 source.n226 a_n2102_n5888# 0.016506f
C405 source.n227 a_n2102_n5888# 0.015589f
C406 source.n228 a_n2102_n5888# 0.029011f
C407 source.n229 a_n2102_n5888# 0.029011f
C408 source.n230 a_n2102_n5888# 0.015589f
C409 source.n231 a_n2102_n5888# 0.016506f
C410 source.n232 a_n2102_n5888# 0.036847f
C411 source.n233 a_n2102_n5888# 0.036847f
C412 source.n234 a_n2102_n5888# 0.016506f
C413 source.n235 a_n2102_n5888# 0.015589f
C414 source.n236 a_n2102_n5888# 0.029011f
C415 source.n237 a_n2102_n5888# 0.029011f
C416 source.n238 a_n2102_n5888# 0.015589f
C417 source.n239 a_n2102_n5888# 0.016506f
C418 source.n240 a_n2102_n5888# 0.036847f
C419 source.n241 a_n2102_n5888# 0.036847f
C420 source.n242 a_n2102_n5888# 0.016506f
C421 source.n243 a_n2102_n5888# 0.015589f
C422 source.n244 a_n2102_n5888# 0.029011f
C423 source.n245 a_n2102_n5888# 0.029011f
C424 source.n246 a_n2102_n5888# 0.015589f
C425 source.n247 a_n2102_n5888# 0.016506f
C426 source.n248 a_n2102_n5888# 0.036847f
C427 source.n249 a_n2102_n5888# 0.036847f
C428 source.n250 a_n2102_n5888# 0.016506f
C429 source.n251 a_n2102_n5888# 0.015589f
C430 source.n252 a_n2102_n5888# 0.029011f
C431 source.n253 a_n2102_n5888# 0.029011f
C432 source.n254 a_n2102_n5888# 0.015589f
C433 source.n255 a_n2102_n5888# 0.016506f
C434 source.n256 a_n2102_n5888# 0.036847f
C435 source.n257 a_n2102_n5888# 0.036847f
C436 source.n258 a_n2102_n5888# 0.016506f
C437 source.n259 a_n2102_n5888# 0.015589f
C438 source.n260 a_n2102_n5888# 0.029011f
C439 source.n261 a_n2102_n5888# 0.029011f
C440 source.n262 a_n2102_n5888# 0.015589f
C441 source.n263 a_n2102_n5888# 0.016048f
C442 source.n264 a_n2102_n5888# 0.016048f
C443 source.n265 a_n2102_n5888# 0.036847f
C444 source.n266 a_n2102_n5888# 0.036847f
C445 source.n267 a_n2102_n5888# 0.016506f
C446 source.n268 a_n2102_n5888# 0.015589f
C447 source.n269 a_n2102_n5888# 0.029011f
C448 source.n270 a_n2102_n5888# 0.029011f
C449 source.n271 a_n2102_n5888# 0.015589f
C450 source.n272 a_n2102_n5888# 0.016506f
C451 source.n273 a_n2102_n5888# 0.036847f
C452 source.n274 a_n2102_n5888# 0.036847f
C453 source.n275 a_n2102_n5888# 0.016506f
C454 source.n276 a_n2102_n5888# 0.015589f
C455 source.n277 a_n2102_n5888# 0.029011f
C456 source.n278 a_n2102_n5888# 0.029011f
C457 source.n279 a_n2102_n5888# 0.015589f
C458 source.n280 a_n2102_n5888# 0.016506f
C459 source.n281 a_n2102_n5888# 0.036847f
C460 source.n282 a_n2102_n5888# 0.078383f
C461 source.n283 a_n2102_n5888# 0.016506f
C462 source.n284 a_n2102_n5888# 0.015589f
C463 source.n285 a_n2102_n5888# 0.063887f
C464 source.n286 a_n2102_n5888# 0.043617f
C465 source.n287 a_n2102_n5888# 0.117678f
C466 source.n288 a_n2102_n5888# 0.039994f
C467 source.n289 a_n2102_n5888# 0.029011f
C468 source.n290 a_n2102_n5888# 0.015589f
C469 source.n291 a_n2102_n5888# 0.036847f
C470 source.n292 a_n2102_n5888# 0.016506f
C471 source.n293 a_n2102_n5888# 0.029011f
C472 source.n294 a_n2102_n5888# 0.015589f
C473 source.n295 a_n2102_n5888# 0.036847f
C474 source.n296 a_n2102_n5888# 0.016506f
C475 source.n297 a_n2102_n5888# 0.029011f
C476 source.n298 a_n2102_n5888# 0.015589f
C477 source.n299 a_n2102_n5888# 0.036847f
C478 source.n300 a_n2102_n5888# 0.016506f
C479 source.n301 a_n2102_n5888# 0.029011f
C480 source.n302 a_n2102_n5888# 0.015589f
C481 source.n303 a_n2102_n5888# 0.036847f
C482 source.n304 a_n2102_n5888# 0.036847f
C483 source.n305 a_n2102_n5888# 0.016506f
C484 source.n306 a_n2102_n5888# 0.029011f
C485 source.n307 a_n2102_n5888# 0.015589f
C486 source.n308 a_n2102_n5888# 0.036847f
C487 source.n309 a_n2102_n5888# 0.016506f
C488 source.n310 a_n2102_n5888# 0.029011f
C489 source.n311 a_n2102_n5888# 0.015589f
C490 source.n312 a_n2102_n5888# 0.036847f
C491 source.n313 a_n2102_n5888# 0.016506f
C492 source.n314 a_n2102_n5888# 0.029011f
C493 source.n315 a_n2102_n5888# 0.015589f
C494 source.n316 a_n2102_n5888# 0.036847f
C495 source.n317 a_n2102_n5888# 0.016506f
C496 source.n318 a_n2102_n5888# 0.029011f
C497 source.n319 a_n2102_n5888# 0.015589f
C498 source.n320 a_n2102_n5888# 0.036847f
C499 source.n321 a_n2102_n5888# 0.016506f
C500 source.n322 a_n2102_n5888# 0.029011f
C501 source.n323 a_n2102_n5888# 0.016048f
C502 source.n324 a_n2102_n5888# 0.036847f
C503 source.n325 a_n2102_n5888# 0.015589f
C504 source.n326 a_n2102_n5888# 0.016506f
C505 source.n327 a_n2102_n5888# 0.029011f
C506 source.n328 a_n2102_n5888# 0.015589f
C507 source.n329 a_n2102_n5888# 0.036847f
C508 source.n330 a_n2102_n5888# 0.016506f
C509 source.n331 a_n2102_n5888# 0.029011f
C510 source.n332 a_n2102_n5888# 0.015589f
C511 source.n333 a_n2102_n5888# 0.027635f
C512 source.n334 a_n2102_n5888# 0.026048f
C513 source.t2 a_n2102_n5888# 0.064263f
C514 source.n335 a_n2102_n5888# 0.353956f
C515 source.n336 a_n2102_n5888# 3.14101f
C516 source.n337 a_n2102_n5888# 0.015589f
C517 source.n338 a_n2102_n5888# 0.016506f
C518 source.n339 a_n2102_n5888# 0.036847f
C519 source.n340 a_n2102_n5888# 0.036847f
C520 source.n341 a_n2102_n5888# 0.016506f
C521 source.n342 a_n2102_n5888# 0.015589f
C522 source.n343 a_n2102_n5888# 0.029011f
C523 source.n344 a_n2102_n5888# 0.029011f
C524 source.n345 a_n2102_n5888# 0.015589f
C525 source.n346 a_n2102_n5888# 0.016506f
C526 source.n347 a_n2102_n5888# 0.036847f
C527 source.n348 a_n2102_n5888# 0.036847f
C528 source.n349 a_n2102_n5888# 0.016506f
C529 source.n350 a_n2102_n5888# 0.015589f
C530 source.n351 a_n2102_n5888# 0.029011f
C531 source.n352 a_n2102_n5888# 0.029011f
C532 source.n353 a_n2102_n5888# 0.015589f
C533 source.n354 a_n2102_n5888# 0.016506f
C534 source.n355 a_n2102_n5888# 0.036847f
C535 source.n356 a_n2102_n5888# 0.036847f
C536 source.n357 a_n2102_n5888# 0.036847f
C537 source.n358 a_n2102_n5888# 0.016048f
C538 source.n359 a_n2102_n5888# 0.015589f
C539 source.n360 a_n2102_n5888# 0.029011f
C540 source.n361 a_n2102_n5888# 0.029011f
C541 source.n362 a_n2102_n5888# 0.015589f
C542 source.n363 a_n2102_n5888# 0.016506f
C543 source.n364 a_n2102_n5888# 0.036847f
C544 source.n365 a_n2102_n5888# 0.036847f
C545 source.n366 a_n2102_n5888# 0.016506f
C546 source.n367 a_n2102_n5888# 0.015589f
C547 source.n368 a_n2102_n5888# 0.029011f
C548 source.n369 a_n2102_n5888# 0.029011f
C549 source.n370 a_n2102_n5888# 0.015589f
C550 source.n371 a_n2102_n5888# 0.016506f
C551 source.n372 a_n2102_n5888# 0.036847f
C552 source.n373 a_n2102_n5888# 0.036847f
C553 source.n374 a_n2102_n5888# 0.016506f
C554 source.n375 a_n2102_n5888# 0.015589f
C555 source.n376 a_n2102_n5888# 0.029011f
C556 source.n377 a_n2102_n5888# 0.029011f
C557 source.n378 a_n2102_n5888# 0.015589f
C558 source.n379 a_n2102_n5888# 0.016506f
C559 source.n380 a_n2102_n5888# 0.036847f
C560 source.n381 a_n2102_n5888# 0.036847f
C561 source.n382 a_n2102_n5888# 0.016506f
C562 source.n383 a_n2102_n5888# 0.015589f
C563 source.n384 a_n2102_n5888# 0.029011f
C564 source.n385 a_n2102_n5888# 0.029011f
C565 source.n386 a_n2102_n5888# 0.015589f
C566 source.n387 a_n2102_n5888# 0.016506f
C567 source.n388 a_n2102_n5888# 0.036847f
C568 source.n389 a_n2102_n5888# 0.036847f
C569 source.n390 a_n2102_n5888# 0.016506f
C570 source.n391 a_n2102_n5888# 0.015589f
C571 source.n392 a_n2102_n5888# 0.029011f
C572 source.n393 a_n2102_n5888# 0.029011f
C573 source.n394 a_n2102_n5888# 0.015589f
C574 source.n395 a_n2102_n5888# 0.016506f
C575 source.n396 a_n2102_n5888# 0.036847f
C576 source.n397 a_n2102_n5888# 0.036847f
C577 source.n398 a_n2102_n5888# 0.016506f
C578 source.n399 a_n2102_n5888# 0.015589f
C579 source.n400 a_n2102_n5888# 0.029011f
C580 source.n401 a_n2102_n5888# 0.029011f
C581 source.n402 a_n2102_n5888# 0.015589f
C582 source.n403 a_n2102_n5888# 0.016048f
C583 source.n404 a_n2102_n5888# 0.016048f
C584 source.n405 a_n2102_n5888# 0.036847f
C585 source.n406 a_n2102_n5888# 0.036847f
C586 source.n407 a_n2102_n5888# 0.016506f
C587 source.n408 a_n2102_n5888# 0.015589f
C588 source.n409 a_n2102_n5888# 0.029011f
C589 source.n410 a_n2102_n5888# 0.029011f
C590 source.n411 a_n2102_n5888# 0.015589f
C591 source.n412 a_n2102_n5888# 0.016506f
C592 source.n413 a_n2102_n5888# 0.036847f
C593 source.n414 a_n2102_n5888# 0.036847f
C594 source.n415 a_n2102_n5888# 0.016506f
C595 source.n416 a_n2102_n5888# 0.015589f
C596 source.n417 a_n2102_n5888# 0.029011f
C597 source.n418 a_n2102_n5888# 0.029011f
C598 source.n419 a_n2102_n5888# 0.015589f
C599 source.n420 a_n2102_n5888# 0.016506f
C600 source.n421 a_n2102_n5888# 0.036847f
C601 source.n422 a_n2102_n5888# 0.078383f
C602 source.n423 a_n2102_n5888# 0.016506f
C603 source.n424 a_n2102_n5888# 0.015589f
C604 source.n425 a_n2102_n5888# 0.063887f
C605 source.n426 a_n2102_n5888# 0.043617f
C606 source.n427 a_n2102_n5888# 0.117678f
C607 source.t1 a_n2102_n5888# 0.57313f
C608 source.t5 a_n2102_n5888# 0.57313f
C609 source.n428 a_n2102_n5888# 5.18691f
C610 source.n429 a_n2102_n5888# 0.402437f
C611 source.t12 a_n2102_n5888# 0.57313f
C612 source.t0 a_n2102_n5888# 0.57313f
C613 source.n430 a_n2102_n5888# 5.18691f
C614 source.n431 a_n2102_n5888# 0.402437f
C615 source.t9 a_n2102_n5888# 0.57313f
C616 source.t8 a_n2102_n5888# 0.57313f
C617 source.n432 a_n2102_n5888# 5.18691f
C618 source.n433 a_n2102_n5888# 0.402437f
C619 source.t4 a_n2102_n5888# 0.57313f
C620 source.t7 a_n2102_n5888# 0.57313f
C621 source.n434 a_n2102_n5888# 5.18691f
C622 source.n435 a_n2102_n5888# 0.402437f
C623 source.n436 a_n2102_n5888# 0.039994f
C624 source.n437 a_n2102_n5888# 0.029011f
C625 source.n438 a_n2102_n5888# 0.015589f
C626 source.n439 a_n2102_n5888# 0.036847f
C627 source.n440 a_n2102_n5888# 0.016506f
C628 source.n441 a_n2102_n5888# 0.029011f
C629 source.n442 a_n2102_n5888# 0.015589f
C630 source.n443 a_n2102_n5888# 0.036847f
C631 source.n444 a_n2102_n5888# 0.016506f
C632 source.n445 a_n2102_n5888# 0.029011f
C633 source.n446 a_n2102_n5888# 0.015589f
C634 source.n447 a_n2102_n5888# 0.036847f
C635 source.n448 a_n2102_n5888# 0.016506f
C636 source.n449 a_n2102_n5888# 0.029011f
C637 source.n450 a_n2102_n5888# 0.015589f
C638 source.n451 a_n2102_n5888# 0.036847f
C639 source.n452 a_n2102_n5888# 0.036847f
C640 source.n453 a_n2102_n5888# 0.016506f
C641 source.n454 a_n2102_n5888# 0.029011f
C642 source.n455 a_n2102_n5888# 0.015589f
C643 source.n456 a_n2102_n5888# 0.036847f
C644 source.n457 a_n2102_n5888# 0.016506f
C645 source.n458 a_n2102_n5888# 0.029011f
C646 source.n459 a_n2102_n5888# 0.015589f
C647 source.n460 a_n2102_n5888# 0.036847f
C648 source.n461 a_n2102_n5888# 0.016506f
C649 source.n462 a_n2102_n5888# 0.029011f
C650 source.n463 a_n2102_n5888# 0.015589f
C651 source.n464 a_n2102_n5888# 0.036847f
C652 source.n465 a_n2102_n5888# 0.016506f
C653 source.n466 a_n2102_n5888# 0.029011f
C654 source.n467 a_n2102_n5888# 0.015589f
C655 source.n468 a_n2102_n5888# 0.036847f
C656 source.n469 a_n2102_n5888# 0.016506f
C657 source.n470 a_n2102_n5888# 0.029011f
C658 source.n471 a_n2102_n5888# 0.016048f
C659 source.n472 a_n2102_n5888# 0.036847f
C660 source.n473 a_n2102_n5888# 0.015589f
C661 source.n474 a_n2102_n5888# 0.016506f
C662 source.n475 a_n2102_n5888# 0.029011f
C663 source.n476 a_n2102_n5888# 0.015589f
C664 source.n477 a_n2102_n5888# 0.036847f
C665 source.n478 a_n2102_n5888# 0.016506f
C666 source.n479 a_n2102_n5888# 0.029011f
C667 source.n480 a_n2102_n5888# 0.015589f
C668 source.n481 a_n2102_n5888# 0.027635f
C669 source.n482 a_n2102_n5888# 0.026048f
C670 source.t38 a_n2102_n5888# 0.064263f
C671 source.n483 a_n2102_n5888# 0.353956f
C672 source.n484 a_n2102_n5888# 3.14101f
C673 source.n485 a_n2102_n5888# 0.015589f
C674 source.n486 a_n2102_n5888# 0.016506f
C675 source.n487 a_n2102_n5888# 0.036847f
C676 source.n488 a_n2102_n5888# 0.036847f
C677 source.n489 a_n2102_n5888# 0.016506f
C678 source.n490 a_n2102_n5888# 0.015589f
C679 source.n491 a_n2102_n5888# 0.029011f
C680 source.n492 a_n2102_n5888# 0.029011f
C681 source.n493 a_n2102_n5888# 0.015589f
C682 source.n494 a_n2102_n5888# 0.016506f
C683 source.n495 a_n2102_n5888# 0.036847f
C684 source.n496 a_n2102_n5888# 0.036847f
C685 source.n497 a_n2102_n5888# 0.016506f
C686 source.n498 a_n2102_n5888# 0.015589f
C687 source.n499 a_n2102_n5888# 0.029011f
C688 source.n500 a_n2102_n5888# 0.029011f
C689 source.n501 a_n2102_n5888# 0.015589f
C690 source.n502 a_n2102_n5888# 0.016506f
C691 source.n503 a_n2102_n5888# 0.036847f
C692 source.n504 a_n2102_n5888# 0.036847f
C693 source.n505 a_n2102_n5888# 0.036847f
C694 source.n506 a_n2102_n5888# 0.016048f
C695 source.n507 a_n2102_n5888# 0.015589f
C696 source.n508 a_n2102_n5888# 0.029011f
C697 source.n509 a_n2102_n5888# 0.029011f
C698 source.n510 a_n2102_n5888# 0.015589f
C699 source.n511 a_n2102_n5888# 0.016506f
C700 source.n512 a_n2102_n5888# 0.036847f
C701 source.n513 a_n2102_n5888# 0.036847f
C702 source.n514 a_n2102_n5888# 0.016506f
C703 source.n515 a_n2102_n5888# 0.015589f
C704 source.n516 a_n2102_n5888# 0.029011f
C705 source.n517 a_n2102_n5888# 0.029011f
C706 source.n518 a_n2102_n5888# 0.015589f
C707 source.n519 a_n2102_n5888# 0.016506f
C708 source.n520 a_n2102_n5888# 0.036847f
C709 source.n521 a_n2102_n5888# 0.036847f
C710 source.n522 a_n2102_n5888# 0.016506f
C711 source.n523 a_n2102_n5888# 0.015589f
C712 source.n524 a_n2102_n5888# 0.029011f
C713 source.n525 a_n2102_n5888# 0.029011f
C714 source.n526 a_n2102_n5888# 0.015589f
C715 source.n527 a_n2102_n5888# 0.016506f
C716 source.n528 a_n2102_n5888# 0.036847f
C717 source.n529 a_n2102_n5888# 0.036847f
C718 source.n530 a_n2102_n5888# 0.016506f
C719 source.n531 a_n2102_n5888# 0.015589f
C720 source.n532 a_n2102_n5888# 0.029011f
C721 source.n533 a_n2102_n5888# 0.029011f
C722 source.n534 a_n2102_n5888# 0.015589f
C723 source.n535 a_n2102_n5888# 0.016506f
C724 source.n536 a_n2102_n5888# 0.036847f
C725 source.n537 a_n2102_n5888# 0.036847f
C726 source.n538 a_n2102_n5888# 0.016506f
C727 source.n539 a_n2102_n5888# 0.015589f
C728 source.n540 a_n2102_n5888# 0.029011f
C729 source.n541 a_n2102_n5888# 0.029011f
C730 source.n542 a_n2102_n5888# 0.015589f
C731 source.n543 a_n2102_n5888# 0.016506f
C732 source.n544 a_n2102_n5888# 0.036847f
C733 source.n545 a_n2102_n5888# 0.036847f
C734 source.n546 a_n2102_n5888# 0.016506f
C735 source.n547 a_n2102_n5888# 0.015589f
C736 source.n548 a_n2102_n5888# 0.029011f
C737 source.n549 a_n2102_n5888# 0.029011f
C738 source.n550 a_n2102_n5888# 0.015589f
C739 source.n551 a_n2102_n5888# 0.016048f
C740 source.n552 a_n2102_n5888# 0.016048f
C741 source.n553 a_n2102_n5888# 0.036847f
C742 source.n554 a_n2102_n5888# 0.036847f
C743 source.n555 a_n2102_n5888# 0.016506f
C744 source.n556 a_n2102_n5888# 0.015589f
C745 source.n557 a_n2102_n5888# 0.029011f
C746 source.n558 a_n2102_n5888# 0.029011f
C747 source.n559 a_n2102_n5888# 0.015589f
C748 source.n560 a_n2102_n5888# 0.016506f
C749 source.n561 a_n2102_n5888# 0.036847f
C750 source.n562 a_n2102_n5888# 0.036847f
C751 source.n563 a_n2102_n5888# 0.016506f
C752 source.n564 a_n2102_n5888# 0.015589f
C753 source.n565 a_n2102_n5888# 0.029011f
C754 source.n566 a_n2102_n5888# 0.029011f
C755 source.n567 a_n2102_n5888# 0.015589f
C756 source.n568 a_n2102_n5888# 0.016506f
C757 source.n569 a_n2102_n5888# 0.036847f
C758 source.n570 a_n2102_n5888# 0.078383f
C759 source.n571 a_n2102_n5888# 0.016506f
C760 source.n572 a_n2102_n5888# 0.015589f
C761 source.n573 a_n2102_n5888# 0.063887f
C762 source.n574 a_n2102_n5888# 0.043617f
C763 source.n575 a_n2102_n5888# 2.81671f
C764 source.n576 a_n2102_n5888# 0.039994f
C765 source.n577 a_n2102_n5888# 0.029011f
C766 source.n578 a_n2102_n5888# 0.015589f
C767 source.n579 a_n2102_n5888# 0.036847f
C768 source.n580 a_n2102_n5888# 0.016506f
C769 source.n581 a_n2102_n5888# 0.029011f
C770 source.n582 a_n2102_n5888# 0.015589f
C771 source.n583 a_n2102_n5888# 0.036847f
C772 source.n584 a_n2102_n5888# 0.016506f
C773 source.n585 a_n2102_n5888# 0.029011f
C774 source.n586 a_n2102_n5888# 0.015589f
C775 source.n587 a_n2102_n5888# 0.036847f
C776 source.n588 a_n2102_n5888# 0.016506f
C777 source.n589 a_n2102_n5888# 0.029011f
C778 source.n590 a_n2102_n5888# 0.015589f
C779 source.n591 a_n2102_n5888# 0.036847f
C780 source.n592 a_n2102_n5888# 0.016506f
C781 source.n593 a_n2102_n5888# 0.029011f
C782 source.n594 a_n2102_n5888# 0.015589f
C783 source.n595 a_n2102_n5888# 0.036847f
C784 source.n596 a_n2102_n5888# 0.016506f
C785 source.n597 a_n2102_n5888# 0.029011f
C786 source.n598 a_n2102_n5888# 0.015589f
C787 source.n599 a_n2102_n5888# 0.036847f
C788 source.n600 a_n2102_n5888# 0.016506f
C789 source.n601 a_n2102_n5888# 0.029011f
C790 source.n602 a_n2102_n5888# 0.015589f
C791 source.n603 a_n2102_n5888# 0.036847f
C792 source.n604 a_n2102_n5888# 0.016506f
C793 source.n605 a_n2102_n5888# 0.029011f
C794 source.n606 a_n2102_n5888# 0.015589f
C795 source.n607 a_n2102_n5888# 0.036847f
C796 source.n608 a_n2102_n5888# 0.016506f
C797 source.n609 a_n2102_n5888# 0.029011f
C798 source.n610 a_n2102_n5888# 0.016048f
C799 source.n611 a_n2102_n5888# 0.036847f
C800 source.n612 a_n2102_n5888# 0.016506f
C801 source.n613 a_n2102_n5888# 0.029011f
C802 source.n614 a_n2102_n5888# 0.015589f
C803 source.n615 a_n2102_n5888# 0.036847f
C804 source.n616 a_n2102_n5888# 0.016506f
C805 source.n617 a_n2102_n5888# 0.029011f
C806 source.n618 a_n2102_n5888# 0.015589f
C807 source.n619 a_n2102_n5888# 0.027635f
C808 source.n620 a_n2102_n5888# 0.026048f
C809 source.t26 a_n2102_n5888# 0.064264f
C810 source.n621 a_n2102_n5888# 0.353956f
C811 source.n622 a_n2102_n5888# 3.14101f
C812 source.n623 a_n2102_n5888# 0.015589f
C813 source.n624 a_n2102_n5888# 0.016506f
C814 source.n625 a_n2102_n5888# 0.036847f
C815 source.n626 a_n2102_n5888# 0.036847f
C816 source.n627 a_n2102_n5888# 0.016506f
C817 source.n628 a_n2102_n5888# 0.015589f
C818 source.n629 a_n2102_n5888# 0.029011f
C819 source.n630 a_n2102_n5888# 0.029011f
C820 source.n631 a_n2102_n5888# 0.015589f
C821 source.n632 a_n2102_n5888# 0.016506f
C822 source.n633 a_n2102_n5888# 0.036847f
C823 source.n634 a_n2102_n5888# 0.036847f
C824 source.n635 a_n2102_n5888# 0.016506f
C825 source.n636 a_n2102_n5888# 0.015589f
C826 source.n637 a_n2102_n5888# 0.029011f
C827 source.n638 a_n2102_n5888# 0.029011f
C828 source.n639 a_n2102_n5888# 0.015589f
C829 source.n640 a_n2102_n5888# 0.015589f
C830 source.n641 a_n2102_n5888# 0.016506f
C831 source.n642 a_n2102_n5888# 0.036847f
C832 source.n643 a_n2102_n5888# 0.036847f
C833 source.n644 a_n2102_n5888# 0.036847f
C834 source.n645 a_n2102_n5888# 0.016048f
C835 source.n646 a_n2102_n5888# 0.015589f
C836 source.n647 a_n2102_n5888# 0.029011f
C837 source.n648 a_n2102_n5888# 0.029011f
C838 source.n649 a_n2102_n5888# 0.015589f
C839 source.n650 a_n2102_n5888# 0.016506f
C840 source.n651 a_n2102_n5888# 0.036847f
C841 source.n652 a_n2102_n5888# 0.036847f
C842 source.n653 a_n2102_n5888# 0.016506f
C843 source.n654 a_n2102_n5888# 0.015589f
C844 source.n655 a_n2102_n5888# 0.029011f
C845 source.n656 a_n2102_n5888# 0.029011f
C846 source.n657 a_n2102_n5888# 0.015589f
C847 source.n658 a_n2102_n5888# 0.016506f
C848 source.n659 a_n2102_n5888# 0.036847f
C849 source.n660 a_n2102_n5888# 0.036847f
C850 source.n661 a_n2102_n5888# 0.016506f
C851 source.n662 a_n2102_n5888# 0.015589f
C852 source.n663 a_n2102_n5888# 0.029011f
C853 source.n664 a_n2102_n5888# 0.029011f
C854 source.n665 a_n2102_n5888# 0.015589f
C855 source.n666 a_n2102_n5888# 0.016506f
C856 source.n667 a_n2102_n5888# 0.036847f
C857 source.n668 a_n2102_n5888# 0.036847f
C858 source.n669 a_n2102_n5888# 0.016506f
C859 source.n670 a_n2102_n5888# 0.015589f
C860 source.n671 a_n2102_n5888# 0.029011f
C861 source.n672 a_n2102_n5888# 0.029011f
C862 source.n673 a_n2102_n5888# 0.015589f
C863 source.n674 a_n2102_n5888# 0.016506f
C864 source.n675 a_n2102_n5888# 0.036847f
C865 source.n676 a_n2102_n5888# 0.036847f
C866 source.n677 a_n2102_n5888# 0.016506f
C867 source.n678 a_n2102_n5888# 0.015589f
C868 source.n679 a_n2102_n5888# 0.029011f
C869 source.n680 a_n2102_n5888# 0.029011f
C870 source.n681 a_n2102_n5888# 0.015589f
C871 source.n682 a_n2102_n5888# 0.016506f
C872 source.n683 a_n2102_n5888# 0.036847f
C873 source.n684 a_n2102_n5888# 0.036847f
C874 source.n685 a_n2102_n5888# 0.036847f
C875 source.n686 a_n2102_n5888# 0.016506f
C876 source.n687 a_n2102_n5888# 0.015589f
C877 source.n688 a_n2102_n5888# 0.029011f
C878 source.n689 a_n2102_n5888# 0.029011f
C879 source.n690 a_n2102_n5888# 0.015589f
C880 source.n691 a_n2102_n5888# 0.016048f
C881 source.n692 a_n2102_n5888# 0.016048f
C882 source.n693 a_n2102_n5888# 0.036847f
C883 source.n694 a_n2102_n5888# 0.036847f
C884 source.n695 a_n2102_n5888# 0.016506f
C885 source.n696 a_n2102_n5888# 0.015589f
C886 source.n697 a_n2102_n5888# 0.029011f
C887 source.n698 a_n2102_n5888# 0.029011f
C888 source.n699 a_n2102_n5888# 0.015589f
C889 source.n700 a_n2102_n5888# 0.016506f
C890 source.n701 a_n2102_n5888# 0.036847f
C891 source.n702 a_n2102_n5888# 0.036847f
C892 source.n703 a_n2102_n5888# 0.016506f
C893 source.n704 a_n2102_n5888# 0.015589f
C894 source.n705 a_n2102_n5888# 0.029011f
C895 source.n706 a_n2102_n5888# 0.029011f
C896 source.n707 a_n2102_n5888# 0.015589f
C897 source.n708 a_n2102_n5888# 0.016506f
C898 source.n709 a_n2102_n5888# 0.036847f
C899 source.n710 a_n2102_n5888# 0.078383f
C900 source.n711 a_n2102_n5888# 0.016506f
C901 source.n712 a_n2102_n5888# 0.015589f
C902 source.n713 a_n2102_n5888# 0.063887f
C903 source.n714 a_n2102_n5888# 0.043617f
C904 source.n715 a_n2102_n5888# 2.81671f
C905 source.t30 a_n2102_n5888# 0.57313f
C906 source.t29 a_n2102_n5888# 0.57313f
C907 source.n716 a_n2102_n5888# 5.18691f
C908 source.n717 a_n2102_n5888# 0.402439f
C909 source.t21 a_n2102_n5888# 0.57313f
C910 source.t25 a_n2102_n5888# 0.57313f
C911 source.n718 a_n2102_n5888# 5.18691f
C912 source.n719 a_n2102_n5888# 0.402439f
C913 source.t22 a_n2102_n5888# 0.57313f
C914 source.t27 a_n2102_n5888# 0.57313f
C915 source.n720 a_n2102_n5888# 5.18691f
C916 source.n721 a_n2102_n5888# 0.402439f
C917 source.t36 a_n2102_n5888# 0.57313f
C918 source.t24 a_n2102_n5888# 0.57313f
C919 source.n722 a_n2102_n5888# 5.18691f
C920 source.n723 a_n2102_n5888# 0.402439f
C921 source.n724 a_n2102_n5888# 0.039994f
C922 source.n725 a_n2102_n5888# 0.029011f
C923 source.n726 a_n2102_n5888# 0.015589f
C924 source.n727 a_n2102_n5888# 0.036847f
C925 source.n728 a_n2102_n5888# 0.016506f
C926 source.n729 a_n2102_n5888# 0.029011f
C927 source.n730 a_n2102_n5888# 0.015589f
C928 source.n731 a_n2102_n5888# 0.036847f
C929 source.n732 a_n2102_n5888# 0.016506f
C930 source.n733 a_n2102_n5888# 0.029011f
C931 source.n734 a_n2102_n5888# 0.015589f
C932 source.n735 a_n2102_n5888# 0.036847f
C933 source.n736 a_n2102_n5888# 0.016506f
C934 source.n737 a_n2102_n5888# 0.029011f
C935 source.n738 a_n2102_n5888# 0.015589f
C936 source.n739 a_n2102_n5888# 0.036847f
C937 source.n740 a_n2102_n5888# 0.016506f
C938 source.n741 a_n2102_n5888# 0.029011f
C939 source.n742 a_n2102_n5888# 0.015589f
C940 source.n743 a_n2102_n5888# 0.036847f
C941 source.n744 a_n2102_n5888# 0.016506f
C942 source.n745 a_n2102_n5888# 0.029011f
C943 source.n746 a_n2102_n5888# 0.015589f
C944 source.n747 a_n2102_n5888# 0.036847f
C945 source.n748 a_n2102_n5888# 0.016506f
C946 source.n749 a_n2102_n5888# 0.029011f
C947 source.n750 a_n2102_n5888# 0.015589f
C948 source.n751 a_n2102_n5888# 0.036847f
C949 source.n752 a_n2102_n5888# 0.016506f
C950 source.n753 a_n2102_n5888# 0.029011f
C951 source.n754 a_n2102_n5888# 0.015589f
C952 source.n755 a_n2102_n5888# 0.036847f
C953 source.n756 a_n2102_n5888# 0.016506f
C954 source.n757 a_n2102_n5888# 0.029011f
C955 source.n758 a_n2102_n5888# 0.016048f
C956 source.n759 a_n2102_n5888# 0.036847f
C957 source.n760 a_n2102_n5888# 0.016506f
C958 source.n761 a_n2102_n5888# 0.029011f
C959 source.n762 a_n2102_n5888# 0.015589f
C960 source.n763 a_n2102_n5888# 0.036847f
C961 source.n764 a_n2102_n5888# 0.016506f
C962 source.n765 a_n2102_n5888# 0.029011f
C963 source.n766 a_n2102_n5888# 0.015589f
C964 source.n767 a_n2102_n5888# 0.027635f
C965 source.n768 a_n2102_n5888# 0.026048f
C966 source.t35 a_n2102_n5888# 0.064264f
C967 source.n769 a_n2102_n5888# 0.353956f
C968 source.n770 a_n2102_n5888# 3.14101f
C969 source.n771 a_n2102_n5888# 0.015589f
C970 source.n772 a_n2102_n5888# 0.016506f
C971 source.n773 a_n2102_n5888# 0.036847f
C972 source.n774 a_n2102_n5888# 0.036847f
C973 source.n775 a_n2102_n5888# 0.016506f
C974 source.n776 a_n2102_n5888# 0.015589f
C975 source.n777 a_n2102_n5888# 0.029011f
C976 source.n778 a_n2102_n5888# 0.029011f
C977 source.n779 a_n2102_n5888# 0.015589f
C978 source.n780 a_n2102_n5888# 0.016506f
C979 source.n781 a_n2102_n5888# 0.036847f
C980 source.n782 a_n2102_n5888# 0.036847f
C981 source.n783 a_n2102_n5888# 0.016506f
C982 source.n784 a_n2102_n5888# 0.015589f
C983 source.n785 a_n2102_n5888# 0.029011f
C984 source.n786 a_n2102_n5888# 0.029011f
C985 source.n787 a_n2102_n5888# 0.015589f
C986 source.n788 a_n2102_n5888# 0.015589f
C987 source.n789 a_n2102_n5888# 0.016506f
C988 source.n790 a_n2102_n5888# 0.036847f
C989 source.n791 a_n2102_n5888# 0.036847f
C990 source.n792 a_n2102_n5888# 0.036847f
C991 source.n793 a_n2102_n5888# 0.016048f
C992 source.n794 a_n2102_n5888# 0.015589f
C993 source.n795 a_n2102_n5888# 0.029011f
C994 source.n796 a_n2102_n5888# 0.029011f
C995 source.n797 a_n2102_n5888# 0.015589f
C996 source.n798 a_n2102_n5888# 0.016506f
C997 source.n799 a_n2102_n5888# 0.036847f
C998 source.n800 a_n2102_n5888# 0.036847f
C999 source.n801 a_n2102_n5888# 0.016506f
C1000 source.n802 a_n2102_n5888# 0.015589f
C1001 source.n803 a_n2102_n5888# 0.029011f
C1002 source.n804 a_n2102_n5888# 0.029011f
C1003 source.n805 a_n2102_n5888# 0.015589f
C1004 source.n806 a_n2102_n5888# 0.016506f
C1005 source.n807 a_n2102_n5888# 0.036847f
C1006 source.n808 a_n2102_n5888# 0.036847f
C1007 source.n809 a_n2102_n5888# 0.016506f
C1008 source.n810 a_n2102_n5888# 0.015589f
C1009 source.n811 a_n2102_n5888# 0.029011f
C1010 source.n812 a_n2102_n5888# 0.029011f
C1011 source.n813 a_n2102_n5888# 0.015589f
C1012 source.n814 a_n2102_n5888# 0.016506f
C1013 source.n815 a_n2102_n5888# 0.036847f
C1014 source.n816 a_n2102_n5888# 0.036847f
C1015 source.n817 a_n2102_n5888# 0.016506f
C1016 source.n818 a_n2102_n5888# 0.015589f
C1017 source.n819 a_n2102_n5888# 0.029011f
C1018 source.n820 a_n2102_n5888# 0.029011f
C1019 source.n821 a_n2102_n5888# 0.015589f
C1020 source.n822 a_n2102_n5888# 0.016506f
C1021 source.n823 a_n2102_n5888# 0.036847f
C1022 source.n824 a_n2102_n5888# 0.036847f
C1023 source.n825 a_n2102_n5888# 0.016506f
C1024 source.n826 a_n2102_n5888# 0.015589f
C1025 source.n827 a_n2102_n5888# 0.029011f
C1026 source.n828 a_n2102_n5888# 0.029011f
C1027 source.n829 a_n2102_n5888# 0.015589f
C1028 source.n830 a_n2102_n5888# 0.016506f
C1029 source.n831 a_n2102_n5888# 0.036847f
C1030 source.n832 a_n2102_n5888# 0.036847f
C1031 source.n833 a_n2102_n5888# 0.036847f
C1032 source.n834 a_n2102_n5888# 0.016506f
C1033 source.n835 a_n2102_n5888# 0.015589f
C1034 source.n836 a_n2102_n5888# 0.029011f
C1035 source.n837 a_n2102_n5888# 0.029011f
C1036 source.n838 a_n2102_n5888# 0.015589f
C1037 source.n839 a_n2102_n5888# 0.016048f
C1038 source.n840 a_n2102_n5888# 0.016048f
C1039 source.n841 a_n2102_n5888# 0.036847f
C1040 source.n842 a_n2102_n5888# 0.036847f
C1041 source.n843 a_n2102_n5888# 0.016506f
C1042 source.n844 a_n2102_n5888# 0.015589f
C1043 source.n845 a_n2102_n5888# 0.029011f
C1044 source.n846 a_n2102_n5888# 0.029011f
C1045 source.n847 a_n2102_n5888# 0.015589f
C1046 source.n848 a_n2102_n5888# 0.016506f
C1047 source.n849 a_n2102_n5888# 0.036847f
C1048 source.n850 a_n2102_n5888# 0.036847f
C1049 source.n851 a_n2102_n5888# 0.016506f
C1050 source.n852 a_n2102_n5888# 0.015589f
C1051 source.n853 a_n2102_n5888# 0.029011f
C1052 source.n854 a_n2102_n5888# 0.029011f
C1053 source.n855 a_n2102_n5888# 0.015589f
C1054 source.n856 a_n2102_n5888# 0.016506f
C1055 source.n857 a_n2102_n5888# 0.036847f
C1056 source.n858 a_n2102_n5888# 0.078383f
C1057 source.n859 a_n2102_n5888# 0.016506f
C1058 source.n860 a_n2102_n5888# 0.015589f
C1059 source.n861 a_n2102_n5888# 0.063887f
C1060 source.n862 a_n2102_n5888# 0.043617f
C1061 source.n863 a_n2102_n5888# 0.117678f
C1062 source.n864 a_n2102_n5888# 0.039994f
C1063 source.n865 a_n2102_n5888# 0.029011f
C1064 source.n866 a_n2102_n5888# 0.015589f
C1065 source.n867 a_n2102_n5888# 0.036847f
C1066 source.n868 a_n2102_n5888# 0.016506f
C1067 source.n869 a_n2102_n5888# 0.029011f
C1068 source.n870 a_n2102_n5888# 0.015589f
C1069 source.n871 a_n2102_n5888# 0.036847f
C1070 source.n872 a_n2102_n5888# 0.016506f
C1071 source.n873 a_n2102_n5888# 0.029011f
C1072 source.n874 a_n2102_n5888# 0.015589f
C1073 source.n875 a_n2102_n5888# 0.036847f
C1074 source.n876 a_n2102_n5888# 0.016506f
C1075 source.n877 a_n2102_n5888# 0.029011f
C1076 source.n878 a_n2102_n5888# 0.015589f
C1077 source.n879 a_n2102_n5888# 0.036847f
C1078 source.n880 a_n2102_n5888# 0.016506f
C1079 source.n881 a_n2102_n5888# 0.029011f
C1080 source.n882 a_n2102_n5888# 0.015589f
C1081 source.n883 a_n2102_n5888# 0.036847f
C1082 source.n884 a_n2102_n5888# 0.016506f
C1083 source.n885 a_n2102_n5888# 0.029011f
C1084 source.n886 a_n2102_n5888# 0.015589f
C1085 source.n887 a_n2102_n5888# 0.036847f
C1086 source.n888 a_n2102_n5888# 0.016506f
C1087 source.n889 a_n2102_n5888# 0.029011f
C1088 source.n890 a_n2102_n5888# 0.015589f
C1089 source.n891 a_n2102_n5888# 0.036847f
C1090 source.n892 a_n2102_n5888# 0.016506f
C1091 source.n893 a_n2102_n5888# 0.029011f
C1092 source.n894 a_n2102_n5888# 0.015589f
C1093 source.n895 a_n2102_n5888# 0.036847f
C1094 source.n896 a_n2102_n5888# 0.016506f
C1095 source.n897 a_n2102_n5888# 0.029011f
C1096 source.n898 a_n2102_n5888# 0.016048f
C1097 source.n899 a_n2102_n5888# 0.036847f
C1098 source.n900 a_n2102_n5888# 0.016506f
C1099 source.n901 a_n2102_n5888# 0.029011f
C1100 source.n902 a_n2102_n5888# 0.015589f
C1101 source.n903 a_n2102_n5888# 0.036847f
C1102 source.n904 a_n2102_n5888# 0.016506f
C1103 source.n905 a_n2102_n5888# 0.029011f
C1104 source.n906 a_n2102_n5888# 0.015589f
C1105 source.n907 a_n2102_n5888# 0.027635f
C1106 source.n908 a_n2102_n5888# 0.026048f
C1107 source.t13 a_n2102_n5888# 0.064264f
C1108 source.n909 a_n2102_n5888# 0.353956f
C1109 source.n910 a_n2102_n5888# 3.14101f
C1110 source.n911 a_n2102_n5888# 0.015589f
C1111 source.n912 a_n2102_n5888# 0.016506f
C1112 source.n913 a_n2102_n5888# 0.036847f
C1113 source.n914 a_n2102_n5888# 0.036847f
C1114 source.n915 a_n2102_n5888# 0.016506f
C1115 source.n916 a_n2102_n5888# 0.015589f
C1116 source.n917 a_n2102_n5888# 0.029011f
C1117 source.n918 a_n2102_n5888# 0.029011f
C1118 source.n919 a_n2102_n5888# 0.015589f
C1119 source.n920 a_n2102_n5888# 0.016506f
C1120 source.n921 a_n2102_n5888# 0.036847f
C1121 source.n922 a_n2102_n5888# 0.036847f
C1122 source.n923 a_n2102_n5888# 0.016506f
C1123 source.n924 a_n2102_n5888# 0.015589f
C1124 source.n925 a_n2102_n5888# 0.029011f
C1125 source.n926 a_n2102_n5888# 0.029011f
C1126 source.n927 a_n2102_n5888# 0.015589f
C1127 source.n928 a_n2102_n5888# 0.015589f
C1128 source.n929 a_n2102_n5888# 0.016506f
C1129 source.n930 a_n2102_n5888# 0.036847f
C1130 source.n931 a_n2102_n5888# 0.036847f
C1131 source.n932 a_n2102_n5888# 0.036847f
C1132 source.n933 a_n2102_n5888# 0.016048f
C1133 source.n934 a_n2102_n5888# 0.015589f
C1134 source.n935 a_n2102_n5888# 0.029011f
C1135 source.n936 a_n2102_n5888# 0.029011f
C1136 source.n937 a_n2102_n5888# 0.015589f
C1137 source.n938 a_n2102_n5888# 0.016506f
C1138 source.n939 a_n2102_n5888# 0.036847f
C1139 source.n940 a_n2102_n5888# 0.036847f
C1140 source.n941 a_n2102_n5888# 0.016506f
C1141 source.n942 a_n2102_n5888# 0.015589f
C1142 source.n943 a_n2102_n5888# 0.029011f
C1143 source.n944 a_n2102_n5888# 0.029011f
C1144 source.n945 a_n2102_n5888# 0.015589f
C1145 source.n946 a_n2102_n5888# 0.016506f
C1146 source.n947 a_n2102_n5888# 0.036847f
C1147 source.n948 a_n2102_n5888# 0.036847f
C1148 source.n949 a_n2102_n5888# 0.016506f
C1149 source.n950 a_n2102_n5888# 0.015589f
C1150 source.n951 a_n2102_n5888# 0.029011f
C1151 source.n952 a_n2102_n5888# 0.029011f
C1152 source.n953 a_n2102_n5888# 0.015589f
C1153 source.n954 a_n2102_n5888# 0.016506f
C1154 source.n955 a_n2102_n5888# 0.036847f
C1155 source.n956 a_n2102_n5888# 0.036847f
C1156 source.n957 a_n2102_n5888# 0.016506f
C1157 source.n958 a_n2102_n5888# 0.015589f
C1158 source.n959 a_n2102_n5888# 0.029011f
C1159 source.n960 a_n2102_n5888# 0.029011f
C1160 source.n961 a_n2102_n5888# 0.015589f
C1161 source.n962 a_n2102_n5888# 0.016506f
C1162 source.n963 a_n2102_n5888# 0.036847f
C1163 source.n964 a_n2102_n5888# 0.036847f
C1164 source.n965 a_n2102_n5888# 0.016506f
C1165 source.n966 a_n2102_n5888# 0.015589f
C1166 source.n967 a_n2102_n5888# 0.029011f
C1167 source.n968 a_n2102_n5888# 0.029011f
C1168 source.n969 a_n2102_n5888# 0.015589f
C1169 source.n970 a_n2102_n5888# 0.016506f
C1170 source.n971 a_n2102_n5888# 0.036847f
C1171 source.n972 a_n2102_n5888# 0.036847f
C1172 source.n973 a_n2102_n5888# 0.036847f
C1173 source.n974 a_n2102_n5888# 0.016506f
C1174 source.n975 a_n2102_n5888# 0.015589f
C1175 source.n976 a_n2102_n5888# 0.029011f
C1176 source.n977 a_n2102_n5888# 0.029011f
C1177 source.n978 a_n2102_n5888# 0.015589f
C1178 source.n979 a_n2102_n5888# 0.016048f
C1179 source.n980 a_n2102_n5888# 0.016048f
C1180 source.n981 a_n2102_n5888# 0.036847f
C1181 source.n982 a_n2102_n5888# 0.036847f
C1182 source.n983 a_n2102_n5888# 0.016506f
C1183 source.n984 a_n2102_n5888# 0.015589f
C1184 source.n985 a_n2102_n5888# 0.029011f
C1185 source.n986 a_n2102_n5888# 0.029011f
C1186 source.n987 a_n2102_n5888# 0.015589f
C1187 source.n988 a_n2102_n5888# 0.016506f
C1188 source.n989 a_n2102_n5888# 0.036847f
C1189 source.n990 a_n2102_n5888# 0.036847f
C1190 source.n991 a_n2102_n5888# 0.016506f
C1191 source.n992 a_n2102_n5888# 0.015589f
C1192 source.n993 a_n2102_n5888# 0.029011f
C1193 source.n994 a_n2102_n5888# 0.029011f
C1194 source.n995 a_n2102_n5888# 0.015589f
C1195 source.n996 a_n2102_n5888# 0.016506f
C1196 source.n997 a_n2102_n5888# 0.036847f
C1197 source.n998 a_n2102_n5888# 0.078383f
C1198 source.n999 a_n2102_n5888# 0.016506f
C1199 source.n1000 a_n2102_n5888# 0.015589f
C1200 source.n1001 a_n2102_n5888# 0.063887f
C1201 source.n1002 a_n2102_n5888# 0.043617f
C1202 source.n1003 a_n2102_n5888# 0.117678f
C1203 source.t10 a_n2102_n5888# 0.57313f
C1204 source.t11 a_n2102_n5888# 0.57313f
C1205 source.n1004 a_n2102_n5888# 5.18691f
C1206 source.n1005 a_n2102_n5888# 0.402439f
C1207 source.t16 a_n2102_n5888# 0.57313f
C1208 source.t3 a_n2102_n5888# 0.57313f
C1209 source.n1006 a_n2102_n5888# 5.18691f
C1210 source.n1007 a_n2102_n5888# 0.402439f
C1211 source.t17 a_n2102_n5888# 0.57313f
C1212 source.t39 a_n2102_n5888# 0.57313f
C1213 source.n1008 a_n2102_n5888# 5.18691f
C1214 source.n1009 a_n2102_n5888# 0.402439f
C1215 source.t15 a_n2102_n5888# 0.57313f
C1216 source.t6 a_n2102_n5888# 0.57313f
C1217 source.n1010 a_n2102_n5888# 5.18691f
C1218 source.n1011 a_n2102_n5888# 0.402439f
C1219 source.n1012 a_n2102_n5888# 0.039994f
C1220 source.n1013 a_n2102_n5888# 0.029011f
C1221 source.n1014 a_n2102_n5888# 0.015589f
C1222 source.n1015 a_n2102_n5888# 0.036847f
C1223 source.n1016 a_n2102_n5888# 0.016506f
C1224 source.n1017 a_n2102_n5888# 0.029011f
C1225 source.n1018 a_n2102_n5888# 0.015589f
C1226 source.n1019 a_n2102_n5888# 0.036847f
C1227 source.n1020 a_n2102_n5888# 0.016506f
C1228 source.n1021 a_n2102_n5888# 0.029011f
C1229 source.n1022 a_n2102_n5888# 0.015589f
C1230 source.n1023 a_n2102_n5888# 0.036847f
C1231 source.n1024 a_n2102_n5888# 0.016506f
C1232 source.n1025 a_n2102_n5888# 0.029011f
C1233 source.n1026 a_n2102_n5888# 0.015589f
C1234 source.n1027 a_n2102_n5888# 0.036847f
C1235 source.n1028 a_n2102_n5888# 0.016506f
C1236 source.n1029 a_n2102_n5888# 0.029011f
C1237 source.n1030 a_n2102_n5888# 0.015589f
C1238 source.n1031 a_n2102_n5888# 0.036847f
C1239 source.n1032 a_n2102_n5888# 0.016506f
C1240 source.n1033 a_n2102_n5888# 0.029011f
C1241 source.n1034 a_n2102_n5888# 0.015589f
C1242 source.n1035 a_n2102_n5888# 0.036847f
C1243 source.n1036 a_n2102_n5888# 0.016506f
C1244 source.n1037 a_n2102_n5888# 0.029011f
C1245 source.n1038 a_n2102_n5888# 0.015589f
C1246 source.n1039 a_n2102_n5888# 0.036847f
C1247 source.n1040 a_n2102_n5888# 0.016506f
C1248 source.n1041 a_n2102_n5888# 0.029011f
C1249 source.n1042 a_n2102_n5888# 0.015589f
C1250 source.n1043 a_n2102_n5888# 0.036847f
C1251 source.n1044 a_n2102_n5888# 0.016506f
C1252 source.n1045 a_n2102_n5888# 0.029011f
C1253 source.n1046 a_n2102_n5888# 0.016048f
C1254 source.n1047 a_n2102_n5888# 0.036847f
C1255 source.n1048 a_n2102_n5888# 0.016506f
C1256 source.n1049 a_n2102_n5888# 0.029011f
C1257 source.n1050 a_n2102_n5888# 0.015589f
C1258 source.n1051 a_n2102_n5888# 0.036847f
C1259 source.n1052 a_n2102_n5888# 0.016506f
C1260 source.n1053 a_n2102_n5888# 0.029011f
C1261 source.n1054 a_n2102_n5888# 0.015589f
C1262 source.n1055 a_n2102_n5888# 0.027635f
C1263 source.n1056 a_n2102_n5888# 0.026048f
C1264 source.t14 a_n2102_n5888# 0.064264f
C1265 source.n1057 a_n2102_n5888# 0.353956f
C1266 source.n1058 a_n2102_n5888# 3.14101f
C1267 source.n1059 a_n2102_n5888# 0.015589f
C1268 source.n1060 a_n2102_n5888# 0.016506f
C1269 source.n1061 a_n2102_n5888# 0.036847f
C1270 source.n1062 a_n2102_n5888# 0.036847f
C1271 source.n1063 a_n2102_n5888# 0.016506f
C1272 source.n1064 a_n2102_n5888# 0.015589f
C1273 source.n1065 a_n2102_n5888# 0.029011f
C1274 source.n1066 a_n2102_n5888# 0.029011f
C1275 source.n1067 a_n2102_n5888# 0.015589f
C1276 source.n1068 a_n2102_n5888# 0.016506f
C1277 source.n1069 a_n2102_n5888# 0.036847f
C1278 source.n1070 a_n2102_n5888# 0.036847f
C1279 source.n1071 a_n2102_n5888# 0.016506f
C1280 source.n1072 a_n2102_n5888# 0.015589f
C1281 source.n1073 a_n2102_n5888# 0.029011f
C1282 source.n1074 a_n2102_n5888# 0.029011f
C1283 source.n1075 a_n2102_n5888# 0.015589f
C1284 source.n1076 a_n2102_n5888# 0.015589f
C1285 source.n1077 a_n2102_n5888# 0.016506f
C1286 source.n1078 a_n2102_n5888# 0.036847f
C1287 source.n1079 a_n2102_n5888# 0.036847f
C1288 source.n1080 a_n2102_n5888# 0.036847f
C1289 source.n1081 a_n2102_n5888# 0.016048f
C1290 source.n1082 a_n2102_n5888# 0.015589f
C1291 source.n1083 a_n2102_n5888# 0.029011f
C1292 source.n1084 a_n2102_n5888# 0.029011f
C1293 source.n1085 a_n2102_n5888# 0.015589f
C1294 source.n1086 a_n2102_n5888# 0.016506f
C1295 source.n1087 a_n2102_n5888# 0.036847f
C1296 source.n1088 a_n2102_n5888# 0.036847f
C1297 source.n1089 a_n2102_n5888# 0.016506f
C1298 source.n1090 a_n2102_n5888# 0.015589f
C1299 source.n1091 a_n2102_n5888# 0.029011f
C1300 source.n1092 a_n2102_n5888# 0.029011f
C1301 source.n1093 a_n2102_n5888# 0.015589f
C1302 source.n1094 a_n2102_n5888# 0.016506f
C1303 source.n1095 a_n2102_n5888# 0.036847f
C1304 source.n1096 a_n2102_n5888# 0.036847f
C1305 source.n1097 a_n2102_n5888# 0.016506f
C1306 source.n1098 a_n2102_n5888# 0.015589f
C1307 source.n1099 a_n2102_n5888# 0.029011f
C1308 source.n1100 a_n2102_n5888# 0.029011f
C1309 source.n1101 a_n2102_n5888# 0.015589f
C1310 source.n1102 a_n2102_n5888# 0.016506f
C1311 source.n1103 a_n2102_n5888# 0.036847f
C1312 source.n1104 a_n2102_n5888# 0.036847f
C1313 source.n1105 a_n2102_n5888# 0.016506f
C1314 source.n1106 a_n2102_n5888# 0.015589f
C1315 source.n1107 a_n2102_n5888# 0.029011f
C1316 source.n1108 a_n2102_n5888# 0.029011f
C1317 source.n1109 a_n2102_n5888# 0.015589f
C1318 source.n1110 a_n2102_n5888# 0.016506f
C1319 source.n1111 a_n2102_n5888# 0.036847f
C1320 source.n1112 a_n2102_n5888# 0.036847f
C1321 source.n1113 a_n2102_n5888# 0.016506f
C1322 source.n1114 a_n2102_n5888# 0.015589f
C1323 source.n1115 a_n2102_n5888# 0.029011f
C1324 source.n1116 a_n2102_n5888# 0.029011f
C1325 source.n1117 a_n2102_n5888# 0.015589f
C1326 source.n1118 a_n2102_n5888# 0.016506f
C1327 source.n1119 a_n2102_n5888# 0.036847f
C1328 source.n1120 a_n2102_n5888# 0.036847f
C1329 source.n1121 a_n2102_n5888# 0.036847f
C1330 source.n1122 a_n2102_n5888# 0.016506f
C1331 source.n1123 a_n2102_n5888# 0.015589f
C1332 source.n1124 a_n2102_n5888# 0.029011f
C1333 source.n1125 a_n2102_n5888# 0.029011f
C1334 source.n1126 a_n2102_n5888# 0.015589f
C1335 source.n1127 a_n2102_n5888# 0.016048f
C1336 source.n1128 a_n2102_n5888# 0.016048f
C1337 source.n1129 a_n2102_n5888# 0.036847f
C1338 source.n1130 a_n2102_n5888# 0.036847f
C1339 source.n1131 a_n2102_n5888# 0.016506f
C1340 source.n1132 a_n2102_n5888# 0.015589f
C1341 source.n1133 a_n2102_n5888# 0.029011f
C1342 source.n1134 a_n2102_n5888# 0.029011f
C1343 source.n1135 a_n2102_n5888# 0.015589f
C1344 source.n1136 a_n2102_n5888# 0.016506f
C1345 source.n1137 a_n2102_n5888# 0.036847f
C1346 source.n1138 a_n2102_n5888# 0.036847f
C1347 source.n1139 a_n2102_n5888# 0.016506f
C1348 source.n1140 a_n2102_n5888# 0.015589f
C1349 source.n1141 a_n2102_n5888# 0.029011f
C1350 source.n1142 a_n2102_n5888# 0.029011f
C1351 source.n1143 a_n2102_n5888# 0.015589f
C1352 source.n1144 a_n2102_n5888# 0.016506f
C1353 source.n1145 a_n2102_n5888# 0.036847f
C1354 source.n1146 a_n2102_n5888# 0.078383f
C1355 source.n1147 a_n2102_n5888# 0.016506f
C1356 source.n1148 a_n2102_n5888# 0.015589f
C1357 source.n1149 a_n2102_n5888# 0.063887f
C1358 source.n1150 a_n2102_n5888# 0.043617f
C1359 source.n1151 a_n2102_n5888# 0.281444f
C1360 source.n1152 a_n2102_n5888# 3.09259f
C1361 plus.n0 a_n2102_n5888# 0.050015f
C1362 plus.t7 a_n2102_n5888# 1.05545f
C1363 plus.t0 a_n2102_n5888# 1.05545f
C1364 plus.n1 a_n2102_n5888# 0.018288f
C1365 plus.n2 a_n2102_n5888# 0.050015f
C1366 plus.t9 a_n2102_n5888# 1.05545f
C1367 plus.t5 a_n2102_n5888# 1.05545f
C1368 plus.t17 a_n2102_n5888# 1.05545f
C1369 plus.n3 a_n2102_n5888# 0.384054f
C1370 plus.n4 a_n2102_n5888# 0.050015f
C1371 plus.t11 a_n2102_n5888# 1.05545f
C1372 plus.t6 a_n2102_n5888# 1.05545f
C1373 plus.n5 a_n2102_n5888# 0.384054f
C1374 plus.t1 a_n2102_n5888# 1.06424f
C1375 plus.n6 a_n2102_n5888# 0.400106f
C1376 plus.n7 a_n2102_n5888# 0.114448f
C1377 plus.n8 a_n2102_n5888# 0.0206f
C1378 plus.n9 a_n2102_n5888# 0.384054f
C1379 plus.n10 a_n2102_n5888# 0.018904f
C1380 plus.n11 a_n2102_n5888# 0.018288f
C1381 plus.n12 a_n2102_n5888# 0.050015f
C1382 plus.n13 a_n2102_n5888# 0.050015f
C1383 plus.n14 a_n2102_n5888# 0.0206f
C1384 plus.n15 a_n2102_n5888# 0.384054f
C1385 plus.n16 a_n2102_n5888# 0.0206f
C1386 plus.n17 a_n2102_n5888# 0.384054f
C1387 plus.t16 a_n2102_n5888# 1.05545f
C1388 plus.n18 a_n2102_n5888# 0.384054f
C1389 plus.n19 a_n2102_n5888# 0.0206f
C1390 plus.n20 a_n2102_n5888# 0.050015f
C1391 plus.n21 a_n2102_n5888# 0.050015f
C1392 plus.n22 a_n2102_n5888# 0.050015f
C1393 plus.n23 a_n2102_n5888# 0.018904f
C1394 plus.n24 a_n2102_n5888# 0.384054f
C1395 plus.n25 a_n2102_n5888# 0.0206f
C1396 plus.n26 a_n2102_n5888# 0.384054f
C1397 plus.t13 a_n2102_n5888# 1.06424f
C1398 plus.n27 a_n2102_n5888# 0.40003f
C1399 plus.n28 a_n2102_n5888# 0.894561f
C1400 plus.n29 a_n2102_n5888# 0.050015f
C1401 plus.t15 a_n2102_n5888# 1.06424f
C1402 plus.t2 a_n2102_n5888# 1.05545f
C1403 plus.t14 a_n2102_n5888# 1.05545f
C1404 plus.n30 a_n2102_n5888# 0.018288f
C1405 plus.n31 a_n2102_n5888# 0.050015f
C1406 plus.t4 a_n2102_n5888# 1.05545f
C1407 plus.n32 a_n2102_n5888# 0.384054f
C1408 plus.t12 a_n2102_n5888# 1.05545f
C1409 plus.t3 a_n2102_n5888# 1.05545f
C1410 plus.t10 a_n2102_n5888# 1.05545f
C1411 plus.n33 a_n2102_n5888# 0.384054f
C1412 plus.n34 a_n2102_n5888# 0.050015f
C1413 plus.t19 a_n2102_n5888# 1.05545f
C1414 plus.t8 a_n2102_n5888# 1.05545f
C1415 plus.n35 a_n2102_n5888# 0.384054f
C1416 plus.t18 a_n2102_n5888# 1.06424f
C1417 plus.n36 a_n2102_n5888# 0.400106f
C1418 plus.n37 a_n2102_n5888# 0.114448f
C1419 plus.n38 a_n2102_n5888# 0.0206f
C1420 plus.n39 a_n2102_n5888# 0.384054f
C1421 plus.n40 a_n2102_n5888# 0.018904f
C1422 plus.n41 a_n2102_n5888# 0.018288f
C1423 plus.n42 a_n2102_n5888# 0.050015f
C1424 plus.n43 a_n2102_n5888# 0.050015f
C1425 plus.n44 a_n2102_n5888# 0.0206f
C1426 plus.n45 a_n2102_n5888# 0.384054f
C1427 plus.n46 a_n2102_n5888# 0.0206f
C1428 plus.n47 a_n2102_n5888# 0.384054f
C1429 plus.n48 a_n2102_n5888# 0.0206f
C1430 plus.n49 a_n2102_n5888# 0.050015f
C1431 plus.n50 a_n2102_n5888# 0.050015f
C1432 plus.n51 a_n2102_n5888# 0.050015f
C1433 plus.n52 a_n2102_n5888# 0.018904f
C1434 plus.n53 a_n2102_n5888# 0.384054f
C1435 plus.n54 a_n2102_n5888# 0.0206f
C1436 plus.n55 a_n2102_n5888# 0.384054f
C1437 plus.n56 a_n2102_n5888# 0.40003f
C1438 plus.n57 a_n2102_n5888# 1.99953f
.ends

