* NGSPICE file created from diffpair644.ext - technology: sky130A

.subckt diffpair644 minus drain_right drain_left source plus
X0 source.t17 minus.t0 drain_right.t7 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 drain_right.t5 minus.t1 source.t16 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X2 drain_left.t9 plus.t0 source.t5 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X3 a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X4 a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X5 source.t15 minus.t2 drain_right.t4 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X6 source.t7 plus.t1 drain_left.t8 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X7 drain_right.t8 minus.t3 source.t14 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X8 drain_right.t2 minus.t4 source.t13 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X9 drain_right.t0 minus.t5 source.t12 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X10 drain_left.t7 plus.t2 source.t6 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X11 source.t11 minus.t6 drain_right.t1 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X12 a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X13 drain_left.t6 plus.t3 source.t0 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X14 drain_left.t5 plus.t4 source.t4 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X15 drain_right.t3 minus.t7 source.t10 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X16 source.t9 minus.t8 drain_right.t6 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 source.t1 plus.t5 drain_left.t4 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X18 source.t3 plus.t6 drain_left.t3 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 drain_left.t2 plus.t7 source.t2 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X20 source.t18 plus.t8 drain_left.t1 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X21 drain_right.t9 minus.t9 source.t8 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 drain_left.t0 plus.t9 source.t19 a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X23 a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# a_n1496_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
R0 minus.n9 minus.t4 4269.35
R1 minus.n3 minus.t3 4269.35
R2 minus.n20 minus.t5 4269.35
R3 minus.n14 minus.t1 4269.35
R4 minus.n6 minus.t7 4225.53
R5 minus.n8 minus.t6 4225.53
R6 minus.n2 minus.t2 4225.53
R7 minus.n17 minus.t9 4225.53
R8 minus.n19 minus.t0 4225.53
R9 minus.n13 minus.t8 4225.53
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 44.6501
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t5 60.4756
R42 drain_right.n7 drain_right.t2 59.9154
R43 drain_right.n6 drain_right.n4 59.2756
R44 drain_right.n3 drain_right.n2 59.0803
R45 drain_right.n1 drain_right.n0 58.7154
R46 drain_right.n6 drain_right.n5 58.7154
R47 drain_right drain_right.n3 39.0438
R48 drain_right drain_right.n7 5.93339
R49 drain_right.n2 drain_right.t7 1.2005
R50 drain_right.n2 drain_right.t0 1.2005
R51 drain_right.n0 drain_right.t6 1.2005
R52 drain_right.n0 drain_right.t9 1.2005
R53 drain_right.n4 drain_right.t4 1.2005
R54 drain_right.n4 drain_right.t8 1.2005
R55 drain_right.n5 drain_right.t1 1.2005
R56 drain_right.n5 drain_right.t3 1.2005
R57 drain_right.n7 drain_right.n6 0.560845
R58 drain_right.n3 drain_right.n1 0.0852402
R59 source.n5 source.t14 43.2366
R60 source.n19 source.t12 43.2365
R61 source.n14 source.t6 43.2365
R62 source.n0 source.t19 43.2365
R63 source.n18 source.n17 42.0366
R64 source.n16 source.n15 42.0366
R65 source.n13 source.n12 42.0366
R66 source.n11 source.n10 42.0366
R67 source.n2 source.n1 42.0366
R68 source.n4 source.n3 42.0366
R69 source.n7 source.n6 42.0366
R70 source.n9 source.n8 42.0366
R71 source.n11 source.n9 32.2569
R72 source.n20 source.n0 26.1535
R73 source.n20 source.n19 5.5436
R74 source.n17 source.t8 1.2005
R75 source.n17 source.t17 1.2005
R76 source.n15 source.t16 1.2005
R77 source.n15 source.t9 1.2005
R78 source.n12 source.t5 1.2005
R79 source.n12 source.t3 1.2005
R80 source.n10 source.t0 1.2005
R81 source.n10 source.t7 1.2005
R82 source.n1 source.t2 1.2005
R83 source.n1 source.t1 1.2005
R84 source.n3 source.t4 1.2005
R85 source.n3 source.t18 1.2005
R86 source.n6 source.t10 1.2005
R87 source.n6 source.t15 1.2005
R88 source.n8 source.t13 1.2005
R89 source.n8 source.t11 1.2005
R90 source.n5 source.n4 0.7505
R91 source.n16 source.n14 0.7505
R92 source.n9 source.n7 0.560845
R93 source.n7 source.n5 0.560845
R94 source.n4 source.n2 0.560845
R95 source.n2 source.n0 0.560845
R96 source.n13 source.n11 0.560845
R97 source.n14 source.n13 0.560845
R98 source.n18 source.n16 0.560845
R99 source.n19 source.n18 0.560845
R100 source source.n20 0.188
R101 plus.n3 plus.t4 4269.35
R102 plus.n9 plus.t9 4269.35
R103 plus.n14 plus.t2 4269.35
R104 plus.n20 plus.t3 4269.35
R105 plus.n6 plus.t7 4225.53
R106 plus.n2 plus.t8 4225.53
R107 plus.n8 plus.t5 4225.53
R108 plus.n17 plus.t0 4225.53
R109 plus.n13 plus.t6 4225.53
R110 plus.n19 plus.t1 4225.53
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 33.607
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 17.0819
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t5 60.4758
R142 drain_left.n1 drain_left.t6 60.4756
R143 drain_left.n3 drain_left.n2 59.0803
R144 drain_left.n1 drain_left.n0 58.7154
R145 drain_left.n5 drain_left.n4 58.7154
R146 drain_left.n7 drain_left.n6 58.7153
R147 drain_left drain_left.n3 39.597
R148 drain_left drain_left.n7 6.21356
R149 drain_left.n2 drain_left.t3 1.2005
R150 drain_left.n2 drain_left.t7 1.2005
R151 drain_left.n0 drain_left.t8 1.2005
R152 drain_left.n0 drain_left.t9 1.2005
R153 drain_left.n6 drain_left.t4 1.2005
R154 drain_left.n6 drain_left.t0 1.2005
R155 drain_left.n4 drain_left.t1 1.2005
R156 drain_left.n4 drain_left.t2 1.2005
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 source plus 3.68136f
C1 plus minus 7.41088f
C2 drain_right plus 0.300949f
C3 source drain_left 42.3408f
C4 minus drain_left 0.170828f
C5 drain_right drain_left 0.741659f
C6 source minus 3.66598f
C7 drain_right source 42.319702f
C8 plus drain_left 4.96057f
C9 drain_right minus 4.82342f
C10 drain_right a_n1496_n5888# 10.12675f
C11 drain_left a_n1496_n5888# 10.3683f
C12 source a_n1496_n5888# 10.689644f
C13 minus a_n1496_n5888# 6.377497f
C14 plus a_n1496_n5888# 9.57259f
C15 drain_left.t6 a_n1496_n5888# 6.40384f
C16 drain_left.t8 a_n1496_n5888# 0.760928f
C17 drain_left.t9 a_n1496_n5888# 0.760928f
C18 drain_left.n0 a_n1496_n5888# 5.14586f
C19 drain_left.n1 a_n1496_n5888# 0.657384f
C20 drain_left.t3 a_n1496_n5888# 0.760928f
C21 drain_left.t7 a_n1496_n5888# 0.760928f
C22 drain_left.n2 a_n1496_n5888# 5.14773f
C23 drain_left.n3 a_n1496_n5888# 2.28529f
C24 drain_left.t5 a_n1496_n5888# 6.40385f
C25 drain_left.t1 a_n1496_n5888# 0.760928f
C26 drain_left.t2 a_n1496_n5888# 0.760928f
C27 drain_left.n4 a_n1496_n5888# 5.14586f
C28 drain_left.n5 a_n1496_n5888# 0.689374f
C29 drain_left.t4 a_n1496_n5888# 0.760928f
C30 drain_left.t0 a_n1496_n5888# 0.760928f
C31 drain_left.n6 a_n1496_n5888# 5.14585f
C32 drain_left.n7 a_n1496_n5888# 0.518983f
C33 plus.n0 a_n1496_n5888# 0.059917f
C34 plus.t5 a_n1496_n5888# 0.6322f
C35 plus.t7 a_n1496_n5888# 0.6322f
C36 plus.n1 a_n1496_n5888# 0.025418f
C37 plus.t4 a_n1496_n5888# 0.634637f
C38 plus.t8 a_n1496_n5888# 0.6322f
C39 plus.n2 a_n1496_n5888# 0.239279f
C40 plus.n3 a_n1496_n5888# 0.260493f
C41 plus.n4 a_n1496_n5888# 0.128988f
C42 plus.n5 a_n1496_n5888# 0.059917f
C43 plus.n6 a_n1496_n5888# 0.259155f
C44 plus.n7 a_n1496_n5888# 0.025418f
C45 plus.n8 a_n1496_n5888# 0.239279f
C46 plus.t9 a_n1496_n5888# 0.634637f
C47 plus.n9 a_n1496_n5888# 0.260412f
C48 plus.n10 a_n1496_n5888# 1.07141f
C49 plus.n11 a_n1496_n5888# 0.059917f
C50 plus.t3 a_n1496_n5888# 0.634637f
C51 plus.t1 a_n1496_n5888# 0.6322f
C52 plus.t0 a_n1496_n5888# 0.6322f
C53 plus.n12 a_n1496_n5888# 0.025418f
C54 plus.t6 a_n1496_n5888# 0.6322f
C55 plus.n13 a_n1496_n5888# 0.239279f
C56 plus.t2 a_n1496_n5888# 0.634637f
C57 plus.n14 a_n1496_n5888# 0.260493f
C58 plus.n15 a_n1496_n5888# 0.128988f
C59 plus.n16 a_n1496_n5888# 0.059917f
C60 plus.n17 a_n1496_n5888# 0.259155f
C61 plus.n18 a_n1496_n5888# 0.025418f
C62 plus.n19 a_n1496_n5888# 0.239279f
C63 plus.n20 a_n1496_n5888# 0.260412f
C64 plus.n21 a_n1496_n5888# 2.20714f
C65 source.t19 a_n1496_n5888# 6.25299f
C66 source.n0 a_n1496_n5888# 2.39269f
C67 source.t2 a_n1496_n5888# 0.758287f
C68 source.t1 a_n1496_n5888# 0.758287f
C69 source.n1 a_n1496_n5888# 5.04495f
C70 source.n2 a_n1496_n5888# 0.354231f
C71 source.t4 a_n1496_n5888# 0.758287f
C72 source.t18 a_n1496_n5888# 0.758287f
C73 source.n3 a_n1496_n5888# 5.04495f
C74 source.n4 a_n1496_n5888# 0.369713f
C75 source.t14 a_n1496_n5888# 6.25301f
C76 source.n5 a_n1496_n5888# 0.52657f
C77 source.t10 a_n1496_n5888# 0.758287f
C78 source.t15 a_n1496_n5888# 0.758287f
C79 source.n6 a_n1496_n5888# 5.04495f
C80 source.n7 a_n1496_n5888# 0.354231f
C81 source.t13 a_n1496_n5888# 0.758287f
C82 source.t11 a_n1496_n5888# 0.758287f
C83 source.n8 a_n1496_n5888# 5.04495f
C84 source.n9 a_n1496_n5888# 2.75084f
C85 source.t0 a_n1496_n5888# 0.758287f
C86 source.t7 a_n1496_n5888# 0.758287f
C87 source.n10 a_n1496_n5888# 5.04495f
C88 source.n11 a_n1496_n5888# 2.75084f
C89 source.t5 a_n1496_n5888# 0.758287f
C90 source.t3 a_n1496_n5888# 0.758287f
C91 source.n12 a_n1496_n5888# 5.04495f
C92 source.n13 a_n1496_n5888# 0.354233f
C93 source.t6 a_n1496_n5888# 6.25299f
C94 source.n14 a_n1496_n5888# 0.526586f
C95 source.t16 a_n1496_n5888# 0.758287f
C96 source.t9 a_n1496_n5888# 0.758287f
C97 source.n15 a_n1496_n5888# 5.04495f
C98 source.n16 a_n1496_n5888# 0.369714f
C99 source.t8 a_n1496_n5888# 0.758287f
C100 source.t17 a_n1496_n5888# 0.758287f
C101 source.n17 a_n1496_n5888# 5.04495f
C102 source.n18 a_n1496_n5888# 0.354233f
C103 source.t12 a_n1496_n5888# 6.25299f
C104 source.n19 a_n1496_n5888# 0.647844f
C105 source.n20 a_n1496_n5888# 2.70144f
C106 drain_right.t5 a_n1496_n5888# 6.3902f
C107 drain_right.t6 a_n1496_n5888# 0.759307f
C108 drain_right.t9 a_n1496_n5888# 0.759307f
C109 drain_right.n0 a_n1496_n5888# 5.1349f
C110 drain_right.n1 a_n1496_n5888# 0.655983f
C111 drain_right.t7 a_n1496_n5888# 0.759307f
C112 drain_right.t0 a_n1496_n5888# 0.759307f
C113 drain_right.n2 a_n1496_n5888# 5.13676f
C114 drain_right.n3 a_n1496_n5888# 2.22759f
C115 drain_right.t4 a_n1496_n5888# 0.759307f
C116 drain_right.t8 a_n1496_n5888# 0.759307f
C117 drain_right.n4 a_n1496_n5888# 5.13787f
C118 drain_right.t1 a_n1496_n5888# 0.759307f
C119 drain_right.t3 a_n1496_n5888# 0.759307f
C120 drain_right.n5 a_n1496_n5888# 5.1349f
C121 drain_right.n6 a_n1496_n5888# 0.61929f
C122 drain_right.t2 a_n1496_n5888# 6.38664f
C123 drain_right.n7 a_n1496_n5888# 0.59816f
C124 minus.n0 a_n1496_n5888# 0.05873f
C125 minus.t4 a_n1496_n5888# 0.622071f
C126 minus.t6 a_n1496_n5888# 0.619683f
C127 minus.t7 a_n1496_n5888# 0.619683f
C128 minus.n1 a_n1496_n5888# 0.024914f
C129 minus.t2 a_n1496_n5888# 0.619683f
C130 minus.n2 a_n1496_n5888# 0.234541f
C131 minus.t3 a_n1496_n5888# 0.622071f
C132 minus.n3 a_n1496_n5888# 0.255336f
C133 minus.n4 a_n1496_n5888# 0.126434f
C134 minus.n5 a_n1496_n5888# 0.05873f
C135 minus.n6 a_n1496_n5888# 0.254024f
C136 minus.n7 a_n1496_n5888# 0.024914f
C137 minus.n8 a_n1496_n5888# 0.234541f
C138 minus.n9 a_n1496_n5888# 0.255257f
C139 minus.n10 a_n1496_n5888# 2.84383f
C140 minus.n11 a_n1496_n5888# 0.05873f
C141 minus.t0 a_n1496_n5888# 0.619683f
C142 minus.t9 a_n1496_n5888# 0.619683f
C143 minus.n12 a_n1496_n5888# 0.024914f
C144 minus.t1 a_n1496_n5888# 0.622071f
C145 minus.t8 a_n1496_n5888# 0.619683f
C146 minus.n13 a_n1496_n5888# 0.234541f
C147 minus.n14 a_n1496_n5888# 0.255336f
C148 minus.n15 a_n1496_n5888# 0.126434f
C149 minus.n16 a_n1496_n5888# 0.05873f
C150 minus.n17 a_n1496_n5888# 0.254024f
C151 minus.n18 a_n1496_n5888# 0.024914f
C152 minus.n19 a_n1496_n5888# 0.234541f
C153 minus.t5 a_n1496_n5888# 0.622071f
C154 minus.n20 a_n1496_n5888# 0.255257f
C155 minus.n21 a_n1496_n5888# 0.385867f
C156 minus.n22 a_n1496_n5888# 3.37051f
.ends

