* NGSPICE file created from diffpair236.ext - technology: sky130A

.subckt diffpair236 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t14 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X1 drain_right.t12 minus.t1 source.t23 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X2 drain_left.t13 plus.t0 source.t0 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X3 drain_left.t12 plus.t1 source.t1 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X4 drain_right.t11 minus.t2 source.t16 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X5 a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X6 drain_right.t10 minus.t3 source.t22 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X7 a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X8 drain_left.t11 plus.t2 source.t25 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X9 a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X10 drain_left.t10 plus.t3 source.t26 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X11 drain_right.t9 minus.t4 source.t15 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X12 source.t17 minus.t5 drain_right.t8 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X13 source.t18 minus.t6 drain_right.t7 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X14 source.t11 minus.t7 drain_right.t6 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X15 drain_right.t5 minus.t8 source.t19 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X16 drain_right.t4 minus.t9 source.t20 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X17 source.t21 minus.t10 drain_right.t3 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X18 source.t13 minus.t11 drain_right.t2 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 source.t27 plus.t4 drain_left.t9 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X20 source.t12 minus.t12 drain_right.t1 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X21 source.t4 plus.t5 drain_left.t8 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X22 source.t3 plus.t6 drain_left.t7 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X23 drain_right.t0 minus.t13 source.t10 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X24 drain_left.t6 plus.t7 source.t8 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X25 source.t24 plus.t8 drain_left.t5 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X26 source.t7 plus.t9 drain_left.t4 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X27 drain_left.t3 plus.t10 source.t5 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X28 drain_left.t2 plus.t11 source.t6 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X29 source.t9 plus.t12 drain_left.t1 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X30 a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X31 drain_left.t0 plus.t13 source.t2 a_n2524_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
R0 minus.n5 minus.t9 163.326
R1 minus.n23 minus.t2 163.326
R2 minus.n17 minus.n16 161.3
R3 minus.n15 minus.n0 161.3
R4 minus.n14 minus.n13 161.3
R5 minus.n12 minus.n1 161.3
R6 minus.n6 minus.n3 161.3
R7 minus.n35 minus.n34 161.3
R8 minus.n33 minus.n18 161.3
R9 minus.n32 minus.n31 161.3
R10 minus.n30 minus.n19 161.3
R11 minus.n24 minus.n21 161.3
R12 minus.n4 minus.t6 139.48
R13 minus.n8 minus.t4 139.48
R14 minus.n9 minus.t12 139.48
R15 minus.n10 minus.t13 139.48
R16 minus.n14 minus.t10 139.48
R17 minus.n16 minus.t8 139.48
R18 minus.n22 minus.t5 139.48
R19 minus.n26 minus.t3 139.48
R20 minus.n27 minus.t7 139.48
R21 minus.n28 minus.t0 139.48
R22 minus.n32 minus.t11 139.48
R23 minus.n34 minus.t1 139.48
R24 minus.n11 minus.n10 80.6037
R25 minus.n9 minus.n2 80.6037
R26 minus.n8 minus.n7 80.6037
R27 minus.n29 minus.n28 80.6037
R28 minus.n27 minus.n20 80.6037
R29 minus.n26 minus.n25 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n6 minus.n5 44.9119
R35 minus.n24 minus.n23 44.9119
R36 minus.n16 minus.n15 35.055
R37 minus.n34 minus.n33 35.055
R38 minus.n8 minus.n3 32.1338
R39 minus.n10 minus.n1 32.1338
R40 minus.n26 minus.n21 32.1338
R41 minus.n28 minus.n19 32.1338
R42 minus.n36 minus.n17 32.0895
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n4 minus.n3 16.0672
R46 minus.n14 minus.n1 16.0672
R47 minus.n22 minus.n21 16.0672
R48 minus.n32 minus.n19 16.0672
R49 minus.n15 minus.n14 13.146
R50 minus.n33 minus.n32 13.146
R51 minus.n36 minus.n35 6.72588
R52 minus.n11 minus.n2 0.380177
R53 minus.n7 minus.n2 0.380177
R54 minus.n25 minus.n20 0.380177
R55 minus.n29 minus.n20 0.380177
R56 minus.n12 minus.n11 0.285035
R57 minus.n7 minus.n6 0.285035
R58 minus.n25 minus.n24 0.285035
R59 minus.n30 minus.n29 0.285035
R60 minus.n17 minus.n0 0.189894
R61 minus.n13 minus.n0 0.189894
R62 minus.n13 minus.n12 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 source.n0 source.t8 69.6943
R68 source.n7 source.t20 69.6943
R69 source.n27 source.t23 69.6942
R70 source.n20 source.t25 69.6942
R71 source.n2 source.n1 63.0943
R72 source.n4 source.n3 63.0943
R73 source.n6 source.n5 63.0943
R74 source.n9 source.n8 63.0943
R75 source.n11 source.n10 63.0943
R76 source.n13 source.n12 63.0943
R77 source.n26 source.n25 63.0942
R78 source.n24 source.n23 63.0942
R79 source.n22 source.n21 63.0942
R80 source.n19 source.n18 63.0942
R81 source.n17 source.n16 63.0942
R82 source.n15 source.n14 63.0942
R83 source.n15 source.n13 16.4178
R84 source.n28 source.n0 9.69368
R85 source.n25 source.t14 6.6005
R86 source.n25 source.t13 6.6005
R87 source.n23 source.t22 6.6005
R88 source.n23 source.t11 6.6005
R89 source.n21 source.t16 6.6005
R90 source.n21 source.t17 6.6005
R91 source.n18 source.t26 6.6005
R92 source.n18 source.t27 6.6005
R93 source.n16 source.t0 6.6005
R94 source.n16 source.t4 6.6005
R95 source.n14 source.t1 6.6005
R96 source.n14 source.t3 6.6005
R97 source.n1 source.t6 6.6005
R98 source.n1 source.t24 6.6005
R99 source.n3 source.t5 6.6005
R100 source.n3 source.t7 6.6005
R101 source.n5 source.t2 6.6005
R102 source.n5 source.t9 6.6005
R103 source.n8 source.t15 6.6005
R104 source.n8 source.t18 6.6005
R105 source.n10 source.t10 6.6005
R106 source.n10 source.t12 6.6005
R107 source.n12 source.t19 6.6005
R108 source.n12 source.t21 6.6005
R109 source.n28 source.n27 5.7505
R110 source.n13 source.n11 0.974638
R111 source.n11 source.n9 0.974638
R112 source.n9 source.n7 0.974638
R113 source.n6 source.n4 0.974638
R114 source.n4 source.n2 0.974638
R115 source.n2 source.n0 0.974638
R116 source.n17 source.n15 0.974638
R117 source.n19 source.n17 0.974638
R118 source.n20 source.n19 0.974638
R119 source.n24 source.n22 0.974638
R120 source.n26 source.n24 0.974638
R121 source.n27 source.n26 0.974638
R122 source.n7 source.n6 0.957397
R123 source.n22 source.n20 0.957397
R124 source source.n28 0.188
R125 drain_right.n1 drain_right.t11 87.3471
R126 drain_right.n11 drain_right.t5 86.3731
R127 drain_right.n8 drain_right.n6 80.7472
R128 drain_right.n4 drain_right.n2 80.7471
R129 drain_right.n8 drain_right.n7 79.7731
R130 drain_right.n10 drain_right.n9 79.7731
R131 drain_right.n4 drain_right.n3 79.773
R132 drain_right.n1 drain_right.n0 79.773
R133 drain_right drain_right.n5 25.597
R134 drain_right.n2 drain_right.t2 6.6005
R135 drain_right.n2 drain_right.t12 6.6005
R136 drain_right.n3 drain_right.t6 6.6005
R137 drain_right.n3 drain_right.t13 6.6005
R138 drain_right.n0 drain_right.t8 6.6005
R139 drain_right.n0 drain_right.t10 6.6005
R140 drain_right.n6 drain_right.t7 6.6005
R141 drain_right.n6 drain_right.t4 6.6005
R142 drain_right.n7 drain_right.t1 6.6005
R143 drain_right.n7 drain_right.t9 6.6005
R144 drain_right.n9 drain_right.t3 6.6005
R145 drain_right.n9 drain_right.t0 6.6005
R146 drain_right drain_right.n11 6.14028
R147 drain_right.n11 drain_right.n10 0.974638
R148 drain_right.n10 drain_right.n8 0.974638
R149 drain_right.n5 drain_right.n1 0.675757
R150 drain_right.n5 drain_right.n4 0.188688
R151 plus.n5 plus.t13 163.326
R152 plus.n23 plus.t2 163.326
R153 plus.n7 plus.n6 161.3
R154 plus.n13 plus.n12 161.3
R155 plus.n14 plus.n1 161.3
R156 plus.n15 plus.n0 161.3
R157 plus.n17 plus.n16 161.3
R158 plus.n25 plus.n24 161.3
R159 plus.n31 plus.n30 161.3
R160 plus.n32 plus.n19 161.3
R161 plus.n33 plus.n18 161.3
R162 plus.n35 plus.n34 161.3
R163 plus.n16 plus.t7 139.48
R164 plus.n14 plus.t8 139.48
R165 plus.n2 plus.t11 139.48
R166 plus.n9 plus.t9 139.48
R167 plus.n8 plus.t10 139.48
R168 plus.n4 plus.t12 139.48
R169 plus.n34 plus.t1 139.48
R170 plus.n32 plus.t6 139.48
R171 plus.n20 plus.t0 139.48
R172 plus.n27 plus.t5 139.48
R173 plus.n26 plus.t3 139.48
R174 plus.n22 plus.t4 139.48
R175 plus.n8 plus.n3 80.6037
R176 plus.n10 plus.n9 80.6037
R177 plus.n11 plus.n2 80.6037
R178 plus.n26 plus.n21 80.6037
R179 plus.n28 plus.n27 80.6037
R180 plus.n29 plus.n20 80.6037
R181 plus.n9 plus.n2 48.2005
R182 plus.n9 plus.n8 48.2005
R183 plus.n27 plus.n20 48.2005
R184 plus.n27 plus.n26 48.2005
R185 plus.n24 plus.n23 44.9119
R186 plus.n6 plus.n5 44.9119
R187 plus.n16 plus.n15 35.055
R188 plus.n34 plus.n33 35.055
R189 plus.n13 plus.n2 32.1338
R190 plus.n8 plus.n7 32.1338
R191 plus.n31 plus.n20 32.1338
R192 plus.n26 plus.n25 32.1338
R193 plus plus.n35 29.3797
R194 plus.n23 plus.n22 17.739
R195 plus.n5 plus.n4 17.739
R196 plus.n14 plus.n13 16.0672
R197 plus.n7 plus.n4 16.0672
R198 plus.n32 plus.n31 16.0672
R199 plus.n25 plus.n22 16.0672
R200 plus.n15 plus.n14 13.146
R201 plus.n33 plus.n32 13.146
R202 plus plus.n17 8.96073
R203 plus.n10 plus.n3 0.380177
R204 plus.n11 plus.n10 0.380177
R205 plus.n29 plus.n28 0.380177
R206 plus.n28 plus.n21 0.380177
R207 plus.n6 plus.n3 0.285035
R208 plus.n12 plus.n11 0.285035
R209 plus.n30 plus.n29 0.285035
R210 plus.n24 plus.n21 0.285035
R211 plus.n12 plus.n1 0.189894
R212 plus.n1 plus.n0 0.189894
R213 plus.n17 plus.n0 0.189894
R214 plus.n35 plus.n18 0.189894
R215 plus.n19 plus.n18 0.189894
R216 plus.n30 plus.n19 0.189894
R217 drain_left.n7 drain_left.t0 87.3472
R218 drain_left.n1 drain_left.t12 87.3471
R219 drain_left.n4 drain_left.n2 80.7471
R220 drain_left.n11 drain_left.n10 79.7731
R221 drain_left.n9 drain_left.n8 79.7731
R222 drain_left.n7 drain_left.n6 79.7731
R223 drain_left.n4 drain_left.n3 79.773
R224 drain_left.n1 drain_left.n0 79.773
R225 drain_left drain_left.n5 26.1502
R226 drain_left drain_left.n11 6.62735
R227 drain_left.n2 drain_left.t9 6.6005
R228 drain_left.n2 drain_left.t11 6.6005
R229 drain_left.n3 drain_left.t8 6.6005
R230 drain_left.n3 drain_left.t10 6.6005
R231 drain_left.n0 drain_left.t7 6.6005
R232 drain_left.n0 drain_left.t13 6.6005
R233 drain_left.n10 drain_left.t5 6.6005
R234 drain_left.n10 drain_left.t6 6.6005
R235 drain_left.n8 drain_left.t4 6.6005
R236 drain_left.n8 drain_left.t2 6.6005
R237 drain_left.n6 drain_left.t1 6.6005
R238 drain_left.n6 drain_left.t3 6.6005
R239 drain_left.n9 drain_left.n7 0.974638
R240 drain_left.n11 drain_left.n9 0.974638
R241 drain_left.n5 drain_left.n1 0.675757
R242 drain_left.n5 drain_left.n4 0.188688
C0 plus minus 4.62663f
C1 source plus 3.37679f
C2 drain_left plus 3.0914f
C3 drain_right minus 2.84223f
C4 source drain_right 6.91818f
C5 drain_left drain_right 1.31433f
C6 source minus 3.36267f
C7 drain_left minus 0.178503f
C8 source drain_left 6.91815f
C9 drain_right plus 0.412802f
C10 drain_right a_n2524_n1488# 5.15621f
C11 drain_left a_n2524_n1488# 5.55276f
C12 source a_n2524_n1488# 3.238639f
C13 minus a_n2524_n1488# 9.280962f
C14 plus a_n2524_n1488# 10.5765f
C15 drain_left.t12 a_n2524_n1488# 0.553279f
C16 drain_left.t7 a_n2524_n1488# 0.059377f
C17 drain_left.t13 a_n2524_n1488# 0.059377f
C18 drain_left.n0 a_n2524_n1488# 0.428222f
C19 drain_left.n1 a_n2524_n1488# 0.660546f
C20 drain_left.t9 a_n2524_n1488# 0.059377f
C21 drain_left.t11 a_n2524_n1488# 0.059377f
C22 drain_left.n2 a_n2524_n1488# 0.43266f
C23 drain_left.t8 a_n2524_n1488# 0.059377f
C24 drain_left.t10 a_n2524_n1488# 0.059377f
C25 drain_left.n3 a_n2524_n1488# 0.428222f
C26 drain_left.n4 a_n2524_n1488# 0.660762f
C27 drain_left.n5 a_n2524_n1488# 0.955277f
C28 drain_left.t0 a_n2524_n1488# 0.553281f
C29 drain_left.t1 a_n2524_n1488# 0.059377f
C30 drain_left.t3 a_n2524_n1488# 0.059377f
C31 drain_left.n6 a_n2524_n1488# 0.428224f
C32 drain_left.n7 a_n2524_n1488# 0.683804f
C33 drain_left.t4 a_n2524_n1488# 0.059377f
C34 drain_left.t2 a_n2524_n1488# 0.059377f
C35 drain_left.n8 a_n2524_n1488# 0.428224f
C36 drain_left.n9 a_n2524_n1488# 0.357726f
C37 drain_left.t5 a_n2524_n1488# 0.059377f
C38 drain_left.t6 a_n2524_n1488# 0.059377f
C39 drain_left.n10 a_n2524_n1488# 0.428224f
C40 drain_left.n11 a_n2524_n1488# 0.582315f
C41 plus.n0 a_n2524_n1488# 0.042829f
C42 plus.t7 a_n2524_n1488# 0.308225f
C43 plus.t8 a_n2524_n1488# 0.308225f
C44 plus.n1 a_n2524_n1488# 0.042829f
C45 plus.t11 a_n2524_n1488# 0.308225f
C46 plus.n2 a_n2524_n1488# 0.185849f
C47 plus.n3 a_n2524_n1488# 0.071336f
C48 plus.t9 a_n2524_n1488# 0.308225f
C49 plus.t10 a_n2524_n1488# 0.308225f
C50 plus.t12 a_n2524_n1488# 0.308225f
C51 plus.n4 a_n2524_n1488# 0.180907f
C52 plus.t13 a_n2524_n1488# 0.334258f
C53 plus.n5 a_n2524_n1488# 0.155974f
C54 plus.n6 a_n2524_n1488# 0.200015f
C55 plus.n7 a_n2524_n1488# 0.009719f
C56 plus.n8 a_n2524_n1488# 0.185849f
C57 plus.n9 a_n2524_n1488# 0.188753f
C58 plus.n10 a_n2524_n1488# 0.085657f
C59 plus.n11 a_n2524_n1488# 0.071336f
C60 plus.n12 a_n2524_n1488# 0.057149f
C61 plus.n13 a_n2524_n1488# 0.009719f
C62 plus.n14 a_n2524_n1488# 0.175602f
C63 plus.n15 a_n2524_n1488# 0.009719f
C64 plus.n16 a_n2524_n1488# 0.176658f
C65 plus.n17 a_n2524_n1488# 0.343701f
C66 plus.n18 a_n2524_n1488# 0.042829f
C67 plus.t1 a_n2524_n1488# 0.308225f
C68 plus.n19 a_n2524_n1488# 0.042829f
C69 plus.t6 a_n2524_n1488# 0.308225f
C70 plus.t0 a_n2524_n1488# 0.308225f
C71 plus.n20 a_n2524_n1488# 0.185849f
C72 plus.n21 a_n2524_n1488# 0.071336f
C73 plus.t5 a_n2524_n1488# 0.308225f
C74 plus.t3 a_n2524_n1488# 0.308225f
C75 plus.t4 a_n2524_n1488# 0.308225f
C76 plus.n22 a_n2524_n1488# 0.180907f
C77 plus.t2 a_n2524_n1488# 0.334258f
C78 plus.n23 a_n2524_n1488# 0.155974f
C79 plus.n24 a_n2524_n1488# 0.200015f
C80 plus.n25 a_n2524_n1488# 0.009719f
C81 plus.n26 a_n2524_n1488# 0.185849f
C82 plus.n27 a_n2524_n1488# 0.188753f
C83 plus.n28 a_n2524_n1488# 0.085657f
C84 plus.n29 a_n2524_n1488# 0.071336f
C85 plus.n30 a_n2524_n1488# 0.057149f
C86 plus.n31 a_n2524_n1488# 0.009719f
C87 plus.n32 a_n2524_n1488# 0.175602f
C88 plus.n33 a_n2524_n1488# 0.009719f
C89 plus.n34 a_n2524_n1488# 0.176658f
C90 plus.n35 a_n2524_n1488# 1.17973f
C91 drain_right.t11 a_n2524_n1488# 0.541991f
C92 drain_right.t8 a_n2524_n1488# 0.058166f
C93 drain_right.t10 a_n2524_n1488# 0.058166f
C94 drain_right.n0 a_n2524_n1488# 0.419486f
C95 drain_right.n1 a_n2524_n1488# 0.64707f
C96 drain_right.t2 a_n2524_n1488# 0.058166f
C97 drain_right.t12 a_n2524_n1488# 0.058166f
C98 drain_right.n2 a_n2524_n1488# 0.423833f
C99 drain_right.t6 a_n2524_n1488# 0.058166f
C100 drain_right.t13 a_n2524_n1488# 0.058166f
C101 drain_right.n3 a_n2524_n1488# 0.419486f
C102 drain_right.n4 a_n2524_n1488# 0.647281f
C103 drain_right.n5 a_n2524_n1488# 0.887553f
C104 drain_right.t7 a_n2524_n1488# 0.058166f
C105 drain_right.t4 a_n2524_n1488# 0.058166f
C106 drain_right.n6 a_n2524_n1488# 0.423835f
C107 drain_right.t1 a_n2524_n1488# 0.058166f
C108 drain_right.t9 a_n2524_n1488# 0.058166f
C109 drain_right.n7 a_n2524_n1488# 0.419488f
C110 drain_right.n8 a_n2524_n1488# 0.706391f
C111 drain_right.t3 a_n2524_n1488# 0.058166f
C112 drain_right.t0 a_n2524_n1488# 0.058166f
C113 drain_right.n9 a_n2524_n1488# 0.419488f
C114 drain_right.n10 a_n2524_n1488# 0.350428f
C115 drain_right.t5 a_n2524_n1488# 0.53839f
C116 drain_right.n11 a_n2524_n1488# 0.55366f
C117 source.t8 a_n2524_n1488# 0.610206f
C118 source.n0 a_n2524_n1488# 0.908098f
C119 source.t6 a_n2524_n1488# 0.073485f
C120 source.t24 a_n2524_n1488# 0.073485f
C121 source.n1 a_n2524_n1488# 0.465936f
C122 source.n2 a_n2524_n1488# 0.46462f
C123 source.t5 a_n2524_n1488# 0.073485f
C124 source.t7 a_n2524_n1488# 0.073485f
C125 source.n3 a_n2524_n1488# 0.465936f
C126 source.n4 a_n2524_n1488# 0.46462f
C127 source.t2 a_n2524_n1488# 0.073485f
C128 source.t9 a_n2524_n1488# 0.073485f
C129 source.n5 a_n2524_n1488# 0.465936f
C130 source.n6 a_n2524_n1488# 0.462898f
C131 source.t20 a_n2524_n1488# 0.610206f
C132 source.n7 a_n2524_n1488# 0.519042f
C133 source.t15 a_n2524_n1488# 0.073485f
C134 source.t18 a_n2524_n1488# 0.073485f
C135 source.n8 a_n2524_n1488# 0.465936f
C136 source.n9 a_n2524_n1488# 0.46462f
C137 source.t10 a_n2524_n1488# 0.073485f
C138 source.t12 a_n2524_n1488# 0.073485f
C139 source.n10 a_n2524_n1488# 0.465936f
C140 source.n11 a_n2524_n1488# 0.46462f
C141 source.t19 a_n2524_n1488# 0.073485f
C142 source.t21 a_n2524_n1488# 0.073485f
C143 source.n12 a_n2524_n1488# 0.465936f
C144 source.n13 a_n2524_n1488# 1.28289f
C145 source.t1 a_n2524_n1488# 0.073485f
C146 source.t3 a_n2524_n1488# 0.073485f
C147 source.n14 a_n2524_n1488# 0.465933f
C148 source.n15 a_n2524_n1488# 1.28289f
C149 source.t0 a_n2524_n1488# 0.073485f
C150 source.t4 a_n2524_n1488# 0.073485f
C151 source.n16 a_n2524_n1488# 0.465933f
C152 source.n17 a_n2524_n1488# 0.464623f
C153 source.t26 a_n2524_n1488# 0.073485f
C154 source.t27 a_n2524_n1488# 0.073485f
C155 source.n18 a_n2524_n1488# 0.465933f
C156 source.n19 a_n2524_n1488# 0.464623f
C157 source.t25 a_n2524_n1488# 0.610202f
C158 source.n20 a_n2524_n1488# 0.519045f
C159 source.t16 a_n2524_n1488# 0.073485f
C160 source.t17 a_n2524_n1488# 0.073485f
C161 source.n21 a_n2524_n1488# 0.465933f
C162 source.n22 a_n2524_n1488# 0.462901f
C163 source.t22 a_n2524_n1488# 0.073485f
C164 source.t11 a_n2524_n1488# 0.073485f
C165 source.n23 a_n2524_n1488# 0.465933f
C166 source.n24 a_n2524_n1488# 0.464623f
C167 source.t14 a_n2524_n1488# 0.073485f
C168 source.t13 a_n2524_n1488# 0.073485f
C169 source.n25 a_n2524_n1488# 0.465933f
C170 source.n26 a_n2524_n1488# 0.464623f
C171 source.t23 a_n2524_n1488# 0.610202f
C172 source.n27 a_n2524_n1488# 0.679304f
C173 source.n28 a_n2524_n1488# 0.918115f
C174 minus.n0 a_n2524_n1488# 0.041348f
C175 minus.n1 a_n2524_n1488# 0.009383f
C176 minus.t10 a_n2524_n1488# 0.297573f
C177 minus.n2 a_n2524_n1488# 0.082697f
C178 minus.n3 a_n2524_n1488# 0.009383f
C179 minus.t4 a_n2524_n1488# 0.297573f
C180 minus.t9 a_n2524_n1488# 0.322706f
C181 minus.t6 a_n2524_n1488# 0.297573f
C182 minus.n4 a_n2524_n1488# 0.174655f
C183 minus.n5 a_n2524_n1488# 0.150583f
C184 minus.n6 a_n2524_n1488# 0.193102f
C185 minus.n7 a_n2524_n1488# 0.068871f
C186 minus.n8 a_n2524_n1488# 0.179426f
C187 minus.t12 a_n2524_n1488# 0.297573f
C188 minus.n9 a_n2524_n1488# 0.18223f
C189 minus.t13 a_n2524_n1488# 0.297573f
C190 minus.n10 a_n2524_n1488# 0.179426f
C191 minus.n11 a_n2524_n1488# 0.068871f
C192 minus.n12 a_n2524_n1488# 0.055174f
C193 minus.n13 a_n2524_n1488# 0.041348f
C194 minus.n14 a_n2524_n1488# 0.169533f
C195 minus.n15 a_n2524_n1488# 0.009383f
C196 minus.t8 a_n2524_n1488# 0.297573f
C197 minus.n16 a_n2524_n1488# 0.170553f
C198 minus.n17 a_n2524_n1488# 1.21252f
C199 minus.n18 a_n2524_n1488# 0.041348f
C200 minus.n19 a_n2524_n1488# 0.009383f
C201 minus.n20 a_n2524_n1488# 0.082697f
C202 minus.n21 a_n2524_n1488# 0.009383f
C203 minus.t2 a_n2524_n1488# 0.322706f
C204 minus.t5 a_n2524_n1488# 0.297573f
C205 minus.n22 a_n2524_n1488# 0.174655f
C206 minus.n23 a_n2524_n1488# 0.150583f
C207 minus.n24 a_n2524_n1488# 0.193102f
C208 minus.n25 a_n2524_n1488# 0.068871f
C209 minus.t3 a_n2524_n1488# 0.297573f
C210 minus.n26 a_n2524_n1488# 0.179426f
C211 minus.t7 a_n2524_n1488# 0.297573f
C212 minus.n27 a_n2524_n1488# 0.18223f
C213 minus.t0 a_n2524_n1488# 0.297573f
C214 minus.n28 a_n2524_n1488# 0.179426f
C215 minus.n29 a_n2524_n1488# 0.068871f
C216 minus.n30 a_n2524_n1488# 0.055174f
C217 minus.n31 a_n2524_n1488# 0.041348f
C218 minus.t11 a_n2524_n1488# 0.297573f
C219 minus.n32 a_n2524_n1488# 0.169533f
C220 minus.n33 a_n2524_n1488# 0.009383f
C221 minus.t1 a_n2524_n1488# 0.297573f
C222 minus.n34 a_n2524_n1488# 0.170553f
C223 minus.n35 a_n2524_n1488# 0.2921f
C224 minus.n36 a_n2524_n1488# 1.48001f
.ends

