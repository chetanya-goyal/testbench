* NGSPICE file created from diffpair525.ext - technology: sky130A

.subckt diffpair525 minus drain_right drain_left source plus
X0 a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X1 source.t20 plus.t0 drain_left.t6 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X2 drain_left.t9 plus.t1 source.t19 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X3 source.t2 minus.t0 drain_right.t11 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X4 source.t18 plus.t2 drain_left.t5 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X5 source.t17 plus.t3 drain_left.t10 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X6 drain_left.t2 plus.t4 source.t16 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X7 drain_right.t10 minus.t1 source.t7 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X8 drain_right.t9 minus.t2 source.t1 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X9 source.t5 minus.t3 drain_right.t8 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X10 drain_right.t7 minus.t4 source.t6 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X11 a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X12 drain_left.t8 plus.t5 source.t15 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X13 source.t22 minus.t5 drain_right.t6 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X14 drain_left.t11 plus.t6 source.t14 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 source.t8 minus.t6 drain_right.t5 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X16 a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X17 source.t13 plus.t7 drain_left.t0 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X18 drain_right.t4 minus.t7 source.t0 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X19 drain_right.t3 minus.t8 source.t23 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X20 source.t4 minus.t9 drain_right.t2 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X21 drain_left.t7 plus.t8 source.t12 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X22 a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X23 source.t3 minus.t10 drain_right.t1 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X24 drain_right.t0 minus.t11 source.t21 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X25 source.t11 plus.t9 drain_left.t4 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X26 source.t10 plus.t10 drain_left.t3 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X27 drain_left.t1 plus.t11 source.t9 a_n1878_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
R0 plus.n5 plus.t2 828.236
R1 plus.n19 plus.t1 828.236
R2 plus.n12 plus.t11 801.567
R3 plus.n10 plus.t9 801.567
R4 plus.n9 plus.t5 801.567
R5 plus.n3 plus.t10 801.567
R6 plus.n4 plus.t8 801.567
R7 plus.n26 plus.t7 801.567
R8 plus.n24 plus.t4 801.567
R9 plus.n23 plus.t3 801.567
R10 plus.n17 plus.t6 801.567
R11 plus.n18 plus.t0 801.567
R12 plus.n6 plus.n3 161.3
R13 plus.n8 plus.n7 161.3
R14 plus.n9 plus.n2 161.3
R15 plus.n10 plus.n1 161.3
R16 plus.n11 plus.n0 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n20 plus.n17 161.3
R19 plus.n22 plus.n21 161.3
R20 plus.n23 plus.n16 161.3
R21 plus.n24 plus.n15 161.3
R22 plus.n25 plus.n14 161.3
R23 plus.n27 plus.n26 161.3
R24 plus.n10 plus.n9 48.2005
R25 plus.n4 plus.n3 48.2005
R26 plus.n24 plus.n23 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n12 plus.n11 47.4702
R29 plus.n26 plus.n25 47.4702
R30 plus.n6 plus.n5 45.1192
R31 plus.n20 plus.n19 45.1192
R32 plus plus.n27 31.2831
R33 plus.n8 plus.n3 24.1005
R34 plus.n9 plus.n8 24.1005
R35 plus.n23 plus.n22 24.1005
R36 plus.n22 plus.n17 24.1005
R37 plus.n5 plus.n4 13.6377
R38 plus.n19 plus.n18 13.6377
R39 plus plus.n13 13.3111
R40 plus.n11 plus.n10 0.730803
R41 plus.n25 plus.n24 0.730803
R42 plus.n7 plus.n6 0.189894
R43 plus.n7 plus.n2 0.189894
R44 plus.n2 plus.n1 0.189894
R45 plus.n1 plus.n0 0.189894
R46 plus.n13 plus.n0 0.189894
R47 plus.n27 plus.n14 0.189894
R48 plus.n15 plus.n14 0.189894
R49 plus.n16 plus.n15 0.189894
R50 plus.n21 plus.n16 0.189894
R51 plus.n21 plus.n20 0.189894
R52 drain_left.n6 drain_left.n4 61.5953
R53 drain_left.n3 drain_left.n2 61.5397
R54 drain_left.n3 drain_left.n0 61.5397
R55 drain_left.n6 drain_left.n5 60.8798
R56 drain_left.n8 drain_left.n7 60.8796
R57 drain_left.n3 drain_left.n1 60.8796
R58 drain_left drain_left.n3 33.2174
R59 drain_left drain_left.n8 6.36873
R60 drain_left.n1 drain_left.t10 1.3205
R61 drain_left.n1 drain_left.t11 1.3205
R62 drain_left.n2 drain_left.t6 1.3205
R63 drain_left.n2 drain_left.t9 1.3205
R64 drain_left.n0 drain_left.t0 1.3205
R65 drain_left.n0 drain_left.t2 1.3205
R66 drain_left.n7 drain_left.t4 1.3205
R67 drain_left.n7 drain_left.t1 1.3205
R68 drain_left.n5 drain_left.t3 1.3205
R69 drain_left.n5 drain_left.t8 1.3205
R70 drain_left.n4 drain_left.t5 1.3205
R71 drain_left.n4 drain_left.t7 1.3205
R72 drain_left.n8 drain_left.n6 0.716017
R73 source.n5 source.t18 45.521
R74 source.n6 source.t0 45.521
R75 source.n11 source.t8 45.521
R76 source.n23 source.t21 45.5208
R77 source.n18 source.t5 45.5208
R78 source.n17 source.t19 45.5208
R79 source.n12 source.t13 45.5208
R80 source.n0 source.t9 45.5208
R81 source.n2 source.n1 44.201
R82 source.n4 source.n3 44.201
R83 source.n8 source.n7 44.201
R84 source.n10 source.n9 44.201
R85 source.n22 source.n21 44.2008
R86 source.n20 source.n19 44.2008
R87 source.n16 source.n15 44.2008
R88 source.n14 source.n13 44.2008
R89 source.n12 source.n11 24.276
R90 source.n24 source.n0 18.6553
R91 source.n24 source.n23 5.62119
R92 source.n21 source.t23 1.3205
R93 source.n21 source.t22 1.3205
R94 source.n19 source.t1 1.3205
R95 source.n19 source.t4 1.3205
R96 source.n15 source.t14 1.3205
R97 source.n15 source.t20 1.3205
R98 source.n13 source.t16 1.3205
R99 source.n13 source.t17 1.3205
R100 source.n1 source.t15 1.3205
R101 source.n1 source.t11 1.3205
R102 source.n3 source.t12 1.3205
R103 source.n3 source.t10 1.3205
R104 source.n7 source.t6 1.3205
R105 source.n7 source.t2 1.3205
R106 source.n9 source.t7 1.3205
R107 source.n9 source.t3 1.3205
R108 source.n11 source.n10 0.716017
R109 source.n10 source.n8 0.716017
R110 source.n8 source.n6 0.716017
R111 source.n5 source.n4 0.716017
R112 source.n4 source.n2 0.716017
R113 source.n2 source.n0 0.716017
R114 source.n14 source.n12 0.716017
R115 source.n16 source.n14 0.716017
R116 source.n17 source.n16 0.716017
R117 source.n20 source.n18 0.716017
R118 source.n22 source.n20 0.716017
R119 source.n23 source.n22 0.716017
R120 source.n6 source.n5 0.470328
R121 source.n18 source.n17 0.470328
R122 source source.n24 0.188
R123 minus.n3 minus.t7 828.236
R124 minus.n17 minus.t3 828.236
R125 minus.n4 minus.t0 801.567
R126 minus.n5 minus.t4 801.567
R127 minus.n1 minus.t10 801.567
R128 minus.n10 minus.t1 801.567
R129 minus.n12 minus.t6 801.567
R130 minus.n18 minus.t2 801.567
R131 minus.n19 minus.t9 801.567
R132 minus.n15 minus.t8 801.567
R133 minus.n24 minus.t5 801.567
R134 minus.n26 minus.t11 801.567
R135 minus.n13 minus.n12 161.3
R136 minus.n11 minus.n0 161.3
R137 minus.n10 minus.n9 161.3
R138 minus.n8 minus.n1 161.3
R139 minus.n7 minus.n6 161.3
R140 minus.n5 minus.n2 161.3
R141 minus.n27 minus.n26 161.3
R142 minus.n25 minus.n14 161.3
R143 minus.n24 minus.n23 161.3
R144 minus.n22 minus.n15 161.3
R145 minus.n21 minus.n20 161.3
R146 minus.n19 minus.n16 161.3
R147 minus.n5 minus.n4 48.2005
R148 minus.n10 minus.n1 48.2005
R149 minus.n19 minus.n18 48.2005
R150 minus.n24 minus.n15 48.2005
R151 minus.n12 minus.n11 47.4702
R152 minus.n26 minus.n25 47.4702
R153 minus.n3 minus.n2 45.1192
R154 minus.n17 minus.n16 45.1192
R155 minus.n28 minus.n13 38.5384
R156 minus.n6 minus.n1 24.1005
R157 minus.n6 minus.n5 24.1005
R158 minus.n20 minus.n19 24.1005
R159 minus.n20 minus.n15 24.1005
R160 minus.n4 minus.n3 13.6377
R161 minus.n18 minus.n17 13.6377
R162 minus.n28 minus.n27 6.5308
R163 minus.n11 minus.n10 0.730803
R164 minus.n25 minus.n24 0.730803
R165 minus.n13 minus.n0 0.189894
R166 minus.n9 minus.n0 0.189894
R167 minus.n9 minus.n8 0.189894
R168 minus.n8 minus.n7 0.189894
R169 minus.n7 minus.n2 0.189894
R170 minus.n21 minus.n16 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n14 0.189894
R174 minus.n27 minus.n14 0.189894
R175 minus minus.n28 0.188
R176 drain_right.n6 drain_right.n4 61.5952
R177 drain_right.n3 drain_right.n2 61.5397
R178 drain_right.n3 drain_right.n0 61.5397
R179 drain_right.n6 drain_right.n5 60.8798
R180 drain_right.n8 drain_right.n7 60.8798
R181 drain_right.n3 drain_right.n1 60.8796
R182 drain_right drain_right.n3 32.6642
R183 drain_right drain_right.n8 6.36873
R184 drain_right.n1 drain_right.t2 1.3205
R185 drain_right.n1 drain_right.t3 1.3205
R186 drain_right.n2 drain_right.t6 1.3205
R187 drain_right.n2 drain_right.t0 1.3205
R188 drain_right.n0 drain_right.t8 1.3205
R189 drain_right.n0 drain_right.t9 1.3205
R190 drain_right.n4 drain_right.t11 1.3205
R191 drain_right.n4 drain_right.t4 1.3205
R192 drain_right.n5 drain_right.t1 1.3205
R193 drain_right.n5 drain_right.t7 1.3205
R194 drain_right.n7 drain_right.t5 1.3205
R195 drain_right.n7 drain_right.t10 1.3205
R196 drain_right.n8 drain_right.n6 0.716017
C0 drain_left plus 8.165359f
C1 source plus 7.64631f
C2 drain_right minus 7.982759f
C3 drain_right drain_left 0.936346f
C4 drain_right source 22.242699f
C5 minus drain_left 0.171641f
C6 minus source 7.63227f
C7 drain_right plus 0.337327f
C8 minus plus 6.04879f
C9 source drain_left 22.2417f
C10 drain_right a_n1878_n3888# 6.67138f
C11 drain_left a_n1878_n3888# 6.953031f
C12 source a_n1878_n3888# 10.544842f
C13 minus a_n1878_n3888# 7.563513f
C14 plus a_n1878_n3888# 9.55871f
C15 drain_right.t8 a_n1878_n3888# 0.346507f
C16 drain_right.t9 a_n1878_n3888# 0.346507f
C17 drain_right.n0 a_n1878_n3888# 3.13611f
C18 drain_right.t2 a_n1878_n3888# 0.346507f
C19 drain_right.t3 a_n1878_n3888# 0.346507f
C20 drain_right.n1 a_n1878_n3888# 3.13202f
C21 drain_right.t6 a_n1878_n3888# 0.346507f
C22 drain_right.t0 a_n1878_n3888# 0.346507f
C23 drain_right.n2 a_n1878_n3888# 3.13611f
C24 drain_right.n3 a_n1878_n3888# 2.6676f
C25 drain_right.t11 a_n1878_n3888# 0.346507f
C26 drain_right.t4 a_n1878_n3888# 0.346507f
C27 drain_right.n4 a_n1878_n3888# 3.13649f
C28 drain_right.t1 a_n1878_n3888# 0.346507f
C29 drain_right.t7 a_n1878_n3888# 0.346507f
C30 drain_right.n5 a_n1878_n3888# 3.13202f
C31 drain_right.n6 a_n1878_n3888# 0.75575f
C32 drain_right.t5 a_n1878_n3888# 0.346507f
C33 drain_right.t10 a_n1878_n3888# 0.346507f
C34 drain_right.n7 a_n1878_n3888# 3.13202f
C35 drain_right.n8 a_n1878_n3888# 0.625373f
C36 minus.n0 a_n1878_n3888# 0.046299f
C37 minus.t10 a_n1878_n3888# 0.986752f
C38 minus.n1 a_n1878_n3888# 0.389113f
C39 minus.t1 a_n1878_n3888# 0.986752f
C40 minus.n2 a_n1878_n3888# 0.188557f
C41 minus.t7 a_n1878_n3888# 0.999131f
C42 minus.n3 a_n1878_n3888# 0.373159f
C43 minus.t0 a_n1878_n3888# 0.986752f
C44 minus.n4 a_n1878_n3888# 0.394694f
C45 minus.t4 a_n1878_n3888# 0.986752f
C46 minus.n5 a_n1878_n3888# 0.389113f
C47 minus.n6 a_n1878_n3888# 0.010506f
C48 minus.n7 a_n1878_n3888# 0.046299f
C49 minus.n8 a_n1878_n3888# 0.046299f
C50 minus.n9 a_n1878_n3888# 0.046299f
C51 minus.n10 a_n1878_n3888# 0.384546f
C52 minus.n11 a_n1878_n3888# 0.010506f
C53 minus.t6 a_n1878_n3888# 0.986752f
C54 minus.n12 a_n1878_n3888# 0.384261f
C55 minus.n13 a_n1878_n3888# 1.80367f
C56 minus.n14 a_n1878_n3888# 0.046299f
C57 minus.t8 a_n1878_n3888# 0.986752f
C58 minus.n15 a_n1878_n3888# 0.389113f
C59 minus.n16 a_n1878_n3888# 0.188557f
C60 minus.t3 a_n1878_n3888# 0.999131f
C61 minus.n17 a_n1878_n3888# 0.373159f
C62 minus.t2 a_n1878_n3888# 0.986752f
C63 minus.n18 a_n1878_n3888# 0.394694f
C64 minus.t9 a_n1878_n3888# 0.986752f
C65 minus.n19 a_n1878_n3888# 0.389113f
C66 minus.n20 a_n1878_n3888# 0.010506f
C67 minus.n21 a_n1878_n3888# 0.046299f
C68 minus.n22 a_n1878_n3888# 0.046299f
C69 minus.n23 a_n1878_n3888# 0.046299f
C70 minus.t5 a_n1878_n3888# 0.986752f
C71 minus.n24 a_n1878_n3888# 0.384546f
C72 minus.n25 a_n1878_n3888# 0.010506f
C73 minus.t11 a_n1878_n3888# 0.986752f
C74 minus.n26 a_n1878_n3888# 0.384261f
C75 minus.n27 a_n1878_n3888# 0.306043f
C76 minus.n28 a_n1878_n3888# 2.1748f
C77 source.t9 a_n1878_n3888# 3.05726f
C78 source.n0 a_n1878_n3888# 1.43668f
C79 source.t15 a_n1878_n3888# 0.272808f
C80 source.t11 a_n1878_n3888# 0.272808f
C81 source.n1 a_n1878_n3888# 2.39639f
C82 source.n2 a_n1878_n3888# 0.332826f
C83 source.t12 a_n1878_n3888# 0.272808f
C84 source.t10 a_n1878_n3888# 0.272808f
C85 source.n3 a_n1878_n3888# 2.39639f
C86 source.n4 a_n1878_n3888# 0.332826f
C87 source.t18 a_n1878_n3888# 3.05726f
C88 source.n5 a_n1878_n3888# 0.397761f
C89 source.t0 a_n1878_n3888# 3.05726f
C90 source.n6 a_n1878_n3888# 0.397761f
C91 source.t6 a_n1878_n3888# 0.272808f
C92 source.t2 a_n1878_n3888# 0.272808f
C93 source.n7 a_n1878_n3888# 2.39639f
C94 source.n8 a_n1878_n3888# 0.332826f
C95 source.t7 a_n1878_n3888# 0.272808f
C96 source.t3 a_n1878_n3888# 0.272808f
C97 source.n9 a_n1878_n3888# 2.39639f
C98 source.n10 a_n1878_n3888# 0.332826f
C99 source.t8 a_n1878_n3888# 3.05726f
C100 source.n11 a_n1878_n3888# 1.82428f
C101 source.t13 a_n1878_n3888# 3.05726f
C102 source.n12 a_n1878_n3888# 1.82428f
C103 source.t16 a_n1878_n3888# 0.272808f
C104 source.t17 a_n1878_n3888# 0.272808f
C105 source.n13 a_n1878_n3888# 2.39639f
C106 source.n14 a_n1878_n3888# 0.33283f
C107 source.t14 a_n1878_n3888# 0.272808f
C108 source.t20 a_n1878_n3888# 0.272808f
C109 source.n15 a_n1878_n3888# 2.39639f
C110 source.n16 a_n1878_n3888# 0.33283f
C111 source.t19 a_n1878_n3888# 3.05726f
C112 source.n17 a_n1878_n3888# 0.397764f
C113 source.t5 a_n1878_n3888# 3.05726f
C114 source.n18 a_n1878_n3888# 0.397764f
C115 source.t1 a_n1878_n3888# 0.272808f
C116 source.t4 a_n1878_n3888# 0.272808f
C117 source.n19 a_n1878_n3888# 2.39639f
C118 source.n20 a_n1878_n3888# 0.33283f
C119 source.t23 a_n1878_n3888# 0.272808f
C120 source.t22 a_n1878_n3888# 0.272808f
C121 source.n21 a_n1878_n3888# 2.39639f
C122 source.n22 a_n1878_n3888# 0.33283f
C123 source.t21 a_n1878_n3888# 3.05726f
C124 source.n23 a_n1878_n3888# 0.537845f
C125 source.n24 a_n1878_n3888# 1.69041f
C126 drain_left.t0 a_n1878_n3888# 0.347486f
C127 drain_left.t2 a_n1878_n3888# 0.347486f
C128 drain_left.n0 a_n1878_n3888# 3.14497f
C129 drain_left.t10 a_n1878_n3888# 0.347486f
C130 drain_left.t11 a_n1878_n3888# 0.347486f
C131 drain_left.n1 a_n1878_n3888# 3.14087f
C132 drain_left.t6 a_n1878_n3888# 0.347486f
C133 drain_left.t9 a_n1878_n3888# 0.347486f
C134 drain_left.n2 a_n1878_n3888# 3.14497f
C135 drain_left.n3 a_n1878_n3888# 2.73612f
C136 drain_left.t5 a_n1878_n3888# 0.347486f
C137 drain_left.t7 a_n1878_n3888# 0.347486f
C138 drain_left.n4 a_n1878_n3888# 3.14536f
C139 drain_left.t3 a_n1878_n3888# 0.347486f
C140 drain_left.t8 a_n1878_n3888# 0.347486f
C141 drain_left.n5 a_n1878_n3888# 3.14087f
C142 drain_left.n6 a_n1878_n3888# 0.757875f
C143 drain_left.t4 a_n1878_n3888# 0.347486f
C144 drain_left.t1 a_n1878_n3888# 0.347486f
C145 drain_left.n7 a_n1878_n3888# 3.14086f
C146 drain_left.n8 a_n1878_n3888# 0.627151f
C147 plus.n0 a_n1878_n3888# 0.046931f
C148 plus.t11 a_n1878_n3888# 1.00022f
C149 plus.t9 a_n1878_n3888# 1.00022f
C150 plus.n1 a_n1878_n3888# 0.046931f
C151 plus.t5 a_n1878_n3888# 1.00022f
C152 plus.n2 a_n1878_n3888# 0.046931f
C153 plus.t10 a_n1878_n3888# 1.00022f
C154 plus.n3 a_n1878_n3888# 0.394426f
C155 plus.t8 a_n1878_n3888# 1.00022f
C156 plus.n4 a_n1878_n3888# 0.400083f
C157 plus.t2 a_n1878_n3888# 1.01277f
C158 plus.n5 a_n1878_n3888# 0.378253f
C159 plus.n6 a_n1878_n3888# 0.191132f
C160 plus.n7 a_n1878_n3888# 0.046931f
C161 plus.n8 a_n1878_n3888# 0.01065f
C162 plus.n9 a_n1878_n3888# 0.394426f
C163 plus.n10 a_n1878_n3888# 0.389796f
C164 plus.n11 a_n1878_n3888# 0.01065f
C165 plus.n12 a_n1878_n3888# 0.389507f
C166 plus.n13 a_n1878_n3888# 0.596459f
C167 plus.n14 a_n1878_n3888# 0.046931f
C168 plus.t7 a_n1878_n3888# 1.00022f
C169 plus.n15 a_n1878_n3888# 0.046931f
C170 plus.t4 a_n1878_n3888# 1.00022f
C171 plus.n16 a_n1878_n3888# 0.046931f
C172 plus.t3 a_n1878_n3888# 1.00022f
C173 plus.t6 a_n1878_n3888# 1.00022f
C174 plus.n17 a_n1878_n3888# 0.394426f
C175 plus.t1 a_n1878_n3888# 1.01277f
C176 plus.t0 a_n1878_n3888# 1.00022f
C177 plus.n18 a_n1878_n3888# 0.400083f
C178 plus.n19 a_n1878_n3888# 0.378253f
C179 plus.n20 a_n1878_n3888# 0.191132f
C180 plus.n21 a_n1878_n3888# 0.046931f
C181 plus.n22 a_n1878_n3888# 0.01065f
C182 plus.n23 a_n1878_n3888# 0.394426f
C183 plus.n24 a_n1878_n3888# 0.389796f
C184 plus.n25 a_n1878_n3888# 0.01065f
C185 plus.n26 a_n1878_n3888# 0.389507f
C186 plus.n27 a_n1878_n3888# 1.50529f
.ends

