* NGSPICE file created from diffpair531.ext - technology: sky130A

.subckt diffpair531 minus drain_right drain_left source plus
X0 a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.6
X1 drain_left plus source a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X2 a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X3 drain_right minus source a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X4 a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X5 source plus drain_left a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X6 source minus drain_right a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X7 drain_right minus source a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X8 drain_left plus source a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X9 source plus drain_left a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X10 source minus drain_right a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X11 a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# a_n1274_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
.ends

