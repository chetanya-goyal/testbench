* NGSPICE file created from diffpair155.ext - technology: sky130A

.subckt diffpair155 minus drain_right drain_left source plus
X0 a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X1 drain_right.t11 minus.t0 source.t13 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X2 drain_right.t10 minus.t1 source.t12 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 drain_right.t9 minus.t2 source.t14 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X4 a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X5 source.t4 plus.t0 drain_left.t11 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X6 source.t1 plus.t1 drain_left.t10 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X7 source.t3 plus.t2 drain_left.t9 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X8 a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X9 drain_right.t8 minus.t3 source.t19 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X10 source.t22 minus.t4 drain_right.t7 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X11 drain_right.t6 minus.t5 source.t17 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X12 source.t15 minus.t6 drain_right.t5 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X13 source.t16 minus.t7 drain_right.t4 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X14 drain_left.t8 plus.t3 source.t8 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X15 source.t18 minus.t8 drain_right.t3 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X16 drain_right.t2 minus.t9 source.t21 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X17 drain_left.t7 plus.t4 source.t9 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X18 drain_left.t6 plus.t5 source.t5 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X19 source.t23 minus.t10 drain_right.t1 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X20 source.t7 plus.t6 drain_left.t5 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X21 source.t20 minus.t11 drain_right.t0 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X22 source.t2 plus.t7 drain_left.t4 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X23 drain_left.t3 plus.t8 source.t10 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X24 a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X25 drain_left.t2 plus.t9 source.t11 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X26 source.t6 plus.t10 drain_left.t1 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X27 drain_left.t0 plus.t11 source.t0 a_n2298_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n15 minus.n14 161.3
R1 minus.n13 minus.n0 161.3
R2 minus.n12 minus.n11 161.3
R3 minus.n10 minus.n1 161.3
R4 minus.n6 minus.n5 161.3
R5 minus.n31 minus.n30 161.3
R6 minus.n29 minus.n16 161.3
R7 minus.n28 minus.n27 161.3
R8 minus.n26 minus.n17 161.3
R9 minus.n22 minus.n21 161.3
R10 minus.n4 minus.t5 130.75
R11 minus.n20 minus.t10 130.75
R12 minus.n3 minus.t4 109.355
R13 minus.n7 minus.t3 109.355
R14 minus.n8 minus.t8 109.355
R15 minus.n12 minus.t9 109.355
R16 minus.n14 minus.t7 109.355
R17 minus.n19 minus.t0 109.355
R18 minus.n23 minus.t11 109.355
R19 minus.n24 minus.t1 109.355
R20 minus.n28 minus.t6 109.355
R21 minus.n30 minus.t2 109.355
R22 minus.n9 minus.n8 80.6037
R23 minus.n7 minus.n2 80.6037
R24 minus.n25 minus.n24 80.6037
R25 minus.n23 minus.n18 80.6037
R26 minus.n8 minus.n7 48.2005
R27 minus.n24 minus.n23 48.2005
R28 minus.n5 minus.n4 44.853
R29 minus.n21 minus.n20 44.853
R30 minus.n7 minus.n6 41.6278
R31 minus.n8 minus.n1 41.6278
R32 minus.n23 minus.n22 41.6278
R33 minus.n24 minus.n17 41.6278
R34 minus.n32 minus.n15 30.4513
R35 minus.n14 minus.n13 25.5611
R36 minus.n30 minus.n29 25.5611
R37 minus.n13 minus.n12 22.6399
R38 minus.n29 minus.n28 22.6399
R39 minus.n4 minus.n3 20.5405
R40 minus.n20 minus.n19 20.5405
R41 minus.n32 minus.n31 6.70126
R42 minus.n6 minus.n3 6.57323
R43 minus.n12 minus.n1 6.57323
R44 minus.n22 minus.n19 6.57323
R45 minus.n28 minus.n17 6.57323
R46 minus.n9 minus.n2 0.380177
R47 minus.n25 minus.n18 0.380177
R48 minus.n10 minus.n9 0.285035
R49 minus.n5 minus.n2 0.285035
R50 minus.n21 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n27 minus.n26 0.189894
R56 minus.n27 minus.n16 0.189894
R57 minus.n31 minus.n16 0.189894
R58 minus minus.n32 0.188
R59 source.n74 source.n72 289.615
R60 source.n62 source.n60 289.615
R61 source.n54 source.n52 289.615
R62 source.n42 source.n40 289.615
R63 source.n2 source.n0 289.615
R64 source.n14 source.n12 289.615
R65 source.n22 source.n20 289.615
R66 source.n34 source.n32 289.615
R67 source.n75 source.n74 185
R68 source.n63 source.n62 185
R69 source.n55 source.n54 185
R70 source.n43 source.n42 185
R71 source.n3 source.n2 185
R72 source.n15 source.n14 185
R73 source.n23 source.n22 185
R74 source.n35 source.n34 185
R75 source.t14 source.n73 167.117
R76 source.t23 source.n61 167.117
R77 source.t11 source.n53 167.117
R78 source.t3 source.n41 167.117
R79 source.t9 source.n1 167.117
R80 source.t6 source.n13 167.117
R81 source.t17 source.n21 167.117
R82 source.t16 source.n33 167.117
R83 source.n9 source.n8 84.1169
R84 source.n11 source.n10 84.1169
R85 source.n29 source.n28 84.1169
R86 source.n31 source.n30 84.1169
R87 source.n71 source.n70 84.1168
R88 source.n69 source.n68 84.1168
R89 source.n51 source.n50 84.1168
R90 source.n49 source.n48 84.1168
R91 source.n74 source.t14 52.3082
R92 source.n62 source.t23 52.3082
R93 source.n54 source.t11 52.3082
R94 source.n42 source.t3 52.3082
R95 source.n2 source.t9 52.3082
R96 source.n14 source.t6 52.3082
R97 source.n22 source.t17 52.3082
R98 source.n34 source.t16 52.3082
R99 source.n79 source.n78 31.4096
R100 source.n67 source.n66 31.4096
R101 source.n59 source.n58 31.4096
R102 source.n47 source.n46 31.4096
R103 source.n7 source.n6 31.4096
R104 source.n19 source.n18 31.4096
R105 source.n27 source.n26 31.4096
R106 source.n39 source.n38 31.4096
R107 source.n47 source.n39 14.6861
R108 source.n70 source.t12 9.9005
R109 source.n70 source.t15 9.9005
R110 source.n68 source.t13 9.9005
R111 source.n68 source.t20 9.9005
R112 source.n50 source.t0 9.9005
R113 source.n50 source.t4 9.9005
R114 source.n48 source.t8 9.9005
R115 source.n48 source.t1 9.9005
R116 source.n8 source.t5 9.9005
R117 source.n8 source.t2 9.9005
R118 source.n10 source.t10 9.9005
R119 source.n10 source.t7 9.9005
R120 source.n28 source.t19 9.9005
R121 source.n28 source.t22 9.9005
R122 source.n30 source.t21 9.9005
R123 source.n30 source.t18 9.9005
R124 source.n75 source.n73 9.71174
R125 source.n63 source.n61 9.71174
R126 source.n55 source.n53 9.71174
R127 source.n43 source.n41 9.71174
R128 source.n3 source.n1 9.71174
R129 source.n15 source.n13 9.71174
R130 source.n23 source.n21 9.71174
R131 source.n35 source.n33 9.71174
R132 source.n78 source.n77 9.45567
R133 source.n66 source.n65 9.45567
R134 source.n58 source.n57 9.45567
R135 source.n46 source.n45 9.45567
R136 source.n6 source.n5 9.45567
R137 source.n18 source.n17 9.45567
R138 source.n26 source.n25 9.45567
R139 source.n38 source.n37 9.45567
R140 source.n77 source.n76 9.3005
R141 source.n65 source.n64 9.3005
R142 source.n57 source.n56 9.3005
R143 source.n45 source.n44 9.3005
R144 source.n5 source.n4 9.3005
R145 source.n17 source.n16 9.3005
R146 source.n25 source.n24 9.3005
R147 source.n37 source.n36 9.3005
R148 source.n80 source.n7 8.93611
R149 source.n78 source.n72 8.14595
R150 source.n66 source.n60 8.14595
R151 source.n58 source.n52 8.14595
R152 source.n46 source.n40 8.14595
R153 source.n6 source.n0 8.14595
R154 source.n18 source.n12 8.14595
R155 source.n26 source.n20 8.14595
R156 source.n38 source.n32 8.14595
R157 source.n76 source.n75 7.3702
R158 source.n64 source.n63 7.3702
R159 source.n56 source.n55 7.3702
R160 source.n44 source.n43 7.3702
R161 source.n4 source.n3 7.3702
R162 source.n16 source.n15 7.3702
R163 source.n24 source.n23 7.3702
R164 source.n36 source.n35 7.3702
R165 source.n76 source.n72 5.81868
R166 source.n64 source.n60 5.81868
R167 source.n56 source.n52 5.81868
R168 source.n44 source.n40 5.81868
R169 source.n4 source.n0 5.81868
R170 source.n16 source.n12 5.81868
R171 source.n24 source.n20 5.81868
R172 source.n36 source.n32 5.81868
R173 source.n80 source.n79 5.7505
R174 source.n77 source.n73 3.44771
R175 source.n65 source.n61 3.44771
R176 source.n57 source.n53 3.44771
R177 source.n45 source.n41 3.44771
R178 source.n5 source.n1 3.44771
R179 source.n17 source.n13 3.44771
R180 source.n25 source.n21 3.44771
R181 source.n37 source.n33 3.44771
R182 source.n39 source.n31 0.974638
R183 source.n31 source.n29 0.974638
R184 source.n29 source.n27 0.974638
R185 source.n19 source.n11 0.974638
R186 source.n11 source.n9 0.974638
R187 source.n9 source.n7 0.974638
R188 source.n49 source.n47 0.974638
R189 source.n51 source.n49 0.974638
R190 source.n59 source.n51 0.974638
R191 source.n69 source.n67 0.974638
R192 source.n71 source.n69 0.974638
R193 source.n79 source.n71 0.974638
R194 source.n27 source.n19 0.470328
R195 source.n67 source.n59 0.470328
R196 source source.n80 0.188
R197 drain_right.n6 drain_right.n4 101.769
R198 drain_right.n3 drain_right.n2 101.715
R199 drain_right.n3 drain_right.n0 101.715
R200 drain_right.n6 drain_right.n5 100.796
R201 drain_right.n8 drain_right.n7 100.796
R202 drain_right.n3 drain_right.n1 100.796
R203 drain_right drain_right.n3 24.1088
R204 drain_right.n1 drain_right.t0 9.9005
R205 drain_right.n1 drain_right.t10 9.9005
R206 drain_right.n2 drain_right.t5 9.9005
R207 drain_right.n2 drain_right.t9 9.9005
R208 drain_right.n0 drain_right.t1 9.9005
R209 drain_right.n0 drain_right.t11 9.9005
R210 drain_right.n4 drain_right.t7 9.9005
R211 drain_right.n4 drain_right.t6 9.9005
R212 drain_right.n5 drain_right.t3 9.9005
R213 drain_right.n5 drain_right.t8 9.9005
R214 drain_right.n7 drain_right.t4 9.9005
R215 drain_right.n7 drain_right.t2 9.9005
R216 drain_right drain_right.n8 6.62735
R217 drain_right.n8 drain_right.n6 0.974638
R218 plus.n6 plus.n3 161.3
R219 plus.n11 plus.n10 161.3
R220 plus.n12 plus.n1 161.3
R221 plus.n13 plus.n0 161.3
R222 plus.n15 plus.n14 161.3
R223 plus.n22 plus.n19 161.3
R224 plus.n27 plus.n26 161.3
R225 plus.n28 plus.n17 161.3
R226 plus.n29 plus.n16 161.3
R227 plus.n31 plus.n30 161.3
R228 plus.n4 plus.t10 130.75
R229 plus.n20 plus.t9 130.75
R230 plus.n14 plus.t4 109.355
R231 plus.n12 plus.t7 109.355
R232 plus.n2 plus.t5 109.355
R233 plus.n7 plus.t6 109.355
R234 plus.n5 plus.t8 109.355
R235 plus.n30 plus.t2 109.355
R236 plus.n28 plus.t3 109.355
R237 plus.n18 plus.t1 109.355
R238 plus.n23 plus.t11 109.355
R239 plus.n21 plus.t0 109.355
R240 plus.n8 plus.n7 80.6037
R241 plus.n9 plus.n2 80.6037
R242 plus.n24 plus.n23 80.6037
R243 plus.n25 plus.n18 80.6037
R244 plus.n7 plus.n2 48.2005
R245 plus.n23 plus.n18 48.2005
R246 plus.n4 plus.n3 44.853
R247 plus.n20 plus.n19 44.853
R248 plus.n11 plus.n2 41.6278
R249 plus.n7 plus.n6 41.6278
R250 plus.n27 plus.n18 41.6278
R251 plus.n23 plus.n22 41.6278
R252 plus plus.n31 28.1202
R253 plus.n14 plus.n13 25.5611
R254 plus.n30 plus.n29 25.5611
R255 plus.n13 plus.n12 22.6399
R256 plus.n29 plus.n28 22.6399
R257 plus.n5 plus.n4 20.5405
R258 plus.n21 plus.n20 20.5405
R259 plus plus.n15 8.55732
R260 plus.n12 plus.n11 6.57323
R261 plus.n6 plus.n5 6.57323
R262 plus.n28 plus.n27 6.57323
R263 plus.n22 plus.n21 6.57323
R264 plus.n9 plus.n8 0.380177
R265 plus.n25 plus.n24 0.380177
R266 plus.n8 plus.n3 0.285035
R267 plus.n10 plus.n9 0.285035
R268 plus.n26 plus.n25 0.285035
R269 plus.n24 plus.n19 0.285035
R270 plus.n10 plus.n1 0.189894
R271 plus.n1 plus.n0 0.189894
R272 plus.n15 plus.n0 0.189894
R273 plus.n31 plus.n16 0.189894
R274 plus.n17 plus.n16 0.189894
R275 plus.n26 plus.n17 0.189894
R276 drain_left.n6 drain_left.n4 101.769
R277 drain_left.n3 drain_left.n2 101.715
R278 drain_left.n3 drain_left.n0 101.715
R279 drain_left.n8 drain_left.n7 100.796
R280 drain_left.n6 drain_left.n5 100.796
R281 drain_left.n3 drain_left.n1 100.796
R282 drain_left drain_left.n3 24.662
R283 drain_left.n1 drain_left.t10 9.9005
R284 drain_left.n1 drain_left.t0 9.9005
R285 drain_left.n2 drain_left.t11 9.9005
R286 drain_left.n2 drain_left.t2 9.9005
R287 drain_left.n0 drain_left.t9 9.9005
R288 drain_left.n0 drain_left.t8 9.9005
R289 drain_left.n7 drain_left.t4 9.9005
R290 drain_left.n7 drain_left.t7 9.9005
R291 drain_left.n5 drain_left.t5 9.9005
R292 drain_left.n5 drain_left.t6 9.9005
R293 drain_left.n4 drain_left.t1 9.9005
R294 drain_left.n4 drain_left.t3 9.9005
R295 drain_left drain_left.n8 6.62735
R296 drain_left.n8 drain_left.n6 0.974638
C0 drain_right plus 0.388551f
C1 drain_left minus 0.178088f
C2 drain_left drain_right 1.1621f
C3 drain_left plus 2.05538f
C4 source minus 2.31636f
C5 source drain_right 4.88724f
C6 drain_right minus 1.82918f
C7 source plus 2.33032f
C8 plus minus 4.16143f
C9 source drain_left 4.88468f
C10 drain_right a_n2298_n1288# 3.94346f
C11 drain_left a_n2298_n1288# 4.714129f
C12 source a_n2298_n1288# 3.278924f
C13 minus a_n2298_n1288# 8.247768f
C14 plus a_n2298_n1288# 9.48837f
C15 drain_left.t9 a_n2298_n1288# 0.041871f
C16 drain_left.t8 a_n2298_n1288# 0.041871f
C17 drain_left.n0 a_n2298_n1288# 0.266444f
C18 drain_left.t10 a_n2298_n1288# 0.041871f
C19 drain_left.t0 a_n2298_n1288# 0.041871f
C20 drain_left.n1 a_n2298_n1288# 0.26305f
C21 drain_left.t11 a_n2298_n1288# 0.041871f
C22 drain_left.t2 a_n2298_n1288# 0.041871f
C23 drain_left.n2 a_n2298_n1288# 0.266444f
C24 drain_left.n3 a_n2298_n1288# 1.93699f
C25 drain_left.t1 a_n2298_n1288# 0.041871f
C26 drain_left.t3 a_n2298_n1288# 0.041871f
C27 drain_left.n4 a_n2298_n1288# 0.266686f
C28 drain_left.t5 a_n2298_n1288# 0.041871f
C29 drain_left.t6 a_n2298_n1288# 0.041871f
C30 drain_left.n5 a_n2298_n1288# 0.263051f
C31 drain_left.n6 a_n2298_n1288# 0.745225f
C32 drain_left.t4 a_n2298_n1288# 0.041871f
C33 drain_left.t7 a_n2298_n1288# 0.041871f
C34 drain_left.n7 a_n2298_n1288# 0.263051f
C35 drain_left.n8 a_n2298_n1288# 0.606658f
C36 plus.n0 a_n2298_n1288# 0.045139f
C37 plus.t4 a_n2298_n1288# 0.223656f
C38 plus.t7 a_n2298_n1288# 0.223656f
C39 plus.n1 a_n2298_n1288# 0.045139f
C40 plus.t5 a_n2298_n1288# 0.223656f
C41 plus.n2 a_n2298_n1288# 0.163952f
C42 plus.n3 a_n2298_n1288# 0.207225f
C43 plus.t6 a_n2298_n1288# 0.223656f
C44 plus.t8 a_n2298_n1288# 0.223656f
C45 plus.t10 a_n2298_n1288# 0.248829f
C46 plus.n4 a_n2298_n1288# 0.133151f
C47 plus.n5 a_n2298_n1288# 0.15486f
C48 plus.n6 a_n2298_n1288# 0.010243f
C49 plus.n7 a_n2298_n1288# 0.163952f
C50 plus.n8 a_n2298_n1288# 0.075186f
C51 plus.n9 a_n2298_n1288# 0.075186f
C52 plus.n10 a_n2298_n1288# 0.060233f
C53 plus.n11 a_n2298_n1288# 0.010243f
C54 plus.n12 a_n2298_n1288# 0.151344f
C55 plus.n13 a_n2298_n1288# 0.010243f
C56 plus.n14 a_n2298_n1288# 0.150648f
C57 plus.n15 a_n2298_n1288# 0.345069f
C58 plus.n16 a_n2298_n1288# 0.045139f
C59 plus.t2 a_n2298_n1288# 0.223656f
C60 plus.n17 a_n2298_n1288# 0.045139f
C61 plus.t3 a_n2298_n1288# 0.223656f
C62 plus.t1 a_n2298_n1288# 0.223656f
C63 plus.n18 a_n2298_n1288# 0.163952f
C64 plus.n19 a_n2298_n1288# 0.207225f
C65 plus.t11 a_n2298_n1288# 0.223656f
C66 plus.t9 a_n2298_n1288# 0.248829f
C67 plus.n20 a_n2298_n1288# 0.133151f
C68 plus.t0 a_n2298_n1288# 0.223656f
C69 plus.n21 a_n2298_n1288# 0.15486f
C70 plus.n22 a_n2298_n1288# 0.010243f
C71 plus.n23 a_n2298_n1288# 0.163952f
C72 plus.n24 a_n2298_n1288# 0.075186f
C73 plus.n25 a_n2298_n1288# 0.075186f
C74 plus.n26 a_n2298_n1288# 0.060233f
C75 plus.n27 a_n2298_n1288# 0.010243f
C76 plus.n28 a_n2298_n1288# 0.151344f
C77 plus.n29 a_n2298_n1288# 0.010243f
C78 plus.n30 a_n2298_n1288# 0.150648f
C79 plus.n31 a_n2298_n1288# 1.15531f
C80 drain_right.t1 a_n2298_n1288# 0.02975f
C81 drain_right.t11 a_n2298_n1288# 0.02975f
C82 drain_right.n0 a_n2298_n1288# 0.189313f
C83 drain_right.t0 a_n2298_n1288# 0.02975f
C84 drain_right.t10 a_n2298_n1288# 0.02975f
C85 drain_right.n1 a_n2298_n1288# 0.186902f
C86 drain_right.t5 a_n2298_n1288# 0.02975f
C87 drain_right.t9 a_n2298_n1288# 0.02975f
C88 drain_right.n2 a_n2298_n1288# 0.189313f
C89 drain_right.n3 a_n2298_n1288# 1.33955f
C90 drain_right.t7 a_n2298_n1288# 0.02975f
C91 drain_right.t6 a_n2298_n1288# 0.02975f
C92 drain_right.n4 a_n2298_n1288# 0.189486f
C93 drain_right.t3 a_n2298_n1288# 0.02975f
C94 drain_right.t8 a_n2298_n1288# 0.02975f
C95 drain_right.n5 a_n2298_n1288# 0.186903f
C96 drain_right.n6 a_n2298_n1288# 0.529497f
C97 drain_right.t4 a_n2298_n1288# 0.02975f
C98 drain_right.t2 a_n2298_n1288# 0.02975f
C99 drain_right.n7 a_n2298_n1288# 0.186903f
C100 drain_right.n8 a_n2298_n1288# 0.431042f
C101 source.n0 a_n2298_n1288# 0.042368f
C102 source.n1 a_n2298_n1288# 0.093743f
C103 source.t9 a_n2298_n1288# 0.07035f
C104 source.n2 a_n2298_n1288# 0.073367f
C105 source.n3 a_n2298_n1288# 0.023651f
C106 source.n4 a_n2298_n1288# 0.015598f
C107 source.n5 a_n2298_n1288# 0.206633f
C108 source.n6 a_n2298_n1288# 0.046445f
C109 source.n7 a_n2298_n1288# 0.509646f
C110 source.t5 a_n2298_n1288# 0.045877f
C111 source.t2 a_n2298_n1288# 0.045877f
C112 source.n8 a_n2298_n1288# 0.245257f
C113 source.n9 a_n2298_n1288# 0.407905f
C114 source.t10 a_n2298_n1288# 0.045877f
C115 source.t7 a_n2298_n1288# 0.045877f
C116 source.n10 a_n2298_n1288# 0.245257f
C117 source.n11 a_n2298_n1288# 0.407905f
C118 source.n12 a_n2298_n1288# 0.042368f
C119 source.n13 a_n2298_n1288# 0.093743f
C120 source.t6 a_n2298_n1288# 0.07035f
C121 source.n14 a_n2298_n1288# 0.073367f
C122 source.n15 a_n2298_n1288# 0.023651f
C123 source.n16 a_n2298_n1288# 0.015598f
C124 source.n17 a_n2298_n1288# 0.206633f
C125 source.n18 a_n2298_n1288# 0.046445f
C126 source.n19 a_n2298_n1288# 0.158956f
C127 source.n20 a_n2298_n1288# 0.042368f
C128 source.n21 a_n2298_n1288# 0.093743f
C129 source.t17 a_n2298_n1288# 0.07035f
C130 source.n22 a_n2298_n1288# 0.073367f
C131 source.n23 a_n2298_n1288# 0.023651f
C132 source.n24 a_n2298_n1288# 0.015598f
C133 source.n25 a_n2298_n1288# 0.206633f
C134 source.n26 a_n2298_n1288# 0.046445f
C135 source.n27 a_n2298_n1288# 0.158956f
C136 source.t19 a_n2298_n1288# 0.045877f
C137 source.t22 a_n2298_n1288# 0.045877f
C138 source.n28 a_n2298_n1288# 0.245257f
C139 source.n29 a_n2298_n1288# 0.407905f
C140 source.t21 a_n2298_n1288# 0.045877f
C141 source.t18 a_n2298_n1288# 0.045877f
C142 source.n30 a_n2298_n1288# 0.245257f
C143 source.n31 a_n2298_n1288# 0.407905f
C144 source.n32 a_n2298_n1288# 0.042368f
C145 source.n33 a_n2298_n1288# 0.093743f
C146 source.t16 a_n2298_n1288# 0.07035f
C147 source.n34 a_n2298_n1288# 0.073367f
C148 source.n35 a_n2298_n1288# 0.023651f
C149 source.n36 a_n2298_n1288# 0.015598f
C150 source.n37 a_n2298_n1288# 0.206633f
C151 source.n38 a_n2298_n1288# 0.046445f
C152 source.n39 a_n2298_n1288# 0.789526f
C153 source.n40 a_n2298_n1288# 0.042368f
C154 source.n41 a_n2298_n1288# 0.093743f
C155 source.t3 a_n2298_n1288# 0.07035f
C156 source.n42 a_n2298_n1288# 0.073367f
C157 source.n43 a_n2298_n1288# 0.023651f
C158 source.n44 a_n2298_n1288# 0.015598f
C159 source.n45 a_n2298_n1288# 0.206633f
C160 source.n46 a_n2298_n1288# 0.046445f
C161 source.n47 a_n2298_n1288# 0.789526f
C162 source.t8 a_n2298_n1288# 0.045877f
C163 source.t1 a_n2298_n1288# 0.045877f
C164 source.n48 a_n2298_n1288# 0.245255f
C165 source.n49 a_n2298_n1288# 0.407906f
C166 source.t0 a_n2298_n1288# 0.045877f
C167 source.t4 a_n2298_n1288# 0.045877f
C168 source.n50 a_n2298_n1288# 0.245255f
C169 source.n51 a_n2298_n1288# 0.407906f
C170 source.n52 a_n2298_n1288# 0.042368f
C171 source.n53 a_n2298_n1288# 0.093743f
C172 source.t11 a_n2298_n1288# 0.07035f
C173 source.n54 a_n2298_n1288# 0.073367f
C174 source.n55 a_n2298_n1288# 0.023651f
C175 source.n56 a_n2298_n1288# 0.015598f
C176 source.n57 a_n2298_n1288# 0.206633f
C177 source.n58 a_n2298_n1288# 0.046445f
C178 source.n59 a_n2298_n1288# 0.158956f
C179 source.n60 a_n2298_n1288# 0.042368f
C180 source.n61 a_n2298_n1288# 0.093743f
C181 source.t23 a_n2298_n1288# 0.07035f
C182 source.n62 a_n2298_n1288# 0.073367f
C183 source.n63 a_n2298_n1288# 0.023651f
C184 source.n64 a_n2298_n1288# 0.015598f
C185 source.n65 a_n2298_n1288# 0.206633f
C186 source.n66 a_n2298_n1288# 0.046445f
C187 source.n67 a_n2298_n1288# 0.158956f
C188 source.t13 a_n2298_n1288# 0.045877f
C189 source.t20 a_n2298_n1288# 0.045877f
C190 source.n68 a_n2298_n1288# 0.245255f
C191 source.n69 a_n2298_n1288# 0.407906f
C192 source.t12 a_n2298_n1288# 0.045877f
C193 source.t15 a_n2298_n1288# 0.045877f
C194 source.n70 a_n2298_n1288# 0.245255f
C195 source.n71 a_n2298_n1288# 0.407906f
C196 source.n72 a_n2298_n1288# 0.042368f
C197 source.n73 a_n2298_n1288# 0.093743f
C198 source.t14 a_n2298_n1288# 0.07035f
C199 source.n74 a_n2298_n1288# 0.073367f
C200 source.n75 a_n2298_n1288# 0.023651f
C201 source.n76 a_n2298_n1288# 0.015598f
C202 source.n77 a_n2298_n1288# 0.206633f
C203 source.n78 a_n2298_n1288# 0.046445f
C204 source.n79 a_n2298_n1288# 0.354588f
C205 source.n80 a_n2298_n1288# 0.735466f
C206 minus.n0 a_n2298_n1288# 0.033759f
C207 minus.n1 a_n2298_n1288# 0.007661f
C208 minus.t9 a_n2298_n1288# 0.167267f
C209 minus.n2 a_n2298_n1288# 0.056229f
C210 minus.t4 a_n2298_n1288# 0.167267f
C211 minus.n3 a_n2298_n1288# 0.115816f
C212 minus.t5 a_n2298_n1288# 0.186093f
C213 minus.n4 a_n2298_n1288# 0.09958f
C214 minus.n5 a_n2298_n1288# 0.154978f
C215 minus.n6 a_n2298_n1288# 0.007661f
C216 minus.t3 a_n2298_n1288# 0.167267f
C217 minus.n7 a_n2298_n1288# 0.122616f
C218 minus.t8 a_n2298_n1288# 0.167267f
C219 minus.n8 a_n2298_n1288# 0.122616f
C220 minus.n9 a_n2298_n1288# 0.056229f
C221 minus.n10 a_n2298_n1288# 0.045047f
C222 minus.n11 a_n2298_n1288# 0.033759f
C223 minus.n12 a_n2298_n1288# 0.113186f
C224 minus.n13 a_n2298_n1288# 0.007661f
C225 minus.t7 a_n2298_n1288# 0.167267f
C226 minus.n14 a_n2298_n1288# 0.112666f
C227 minus.n15 a_n2298_n1288# 0.907026f
C228 minus.n16 a_n2298_n1288# 0.033759f
C229 minus.n17 a_n2298_n1288# 0.007661f
C230 minus.n18 a_n2298_n1288# 0.056229f
C231 minus.t0 a_n2298_n1288# 0.167267f
C232 minus.n19 a_n2298_n1288# 0.115816f
C233 minus.t10 a_n2298_n1288# 0.186093f
C234 minus.n20 a_n2298_n1288# 0.09958f
C235 minus.n21 a_n2298_n1288# 0.154978f
C236 minus.n22 a_n2298_n1288# 0.007661f
C237 minus.t11 a_n2298_n1288# 0.167267f
C238 minus.n23 a_n2298_n1288# 0.122616f
C239 minus.t1 a_n2298_n1288# 0.167267f
C240 minus.n24 a_n2298_n1288# 0.122616f
C241 minus.n25 a_n2298_n1288# 0.056229f
C242 minus.n26 a_n2298_n1288# 0.045047f
C243 minus.n27 a_n2298_n1288# 0.033759f
C244 minus.t6 a_n2298_n1288# 0.167267f
C245 minus.n28 a_n2298_n1288# 0.113186f
C246 minus.n29 a_n2298_n1288# 0.007661f
C247 minus.t2 a_n2298_n1288# 0.167267f
C248 minus.n30 a_n2298_n1288# 0.112666f
C249 minus.n31 a_n2298_n1288# 0.236564f
C250 minus.n32 a_n2298_n1288# 1.11046f
.ends

