* NGSPICE file created from diffpair416.ext - technology: sky130A

.subckt diffpair416 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t26 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X1 drain_right.t12 minus.t1 source.t24 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X2 drain_right.t11 minus.t2 source.t22 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X3 drain_right.t10 minus.t3 source.t19 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X4 a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X5 drain_left.t13 plus.t0 source.t7 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X6 source.t2 plus.t1 drain_left.t12 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X7 source.t18 minus.t4 drain_right.t9 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X8 source.t27 minus.t5 drain_right.t8 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X9 source.t25 minus.t6 drain_right.t7 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X10 source.t17 minus.t7 drain_right.t6 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X11 source.t14 minus.t8 drain_right.t5 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X12 a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X13 drain_right.t4 minus.t9 source.t20 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X14 source.t1 plus.t2 drain_left.t11 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X15 drain_left.t10 plus.t3 source.t3 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X16 drain_right.t3 minus.t10 source.t15 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X17 drain_right.t2 minus.t11 source.t16 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X18 drain_right.t1 minus.t12 source.t23 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X19 source.t6 plus.t4 drain_left.t9 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X20 source.t8 plus.t5 drain_left.t8 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X21 a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X22 a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X23 drain_left.t7 plus.t6 source.t9 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X24 source.t0 plus.t7 drain_left.t6 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X25 drain_left.t5 plus.t8 source.t11 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X26 drain_left.t4 plus.t9 source.t4 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X27 drain_left.t3 plus.t10 source.t10 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X28 source.t21 minus.t13 drain_right.t0 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X29 drain_left.t2 plus.t11 source.t13 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X30 drain_left.t1 plus.t12 source.t5 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X31 source.t12 plus.t13 drain_left.t0 a_n1564_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 minus.n14 minus.t1 1652.31
R1 minus.n3 minus.t11 1652.31
R2 minus.n30 minus.t9 1652.31
R3 minus.n19 minus.t3 1652.31
R4 minus.n13 minus.t7 1602.65
R5 minus.n11 minus.t12 1602.65
R6 minus.n1 minus.t13 1602.65
R7 minus.n6 minus.t0 1602.65
R8 minus.n4 minus.t8 1602.65
R9 minus.n29 minus.t6 1602.65
R10 minus.n27 minus.t10 1602.65
R11 minus.n17 minus.t4 1602.65
R12 minus.n22 minus.t2 1602.65
R13 minus.n20 minus.t5 1602.65
R14 minus.n3 minus.n2 161.489
R15 minus.n19 minus.n18 161.489
R16 minus.n15 minus.n14 161.3
R17 minus.n12 minus.n0 161.3
R18 minus.n10 minus.n9 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n5 minus.n2 161.3
R21 minus.n31 minus.n30 161.3
R22 minus.n28 minus.n16 161.3
R23 minus.n26 minus.n25 161.3
R24 minus.n24 minus.n23 161.3
R25 minus.n21 minus.n18 161.3
R26 minus.n13 minus.n12 45.2793
R27 minus.n5 minus.n4 45.2793
R28 minus.n21 minus.n20 45.2793
R29 minus.n29 minus.n28 45.2793
R30 minus.n11 minus.n10 40.8975
R31 minus.n7 minus.n6 40.8975
R32 minus.n23 minus.n22 40.8975
R33 minus.n27 minus.n26 40.8975
R34 minus.n10 minus.n1 36.5157
R35 minus.n7 minus.n1 36.5157
R36 minus.n23 minus.n17 36.5157
R37 minus.n26 minus.n17 36.5157
R38 minus.n32 minus.n15 35.0062
R39 minus.n12 minus.n11 32.1338
R40 minus.n6 minus.n5 32.1338
R41 minus.n22 minus.n21 32.1338
R42 minus.n28 minus.n27 32.1338
R43 minus.n14 minus.n13 27.752
R44 minus.n4 minus.n3 27.752
R45 minus.n20 minus.n19 27.752
R46 minus.n30 minus.n29 27.752
R47 minus.n32 minus.n31 6.46073
R48 minus.n15 minus.n0 0.189894
R49 minus.n9 minus.n0 0.189894
R50 minus.n9 minus.n8 0.189894
R51 minus.n8 minus.n2 0.189894
R52 minus.n24 minus.n18 0.189894
R53 minus.n25 minus.n24 0.189894
R54 minus.n25 minus.n16 0.189894
R55 minus.n31 minus.n16 0.189894
R56 minus minus.n32 0.188
R57 source.n282 source.n222 289.615
R58 source.n210 source.n150 289.615
R59 source.n60 source.n0 289.615
R60 source.n132 source.n72 289.615
R61 source.n242 source.n241 185
R62 source.n247 source.n246 185
R63 source.n249 source.n248 185
R64 source.n238 source.n237 185
R65 source.n255 source.n254 185
R66 source.n257 source.n256 185
R67 source.n234 source.n233 185
R68 source.n264 source.n263 185
R69 source.n265 source.n232 185
R70 source.n267 source.n266 185
R71 source.n230 source.n229 185
R72 source.n273 source.n272 185
R73 source.n275 source.n274 185
R74 source.n226 source.n225 185
R75 source.n281 source.n280 185
R76 source.n283 source.n282 185
R77 source.n170 source.n169 185
R78 source.n175 source.n174 185
R79 source.n177 source.n176 185
R80 source.n166 source.n165 185
R81 source.n183 source.n182 185
R82 source.n185 source.n184 185
R83 source.n162 source.n161 185
R84 source.n192 source.n191 185
R85 source.n193 source.n160 185
R86 source.n195 source.n194 185
R87 source.n158 source.n157 185
R88 source.n201 source.n200 185
R89 source.n203 source.n202 185
R90 source.n154 source.n153 185
R91 source.n209 source.n208 185
R92 source.n211 source.n210 185
R93 source.n61 source.n60 185
R94 source.n59 source.n58 185
R95 source.n4 source.n3 185
R96 source.n53 source.n52 185
R97 source.n51 source.n50 185
R98 source.n8 source.n7 185
R99 source.n45 source.n44 185
R100 source.n43 source.n10 185
R101 source.n42 source.n41 185
R102 source.n13 source.n11 185
R103 source.n36 source.n35 185
R104 source.n34 source.n33 185
R105 source.n17 source.n16 185
R106 source.n28 source.n27 185
R107 source.n26 source.n25 185
R108 source.n21 source.n20 185
R109 source.n133 source.n132 185
R110 source.n131 source.n130 185
R111 source.n76 source.n75 185
R112 source.n125 source.n124 185
R113 source.n123 source.n122 185
R114 source.n80 source.n79 185
R115 source.n117 source.n116 185
R116 source.n115 source.n82 185
R117 source.n114 source.n113 185
R118 source.n85 source.n83 185
R119 source.n108 source.n107 185
R120 source.n106 source.n105 185
R121 source.n89 source.n88 185
R122 source.n100 source.n99 185
R123 source.n98 source.n97 185
R124 source.n93 source.n92 185
R125 source.n243 source.t20 149.524
R126 source.n171 source.t13 149.524
R127 source.n22 source.t7 149.524
R128 source.n94 source.t16 149.524
R129 source.n247 source.n241 104.615
R130 source.n248 source.n247 104.615
R131 source.n248 source.n237 104.615
R132 source.n255 source.n237 104.615
R133 source.n256 source.n255 104.615
R134 source.n256 source.n233 104.615
R135 source.n264 source.n233 104.615
R136 source.n265 source.n264 104.615
R137 source.n266 source.n265 104.615
R138 source.n266 source.n229 104.615
R139 source.n273 source.n229 104.615
R140 source.n274 source.n273 104.615
R141 source.n274 source.n225 104.615
R142 source.n281 source.n225 104.615
R143 source.n282 source.n281 104.615
R144 source.n175 source.n169 104.615
R145 source.n176 source.n175 104.615
R146 source.n176 source.n165 104.615
R147 source.n183 source.n165 104.615
R148 source.n184 source.n183 104.615
R149 source.n184 source.n161 104.615
R150 source.n192 source.n161 104.615
R151 source.n193 source.n192 104.615
R152 source.n194 source.n193 104.615
R153 source.n194 source.n157 104.615
R154 source.n201 source.n157 104.615
R155 source.n202 source.n201 104.615
R156 source.n202 source.n153 104.615
R157 source.n209 source.n153 104.615
R158 source.n210 source.n209 104.615
R159 source.n60 source.n59 104.615
R160 source.n59 source.n3 104.615
R161 source.n52 source.n3 104.615
R162 source.n52 source.n51 104.615
R163 source.n51 source.n7 104.615
R164 source.n44 source.n7 104.615
R165 source.n44 source.n43 104.615
R166 source.n43 source.n42 104.615
R167 source.n42 source.n11 104.615
R168 source.n35 source.n11 104.615
R169 source.n35 source.n34 104.615
R170 source.n34 source.n16 104.615
R171 source.n27 source.n16 104.615
R172 source.n27 source.n26 104.615
R173 source.n26 source.n20 104.615
R174 source.n132 source.n131 104.615
R175 source.n131 source.n75 104.615
R176 source.n124 source.n75 104.615
R177 source.n124 source.n123 104.615
R178 source.n123 source.n79 104.615
R179 source.n116 source.n79 104.615
R180 source.n116 source.n115 104.615
R181 source.n115 source.n114 104.615
R182 source.n114 source.n83 104.615
R183 source.n107 source.n83 104.615
R184 source.n107 source.n106 104.615
R185 source.n106 source.n88 104.615
R186 source.n99 source.n88 104.615
R187 source.n99 source.n98 104.615
R188 source.n98 source.n92 104.615
R189 source.t20 source.n241 52.3082
R190 source.t13 source.n169 52.3082
R191 source.t7 source.n20 52.3082
R192 source.t16 source.n92 52.3082
R193 source.n67 source.n66 42.8739
R194 source.n69 source.n68 42.8739
R195 source.n71 source.n70 42.8739
R196 source.n139 source.n138 42.8739
R197 source.n141 source.n140 42.8739
R198 source.n143 source.n142 42.8739
R199 source.n221 source.n220 42.8737
R200 source.n219 source.n218 42.8737
R201 source.n217 source.n216 42.8737
R202 source.n149 source.n148 42.8737
R203 source.n147 source.n146 42.8737
R204 source.n145 source.n144 42.8737
R205 source.n287 source.n286 29.8581
R206 source.n215 source.n214 29.8581
R207 source.n65 source.n64 29.8581
R208 source.n137 source.n136 29.8581
R209 source.n145 source.n143 22.2015
R210 source.n288 source.n65 16.2532
R211 source.n267 source.n232 13.1884
R212 source.n195 source.n160 13.1884
R213 source.n45 source.n10 13.1884
R214 source.n117 source.n82 13.1884
R215 source.n263 source.n262 12.8005
R216 source.n268 source.n230 12.8005
R217 source.n191 source.n190 12.8005
R218 source.n196 source.n158 12.8005
R219 source.n46 source.n8 12.8005
R220 source.n41 source.n12 12.8005
R221 source.n118 source.n80 12.8005
R222 source.n113 source.n84 12.8005
R223 source.n261 source.n234 12.0247
R224 source.n272 source.n271 12.0247
R225 source.n189 source.n162 12.0247
R226 source.n200 source.n199 12.0247
R227 source.n50 source.n49 12.0247
R228 source.n40 source.n13 12.0247
R229 source.n122 source.n121 12.0247
R230 source.n112 source.n85 12.0247
R231 source.n258 source.n257 11.249
R232 source.n275 source.n228 11.249
R233 source.n186 source.n185 11.249
R234 source.n203 source.n156 11.249
R235 source.n53 source.n6 11.249
R236 source.n37 source.n36 11.249
R237 source.n125 source.n78 11.249
R238 source.n109 source.n108 11.249
R239 source.n254 source.n236 10.4732
R240 source.n276 source.n226 10.4732
R241 source.n182 source.n164 10.4732
R242 source.n204 source.n154 10.4732
R243 source.n54 source.n4 10.4732
R244 source.n33 source.n15 10.4732
R245 source.n126 source.n76 10.4732
R246 source.n105 source.n87 10.4732
R247 source.n243 source.n242 10.2747
R248 source.n171 source.n170 10.2747
R249 source.n22 source.n21 10.2747
R250 source.n94 source.n93 10.2747
R251 source.n253 source.n238 9.69747
R252 source.n280 source.n279 9.69747
R253 source.n181 source.n166 9.69747
R254 source.n208 source.n207 9.69747
R255 source.n58 source.n57 9.69747
R256 source.n32 source.n17 9.69747
R257 source.n130 source.n129 9.69747
R258 source.n104 source.n89 9.69747
R259 source.n286 source.n285 9.45567
R260 source.n214 source.n213 9.45567
R261 source.n64 source.n63 9.45567
R262 source.n136 source.n135 9.45567
R263 source.n285 source.n284 9.3005
R264 source.n224 source.n223 9.3005
R265 source.n279 source.n278 9.3005
R266 source.n277 source.n276 9.3005
R267 source.n228 source.n227 9.3005
R268 source.n271 source.n270 9.3005
R269 source.n269 source.n268 9.3005
R270 source.n245 source.n244 9.3005
R271 source.n240 source.n239 9.3005
R272 source.n251 source.n250 9.3005
R273 source.n253 source.n252 9.3005
R274 source.n236 source.n235 9.3005
R275 source.n259 source.n258 9.3005
R276 source.n261 source.n260 9.3005
R277 source.n262 source.n231 9.3005
R278 source.n213 source.n212 9.3005
R279 source.n152 source.n151 9.3005
R280 source.n207 source.n206 9.3005
R281 source.n205 source.n204 9.3005
R282 source.n156 source.n155 9.3005
R283 source.n199 source.n198 9.3005
R284 source.n197 source.n196 9.3005
R285 source.n173 source.n172 9.3005
R286 source.n168 source.n167 9.3005
R287 source.n179 source.n178 9.3005
R288 source.n181 source.n180 9.3005
R289 source.n164 source.n163 9.3005
R290 source.n187 source.n186 9.3005
R291 source.n189 source.n188 9.3005
R292 source.n190 source.n159 9.3005
R293 source.n24 source.n23 9.3005
R294 source.n19 source.n18 9.3005
R295 source.n30 source.n29 9.3005
R296 source.n32 source.n31 9.3005
R297 source.n15 source.n14 9.3005
R298 source.n38 source.n37 9.3005
R299 source.n40 source.n39 9.3005
R300 source.n12 source.n9 9.3005
R301 source.n63 source.n62 9.3005
R302 source.n2 source.n1 9.3005
R303 source.n57 source.n56 9.3005
R304 source.n55 source.n54 9.3005
R305 source.n6 source.n5 9.3005
R306 source.n49 source.n48 9.3005
R307 source.n47 source.n46 9.3005
R308 source.n96 source.n95 9.3005
R309 source.n91 source.n90 9.3005
R310 source.n102 source.n101 9.3005
R311 source.n104 source.n103 9.3005
R312 source.n87 source.n86 9.3005
R313 source.n110 source.n109 9.3005
R314 source.n112 source.n111 9.3005
R315 source.n84 source.n81 9.3005
R316 source.n135 source.n134 9.3005
R317 source.n74 source.n73 9.3005
R318 source.n129 source.n128 9.3005
R319 source.n127 source.n126 9.3005
R320 source.n78 source.n77 9.3005
R321 source.n121 source.n120 9.3005
R322 source.n119 source.n118 9.3005
R323 source.n250 source.n249 8.92171
R324 source.n283 source.n224 8.92171
R325 source.n178 source.n177 8.92171
R326 source.n211 source.n152 8.92171
R327 source.n61 source.n2 8.92171
R328 source.n29 source.n28 8.92171
R329 source.n133 source.n74 8.92171
R330 source.n101 source.n100 8.92171
R331 source.n246 source.n240 8.14595
R332 source.n284 source.n222 8.14595
R333 source.n174 source.n168 8.14595
R334 source.n212 source.n150 8.14595
R335 source.n62 source.n0 8.14595
R336 source.n25 source.n19 8.14595
R337 source.n134 source.n72 8.14595
R338 source.n97 source.n91 8.14595
R339 source.n245 source.n242 7.3702
R340 source.n173 source.n170 7.3702
R341 source.n24 source.n21 7.3702
R342 source.n96 source.n93 7.3702
R343 source.n246 source.n245 5.81868
R344 source.n286 source.n222 5.81868
R345 source.n174 source.n173 5.81868
R346 source.n214 source.n150 5.81868
R347 source.n64 source.n0 5.81868
R348 source.n25 source.n24 5.81868
R349 source.n136 source.n72 5.81868
R350 source.n97 source.n96 5.81868
R351 source.n288 source.n287 5.49188
R352 source.n249 source.n240 5.04292
R353 source.n284 source.n283 5.04292
R354 source.n177 source.n168 5.04292
R355 source.n212 source.n211 5.04292
R356 source.n62 source.n61 5.04292
R357 source.n28 source.n19 5.04292
R358 source.n134 source.n133 5.04292
R359 source.n100 source.n91 5.04292
R360 source.n250 source.n238 4.26717
R361 source.n280 source.n224 4.26717
R362 source.n178 source.n166 4.26717
R363 source.n208 source.n152 4.26717
R364 source.n58 source.n2 4.26717
R365 source.n29 source.n17 4.26717
R366 source.n130 source.n74 4.26717
R367 source.n101 source.n89 4.26717
R368 source.n254 source.n253 3.49141
R369 source.n279 source.n226 3.49141
R370 source.n182 source.n181 3.49141
R371 source.n207 source.n154 3.49141
R372 source.n57 source.n4 3.49141
R373 source.n33 source.n32 3.49141
R374 source.n129 source.n76 3.49141
R375 source.n105 source.n104 3.49141
R376 source.n244 source.n243 2.84303
R377 source.n172 source.n171 2.84303
R378 source.n23 source.n22 2.84303
R379 source.n95 source.n94 2.84303
R380 source.n257 source.n236 2.71565
R381 source.n276 source.n275 2.71565
R382 source.n185 source.n164 2.71565
R383 source.n204 source.n203 2.71565
R384 source.n54 source.n53 2.71565
R385 source.n36 source.n15 2.71565
R386 source.n126 source.n125 2.71565
R387 source.n108 source.n87 2.71565
R388 source.n258 source.n234 1.93989
R389 source.n272 source.n228 1.93989
R390 source.n186 source.n162 1.93989
R391 source.n200 source.n156 1.93989
R392 source.n50 source.n6 1.93989
R393 source.n37 source.n13 1.93989
R394 source.n122 source.n78 1.93989
R395 source.n109 source.n85 1.93989
R396 source.n220 source.t15 1.6505
R397 source.n220 source.t25 1.6505
R398 source.n218 source.t22 1.6505
R399 source.n218 source.t18 1.6505
R400 source.n216 source.t19 1.6505
R401 source.n216 source.t27 1.6505
R402 source.n148 source.t4 1.6505
R403 source.n148 source.t12 1.6505
R404 source.n146 source.t10 1.6505
R405 source.n146 source.t8 1.6505
R406 source.n144 source.t11 1.6505
R407 source.n144 source.t6 1.6505
R408 source.n66 source.t9 1.6505
R409 source.n66 source.t1 1.6505
R410 source.n68 source.t5 1.6505
R411 source.n68 source.t0 1.6505
R412 source.n70 source.t3 1.6505
R413 source.n70 source.t2 1.6505
R414 source.n138 source.t26 1.6505
R415 source.n138 source.t14 1.6505
R416 source.n140 source.t23 1.6505
R417 source.n140 source.t21 1.6505
R418 source.n142 source.t24 1.6505
R419 source.n142 source.t17 1.6505
R420 source.n263 source.n261 1.16414
R421 source.n271 source.n230 1.16414
R422 source.n191 source.n189 1.16414
R423 source.n199 source.n158 1.16414
R424 source.n49 source.n8 1.16414
R425 source.n41 source.n40 1.16414
R426 source.n121 source.n80 1.16414
R427 source.n113 source.n112 1.16414
R428 source.n137 source.n71 0.698776
R429 source.n217 source.n215 0.698776
R430 source.n143 source.n141 0.457397
R431 source.n141 source.n139 0.457397
R432 source.n139 source.n137 0.457397
R433 source.n71 source.n69 0.457397
R434 source.n69 source.n67 0.457397
R435 source.n67 source.n65 0.457397
R436 source.n147 source.n145 0.457397
R437 source.n149 source.n147 0.457397
R438 source.n215 source.n149 0.457397
R439 source.n219 source.n217 0.457397
R440 source.n221 source.n219 0.457397
R441 source.n287 source.n221 0.457397
R442 source.n262 source.n232 0.388379
R443 source.n268 source.n267 0.388379
R444 source.n190 source.n160 0.388379
R445 source.n196 source.n195 0.388379
R446 source.n46 source.n45 0.388379
R447 source.n12 source.n10 0.388379
R448 source.n118 source.n117 0.388379
R449 source.n84 source.n82 0.388379
R450 source source.n288 0.188
R451 source.n244 source.n239 0.155672
R452 source.n251 source.n239 0.155672
R453 source.n252 source.n251 0.155672
R454 source.n252 source.n235 0.155672
R455 source.n259 source.n235 0.155672
R456 source.n260 source.n259 0.155672
R457 source.n260 source.n231 0.155672
R458 source.n269 source.n231 0.155672
R459 source.n270 source.n269 0.155672
R460 source.n270 source.n227 0.155672
R461 source.n277 source.n227 0.155672
R462 source.n278 source.n277 0.155672
R463 source.n278 source.n223 0.155672
R464 source.n285 source.n223 0.155672
R465 source.n172 source.n167 0.155672
R466 source.n179 source.n167 0.155672
R467 source.n180 source.n179 0.155672
R468 source.n180 source.n163 0.155672
R469 source.n187 source.n163 0.155672
R470 source.n188 source.n187 0.155672
R471 source.n188 source.n159 0.155672
R472 source.n197 source.n159 0.155672
R473 source.n198 source.n197 0.155672
R474 source.n198 source.n155 0.155672
R475 source.n205 source.n155 0.155672
R476 source.n206 source.n205 0.155672
R477 source.n206 source.n151 0.155672
R478 source.n213 source.n151 0.155672
R479 source.n63 source.n1 0.155672
R480 source.n56 source.n1 0.155672
R481 source.n56 source.n55 0.155672
R482 source.n55 source.n5 0.155672
R483 source.n48 source.n5 0.155672
R484 source.n48 source.n47 0.155672
R485 source.n47 source.n9 0.155672
R486 source.n39 source.n9 0.155672
R487 source.n39 source.n38 0.155672
R488 source.n38 source.n14 0.155672
R489 source.n31 source.n14 0.155672
R490 source.n31 source.n30 0.155672
R491 source.n30 source.n18 0.155672
R492 source.n23 source.n18 0.155672
R493 source.n135 source.n73 0.155672
R494 source.n128 source.n73 0.155672
R495 source.n128 source.n127 0.155672
R496 source.n127 source.n77 0.155672
R497 source.n120 source.n77 0.155672
R498 source.n120 source.n119 0.155672
R499 source.n119 source.n81 0.155672
R500 source.n111 source.n81 0.155672
R501 source.n111 source.n110 0.155672
R502 source.n110 source.n86 0.155672
R503 source.n103 source.n86 0.155672
R504 source.n103 source.n102 0.155672
R505 source.n102 source.n90 0.155672
R506 source.n95 source.n90 0.155672
R507 drain_right.n60 drain_right.n0 289.615
R508 drain_right.n136 drain_right.n76 289.615
R509 drain_right.n20 drain_right.n19 185
R510 drain_right.n25 drain_right.n24 185
R511 drain_right.n27 drain_right.n26 185
R512 drain_right.n16 drain_right.n15 185
R513 drain_right.n33 drain_right.n32 185
R514 drain_right.n35 drain_right.n34 185
R515 drain_right.n12 drain_right.n11 185
R516 drain_right.n42 drain_right.n41 185
R517 drain_right.n43 drain_right.n10 185
R518 drain_right.n45 drain_right.n44 185
R519 drain_right.n8 drain_right.n7 185
R520 drain_right.n51 drain_right.n50 185
R521 drain_right.n53 drain_right.n52 185
R522 drain_right.n4 drain_right.n3 185
R523 drain_right.n59 drain_right.n58 185
R524 drain_right.n61 drain_right.n60 185
R525 drain_right.n137 drain_right.n136 185
R526 drain_right.n135 drain_right.n134 185
R527 drain_right.n80 drain_right.n79 185
R528 drain_right.n129 drain_right.n128 185
R529 drain_right.n127 drain_right.n126 185
R530 drain_right.n84 drain_right.n83 185
R531 drain_right.n121 drain_right.n120 185
R532 drain_right.n119 drain_right.n86 185
R533 drain_right.n118 drain_right.n117 185
R534 drain_right.n89 drain_right.n87 185
R535 drain_right.n112 drain_right.n111 185
R536 drain_right.n110 drain_right.n109 185
R537 drain_right.n93 drain_right.n92 185
R538 drain_right.n104 drain_right.n103 185
R539 drain_right.n102 drain_right.n101 185
R540 drain_right.n97 drain_right.n96 185
R541 drain_right.n21 drain_right.t10 149.524
R542 drain_right.n98 drain_right.t12 149.524
R543 drain_right.n25 drain_right.n19 104.615
R544 drain_right.n26 drain_right.n25 104.615
R545 drain_right.n26 drain_right.n15 104.615
R546 drain_right.n33 drain_right.n15 104.615
R547 drain_right.n34 drain_right.n33 104.615
R548 drain_right.n34 drain_right.n11 104.615
R549 drain_right.n42 drain_right.n11 104.615
R550 drain_right.n43 drain_right.n42 104.615
R551 drain_right.n44 drain_right.n43 104.615
R552 drain_right.n44 drain_right.n7 104.615
R553 drain_right.n51 drain_right.n7 104.615
R554 drain_right.n52 drain_right.n51 104.615
R555 drain_right.n52 drain_right.n3 104.615
R556 drain_right.n59 drain_right.n3 104.615
R557 drain_right.n60 drain_right.n59 104.615
R558 drain_right.n136 drain_right.n135 104.615
R559 drain_right.n135 drain_right.n79 104.615
R560 drain_right.n128 drain_right.n79 104.615
R561 drain_right.n128 drain_right.n127 104.615
R562 drain_right.n127 drain_right.n83 104.615
R563 drain_right.n120 drain_right.n83 104.615
R564 drain_right.n120 drain_right.n119 104.615
R565 drain_right.n119 drain_right.n118 104.615
R566 drain_right.n118 drain_right.n87 104.615
R567 drain_right.n111 drain_right.n87 104.615
R568 drain_right.n111 drain_right.n110 104.615
R569 drain_right.n110 drain_right.n92 104.615
R570 drain_right.n103 drain_right.n92 104.615
R571 drain_right.n103 drain_right.n102 104.615
R572 drain_right.n102 drain_right.n96 104.615
R573 drain_right.n69 drain_right.n67 60.0094
R574 drain_right.n73 drain_right.n71 60.0094
R575 drain_right.n73 drain_right.n72 59.5527
R576 drain_right.n75 drain_right.n74 59.5527
R577 drain_right.n69 drain_right.n68 59.5525
R578 drain_right.n66 drain_right.n65 59.5525
R579 drain_right.t10 drain_right.n19 52.3082
R580 drain_right.t12 drain_right.n96 52.3082
R581 drain_right.n66 drain_right.n64 46.9938
R582 drain_right.n141 drain_right.n140 46.5369
R583 drain_right drain_right.n70 29.441
R584 drain_right.n45 drain_right.n10 13.1884
R585 drain_right.n121 drain_right.n86 13.1884
R586 drain_right.n41 drain_right.n40 12.8005
R587 drain_right.n46 drain_right.n8 12.8005
R588 drain_right.n122 drain_right.n84 12.8005
R589 drain_right.n117 drain_right.n88 12.8005
R590 drain_right.n39 drain_right.n12 12.0247
R591 drain_right.n50 drain_right.n49 12.0247
R592 drain_right.n126 drain_right.n125 12.0247
R593 drain_right.n116 drain_right.n89 12.0247
R594 drain_right.n36 drain_right.n35 11.249
R595 drain_right.n53 drain_right.n6 11.249
R596 drain_right.n129 drain_right.n82 11.249
R597 drain_right.n113 drain_right.n112 11.249
R598 drain_right.n32 drain_right.n14 10.4732
R599 drain_right.n54 drain_right.n4 10.4732
R600 drain_right.n130 drain_right.n80 10.4732
R601 drain_right.n109 drain_right.n91 10.4732
R602 drain_right.n21 drain_right.n20 10.2747
R603 drain_right.n98 drain_right.n97 10.2747
R604 drain_right.n31 drain_right.n16 9.69747
R605 drain_right.n58 drain_right.n57 9.69747
R606 drain_right.n134 drain_right.n133 9.69747
R607 drain_right.n108 drain_right.n93 9.69747
R608 drain_right.n64 drain_right.n63 9.45567
R609 drain_right.n140 drain_right.n139 9.45567
R610 drain_right.n63 drain_right.n62 9.3005
R611 drain_right.n2 drain_right.n1 9.3005
R612 drain_right.n57 drain_right.n56 9.3005
R613 drain_right.n55 drain_right.n54 9.3005
R614 drain_right.n6 drain_right.n5 9.3005
R615 drain_right.n49 drain_right.n48 9.3005
R616 drain_right.n47 drain_right.n46 9.3005
R617 drain_right.n23 drain_right.n22 9.3005
R618 drain_right.n18 drain_right.n17 9.3005
R619 drain_right.n29 drain_right.n28 9.3005
R620 drain_right.n31 drain_right.n30 9.3005
R621 drain_right.n14 drain_right.n13 9.3005
R622 drain_right.n37 drain_right.n36 9.3005
R623 drain_right.n39 drain_right.n38 9.3005
R624 drain_right.n40 drain_right.n9 9.3005
R625 drain_right.n100 drain_right.n99 9.3005
R626 drain_right.n95 drain_right.n94 9.3005
R627 drain_right.n106 drain_right.n105 9.3005
R628 drain_right.n108 drain_right.n107 9.3005
R629 drain_right.n91 drain_right.n90 9.3005
R630 drain_right.n114 drain_right.n113 9.3005
R631 drain_right.n116 drain_right.n115 9.3005
R632 drain_right.n88 drain_right.n85 9.3005
R633 drain_right.n139 drain_right.n138 9.3005
R634 drain_right.n78 drain_right.n77 9.3005
R635 drain_right.n133 drain_right.n132 9.3005
R636 drain_right.n131 drain_right.n130 9.3005
R637 drain_right.n82 drain_right.n81 9.3005
R638 drain_right.n125 drain_right.n124 9.3005
R639 drain_right.n123 drain_right.n122 9.3005
R640 drain_right.n28 drain_right.n27 8.92171
R641 drain_right.n61 drain_right.n2 8.92171
R642 drain_right.n137 drain_right.n78 8.92171
R643 drain_right.n105 drain_right.n104 8.92171
R644 drain_right.n24 drain_right.n18 8.14595
R645 drain_right.n62 drain_right.n0 8.14595
R646 drain_right.n138 drain_right.n76 8.14595
R647 drain_right.n101 drain_right.n95 8.14595
R648 drain_right.n23 drain_right.n20 7.3702
R649 drain_right.n100 drain_right.n97 7.3702
R650 drain_right drain_right.n141 5.88166
R651 drain_right.n24 drain_right.n23 5.81868
R652 drain_right.n64 drain_right.n0 5.81868
R653 drain_right.n140 drain_right.n76 5.81868
R654 drain_right.n101 drain_right.n100 5.81868
R655 drain_right.n27 drain_right.n18 5.04292
R656 drain_right.n62 drain_right.n61 5.04292
R657 drain_right.n138 drain_right.n137 5.04292
R658 drain_right.n104 drain_right.n95 5.04292
R659 drain_right.n28 drain_right.n16 4.26717
R660 drain_right.n58 drain_right.n2 4.26717
R661 drain_right.n134 drain_right.n78 4.26717
R662 drain_right.n105 drain_right.n93 4.26717
R663 drain_right.n32 drain_right.n31 3.49141
R664 drain_right.n57 drain_right.n4 3.49141
R665 drain_right.n133 drain_right.n80 3.49141
R666 drain_right.n109 drain_right.n108 3.49141
R667 drain_right.n22 drain_right.n21 2.84303
R668 drain_right.n99 drain_right.n98 2.84303
R669 drain_right.n35 drain_right.n14 2.71565
R670 drain_right.n54 drain_right.n53 2.71565
R671 drain_right.n130 drain_right.n129 2.71565
R672 drain_right.n112 drain_right.n91 2.71565
R673 drain_right.n36 drain_right.n12 1.93989
R674 drain_right.n50 drain_right.n6 1.93989
R675 drain_right.n126 drain_right.n82 1.93989
R676 drain_right.n113 drain_right.n89 1.93989
R677 drain_right.n67 drain_right.t7 1.6505
R678 drain_right.n67 drain_right.t4 1.6505
R679 drain_right.n68 drain_right.t9 1.6505
R680 drain_right.n68 drain_right.t3 1.6505
R681 drain_right.n65 drain_right.t8 1.6505
R682 drain_right.n65 drain_right.t11 1.6505
R683 drain_right.n71 drain_right.t5 1.6505
R684 drain_right.n71 drain_right.t2 1.6505
R685 drain_right.n72 drain_right.t0 1.6505
R686 drain_right.n72 drain_right.t13 1.6505
R687 drain_right.n74 drain_right.t6 1.6505
R688 drain_right.n74 drain_right.t1 1.6505
R689 drain_right.n41 drain_right.n39 1.16414
R690 drain_right.n49 drain_right.n8 1.16414
R691 drain_right.n125 drain_right.n84 1.16414
R692 drain_right.n117 drain_right.n116 1.16414
R693 drain_right.n141 drain_right.n75 0.457397
R694 drain_right.n75 drain_right.n73 0.457397
R695 drain_right.n40 drain_right.n10 0.388379
R696 drain_right.n46 drain_right.n45 0.388379
R697 drain_right.n122 drain_right.n121 0.388379
R698 drain_right.n88 drain_right.n86 0.388379
R699 drain_right.n70 drain_right.n66 0.287826
R700 drain_right.n22 drain_right.n17 0.155672
R701 drain_right.n29 drain_right.n17 0.155672
R702 drain_right.n30 drain_right.n29 0.155672
R703 drain_right.n30 drain_right.n13 0.155672
R704 drain_right.n37 drain_right.n13 0.155672
R705 drain_right.n38 drain_right.n37 0.155672
R706 drain_right.n38 drain_right.n9 0.155672
R707 drain_right.n47 drain_right.n9 0.155672
R708 drain_right.n48 drain_right.n47 0.155672
R709 drain_right.n48 drain_right.n5 0.155672
R710 drain_right.n55 drain_right.n5 0.155672
R711 drain_right.n56 drain_right.n55 0.155672
R712 drain_right.n56 drain_right.n1 0.155672
R713 drain_right.n63 drain_right.n1 0.155672
R714 drain_right.n139 drain_right.n77 0.155672
R715 drain_right.n132 drain_right.n77 0.155672
R716 drain_right.n132 drain_right.n131 0.155672
R717 drain_right.n131 drain_right.n81 0.155672
R718 drain_right.n124 drain_right.n81 0.155672
R719 drain_right.n124 drain_right.n123 0.155672
R720 drain_right.n123 drain_right.n85 0.155672
R721 drain_right.n115 drain_right.n85 0.155672
R722 drain_right.n115 drain_right.n114 0.155672
R723 drain_right.n114 drain_right.n90 0.155672
R724 drain_right.n107 drain_right.n90 0.155672
R725 drain_right.n107 drain_right.n106 0.155672
R726 drain_right.n106 drain_right.n94 0.155672
R727 drain_right.n99 drain_right.n94 0.155672
R728 drain_right.n70 drain_right.n69 0.0593781
R729 plus.n3 plus.t3 1652.31
R730 plus.n14 plus.t0 1652.31
R731 plus.n19 plus.t11 1652.31
R732 plus.n30 plus.t8 1652.31
R733 plus.n4 plus.t1 1602.65
R734 plus.n6 plus.t12 1602.65
R735 plus.n1 plus.t7 1602.65
R736 plus.n11 plus.t6 1602.65
R737 plus.n13 plus.t2 1602.65
R738 plus.n20 plus.t13 1602.65
R739 plus.n22 plus.t9 1602.65
R740 plus.n17 plus.t5 1602.65
R741 plus.n27 plus.t10 1602.65
R742 plus.n29 plus.t4 1602.65
R743 plus.n3 plus.n2 161.489
R744 plus.n19 plus.n18 161.489
R745 plus.n5 plus.n2 161.3
R746 plus.n8 plus.n7 161.3
R747 plus.n10 plus.n9 161.3
R748 plus.n12 plus.n0 161.3
R749 plus.n15 plus.n14 161.3
R750 plus.n21 plus.n18 161.3
R751 plus.n24 plus.n23 161.3
R752 plus.n26 plus.n25 161.3
R753 plus.n28 plus.n16 161.3
R754 plus.n31 plus.n30 161.3
R755 plus.n5 plus.n4 45.2793
R756 plus.n13 plus.n12 45.2793
R757 plus.n29 plus.n28 45.2793
R758 plus.n21 plus.n20 45.2793
R759 plus.n7 plus.n6 40.8975
R760 plus.n11 plus.n10 40.8975
R761 plus.n27 plus.n26 40.8975
R762 plus.n23 plus.n22 40.8975
R763 plus.n7 plus.n1 36.5157
R764 plus.n10 plus.n1 36.5157
R765 plus.n26 plus.n17 36.5157
R766 plus.n23 plus.n17 36.5157
R767 plus.n6 plus.n5 32.1338
R768 plus.n12 plus.n11 32.1338
R769 plus.n28 plus.n27 32.1338
R770 plus.n22 plus.n21 32.1338
R771 plus plus.n31 28.8873
R772 plus.n4 plus.n3 27.752
R773 plus.n14 plus.n13 27.752
R774 plus.n30 plus.n29 27.752
R775 plus.n20 plus.n19 27.752
R776 plus plus.n15 12.1047
R777 plus.n8 plus.n2 0.189894
R778 plus.n9 plus.n8 0.189894
R779 plus.n9 plus.n0 0.189894
R780 plus.n15 plus.n0 0.189894
R781 plus.n31 plus.n16 0.189894
R782 plus.n25 plus.n16 0.189894
R783 plus.n25 plus.n24 0.189894
R784 plus.n24 plus.n18 0.189894
R785 drain_left.n60 drain_left.n0 289.615
R786 drain_left.n131 drain_left.n71 289.615
R787 drain_left.n20 drain_left.n19 185
R788 drain_left.n25 drain_left.n24 185
R789 drain_left.n27 drain_left.n26 185
R790 drain_left.n16 drain_left.n15 185
R791 drain_left.n33 drain_left.n32 185
R792 drain_left.n35 drain_left.n34 185
R793 drain_left.n12 drain_left.n11 185
R794 drain_left.n42 drain_left.n41 185
R795 drain_left.n43 drain_left.n10 185
R796 drain_left.n45 drain_left.n44 185
R797 drain_left.n8 drain_left.n7 185
R798 drain_left.n51 drain_left.n50 185
R799 drain_left.n53 drain_left.n52 185
R800 drain_left.n4 drain_left.n3 185
R801 drain_left.n59 drain_left.n58 185
R802 drain_left.n61 drain_left.n60 185
R803 drain_left.n132 drain_left.n131 185
R804 drain_left.n130 drain_left.n129 185
R805 drain_left.n75 drain_left.n74 185
R806 drain_left.n124 drain_left.n123 185
R807 drain_left.n122 drain_left.n121 185
R808 drain_left.n79 drain_left.n78 185
R809 drain_left.n116 drain_left.n115 185
R810 drain_left.n114 drain_left.n81 185
R811 drain_left.n113 drain_left.n112 185
R812 drain_left.n84 drain_left.n82 185
R813 drain_left.n107 drain_left.n106 185
R814 drain_left.n105 drain_left.n104 185
R815 drain_left.n88 drain_left.n87 185
R816 drain_left.n99 drain_left.n98 185
R817 drain_left.n97 drain_left.n96 185
R818 drain_left.n92 drain_left.n91 185
R819 drain_left.n21 drain_left.t5 149.524
R820 drain_left.n93 drain_left.t10 149.524
R821 drain_left.n25 drain_left.n19 104.615
R822 drain_left.n26 drain_left.n25 104.615
R823 drain_left.n26 drain_left.n15 104.615
R824 drain_left.n33 drain_left.n15 104.615
R825 drain_left.n34 drain_left.n33 104.615
R826 drain_left.n34 drain_left.n11 104.615
R827 drain_left.n42 drain_left.n11 104.615
R828 drain_left.n43 drain_left.n42 104.615
R829 drain_left.n44 drain_left.n43 104.615
R830 drain_left.n44 drain_left.n7 104.615
R831 drain_left.n51 drain_left.n7 104.615
R832 drain_left.n52 drain_left.n51 104.615
R833 drain_left.n52 drain_left.n3 104.615
R834 drain_left.n59 drain_left.n3 104.615
R835 drain_left.n60 drain_left.n59 104.615
R836 drain_left.n131 drain_left.n130 104.615
R837 drain_left.n130 drain_left.n74 104.615
R838 drain_left.n123 drain_left.n74 104.615
R839 drain_left.n123 drain_left.n122 104.615
R840 drain_left.n122 drain_left.n78 104.615
R841 drain_left.n115 drain_left.n78 104.615
R842 drain_left.n115 drain_left.n114 104.615
R843 drain_left.n114 drain_left.n113 104.615
R844 drain_left.n113 drain_left.n82 104.615
R845 drain_left.n106 drain_left.n82 104.615
R846 drain_left.n106 drain_left.n105 104.615
R847 drain_left.n105 drain_left.n87 104.615
R848 drain_left.n98 drain_left.n87 104.615
R849 drain_left.n98 drain_left.n97 104.615
R850 drain_left.n97 drain_left.n91 104.615
R851 drain_left.n69 drain_left.n67 60.0094
R852 drain_left.n139 drain_left.n138 59.5527
R853 drain_left.n137 drain_left.n136 59.5527
R854 drain_left.n69 drain_left.n68 59.5525
R855 drain_left.n66 drain_left.n65 59.5525
R856 drain_left.n141 drain_left.n140 59.5525
R857 drain_left.t5 drain_left.n19 52.3082
R858 drain_left.t10 drain_left.n91 52.3082
R859 drain_left.n66 drain_left.n64 46.9938
R860 drain_left.n137 drain_left.n135 46.9938
R861 drain_left drain_left.n70 29.9942
R862 drain_left.n45 drain_left.n10 13.1884
R863 drain_left.n116 drain_left.n81 13.1884
R864 drain_left.n41 drain_left.n40 12.8005
R865 drain_left.n46 drain_left.n8 12.8005
R866 drain_left.n117 drain_left.n79 12.8005
R867 drain_left.n112 drain_left.n83 12.8005
R868 drain_left.n39 drain_left.n12 12.0247
R869 drain_left.n50 drain_left.n49 12.0247
R870 drain_left.n121 drain_left.n120 12.0247
R871 drain_left.n111 drain_left.n84 12.0247
R872 drain_left.n36 drain_left.n35 11.249
R873 drain_left.n53 drain_left.n6 11.249
R874 drain_left.n124 drain_left.n77 11.249
R875 drain_left.n108 drain_left.n107 11.249
R876 drain_left.n32 drain_left.n14 10.4732
R877 drain_left.n54 drain_left.n4 10.4732
R878 drain_left.n125 drain_left.n75 10.4732
R879 drain_left.n104 drain_left.n86 10.4732
R880 drain_left.n21 drain_left.n20 10.2747
R881 drain_left.n93 drain_left.n92 10.2747
R882 drain_left.n31 drain_left.n16 9.69747
R883 drain_left.n58 drain_left.n57 9.69747
R884 drain_left.n129 drain_left.n128 9.69747
R885 drain_left.n103 drain_left.n88 9.69747
R886 drain_left.n64 drain_left.n63 9.45567
R887 drain_left.n135 drain_left.n134 9.45567
R888 drain_left.n63 drain_left.n62 9.3005
R889 drain_left.n2 drain_left.n1 9.3005
R890 drain_left.n57 drain_left.n56 9.3005
R891 drain_left.n55 drain_left.n54 9.3005
R892 drain_left.n6 drain_left.n5 9.3005
R893 drain_left.n49 drain_left.n48 9.3005
R894 drain_left.n47 drain_left.n46 9.3005
R895 drain_left.n23 drain_left.n22 9.3005
R896 drain_left.n18 drain_left.n17 9.3005
R897 drain_left.n29 drain_left.n28 9.3005
R898 drain_left.n31 drain_left.n30 9.3005
R899 drain_left.n14 drain_left.n13 9.3005
R900 drain_left.n37 drain_left.n36 9.3005
R901 drain_left.n39 drain_left.n38 9.3005
R902 drain_left.n40 drain_left.n9 9.3005
R903 drain_left.n95 drain_left.n94 9.3005
R904 drain_left.n90 drain_left.n89 9.3005
R905 drain_left.n101 drain_left.n100 9.3005
R906 drain_left.n103 drain_left.n102 9.3005
R907 drain_left.n86 drain_left.n85 9.3005
R908 drain_left.n109 drain_left.n108 9.3005
R909 drain_left.n111 drain_left.n110 9.3005
R910 drain_left.n83 drain_left.n80 9.3005
R911 drain_left.n134 drain_left.n133 9.3005
R912 drain_left.n73 drain_left.n72 9.3005
R913 drain_left.n128 drain_left.n127 9.3005
R914 drain_left.n126 drain_left.n125 9.3005
R915 drain_left.n77 drain_left.n76 9.3005
R916 drain_left.n120 drain_left.n119 9.3005
R917 drain_left.n118 drain_left.n117 9.3005
R918 drain_left.n28 drain_left.n27 8.92171
R919 drain_left.n61 drain_left.n2 8.92171
R920 drain_left.n132 drain_left.n73 8.92171
R921 drain_left.n100 drain_left.n99 8.92171
R922 drain_left.n24 drain_left.n18 8.14595
R923 drain_left.n62 drain_left.n0 8.14595
R924 drain_left.n133 drain_left.n71 8.14595
R925 drain_left.n96 drain_left.n90 8.14595
R926 drain_left.n23 drain_left.n20 7.3702
R927 drain_left.n95 drain_left.n92 7.3702
R928 drain_left drain_left.n141 6.11011
R929 drain_left.n24 drain_left.n23 5.81868
R930 drain_left.n64 drain_left.n0 5.81868
R931 drain_left.n135 drain_left.n71 5.81868
R932 drain_left.n96 drain_left.n95 5.81868
R933 drain_left.n27 drain_left.n18 5.04292
R934 drain_left.n62 drain_left.n61 5.04292
R935 drain_left.n133 drain_left.n132 5.04292
R936 drain_left.n99 drain_left.n90 5.04292
R937 drain_left.n28 drain_left.n16 4.26717
R938 drain_left.n58 drain_left.n2 4.26717
R939 drain_left.n129 drain_left.n73 4.26717
R940 drain_left.n100 drain_left.n88 4.26717
R941 drain_left.n32 drain_left.n31 3.49141
R942 drain_left.n57 drain_left.n4 3.49141
R943 drain_left.n128 drain_left.n75 3.49141
R944 drain_left.n104 drain_left.n103 3.49141
R945 drain_left.n22 drain_left.n21 2.84303
R946 drain_left.n94 drain_left.n93 2.84303
R947 drain_left.n35 drain_left.n14 2.71565
R948 drain_left.n54 drain_left.n53 2.71565
R949 drain_left.n125 drain_left.n124 2.71565
R950 drain_left.n107 drain_left.n86 2.71565
R951 drain_left.n36 drain_left.n12 1.93989
R952 drain_left.n50 drain_left.n6 1.93989
R953 drain_left.n121 drain_left.n77 1.93989
R954 drain_left.n108 drain_left.n84 1.93989
R955 drain_left.n67 drain_left.t0 1.6505
R956 drain_left.n67 drain_left.t2 1.6505
R957 drain_left.n68 drain_left.t8 1.6505
R958 drain_left.n68 drain_left.t4 1.6505
R959 drain_left.n65 drain_left.t9 1.6505
R960 drain_left.n65 drain_left.t3 1.6505
R961 drain_left.n140 drain_left.t11 1.6505
R962 drain_left.n140 drain_left.t13 1.6505
R963 drain_left.n138 drain_left.t6 1.6505
R964 drain_left.n138 drain_left.t7 1.6505
R965 drain_left.n136 drain_left.t12 1.6505
R966 drain_left.n136 drain_left.t1 1.6505
R967 drain_left.n41 drain_left.n39 1.16414
R968 drain_left.n49 drain_left.n8 1.16414
R969 drain_left.n120 drain_left.n79 1.16414
R970 drain_left.n112 drain_left.n111 1.16414
R971 drain_left.n139 drain_left.n137 0.457397
R972 drain_left.n141 drain_left.n139 0.457397
R973 drain_left.n40 drain_left.n10 0.388379
R974 drain_left.n46 drain_left.n45 0.388379
R975 drain_left.n117 drain_left.n116 0.388379
R976 drain_left.n83 drain_left.n81 0.388379
R977 drain_left.n70 drain_left.n66 0.287826
R978 drain_left.n22 drain_left.n17 0.155672
R979 drain_left.n29 drain_left.n17 0.155672
R980 drain_left.n30 drain_left.n29 0.155672
R981 drain_left.n30 drain_left.n13 0.155672
R982 drain_left.n37 drain_left.n13 0.155672
R983 drain_left.n38 drain_left.n37 0.155672
R984 drain_left.n38 drain_left.n9 0.155672
R985 drain_left.n47 drain_left.n9 0.155672
R986 drain_left.n48 drain_left.n47 0.155672
R987 drain_left.n48 drain_left.n5 0.155672
R988 drain_left.n55 drain_left.n5 0.155672
R989 drain_left.n56 drain_left.n55 0.155672
R990 drain_left.n56 drain_left.n1 0.155672
R991 drain_left.n63 drain_left.n1 0.155672
R992 drain_left.n134 drain_left.n72 0.155672
R993 drain_left.n127 drain_left.n72 0.155672
R994 drain_left.n127 drain_left.n126 0.155672
R995 drain_left.n126 drain_left.n76 0.155672
R996 drain_left.n119 drain_left.n76 0.155672
R997 drain_left.n119 drain_left.n118 0.155672
R998 drain_left.n118 drain_left.n80 0.155672
R999 drain_left.n110 drain_left.n80 0.155672
R1000 drain_left.n110 drain_left.n109 0.155672
R1001 drain_left.n109 drain_left.n85 0.155672
R1002 drain_left.n102 drain_left.n85 0.155672
R1003 drain_left.n102 drain_left.n101 0.155672
R1004 drain_left.n101 drain_left.n89 0.155672
R1005 drain_left.n94 drain_left.n89 0.155672
R1006 drain_left.n70 drain_left.n69 0.0593781
C0 source drain_right 33.4249f
C1 source drain_left 33.4367f
C2 minus plus 5.105f
C3 drain_right plus 0.30613f
C4 drain_left plus 4.12235f
C5 source plus 3.56581f
C6 minus drain_right 3.9753f
C7 minus drain_left 0.171065f
C8 source minus 3.55107f
C9 drain_left drain_right 0.795404f
C10 drain_right a_n1564_n3288# 7.535531f
C11 drain_left a_n1564_n3288# 7.79546f
C12 source a_n1564_n3288# 6.033535f
C13 minus a_n1564_n3288# 6.052875f
C14 plus a_n1564_n3288# 8.123601f
C15 drain_left.n0 a_n1564_n3288# 0.0461f
C16 drain_left.n1 a_n1564_n3288# 0.034803f
C17 drain_left.n2 a_n1564_n3288# 0.018701f
C18 drain_left.n3 a_n1564_n3288# 0.044203f
C19 drain_left.n4 a_n1564_n3288# 0.019802f
C20 drain_left.n5 a_n1564_n3288# 0.034803f
C21 drain_left.n6 a_n1564_n3288# 0.018701f
C22 drain_left.n7 a_n1564_n3288# 0.044203f
C23 drain_left.n8 a_n1564_n3288# 0.019802f
C24 drain_left.n9 a_n1564_n3288# 0.034803f
C25 drain_left.n10 a_n1564_n3288# 0.019251f
C26 drain_left.n11 a_n1564_n3288# 0.044203f
C27 drain_left.n12 a_n1564_n3288# 0.019802f
C28 drain_left.n13 a_n1564_n3288# 0.034803f
C29 drain_left.n14 a_n1564_n3288# 0.018701f
C30 drain_left.n15 a_n1564_n3288# 0.044203f
C31 drain_left.n16 a_n1564_n3288# 0.019802f
C32 drain_left.n17 a_n1564_n3288# 0.034803f
C33 drain_left.n18 a_n1564_n3288# 0.018701f
C34 drain_left.n19 a_n1564_n3288# 0.033152f
C35 drain_left.n20 a_n1564_n3288# 0.031248f
C36 drain_left.t5 a_n1564_n3288# 0.074656f
C37 drain_left.n21 a_n1564_n3288# 0.250922f
C38 drain_left.n22 a_n1564_n3288# 1.75573f
C39 drain_left.n23 a_n1564_n3288# 0.018701f
C40 drain_left.n24 a_n1564_n3288# 0.019802f
C41 drain_left.n25 a_n1564_n3288# 0.044203f
C42 drain_left.n26 a_n1564_n3288# 0.044203f
C43 drain_left.n27 a_n1564_n3288# 0.019802f
C44 drain_left.n28 a_n1564_n3288# 0.018701f
C45 drain_left.n29 a_n1564_n3288# 0.034803f
C46 drain_left.n30 a_n1564_n3288# 0.034803f
C47 drain_left.n31 a_n1564_n3288# 0.018701f
C48 drain_left.n32 a_n1564_n3288# 0.019802f
C49 drain_left.n33 a_n1564_n3288# 0.044203f
C50 drain_left.n34 a_n1564_n3288# 0.044203f
C51 drain_left.n35 a_n1564_n3288# 0.019802f
C52 drain_left.n36 a_n1564_n3288# 0.018701f
C53 drain_left.n37 a_n1564_n3288# 0.034803f
C54 drain_left.n38 a_n1564_n3288# 0.034803f
C55 drain_left.n39 a_n1564_n3288# 0.018701f
C56 drain_left.n40 a_n1564_n3288# 0.018701f
C57 drain_left.n41 a_n1564_n3288# 0.019802f
C58 drain_left.n42 a_n1564_n3288# 0.044203f
C59 drain_left.n43 a_n1564_n3288# 0.044203f
C60 drain_left.n44 a_n1564_n3288# 0.044203f
C61 drain_left.n45 a_n1564_n3288# 0.019251f
C62 drain_left.n46 a_n1564_n3288# 0.018701f
C63 drain_left.n47 a_n1564_n3288# 0.034803f
C64 drain_left.n48 a_n1564_n3288# 0.034803f
C65 drain_left.n49 a_n1564_n3288# 0.018701f
C66 drain_left.n50 a_n1564_n3288# 0.019802f
C67 drain_left.n51 a_n1564_n3288# 0.044203f
C68 drain_left.n52 a_n1564_n3288# 0.044203f
C69 drain_left.n53 a_n1564_n3288# 0.019802f
C70 drain_left.n54 a_n1564_n3288# 0.018701f
C71 drain_left.n55 a_n1564_n3288# 0.034803f
C72 drain_left.n56 a_n1564_n3288# 0.034803f
C73 drain_left.n57 a_n1564_n3288# 0.018701f
C74 drain_left.n58 a_n1564_n3288# 0.019802f
C75 drain_left.n59 a_n1564_n3288# 0.044203f
C76 drain_left.n60 a_n1564_n3288# 0.09071f
C77 drain_left.n61 a_n1564_n3288# 0.019802f
C78 drain_left.n62 a_n1564_n3288# 0.018701f
C79 drain_left.n63 a_n1564_n3288# 0.074739f
C80 drain_left.n64 a_n1564_n3288# 0.07526f
C81 drain_left.t9 a_n1564_n3288# 0.330024f
C82 drain_left.t3 a_n1564_n3288# 0.330024f
C83 drain_left.n65 a_n1564_n3288# 2.93671f
C84 drain_left.n66 a_n1564_n3288# 0.492219f
C85 drain_left.t0 a_n1564_n3288# 0.330024f
C86 drain_left.t2 a_n1564_n3288# 0.330024f
C87 drain_left.n67 a_n1564_n3288# 2.93982f
C88 drain_left.t8 a_n1564_n3288# 0.330024f
C89 drain_left.t4 a_n1564_n3288# 0.330024f
C90 drain_left.n68 a_n1564_n3288# 2.93671f
C91 drain_left.n69 a_n1564_n3288# 0.76909f
C92 drain_left.n70 a_n1564_n3288# 1.58617f
C93 drain_left.n71 a_n1564_n3288# 0.0461f
C94 drain_left.n72 a_n1564_n3288# 0.034803f
C95 drain_left.n73 a_n1564_n3288# 0.018701f
C96 drain_left.n74 a_n1564_n3288# 0.044203f
C97 drain_left.n75 a_n1564_n3288# 0.019802f
C98 drain_left.n76 a_n1564_n3288# 0.034803f
C99 drain_left.n77 a_n1564_n3288# 0.018701f
C100 drain_left.n78 a_n1564_n3288# 0.044203f
C101 drain_left.n79 a_n1564_n3288# 0.019802f
C102 drain_left.n80 a_n1564_n3288# 0.034803f
C103 drain_left.n81 a_n1564_n3288# 0.019251f
C104 drain_left.n82 a_n1564_n3288# 0.044203f
C105 drain_left.n83 a_n1564_n3288# 0.018701f
C106 drain_left.n84 a_n1564_n3288# 0.019802f
C107 drain_left.n85 a_n1564_n3288# 0.034803f
C108 drain_left.n86 a_n1564_n3288# 0.018701f
C109 drain_left.n87 a_n1564_n3288# 0.044203f
C110 drain_left.n88 a_n1564_n3288# 0.019802f
C111 drain_left.n89 a_n1564_n3288# 0.034803f
C112 drain_left.n90 a_n1564_n3288# 0.018701f
C113 drain_left.n91 a_n1564_n3288# 0.033152f
C114 drain_left.n92 a_n1564_n3288# 0.031248f
C115 drain_left.t10 a_n1564_n3288# 0.074656f
C116 drain_left.n93 a_n1564_n3288# 0.250922f
C117 drain_left.n94 a_n1564_n3288# 1.75573f
C118 drain_left.n95 a_n1564_n3288# 0.018701f
C119 drain_left.n96 a_n1564_n3288# 0.019802f
C120 drain_left.n97 a_n1564_n3288# 0.044203f
C121 drain_left.n98 a_n1564_n3288# 0.044203f
C122 drain_left.n99 a_n1564_n3288# 0.019802f
C123 drain_left.n100 a_n1564_n3288# 0.018701f
C124 drain_left.n101 a_n1564_n3288# 0.034803f
C125 drain_left.n102 a_n1564_n3288# 0.034803f
C126 drain_left.n103 a_n1564_n3288# 0.018701f
C127 drain_left.n104 a_n1564_n3288# 0.019802f
C128 drain_left.n105 a_n1564_n3288# 0.044203f
C129 drain_left.n106 a_n1564_n3288# 0.044203f
C130 drain_left.n107 a_n1564_n3288# 0.019802f
C131 drain_left.n108 a_n1564_n3288# 0.018701f
C132 drain_left.n109 a_n1564_n3288# 0.034803f
C133 drain_left.n110 a_n1564_n3288# 0.034803f
C134 drain_left.n111 a_n1564_n3288# 0.018701f
C135 drain_left.n112 a_n1564_n3288# 0.019802f
C136 drain_left.n113 a_n1564_n3288# 0.044203f
C137 drain_left.n114 a_n1564_n3288# 0.044203f
C138 drain_left.n115 a_n1564_n3288# 0.044203f
C139 drain_left.n116 a_n1564_n3288# 0.019251f
C140 drain_left.n117 a_n1564_n3288# 0.018701f
C141 drain_left.n118 a_n1564_n3288# 0.034803f
C142 drain_left.n119 a_n1564_n3288# 0.034803f
C143 drain_left.n120 a_n1564_n3288# 0.018701f
C144 drain_left.n121 a_n1564_n3288# 0.019802f
C145 drain_left.n122 a_n1564_n3288# 0.044203f
C146 drain_left.n123 a_n1564_n3288# 0.044203f
C147 drain_left.n124 a_n1564_n3288# 0.019802f
C148 drain_left.n125 a_n1564_n3288# 0.018701f
C149 drain_left.n126 a_n1564_n3288# 0.034803f
C150 drain_left.n127 a_n1564_n3288# 0.034803f
C151 drain_left.n128 a_n1564_n3288# 0.018701f
C152 drain_left.n129 a_n1564_n3288# 0.019802f
C153 drain_left.n130 a_n1564_n3288# 0.044203f
C154 drain_left.n131 a_n1564_n3288# 0.09071f
C155 drain_left.n132 a_n1564_n3288# 0.019802f
C156 drain_left.n133 a_n1564_n3288# 0.018701f
C157 drain_left.n134 a_n1564_n3288# 0.074739f
C158 drain_left.n135 a_n1564_n3288# 0.07526f
C159 drain_left.t12 a_n1564_n3288# 0.330024f
C160 drain_left.t1 a_n1564_n3288# 0.330024f
C161 drain_left.n136 a_n1564_n3288# 2.93672f
C162 drain_left.n137 a_n1564_n3288# 0.508415f
C163 drain_left.t6 a_n1564_n3288# 0.330024f
C164 drain_left.t7 a_n1564_n3288# 0.330024f
C165 drain_left.n138 a_n1564_n3288# 2.93672f
C166 drain_left.n139 a_n1564_n3288# 0.394545f
C167 drain_left.t11 a_n1564_n3288# 0.330024f
C168 drain_left.t13 a_n1564_n3288# 0.330024f
C169 drain_left.n140 a_n1564_n3288# 2.93671f
C170 drain_left.n141 a_n1564_n3288# 0.679383f
C171 plus.n0 a_n1564_n3288# 0.056074f
C172 plus.t2 a_n1564_n3288# 0.380292f
C173 plus.t6 a_n1564_n3288# 0.380292f
C174 plus.t7 a_n1564_n3288# 0.380292f
C175 plus.n1 a_n1564_n3288# 0.156622f
C176 plus.n2 a_n1564_n3288# 0.125204f
C177 plus.t12 a_n1564_n3288# 0.380292f
C178 plus.t1 a_n1564_n3288# 0.380292f
C179 plus.t3 a_n1564_n3288# 0.385041f
C180 plus.n3 a_n1564_n3288# 0.172976f
C181 plus.n4 a_n1564_n3288# 0.156622f
C182 plus.n5 a_n1564_n3288# 0.019639f
C183 plus.n6 a_n1564_n3288# 0.156622f
C184 plus.n7 a_n1564_n3288# 0.019639f
C185 plus.n8 a_n1564_n3288# 0.056074f
C186 plus.n9 a_n1564_n3288# 0.056074f
C187 plus.n10 a_n1564_n3288# 0.019639f
C188 plus.n11 a_n1564_n3288# 0.156622f
C189 plus.n12 a_n1564_n3288# 0.019639f
C190 plus.n13 a_n1564_n3288# 0.156622f
C191 plus.t0 a_n1564_n3288# 0.385041f
C192 plus.n14 a_n1564_n3288# 0.172894f
C193 plus.n15 a_n1564_n3288# 0.622111f
C194 plus.n16 a_n1564_n3288# 0.056074f
C195 plus.t8 a_n1564_n3288# 0.385041f
C196 plus.t4 a_n1564_n3288# 0.380292f
C197 plus.t10 a_n1564_n3288# 0.380292f
C198 plus.t5 a_n1564_n3288# 0.380292f
C199 plus.n17 a_n1564_n3288# 0.156622f
C200 plus.n18 a_n1564_n3288# 0.125204f
C201 plus.t9 a_n1564_n3288# 0.380292f
C202 plus.t13 a_n1564_n3288# 0.380292f
C203 plus.t11 a_n1564_n3288# 0.385041f
C204 plus.n19 a_n1564_n3288# 0.172976f
C205 plus.n20 a_n1564_n3288# 0.156622f
C206 plus.n21 a_n1564_n3288# 0.019639f
C207 plus.n22 a_n1564_n3288# 0.156622f
C208 plus.n23 a_n1564_n3288# 0.019639f
C209 plus.n24 a_n1564_n3288# 0.056074f
C210 plus.n25 a_n1564_n3288# 0.056074f
C211 plus.n26 a_n1564_n3288# 0.019639f
C212 plus.n27 a_n1564_n3288# 0.156622f
C213 plus.n28 a_n1564_n3288# 0.019639f
C214 plus.n29 a_n1564_n3288# 0.156622f
C215 plus.n30 a_n1564_n3288# 0.172894f
C216 plus.n31 a_n1564_n3288# 1.58428f
C217 drain_right.n0 a_n1564_n3288# 0.046145f
C218 drain_right.n1 a_n1564_n3288# 0.034836f
C219 drain_right.n2 a_n1564_n3288# 0.018719f
C220 drain_right.n3 a_n1564_n3288# 0.044246f
C221 drain_right.n4 a_n1564_n3288# 0.019821f
C222 drain_right.n5 a_n1564_n3288# 0.034836f
C223 drain_right.n6 a_n1564_n3288# 0.018719f
C224 drain_right.n7 a_n1564_n3288# 0.044246f
C225 drain_right.n8 a_n1564_n3288# 0.019821f
C226 drain_right.n9 a_n1564_n3288# 0.034836f
C227 drain_right.n10 a_n1564_n3288# 0.01927f
C228 drain_right.n11 a_n1564_n3288# 0.044246f
C229 drain_right.n12 a_n1564_n3288# 0.019821f
C230 drain_right.n13 a_n1564_n3288# 0.034836f
C231 drain_right.n14 a_n1564_n3288# 0.018719f
C232 drain_right.n15 a_n1564_n3288# 0.044246f
C233 drain_right.n16 a_n1564_n3288# 0.019821f
C234 drain_right.n17 a_n1564_n3288# 0.034836f
C235 drain_right.n18 a_n1564_n3288# 0.018719f
C236 drain_right.n19 a_n1564_n3288# 0.033185f
C237 drain_right.n20 a_n1564_n3288# 0.031278f
C238 drain_right.t10 a_n1564_n3288# 0.074729f
C239 drain_right.n21 a_n1564_n3288# 0.251165f
C240 drain_right.n22 a_n1564_n3288# 1.75743f
C241 drain_right.n23 a_n1564_n3288# 0.018719f
C242 drain_right.n24 a_n1564_n3288# 0.019821f
C243 drain_right.n25 a_n1564_n3288# 0.044246f
C244 drain_right.n26 a_n1564_n3288# 0.044246f
C245 drain_right.n27 a_n1564_n3288# 0.019821f
C246 drain_right.n28 a_n1564_n3288# 0.018719f
C247 drain_right.n29 a_n1564_n3288# 0.034836f
C248 drain_right.n30 a_n1564_n3288# 0.034836f
C249 drain_right.n31 a_n1564_n3288# 0.018719f
C250 drain_right.n32 a_n1564_n3288# 0.019821f
C251 drain_right.n33 a_n1564_n3288# 0.044246f
C252 drain_right.n34 a_n1564_n3288# 0.044246f
C253 drain_right.n35 a_n1564_n3288# 0.019821f
C254 drain_right.n36 a_n1564_n3288# 0.018719f
C255 drain_right.n37 a_n1564_n3288# 0.034836f
C256 drain_right.n38 a_n1564_n3288# 0.034836f
C257 drain_right.n39 a_n1564_n3288# 0.018719f
C258 drain_right.n40 a_n1564_n3288# 0.018719f
C259 drain_right.n41 a_n1564_n3288# 0.019821f
C260 drain_right.n42 a_n1564_n3288# 0.044246f
C261 drain_right.n43 a_n1564_n3288# 0.044246f
C262 drain_right.n44 a_n1564_n3288# 0.044246f
C263 drain_right.n45 a_n1564_n3288# 0.01927f
C264 drain_right.n46 a_n1564_n3288# 0.018719f
C265 drain_right.n47 a_n1564_n3288# 0.034836f
C266 drain_right.n48 a_n1564_n3288# 0.034836f
C267 drain_right.n49 a_n1564_n3288# 0.018719f
C268 drain_right.n50 a_n1564_n3288# 0.019821f
C269 drain_right.n51 a_n1564_n3288# 0.044246f
C270 drain_right.n52 a_n1564_n3288# 0.044246f
C271 drain_right.n53 a_n1564_n3288# 0.019821f
C272 drain_right.n54 a_n1564_n3288# 0.018719f
C273 drain_right.n55 a_n1564_n3288# 0.034836f
C274 drain_right.n56 a_n1564_n3288# 0.034836f
C275 drain_right.n57 a_n1564_n3288# 0.018719f
C276 drain_right.n58 a_n1564_n3288# 0.019821f
C277 drain_right.n59 a_n1564_n3288# 0.044246f
C278 drain_right.n60 a_n1564_n3288# 0.090797f
C279 drain_right.n61 a_n1564_n3288# 0.019821f
C280 drain_right.n62 a_n1564_n3288# 0.018719f
C281 drain_right.n63 a_n1564_n3288# 0.074811f
C282 drain_right.n64 a_n1564_n3288# 0.075333f
C283 drain_right.t8 a_n1564_n3288# 0.330344f
C284 drain_right.t11 a_n1564_n3288# 0.330344f
C285 drain_right.n65 a_n1564_n3288# 2.93955f
C286 drain_right.n66 a_n1564_n3288# 0.492695f
C287 drain_right.t7 a_n1564_n3288# 0.330344f
C288 drain_right.t4 a_n1564_n3288# 0.330344f
C289 drain_right.n67 a_n1564_n3288# 2.94266f
C290 drain_right.t9 a_n1564_n3288# 0.330344f
C291 drain_right.t3 a_n1564_n3288# 0.330344f
C292 drain_right.n68 a_n1564_n3288# 2.93955f
C293 drain_right.n69 a_n1564_n3288# 0.769834f
C294 drain_right.n70 a_n1564_n3288# 1.51509f
C295 drain_right.t5 a_n1564_n3288# 0.330344f
C296 drain_right.t2 a_n1564_n3288# 0.330344f
C297 drain_right.n71 a_n1564_n3288# 2.94266f
C298 drain_right.t0 a_n1564_n3288# 0.330344f
C299 drain_right.t13 a_n1564_n3288# 0.330344f
C300 drain_right.n72 a_n1564_n3288# 2.93956f
C301 drain_right.n73 a_n1564_n3288# 0.800782f
C302 drain_right.t6 a_n1564_n3288# 0.330344f
C303 drain_right.t1 a_n1564_n3288# 0.330344f
C304 drain_right.n74 a_n1564_n3288# 2.93956f
C305 drain_right.n75 a_n1564_n3288# 0.394926f
C306 drain_right.n76 a_n1564_n3288# 0.046145f
C307 drain_right.n77 a_n1564_n3288# 0.034836f
C308 drain_right.n78 a_n1564_n3288# 0.018719f
C309 drain_right.n79 a_n1564_n3288# 0.044246f
C310 drain_right.n80 a_n1564_n3288# 0.019821f
C311 drain_right.n81 a_n1564_n3288# 0.034836f
C312 drain_right.n82 a_n1564_n3288# 0.018719f
C313 drain_right.n83 a_n1564_n3288# 0.044246f
C314 drain_right.n84 a_n1564_n3288# 0.019821f
C315 drain_right.n85 a_n1564_n3288# 0.034836f
C316 drain_right.n86 a_n1564_n3288# 0.01927f
C317 drain_right.n87 a_n1564_n3288# 0.044246f
C318 drain_right.n88 a_n1564_n3288# 0.018719f
C319 drain_right.n89 a_n1564_n3288# 0.019821f
C320 drain_right.n90 a_n1564_n3288# 0.034836f
C321 drain_right.n91 a_n1564_n3288# 0.018719f
C322 drain_right.n92 a_n1564_n3288# 0.044246f
C323 drain_right.n93 a_n1564_n3288# 0.019821f
C324 drain_right.n94 a_n1564_n3288# 0.034836f
C325 drain_right.n95 a_n1564_n3288# 0.018719f
C326 drain_right.n96 a_n1564_n3288# 0.033185f
C327 drain_right.n97 a_n1564_n3288# 0.031278f
C328 drain_right.t12 a_n1564_n3288# 0.074729f
C329 drain_right.n98 a_n1564_n3288# 0.251165f
C330 drain_right.n99 a_n1564_n3288# 1.75743f
C331 drain_right.n100 a_n1564_n3288# 0.018719f
C332 drain_right.n101 a_n1564_n3288# 0.019821f
C333 drain_right.n102 a_n1564_n3288# 0.044246f
C334 drain_right.n103 a_n1564_n3288# 0.044246f
C335 drain_right.n104 a_n1564_n3288# 0.019821f
C336 drain_right.n105 a_n1564_n3288# 0.018719f
C337 drain_right.n106 a_n1564_n3288# 0.034836f
C338 drain_right.n107 a_n1564_n3288# 0.034836f
C339 drain_right.n108 a_n1564_n3288# 0.018719f
C340 drain_right.n109 a_n1564_n3288# 0.019821f
C341 drain_right.n110 a_n1564_n3288# 0.044246f
C342 drain_right.n111 a_n1564_n3288# 0.044246f
C343 drain_right.n112 a_n1564_n3288# 0.019821f
C344 drain_right.n113 a_n1564_n3288# 0.018719f
C345 drain_right.n114 a_n1564_n3288# 0.034836f
C346 drain_right.n115 a_n1564_n3288# 0.034836f
C347 drain_right.n116 a_n1564_n3288# 0.018719f
C348 drain_right.n117 a_n1564_n3288# 0.019821f
C349 drain_right.n118 a_n1564_n3288# 0.044246f
C350 drain_right.n119 a_n1564_n3288# 0.044246f
C351 drain_right.n120 a_n1564_n3288# 0.044246f
C352 drain_right.n121 a_n1564_n3288# 0.01927f
C353 drain_right.n122 a_n1564_n3288# 0.018719f
C354 drain_right.n123 a_n1564_n3288# 0.034836f
C355 drain_right.n124 a_n1564_n3288# 0.034836f
C356 drain_right.n125 a_n1564_n3288# 0.018719f
C357 drain_right.n126 a_n1564_n3288# 0.019821f
C358 drain_right.n127 a_n1564_n3288# 0.044246f
C359 drain_right.n128 a_n1564_n3288# 0.044246f
C360 drain_right.n129 a_n1564_n3288# 0.019821f
C361 drain_right.n130 a_n1564_n3288# 0.018719f
C362 drain_right.n131 a_n1564_n3288# 0.034836f
C363 drain_right.n132 a_n1564_n3288# 0.034836f
C364 drain_right.n133 a_n1564_n3288# 0.018719f
C365 drain_right.n134 a_n1564_n3288# 0.019821f
C366 drain_right.n135 a_n1564_n3288# 0.044246f
C367 drain_right.n136 a_n1564_n3288# 0.090797f
C368 drain_right.n137 a_n1564_n3288# 0.019821f
C369 drain_right.n138 a_n1564_n3288# 0.018719f
C370 drain_right.n139 a_n1564_n3288# 0.074811f
C371 drain_right.n140 a_n1564_n3288# 0.074214f
C372 drain_right.n141 a_n1564_n3288# 0.39824f
C373 source.n0 a_n1564_n3288# 0.047675f
C374 source.n1 a_n1564_n3288# 0.035991f
C375 source.n2 a_n1564_n3288# 0.01934f
C376 source.n3 a_n1564_n3288# 0.045713f
C377 source.n4 a_n1564_n3288# 0.020478f
C378 source.n5 a_n1564_n3288# 0.035991f
C379 source.n6 a_n1564_n3288# 0.01934f
C380 source.n7 a_n1564_n3288# 0.045713f
C381 source.n8 a_n1564_n3288# 0.020478f
C382 source.n9 a_n1564_n3288# 0.035991f
C383 source.n10 a_n1564_n3288# 0.019909f
C384 source.n11 a_n1564_n3288# 0.045713f
C385 source.n12 a_n1564_n3288# 0.01934f
C386 source.n13 a_n1564_n3288# 0.020478f
C387 source.n14 a_n1564_n3288# 0.035991f
C388 source.n15 a_n1564_n3288# 0.01934f
C389 source.n16 a_n1564_n3288# 0.045713f
C390 source.n17 a_n1564_n3288# 0.020478f
C391 source.n18 a_n1564_n3288# 0.035991f
C392 source.n19 a_n1564_n3288# 0.01934f
C393 source.n20 a_n1564_n3288# 0.034284f
C394 source.n21 a_n1564_n3288# 0.032315f
C395 source.t7 a_n1564_n3288# 0.077206f
C396 source.n22 a_n1564_n3288# 0.259491f
C397 source.n23 a_n1564_n3288# 1.81568f
C398 source.n24 a_n1564_n3288# 0.01934f
C399 source.n25 a_n1564_n3288# 0.020478f
C400 source.n26 a_n1564_n3288# 0.045713f
C401 source.n27 a_n1564_n3288# 0.045713f
C402 source.n28 a_n1564_n3288# 0.020478f
C403 source.n29 a_n1564_n3288# 0.01934f
C404 source.n30 a_n1564_n3288# 0.035991f
C405 source.n31 a_n1564_n3288# 0.035991f
C406 source.n32 a_n1564_n3288# 0.01934f
C407 source.n33 a_n1564_n3288# 0.020478f
C408 source.n34 a_n1564_n3288# 0.045713f
C409 source.n35 a_n1564_n3288# 0.045713f
C410 source.n36 a_n1564_n3288# 0.020478f
C411 source.n37 a_n1564_n3288# 0.01934f
C412 source.n38 a_n1564_n3288# 0.035991f
C413 source.n39 a_n1564_n3288# 0.035991f
C414 source.n40 a_n1564_n3288# 0.01934f
C415 source.n41 a_n1564_n3288# 0.020478f
C416 source.n42 a_n1564_n3288# 0.045713f
C417 source.n43 a_n1564_n3288# 0.045713f
C418 source.n44 a_n1564_n3288# 0.045713f
C419 source.n45 a_n1564_n3288# 0.019909f
C420 source.n46 a_n1564_n3288# 0.01934f
C421 source.n47 a_n1564_n3288# 0.035991f
C422 source.n48 a_n1564_n3288# 0.035991f
C423 source.n49 a_n1564_n3288# 0.01934f
C424 source.n50 a_n1564_n3288# 0.020478f
C425 source.n51 a_n1564_n3288# 0.045713f
C426 source.n52 a_n1564_n3288# 0.045713f
C427 source.n53 a_n1564_n3288# 0.020478f
C428 source.n54 a_n1564_n3288# 0.01934f
C429 source.n55 a_n1564_n3288# 0.035991f
C430 source.n56 a_n1564_n3288# 0.035991f
C431 source.n57 a_n1564_n3288# 0.01934f
C432 source.n58 a_n1564_n3288# 0.020478f
C433 source.n59 a_n1564_n3288# 0.045713f
C434 source.n60 a_n1564_n3288# 0.093807f
C435 source.n61 a_n1564_n3288# 0.020478f
C436 source.n62 a_n1564_n3288# 0.01934f
C437 source.n63 a_n1564_n3288# 0.077291f
C438 source.n64 a_n1564_n3288# 0.051771f
C439 source.n65 a_n1564_n3288# 1.43205f
C440 source.t9 a_n1564_n3288# 0.341294f
C441 source.t1 a_n1564_n3288# 0.341294f
C442 source.n66 a_n1564_n3288# 2.92217f
C443 source.n67 a_n1564_n3288# 0.473935f
C444 source.t5 a_n1564_n3288# 0.341294f
C445 source.t0 a_n1564_n3288# 0.341294f
C446 source.n68 a_n1564_n3288# 2.92217f
C447 source.n69 a_n1564_n3288# 0.473935f
C448 source.t3 a_n1564_n3288# 0.341294f
C449 source.t2 a_n1564_n3288# 0.341294f
C450 source.n70 a_n1564_n3288# 2.92217f
C451 source.n71 a_n1564_n3288# 0.501928f
C452 source.n72 a_n1564_n3288# 0.047675f
C453 source.n73 a_n1564_n3288# 0.035991f
C454 source.n74 a_n1564_n3288# 0.01934f
C455 source.n75 a_n1564_n3288# 0.045713f
C456 source.n76 a_n1564_n3288# 0.020478f
C457 source.n77 a_n1564_n3288# 0.035991f
C458 source.n78 a_n1564_n3288# 0.01934f
C459 source.n79 a_n1564_n3288# 0.045713f
C460 source.n80 a_n1564_n3288# 0.020478f
C461 source.n81 a_n1564_n3288# 0.035991f
C462 source.n82 a_n1564_n3288# 0.019909f
C463 source.n83 a_n1564_n3288# 0.045713f
C464 source.n84 a_n1564_n3288# 0.01934f
C465 source.n85 a_n1564_n3288# 0.020478f
C466 source.n86 a_n1564_n3288# 0.035991f
C467 source.n87 a_n1564_n3288# 0.01934f
C468 source.n88 a_n1564_n3288# 0.045713f
C469 source.n89 a_n1564_n3288# 0.020478f
C470 source.n90 a_n1564_n3288# 0.035991f
C471 source.n91 a_n1564_n3288# 0.01934f
C472 source.n92 a_n1564_n3288# 0.034284f
C473 source.n93 a_n1564_n3288# 0.032315f
C474 source.t16 a_n1564_n3288# 0.077206f
C475 source.n94 a_n1564_n3288# 0.259491f
C476 source.n95 a_n1564_n3288# 1.81568f
C477 source.n96 a_n1564_n3288# 0.01934f
C478 source.n97 a_n1564_n3288# 0.020478f
C479 source.n98 a_n1564_n3288# 0.045713f
C480 source.n99 a_n1564_n3288# 0.045713f
C481 source.n100 a_n1564_n3288# 0.020478f
C482 source.n101 a_n1564_n3288# 0.01934f
C483 source.n102 a_n1564_n3288# 0.035991f
C484 source.n103 a_n1564_n3288# 0.035991f
C485 source.n104 a_n1564_n3288# 0.01934f
C486 source.n105 a_n1564_n3288# 0.020478f
C487 source.n106 a_n1564_n3288# 0.045713f
C488 source.n107 a_n1564_n3288# 0.045713f
C489 source.n108 a_n1564_n3288# 0.020478f
C490 source.n109 a_n1564_n3288# 0.01934f
C491 source.n110 a_n1564_n3288# 0.035991f
C492 source.n111 a_n1564_n3288# 0.035991f
C493 source.n112 a_n1564_n3288# 0.01934f
C494 source.n113 a_n1564_n3288# 0.020478f
C495 source.n114 a_n1564_n3288# 0.045713f
C496 source.n115 a_n1564_n3288# 0.045713f
C497 source.n116 a_n1564_n3288# 0.045713f
C498 source.n117 a_n1564_n3288# 0.019909f
C499 source.n118 a_n1564_n3288# 0.01934f
C500 source.n119 a_n1564_n3288# 0.035991f
C501 source.n120 a_n1564_n3288# 0.035991f
C502 source.n121 a_n1564_n3288# 0.01934f
C503 source.n122 a_n1564_n3288# 0.020478f
C504 source.n123 a_n1564_n3288# 0.045713f
C505 source.n124 a_n1564_n3288# 0.045713f
C506 source.n125 a_n1564_n3288# 0.020478f
C507 source.n126 a_n1564_n3288# 0.01934f
C508 source.n127 a_n1564_n3288# 0.035991f
C509 source.n128 a_n1564_n3288# 0.035991f
C510 source.n129 a_n1564_n3288# 0.01934f
C511 source.n130 a_n1564_n3288# 0.020478f
C512 source.n131 a_n1564_n3288# 0.045713f
C513 source.n132 a_n1564_n3288# 0.093807f
C514 source.n133 a_n1564_n3288# 0.020478f
C515 source.n134 a_n1564_n3288# 0.01934f
C516 source.n135 a_n1564_n3288# 0.077291f
C517 source.n136 a_n1564_n3288# 0.051771f
C518 source.n137 a_n1564_n3288# 0.161382f
C519 source.t26 a_n1564_n3288# 0.341294f
C520 source.t14 a_n1564_n3288# 0.341294f
C521 source.n138 a_n1564_n3288# 2.92217f
C522 source.n139 a_n1564_n3288# 0.473935f
C523 source.t23 a_n1564_n3288# 0.341294f
C524 source.t21 a_n1564_n3288# 0.341294f
C525 source.n140 a_n1564_n3288# 2.92217f
C526 source.n141 a_n1564_n3288# 0.473935f
C527 source.t24 a_n1564_n3288# 0.341294f
C528 source.t17 a_n1564_n3288# 0.341294f
C529 source.n142 a_n1564_n3288# 2.92217f
C530 source.n143 a_n1564_n3288# 2.38792f
C531 source.t11 a_n1564_n3288# 0.341294f
C532 source.t6 a_n1564_n3288# 0.341294f
C533 source.n144 a_n1564_n3288# 2.92215f
C534 source.n145 a_n1564_n3288# 2.38794f
C535 source.t10 a_n1564_n3288# 0.341294f
C536 source.t8 a_n1564_n3288# 0.341294f
C537 source.n146 a_n1564_n3288# 2.92215f
C538 source.n147 a_n1564_n3288# 0.473953f
C539 source.t4 a_n1564_n3288# 0.341294f
C540 source.t12 a_n1564_n3288# 0.341294f
C541 source.n148 a_n1564_n3288# 2.92215f
C542 source.n149 a_n1564_n3288# 0.473953f
C543 source.n150 a_n1564_n3288# 0.047675f
C544 source.n151 a_n1564_n3288# 0.035991f
C545 source.n152 a_n1564_n3288# 0.01934f
C546 source.n153 a_n1564_n3288# 0.045713f
C547 source.n154 a_n1564_n3288# 0.020478f
C548 source.n155 a_n1564_n3288# 0.035991f
C549 source.n156 a_n1564_n3288# 0.01934f
C550 source.n157 a_n1564_n3288# 0.045713f
C551 source.n158 a_n1564_n3288# 0.020478f
C552 source.n159 a_n1564_n3288# 0.035991f
C553 source.n160 a_n1564_n3288# 0.019909f
C554 source.n161 a_n1564_n3288# 0.045713f
C555 source.n162 a_n1564_n3288# 0.020478f
C556 source.n163 a_n1564_n3288# 0.035991f
C557 source.n164 a_n1564_n3288# 0.01934f
C558 source.n165 a_n1564_n3288# 0.045713f
C559 source.n166 a_n1564_n3288# 0.020478f
C560 source.n167 a_n1564_n3288# 0.035991f
C561 source.n168 a_n1564_n3288# 0.01934f
C562 source.n169 a_n1564_n3288# 0.034284f
C563 source.n170 a_n1564_n3288# 0.032315f
C564 source.t13 a_n1564_n3288# 0.077206f
C565 source.n171 a_n1564_n3288# 0.259491f
C566 source.n172 a_n1564_n3288# 1.81568f
C567 source.n173 a_n1564_n3288# 0.01934f
C568 source.n174 a_n1564_n3288# 0.020478f
C569 source.n175 a_n1564_n3288# 0.045713f
C570 source.n176 a_n1564_n3288# 0.045713f
C571 source.n177 a_n1564_n3288# 0.020478f
C572 source.n178 a_n1564_n3288# 0.01934f
C573 source.n179 a_n1564_n3288# 0.035991f
C574 source.n180 a_n1564_n3288# 0.035991f
C575 source.n181 a_n1564_n3288# 0.01934f
C576 source.n182 a_n1564_n3288# 0.020478f
C577 source.n183 a_n1564_n3288# 0.045713f
C578 source.n184 a_n1564_n3288# 0.045713f
C579 source.n185 a_n1564_n3288# 0.020478f
C580 source.n186 a_n1564_n3288# 0.01934f
C581 source.n187 a_n1564_n3288# 0.035991f
C582 source.n188 a_n1564_n3288# 0.035991f
C583 source.n189 a_n1564_n3288# 0.01934f
C584 source.n190 a_n1564_n3288# 0.01934f
C585 source.n191 a_n1564_n3288# 0.020478f
C586 source.n192 a_n1564_n3288# 0.045713f
C587 source.n193 a_n1564_n3288# 0.045713f
C588 source.n194 a_n1564_n3288# 0.045713f
C589 source.n195 a_n1564_n3288# 0.019909f
C590 source.n196 a_n1564_n3288# 0.01934f
C591 source.n197 a_n1564_n3288# 0.035991f
C592 source.n198 a_n1564_n3288# 0.035991f
C593 source.n199 a_n1564_n3288# 0.01934f
C594 source.n200 a_n1564_n3288# 0.020478f
C595 source.n201 a_n1564_n3288# 0.045713f
C596 source.n202 a_n1564_n3288# 0.045713f
C597 source.n203 a_n1564_n3288# 0.020478f
C598 source.n204 a_n1564_n3288# 0.01934f
C599 source.n205 a_n1564_n3288# 0.035991f
C600 source.n206 a_n1564_n3288# 0.035991f
C601 source.n207 a_n1564_n3288# 0.01934f
C602 source.n208 a_n1564_n3288# 0.020478f
C603 source.n209 a_n1564_n3288# 0.045713f
C604 source.n210 a_n1564_n3288# 0.093807f
C605 source.n211 a_n1564_n3288# 0.020478f
C606 source.n212 a_n1564_n3288# 0.01934f
C607 source.n213 a_n1564_n3288# 0.077291f
C608 source.n214 a_n1564_n3288# 0.051771f
C609 source.n215 a_n1564_n3288# 0.161382f
C610 source.t19 a_n1564_n3288# 0.341294f
C611 source.t27 a_n1564_n3288# 0.341294f
C612 source.n216 a_n1564_n3288# 2.92215f
C613 source.n217 a_n1564_n3288# 0.501946f
C614 source.t22 a_n1564_n3288# 0.341294f
C615 source.t18 a_n1564_n3288# 0.341294f
C616 source.n218 a_n1564_n3288# 2.92215f
C617 source.n219 a_n1564_n3288# 0.473953f
C618 source.t15 a_n1564_n3288# 0.341294f
C619 source.t25 a_n1564_n3288# 0.341294f
C620 source.n220 a_n1564_n3288# 2.92215f
C621 source.n221 a_n1564_n3288# 0.473953f
C622 source.n222 a_n1564_n3288# 0.047675f
C623 source.n223 a_n1564_n3288# 0.035991f
C624 source.n224 a_n1564_n3288# 0.01934f
C625 source.n225 a_n1564_n3288# 0.045713f
C626 source.n226 a_n1564_n3288# 0.020478f
C627 source.n227 a_n1564_n3288# 0.035991f
C628 source.n228 a_n1564_n3288# 0.01934f
C629 source.n229 a_n1564_n3288# 0.045713f
C630 source.n230 a_n1564_n3288# 0.020478f
C631 source.n231 a_n1564_n3288# 0.035991f
C632 source.n232 a_n1564_n3288# 0.019909f
C633 source.n233 a_n1564_n3288# 0.045713f
C634 source.n234 a_n1564_n3288# 0.020478f
C635 source.n235 a_n1564_n3288# 0.035991f
C636 source.n236 a_n1564_n3288# 0.01934f
C637 source.n237 a_n1564_n3288# 0.045713f
C638 source.n238 a_n1564_n3288# 0.020478f
C639 source.n239 a_n1564_n3288# 0.035991f
C640 source.n240 a_n1564_n3288# 0.01934f
C641 source.n241 a_n1564_n3288# 0.034284f
C642 source.n242 a_n1564_n3288# 0.032315f
C643 source.t20 a_n1564_n3288# 0.077206f
C644 source.n243 a_n1564_n3288# 0.259491f
C645 source.n244 a_n1564_n3288# 1.81568f
C646 source.n245 a_n1564_n3288# 0.01934f
C647 source.n246 a_n1564_n3288# 0.020478f
C648 source.n247 a_n1564_n3288# 0.045713f
C649 source.n248 a_n1564_n3288# 0.045713f
C650 source.n249 a_n1564_n3288# 0.020478f
C651 source.n250 a_n1564_n3288# 0.01934f
C652 source.n251 a_n1564_n3288# 0.035991f
C653 source.n252 a_n1564_n3288# 0.035991f
C654 source.n253 a_n1564_n3288# 0.01934f
C655 source.n254 a_n1564_n3288# 0.020478f
C656 source.n255 a_n1564_n3288# 0.045713f
C657 source.n256 a_n1564_n3288# 0.045713f
C658 source.n257 a_n1564_n3288# 0.020478f
C659 source.n258 a_n1564_n3288# 0.01934f
C660 source.n259 a_n1564_n3288# 0.035991f
C661 source.n260 a_n1564_n3288# 0.035991f
C662 source.n261 a_n1564_n3288# 0.01934f
C663 source.n262 a_n1564_n3288# 0.01934f
C664 source.n263 a_n1564_n3288# 0.020478f
C665 source.n264 a_n1564_n3288# 0.045713f
C666 source.n265 a_n1564_n3288# 0.045713f
C667 source.n266 a_n1564_n3288# 0.045713f
C668 source.n267 a_n1564_n3288# 0.019909f
C669 source.n268 a_n1564_n3288# 0.01934f
C670 source.n269 a_n1564_n3288# 0.035991f
C671 source.n270 a_n1564_n3288# 0.035991f
C672 source.n271 a_n1564_n3288# 0.01934f
C673 source.n272 a_n1564_n3288# 0.020478f
C674 source.n273 a_n1564_n3288# 0.045713f
C675 source.n274 a_n1564_n3288# 0.045713f
C676 source.n275 a_n1564_n3288# 0.020478f
C677 source.n276 a_n1564_n3288# 0.01934f
C678 source.n277 a_n1564_n3288# 0.035991f
C679 source.n278 a_n1564_n3288# 0.035991f
C680 source.n279 a_n1564_n3288# 0.01934f
C681 source.n280 a_n1564_n3288# 0.020478f
C682 source.n281 a_n1564_n3288# 0.045713f
C683 source.n282 a_n1564_n3288# 0.093807f
C684 source.n283 a_n1564_n3288# 0.020478f
C685 source.n284 a_n1564_n3288# 0.01934f
C686 source.n285 a_n1564_n3288# 0.077291f
C687 source.n286 a_n1564_n3288# 0.051771f
C688 source.n287 a_n1564_n3288# 0.330043f
C689 source.n288 a_n1564_n3288# 2.25229f
C690 minus.n0 a_n1564_n3288# 0.055147f
C691 minus.t1 a_n1564_n3288# 0.378678f
C692 minus.t7 a_n1564_n3288# 0.374008f
C693 minus.t12 a_n1564_n3288# 0.374008f
C694 minus.t13 a_n1564_n3288# 0.374008f
C695 minus.n1 a_n1564_n3288# 0.154033f
C696 minus.n2 a_n1564_n3288# 0.123135f
C697 minus.t0 a_n1564_n3288# 0.374008f
C698 minus.t8 a_n1564_n3288# 0.374008f
C699 minus.t11 a_n1564_n3288# 0.378678f
C700 minus.n3 a_n1564_n3288# 0.170117f
C701 minus.n4 a_n1564_n3288# 0.154033f
C702 minus.n5 a_n1564_n3288# 0.019314f
C703 minus.n6 a_n1564_n3288# 0.154033f
C704 minus.n7 a_n1564_n3288# 0.019314f
C705 minus.n8 a_n1564_n3288# 0.055147f
C706 minus.n9 a_n1564_n3288# 0.055147f
C707 minus.n10 a_n1564_n3288# 0.019314f
C708 minus.n11 a_n1564_n3288# 0.154033f
C709 minus.n12 a_n1564_n3288# 0.019314f
C710 minus.n13 a_n1564_n3288# 0.154033f
C711 minus.n14 a_n1564_n3288# 0.170037f
C712 minus.n15 a_n1564_n3288# 1.84748f
C713 minus.n16 a_n1564_n3288# 0.055147f
C714 minus.t6 a_n1564_n3288# 0.374008f
C715 minus.t10 a_n1564_n3288# 0.374008f
C716 minus.t4 a_n1564_n3288# 0.374008f
C717 minus.n17 a_n1564_n3288# 0.154033f
C718 minus.n18 a_n1564_n3288# 0.123135f
C719 minus.t2 a_n1564_n3288# 0.374008f
C720 minus.t5 a_n1564_n3288# 0.374008f
C721 minus.t3 a_n1564_n3288# 0.378678f
C722 minus.n19 a_n1564_n3288# 0.170117f
C723 minus.n20 a_n1564_n3288# 0.154033f
C724 minus.n21 a_n1564_n3288# 0.019314f
C725 minus.n22 a_n1564_n3288# 0.154033f
C726 minus.n23 a_n1564_n3288# 0.019314f
C727 minus.n24 a_n1564_n3288# 0.055147f
C728 minus.n25 a_n1564_n3288# 0.055147f
C729 minus.n26 a_n1564_n3288# 0.019314f
C730 minus.n27 a_n1564_n3288# 0.154033f
C731 minus.n28 a_n1564_n3288# 0.019314f
C732 minus.n29 a_n1564_n3288# 0.154033f
C733 minus.t9 a_n1564_n3288# 0.378678f
C734 minus.n30 a_n1564_n3288# 0.170037f
C735 minus.n31 a_n1564_n3288# 0.355427f
C736 minus.n32 a_n1564_n3288# 2.25378f
.ends

