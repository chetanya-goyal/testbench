* NGSPICE file created from diffpair229.ext - technology: sky130A

.subckt diffpair229 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t32 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 source.t41 minus.t1 drain_right.t22 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X3 drain_left.t23 plus.t0 source.t10 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X4 source.t16 plus.t1 drain_left.t22 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 source.t7 plus.t2 drain_left.t21 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X6 source.t47 minus.t2 drain_right.t21 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X7 drain_left.t20 plus.t3 source.t9 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X8 a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X9 source.t15 plus.t4 drain_left.t19 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X10 source.t1 plus.t5 drain_left.t18 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X11 source.t3 plus.t6 drain_left.t17 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X12 drain_right.t20 minus.t3 source.t42 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X13 drain_right.t19 minus.t4 source.t40 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X14 source.t39 minus.t5 drain_right.t18 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X15 drain_right.t17 minus.t6 source.t43 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 source.t45 minus.t7 drain_right.t16 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X17 drain_right.t15 minus.t8 source.t46 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X18 drain_left.t16 plus.t7 source.t11 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X19 source.t17 plus.t8 drain_left.t15 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X20 a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X21 drain_left.t14 plus.t9 source.t8 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X22 source.t5 plus.t10 drain_left.t13 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 drain_right.t14 minus.t9 source.t44 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X24 drain_right.t13 minus.t10 source.t33 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X25 drain_right.t12 minus.t11 source.t25 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X26 source.t34 minus.t12 drain_right.t11 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X27 drain_left.t12 plus.t11 source.t6 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X28 source.t37 minus.t13 drain_right.t10 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X29 drain_right.t9 minus.t14 source.t35 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X30 drain_left.t11 plus.t12 source.t2 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X31 drain_right.t8 minus.t15 source.t30 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X32 drain_left.t10 plus.t13 source.t4 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X33 source.t13 plus.t14 drain_left.t9 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X34 drain_left.t8 plus.t15 source.t21 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X35 drain_right.t7 minus.t16 source.t36 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X36 a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X37 drain_left.t7 plus.t16 source.t20 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X38 source.t38 minus.t17 drain_right.t6 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X39 source.t27 minus.t18 drain_right.t5 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X40 drain_left.t6 plus.t17 source.t12 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X41 source.t18 plus.t18 drain_left.t5 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X42 drain_right.t4 minus.t19 source.t24 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X43 drain_left.t4 plus.t19 source.t22 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X44 source.t26 minus.t20 drain_right.t3 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X45 source.t0 plus.t20 drain_left.t3 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X46 source.t29 minus.t21 drain_right.t2 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X47 drain_left.t2 plus.t21 source.t19 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X48 source.t28 minus.t22 drain_right.t1 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X49 source.t31 minus.t23 drain_right.t0 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X50 source.t14 plus.t22 drain_left.t1 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X51 source.t23 plus.t23 drain_left.t0 a_n3394_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n11 minus.t16 185.763
R1 minus.n53 minus.t1 185.763
R2 minus.n41 minus.n40 161.3
R3 minus.n39 minus.n0 161.3
R4 minus.n38 minus.n37 161.3
R5 minus.n36 minus.n1 161.3
R6 minus.n35 minus.n34 161.3
R7 minus.n33 minus.n2 161.3
R8 minus.n32 minus.n31 161.3
R9 minus.n30 minus.n3 161.3
R10 minus.n29 minus.n28 161.3
R11 minus.n27 minus.n4 161.3
R12 minus.n26 minus.n25 161.3
R13 minus.n24 minus.n5 161.3
R14 minus.n23 minus.n22 161.3
R15 minus.n21 minus.n6 161.3
R16 minus.n20 minus.n19 161.3
R17 minus.n18 minus.n7 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n8 161.3
R20 minus.n14 minus.n13 161.3
R21 minus.n12 minus.n9 161.3
R22 minus.n83 minus.n82 161.3
R23 minus.n81 minus.n42 161.3
R24 minus.n80 minus.n79 161.3
R25 minus.n78 minus.n43 161.3
R26 minus.n77 minus.n76 161.3
R27 minus.n75 minus.n44 161.3
R28 minus.n74 minus.n73 161.3
R29 minus.n72 minus.n45 161.3
R30 minus.n71 minus.n70 161.3
R31 minus.n69 minus.n46 161.3
R32 minus.n68 minus.n67 161.3
R33 minus.n66 minus.n47 161.3
R34 minus.n65 minus.n64 161.3
R35 minus.n63 minus.n48 161.3
R36 minus.n62 minus.n61 161.3
R37 minus.n60 minus.n49 161.3
R38 minus.n59 minus.n58 161.3
R39 minus.n57 minus.n50 161.3
R40 minus.n56 minus.n55 161.3
R41 minus.n54 minus.n51 161.3
R42 minus.n10 minus.t2 159.405
R43 minus.n14 minus.t15 159.405
R44 minus.n16 minus.t22 159.405
R45 minus.n20 minus.t10 159.405
R46 minus.n22 minus.t23 159.405
R47 minus.n26 minus.t9 159.405
R48 minus.n28 minus.t21 159.405
R49 minus.n32 minus.t8 159.405
R50 minus.n34 minus.t20 159.405
R51 minus.n38 minus.t3 159.405
R52 minus.n40 minus.t17 159.405
R53 minus.n52 minus.t0 159.405
R54 minus.n56 minus.t5 159.405
R55 minus.n58 minus.t4 159.405
R56 minus.n62 minus.t7 159.405
R57 minus.n64 minus.t14 159.405
R58 minus.n68 minus.t12 159.405
R59 minus.n70 minus.t19 159.405
R60 minus.n74 minus.t18 159.405
R61 minus.n76 minus.t6 159.405
R62 minus.n80 minus.t13 159.405
R63 minus.n82 minus.t11 159.405
R64 minus.n40 minus.n39 46.0096
R65 minus.n82 minus.n81 46.0096
R66 minus.n12 minus.n11 45.0871
R67 minus.n54 minus.n53 45.0871
R68 minus.n10 minus.n9 41.6278
R69 minus.n38 minus.n1 41.6278
R70 minus.n52 minus.n51 41.6278
R71 minus.n80 minus.n43 41.6278
R72 minus.n15 minus.n14 37.246
R73 minus.n34 minus.n33 37.246
R74 minus.n57 minus.n56 37.246
R75 minus.n76 minus.n75 37.246
R76 minus.n84 minus.n41 35.3376
R77 minus.n16 minus.n7 32.8641
R78 minus.n32 minus.n3 32.8641
R79 minus.n58 minus.n49 32.8641
R80 minus.n74 minus.n45 32.8641
R81 minus.n21 minus.n20 28.4823
R82 minus.n28 minus.n27 28.4823
R83 minus.n63 minus.n62 28.4823
R84 minus.n70 minus.n69 28.4823
R85 minus.n26 minus.n5 24.1005
R86 minus.n22 minus.n5 24.1005
R87 minus.n64 minus.n47 24.1005
R88 minus.n68 minus.n47 24.1005
R89 minus.n22 minus.n21 19.7187
R90 minus.n27 minus.n26 19.7187
R91 minus.n64 minus.n63 19.7187
R92 minus.n69 minus.n68 19.7187
R93 minus.n20 minus.n7 15.3369
R94 minus.n28 minus.n3 15.3369
R95 minus.n62 minus.n49 15.3369
R96 minus.n70 minus.n45 15.3369
R97 minus.n11 minus.n10 14.1472
R98 minus.n53 minus.n52 14.1472
R99 minus.n16 minus.n15 10.955
R100 minus.n33 minus.n32 10.955
R101 minus.n58 minus.n57 10.955
R102 minus.n75 minus.n74 10.955
R103 minus.n84 minus.n83 6.67853
R104 minus.n14 minus.n9 6.57323
R105 minus.n34 minus.n1 6.57323
R106 minus.n56 minus.n51 6.57323
R107 minus.n76 minus.n43 6.57323
R108 minus.n39 minus.n38 2.19141
R109 minus.n81 minus.n80 2.19141
R110 minus.n41 minus.n0 0.189894
R111 minus.n37 minus.n0 0.189894
R112 minus.n37 minus.n36 0.189894
R113 minus.n36 minus.n35 0.189894
R114 minus.n35 minus.n2 0.189894
R115 minus.n31 minus.n2 0.189894
R116 minus.n31 minus.n30 0.189894
R117 minus.n30 minus.n29 0.189894
R118 minus.n29 minus.n4 0.189894
R119 minus.n25 minus.n4 0.189894
R120 minus.n25 minus.n24 0.189894
R121 minus.n24 minus.n23 0.189894
R122 minus.n23 minus.n6 0.189894
R123 minus.n19 minus.n6 0.189894
R124 minus.n19 minus.n18 0.189894
R125 minus.n18 minus.n17 0.189894
R126 minus.n17 minus.n8 0.189894
R127 minus.n13 minus.n8 0.189894
R128 minus.n13 minus.n12 0.189894
R129 minus.n55 minus.n54 0.189894
R130 minus.n55 minus.n50 0.189894
R131 minus.n59 minus.n50 0.189894
R132 minus.n60 minus.n59 0.189894
R133 minus.n61 minus.n60 0.189894
R134 minus.n61 minus.n48 0.189894
R135 minus.n65 minus.n48 0.189894
R136 minus.n66 minus.n65 0.189894
R137 minus.n67 minus.n66 0.189894
R138 minus.n67 minus.n46 0.189894
R139 minus.n71 minus.n46 0.189894
R140 minus.n72 minus.n71 0.189894
R141 minus.n73 minus.n72 0.189894
R142 minus.n73 minus.n44 0.189894
R143 minus.n77 minus.n44 0.189894
R144 minus.n78 minus.n77 0.189894
R145 minus.n79 minus.n78 0.189894
R146 minus.n79 minus.n42 0.189894
R147 minus.n83 minus.n42 0.189894
R148 minus minus.n84 0.188
R149 source.n0 source.t10 69.6943
R150 source.n11 source.t3 69.6943
R151 source.n12 source.t36 69.6943
R152 source.n23 source.t38 69.6943
R153 source.n47 source.t25 69.6942
R154 source.n36 source.t41 69.6942
R155 source.n35 source.t11 69.6942
R156 source.n24 source.t18 69.6942
R157 source.n2 source.n1 63.0943
R158 source.n4 source.n3 63.0943
R159 source.n6 source.n5 63.0943
R160 source.n8 source.n7 63.0943
R161 source.n10 source.n9 63.0943
R162 source.n14 source.n13 63.0943
R163 source.n16 source.n15 63.0943
R164 source.n18 source.n17 63.0943
R165 source.n20 source.n19 63.0943
R166 source.n22 source.n21 63.0943
R167 source.n46 source.n45 63.0942
R168 source.n44 source.n43 63.0942
R169 source.n42 source.n41 63.0942
R170 source.n40 source.n39 63.0942
R171 source.n38 source.n37 63.0942
R172 source.n34 source.n33 63.0942
R173 source.n32 source.n31 63.0942
R174 source.n30 source.n29 63.0942
R175 source.n28 source.n27 63.0942
R176 source.n26 source.n25 63.0942
R177 source.n24 source.n23 15.3575
R178 source.n48 source.n0 9.65058
R179 source.n45 source.t43 6.6005
R180 source.n45 source.t37 6.6005
R181 source.n43 source.t24 6.6005
R182 source.n43 source.t27 6.6005
R183 source.n41 source.t35 6.6005
R184 source.n41 source.t34 6.6005
R185 source.n39 source.t40 6.6005
R186 source.n39 source.t45 6.6005
R187 source.n37 source.t32 6.6005
R188 source.n37 source.t39 6.6005
R189 source.n33 source.t2 6.6005
R190 source.n33 source.t17 6.6005
R191 source.n31 source.t22 6.6005
R192 source.n31 source.t0 6.6005
R193 source.n29 source.t19 6.6005
R194 source.n29 source.t14 6.6005
R195 source.n27 source.t8 6.6005
R196 source.n27 source.t15 6.6005
R197 source.n25 source.t12 6.6005
R198 source.n25 source.t5 6.6005
R199 source.n1 source.t9 6.6005
R200 source.n1 source.t13 6.6005
R201 source.n3 source.t6 6.6005
R202 source.n3 source.t23 6.6005
R203 source.n5 source.t21 6.6005
R204 source.n5 source.t16 6.6005
R205 source.n7 source.t4 6.6005
R206 source.n7 source.t1 6.6005
R207 source.n9 source.t20 6.6005
R208 source.n9 source.t7 6.6005
R209 source.n13 source.t30 6.6005
R210 source.n13 source.t47 6.6005
R211 source.n15 source.t33 6.6005
R212 source.n15 source.t28 6.6005
R213 source.n17 source.t44 6.6005
R214 source.n17 source.t31 6.6005
R215 source.n19 source.t46 6.6005
R216 source.n19 source.t29 6.6005
R217 source.n21 source.t42 6.6005
R218 source.n21 source.t26 6.6005
R219 source.n48 source.n47 5.7074
R220 source.n23 source.n22 0.888431
R221 source.n22 source.n20 0.888431
R222 source.n20 source.n18 0.888431
R223 source.n18 source.n16 0.888431
R224 source.n16 source.n14 0.888431
R225 source.n14 source.n12 0.888431
R226 source.n11 source.n10 0.888431
R227 source.n10 source.n8 0.888431
R228 source.n8 source.n6 0.888431
R229 source.n6 source.n4 0.888431
R230 source.n4 source.n2 0.888431
R231 source.n2 source.n0 0.888431
R232 source.n26 source.n24 0.888431
R233 source.n28 source.n26 0.888431
R234 source.n30 source.n28 0.888431
R235 source.n32 source.n30 0.888431
R236 source.n34 source.n32 0.888431
R237 source.n35 source.n34 0.888431
R238 source.n38 source.n36 0.888431
R239 source.n40 source.n38 0.888431
R240 source.n42 source.n40 0.888431
R241 source.n44 source.n42 0.888431
R242 source.n46 source.n44 0.888431
R243 source.n47 source.n46 0.888431
R244 source.n12 source.n11 0.470328
R245 source.n36 source.n35 0.470328
R246 source source.n48 0.188
R247 drain_right.n13 drain_right.n11 80.661
R248 drain_right.n7 drain_right.n5 80.6609
R249 drain_right.n2 drain_right.n0 80.6609
R250 drain_right.n13 drain_right.n12 79.7731
R251 drain_right.n15 drain_right.n14 79.7731
R252 drain_right.n17 drain_right.n16 79.7731
R253 drain_right.n19 drain_right.n18 79.7731
R254 drain_right.n21 drain_right.n20 79.7731
R255 drain_right.n7 drain_right.n6 79.773
R256 drain_right.n9 drain_right.n8 79.773
R257 drain_right.n4 drain_right.n3 79.773
R258 drain_right.n2 drain_right.n1 79.773
R259 drain_right drain_right.n10 28.431
R260 drain_right.n5 drain_right.t10 6.6005
R261 drain_right.n5 drain_right.t12 6.6005
R262 drain_right.n6 drain_right.t5 6.6005
R263 drain_right.n6 drain_right.t17 6.6005
R264 drain_right.n8 drain_right.t11 6.6005
R265 drain_right.n8 drain_right.t4 6.6005
R266 drain_right.n3 drain_right.t16 6.6005
R267 drain_right.n3 drain_right.t9 6.6005
R268 drain_right.n1 drain_right.t18 6.6005
R269 drain_right.n1 drain_right.t19 6.6005
R270 drain_right.n0 drain_right.t22 6.6005
R271 drain_right.n0 drain_right.t23 6.6005
R272 drain_right.n11 drain_right.t21 6.6005
R273 drain_right.n11 drain_right.t7 6.6005
R274 drain_right.n12 drain_right.t1 6.6005
R275 drain_right.n12 drain_right.t8 6.6005
R276 drain_right.n14 drain_right.t0 6.6005
R277 drain_right.n14 drain_right.t13 6.6005
R278 drain_right.n16 drain_right.t2 6.6005
R279 drain_right.n16 drain_right.t14 6.6005
R280 drain_right.n18 drain_right.t3 6.6005
R281 drain_right.n18 drain_right.t15 6.6005
R282 drain_right.n20 drain_right.t6 6.6005
R283 drain_right.n20 drain_right.t20 6.6005
R284 drain_right drain_right.n21 6.54115
R285 drain_right.n9 drain_right.n7 0.888431
R286 drain_right.n4 drain_right.n2 0.888431
R287 drain_right.n21 drain_right.n19 0.888431
R288 drain_right.n19 drain_right.n17 0.888431
R289 drain_right.n17 drain_right.n15 0.888431
R290 drain_right.n15 drain_right.n13 0.888431
R291 drain_right.n10 drain_right.n9 0.389119
R292 drain_right.n10 drain_right.n4 0.389119
R293 plus.n11 plus.t6 185.763
R294 plus.n53 plus.t7 185.763
R295 plus.n13 plus.n12 161.3
R296 plus.n14 plus.n9 161.3
R297 plus.n16 plus.n15 161.3
R298 plus.n17 plus.n8 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n7 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n23 plus.n6 161.3
R303 plus.n25 plus.n24 161.3
R304 plus.n26 plus.n5 161.3
R305 plus.n28 plus.n27 161.3
R306 plus.n29 plus.n4 161.3
R307 plus.n31 plus.n30 161.3
R308 plus.n32 plus.n3 161.3
R309 plus.n34 plus.n33 161.3
R310 plus.n35 plus.n2 161.3
R311 plus.n37 plus.n36 161.3
R312 plus.n38 plus.n1 161.3
R313 plus.n39 plus.n0 161.3
R314 plus.n41 plus.n40 161.3
R315 plus.n55 plus.n54 161.3
R316 plus.n56 plus.n51 161.3
R317 plus.n58 plus.n57 161.3
R318 plus.n59 plus.n50 161.3
R319 plus.n61 plus.n60 161.3
R320 plus.n62 plus.n49 161.3
R321 plus.n64 plus.n63 161.3
R322 plus.n65 plus.n48 161.3
R323 plus.n67 plus.n66 161.3
R324 plus.n68 plus.n47 161.3
R325 plus.n70 plus.n69 161.3
R326 plus.n71 plus.n46 161.3
R327 plus.n73 plus.n72 161.3
R328 plus.n74 plus.n45 161.3
R329 plus.n76 plus.n75 161.3
R330 plus.n77 plus.n44 161.3
R331 plus.n79 plus.n78 161.3
R332 plus.n80 plus.n43 161.3
R333 plus.n81 plus.n42 161.3
R334 plus.n83 plus.n82 161.3
R335 plus.n40 plus.t0 159.405
R336 plus.n38 plus.t14 159.405
R337 plus.n2 plus.t3 159.405
R338 plus.n32 plus.t23 159.405
R339 plus.n4 plus.t11 159.405
R340 plus.n26 plus.t1 159.405
R341 plus.n6 plus.t15 159.405
R342 plus.n20 plus.t5 159.405
R343 plus.n8 plus.t13 159.405
R344 plus.n14 plus.t2 159.405
R345 plus.n10 plus.t16 159.405
R346 plus.n82 plus.t18 159.405
R347 plus.n80 plus.t17 159.405
R348 plus.n44 plus.t10 159.405
R349 plus.n74 plus.t9 159.405
R350 plus.n46 plus.t4 159.405
R351 plus.n68 plus.t21 159.405
R352 plus.n48 plus.t22 159.405
R353 plus.n62 plus.t19 159.405
R354 plus.n50 plus.t20 159.405
R355 plus.n56 plus.t12 159.405
R356 plus.n52 plus.t8 159.405
R357 plus.n40 plus.n39 46.0096
R358 plus.n82 plus.n81 46.0096
R359 plus.n12 plus.n11 45.0871
R360 plus.n54 plus.n53 45.0871
R361 plus.n38 plus.n37 41.6278
R362 plus.n13 plus.n10 41.6278
R363 plus.n80 plus.n79 41.6278
R364 plus.n55 plus.n52 41.6278
R365 plus.n33 plus.n2 37.246
R366 plus.n15 plus.n14 37.246
R367 plus.n75 plus.n44 37.246
R368 plus.n57 plus.n56 37.246
R369 plus.n32 plus.n31 32.8641
R370 plus.n19 plus.n8 32.8641
R371 plus.n74 plus.n73 32.8641
R372 plus.n61 plus.n50 32.8641
R373 plus plus.n83 32.6278
R374 plus.n27 plus.n4 28.4823
R375 plus.n21 plus.n20 28.4823
R376 plus.n69 plus.n46 28.4823
R377 plus.n63 plus.n62 28.4823
R378 plus.n25 plus.n6 24.1005
R379 plus.n26 plus.n25 24.1005
R380 plus.n68 plus.n67 24.1005
R381 plus.n67 plus.n48 24.1005
R382 plus.n27 plus.n26 19.7187
R383 plus.n21 plus.n6 19.7187
R384 plus.n69 plus.n68 19.7187
R385 plus.n63 plus.n48 19.7187
R386 plus.n31 plus.n4 15.3369
R387 plus.n20 plus.n19 15.3369
R388 plus.n73 plus.n46 15.3369
R389 plus.n62 plus.n61 15.3369
R390 plus.n11 plus.n10 14.1472
R391 plus.n53 plus.n52 14.1472
R392 plus.n33 plus.n32 10.955
R393 plus.n15 plus.n8 10.955
R394 plus.n75 plus.n74 10.955
R395 plus.n57 plus.n50 10.955
R396 plus plus.n41 8.91338
R397 plus.n37 plus.n2 6.57323
R398 plus.n14 plus.n13 6.57323
R399 plus.n79 plus.n44 6.57323
R400 plus.n56 plus.n55 6.57323
R401 plus.n39 plus.n38 2.19141
R402 plus.n81 plus.n80 2.19141
R403 plus.n12 plus.n9 0.189894
R404 plus.n16 plus.n9 0.189894
R405 plus.n17 plus.n16 0.189894
R406 plus.n18 plus.n17 0.189894
R407 plus.n18 plus.n7 0.189894
R408 plus.n22 plus.n7 0.189894
R409 plus.n23 plus.n22 0.189894
R410 plus.n24 plus.n23 0.189894
R411 plus.n24 plus.n5 0.189894
R412 plus.n28 plus.n5 0.189894
R413 plus.n29 plus.n28 0.189894
R414 plus.n30 plus.n29 0.189894
R415 plus.n30 plus.n3 0.189894
R416 plus.n34 plus.n3 0.189894
R417 plus.n35 plus.n34 0.189894
R418 plus.n36 plus.n35 0.189894
R419 plus.n36 plus.n1 0.189894
R420 plus.n1 plus.n0 0.189894
R421 plus.n41 plus.n0 0.189894
R422 plus.n83 plus.n42 0.189894
R423 plus.n43 plus.n42 0.189894
R424 plus.n78 plus.n43 0.189894
R425 plus.n78 plus.n77 0.189894
R426 plus.n77 plus.n76 0.189894
R427 plus.n76 plus.n45 0.189894
R428 plus.n72 plus.n45 0.189894
R429 plus.n72 plus.n71 0.189894
R430 plus.n71 plus.n70 0.189894
R431 plus.n70 plus.n47 0.189894
R432 plus.n66 plus.n47 0.189894
R433 plus.n66 plus.n65 0.189894
R434 plus.n65 plus.n64 0.189894
R435 plus.n64 plus.n49 0.189894
R436 plus.n60 plus.n49 0.189894
R437 plus.n60 plus.n59 0.189894
R438 plus.n59 plus.n58 0.189894
R439 plus.n58 plus.n51 0.189894
R440 plus.n54 plus.n51 0.189894
R441 drain_left.n13 drain_left.n11 80.661
R442 drain_left.n7 drain_left.n5 80.6609
R443 drain_left.n2 drain_left.n0 80.6609
R444 drain_left.n21 drain_left.n20 79.7731
R445 drain_left.n19 drain_left.n18 79.7731
R446 drain_left.n17 drain_left.n16 79.7731
R447 drain_left.n15 drain_left.n14 79.7731
R448 drain_left.n13 drain_left.n12 79.7731
R449 drain_left.n7 drain_left.n6 79.773
R450 drain_left.n9 drain_left.n8 79.773
R451 drain_left.n4 drain_left.n3 79.773
R452 drain_left.n2 drain_left.n1 79.773
R453 drain_left drain_left.n10 28.9842
R454 drain_left.n5 drain_left.t15 6.6005
R455 drain_left.n5 drain_left.t16 6.6005
R456 drain_left.n6 drain_left.t3 6.6005
R457 drain_left.n6 drain_left.t11 6.6005
R458 drain_left.n8 drain_left.t1 6.6005
R459 drain_left.n8 drain_left.t4 6.6005
R460 drain_left.n3 drain_left.t19 6.6005
R461 drain_left.n3 drain_left.t2 6.6005
R462 drain_left.n1 drain_left.t13 6.6005
R463 drain_left.n1 drain_left.t14 6.6005
R464 drain_left.n0 drain_left.t5 6.6005
R465 drain_left.n0 drain_left.t6 6.6005
R466 drain_left.n20 drain_left.t9 6.6005
R467 drain_left.n20 drain_left.t23 6.6005
R468 drain_left.n18 drain_left.t0 6.6005
R469 drain_left.n18 drain_left.t20 6.6005
R470 drain_left.n16 drain_left.t22 6.6005
R471 drain_left.n16 drain_left.t12 6.6005
R472 drain_left.n14 drain_left.t18 6.6005
R473 drain_left.n14 drain_left.t8 6.6005
R474 drain_left.n12 drain_left.t21 6.6005
R475 drain_left.n12 drain_left.t10 6.6005
R476 drain_left.n11 drain_left.t17 6.6005
R477 drain_left.n11 drain_left.t7 6.6005
R478 drain_left drain_left.n21 6.54115
R479 drain_left.n9 drain_left.n7 0.888431
R480 drain_left.n4 drain_left.n2 0.888431
R481 drain_left.n15 drain_left.n13 0.888431
R482 drain_left.n17 drain_left.n15 0.888431
R483 drain_left.n19 drain_left.n17 0.888431
R484 drain_left.n21 drain_left.n19 0.888431
R485 drain_left.n10 drain_left.n9 0.389119
R486 drain_left.n10 drain_left.n4 0.389119
C0 drain_left plus 4.66759f
C1 source minus 5.14187f
C2 drain_left minus 0.179641f
C3 drain_right plus 0.50453f
C4 drain_right minus 4.32726f
C5 drain_left source 10.6568f
C6 drain_right source 10.659401f
C7 minus plus 5.72115f
C8 drain_right drain_left 1.87044f
C9 source plus 5.15586f
C10 drain_right a_n3394_n1488# 6.1775f
C11 drain_left a_n3394_n1488# 6.674731f
C12 source a_n3394_n1488# 4.245335f
C13 minus a_n3394_n1488# 12.961848f
C14 plus a_n3394_n1488# 14.45839f
C15 drain_left.t5 a_n3394_n1488# 0.06544f
C16 drain_left.t6 a_n3394_n1488# 0.06544f
C17 drain_left.n0 a_n3394_n1488# 0.476242f
C18 drain_left.t13 a_n3394_n1488# 0.06544f
C19 drain_left.t14 a_n3394_n1488# 0.06544f
C20 drain_left.n1 a_n3394_n1488# 0.471948f
C21 drain_left.n2 a_n3394_n1488# 0.764665f
C22 drain_left.t19 a_n3394_n1488# 0.06544f
C23 drain_left.t2 a_n3394_n1488# 0.06544f
C24 drain_left.n3 a_n3394_n1488# 0.471948f
C25 drain_left.n4 a_n3394_n1488# 0.336155f
C26 drain_left.t15 a_n3394_n1488# 0.06544f
C27 drain_left.t16 a_n3394_n1488# 0.06544f
C28 drain_left.n5 a_n3394_n1488# 0.476242f
C29 drain_left.t3 a_n3394_n1488# 0.06544f
C30 drain_left.t11 a_n3394_n1488# 0.06544f
C31 drain_left.n6 a_n3394_n1488# 0.471948f
C32 drain_left.n7 a_n3394_n1488# 0.764665f
C33 drain_left.t1 a_n3394_n1488# 0.06544f
C34 drain_left.t4 a_n3394_n1488# 0.06544f
C35 drain_left.n8 a_n3394_n1488# 0.471948f
C36 drain_left.n9 a_n3394_n1488# 0.336155f
C37 drain_left.n10 a_n3394_n1488# 1.28955f
C38 drain_left.t17 a_n3394_n1488# 0.06544f
C39 drain_left.t7 a_n3394_n1488# 0.06544f
C40 drain_left.n11 a_n3394_n1488# 0.476244f
C41 drain_left.t21 a_n3394_n1488# 0.06544f
C42 drain_left.t10 a_n3394_n1488# 0.06544f
C43 drain_left.n12 a_n3394_n1488# 0.47195f
C44 drain_left.n13 a_n3394_n1488# 0.76466f
C45 drain_left.t18 a_n3394_n1488# 0.06544f
C46 drain_left.t8 a_n3394_n1488# 0.06544f
C47 drain_left.n14 a_n3394_n1488# 0.47195f
C48 drain_left.n15 a_n3394_n1488# 0.378918f
C49 drain_left.t22 a_n3394_n1488# 0.06544f
C50 drain_left.t12 a_n3394_n1488# 0.06544f
C51 drain_left.n16 a_n3394_n1488# 0.47195f
C52 drain_left.n17 a_n3394_n1488# 0.378918f
C53 drain_left.t0 a_n3394_n1488# 0.06544f
C54 drain_left.t20 a_n3394_n1488# 0.06544f
C55 drain_left.n18 a_n3394_n1488# 0.47195f
C56 drain_left.n19 a_n3394_n1488# 0.378918f
C57 drain_left.t9 a_n3394_n1488# 0.06544f
C58 drain_left.t23 a_n3394_n1488# 0.06544f
C59 drain_left.n20 a_n3394_n1488# 0.47195f
C60 drain_left.n21 a_n3394_n1488# 0.623076f
C61 plus.n0 a_n3394_n1488# 0.042154f
C62 plus.t0 a_n3394_n1488# 0.265449f
C63 plus.t14 a_n3394_n1488# 0.265449f
C64 plus.n1 a_n3394_n1488# 0.042154f
C65 plus.t3 a_n3394_n1488# 0.265449f
C66 plus.n2 a_n3394_n1488# 0.154603f
C67 plus.n3 a_n3394_n1488# 0.042154f
C68 plus.t23 a_n3394_n1488# 0.265449f
C69 plus.t11 a_n3394_n1488# 0.265449f
C70 plus.n4 a_n3394_n1488# 0.154603f
C71 plus.n5 a_n3394_n1488# 0.042154f
C72 plus.t1 a_n3394_n1488# 0.265449f
C73 plus.t15 a_n3394_n1488# 0.265449f
C74 plus.n6 a_n3394_n1488# 0.154603f
C75 plus.n7 a_n3394_n1488# 0.042154f
C76 plus.t5 a_n3394_n1488# 0.265449f
C77 plus.t13 a_n3394_n1488# 0.265449f
C78 plus.n8 a_n3394_n1488# 0.154603f
C79 plus.n9 a_n3394_n1488# 0.042154f
C80 plus.t2 a_n3394_n1488# 0.265449f
C81 plus.t16 a_n3394_n1488# 0.265449f
C82 plus.n10 a_n3394_n1488# 0.16323f
C83 plus.t6 a_n3394_n1488# 0.287491f
C84 plus.n11 a_n3394_n1488# 0.134806f
C85 plus.n12 a_n3394_n1488# 0.181474f
C86 plus.n13 a_n3394_n1488# 0.009566f
C87 plus.n14 a_n3394_n1488# 0.154603f
C88 plus.n15 a_n3394_n1488# 0.009566f
C89 plus.n16 a_n3394_n1488# 0.042154f
C90 plus.n17 a_n3394_n1488# 0.042154f
C91 plus.n18 a_n3394_n1488# 0.042154f
C92 plus.n19 a_n3394_n1488# 0.009566f
C93 plus.n20 a_n3394_n1488# 0.154603f
C94 plus.n21 a_n3394_n1488# 0.009566f
C95 plus.n22 a_n3394_n1488# 0.042154f
C96 plus.n23 a_n3394_n1488# 0.042154f
C97 plus.n24 a_n3394_n1488# 0.042154f
C98 plus.n25 a_n3394_n1488# 0.009566f
C99 plus.n26 a_n3394_n1488# 0.154603f
C100 plus.n27 a_n3394_n1488# 0.009566f
C101 plus.n28 a_n3394_n1488# 0.042154f
C102 plus.n29 a_n3394_n1488# 0.042154f
C103 plus.n30 a_n3394_n1488# 0.042154f
C104 plus.n31 a_n3394_n1488# 0.009566f
C105 plus.n32 a_n3394_n1488# 0.154603f
C106 plus.n33 a_n3394_n1488# 0.009566f
C107 plus.n34 a_n3394_n1488# 0.042154f
C108 plus.n35 a_n3394_n1488# 0.042154f
C109 plus.n36 a_n3394_n1488# 0.042154f
C110 plus.n37 a_n3394_n1488# 0.009566f
C111 plus.n38 a_n3394_n1488# 0.154603f
C112 plus.n39 a_n3394_n1488# 0.009566f
C113 plus.n40 a_n3394_n1488# 0.154993f
C114 plus.n41 a_n3394_n1488# 0.333414f
C115 plus.n42 a_n3394_n1488# 0.042154f
C116 plus.t18 a_n3394_n1488# 0.265449f
C117 plus.n43 a_n3394_n1488# 0.042154f
C118 plus.t17 a_n3394_n1488# 0.265449f
C119 plus.t10 a_n3394_n1488# 0.265449f
C120 plus.n44 a_n3394_n1488# 0.154603f
C121 plus.n45 a_n3394_n1488# 0.042154f
C122 plus.t9 a_n3394_n1488# 0.265449f
C123 plus.t4 a_n3394_n1488# 0.265449f
C124 plus.n46 a_n3394_n1488# 0.154603f
C125 plus.n47 a_n3394_n1488# 0.042154f
C126 plus.t21 a_n3394_n1488# 0.265449f
C127 plus.t22 a_n3394_n1488# 0.265449f
C128 plus.n48 a_n3394_n1488# 0.154603f
C129 plus.n49 a_n3394_n1488# 0.042154f
C130 plus.t19 a_n3394_n1488# 0.265449f
C131 plus.t20 a_n3394_n1488# 0.265449f
C132 plus.n50 a_n3394_n1488# 0.154603f
C133 plus.n51 a_n3394_n1488# 0.042154f
C134 plus.t12 a_n3394_n1488# 0.265449f
C135 plus.t8 a_n3394_n1488# 0.265449f
C136 plus.n52 a_n3394_n1488# 0.16323f
C137 plus.t7 a_n3394_n1488# 0.287491f
C138 plus.n53 a_n3394_n1488# 0.134806f
C139 plus.n54 a_n3394_n1488# 0.181474f
C140 plus.n55 a_n3394_n1488# 0.009566f
C141 plus.n56 a_n3394_n1488# 0.154603f
C142 plus.n57 a_n3394_n1488# 0.009566f
C143 plus.n58 a_n3394_n1488# 0.042154f
C144 plus.n59 a_n3394_n1488# 0.042154f
C145 plus.n60 a_n3394_n1488# 0.042154f
C146 plus.n61 a_n3394_n1488# 0.009566f
C147 plus.n62 a_n3394_n1488# 0.154603f
C148 plus.n63 a_n3394_n1488# 0.009566f
C149 plus.n64 a_n3394_n1488# 0.042154f
C150 plus.n65 a_n3394_n1488# 0.042154f
C151 plus.n66 a_n3394_n1488# 0.042154f
C152 plus.n67 a_n3394_n1488# 0.009566f
C153 plus.n68 a_n3394_n1488# 0.154603f
C154 plus.n69 a_n3394_n1488# 0.009566f
C155 plus.n70 a_n3394_n1488# 0.042154f
C156 plus.n71 a_n3394_n1488# 0.042154f
C157 plus.n72 a_n3394_n1488# 0.042154f
C158 plus.n73 a_n3394_n1488# 0.009566f
C159 plus.n74 a_n3394_n1488# 0.154603f
C160 plus.n75 a_n3394_n1488# 0.009566f
C161 plus.n76 a_n3394_n1488# 0.042154f
C162 plus.n77 a_n3394_n1488# 0.042154f
C163 plus.n78 a_n3394_n1488# 0.042154f
C164 plus.n79 a_n3394_n1488# 0.009566f
C165 plus.n80 a_n3394_n1488# 0.154603f
C166 plus.n81 a_n3394_n1488# 0.009566f
C167 plus.n82 a_n3394_n1488# 0.154993f
C168 plus.n83 a_n3394_n1488# 1.35313f
C169 drain_right.t22 a_n3394_n1488# 0.064191f
C170 drain_right.t23 a_n3394_n1488# 0.064191f
C171 drain_right.n0 a_n3394_n1488# 0.467147f
C172 drain_right.t18 a_n3394_n1488# 0.064191f
C173 drain_right.t19 a_n3394_n1488# 0.064191f
C174 drain_right.n1 a_n3394_n1488# 0.462936f
C175 drain_right.n2 a_n3394_n1488# 0.750063f
C176 drain_right.t16 a_n3394_n1488# 0.064191f
C177 drain_right.t9 a_n3394_n1488# 0.064191f
C178 drain_right.n3 a_n3394_n1488# 0.462936f
C179 drain_right.n4 a_n3394_n1488# 0.329736f
C180 drain_right.t10 a_n3394_n1488# 0.064191f
C181 drain_right.t12 a_n3394_n1488# 0.064191f
C182 drain_right.n5 a_n3394_n1488# 0.467147f
C183 drain_right.t5 a_n3394_n1488# 0.064191f
C184 drain_right.t17 a_n3394_n1488# 0.064191f
C185 drain_right.n6 a_n3394_n1488# 0.462936f
C186 drain_right.n7 a_n3394_n1488# 0.750063f
C187 drain_right.t11 a_n3394_n1488# 0.064191f
C188 drain_right.t4 a_n3394_n1488# 0.064191f
C189 drain_right.n8 a_n3394_n1488# 0.462936f
C190 drain_right.n9 a_n3394_n1488# 0.329736f
C191 drain_right.n10 a_n3394_n1488# 1.21219f
C192 drain_right.t21 a_n3394_n1488# 0.064191f
C193 drain_right.t7 a_n3394_n1488# 0.064191f
C194 drain_right.n11 a_n3394_n1488# 0.46715f
C195 drain_right.t1 a_n3394_n1488# 0.064191f
C196 drain_right.t8 a_n3394_n1488# 0.064191f
C197 drain_right.n12 a_n3394_n1488# 0.462938f
C198 drain_right.n13 a_n3394_n1488# 0.750058f
C199 drain_right.t0 a_n3394_n1488# 0.064191f
C200 drain_right.t13 a_n3394_n1488# 0.064191f
C201 drain_right.n14 a_n3394_n1488# 0.462938f
C202 drain_right.n15 a_n3394_n1488# 0.371682f
C203 drain_right.t2 a_n3394_n1488# 0.064191f
C204 drain_right.t14 a_n3394_n1488# 0.064191f
C205 drain_right.n16 a_n3394_n1488# 0.462938f
C206 drain_right.n17 a_n3394_n1488# 0.371682f
C207 drain_right.t3 a_n3394_n1488# 0.064191f
C208 drain_right.t15 a_n3394_n1488# 0.064191f
C209 drain_right.n18 a_n3394_n1488# 0.462938f
C210 drain_right.n19 a_n3394_n1488# 0.371682f
C211 drain_right.t6 a_n3394_n1488# 0.064191f
C212 drain_right.t20 a_n3394_n1488# 0.064191f
C213 drain_right.n20 a_n3394_n1488# 0.462938f
C214 drain_right.n21 a_n3394_n1488# 0.611177f
C215 source.t10 a_n3394_n1488# 0.587821f
C216 source.n0 a_n3394_n1488# 0.860263f
C217 source.t9 a_n3394_n1488# 0.070789f
C218 source.t13 a_n3394_n1488# 0.070789f
C219 source.n1 a_n3394_n1488# 0.448844f
C220 source.n2 a_n3394_n1488# 0.430987f
C221 source.t6 a_n3394_n1488# 0.070789f
C222 source.t23 a_n3394_n1488# 0.070789f
C223 source.n3 a_n3394_n1488# 0.448844f
C224 source.n4 a_n3394_n1488# 0.430987f
C225 source.t21 a_n3394_n1488# 0.070789f
C226 source.t16 a_n3394_n1488# 0.070789f
C227 source.n5 a_n3394_n1488# 0.448844f
C228 source.n6 a_n3394_n1488# 0.430987f
C229 source.t4 a_n3394_n1488# 0.070789f
C230 source.t1 a_n3394_n1488# 0.070789f
C231 source.n7 a_n3394_n1488# 0.448844f
C232 source.n8 a_n3394_n1488# 0.430987f
C233 source.t20 a_n3394_n1488# 0.070789f
C234 source.t7 a_n3394_n1488# 0.070789f
C235 source.n9 a_n3394_n1488# 0.448844f
C236 source.n10 a_n3394_n1488# 0.430987f
C237 source.t3 a_n3394_n1488# 0.587821f
C238 source.n11 a_n3394_n1488# 0.444843f
C239 source.t36 a_n3394_n1488# 0.587821f
C240 source.n12 a_n3394_n1488# 0.444843f
C241 source.t30 a_n3394_n1488# 0.070789f
C242 source.t47 a_n3394_n1488# 0.070789f
C243 source.n13 a_n3394_n1488# 0.448844f
C244 source.n14 a_n3394_n1488# 0.430987f
C245 source.t33 a_n3394_n1488# 0.070789f
C246 source.t28 a_n3394_n1488# 0.070789f
C247 source.n15 a_n3394_n1488# 0.448844f
C248 source.n16 a_n3394_n1488# 0.430987f
C249 source.t44 a_n3394_n1488# 0.070789f
C250 source.t31 a_n3394_n1488# 0.070789f
C251 source.n17 a_n3394_n1488# 0.448844f
C252 source.n18 a_n3394_n1488# 0.430987f
C253 source.t46 a_n3394_n1488# 0.070789f
C254 source.t29 a_n3394_n1488# 0.070789f
C255 source.n19 a_n3394_n1488# 0.448844f
C256 source.n20 a_n3394_n1488# 0.430987f
C257 source.t42 a_n3394_n1488# 0.070789f
C258 source.t26 a_n3394_n1488# 0.070789f
C259 source.n21 a_n3394_n1488# 0.448844f
C260 source.n22 a_n3394_n1488# 0.430987f
C261 source.t38 a_n3394_n1488# 0.587821f
C262 source.n23 a_n3394_n1488# 1.17959f
C263 source.t18 a_n3394_n1488# 0.587818f
C264 source.n24 a_n3394_n1488# 1.1796f
C265 source.t12 a_n3394_n1488# 0.070789f
C266 source.t5 a_n3394_n1488# 0.070789f
C267 source.n25 a_n3394_n1488# 0.448841f
C268 source.n26 a_n3394_n1488# 0.43099f
C269 source.t8 a_n3394_n1488# 0.070789f
C270 source.t15 a_n3394_n1488# 0.070789f
C271 source.n27 a_n3394_n1488# 0.448841f
C272 source.n28 a_n3394_n1488# 0.43099f
C273 source.t19 a_n3394_n1488# 0.070789f
C274 source.t14 a_n3394_n1488# 0.070789f
C275 source.n29 a_n3394_n1488# 0.448841f
C276 source.n30 a_n3394_n1488# 0.43099f
C277 source.t22 a_n3394_n1488# 0.070789f
C278 source.t0 a_n3394_n1488# 0.070789f
C279 source.n31 a_n3394_n1488# 0.448841f
C280 source.n32 a_n3394_n1488# 0.43099f
C281 source.t2 a_n3394_n1488# 0.070789f
C282 source.t17 a_n3394_n1488# 0.070789f
C283 source.n33 a_n3394_n1488# 0.448841f
C284 source.n34 a_n3394_n1488# 0.43099f
C285 source.t11 a_n3394_n1488# 0.587818f
C286 source.n35 a_n3394_n1488# 0.444846f
C287 source.t41 a_n3394_n1488# 0.587818f
C288 source.n36 a_n3394_n1488# 0.444846f
C289 source.t32 a_n3394_n1488# 0.070789f
C290 source.t39 a_n3394_n1488# 0.070789f
C291 source.n37 a_n3394_n1488# 0.448841f
C292 source.n38 a_n3394_n1488# 0.43099f
C293 source.t40 a_n3394_n1488# 0.070789f
C294 source.t45 a_n3394_n1488# 0.070789f
C295 source.n39 a_n3394_n1488# 0.448841f
C296 source.n40 a_n3394_n1488# 0.43099f
C297 source.t35 a_n3394_n1488# 0.070789f
C298 source.t34 a_n3394_n1488# 0.070789f
C299 source.n41 a_n3394_n1488# 0.448841f
C300 source.n42 a_n3394_n1488# 0.43099f
C301 source.t24 a_n3394_n1488# 0.070789f
C302 source.t27 a_n3394_n1488# 0.070789f
C303 source.n43 a_n3394_n1488# 0.448841f
C304 source.n44 a_n3394_n1488# 0.43099f
C305 source.t43 a_n3394_n1488# 0.070789f
C306 source.t37 a_n3394_n1488# 0.070789f
C307 source.n45 a_n3394_n1488# 0.448841f
C308 source.n46 a_n3394_n1488# 0.43099f
C309 source.t25 a_n3394_n1488# 0.587818f
C310 source.n47 a_n3394_n1488# 0.639625f
C311 source.n48 a_n3394_n1488# 0.880538f
C312 minus.n0 a_n3394_n1488# 0.040581f
C313 minus.n1 a_n3394_n1488# 0.009209f
C314 minus.t3 a_n3394_n1488# 0.255544f
C315 minus.n2 a_n3394_n1488# 0.040581f
C316 minus.n3 a_n3394_n1488# 0.009209f
C317 minus.t8 a_n3394_n1488# 0.255544f
C318 minus.n4 a_n3394_n1488# 0.040581f
C319 minus.n5 a_n3394_n1488# 0.009209f
C320 minus.t9 a_n3394_n1488# 0.255544f
C321 minus.n6 a_n3394_n1488# 0.040581f
C322 minus.n7 a_n3394_n1488# 0.009209f
C323 minus.t10 a_n3394_n1488# 0.255544f
C324 minus.n8 a_n3394_n1488# 0.040581f
C325 minus.n9 a_n3394_n1488# 0.009209f
C326 minus.t15 a_n3394_n1488# 0.255544f
C327 minus.t16 a_n3394_n1488# 0.276764f
C328 minus.t2 a_n3394_n1488# 0.255544f
C329 minus.n10 a_n3394_n1488# 0.157139f
C330 minus.n11 a_n3394_n1488# 0.129776f
C331 minus.n12 a_n3394_n1488# 0.174703f
C332 minus.n13 a_n3394_n1488# 0.040581f
C333 minus.n14 a_n3394_n1488# 0.148835f
C334 minus.n15 a_n3394_n1488# 0.009209f
C335 minus.t22 a_n3394_n1488# 0.255544f
C336 minus.n16 a_n3394_n1488# 0.148835f
C337 minus.n17 a_n3394_n1488# 0.040581f
C338 minus.n18 a_n3394_n1488# 0.040581f
C339 minus.n19 a_n3394_n1488# 0.040581f
C340 minus.n20 a_n3394_n1488# 0.148835f
C341 minus.n21 a_n3394_n1488# 0.009209f
C342 minus.t23 a_n3394_n1488# 0.255544f
C343 minus.n22 a_n3394_n1488# 0.148835f
C344 minus.n23 a_n3394_n1488# 0.040581f
C345 minus.n24 a_n3394_n1488# 0.040581f
C346 minus.n25 a_n3394_n1488# 0.040581f
C347 minus.n26 a_n3394_n1488# 0.148835f
C348 minus.n27 a_n3394_n1488# 0.009209f
C349 minus.t21 a_n3394_n1488# 0.255544f
C350 minus.n28 a_n3394_n1488# 0.148835f
C351 minus.n29 a_n3394_n1488# 0.040581f
C352 minus.n30 a_n3394_n1488# 0.040581f
C353 minus.n31 a_n3394_n1488# 0.040581f
C354 minus.n32 a_n3394_n1488# 0.148835f
C355 minus.n33 a_n3394_n1488# 0.009209f
C356 minus.t20 a_n3394_n1488# 0.255544f
C357 minus.n34 a_n3394_n1488# 0.148835f
C358 minus.n35 a_n3394_n1488# 0.040581f
C359 minus.n36 a_n3394_n1488# 0.040581f
C360 minus.n37 a_n3394_n1488# 0.040581f
C361 minus.n38 a_n3394_n1488# 0.148835f
C362 minus.n39 a_n3394_n1488# 0.009209f
C363 minus.t17 a_n3394_n1488# 0.255544f
C364 minus.n40 a_n3394_n1488# 0.14921f
C365 minus.n41 a_n3394_n1488# 1.38694f
C366 minus.n42 a_n3394_n1488# 0.040581f
C367 minus.n43 a_n3394_n1488# 0.009209f
C368 minus.n44 a_n3394_n1488# 0.040581f
C369 minus.n45 a_n3394_n1488# 0.009209f
C370 minus.n46 a_n3394_n1488# 0.040581f
C371 minus.n47 a_n3394_n1488# 0.009209f
C372 minus.n48 a_n3394_n1488# 0.040581f
C373 minus.n49 a_n3394_n1488# 0.009209f
C374 minus.n50 a_n3394_n1488# 0.040581f
C375 minus.n51 a_n3394_n1488# 0.009209f
C376 minus.t1 a_n3394_n1488# 0.276764f
C377 minus.t0 a_n3394_n1488# 0.255544f
C378 minus.n52 a_n3394_n1488# 0.157139f
C379 minus.n53 a_n3394_n1488# 0.129776f
C380 minus.n54 a_n3394_n1488# 0.174703f
C381 minus.n55 a_n3394_n1488# 0.040581f
C382 minus.t5 a_n3394_n1488# 0.255544f
C383 minus.n56 a_n3394_n1488# 0.148835f
C384 minus.n57 a_n3394_n1488# 0.009209f
C385 minus.t4 a_n3394_n1488# 0.255544f
C386 minus.n58 a_n3394_n1488# 0.148835f
C387 minus.n59 a_n3394_n1488# 0.040581f
C388 minus.n60 a_n3394_n1488# 0.040581f
C389 minus.n61 a_n3394_n1488# 0.040581f
C390 minus.t7 a_n3394_n1488# 0.255544f
C391 minus.n62 a_n3394_n1488# 0.148835f
C392 minus.n63 a_n3394_n1488# 0.009209f
C393 minus.t14 a_n3394_n1488# 0.255544f
C394 minus.n64 a_n3394_n1488# 0.148835f
C395 minus.n65 a_n3394_n1488# 0.040581f
C396 minus.n66 a_n3394_n1488# 0.040581f
C397 minus.n67 a_n3394_n1488# 0.040581f
C398 minus.t12 a_n3394_n1488# 0.255544f
C399 minus.n68 a_n3394_n1488# 0.148835f
C400 minus.n69 a_n3394_n1488# 0.009209f
C401 minus.t19 a_n3394_n1488# 0.255544f
C402 minus.n70 a_n3394_n1488# 0.148835f
C403 minus.n71 a_n3394_n1488# 0.040581f
C404 minus.n72 a_n3394_n1488# 0.040581f
C405 minus.n73 a_n3394_n1488# 0.040581f
C406 minus.t18 a_n3394_n1488# 0.255544f
C407 minus.n74 a_n3394_n1488# 0.148835f
C408 minus.n75 a_n3394_n1488# 0.009209f
C409 minus.t6 a_n3394_n1488# 0.255544f
C410 minus.n76 a_n3394_n1488# 0.148835f
C411 minus.n77 a_n3394_n1488# 0.040581f
C412 minus.n78 a_n3394_n1488# 0.040581f
C413 minus.n79 a_n3394_n1488# 0.040581f
C414 minus.t13 a_n3394_n1488# 0.255544f
C415 minus.n80 a_n3394_n1488# 0.148835f
C416 minus.n81 a_n3394_n1488# 0.009209f
C417 minus.t11 a_n3394_n1488# 0.255544f
C418 minus.n82 a_n3394_n1488# 0.14921f
C419 minus.n83 a_n3394_n1488# 0.282235f
C420 minus.n84 a_n3394_n1488# 1.6829f
.ends

