* NGSPICE file created from diffpair418.ext - technology: sky130A

.subckt diffpair418 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t23 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X1 drain_right.t18 minus.t1 source.t18 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X2 source.t28 minus.t2 drain_right.t17 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X3 source.t26 minus.t3 drain_right.t16 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X4 source.t7 plus.t0 drain_left.t19 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X5 drain_left.t18 plus.t1 source.t10 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X6 drain_right.t15 minus.t4 source.t36 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X7 drain_right.t14 minus.t5 source.t33 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X8 drain_right.t13 minus.t6 source.t22 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X9 a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X10 drain_right.t12 minus.t7 source.t24 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X11 drain_right.t11 minus.t8 source.t20 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X12 source.t19 minus.t9 drain_right.t10 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X13 source.t29 minus.t10 drain_right.t9 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X14 drain_left.t17 plus.t2 source.t12 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X15 source.t27 minus.t11 drain_right.t8 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X16 source.t37 minus.t12 drain_right.t7 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X17 source.t25 minus.t13 drain_right.t6 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X18 source.t16 plus.t3 drain_left.t16 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X19 drain_left.t15 plus.t4 source.t9 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X20 source.t13 plus.t5 drain_left.t14 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X21 source.t32 minus.t14 drain_right.t5 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X22 drain_left.t13 plus.t6 source.t14 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X23 a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X24 drain_right.t4 minus.t15 source.t21 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X25 drain_right.t3 minus.t16 source.t30 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X26 drain_right.t2 minus.t17 source.t34 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X27 source.t17 plus.t7 drain_left.t12 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X28 source.t2 plus.t8 drain_left.t11 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X29 source.t5 plus.t9 drain_left.t10 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X30 source.t1 plus.t10 drain_left.t9 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X31 a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X32 source.t4 plus.t11 drain_left.t8 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X33 drain_left.t7 plus.t12 source.t11 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X34 drain_left.t6 plus.t13 source.t15 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X35 drain_left.t5 plus.t14 source.t8 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X36 drain_left.t4 plus.t15 source.t6 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X37 source.t35 minus.t18 drain_right.t1 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X38 source.t31 minus.t19 drain_right.t0 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X39 drain_left.t3 plus.t16 source.t38 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X40 drain_left.t2 plus.t17 source.t39 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X41 source.t3 plus.t18 drain_left.t1 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X42 a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X43 source.t0 plus.t19 drain_left.t0 a_n1882_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 minus.n23 minus.t12 1658.88
R1 minus.n5 minus.t16 1658.88
R2 minus.n48 minus.t4 1658.88
R3 minus.n30 minus.t3 1658.88
R4 minus.n22 minus.t15 1602.65
R5 minus.n20 minus.t19 1602.65
R6 minus.n1 minus.t1 1602.65
R7 minus.n15 minus.t9 1602.65
R8 minus.n13 minus.t17 1602.65
R9 minus.n3 minus.t18 1602.65
R10 minus.n8 minus.t0 1602.65
R11 minus.n6 minus.t10 1602.65
R12 minus.n47 minus.t11 1602.65
R13 minus.n45 minus.t7 1602.65
R14 minus.n26 minus.t13 1602.65
R15 minus.n40 minus.t8 1602.65
R16 minus.n38 minus.t14 1602.65
R17 minus.n28 minus.t5 1602.65
R18 minus.n33 minus.t2 1602.65
R19 minus.n31 minus.t6 1602.65
R20 minus.n5 minus.n4 161.489
R21 minus.n30 minus.n29 161.489
R22 minus.n24 minus.n23 161.3
R23 minus.n21 minus.n0 161.3
R24 minus.n19 minus.n18 161.3
R25 minus.n17 minus.n16 161.3
R26 minus.n14 minus.n2 161.3
R27 minus.n12 minus.n11 161.3
R28 minus.n10 minus.n9 161.3
R29 minus.n7 minus.n4 161.3
R30 minus.n49 minus.n48 161.3
R31 minus.n46 minus.n25 161.3
R32 minus.n44 minus.n43 161.3
R33 minus.n42 minus.n41 161.3
R34 minus.n39 minus.n27 161.3
R35 minus.n37 minus.n36 161.3
R36 minus.n35 minus.n34 161.3
R37 minus.n32 minus.n29 161.3
R38 minus.n22 minus.n21 51.852
R39 minus.n7 minus.n6 51.852
R40 minus.n32 minus.n31 51.852
R41 minus.n47 minus.n46 51.852
R42 minus.n20 minus.n19 47.4702
R43 minus.n9 minus.n8 47.4702
R44 minus.n34 minus.n33 47.4702
R45 minus.n45 minus.n44 47.4702
R46 minus.n16 minus.n1 43.0884
R47 minus.n12 minus.n3 43.0884
R48 minus.n37 minus.n28 43.0884
R49 minus.n41 minus.n26 43.0884
R50 minus.n15 minus.n14 38.7066
R51 minus.n14 minus.n13 38.7066
R52 minus.n39 minus.n38 38.7066
R53 minus.n40 minus.n39 38.7066
R54 minus.n50 minus.n24 36.2278
R55 minus.n16 minus.n15 34.3247
R56 minus.n13 minus.n12 34.3247
R57 minus.n38 minus.n37 34.3247
R58 minus.n41 minus.n40 34.3247
R59 minus.n19 minus.n1 29.9429
R60 minus.n9 minus.n3 29.9429
R61 minus.n34 minus.n28 29.9429
R62 minus.n44 minus.n26 29.9429
R63 minus.n21 minus.n20 25.5611
R64 minus.n8 minus.n7 25.5611
R65 minus.n33 minus.n32 25.5611
R66 minus.n46 minus.n45 25.5611
R67 minus.n23 minus.n22 21.1793
R68 minus.n6 minus.n5 21.1793
R69 minus.n31 minus.n30 21.1793
R70 minus.n48 minus.n47 21.1793
R71 minus.n50 minus.n49 6.47777
R72 minus.n24 minus.n0 0.189894
R73 minus.n18 minus.n0 0.189894
R74 minus.n18 minus.n17 0.189894
R75 minus.n17 minus.n2 0.189894
R76 minus.n11 minus.n2 0.189894
R77 minus.n11 minus.n10 0.189894
R78 minus.n10 minus.n4 0.189894
R79 minus.n35 minus.n29 0.189894
R80 minus.n36 minus.n35 0.189894
R81 minus.n36 minus.n27 0.189894
R82 minus.n42 minus.n27 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n25 0.189894
R85 minus.n49 minus.n25 0.189894
R86 minus minus.n50 0.188
R87 source.n554 source.n494 289.615
R88 source.n480 source.n420 289.615
R89 source.n414 source.n354 289.615
R90 source.n340 source.n280 289.615
R91 source.n60 source.n0 289.615
R92 source.n134 source.n74 289.615
R93 source.n200 source.n140 289.615
R94 source.n274 source.n214 289.615
R95 source.n514 source.n513 185
R96 source.n519 source.n518 185
R97 source.n521 source.n520 185
R98 source.n510 source.n509 185
R99 source.n527 source.n526 185
R100 source.n529 source.n528 185
R101 source.n506 source.n505 185
R102 source.n536 source.n535 185
R103 source.n537 source.n504 185
R104 source.n539 source.n538 185
R105 source.n502 source.n501 185
R106 source.n545 source.n544 185
R107 source.n547 source.n546 185
R108 source.n498 source.n497 185
R109 source.n553 source.n552 185
R110 source.n555 source.n554 185
R111 source.n440 source.n439 185
R112 source.n445 source.n444 185
R113 source.n447 source.n446 185
R114 source.n436 source.n435 185
R115 source.n453 source.n452 185
R116 source.n455 source.n454 185
R117 source.n432 source.n431 185
R118 source.n462 source.n461 185
R119 source.n463 source.n430 185
R120 source.n465 source.n464 185
R121 source.n428 source.n427 185
R122 source.n471 source.n470 185
R123 source.n473 source.n472 185
R124 source.n424 source.n423 185
R125 source.n479 source.n478 185
R126 source.n481 source.n480 185
R127 source.n374 source.n373 185
R128 source.n379 source.n378 185
R129 source.n381 source.n380 185
R130 source.n370 source.n369 185
R131 source.n387 source.n386 185
R132 source.n389 source.n388 185
R133 source.n366 source.n365 185
R134 source.n396 source.n395 185
R135 source.n397 source.n364 185
R136 source.n399 source.n398 185
R137 source.n362 source.n361 185
R138 source.n405 source.n404 185
R139 source.n407 source.n406 185
R140 source.n358 source.n357 185
R141 source.n413 source.n412 185
R142 source.n415 source.n414 185
R143 source.n300 source.n299 185
R144 source.n305 source.n304 185
R145 source.n307 source.n306 185
R146 source.n296 source.n295 185
R147 source.n313 source.n312 185
R148 source.n315 source.n314 185
R149 source.n292 source.n291 185
R150 source.n322 source.n321 185
R151 source.n323 source.n290 185
R152 source.n325 source.n324 185
R153 source.n288 source.n287 185
R154 source.n331 source.n330 185
R155 source.n333 source.n332 185
R156 source.n284 source.n283 185
R157 source.n339 source.n338 185
R158 source.n341 source.n340 185
R159 source.n61 source.n60 185
R160 source.n59 source.n58 185
R161 source.n4 source.n3 185
R162 source.n53 source.n52 185
R163 source.n51 source.n50 185
R164 source.n8 source.n7 185
R165 source.n45 source.n44 185
R166 source.n43 source.n10 185
R167 source.n42 source.n41 185
R168 source.n13 source.n11 185
R169 source.n36 source.n35 185
R170 source.n34 source.n33 185
R171 source.n17 source.n16 185
R172 source.n28 source.n27 185
R173 source.n26 source.n25 185
R174 source.n21 source.n20 185
R175 source.n135 source.n134 185
R176 source.n133 source.n132 185
R177 source.n78 source.n77 185
R178 source.n127 source.n126 185
R179 source.n125 source.n124 185
R180 source.n82 source.n81 185
R181 source.n119 source.n118 185
R182 source.n117 source.n84 185
R183 source.n116 source.n115 185
R184 source.n87 source.n85 185
R185 source.n110 source.n109 185
R186 source.n108 source.n107 185
R187 source.n91 source.n90 185
R188 source.n102 source.n101 185
R189 source.n100 source.n99 185
R190 source.n95 source.n94 185
R191 source.n201 source.n200 185
R192 source.n199 source.n198 185
R193 source.n144 source.n143 185
R194 source.n193 source.n192 185
R195 source.n191 source.n190 185
R196 source.n148 source.n147 185
R197 source.n185 source.n184 185
R198 source.n183 source.n150 185
R199 source.n182 source.n181 185
R200 source.n153 source.n151 185
R201 source.n176 source.n175 185
R202 source.n174 source.n173 185
R203 source.n157 source.n156 185
R204 source.n168 source.n167 185
R205 source.n166 source.n165 185
R206 source.n161 source.n160 185
R207 source.n275 source.n274 185
R208 source.n273 source.n272 185
R209 source.n218 source.n217 185
R210 source.n267 source.n266 185
R211 source.n265 source.n264 185
R212 source.n222 source.n221 185
R213 source.n259 source.n258 185
R214 source.n257 source.n224 185
R215 source.n256 source.n255 185
R216 source.n227 source.n225 185
R217 source.n250 source.n249 185
R218 source.n248 source.n247 185
R219 source.n231 source.n230 185
R220 source.n242 source.n241 185
R221 source.n240 source.n239 185
R222 source.n235 source.n234 185
R223 source.n515 source.t36 149.524
R224 source.n441 source.t26 149.524
R225 source.n375 source.t38 149.524
R226 source.n301 source.t16 149.524
R227 source.n22 source.t12 149.524
R228 source.n96 source.t13 149.524
R229 source.n162 source.t30 149.524
R230 source.n236 source.t37 149.524
R231 source.n519 source.n513 104.615
R232 source.n520 source.n519 104.615
R233 source.n520 source.n509 104.615
R234 source.n527 source.n509 104.615
R235 source.n528 source.n527 104.615
R236 source.n528 source.n505 104.615
R237 source.n536 source.n505 104.615
R238 source.n537 source.n536 104.615
R239 source.n538 source.n537 104.615
R240 source.n538 source.n501 104.615
R241 source.n545 source.n501 104.615
R242 source.n546 source.n545 104.615
R243 source.n546 source.n497 104.615
R244 source.n553 source.n497 104.615
R245 source.n554 source.n553 104.615
R246 source.n445 source.n439 104.615
R247 source.n446 source.n445 104.615
R248 source.n446 source.n435 104.615
R249 source.n453 source.n435 104.615
R250 source.n454 source.n453 104.615
R251 source.n454 source.n431 104.615
R252 source.n462 source.n431 104.615
R253 source.n463 source.n462 104.615
R254 source.n464 source.n463 104.615
R255 source.n464 source.n427 104.615
R256 source.n471 source.n427 104.615
R257 source.n472 source.n471 104.615
R258 source.n472 source.n423 104.615
R259 source.n479 source.n423 104.615
R260 source.n480 source.n479 104.615
R261 source.n379 source.n373 104.615
R262 source.n380 source.n379 104.615
R263 source.n380 source.n369 104.615
R264 source.n387 source.n369 104.615
R265 source.n388 source.n387 104.615
R266 source.n388 source.n365 104.615
R267 source.n396 source.n365 104.615
R268 source.n397 source.n396 104.615
R269 source.n398 source.n397 104.615
R270 source.n398 source.n361 104.615
R271 source.n405 source.n361 104.615
R272 source.n406 source.n405 104.615
R273 source.n406 source.n357 104.615
R274 source.n413 source.n357 104.615
R275 source.n414 source.n413 104.615
R276 source.n305 source.n299 104.615
R277 source.n306 source.n305 104.615
R278 source.n306 source.n295 104.615
R279 source.n313 source.n295 104.615
R280 source.n314 source.n313 104.615
R281 source.n314 source.n291 104.615
R282 source.n322 source.n291 104.615
R283 source.n323 source.n322 104.615
R284 source.n324 source.n323 104.615
R285 source.n324 source.n287 104.615
R286 source.n331 source.n287 104.615
R287 source.n332 source.n331 104.615
R288 source.n332 source.n283 104.615
R289 source.n339 source.n283 104.615
R290 source.n340 source.n339 104.615
R291 source.n60 source.n59 104.615
R292 source.n59 source.n3 104.615
R293 source.n52 source.n3 104.615
R294 source.n52 source.n51 104.615
R295 source.n51 source.n7 104.615
R296 source.n44 source.n7 104.615
R297 source.n44 source.n43 104.615
R298 source.n43 source.n42 104.615
R299 source.n42 source.n11 104.615
R300 source.n35 source.n11 104.615
R301 source.n35 source.n34 104.615
R302 source.n34 source.n16 104.615
R303 source.n27 source.n16 104.615
R304 source.n27 source.n26 104.615
R305 source.n26 source.n20 104.615
R306 source.n134 source.n133 104.615
R307 source.n133 source.n77 104.615
R308 source.n126 source.n77 104.615
R309 source.n126 source.n125 104.615
R310 source.n125 source.n81 104.615
R311 source.n118 source.n81 104.615
R312 source.n118 source.n117 104.615
R313 source.n117 source.n116 104.615
R314 source.n116 source.n85 104.615
R315 source.n109 source.n85 104.615
R316 source.n109 source.n108 104.615
R317 source.n108 source.n90 104.615
R318 source.n101 source.n90 104.615
R319 source.n101 source.n100 104.615
R320 source.n100 source.n94 104.615
R321 source.n200 source.n199 104.615
R322 source.n199 source.n143 104.615
R323 source.n192 source.n143 104.615
R324 source.n192 source.n191 104.615
R325 source.n191 source.n147 104.615
R326 source.n184 source.n147 104.615
R327 source.n184 source.n183 104.615
R328 source.n183 source.n182 104.615
R329 source.n182 source.n151 104.615
R330 source.n175 source.n151 104.615
R331 source.n175 source.n174 104.615
R332 source.n174 source.n156 104.615
R333 source.n167 source.n156 104.615
R334 source.n167 source.n166 104.615
R335 source.n166 source.n160 104.615
R336 source.n274 source.n273 104.615
R337 source.n273 source.n217 104.615
R338 source.n266 source.n217 104.615
R339 source.n266 source.n265 104.615
R340 source.n265 source.n221 104.615
R341 source.n258 source.n221 104.615
R342 source.n258 source.n257 104.615
R343 source.n257 source.n256 104.615
R344 source.n256 source.n225 104.615
R345 source.n249 source.n225 104.615
R346 source.n249 source.n248 104.615
R347 source.n248 source.n230 104.615
R348 source.n241 source.n230 104.615
R349 source.n241 source.n240 104.615
R350 source.n240 source.n234 104.615
R351 source.t36 source.n513 52.3082
R352 source.t26 source.n439 52.3082
R353 source.t38 source.n373 52.3082
R354 source.t16 source.n299 52.3082
R355 source.t12 source.n20 52.3082
R356 source.t13 source.n94 52.3082
R357 source.t30 source.n160 52.3082
R358 source.t37 source.n234 52.3082
R359 source.n67 source.n66 42.8739
R360 source.n69 source.n68 42.8739
R361 source.n71 source.n70 42.8739
R362 source.n73 source.n72 42.8739
R363 source.n207 source.n206 42.8739
R364 source.n209 source.n208 42.8739
R365 source.n211 source.n210 42.8739
R366 source.n213 source.n212 42.8739
R367 source.n493 source.n492 42.8737
R368 source.n491 source.n490 42.8737
R369 source.n489 source.n488 42.8737
R370 source.n487 source.n486 42.8737
R371 source.n353 source.n352 42.8737
R372 source.n351 source.n350 42.8737
R373 source.n349 source.n348 42.8737
R374 source.n347 source.n346 42.8737
R375 source.n559 source.n558 29.8581
R376 source.n485 source.n484 29.8581
R377 source.n419 source.n418 29.8581
R378 source.n345 source.n344 29.8581
R379 source.n65 source.n64 29.8581
R380 source.n139 source.n138 29.8581
R381 source.n205 source.n204 29.8581
R382 source.n279 source.n278 29.8581
R383 source.n345 source.n279 21.7446
R384 source.n560 source.n65 16.2532
R385 source.n539 source.n504 13.1884
R386 source.n465 source.n430 13.1884
R387 source.n399 source.n364 13.1884
R388 source.n325 source.n290 13.1884
R389 source.n45 source.n10 13.1884
R390 source.n119 source.n84 13.1884
R391 source.n185 source.n150 13.1884
R392 source.n259 source.n224 13.1884
R393 source.n535 source.n534 12.8005
R394 source.n540 source.n502 12.8005
R395 source.n461 source.n460 12.8005
R396 source.n466 source.n428 12.8005
R397 source.n395 source.n394 12.8005
R398 source.n400 source.n362 12.8005
R399 source.n321 source.n320 12.8005
R400 source.n326 source.n288 12.8005
R401 source.n46 source.n8 12.8005
R402 source.n41 source.n12 12.8005
R403 source.n120 source.n82 12.8005
R404 source.n115 source.n86 12.8005
R405 source.n186 source.n148 12.8005
R406 source.n181 source.n152 12.8005
R407 source.n260 source.n222 12.8005
R408 source.n255 source.n226 12.8005
R409 source.n533 source.n506 12.0247
R410 source.n544 source.n543 12.0247
R411 source.n459 source.n432 12.0247
R412 source.n470 source.n469 12.0247
R413 source.n393 source.n366 12.0247
R414 source.n404 source.n403 12.0247
R415 source.n319 source.n292 12.0247
R416 source.n330 source.n329 12.0247
R417 source.n50 source.n49 12.0247
R418 source.n40 source.n13 12.0247
R419 source.n124 source.n123 12.0247
R420 source.n114 source.n87 12.0247
R421 source.n190 source.n189 12.0247
R422 source.n180 source.n153 12.0247
R423 source.n264 source.n263 12.0247
R424 source.n254 source.n227 12.0247
R425 source.n530 source.n529 11.249
R426 source.n547 source.n500 11.249
R427 source.n456 source.n455 11.249
R428 source.n473 source.n426 11.249
R429 source.n390 source.n389 11.249
R430 source.n407 source.n360 11.249
R431 source.n316 source.n315 11.249
R432 source.n333 source.n286 11.249
R433 source.n53 source.n6 11.249
R434 source.n37 source.n36 11.249
R435 source.n127 source.n80 11.249
R436 source.n111 source.n110 11.249
R437 source.n193 source.n146 11.249
R438 source.n177 source.n176 11.249
R439 source.n267 source.n220 11.249
R440 source.n251 source.n250 11.249
R441 source.n526 source.n508 10.4732
R442 source.n548 source.n498 10.4732
R443 source.n452 source.n434 10.4732
R444 source.n474 source.n424 10.4732
R445 source.n386 source.n368 10.4732
R446 source.n408 source.n358 10.4732
R447 source.n312 source.n294 10.4732
R448 source.n334 source.n284 10.4732
R449 source.n54 source.n4 10.4732
R450 source.n33 source.n15 10.4732
R451 source.n128 source.n78 10.4732
R452 source.n107 source.n89 10.4732
R453 source.n194 source.n144 10.4732
R454 source.n173 source.n155 10.4732
R455 source.n268 source.n218 10.4732
R456 source.n247 source.n229 10.4732
R457 source.n515 source.n514 10.2747
R458 source.n441 source.n440 10.2747
R459 source.n375 source.n374 10.2747
R460 source.n301 source.n300 10.2747
R461 source.n22 source.n21 10.2747
R462 source.n96 source.n95 10.2747
R463 source.n162 source.n161 10.2747
R464 source.n236 source.n235 10.2747
R465 source.n525 source.n510 9.69747
R466 source.n552 source.n551 9.69747
R467 source.n451 source.n436 9.69747
R468 source.n478 source.n477 9.69747
R469 source.n385 source.n370 9.69747
R470 source.n412 source.n411 9.69747
R471 source.n311 source.n296 9.69747
R472 source.n338 source.n337 9.69747
R473 source.n58 source.n57 9.69747
R474 source.n32 source.n17 9.69747
R475 source.n132 source.n131 9.69747
R476 source.n106 source.n91 9.69747
R477 source.n198 source.n197 9.69747
R478 source.n172 source.n157 9.69747
R479 source.n272 source.n271 9.69747
R480 source.n246 source.n231 9.69747
R481 source.n558 source.n557 9.45567
R482 source.n484 source.n483 9.45567
R483 source.n418 source.n417 9.45567
R484 source.n344 source.n343 9.45567
R485 source.n64 source.n63 9.45567
R486 source.n138 source.n137 9.45567
R487 source.n204 source.n203 9.45567
R488 source.n278 source.n277 9.45567
R489 source.n557 source.n556 9.3005
R490 source.n496 source.n495 9.3005
R491 source.n551 source.n550 9.3005
R492 source.n549 source.n548 9.3005
R493 source.n500 source.n499 9.3005
R494 source.n543 source.n542 9.3005
R495 source.n541 source.n540 9.3005
R496 source.n517 source.n516 9.3005
R497 source.n512 source.n511 9.3005
R498 source.n523 source.n522 9.3005
R499 source.n525 source.n524 9.3005
R500 source.n508 source.n507 9.3005
R501 source.n531 source.n530 9.3005
R502 source.n533 source.n532 9.3005
R503 source.n534 source.n503 9.3005
R504 source.n483 source.n482 9.3005
R505 source.n422 source.n421 9.3005
R506 source.n477 source.n476 9.3005
R507 source.n475 source.n474 9.3005
R508 source.n426 source.n425 9.3005
R509 source.n469 source.n468 9.3005
R510 source.n467 source.n466 9.3005
R511 source.n443 source.n442 9.3005
R512 source.n438 source.n437 9.3005
R513 source.n449 source.n448 9.3005
R514 source.n451 source.n450 9.3005
R515 source.n434 source.n433 9.3005
R516 source.n457 source.n456 9.3005
R517 source.n459 source.n458 9.3005
R518 source.n460 source.n429 9.3005
R519 source.n417 source.n416 9.3005
R520 source.n356 source.n355 9.3005
R521 source.n411 source.n410 9.3005
R522 source.n409 source.n408 9.3005
R523 source.n360 source.n359 9.3005
R524 source.n403 source.n402 9.3005
R525 source.n401 source.n400 9.3005
R526 source.n377 source.n376 9.3005
R527 source.n372 source.n371 9.3005
R528 source.n383 source.n382 9.3005
R529 source.n385 source.n384 9.3005
R530 source.n368 source.n367 9.3005
R531 source.n391 source.n390 9.3005
R532 source.n393 source.n392 9.3005
R533 source.n394 source.n363 9.3005
R534 source.n343 source.n342 9.3005
R535 source.n282 source.n281 9.3005
R536 source.n337 source.n336 9.3005
R537 source.n335 source.n334 9.3005
R538 source.n286 source.n285 9.3005
R539 source.n329 source.n328 9.3005
R540 source.n327 source.n326 9.3005
R541 source.n303 source.n302 9.3005
R542 source.n298 source.n297 9.3005
R543 source.n309 source.n308 9.3005
R544 source.n311 source.n310 9.3005
R545 source.n294 source.n293 9.3005
R546 source.n317 source.n316 9.3005
R547 source.n319 source.n318 9.3005
R548 source.n320 source.n289 9.3005
R549 source.n24 source.n23 9.3005
R550 source.n19 source.n18 9.3005
R551 source.n30 source.n29 9.3005
R552 source.n32 source.n31 9.3005
R553 source.n15 source.n14 9.3005
R554 source.n38 source.n37 9.3005
R555 source.n40 source.n39 9.3005
R556 source.n12 source.n9 9.3005
R557 source.n63 source.n62 9.3005
R558 source.n2 source.n1 9.3005
R559 source.n57 source.n56 9.3005
R560 source.n55 source.n54 9.3005
R561 source.n6 source.n5 9.3005
R562 source.n49 source.n48 9.3005
R563 source.n47 source.n46 9.3005
R564 source.n98 source.n97 9.3005
R565 source.n93 source.n92 9.3005
R566 source.n104 source.n103 9.3005
R567 source.n106 source.n105 9.3005
R568 source.n89 source.n88 9.3005
R569 source.n112 source.n111 9.3005
R570 source.n114 source.n113 9.3005
R571 source.n86 source.n83 9.3005
R572 source.n137 source.n136 9.3005
R573 source.n76 source.n75 9.3005
R574 source.n131 source.n130 9.3005
R575 source.n129 source.n128 9.3005
R576 source.n80 source.n79 9.3005
R577 source.n123 source.n122 9.3005
R578 source.n121 source.n120 9.3005
R579 source.n164 source.n163 9.3005
R580 source.n159 source.n158 9.3005
R581 source.n170 source.n169 9.3005
R582 source.n172 source.n171 9.3005
R583 source.n155 source.n154 9.3005
R584 source.n178 source.n177 9.3005
R585 source.n180 source.n179 9.3005
R586 source.n152 source.n149 9.3005
R587 source.n203 source.n202 9.3005
R588 source.n142 source.n141 9.3005
R589 source.n197 source.n196 9.3005
R590 source.n195 source.n194 9.3005
R591 source.n146 source.n145 9.3005
R592 source.n189 source.n188 9.3005
R593 source.n187 source.n186 9.3005
R594 source.n238 source.n237 9.3005
R595 source.n233 source.n232 9.3005
R596 source.n244 source.n243 9.3005
R597 source.n246 source.n245 9.3005
R598 source.n229 source.n228 9.3005
R599 source.n252 source.n251 9.3005
R600 source.n254 source.n253 9.3005
R601 source.n226 source.n223 9.3005
R602 source.n277 source.n276 9.3005
R603 source.n216 source.n215 9.3005
R604 source.n271 source.n270 9.3005
R605 source.n269 source.n268 9.3005
R606 source.n220 source.n219 9.3005
R607 source.n263 source.n262 9.3005
R608 source.n261 source.n260 9.3005
R609 source.n522 source.n521 8.92171
R610 source.n555 source.n496 8.92171
R611 source.n448 source.n447 8.92171
R612 source.n481 source.n422 8.92171
R613 source.n382 source.n381 8.92171
R614 source.n415 source.n356 8.92171
R615 source.n308 source.n307 8.92171
R616 source.n341 source.n282 8.92171
R617 source.n61 source.n2 8.92171
R618 source.n29 source.n28 8.92171
R619 source.n135 source.n76 8.92171
R620 source.n103 source.n102 8.92171
R621 source.n201 source.n142 8.92171
R622 source.n169 source.n168 8.92171
R623 source.n275 source.n216 8.92171
R624 source.n243 source.n242 8.92171
R625 source.n518 source.n512 8.14595
R626 source.n556 source.n494 8.14595
R627 source.n444 source.n438 8.14595
R628 source.n482 source.n420 8.14595
R629 source.n378 source.n372 8.14595
R630 source.n416 source.n354 8.14595
R631 source.n304 source.n298 8.14595
R632 source.n342 source.n280 8.14595
R633 source.n62 source.n0 8.14595
R634 source.n25 source.n19 8.14595
R635 source.n136 source.n74 8.14595
R636 source.n99 source.n93 8.14595
R637 source.n202 source.n140 8.14595
R638 source.n165 source.n159 8.14595
R639 source.n276 source.n214 8.14595
R640 source.n239 source.n233 8.14595
R641 source.n517 source.n514 7.3702
R642 source.n443 source.n440 7.3702
R643 source.n377 source.n374 7.3702
R644 source.n303 source.n300 7.3702
R645 source.n24 source.n21 7.3702
R646 source.n98 source.n95 7.3702
R647 source.n164 source.n161 7.3702
R648 source.n238 source.n235 7.3702
R649 source.n518 source.n517 5.81868
R650 source.n558 source.n494 5.81868
R651 source.n444 source.n443 5.81868
R652 source.n484 source.n420 5.81868
R653 source.n378 source.n377 5.81868
R654 source.n418 source.n354 5.81868
R655 source.n304 source.n303 5.81868
R656 source.n344 source.n280 5.81868
R657 source.n64 source.n0 5.81868
R658 source.n25 source.n24 5.81868
R659 source.n138 source.n74 5.81868
R660 source.n99 source.n98 5.81868
R661 source.n204 source.n140 5.81868
R662 source.n165 source.n164 5.81868
R663 source.n278 source.n214 5.81868
R664 source.n239 source.n238 5.81868
R665 source.n560 source.n559 5.49188
R666 source.n521 source.n512 5.04292
R667 source.n556 source.n555 5.04292
R668 source.n447 source.n438 5.04292
R669 source.n482 source.n481 5.04292
R670 source.n381 source.n372 5.04292
R671 source.n416 source.n415 5.04292
R672 source.n307 source.n298 5.04292
R673 source.n342 source.n341 5.04292
R674 source.n62 source.n61 5.04292
R675 source.n28 source.n19 5.04292
R676 source.n136 source.n135 5.04292
R677 source.n102 source.n93 5.04292
R678 source.n202 source.n201 5.04292
R679 source.n168 source.n159 5.04292
R680 source.n276 source.n275 5.04292
R681 source.n242 source.n233 5.04292
R682 source.n522 source.n510 4.26717
R683 source.n552 source.n496 4.26717
R684 source.n448 source.n436 4.26717
R685 source.n478 source.n422 4.26717
R686 source.n382 source.n370 4.26717
R687 source.n412 source.n356 4.26717
R688 source.n308 source.n296 4.26717
R689 source.n338 source.n282 4.26717
R690 source.n58 source.n2 4.26717
R691 source.n29 source.n17 4.26717
R692 source.n132 source.n76 4.26717
R693 source.n103 source.n91 4.26717
R694 source.n198 source.n142 4.26717
R695 source.n169 source.n157 4.26717
R696 source.n272 source.n216 4.26717
R697 source.n243 source.n231 4.26717
R698 source.n526 source.n525 3.49141
R699 source.n551 source.n498 3.49141
R700 source.n452 source.n451 3.49141
R701 source.n477 source.n424 3.49141
R702 source.n386 source.n385 3.49141
R703 source.n411 source.n358 3.49141
R704 source.n312 source.n311 3.49141
R705 source.n337 source.n284 3.49141
R706 source.n57 source.n4 3.49141
R707 source.n33 source.n32 3.49141
R708 source.n131 source.n78 3.49141
R709 source.n107 source.n106 3.49141
R710 source.n197 source.n144 3.49141
R711 source.n173 source.n172 3.49141
R712 source.n271 source.n218 3.49141
R713 source.n247 source.n246 3.49141
R714 source.n516 source.n515 2.84303
R715 source.n442 source.n441 2.84303
R716 source.n376 source.n375 2.84303
R717 source.n302 source.n301 2.84303
R718 source.n23 source.n22 2.84303
R719 source.n97 source.n96 2.84303
R720 source.n163 source.n162 2.84303
R721 source.n237 source.n236 2.84303
R722 source.n529 source.n508 2.71565
R723 source.n548 source.n547 2.71565
R724 source.n455 source.n434 2.71565
R725 source.n474 source.n473 2.71565
R726 source.n389 source.n368 2.71565
R727 source.n408 source.n407 2.71565
R728 source.n315 source.n294 2.71565
R729 source.n334 source.n333 2.71565
R730 source.n54 source.n53 2.71565
R731 source.n36 source.n15 2.71565
R732 source.n128 source.n127 2.71565
R733 source.n110 source.n89 2.71565
R734 source.n194 source.n193 2.71565
R735 source.n176 source.n155 2.71565
R736 source.n268 source.n267 2.71565
R737 source.n250 source.n229 2.71565
R738 source.n530 source.n506 1.93989
R739 source.n544 source.n500 1.93989
R740 source.n456 source.n432 1.93989
R741 source.n470 source.n426 1.93989
R742 source.n390 source.n366 1.93989
R743 source.n404 source.n360 1.93989
R744 source.n316 source.n292 1.93989
R745 source.n330 source.n286 1.93989
R746 source.n50 source.n6 1.93989
R747 source.n37 source.n13 1.93989
R748 source.n124 source.n80 1.93989
R749 source.n111 source.n87 1.93989
R750 source.n190 source.n146 1.93989
R751 source.n177 source.n153 1.93989
R752 source.n264 source.n220 1.93989
R753 source.n251 source.n227 1.93989
R754 source.n492 source.t24 1.6505
R755 source.n492 source.t27 1.6505
R756 source.n490 source.t20 1.6505
R757 source.n490 source.t25 1.6505
R758 source.n488 source.t33 1.6505
R759 source.n488 source.t32 1.6505
R760 source.n486 source.t22 1.6505
R761 source.n486 source.t28 1.6505
R762 source.n352 source.t8 1.6505
R763 source.n352 source.t0 1.6505
R764 source.n350 source.t6 1.6505
R765 source.n350 source.t1 1.6505
R766 source.n348 source.t15 1.6505
R767 source.n348 source.t17 1.6505
R768 source.n346 source.t14 1.6505
R769 source.n346 source.t2 1.6505
R770 source.n66 source.t39 1.6505
R771 source.n66 source.t5 1.6505
R772 source.n68 source.t9 1.6505
R773 source.n68 source.t7 1.6505
R774 source.n70 source.t11 1.6505
R775 source.n70 source.t4 1.6505
R776 source.n72 source.t10 1.6505
R777 source.n72 source.t3 1.6505
R778 source.n206 source.t23 1.6505
R779 source.n206 source.t29 1.6505
R780 source.n208 source.t34 1.6505
R781 source.n208 source.t35 1.6505
R782 source.n210 source.t18 1.6505
R783 source.n210 source.t19 1.6505
R784 source.n212 source.t21 1.6505
R785 source.n212 source.t31 1.6505
R786 source.n535 source.n533 1.16414
R787 source.n543 source.n502 1.16414
R788 source.n461 source.n459 1.16414
R789 source.n469 source.n428 1.16414
R790 source.n395 source.n393 1.16414
R791 source.n403 source.n362 1.16414
R792 source.n321 source.n319 1.16414
R793 source.n329 source.n288 1.16414
R794 source.n49 source.n8 1.16414
R795 source.n41 source.n40 1.16414
R796 source.n123 source.n82 1.16414
R797 source.n115 source.n114 1.16414
R798 source.n189 source.n148 1.16414
R799 source.n181 source.n180 1.16414
R800 source.n263 source.n222 1.16414
R801 source.n255 source.n254 1.16414
R802 source.n205 source.n139 0.470328
R803 source.n485 source.n419 0.470328
R804 source.n279 source.n213 0.457397
R805 source.n213 source.n211 0.457397
R806 source.n211 source.n209 0.457397
R807 source.n209 source.n207 0.457397
R808 source.n207 source.n205 0.457397
R809 source.n139 source.n73 0.457397
R810 source.n73 source.n71 0.457397
R811 source.n71 source.n69 0.457397
R812 source.n69 source.n67 0.457397
R813 source.n67 source.n65 0.457397
R814 source.n347 source.n345 0.457397
R815 source.n349 source.n347 0.457397
R816 source.n351 source.n349 0.457397
R817 source.n353 source.n351 0.457397
R818 source.n419 source.n353 0.457397
R819 source.n487 source.n485 0.457397
R820 source.n489 source.n487 0.457397
R821 source.n491 source.n489 0.457397
R822 source.n493 source.n491 0.457397
R823 source.n559 source.n493 0.457397
R824 source.n534 source.n504 0.388379
R825 source.n540 source.n539 0.388379
R826 source.n460 source.n430 0.388379
R827 source.n466 source.n465 0.388379
R828 source.n394 source.n364 0.388379
R829 source.n400 source.n399 0.388379
R830 source.n320 source.n290 0.388379
R831 source.n326 source.n325 0.388379
R832 source.n46 source.n45 0.388379
R833 source.n12 source.n10 0.388379
R834 source.n120 source.n119 0.388379
R835 source.n86 source.n84 0.388379
R836 source.n186 source.n185 0.388379
R837 source.n152 source.n150 0.388379
R838 source.n260 source.n259 0.388379
R839 source.n226 source.n224 0.388379
R840 source source.n560 0.188
R841 source.n516 source.n511 0.155672
R842 source.n523 source.n511 0.155672
R843 source.n524 source.n523 0.155672
R844 source.n524 source.n507 0.155672
R845 source.n531 source.n507 0.155672
R846 source.n532 source.n531 0.155672
R847 source.n532 source.n503 0.155672
R848 source.n541 source.n503 0.155672
R849 source.n542 source.n541 0.155672
R850 source.n542 source.n499 0.155672
R851 source.n549 source.n499 0.155672
R852 source.n550 source.n549 0.155672
R853 source.n550 source.n495 0.155672
R854 source.n557 source.n495 0.155672
R855 source.n442 source.n437 0.155672
R856 source.n449 source.n437 0.155672
R857 source.n450 source.n449 0.155672
R858 source.n450 source.n433 0.155672
R859 source.n457 source.n433 0.155672
R860 source.n458 source.n457 0.155672
R861 source.n458 source.n429 0.155672
R862 source.n467 source.n429 0.155672
R863 source.n468 source.n467 0.155672
R864 source.n468 source.n425 0.155672
R865 source.n475 source.n425 0.155672
R866 source.n476 source.n475 0.155672
R867 source.n476 source.n421 0.155672
R868 source.n483 source.n421 0.155672
R869 source.n376 source.n371 0.155672
R870 source.n383 source.n371 0.155672
R871 source.n384 source.n383 0.155672
R872 source.n384 source.n367 0.155672
R873 source.n391 source.n367 0.155672
R874 source.n392 source.n391 0.155672
R875 source.n392 source.n363 0.155672
R876 source.n401 source.n363 0.155672
R877 source.n402 source.n401 0.155672
R878 source.n402 source.n359 0.155672
R879 source.n409 source.n359 0.155672
R880 source.n410 source.n409 0.155672
R881 source.n410 source.n355 0.155672
R882 source.n417 source.n355 0.155672
R883 source.n302 source.n297 0.155672
R884 source.n309 source.n297 0.155672
R885 source.n310 source.n309 0.155672
R886 source.n310 source.n293 0.155672
R887 source.n317 source.n293 0.155672
R888 source.n318 source.n317 0.155672
R889 source.n318 source.n289 0.155672
R890 source.n327 source.n289 0.155672
R891 source.n328 source.n327 0.155672
R892 source.n328 source.n285 0.155672
R893 source.n335 source.n285 0.155672
R894 source.n336 source.n335 0.155672
R895 source.n336 source.n281 0.155672
R896 source.n343 source.n281 0.155672
R897 source.n63 source.n1 0.155672
R898 source.n56 source.n1 0.155672
R899 source.n56 source.n55 0.155672
R900 source.n55 source.n5 0.155672
R901 source.n48 source.n5 0.155672
R902 source.n48 source.n47 0.155672
R903 source.n47 source.n9 0.155672
R904 source.n39 source.n9 0.155672
R905 source.n39 source.n38 0.155672
R906 source.n38 source.n14 0.155672
R907 source.n31 source.n14 0.155672
R908 source.n31 source.n30 0.155672
R909 source.n30 source.n18 0.155672
R910 source.n23 source.n18 0.155672
R911 source.n137 source.n75 0.155672
R912 source.n130 source.n75 0.155672
R913 source.n130 source.n129 0.155672
R914 source.n129 source.n79 0.155672
R915 source.n122 source.n79 0.155672
R916 source.n122 source.n121 0.155672
R917 source.n121 source.n83 0.155672
R918 source.n113 source.n83 0.155672
R919 source.n113 source.n112 0.155672
R920 source.n112 source.n88 0.155672
R921 source.n105 source.n88 0.155672
R922 source.n105 source.n104 0.155672
R923 source.n104 source.n92 0.155672
R924 source.n97 source.n92 0.155672
R925 source.n203 source.n141 0.155672
R926 source.n196 source.n141 0.155672
R927 source.n196 source.n195 0.155672
R928 source.n195 source.n145 0.155672
R929 source.n188 source.n145 0.155672
R930 source.n188 source.n187 0.155672
R931 source.n187 source.n149 0.155672
R932 source.n179 source.n149 0.155672
R933 source.n179 source.n178 0.155672
R934 source.n178 source.n154 0.155672
R935 source.n171 source.n154 0.155672
R936 source.n171 source.n170 0.155672
R937 source.n170 source.n158 0.155672
R938 source.n163 source.n158 0.155672
R939 source.n277 source.n215 0.155672
R940 source.n270 source.n215 0.155672
R941 source.n270 source.n269 0.155672
R942 source.n269 source.n219 0.155672
R943 source.n262 source.n219 0.155672
R944 source.n262 source.n261 0.155672
R945 source.n261 source.n223 0.155672
R946 source.n253 source.n223 0.155672
R947 source.n253 source.n252 0.155672
R948 source.n252 source.n228 0.155672
R949 source.n245 source.n228 0.155672
R950 source.n245 source.n244 0.155672
R951 source.n244 source.n232 0.155672
R952 source.n237 source.n232 0.155672
R953 drain_right.n6 drain_right.n4 60.0094
R954 drain_right.n2 drain_right.n0 60.0094
R955 drain_right.n10 drain_right.n8 60.0094
R956 drain_right.n10 drain_right.n9 59.5527
R957 drain_right.n12 drain_right.n11 59.5527
R958 drain_right.n14 drain_right.n13 59.5527
R959 drain_right.n16 drain_right.n15 59.5527
R960 drain_right.n7 drain_right.n3 59.5525
R961 drain_right.n6 drain_right.n5 59.5525
R962 drain_right.n2 drain_right.n1 59.5525
R963 drain_right drain_right.n7 30.469
R964 drain_right drain_right.n16 6.11011
R965 drain_right.n3 drain_right.t5 1.6505
R966 drain_right.n3 drain_right.t11 1.6505
R967 drain_right.n4 drain_right.t8 1.6505
R968 drain_right.n4 drain_right.t15 1.6505
R969 drain_right.n5 drain_right.t6 1.6505
R970 drain_right.n5 drain_right.t12 1.6505
R971 drain_right.n1 drain_right.t17 1.6505
R972 drain_right.n1 drain_right.t14 1.6505
R973 drain_right.n0 drain_right.t16 1.6505
R974 drain_right.n0 drain_right.t13 1.6505
R975 drain_right.n8 drain_right.t9 1.6505
R976 drain_right.n8 drain_right.t3 1.6505
R977 drain_right.n9 drain_right.t1 1.6505
R978 drain_right.n9 drain_right.t19 1.6505
R979 drain_right.n11 drain_right.t10 1.6505
R980 drain_right.n11 drain_right.t2 1.6505
R981 drain_right.n13 drain_right.t0 1.6505
R982 drain_right.n13 drain_right.t18 1.6505
R983 drain_right.n15 drain_right.t7 1.6505
R984 drain_right.n15 drain_right.t4 1.6505
R985 drain_right.n16 drain_right.n14 0.457397
R986 drain_right.n14 drain_right.n12 0.457397
R987 drain_right.n12 drain_right.n10 0.457397
R988 drain_right.n7 drain_right.n6 0.402051
R989 drain_right.n7 drain_right.n2 0.402051
R990 plus.n5 plus.t5 1658.88
R991 plus.n23 plus.t2 1658.88
R992 plus.n30 plus.t16 1658.88
R993 plus.n48 plus.t3 1658.88
R994 plus.n6 plus.t1 1602.65
R995 plus.n8 plus.t18 1602.65
R996 plus.n3 plus.t12 1602.65
R997 plus.n13 plus.t11 1602.65
R998 plus.n15 plus.t4 1602.65
R999 plus.n1 plus.t0 1602.65
R1000 plus.n20 plus.t17 1602.65
R1001 plus.n22 plus.t9 1602.65
R1002 plus.n31 plus.t19 1602.65
R1003 plus.n33 plus.t14 1602.65
R1004 plus.n28 plus.t10 1602.65
R1005 plus.n38 plus.t15 1602.65
R1006 plus.n40 plus.t7 1602.65
R1007 plus.n26 plus.t13 1602.65
R1008 plus.n45 plus.t8 1602.65
R1009 plus.n47 plus.t6 1602.65
R1010 plus.n5 plus.n4 161.489
R1011 plus.n30 plus.n29 161.489
R1012 plus.n7 plus.n4 161.3
R1013 plus.n10 plus.n9 161.3
R1014 plus.n12 plus.n11 161.3
R1015 plus.n14 plus.n2 161.3
R1016 plus.n17 plus.n16 161.3
R1017 plus.n19 plus.n18 161.3
R1018 plus.n21 plus.n0 161.3
R1019 plus.n24 plus.n23 161.3
R1020 plus.n32 plus.n29 161.3
R1021 plus.n35 plus.n34 161.3
R1022 plus.n37 plus.n36 161.3
R1023 plus.n39 plus.n27 161.3
R1024 plus.n42 plus.n41 161.3
R1025 plus.n44 plus.n43 161.3
R1026 plus.n46 plus.n25 161.3
R1027 plus.n49 plus.n48 161.3
R1028 plus.n7 plus.n6 51.852
R1029 plus.n22 plus.n21 51.852
R1030 plus.n47 plus.n46 51.852
R1031 plus.n32 plus.n31 51.852
R1032 plus.n9 plus.n8 47.4702
R1033 plus.n20 plus.n19 47.4702
R1034 plus.n45 plus.n44 47.4702
R1035 plus.n34 plus.n33 47.4702
R1036 plus.n12 plus.n3 43.0884
R1037 plus.n16 plus.n1 43.0884
R1038 plus.n41 plus.n26 43.0884
R1039 plus.n37 plus.n28 43.0884
R1040 plus.n14 plus.n13 38.7066
R1041 plus.n15 plus.n14 38.7066
R1042 plus.n40 plus.n39 38.7066
R1043 plus.n39 plus.n38 38.7066
R1044 plus.n13 plus.n12 34.3247
R1045 plus.n16 plus.n15 34.3247
R1046 plus.n41 plus.n40 34.3247
R1047 plus.n38 plus.n37 34.3247
R1048 plus plus.n49 30.1089
R1049 plus.n9 plus.n3 29.9429
R1050 plus.n19 plus.n1 29.9429
R1051 plus.n44 plus.n26 29.9429
R1052 plus.n34 plus.n28 29.9429
R1053 plus.n8 plus.n7 25.5611
R1054 plus.n21 plus.n20 25.5611
R1055 plus.n46 plus.n45 25.5611
R1056 plus.n33 plus.n32 25.5611
R1057 plus.n6 plus.n5 21.1793
R1058 plus.n23 plus.n22 21.1793
R1059 plus.n48 plus.n47 21.1793
R1060 plus.n31 plus.n30 21.1793
R1061 plus plus.n24 12.1217
R1062 plus.n10 plus.n4 0.189894
R1063 plus.n11 plus.n10 0.189894
R1064 plus.n11 plus.n2 0.189894
R1065 plus.n17 plus.n2 0.189894
R1066 plus.n18 plus.n17 0.189894
R1067 plus.n18 plus.n0 0.189894
R1068 plus.n24 plus.n0 0.189894
R1069 plus.n49 plus.n25 0.189894
R1070 plus.n43 plus.n25 0.189894
R1071 plus.n43 plus.n42 0.189894
R1072 plus.n42 plus.n27 0.189894
R1073 plus.n36 plus.n27 0.189894
R1074 plus.n36 plus.n35 0.189894
R1075 plus.n35 plus.n29 0.189894
R1076 drain_left.n10 drain_left.n8 60.0096
R1077 drain_left.n6 drain_left.n4 60.0094
R1078 drain_left.n2 drain_left.n0 60.0094
R1079 drain_left.n14 drain_left.n13 59.5527
R1080 drain_left.n12 drain_left.n11 59.5527
R1081 drain_left.n10 drain_left.n9 59.5527
R1082 drain_left.n7 drain_left.n3 59.5525
R1083 drain_left.n6 drain_left.n5 59.5525
R1084 drain_left.n2 drain_left.n1 59.5525
R1085 drain_left.n16 drain_left.n15 59.5525
R1086 drain_left drain_left.n7 31.0222
R1087 drain_left drain_left.n16 6.11011
R1088 drain_left.n3 drain_left.t12 1.6505
R1089 drain_left.n3 drain_left.t4 1.6505
R1090 drain_left.n4 drain_left.t0 1.6505
R1091 drain_left.n4 drain_left.t3 1.6505
R1092 drain_left.n5 drain_left.t9 1.6505
R1093 drain_left.n5 drain_left.t5 1.6505
R1094 drain_left.n1 drain_left.t11 1.6505
R1095 drain_left.n1 drain_left.t6 1.6505
R1096 drain_left.n0 drain_left.t16 1.6505
R1097 drain_left.n0 drain_left.t13 1.6505
R1098 drain_left.n15 drain_left.t10 1.6505
R1099 drain_left.n15 drain_left.t17 1.6505
R1100 drain_left.n13 drain_left.t19 1.6505
R1101 drain_left.n13 drain_left.t2 1.6505
R1102 drain_left.n11 drain_left.t8 1.6505
R1103 drain_left.n11 drain_left.t15 1.6505
R1104 drain_left.n9 drain_left.t1 1.6505
R1105 drain_left.n9 drain_left.t7 1.6505
R1106 drain_left.n8 drain_left.t14 1.6505
R1107 drain_left.n8 drain_left.t18 1.6505
R1108 drain_left.n12 drain_left.n10 0.457397
R1109 drain_left.n14 drain_left.n12 0.457397
R1110 drain_left.n16 drain_left.n14 0.457397
R1111 drain_left.n7 drain_left.n6 0.402051
R1112 drain_left.n7 drain_left.n2 0.402051
C0 plus source 4.97249f
C1 minus source 4.95845f
C2 drain_right source 45.2007f
C3 drain_left plus 5.5063f
C4 drain_left minus 0.171252f
C5 drain_right drain_left 0.982035f
C6 plus minus 5.50167f
C7 drain_right plus 0.337271f
C8 drain_right minus 5.32325f
C9 drain_left source 45.2007f
C10 drain_right a_n1882_n3288# 7.1215f
C11 drain_left a_n1882_n3288# 7.42292f
C12 source a_n1882_n3288# 8.614861f
C13 minus a_n1882_n3288# 7.311454f
C14 plus a_n1882_n3288# 9.402691f
C15 drain_left.t16 a_n1882_n3288# 0.369075f
C16 drain_left.t13 a_n1882_n3288# 0.369075f
C17 drain_left.n0 a_n1882_n3288# 3.28767f
C18 drain_left.t11 a_n1882_n3288# 0.369075f
C19 drain_left.t6 a_n1882_n3288# 0.369075f
C20 drain_left.n1 a_n1882_n3288# 3.2842f
C21 drain_left.n2 a_n1882_n3288# 0.889989f
C22 drain_left.t12 a_n1882_n3288# 0.369075f
C23 drain_left.t4 a_n1882_n3288# 0.369075f
C24 drain_left.n3 a_n1882_n3288# 3.2842f
C25 drain_left.t0 a_n1882_n3288# 0.369075f
C26 drain_left.t3 a_n1882_n3288# 0.369075f
C27 drain_left.n4 a_n1882_n3288# 3.28767f
C28 drain_left.t9 a_n1882_n3288# 0.369075f
C29 drain_left.t5 a_n1882_n3288# 0.369075f
C30 drain_left.n5 a_n1882_n3288# 3.2842f
C31 drain_left.n6 a_n1882_n3288# 0.889989f
C32 drain_left.n7 a_n1882_n3288# 2.30034f
C33 drain_left.t14 a_n1882_n3288# 0.369075f
C34 drain_left.t18 a_n1882_n3288# 0.369075f
C35 drain_left.n8 a_n1882_n3288# 3.28769f
C36 drain_left.t1 a_n1882_n3288# 0.369075f
C37 drain_left.t7 a_n1882_n3288# 0.369075f
C38 drain_left.n9 a_n1882_n3288# 3.28421f
C39 drain_left.n10 a_n1882_n3288# 0.894656f
C40 drain_left.t8 a_n1882_n3288# 0.369075f
C41 drain_left.t15 a_n1882_n3288# 0.369075f
C42 drain_left.n11 a_n1882_n3288# 3.28421f
C43 drain_left.n12 a_n1882_n3288# 0.441229f
C44 drain_left.t19 a_n1882_n3288# 0.369075f
C45 drain_left.t2 a_n1882_n3288# 0.369075f
C46 drain_left.n13 a_n1882_n3288# 3.28421f
C47 drain_left.n14 a_n1882_n3288# 0.441229f
C48 drain_left.t10 a_n1882_n3288# 0.369075f
C49 drain_left.t17 a_n1882_n3288# 0.369075f
C50 drain_left.n15 a_n1882_n3288# 3.2842f
C51 drain_left.n16 a_n1882_n3288# 0.759771f
C52 plus.n0 a_n1882_n3288# 0.053677f
C53 plus.t9 a_n1882_n3288# 0.36404f
C54 plus.t17 a_n1882_n3288# 0.36404f
C55 plus.t0 a_n1882_n3288# 0.36404f
C56 plus.n1 a_n1882_n3288# 0.149928f
C57 plus.n2 a_n1882_n3288# 0.053677f
C58 plus.t4 a_n1882_n3288# 0.36404f
C59 plus.t11 a_n1882_n3288# 0.36404f
C60 plus.t12 a_n1882_n3288# 0.36404f
C61 plus.n3 a_n1882_n3288# 0.149928f
C62 plus.n4 a_n1882_n3288# 0.122828f
C63 plus.t18 a_n1882_n3288# 0.36404f
C64 plus.t1 a_n1882_n3288# 0.36404f
C65 plus.t5 a_n1882_n3288# 0.369217f
C66 plus.n5 a_n1882_n3288# 0.166444f
C67 plus.n6 a_n1882_n3288# 0.149928f
C68 plus.n7 a_n1882_n3288# 0.018799f
C69 plus.n8 a_n1882_n3288# 0.149928f
C70 plus.n9 a_n1882_n3288# 0.018799f
C71 plus.n10 a_n1882_n3288# 0.053677f
C72 plus.n11 a_n1882_n3288# 0.053677f
C73 plus.n12 a_n1882_n3288# 0.018799f
C74 plus.n13 a_n1882_n3288# 0.149928f
C75 plus.n14 a_n1882_n3288# 0.018799f
C76 plus.n15 a_n1882_n3288# 0.149928f
C77 plus.n16 a_n1882_n3288# 0.018799f
C78 plus.n17 a_n1882_n3288# 0.053677f
C79 plus.n18 a_n1882_n3288# 0.053677f
C80 plus.n19 a_n1882_n3288# 0.018799f
C81 plus.n20 a_n1882_n3288# 0.149928f
C82 plus.n21 a_n1882_n3288# 0.018799f
C83 plus.n22 a_n1882_n3288# 0.149928f
C84 plus.t2 a_n1882_n3288# 0.369217f
C85 plus.n23 a_n1882_n3288# 0.166363f
C86 plus.n24 a_n1882_n3288# 0.597716f
C87 plus.n25 a_n1882_n3288# 0.053677f
C88 plus.t3 a_n1882_n3288# 0.369217f
C89 plus.t6 a_n1882_n3288# 0.36404f
C90 plus.t8 a_n1882_n3288# 0.36404f
C91 plus.t13 a_n1882_n3288# 0.36404f
C92 plus.n26 a_n1882_n3288# 0.149928f
C93 plus.n27 a_n1882_n3288# 0.053677f
C94 plus.t7 a_n1882_n3288# 0.36404f
C95 plus.t15 a_n1882_n3288# 0.36404f
C96 plus.t10 a_n1882_n3288# 0.36404f
C97 plus.n28 a_n1882_n3288# 0.149928f
C98 plus.n29 a_n1882_n3288# 0.122828f
C99 plus.t14 a_n1882_n3288# 0.36404f
C100 plus.t19 a_n1882_n3288# 0.36404f
C101 plus.t16 a_n1882_n3288# 0.369217f
C102 plus.n30 a_n1882_n3288# 0.166444f
C103 plus.n31 a_n1882_n3288# 0.149928f
C104 plus.n32 a_n1882_n3288# 0.018799f
C105 plus.n33 a_n1882_n3288# 0.149928f
C106 plus.n34 a_n1882_n3288# 0.018799f
C107 plus.n35 a_n1882_n3288# 0.053677f
C108 plus.n36 a_n1882_n3288# 0.053677f
C109 plus.n37 a_n1882_n3288# 0.018799f
C110 plus.n38 a_n1882_n3288# 0.149928f
C111 plus.n39 a_n1882_n3288# 0.018799f
C112 plus.n40 a_n1882_n3288# 0.149928f
C113 plus.n41 a_n1882_n3288# 0.018799f
C114 plus.n42 a_n1882_n3288# 0.053677f
C115 plus.n43 a_n1882_n3288# 0.053677f
C116 plus.n44 a_n1882_n3288# 0.018799f
C117 plus.n45 a_n1882_n3288# 0.149928f
C118 plus.n46 a_n1882_n3288# 0.018799f
C119 plus.n47 a_n1882_n3288# 0.149928f
C120 plus.n48 a_n1882_n3288# 0.166363f
C121 plus.n49 a_n1882_n3288# 1.60573f
C122 drain_right.t16 a_n1882_n3288# 0.368726f
C123 drain_right.t13 a_n1882_n3288# 0.368726f
C124 drain_right.n0 a_n1882_n3288# 3.28457f
C125 drain_right.t17 a_n1882_n3288# 0.368726f
C126 drain_right.t14 a_n1882_n3288# 0.368726f
C127 drain_right.n1 a_n1882_n3288# 3.28109f
C128 drain_right.n2 a_n1882_n3288# 0.889149f
C129 drain_right.t5 a_n1882_n3288# 0.368726f
C130 drain_right.t11 a_n1882_n3288# 0.368726f
C131 drain_right.n3 a_n1882_n3288# 3.28109f
C132 drain_right.t8 a_n1882_n3288# 0.368726f
C133 drain_right.t15 a_n1882_n3288# 0.368726f
C134 drain_right.n4 a_n1882_n3288# 3.28457f
C135 drain_right.t6 a_n1882_n3288# 0.368726f
C136 drain_right.t12 a_n1882_n3288# 0.368726f
C137 drain_right.n5 a_n1882_n3288# 3.28109f
C138 drain_right.n6 a_n1882_n3288# 0.889149f
C139 drain_right.n7 a_n1882_n3288# 2.21759f
C140 drain_right.t9 a_n1882_n3288# 0.368726f
C141 drain_right.t3 a_n1882_n3288# 0.368726f
C142 drain_right.n8 a_n1882_n3288# 3.28457f
C143 drain_right.t1 a_n1882_n3288# 0.368726f
C144 drain_right.t19 a_n1882_n3288# 0.368726f
C145 drain_right.n9 a_n1882_n3288# 3.28111f
C146 drain_right.n10 a_n1882_n3288# 0.893825f
C147 drain_right.t10 a_n1882_n3288# 0.368726f
C148 drain_right.t2 a_n1882_n3288# 0.368726f
C149 drain_right.n11 a_n1882_n3288# 3.28111f
C150 drain_right.n12 a_n1882_n3288# 0.440813f
C151 drain_right.t0 a_n1882_n3288# 0.368726f
C152 drain_right.t18 a_n1882_n3288# 0.368726f
C153 drain_right.n13 a_n1882_n3288# 3.28111f
C154 drain_right.n14 a_n1882_n3288# 0.440813f
C155 drain_right.t7 a_n1882_n3288# 0.368726f
C156 drain_right.t4 a_n1882_n3288# 0.368726f
C157 drain_right.n15 a_n1882_n3288# 3.28111f
C158 drain_right.n16 a_n1882_n3288# 0.75904f
C159 source.n0 a_n1882_n3288# 0.044563f
C160 source.n1 a_n1882_n3288# 0.033642f
C161 source.n2 a_n1882_n3288# 0.018078f
C162 source.n3 a_n1882_n3288# 0.042729f
C163 source.n4 a_n1882_n3288# 0.019141f
C164 source.n5 a_n1882_n3288# 0.033642f
C165 source.n6 a_n1882_n3288# 0.018078f
C166 source.n7 a_n1882_n3288# 0.042729f
C167 source.n8 a_n1882_n3288# 0.019141f
C168 source.n9 a_n1882_n3288# 0.033642f
C169 source.n10 a_n1882_n3288# 0.018609f
C170 source.n11 a_n1882_n3288# 0.042729f
C171 source.n12 a_n1882_n3288# 0.018078f
C172 source.n13 a_n1882_n3288# 0.019141f
C173 source.n14 a_n1882_n3288# 0.033642f
C174 source.n15 a_n1882_n3288# 0.018078f
C175 source.n16 a_n1882_n3288# 0.042729f
C176 source.n17 a_n1882_n3288# 0.019141f
C177 source.n18 a_n1882_n3288# 0.033642f
C178 source.n19 a_n1882_n3288# 0.018078f
C179 source.n20 a_n1882_n3288# 0.032047f
C180 source.n21 a_n1882_n3288# 0.030206f
C181 source.t12 a_n1882_n3288# 0.072167f
C182 source.n22 a_n1882_n3288# 0.242554f
C183 source.n23 a_n1882_n3288# 1.69718f
C184 source.n24 a_n1882_n3288# 0.018078f
C185 source.n25 a_n1882_n3288# 0.019141f
C186 source.n26 a_n1882_n3288# 0.042729f
C187 source.n27 a_n1882_n3288# 0.042729f
C188 source.n28 a_n1882_n3288# 0.019141f
C189 source.n29 a_n1882_n3288# 0.018078f
C190 source.n30 a_n1882_n3288# 0.033642f
C191 source.n31 a_n1882_n3288# 0.033642f
C192 source.n32 a_n1882_n3288# 0.018078f
C193 source.n33 a_n1882_n3288# 0.019141f
C194 source.n34 a_n1882_n3288# 0.042729f
C195 source.n35 a_n1882_n3288# 0.042729f
C196 source.n36 a_n1882_n3288# 0.019141f
C197 source.n37 a_n1882_n3288# 0.018078f
C198 source.n38 a_n1882_n3288# 0.033642f
C199 source.n39 a_n1882_n3288# 0.033642f
C200 source.n40 a_n1882_n3288# 0.018078f
C201 source.n41 a_n1882_n3288# 0.019141f
C202 source.n42 a_n1882_n3288# 0.042729f
C203 source.n43 a_n1882_n3288# 0.042729f
C204 source.n44 a_n1882_n3288# 0.042729f
C205 source.n45 a_n1882_n3288# 0.018609f
C206 source.n46 a_n1882_n3288# 0.018078f
C207 source.n47 a_n1882_n3288# 0.033642f
C208 source.n48 a_n1882_n3288# 0.033642f
C209 source.n49 a_n1882_n3288# 0.018078f
C210 source.n50 a_n1882_n3288# 0.019141f
C211 source.n51 a_n1882_n3288# 0.042729f
C212 source.n52 a_n1882_n3288# 0.042729f
C213 source.n53 a_n1882_n3288# 0.019141f
C214 source.n54 a_n1882_n3288# 0.018078f
C215 source.n55 a_n1882_n3288# 0.033642f
C216 source.n56 a_n1882_n3288# 0.033642f
C217 source.n57 a_n1882_n3288# 0.018078f
C218 source.n58 a_n1882_n3288# 0.019141f
C219 source.n59 a_n1882_n3288# 0.042729f
C220 source.n60 a_n1882_n3288# 0.087685f
C221 source.n61 a_n1882_n3288# 0.019141f
C222 source.n62 a_n1882_n3288# 0.018078f
C223 source.n63 a_n1882_n3288# 0.072247f
C224 source.n64 a_n1882_n3288# 0.048392f
C225 source.n65 a_n1882_n3288# 1.33858f
C226 source.t39 a_n1882_n3288# 0.319019f
C227 source.t5 a_n1882_n3288# 0.319019f
C228 source.n66 a_n1882_n3288# 2.73144f
C229 source.n67 a_n1882_n3288# 0.443003f
C230 source.t9 a_n1882_n3288# 0.319019f
C231 source.t7 a_n1882_n3288# 0.319019f
C232 source.n68 a_n1882_n3288# 2.73144f
C233 source.n69 a_n1882_n3288# 0.443003f
C234 source.t11 a_n1882_n3288# 0.319019f
C235 source.t4 a_n1882_n3288# 0.319019f
C236 source.n70 a_n1882_n3288# 2.73144f
C237 source.n71 a_n1882_n3288# 0.443003f
C238 source.t10 a_n1882_n3288# 0.319019f
C239 source.t3 a_n1882_n3288# 0.319019f
C240 source.n72 a_n1882_n3288# 2.73144f
C241 source.n73 a_n1882_n3288# 0.443003f
C242 source.n74 a_n1882_n3288# 0.044563f
C243 source.n75 a_n1882_n3288# 0.033642f
C244 source.n76 a_n1882_n3288# 0.018078f
C245 source.n77 a_n1882_n3288# 0.042729f
C246 source.n78 a_n1882_n3288# 0.019141f
C247 source.n79 a_n1882_n3288# 0.033642f
C248 source.n80 a_n1882_n3288# 0.018078f
C249 source.n81 a_n1882_n3288# 0.042729f
C250 source.n82 a_n1882_n3288# 0.019141f
C251 source.n83 a_n1882_n3288# 0.033642f
C252 source.n84 a_n1882_n3288# 0.018609f
C253 source.n85 a_n1882_n3288# 0.042729f
C254 source.n86 a_n1882_n3288# 0.018078f
C255 source.n87 a_n1882_n3288# 0.019141f
C256 source.n88 a_n1882_n3288# 0.033642f
C257 source.n89 a_n1882_n3288# 0.018078f
C258 source.n90 a_n1882_n3288# 0.042729f
C259 source.n91 a_n1882_n3288# 0.019141f
C260 source.n92 a_n1882_n3288# 0.033642f
C261 source.n93 a_n1882_n3288# 0.018078f
C262 source.n94 a_n1882_n3288# 0.032047f
C263 source.n95 a_n1882_n3288# 0.030206f
C264 source.t13 a_n1882_n3288# 0.072167f
C265 source.n96 a_n1882_n3288# 0.242554f
C266 source.n97 a_n1882_n3288# 1.69718f
C267 source.n98 a_n1882_n3288# 0.018078f
C268 source.n99 a_n1882_n3288# 0.019141f
C269 source.n100 a_n1882_n3288# 0.042729f
C270 source.n101 a_n1882_n3288# 0.042729f
C271 source.n102 a_n1882_n3288# 0.019141f
C272 source.n103 a_n1882_n3288# 0.018078f
C273 source.n104 a_n1882_n3288# 0.033642f
C274 source.n105 a_n1882_n3288# 0.033642f
C275 source.n106 a_n1882_n3288# 0.018078f
C276 source.n107 a_n1882_n3288# 0.019141f
C277 source.n108 a_n1882_n3288# 0.042729f
C278 source.n109 a_n1882_n3288# 0.042729f
C279 source.n110 a_n1882_n3288# 0.019141f
C280 source.n111 a_n1882_n3288# 0.018078f
C281 source.n112 a_n1882_n3288# 0.033642f
C282 source.n113 a_n1882_n3288# 0.033642f
C283 source.n114 a_n1882_n3288# 0.018078f
C284 source.n115 a_n1882_n3288# 0.019141f
C285 source.n116 a_n1882_n3288# 0.042729f
C286 source.n117 a_n1882_n3288# 0.042729f
C287 source.n118 a_n1882_n3288# 0.042729f
C288 source.n119 a_n1882_n3288# 0.018609f
C289 source.n120 a_n1882_n3288# 0.018078f
C290 source.n121 a_n1882_n3288# 0.033642f
C291 source.n122 a_n1882_n3288# 0.033642f
C292 source.n123 a_n1882_n3288# 0.018078f
C293 source.n124 a_n1882_n3288# 0.019141f
C294 source.n125 a_n1882_n3288# 0.042729f
C295 source.n126 a_n1882_n3288# 0.042729f
C296 source.n127 a_n1882_n3288# 0.019141f
C297 source.n128 a_n1882_n3288# 0.018078f
C298 source.n129 a_n1882_n3288# 0.033642f
C299 source.n130 a_n1882_n3288# 0.033642f
C300 source.n131 a_n1882_n3288# 0.018078f
C301 source.n132 a_n1882_n3288# 0.019141f
C302 source.n133 a_n1882_n3288# 0.042729f
C303 source.n134 a_n1882_n3288# 0.087685f
C304 source.n135 a_n1882_n3288# 0.019141f
C305 source.n136 a_n1882_n3288# 0.018078f
C306 source.n137 a_n1882_n3288# 0.072247f
C307 source.n138 a_n1882_n3288# 0.048392f
C308 source.n139 a_n1882_n3288# 0.126085f
C309 source.n140 a_n1882_n3288# 0.044563f
C310 source.n141 a_n1882_n3288# 0.033642f
C311 source.n142 a_n1882_n3288# 0.018078f
C312 source.n143 a_n1882_n3288# 0.042729f
C313 source.n144 a_n1882_n3288# 0.019141f
C314 source.n145 a_n1882_n3288# 0.033642f
C315 source.n146 a_n1882_n3288# 0.018078f
C316 source.n147 a_n1882_n3288# 0.042729f
C317 source.n148 a_n1882_n3288# 0.019141f
C318 source.n149 a_n1882_n3288# 0.033642f
C319 source.n150 a_n1882_n3288# 0.018609f
C320 source.n151 a_n1882_n3288# 0.042729f
C321 source.n152 a_n1882_n3288# 0.018078f
C322 source.n153 a_n1882_n3288# 0.019141f
C323 source.n154 a_n1882_n3288# 0.033642f
C324 source.n155 a_n1882_n3288# 0.018078f
C325 source.n156 a_n1882_n3288# 0.042729f
C326 source.n157 a_n1882_n3288# 0.019141f
C327 source.n158 a_n1882_n3288# 0.033642f
C328 source.n159 a_n1882_n3288# 0.018078f
C329 source.n160 a_n1882_n3288# 0.032047f
C330 source.n161 a_n1882_n3288# 0.030206f
C331 source.t30 a_n1882_n3288# 0.072167f
C332 source.n162 a_n1882_n3288# 0.242554f
C333 source.n163 a_n1882_n3288# 1.69718f
C334 source.n164 a_n1882_n3288# 0.018078f
C335 source.n165 a_n1882_n3288# 0.019141f
C336 source.n166 a_n1882_n3288# 0.042729f
C337 source.n167 a_n1882_n3288# 0.042729f
C338 source.n168 a_n1882_n3288# 0.019141f
C339 source.n169 a_n1882_n3288# 0.018078f
C340 source.n170 a_n1882_n3288# 0.033642f
C341 source.n171 a_n1882_n3288# 0.033642f
C342 source.n172 a_n1882_n3288# 0.018078f
C343 source.n173 a_n1882_n3288# 0.019141f
C344 source.n174 a_n1882_n3288# 0.042729f
C345 source.n175 a_n1882_n3288# 0.042729f
C346 source.n176 a_n1882_n3288# 0.019141f
C347 source.n177 a_n1882_n3288# 0.018078f
C348 source.n178 a_n1882_n3288# 0.033642f
C349 source.n179 a_n1882_n3288# 0.033642f
C350 source.n180 a_n1882_n3288# 0.018078f
C351 source.n181 a_n1882_n3288# 0.019141f
C352 source.n182 a_n1882_n3288# 0.042729f
C353 source.n183 a_n1882_n3288# 0.042729f
C354 source.n184 a_n1882_n3288# 0.042729f
C355 source.n185 a_n1882_n3288# 0.018609f
C356 source.n186 a_n1882_n3288# 0.018078f
C357 source.n187 a_n1882_n3288# 0.033642f
C358 source.n188 a_n1882_n3288# 0.033642f
C359 source.n189 a_n1882_n3288# 0.018078f
C360 source.n190 a_n1882_n3288# 0.019141f
C361 source.n191 a_n1882_n3288# 0.042729f
C362 source.n192 a_n1882_n3288# 0.042729f
C363 source.n193 a_n1882_n3288# 0.019141f
C364 source.n194 a_n1882_n3288# 0.018078f
C365 source.n195 a_n1882_n3288# 0.033642f
C366 source.n196 a_n1882_n3288# 0.033642f
C367 source.n197 a_n1882_n3288# 0.018078f
C368 source.n198 a_n1882_n3288# 0.019141f
C369 source.n199 a_n1882_n3288# 0.042729f
C370 source.n200 a_n1882_n3288# 0.087685f
C371 source.n201 a_n1882_n3288# 0.019141f
C372 source.n202 a_n1882_n3288# 0.018078f
C373 source.n203 a_n1882_n3288# 0.072247f
C374 source.n204 a_n1882_n3288# 0.048392f
C375 source.n205 a_n1882_n3288# 0.126085f
C376 source.t23 a_n1882_n3288# 0.319019f
C377 source.t29 a_n1882_n3288# 0.319019f
C378 source.n206 a_n1882_n3288# 2.73144f
C379 source.n207 a_n1882_n3288# 0.443003f
C380 source.t34 a_n1882_n3288# 0.319019f
C381 source.t35 a_n1882_n3288# 0.319019f
C382 source.n208 a_n1882_n3288# 2.73144f
C383 source.n209 a_n1882_n3288# 0.443003f
C384 source.t18 a_n1882_n3288# 0.319019f
C385 source.t19 a_n1882_n3288# 0.319019f
C386 source.n210 a_n1882_n3288# 2.73144f
C387 source.n211 a_n1882_n3288# 0.443003f
C388 source.t21 a_n1882_n3288# 0.319019f
C389 source.t31 a_n1882_n3288# 0.319019f
C390 source.n212 a_n1882_n3288# 2.73144f
C391 source.n213 a_n1882_n3288# 0.443003f
C392 source.n214 a_n1882_n3288# 0.044563f
C393 source.n215 a_n1882_n3288# 0.033642f
C394 source.n216 a_n1882_n3288# 0.018078f
C395 source.n217 a_n1882_n3288# 0.042729f
C396 source.n218 a_n1882_n3288# 0.019141f
C397 source.n219 a_n1882_n3288# 0.033642f
C398 source.n220 a_n1882_n3288# 0.018078f
C399 source.n221 a_n1882_n3288# 0.042729f
C400 source.n222 a_n1882_n3288# 0.019141f
C401 source.n223 a_n1882_n3288# 0.033642f
C402 source.n224 a_n1882_n3288# 0.018609f
C403 source.n225 a_n1882_n3288# 0.042729f
C404 source.n226 a_n1882_n3288# 0.018078f
C405 source.n227 a_n1882_n3288# 0.019141f
C406 source.n228 a_n1882_n3288# 0.033642f
C407 source.n229 a_n1882_n3288# 0.018078f
C408 source.n230 a_n1882_n3288# 0.042729f
C409 source.n231 a_n1882_n3288# 0.019141f
C410 source.n232 a_n1882_n3288# 0.033642f
C411 source.n233 a_n1882_n3288# 0.018078f
C412 source.n234 a_n1882_n3288# 0.032047f
C413 source.n235 a_n1882_n3288# 0.030206f
C414 source.t37 a_n1882_n3288# 0.072167f
C415 source.n236 a_n1882_n3288# 0.242554f
C416 source.n237 a_n1882_n3288# 1.69718f
C417 source.n238 a_n1882_n3288# 0.018078f
C418 source.n239 a_n1882_n3288# 0.019141f
C419 source.n240 a_n1882_n3288# 0.042729f
C420 source.n241 a_n1882_n3288# 0.042729f
C421 source.n242 a_n1882_n3288# 0.019141f
C422 source.n243 a_n1882_n3288# 0.018078f
C423 source.n244 a_n1882_n3288# 0.033642f
C424 source.n245 a_n1882_n3288# 0.033642f
C425 source.n246 a_n1882_n3288# 0.018078f
C426 source.n247 a_n1882_n3288# 0.019141f
C427 source.n248 a_n1882_n3288# 0.042729f
C428 source.n249 a_n1882_n3288# 0.042729f
C429 source.n250 a_n1882_n3288# 0.019141f
C430 source.n251 a_n1882_n3288# 0.018078f
C431 source.n252 a_n1882_n3288# 0.033642f
C432 source.n253 a_n1882_n3288# 0.033642f
C433 source.n254 a_n1882_n3288# 0.018078f
C434 source.n255 a_n1882_n3288# 0.019141f
C435 source.n256 a_n1882_n3288# 0.042729f
C436 source.n257 a_n1882_n3288# 0.042729f
C437 source.n258 a_n1882_n3288# 0.042729f
C438 source.n259 a_n1882_n3288# 0.018609f
C439 source.n260 a_n1882_n3288# 0.018078f
C440 source.n261 a_n1882_n3288# 0.033642f
C441 source.n262 a_n1882_n3288# 0.033642f
C442 source.n263 a_n1882_n3288# 0.018078f
C443 source.n264 a_n1882_n3288# 0.019141f
C444 source.n265 a_n1882_n3288# 0.042729f
C445 source.n266 a_n1882_n3288# 0.042729f
C446 source.n267 a_n1882_n3288# 0.019141f
C447 source.n268 a_n1882_n3288# 0.018078f
C448 source.n269 a_n1882_n3288# 0.033642f
C449 source.n270 a_n1882_n3288# 0.033642f
C450 source.n271 a_n1882_n3288# 0.018078f
C451 source.n272 a_n1882_n3288# 0.019141f
C452 source.n273 a_n1882_n3288# 0.042729f
C453 source.n274 a_n1882_n3288# 0.087685f
C454 source.n275 a_n1882_n3288# 0.019141f
C455 source.n276 a_n1882_n3288# 0.018078f
C456 source.n277 a_n1882_n3288# 0.072247f
C457 source.n278 a_n1882_n3288# 0.048392f
C458 source.n279 a_n1882_n3288# 1.86422f
C459 source.n280 a_n1882_n3288# 0.044563f
C460 source.n281 a_n1882_n3288# 0.033642f
C461 source.n282 a_n1882_n3288# 0.018078f
C462 source.n283 a_n1882_n3288# 0.042729f
C463 source.n284 a_n1882_n3288# 0.019141f
C464 source.n285 a_n1882_n3288# 0.033642f
C465 source.n286 a_n1882_n3288# 0.018078f
C466 source.n287 a_n1882_n3288# 0.042729f
C467 source.n288 a_n1882_n3288# 0.019141f
C468 source.n289 a_n1882_n3288# 0.033642f
C469 source.n290 a_n1882_n3288# 0.018609f
C470 source.n291 a_n1882_n3288# 0.042729f
C471 source.n292 a_n1882_n3288# 0.019141f
C472 source.n293 a_n1882_n3288# 0.033642f
C473 source.n294 a_n1882_n3288# 0.018078f
C474 source.n295 a_n1882_n3288# 0.042729f
C475 source.n296 a_n1882_n3288# 0.019141f
C476 source.n297 a_n1882_n3288# 0.033642f
C477 source.n298 a_n1882_n3288# 0.018078f
C478 source.n299 a_n1882_n3288# 0.032047f
C479 source.n300 a_n1882_n3288# 0.030206f
C480 source.t16 a_n1882_n3288# 0.072167f
C481 source.n301 a_n1882_n3288# 0.242554f
C482 source.n302 a_n1882_n3288# 1.69718f
C483 source.n303 a_n1882_n3288# 0.018078f
C484 source.n304 a_n1882_n3288# 0.019141f
C485 source.n305 a_n1882_n3288# 0.042729f
C486 source.n306 a_n1882_n3288# 0.042729f
C487 source.n307 a_n1882_n3288# 0.019141f
C488 source.n308 a_n1882_n3288# 0.018078f
C489 source.n309 a_n1882_n3288# 0.033642f
C490 source.n310 a_n1882_n3288# 0.033642f
C491 source.n311 a_n1882_n3288# 0.018078f
C492 source.n312 a_n1882_n3288# 0.019141f
C493 source.n313 a_n1882_n3288# 0.042729f
C494 source.n314 a_n1882_n3288# 0.042729f
C495 source.n315 a_n1882_n3288# 0.019141f
C496 source.n316 a_n1882_n3288# 0.018078f
C497 source.n317 a_n1882_n3288# 0.033642f
C498 source.n318 a_n1882_n3288# 0.033642f
C499 source.n319 a_n1882_n3288# 0.018078f
C500 source.n320 a_n1882_n3288# 0.018078f
C501 source.n321 a_n1882_n3288# 0.019141f
C502 source.n322 a_n1882_n3288# 0.042729f
C503 source.n323 a_n1882_n3288# 0.042729f
C504 source.n324 a_n1882_n3288# 0.042729f
C505 source.n325 a_n1882_n3288# 0.018609f
C506 source.n326 a_n1882_n3288# 0.018078f
C507 source.n327 a_n1882_n3288# 0.033642f
C508 source.n328 a_n1882_n3288# 0.033642f
C509 source.n329 a_n1882_n3288# 0.018078f
C510 source.n330 a_n1882_n3288# 0.019141f
C511 source.n331 a_n1882_n3288# 0.042729f
C512 source.n332 a_n1882_n3288# 0.042729f
C513 source.n333 a_n1882_n3288# 0.019141f
C514 source.n334 a_n1882_n3288# 0.018078f
C515 source.n335 a_n1882_n3288# 0.033642f
C516 source.n336 a_n1882_n3288# 0.033642f
C517 source.n337 a_n1882_n3288# 0.018078f
C518 source.n338 a_n1882_n3288# 0.019141f
C519 source.n339 a_n1882_n3288# 0.042729f
C520 source.n340 a_n1882_n3288# 0.087685f
C521 source.n341 a_n1882_n3288# 0.019141f
C522 source.n342 a_n1882_n3288# 0.018078f
C523 source.n343 a_n1882_n3288# 0.072247f
C524 source.n344 a_n1882_n3288# 0.048392f
C525 source.n345 a_n1882_n3288# 1.86422f
C526 source.t14 a_n1882_n3288# 0.319019f
C527 source.t2 a_n1882_n3288# 0.319019f
C528 source.n346 a_n1882_n3288# 2.73143f
C529 source.n347 a_n1882_n3288# 0.443019f
C530 source.t15 a_n1882_n3288# 0.319019f
C531 source.t17 a_n1882_n3288# 0.319019f
C532 source.n348 a_n1882_n3288# 2.73143f
C533 source.n349 a_n1882_n3288# 0.443019f
C534 source.t6 a_n1882_n3288# 0.319019f
C535 source.t1 a_n1882_n3288# 0.319019f
C536 source.n350 a_n1882_n3288# 2.73143f
C537 source.n351 a_n1882_n3288# 0.443019f
C538 source.t8 a_n1882_n3288# 0.319019f
C539 source.t0 a_n1882_n3288# 0.319019f
C540 source.n352 a_n1882_n3288# 2.73143f
C541 source.n353 a_n1882_n3288# 0.443019f
C542 source.n354 a_n1882_n3288# 0.044563f
C543 source.n355 a_n1882_n3288# 0.033642f
C544 source.n356 a_n1882_n3288# 0.018078f
C545 source.n357 a_n1882_n3288# 0.042729f
C546 source.n358 a_n1882_n3288# 0.019141f
C547 source.n359 a_n1882_n3288# 0.033642f
C548 source.n360 a_n1882_n3288# 0.018078f
C549 source.n361 a_n1882_n3288# 0.042729f
C550 source.n362 a_n1882_n3288# 0.019141f
C551 source.n363 a_n1882_n3288# 0.033642f
C552 source.n364 a_n1882_n3288# 0.018609f
C553 source.n365 a_n1882_n3288# 0.042729f
C554 source.n366 a_n1882_n3288# 0.019141f
C555 source.n367 a_n1882_n3288# 0.033642f
C556 source.n368 a_n1882_n3288# 0.018078f
C557 source.n369 a_n1882_n3288# 0.042729f
C558 source.n370 a_n1882_n3288# 0.019141f
C559 source.n371 a_n1882_n3288# 0.033642f
C560 source.n372 a_n1882_n3288# 0.018078f
C561 source.n373 a_n1882_n3288# 0.032047f
C562 source.n374 a_n1882_n3288# 0.030206f
C563 source.t38 a_n1882_n3288# 0.072167f
C564 source.n375 a_n1882_n3288# 0.242554f
C565 source.n376 a_n1882_n3288# 1.69718f
C566 source.n377 a_n1882_n3288# 0.018078f
C567 source.n378 a_n1882_n3288# 0.019141f
C568 source.n379 a_n1882_n3288# 0.042729f
C569 source.n380 a_n1882_n3288# 0.042729f
C570 source.n381 a_n1882_n3288# 0.019141f
C571 source.n382 a_n1882_n3288# 0.018078f
C572 source.n383 a_n1882_n3288# 0.033642f
C573 source.n384 a_n1882_n3288# 0.033642f
C574 source.n385 a_n1882_n3288# 0.018078f
C575 source.n386 a_n1882_n3288# 0.019141f
C576 source.n387 a_n1882_n3288# 0.042729f
C577 source.n388 a_n1882_n3288# 0.042729f
C578 source.n389 a_n1882_n3288# 0.019141f
C579 source.n390 a_n1882_n3288# 0.018078f
C580 source.n391 a_n1882_n3288# 0.033642f
C581 source.n392 a_n1882_n3288# 0.033642f
C582 source.n393 a_n1882_n3288# 0.018078f
C583 source.n394 a_n1882_n3288# 0.018078f
C584 source.n395 a_n1882_n3288# 0.019141f
C585 source.n396 a_n1882_n3288# 0.042729f
C586 source.n397 a_n1882_n3288# 0.042729f
C587 source.n398 a_n1882_n3288# 0.042729f
C588 source.n399 a_n1882_n3288# 0.018609f
C589 source.n400 a_n1882_n3288# 0.018078f
C590 source.n401 a_n1882_n3288# 0.033642f
C591 source.n402 a_n1882_n3288# 0.033642f
C592 source.n403 a_n1882_n3288# 0.018078f
C593 source.n404 a_n1882_n3288# 0.019141f
C594 source.n405 a_n1882_n3288# 0.042729f
C595 source.n406 a_n1882_n3288# 0.042729f
C596 source.n407 a_n1882_n3288# 0.019141f
C597 source.n408 a_n1882_n3288# 0.018078f
C598 source.n409 a_n1882_n3288# 0.033642f
C599 source.n410 a_n1882_n3288# 0.033642f
C600 source.n411 a_n1882_n3288# 0.018078f
C601 source.n412 a_n1882_n3288# 0.019141f
C602 source.n413 a_n1882_n3288# 0.042729f
C603 source.n414 a_n1882_n3288# 0.087685f
C604 source.n415 a_n1882_n3288# 0.019141f
C605 source.n416 a_n1882_n3288# 0.018078f
C606 source.n417 a_n1882_n3288# 0.072247f
C607 source.n418 a_n1882_n3288# 0.048392f
C608 source.n419 a_n1882_n3288# 0.126085f
C609 source.n420 a_n1882_n3288# 0.044563f
C610 source.n421 a_n1882_n3288# 0.033642f
C611 source.n422 a_n1882_n3288# 0.018078f
C612 source.n423 a_n1882_n3288# 0.042729f
C613 source.n424 a_n1882_n3288# 0.019141f
C614 source.n425 a_n1882_n3288# 0.033642f
C615 source.n426 a_n1882_n3288# 0.018078f
C616 source.n427 a_n1882_n3288# 0.042729f
C617 source.n428 a_n1882_n3288# 0.019141f
C618 source.n429 a_n1882_n3288# 0.033642f
C619 source.n430 a_n1882_n3288# 0.018609f
C620 source.n431 a_n1882_n3288# 0.042729f
C621 source.n432 a_n1882_n3288# 0.019141f
C622 source.n433 a_n1882_n3288# 0.033642f
C623 source.n434 a_n1882_n3288# 0.018078f
C624 source.n435 a_n1882_n3288# 0.042729f
C625 source.n436 a_n1882_n3288# 0.019141f
C626 source.n437 a_n1882_n3288# 0.033642f
C627 source.n438 a_n1882_n3288# 0.018078f
C628 source.n439 a_n1882_n3288# 0.032047f
C629 source.n440 a_n1882_n3288# 0.030206f
C630 source.t26 a_n1882_n3288# 0.072167f
C631 source.n441 a_n1882_n3288# 0.242554f
C632 source.n442 a_n1882_n3288# 1.69718f
C633 source.n443 a_n1882_n3288# 0.018078f
C634 source.n444 a_n1882_n3288# 0.019141f
C635 source.n445 a_n1882_n3288# 0.042729f
C636 source.n446 a_n1882_n3288# 0.042729f
C637 source.n447 a_n1882_n3288# 0.019141f
C638 source.n448 a_n1882_n3288# 0.018078f
C639 source.n449 a_n1882_n3288# 0.033642f
C640 source.n450 a_n1882_n3288# 0.033642f
C641 source.n451 a_n1882_n3288# 0.018078f
C642 source.n452 a_n1882_n3288# 0.019141f
C643 source.n453 a_n1882_n3288# 0.042729f
C644 source.n454 a_n1882_n3288# 0.042729f
C645 source.n455 a_n1882_n3288# 0.019141f
C646 source.n456 a_n1882_n3288# 0.018078f
C647 source.n457 a_n1882_n3288# 0.033642f
C648 source.n458 a_n1882_n3288# 0.033642f
C649 source.n459 a_n1882_n3288# 0.018078f
C650 source.n460 a_n1882_n3288# 0.018078f
C651 source.n461 a_n1882_n3288# 0.019141f
C652 source.n462 a_n1882_n3288# 0.042729f
C653 source.n463 a_n1882_n3288# 0.042729f
C654 source.n464 a_n1882_n3288# 0.042729f
C655 source.n465 a_n1882_n3288# 0.018609f
C656 source.n466 a_n1882_n3288# 0.018078f
C657 source.n467 a_n1882_n3288# 0.033642f
C658 source.n468 a_n1882_n3288# 0.033642f
C659 source.n469 a_n1882_n3288# 0.018078f
C660 source.n470 a_n1882_n3288# 0.019141f
C661 source.n471 a_n1882_n3288# 0.042729f
C662 source.n472 a_n1882_n3288# 0.042729f
C663 source.n473 a_n1882_n3288# 0.019141f
C664 source.n474 a_n1882_n3288# 0.018078f
C665 source.n475 a_n1882_n3288# 0.033642f
C666 source.n476 a_n1882_n3288# 0.033642f
C667 source.n477 a_n1882_n3288# 0.018078f
C668 source.n478 a_n1882_n3288# 0.019141f
C669 source.n479 a_n1882_n3288# 0.042729f
C670 source.n480 a_n1882_n3288# 0.087685f
C671 source.n481 a_n1882_n3288# 0.019141f
C672 source.n482 a_n1882_n3288# 0.018078f
C673 source.n483 a_n1882_n3288# 0.072247f
C674 source.n484 a_n1882_n3288# 0.048392f
C675 source.n485 a_n1882_n3288# 0.126085f
C676 source.t22 a_n1882_n3288# 0.319019f
C677 source.t28 a_n1882_n3288# 0.319019f
C678 source.n486 a_n1882_n3288# 2.73143f
C679 source.n487 a_n1882_n3288# 0.443019f
C680 source.t33 a_n1882_n3288# 0.319019f
C681 source.t32 a_n1882_n3288# 0.319019f
C682 source.n488 a_n1882_n3288# 2.73143f
C683 source.n489 a_n1882_n3288# 0.443019f
C684 source.t20 a_n1882_n3288# 0.319019f
C685 source.t25 a_n1882_n3288# 0.319019f
C686 source.n490 a_n1882_n3288# 2.73143f
C687 source.n491 a_n1882_n3288# 0.443019f
C688 source.t24 a_n1882_n3288# 0.319019f
C689 source.t27 a_n1882_n3288# 0.319019f
C690 source.n492 a_n1882_n3288# 2.73143f
C691 source.n493 a_n1882_n3288# 0.443019f
C692 source.n494 a_n1882_n3288# 0.044563f
C693 source.n495 a_n1882_n3288# 0.033642f
C694 source.n496 a_n1882_n3288# 0.018078f
C695 source.n497 a_n1882_n3288# 0.042729f
C696 source.n498 a_n1882_n3288# 0.019141f
C697 source.n499 a_n1882_n3288# 0.033642f
C698 source.n500 a_n1882_n3288# 0.018078f
C699 source.n501 a_n1882_n3288# 0.042729f
C700 source.n502 a_n1882_n3288# 0.019141f
C701 source.n503 a_n1882_n3288# 0.033642f
C702 source.n504 a_n1882_n3288# 0.018609f
C703 source.n505 a_n1882_n3288# 0.042729f
C704 source.n506 a_n1882_n3288# 0.019141f
C705 source.n507 a_n1882_n3288# 0.033642f
C706 source.n508 a_n1882_n3288# 0.018078f
C707 source.n509 a_n1882_n3288# 0.042729f
C708 source.n510 a_n1882_n3288# 0.019141f
C709 source.n511 a_n1882_n3288# 0.033642f
C710 source.n512 a_n1882_n3288# 0.018078f
C711 source.n513 a_n1882_n3288# 0.032047f
C712 source.n514 a_n1882_n3288# 0.030206f
C713 source.t36 a_n1882_n3288# 0.072167f
C714 source.n515 a_n1882_n3288# 0.242554f
C715 source.n516 a_n1882_n3288# 1.69718f
C716 source.n517 a_n1882_n3288# 0.018078f
C717 source.n518 a_n1882_n3288# 0.019141f
C718 source.n519 a_n1882_n3288# 0.042729f
C719 source.n520 a_n1882_n3288# 0.042729f
C720 source.n521 a_n1882_n3288# 0.019141f
C721 source.n522 a_n1882_n3288# 0.018078f
C722 source.n523 a_n1882_n3288# 0.033642f
C723 source.n524 a_n1882_n3288# 0.033642f
C724 source.n525 a_n1882_n3288# 0.018078f
C725 source.n526 a_n1882_n3288# 0.019141f
C726 source.n527 a_n1882_n3288# 0.042729f
C727 source.n528 a_n1882_n3288# 0.042729f
C728 source.n529 a_n1882_n3288# 0.019141f
C729 source.n530 a_n1882_n3288# 0.018078f
C730 source.n531 a_n1882_n3288# 0.033642f
C731 source.n532 a_n1882_n3288# 0.033642f
C732 source.n533 a_n1882_n3288# 0.018078f
C733 source.n534 a_n1882_n3288# 0.018078f
C734 source.n535 a_n1882_n3288# 0.019141f
C735 source.n536 a_n1882_n3288# 0.042729f
C736 source.n537 a_n1882_n3288# 0.042729f
C737 source.n538 a_n1882_n3288# 0.042729f
C738 source.n539 a_n1882_n3288# 0.018609f
C739 source.n540 a_n1882_n3288# 0.018078f
C740 source.n541 a_n1882_n3288# 0.033642f
C741 source.n542 a_n1882_n3288# 0.033642f
C742 source.n543 a_n1882_n3288# 0.018078f
C743 source.n544 a_n1882_n3288# 0.019141f
C744 source.n545 a_n1882_n3288# 0.042729f
C745 source.n546 a_n1882_n3288# 0.042729f
C746 source.n547 a_n1882_n3288# 0.019141f
C747 source.n548 a_n1882_n3288# 0.018078f
C748 source.n549 a_n1882_n3288# 0.033642f
C749 source.n550 a_n1882_n3288# 0.033642f
C750 source.n551 a_n1882_n3288# 0.018078f
C751 source.n552 a_n1882_n3288# 0.019141f
C752 source.n553 a_n1882_n3288# 0.042729f
C753 source.n554 a_n1882_n3288# 0.087685f
C754 source.n555 a_n1882_n3288# 0.019141f
C755 source.n556 a_n1882_n3288# 0.018078f
C756 source.n557 a_n1882_n3288# 0.072247f
C757 source.n558 a_n1882_n3288# 0.048392f
C758 source.n559 a_n1882_n3288# 0.308502f
C759 source.n560 a_n1882_n3288# 2.10528f
C760 minus.n0 a_n1882_n3288# 0.052649f
C761 minus.t12 a_n1882_n3288# 0.362145f
C762 minus.t15 a_n1882_n3288# 0.357067f
C763 minus.t19 a_n1882_n3288# 0.357067f
C764 minus.t1 a_n1882_n3288# 0.357067f
C765 minus.n1 a_n1882_n3288# 0.147056f
C766 minus.n2 a_n1882_n3288# 0.052649f
C767 minus.t9 a_n1882_n3288# 0.357067f
C768 minus.t17 a_n1882_n3288# 0.357067f
C769 minus.t18 a_n1882_n3288# 0.357067f
C770 minus.n3 a_n1882_n3288# 0.147056f
C771 minus.n4 a_n1882_n3288# 0.120476f
C772 minus.t0 a_n1882_n3288# 0.357067f
C773 minus.t10 a_n1882_n3288# 0.357067f
C774 minus.t16 a_n1882_n3288# 0.362145f
C775 minus.n5 a_n1882_n3288# 0.163256f
C776 minus.n6 a_n1882_n3288# 0.147056f
C777 minus.n7 a_n1882_n3288# 0.018439f
C778 minus.n8 a_n1882_n3288# 0.147056f
C779 minus.n9 a_n1882_n3288# 0.018439f
C780 minus.n10 a_n1882_n3288# 0.052649f
C781 minus.n11 a_n1882_n3288# 0.052649f
C782 minus.n12 a_n1882_n3288# 0.018439f
C783 minus.n13 a_n1882_n3288# 0.147056f
C784 minus.n14 a_n1882_n3288# 0.018439f
C785 minus.n15 a_n1882_n3288# 0.147056f
C786 minus.n16 a_n1882_n3288# 0.018439f
C787 minus.n17 a_n1882_n3288# 0.052649f
C788 minus.n18 a_n1882_n3288# 0.052649f
C789 minus.n19 a_n1882_n3288# 0.018439f
C790 minus.n20 a_n1882_n3288# 0.147056f
C791 minus.n21 a_n1882_n3288# 0.018439f
C792 minus.n22 a_n1882_n3288# 0.147056f
C793 minus.n23 a_n1882_n3288# 0.163176f
C794 minus.n24 a_n1882_n3288# 1.86252f
C795 minus.n25 a_n1882_n3288# 0.052649f
C796 minus.t11 a_n1882_n3288# 0.357067f
C797 minus.t7 a_n1882_n3288# 0.357067f
C798 minus.t13 a_n1882_n3288# 0.357067f
C799 minus.n26 a_n1882_n3288# 0.147056f
C800 minus.n27 a_n1882_n3288# 0.052649f
C801 minus.t8 a_n1882_n3288# 0.357067f
C802 minus.t14 a_n1882_n3288# 0.357067f
C803 minus.t5 a_n1882_n3288# 0.357067f
C804 minus.n28 a_n1882_n3288# 0.147056f
C805 minus.n29 a_n1882_n3288# 0.120476f
C806 minus.t2 a_n1882_n3288# 0.357067f
C807 minus.t6 a_n1882_n3288# 0.357067f
C808 minus.t3 a_n1882_n3288# 0.362145f
C809 minus.n30 a_n1882_n3288# 0.163256f
C810 minus.n31 a_n1882_n3288# 0.147056f
C811 minus.n32 a_n1882_n3288# 0.018439f
C812 minus.n33 a_n1882_n3288# 0.147056f
C813 minus.n34 a_n1882_n3288# 0.018439f
C814 minus.n35 a_n1882_n3288# 0.052649f
C815 minus.n36 a_n1882_n3288# 0.052649f
C816 minus.n37 a_n1882_n3288# 0.018439f
C817 minus.n38 a_n1882_n3288# 0.147056f
C818 minus.n39 a_n1882_n3288# 0.018439f
C819 minus.n40 a_n1882_n3288# 0.147056f
C820 minus.n41 a_n1882_n3288# 0.018439f
C821 minus.n42 a_n1882_n3288# 0.052649f
C822 minus.n43 a_n1882_n3288# 0.052649f
C823 minus.n44 a_n1882_n3288# 0.018439f
C824 minus.n45 a_n1882_n3288# 0.147056f
C825 minus.n46 a_n1882_n3288# 0.018439f
C826 minus.n47 a_n1882_n3288# 0.147056f
C827 minus.t4 a_n1882_n3288# 0.362145f
C828 minus.n48 a_n1882_n3288# 0.163176f
C829 minus.n49 a_n1882_n3288# 0.341448f
C830 minus.n50 a_n1882_n3288# 2.26315f
.ends

