* NGSPICE file created from diffpair457.ext - technology: sky130A

.subckt diffpair457 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t17 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X1 drain_left.t15 plus.t0 source.t9 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X2 source.t27 minus.t1 drain_right.t14 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X3 drain_right.t13 minus.t2 source.t16 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X4 drain_left.t14 plus.t1 source.t6 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X5 source.t14 plus.t2 drain_left.t13 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X6 source.t15 plus.t3 drain_left.t12 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X7 drain_left.t11 plus.t4 source.t3 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X8 source.t26 minus.t3 drain_right.t12 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X9 a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.6
X10 drain_right.t11 minus.t4 source.t28 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X11 drain_right.t10 minus.t5 source.t24 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X12 source.t29 minus.t6 drain_right.t9 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X13 a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X14 source.t22 minus.t7 drain_right.t8 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X15 source.t10 plus.t5 drain_left.t10 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X16 source.t4 plus.t6 drain_left.t9 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X17 source.t31 minus.t8 drain_right.t7 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X18 source.t21 minus.t9 drain_right.t6 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X19 drain_right.t5 minus.t10 source.t20 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X20 source.t25 minus.t11 drain_right.t4 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X21 a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X22 drain_left.t8 plus.t7 source.t8 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X23 source.t23 minus.t12 drain_right.t3 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X24 source.t11 plus.t8 drain_left.t7 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X25 drain_right.t2 minus.t13 source.t19 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X26 drain_left.t6 plus.t9 source.t0 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X27 drain_left.t5 plus.t10 source.t12 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X28 drain_left.t4 plus.t11 source.t1 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X29 source.t7 plus.t12 drain_left.t3 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X30 a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X31 drain_right.t1 minus.t14 source.t18 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X32 drain_right.t0 minus.t15 source.t30 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X33 drain_left.t2 plus.t13 source.t2 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X34 source.t13 plus.t14 drain_left.t1 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X35 source.t5 plus.t15 drain_left.t0 a_n2390_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
R0 minus.n6 minus.t13 568.453
R1 minus.n30 minus.t11 568.453
R2 minus.n5 minus.t12 547.472
R3 minus.n9 minus.t10 547.472
R4 minus.n3 minus.t8 547.472
R5 minus.n15 minus.t4 547.472
R6 minus.n1 minus.t6 547.472
R7 minus.n21 minus.t5 547.472
R8 minus.n22 minus.t3 547.472
R9 minus.n29 minus.t2 547.472
R10 minus.n33 minus.t7 547.472
R11 minus.n27 minus.t15 547.472
R12 minus.n39 minus.t1 547.472
R13 minus.n25 minus.t0 547.472
R14 minus.n45 minus.t9 547.472
R15 minus.n46 minus.t14 547.472
R16 minus.n23 minus.n22 161.3
R17 minus.n21 minus.n0 161.3
R18 minus.n20 minus.n19 161.3
R19 minus.n18 minus.n1 161.3
R20 minus.n17 minus.n16 161.3
R21 minus.n15 minus.n2 161.3
R22 minus.n14 minus.n13 161.3
R23 minus.n12 minus.n3 161.3
R24 minus.n11 minus.n10 161.3
R25 minus.n9 minus.n4 161.3
R26 minus.n8 minus.n7 161.3
R27 minus.n47 minus.n46 161.3
R28 minus.n45 minus.n24 161.3
R29 minus.n44 minus.n43 161.3
R30 minus.n42 minus.n25 161.3
R31 minus.n41 minus.n40 161.3
R32 minus.n39 minus.n26 161.3
R33 minus.n38 minus.n37 161.3
R34 minus.n36 minus.n27 161.3
R35 minus.n35 minus.n34 161.3
R36 minus.n33 minus.n28 161.3
R37 minus.n32 minus.n31 161.3
R38 minus.n7 minus.n6 70.4033
R39 minus.n31 minus.n30 70.4033
R40 minus.n22 minus.n21 48.2005
R41 minus.n46 minus.n45 48.2005
R42 minus.n9 minus.n8 44.549
R43 minus.n20 minus.n1 44.549
R44 minus.n33 minus.n32 44.549
R45 minus.n44 minus.n25 44.549
R46 minus.n48 minus.n23 38.33
R47 minus.n10 minus.n3 34.3247
R48 minus.n16 minus.n15 34.3247
R49 minus.n34 minus.n27 34.3247
R50 minus.n40 minus.n39 34.3247
R51 minus.n15 minus.n14 24.1005
R52 minus.n14 minus.n3 24.1005
R53 minus.n38 minus.n27 24.1005
R54 minus.n39 minus.n38 24.1005
R55 minus.n6 minus.n5 20.9576
R56 minus.n30 minus.n29 20.9576
R57 minus.n10 minus.n9 13.8763
R58 minus.n16 minus.n1 13.8763
R59 minus.n34 minus.n33 13.8763
R60 minus.n40 minus.n25 13.8763
R61 minus.n48 minus.n47 6.6558
R62 minus.n8 minus.n5 3.65202
R63 minus.n21 minus.n20 3.65202
R64 minus.n32 minus.n29 3.65202
R65 minus.n45 minus.n44 3.65202
R66 minus.n23 minus.n0 0.189894
R67 minus.n19 minus.n0 0.189894
R68 minus.n19 minus.n18 0.189894
R69 minus.n18 minus.n17 0.189894
R70 minus.n17 minus.n2 0.189894
R71 minus.n13 minus.n2 0.189894
R72 minus.n13 minus.n12 0.189894
R73 minus.n12 minus.n11 0.189894
R74 minus.n11 minus.n4 0.189894
R75 minus.n7 minus.n4 0.189894
R76 minus.n31 minus.n28 0.189894
R77 minus.n35 minus.n28 0.189894
R78 minus.n36 minus.n35 0.189894
R79 minus.n37 minus.n36 0.189894
R80 minus.n37 minus.n26 0.189894
R81 minus.n41 minus.n26 0.189894
R82 minus.n42 minus.n41 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n24 0.189894
R85 minus.n47 minus.n24 0.189894
R86 minus minus.n48 0.188
R87 source.n546 source.n486 289.615
R88 source.n474 source.n414 289.615
R89 source.n408 source.n348 289.615
R90 source.n336 source.n276 289.615
R91 source.n60 source.n0 289.615
R92 source.n132 source.n72 289.615
R93 source.n198 source.n138 289.615
R94 source.n270 source.n210 289.615
R95 source.n506 source.n505 185
R96 source.n511 source.n510 185
R97 source.n513 source.n512 185
R98 source.n502 source.n501 185
R99 source.n519 source.n518 185
R100 source.n521 source.n520 185
R101 source.n498 source.n497 185
R102 source.n528 source.n527 185
R103 source.n529 source.n496 185
R104 source.n531 source.n530 185
R105 source.n494 source.n493 185
R106 source.n537 source.n536 185
R107 source.n539 source.n538 185
R108 source.n490 source.n489 185
R109 source.n545 source.n544 185
R110 source.n547 source.n546 185
R111 source.n434 source.n433 185
R112 source.n439 source.n438 185
R113 source.n441 source.n440 185
R114 source.n430 source.n429 185
R115 source.n447 source.n446 185
R116 source.n449 source.n448 185
R117 source.n426 source.n425 185
R118 source.n456 source.n455 185
R119 source.n457 source.n424 185
R120 source.n459 source.n458 185
R121 source.n422 source.n421 185
R122 source.n465 source.n464 185
R123 source.n467 source.n466 185
R124 source.n418 source.n417 185
R125 source.n473 source.n472 185
R126 source.n475 source.n474 185
R127 source.n368 source.n367 185
R128 source.n373 source.n372 185
R129 source.n375 source.n374 185
R130 source.n364 source.n363 185
R131 source.n381 source.n380 185
R132 source.n383 source.n382 185
R133 source.n360 source.n359 185
R134 source.n390 source.n389 185
R135 source.n391 source.n358 185
R136 source.n393 source.n392 185
R137 source.n356 source.n355 185
R138 source.n399 source.n398 185
R139 source.n401 source.n400 185
R140 source.n352 source.n351 185
R141 source.n407 source.n406 185
R142 source.n409 source.n408 185
R143 source.n296 source.n295 185
R144 source.n301 source.n300 185
R145 source.n303 source.n302 185
R146 source.n292 source.n291 185
R147 source.n309 source.n308 185
R148 source.n311 source.n310 185
R149 source.n288 source.n287 185
R150 source.n318 source.n317 185
R151 source.n319 source.n286 185
R152 source.n321 source.n320 185
R153 source.n284 source.n283 185
R154 source.n327 source.n326 185
R155 source.n329 source.n328 185
R156 source.n280 source.n279 185
R157 source.n335 source.n334 185
R158 source.n337 source.n336 185
R159 source.n61 source.n60 185
R160 source.n59 source.n58 185
R161 source.n4 source.n3 185
R162 source.n53 source.n52 185
R163 source.n51 source.n50 185
R164 source.n8 source.n7 185
R165 source.n45 source.n44 185
R166 source.n43 source.n10 185
R167 source.n42 source.n41 185
R168 source.n13 source.n11 185
R169 source.n36 source.n35 185
R170 source.n34 source.n33 185
R171 source.n17 source.n16 185
R172 source.n28 source.n27 185
R173 source.n26 source.n25 185
R174 source.n21 source.n20 185
R175 source.n133 source.n132 185
R176 source.n131 source.n130 185
R177 source.n76 source.n75 185
R178 source.n125 source.n124 185
R179 source.n123 source.n122 185
R180 source.n80 source.n79 185
R181 source.n117 source.n116 185
R182 source.n115 source.n82 185
R183 source.n114 source.n113 185
R184 source.n85 source.n83 185
R185 source.n108 source.n107 185
R186 source.n106 source.n105 185
R187 source.n89 source.n88 185
R188 source.n100 source.n99 185
R189 source.n98 source.n97 185
R190 source.n93 source.n92 185
R191 source.n199 source.n198 185
R192 source.n197 source.n196 185
R193 source.n142 source.n141 185
R194 source.n191 source.n190 185
R195 source.n189 source.n188 185
R196 source.n146 source.n145 185
R197 source.n183 source.n182 185
R198 source.n181 source.n148 185
R199 source.n180 source.n179 185
R200 source.n151 source.n149 185
R201 source.n174 source.n173 185
R202 source.n172 source.n171 185
R203 source.n155 source.n154 185
R204 source.n166 source.n165 185
R205 source.n164 source.n163 185
R206 source.n159 source.n158 185
R207 source.n271 source.n270 185
R208 source.n269 source.n268 185
R209 source.n214 source.n213 185
R210 source.n263 source.n262 185
R211 source.n261 source.n260 185
R212 source.n218 source.n217 185
R213 source.n255 source.n254 185
R214 source.n253 source.n220 185
R215 source.n252 source.n251 185
R216 source.n223 source.n221 185
R217 source.n246 source.n245 185
R218 source.n244 source.n243 185
R219 source.n227 source.n226 185
R220 source.n238 source.n237 185
R221 source.n236 source.n235 185
R222 source.n231 source.n230 185
R223 source.n507 source.t18 149.524
R224 source.n435 source.t25 149.524
R225 source.n369 source.t2 149.524
R226 source.n297 source.t5 149.524
R227 source.n22 source.t6 149.524
R228 source.n94 source.t7 149.524
R229 source.n160 source.t19 149.524
R230 source.n232 source.t26 149.524
R231 source.n511 source.n505 104.615
R232 source.n512 source.n511 104.615
R233 source.n512 source.n501 104.615
R234 source.n519 source.n501 104.615
R235 source.n520 source.n519 104.615
R236 source.n520 source.n497 104.615
R237 source.n528 source.n497 104.615
R238 source.n529 source.n528 104.615
R239 source.n530 source.n529 104.615
R240 source.n530 source.n493 104.615
R241 source.n537 source.n493 104.615
R242 source.n538 source.n537 104.615
R243 source.n538 source.n489 104.615
R244 source.n545 source.n489 104.615
R245 source.n546 source.n545 104.615
R246 source.n439 source.n433 104.615
R247 source.n440 source.n439 104.615
R248 source.n440 source.n429 104.615
R249 source.n447 source.n429 104.615
R250 source.n448 source.n447 104.615
R251 source.n448 source.n425 104.615
R252 source.n456 source.n425 104.615
R253 source.n457 source.n456 104.615
R254 source.n458 source.n457 104.615
R255 source.n458 source.n421 104.615
R256 source.n465 source.n421 104.615
R257 source.n466 source.n465 104.615
R258 source.n466 source.n417 104.615
R259 source.n473 source.n417 104.615
R260 source.n474 source.n473 104.615
R261 source.n373 source.n367 104.615
R262 source.n374 source.n373 104.615
R263 source.n374 source.n363 104.615
R264 source.n381 source.n363 104.615
R265 source.n382 source.n381 104.615
R266 source.n382 source.n359 104.615
R267 source.n390 source.n359 104.615
R268 source.n391 source.n390 104.615
R269 source.n392 source.n391 104.615
R270 source.n392 source.n355 104.615
R271 source.n399 source.n355 104.615
R272 source.n400 source.n399 104.615
R273 source.n400 source.n351 104.615
R274 source.n407 source.n351 104.615
R275 source.n408 source.n407 104.615
R276 source.n301 source.n295 104.615
R277 source.n302 source.n301 104.615
R278 source.n302 source.n291 104.615
R279 source.n309 source.n291 104.615
R280 source.n310 source.n309 104.615
R281 source.n310 source.n287 104.615
R282 source.n318 source.n287 104.615
R283 source.n319 source.n318 104.615
R284 source.n320 source.n319 104.615
R285 source.n320 source.n283 104.615
R286 source.n327 source.n283 104.615
R287 source.n328 source.n327 104.615
R288 source.n328 source.n279 104.615
R289 source.n335 source.n279 104.615
R290 source.n336 source.n335 104.615
R291 source.n60 source.n59 104.615
R292 source.n59 source.n3 104.615
R293 source.n52 source.n3 104.615
R294 source.n52 source.n51 104.615
R295 source.n51 source.n7 104.615
R296 source.n44 source.n7 104.615
R297 source.n44 source.n43 104.615
R298 source.n43 source.n42 104.615
R299 source.n42 source.n11 104.615
R300 source.n35 source.n11 104.615
R301 source.n35 source.n34 104.615
R302 source.n34 source.n16 104.615
R303 source.n27 source.n16 104.615
R304 source.n27 source.n26 104.615
R305 source.n26 source.n20 104.615
R306 source.n132 source.n131 104.615
R307 source.n131 source.n75 104.615
R308 source.n124 source.n75 104.615
R309 source.n124 source.n123 104.615
R310 source.n123 source.n79 104.615
R311 source.n116 source.n79 104.615
R312 source.n116 source.n115 104.615
R313 source.n115 source.n114 104.615
R314 source.n114 source.n83 104.615
R315 source.n107 source.n83 104.615
R316 source.n107 source.n106 104.615
R317 source.n106 source.n88 104.615
R318 source.n99 source.n88 104.615
R319 source.n99 source.n98 104.615
R320 source.n98 source.n92 104.615
R321 source.n198 source.n197 104.615
R322 source.n197 source.n141 104.615
R323 source.n190 source.n141 104.615
R324 source.n190 source.n189 104.615
R325 source.n189 source.n145 104.615
R326 source.n182 source.n145 104.615
R327 source.n182 source.n181 104.615
R328 source.n181 source.n180 104.615
R329 source.n180 source.n149 104.615
R330 source.n173 source.n149 104.615
R331 source.n173 source.n172 104.615
R332 source.n172 source.n154 104.615
R333 source.n165 source.n154 104.615
R334 source.n165 source.n164 104.615
R335 source.n164 source.n158 104.615
R336 source.n270 source.n269 104.615
R337 source.n269 source.n213 104.615
R338 source.n262 source.n213 104.615
R339 source.n262 source.n261 104.615
R340 source.n261 source.n217 104.615
R341 source.n254 source.n217 104.615
R342 source.n254 source.n253 104.615
R343 source.n253 source.n252 104.615
R344 source.n252 source.n221 104.615
R345 source.n245 source.n221 104.615
R346 source.n245 source.n244 104.615
R347 source.n244 source.n226 104.615
R348 source.n237 source.n226 104.615
R349 source.n237 source.n236 104.615
R350 source.n236 source.n230 104.615
R351 source.t18 source.n505 52.3082
R352 source.t25 source.n433 52.3082
R353 source.t2 source.n367 52.3082
R354 source.t5 source.n295 52.3082
R355 source.t6 source.n20 52.3082
R356 source.t7 source.n92 52.3082
R357 source.t19 source.n158 52.3082
R358 source.t26 source.n230 52.3082
R359 source.n67 source.n66 42.8739
R360 source.n69 source.n68 42.8739
R361 source.n71 source.n70 42.8739
R362 source.n205 source.n204 42.8739
R363 source.n207 source.n206 42.8739
R364 source.n209 source.n208 42.8739
R365 source.n485 source.n484 42.8737
R366 source.n483 source.n482 42.8737
R367 source.n481 source.n480 42.8737
R368 source.n347 source.n346 42.8737
R369 source.n345 source.n344 42.8737
R370 source.n343 source.n342 42.8737
R371 source.n551 source.n550 29.8581
R372 source.n479 source.n478 29.8581
R373 source.n413 source.n412 29.8581
R374 source.n341 source.n340 29.8581
R375 source.n65 source.n64 29.8581
R376 source.n137 source.n136 29.8581
R377 source.n203 source.n202 29.8581
R378 source.n275 source.n274 29.8581
R379 source.n341 source.n275 22.0894
R380 source.n552 source.n65 16.4257
R381 source.n531 source.n496 13.1884
R382 source.n459 source.n424 13.1884
R383 source.n393 source.n358 13.1884
R384 source.n321 source.n286 13.1884
R385 source.n45 source.n10 13.1884
R386 source.n117 source.n82 13.1884
R387 source.n183 source.n148 13.1884
R388 source.n255 source.n220 13.1884
R389 source.n527 source.n526 12.8005
R390 source.n532 source.n494 12.8005
R391 source.n455 source.n454 12.8005
R392 source.n460 source.n422 12.8005
R393 source.n389 source.n388 12.8005
R394 source.n394 source.n356 12.8005
R395 source.n317 source.n316 12.8005
R396 source.n322 source.n284 12.8005
R397 source.n46 source.n8 12.8005
R398 source.n41 source.n12 12.8005
R399 source.n118 source.n80 12.8005
R400 source.n113 source.n84 12.8005
R401 source.n184 source.n146 12.8005
R402 source.n179 source.n150 12.8005
R403 source.n256 source.n218 12.8005
R404 source.n251 source.n222 12.8005
R405 source.n525 source.n498 12.0247
R406 source.n536 source.n535 12.0247
R407 source.n453 source.n426 12.0247
R408 source.n464 source.n463 12.0247
R409 source.n387 source.n360 12.0247
R410 source.n398 source.n397 12.0247
R411 source.n315 source.n288 12.0247
R412 source.n326 source.n325 12.0247
R413 source.n50 source.n49 12.0247
R414 source.n40 source.n13 12.0247
R415 source.n122 source.n121 12.0247
R416 source.n112 source.n85 12.0247
R417 source.n188 source.n187 12.0247
R418 source.n178 source.n151 12.0247
R419 source.n260 source.n259 12.0247
R420 source.n250 source.n223 12.0247
R421 source.n522 source.n521 11.249
R422 source.n539 source.n492 11.249
R423 source.n450 source.n449 11.249
R424 source.n467 source.n420 11.249
R425 source.n384 source.n383 11.249
R426 source.n401 source.n354 11.249
R427 source.n312 source.n311 11.249
R428 source.n329 source.n282 11.249
R429 source.n53 source.n6 11.249
R430 source.n37 source.n36 11.249
R431 source.n125 source.n78 11.249
R432 source.n109 source.n108 11.249
R433 source.n191 source.n144 11.249
R434 source.n175 source.n174 11.249
R435 source.n263 source.n216 11.249
R436 source.n247 source.n246 11.249
R437 source.n518 source.n500 10.4732
R438 source.n540 source.n490 10.4732
R439 source.n446 source.n428 10.4732
R440 source.n468 source.n418 10.4732
R441 source.n380 source.n362 10.4732
R442 source.n402 source.n352 10.4732
R443 source.n308 source.n290 10.4732
R444 source.n330 source.n280 10.4732
R445 source.n54 source.n4 10.4732
R446 source.n33 source.n15 10.4732
R447 source.n126 source.n76 10.4732
R448 source.n105 source.n87 10.4732
R449 source.n192 source.n142 10.4732
R450 source.n171 source.n153 10.4732
R451 source.n264 source.n214 10.4732
R452 source.n243 source.n225 10.4732
R453 source.n507 source.n506 10.2747
R454 source.n435 source.n434 10.2747
R455 source.n369 source.n368 10.2747
R456 source.n297 source.n296 10.2747
R457 source.n22 source.n21 10.2747
R458 source.n94 source.n93 10.2747
R459 source.n160 source.n159 10.2747
R460 source.n232 source.n231 10.2747
R461 source.n517 source.n502 9.69747
R462 source.n544 source.n543 9.69747
R463 source.n445 source.n430 9.69747
R464 source.n472 source.n471 9.69747
R465 source.n379 source.n364 9.69747
R466 source.n406 source.n405 9.69747
R467 source.n307 source.n292 9.69747
R468 source.n334 source.n333 9.69747
R469 source.n58 source.n57 9.69747
R470 source.n32 source.n17 9.69747
R471 source.n130 source.n129 9.69747
R472 source.n104 source.n89 9.69747
R473 source.n196 source.n195 9.69747
R474 source.n170 source.n155 9.69747
R475 source.n268 source.n267 9.69747
R476 source.n242 source.n227 9.69747
R477 source.n550 source.n549 9.45567
R478 source.n478 source.n477 9.45567
R479 source.n412 source.n411 9.45567
R480 source.n340 source.n339 9.45567
R481 source.n64 source.n63 9.45567
R482 source.n136 source.n135 9.45567
R483 source.n202 source.n201 9.45567
R484 source.n274 source.n273 9.45567
R485 source.n549 source.n548 9.3005
R486 source.n488 source.n487 9.3005
R487 source.n543 source.n542 9.3005
R488 source.n541 source.n540 9.3005
R489 source.n492 source.n491 9.3005
R490 source.n535 source.n534 9.3005
R491 source.n533 source.n532 9.3005
R492 source.n509 source.n508 9.3005
R493 source.n504 source.n503 9.3005
R494 source.n515 source.n514 9.3005
R495 source.n517 source.n516 9.3005
R496 source.n500 source.n499 9.3005
R497 source.n523 source.n522 9.3005
R498 source.n525 source.n524 9.3005
R499 source.n526 source.n495 9.3005
R500 source.n477 source.n476 9.3005
R501 source.n416 source.n415 9.3005
R502 source.n471 source.n470 9.3005
R503 source.n469 source.n468 9.3005
R504 source.n420 source.n419 9.3005
R505 source.n463 source.n462 9.3005
R506 source.n461 source.n460 9.3005
R507 source.n437 source.n436 9.3005
R508 source.n432 source.n431 9.3005
R509 source.n443 source.n442 9.3005
R510 source.n445 source.n444 9.3005
R511 source.n428 source.n427 9.3005
R512 source.n451 source.n450 9.3005
R513 source.n453 source.n452 9.3005
R514 source.n454 source.n423 9.3005
R515 source.n411 source.n410 9.3005
R516 source.n350 source.n349 9.3005
R517 source.n405 source.n404 9.3005
R518 source.n403 source.n402 9.3005
R519 source.n354 source.n353 9.3005
R520 source.n397 source.n396 9.3005
R521 source.n395 source.n394 9.3005
R522 source.n371 source.n370 9.3005
R523 source.n366 source.n365 9.3005
R524 source.n377 source.n376 9.3005
R525 source.n379 source.n378 9.3005
R526 source.n362 source.n361 9.3005
R527 source.n385 source.n384 9.3005
R528 source.n387 source.n386 9.3005
R529 source.n388 source.n357 9.3005
R530 source.n339 source.n338 9.3005
R531 source.n278 source.n277 9.3005
R532 source.n333 source.n332 9.3005
R533 source.n331 source.n330 9.3005
R534 source.n282 source.n281 9.3005
R535 source.n325 source.n324 9.3005
R536 source.n323 source.n322 9.3005
R537 source.n299 source.n298 9.3005
R538 source.n294 source.n293 9.3005
R539 source.n305 source.n304 9.3005
R540 source.n307 source.n306 9.3005
R541 source.n290 source.n289 9.3005
R542 source.n313 source.n312 9.3005
R543 source.n315 source.n314 9.3005
R544 source.n316 source.n285 9.3005
R545 source.n24 source.n23 9.3005
R546 source.n19 source.n18 9.3005
R547 source.n30 source.n29 9.3005
R548 source.n32 source.n31 9.3005
R549 source.n15 source.n14 9.3005
R550 source.n38 source.n37 9.3005
R551 source.n40 source.n39 9.3005
R552 source.n12 source.n9 9.3005
R553 source.n63 source.n62 9.3005
R554 source.n2 source.n1 9.3005
R555 source.n57 source.n56 9.3005
R556 source.n55 source.n54 9.3005
R557 source.n6 source.n5 9.3005
R558 source.n49 source.n48 9.3005
R559 source.n47 source.n46 9.3005
R560 source.n96 source.n95 9.3005
R561 source.n91 source.n90 9.3005
R562 source.n102 source.n101 9.3005
R563 source.n104 source.n103 9.3005
R564 source.n87 source.n86 9.3005
R565 source.n110 source.n109 9.3005
R566 source.n112 source.n111 9.3005
R567 source.n84 source.n81 9.3005
R568 source.n135 source.n134 9.3005
R569 source.n74 source.n73 9.3005
R570 source.n129 source.n128 9.3005
R571 source.n127 source.n126 9.3005
R572 source.n78 source.n77 9.3005
R573 source.n121 source.n120 9.3005
R574 source.n119 source.n118 9.3005
R575 source.n162 source.n161 9.3005
R576 source.n157 source.n156 9.3005
R577 source.n168 source.n167 9.3005
R578 source.n170 source.n169 9.3005
R579 source.n153 source.n152 9.3005
R580 source.n176 source.n175 9.3005
R581 source.n178 source.n177 9.3005
R582 source.n150 source.n147 9.3005
R583 source.n201 source.n200 9.3005
R584 source.n140 source.n139 9.3005
R585 source.n195 source.n194 9.3005
R586 source.n193 source.n192 9.3005
R587 source.n144 source.n143 9.3005
R588 source.n187 source.n186 9.3005
R589 source.n185 source.n184 9.3005
R590 source.n234 source.n233 9.3005
R591 source.n229 source.n228 9.3005
R592 source.n240 source.n239 9.3005
R593 source.n242 source.n241 9.3005
R594 source.n225 source.n224 9.3005
R595 source.n248 source.n247 9.3005
R596 source.n250 source.n249 9.3005
R597 source.n222 source.n219 9.3005
R598 source.n273 source.n272 9.3005
R599 source.n212 source.n211 9.3005
R600 source.n267 source.n266 9.3005
R601 source.n265 source.n264 9.3005
R602 source.n216 source.n215 9.3005
R603 source.n259 source.n258 9.3005
R604 source.n257 source.n256 9.3005
R605 source.n514 source.n513 8.92171
R606 source.n547 source.n488 8.92171
R607 source.n442 source.n441 8.92171
R608 source.n475 source.n416 8.92171
R609 source.n376 source.n375 8.92171
R610 source.n409 source.n350 8.92171
R611 source.n304 source.n303 8.92171
R612 source.n337 source.n278 8.92171
R613 source.n61 source.n2 8.92171
R614 source.n29 source.n28 8.92171
R615 source.n133 source.n74 8.92171
R616 source.n101 source.n100 8.92171
R617 source.n199 source.n140 8.92171
R618 source.n167 source.n166 8.92171
R619 source.n271 source.n212 8.92171
R620 source.n239 source.n238 8.92171
R621 source.n510 source.n504 8.14595
R622 source.n548 source.n486 8.14595
R623 source.n438 source.n432 8.14595
R624 source.n476 source.n414 8.14595
R625 source.n372 source.n366 8.14595
R626 source.n410 source.n348 8.14595
R627 source.n300 source.n294 8.14595
R628 source.n338 source.n276 8.14595
R629 source.n62 source.n0 8.14595
R630 source.n25 source.n19 8.14595
R631 source.n134 source.n72 8.14595
R632 source.n97 source.n91 8.14595
R633 source.n200 source.n138 8.14595
R634 source.n163 source.n157 8.14595
R635 source.n272 source.n210 8.14595
R636 source.n235 source.n229 8.14595
R637 source.n509 source.n506 7.3702
R638 source.n437 source.n434 7.3702
R639 source.n371 source.n368 7.3702
R640 source.n299 source.n296 7.3702
R641 source.n24 source.n21 7.3702
R642 source.n96 source.n93 7.3702
R643 source.n162 source.n159 7.3702
R644 source.n234 source.n231 7.3702
R645 source.n510 source.n509 5.81868
R646 source.n550 source.n486 5.81868
R647 source.n438 source.n437 5.81868
R648 source.n478 source.n414 5.81868
R649 source.n372 source.n371 5.81868
R650 source.n412 source.n348 5.81868
R651 source.n300 source.n299 5.81868
R652 source.n340 source.n276 5.81868
R653 source.n64 source.n0 5.81868
R654 source.n25 source.n24 5.81868
R655 source.n136 source.n72 5.81868
R656 source.n97 source.n96 5.81868
R657 source.n202 source.n138 5.81868
R658 source.n163 source.n162 5.81868
R659 source.n274 source.n210 5.81868
R660 source.n235 source.n234 5.81868
R661 source.n552 source.n551 5.66429
R662 source.n513 source.n504 5.04292
R663 source.n548 source.n547 5.04292
R664 source.n441 source.n432 5.04292
R665 source.n476 source.n475 5.04292
R666 source.n375 source.n366 5.04292
R667 source.n410 source.n409 5.04292
R668 source.n303 source.n294 5.04292
R669 source.n338 source.n337 5.04292
R670 source.n62 source.n61 5.04292
R671 source.n28 source.n19 5.04292
R672 source.n134 source.n133 5.04292
R673 source.n100 source.n91 5.04292
R674 source.n200 source.n199 5.04292
R675 source.n166 source.n157 5.04292
R676 source.n272 source.n271 5.04292
R677 source.n238 source.n229 5.04292
R678 source.n514 source.n502 4.26717
R679 source.n544 source.n488 4.26717
R680 source.n442 source.n430 4.26717
R681 source.n472 source.n416 4.26717
R682 source.n376 source.n364 4.26717
R683 source.n406 source.n350 4.26717
R684 source.n304 source.n292 4.26717
R685 source.n334 source.n278 4.26717
R686 source.n58 source.n2 4.26717
R687 source.n29 source.n17 4.26717
R688 source.n130 source.n74 4.26717
R689 source.n101 source.n89 4.26717
R690 source.n196 source.n140 4.26717
R691 source.n167 source.n155 4.26717
R692 source.n268 source.n212 4.26717
R693 source.n239 source.n227 4.26717
R694 source.n518 source.n517 3.49141
R695 source.n543 source.n490 3.49141
R696 source.n446 source.n445 3.49141
R697 source.n471 source.n418 3.49141
R698 source.n380 source.n379 3.49141
R699 source.n405 source.n352 3.49141
R700 source.n308 source.n307 3.49141
R701 source.n333 source.n280 3.49141
R702 source.n57 source.n4 3.49141
R703 source.n33 source.n32 3.49141
R704 source.n129 source.n76 3.49141
R705 source.n105 source.n104 3.49141
R706 source.n195 source.n142 3.49141
R707 source.n171 source.n170 3.49141
R708 source.n267 source.n214 3.49141
R709 source.n243 source.n242 3.49141
R710 source.n508 source.n507 2.84303
R711 source.n436 source.n435 2.84303
R712 source.n370 source.n369 2.84303
R713 source.n298 source.n297 2.84303
R714 source.n23 source.n22 2.84303
R715 source.n95 source.n94 2.84303
R716 source.n161 source.n160 2.84303
R717 source.n233 source.n232 2.84303
R718 source.n521 source.n500 2.71565
R719 source.n540 source.n539 2.71565
R720 source.n449 source.n428 2.71565
R721 source.n468 source.n467 2.71565
R722 source.n383 source.n362 2.71565
R723 source.n402 source.n401 2.71565
R724 source.n311 source.n290 2.71565
R725 source.n330 source.n329 2.71565
R726 source.n54 source.n53 2.71565
R727 source.n36 source.n15 2.71565
R728 source.n126 source.n125 2.71565
R729 source.n108 source.n87 2.71565
R730 source.n192 source.n191 2.71565
R731 source.n174 source.n153 2.71565
R732 source.n264 source.n263 2.71565
R733 source.n246 source.n225 2.71565
R734 source.n522 source.n498 1.93989
R735 source.n536 source.n492 1.93989
R736 source.n450 source.n426 1.93989
R737 source.n464 source.n420 1.93989
R738 source.n384 source.n360 1.93989
R739 source.n398 source.n354 1.93989
R740 source.n312 source.n288 1.93989
R741 source.n326 source.n282 1.93989
R742 source.n50 source.n6 1.93989
R743 source.n37 source.n13 1.93989
R744 source.n122 source.n78 1.93989
R745 source.n109 source.n85 1.93989
R746 source.n188 source.n144 1.93989
R747 source.n175 source.n151 1.93989
R748 source.n260 source.n216 1.93989
R749 source.n247 source.n223 1.93989
R750 source.n484 source.t17 1.6505
R751 source.n484 source.t21 1.6505
R752 source.n482 source.t30 1.6505
R753 source.n482 source.t27 1.6505
R754 source.n480 source.t16 1.6505
R755 source.n480 source.t22 1.6505
R756 source.n346 source.t0 1.6505
R757 source.n346 source.t10 1.6505
R758 source.n344 source.t9 1.6505
R759 source.n344 source.t13 1.6505
R760 source.n342 source.t12 1.6505
R761 source.n342 source.t15 1.6505
R762 source.n66 source.t3 1.6505
R763 source.n66 source.t14 1.6505
R764 source.n68 source.t8 1.6505
R765 source.n68 source.t4 1.6505
R766 source.n70 source.t1 1.6505
R767 source.n70 source.t11 1.6505
R768 source.n204 source.t20 1.6505
R769 source.n204 source.t23 1.6505
R770 source.n206 source.t28 1.6505
R771 source.n206 source.t31 1.6505
R772 source.n208 source.t24 1.6505
R773 source.n208 source.t29 1.6505
R774 source.n527 source.n525 1.16414
R775 source.n535 source.n494 1.16414
R776 source.n455 source.n453 1.16414
R777 source.n463 source.n422 1.16414
R778 source.n389 source.n387 1.16414
R779 source.n397 source.n356 1.16414
R780 source.n317 source.n315 1.16414
R781 source.n325 source.n284 1.16414
R782 source.n49 source.n8 1.16414
R783 source.n41 source.n40 1.16414
R784 source.n121 source.n80 1.16414
R785 source.n113 source.n112 1.16414
R786 source.n187 source.n146 1.16414
R787 source.n179 source.n178 1.16414
R788 source.n259 source.n218 1.16414
R789 source.n251 source.n250 1.16414
R790 source.n275 source.n209 0.802224
R791 source.n209 source.n207 0.802224
R792 source.n207 source.n205 0.802224
R793 source.n205 source.n203 0.802224
R794 source.n137 source.n71 0.802224
R795 source.n71 source.n69 0.802224
R796 source.n69 source.n67 0.802224
R797 source.n67 source.n65 0.802224
R798 source.n343 source.n341 0.802224
R799 source.n345 source.n343 0.802224
R800 source.n347 source.n345 0.802224
R801 source.n413 source.n347 0.802224
R802 source.n481 source.n479 0.802224
R803 source.n483 source.n481 0.802224
R804 source.n485 source.n483 0.802224
R805 source.n551 source.n485 0.802224
R806 source.n203 source.n137 0.470328
R807 source.n479 source.n413 0.470328
R808 source.n526 source.n496 0.388379
R809 source.n532 source.n531 0.388379
R810 source.n454 source.n424 0.388379
R811 source.n460 source.n459 0.388379
R812 source.n388 source.n358 0.388379
R813 source.n394 source.n393 0.388379
R814 source.n316 source.n286 0.388379
R815 source.n322 source.n321 0.388379
R816 source.n46 source.n45 0.388379
R817 source.n12 source.n10 0.388379
R818 source.n118 source.n117 0.388379
R819 source.n84 source.n82 0.388379
R820 source.n184 source.n183 0.388379
R821 source.n150 source.n148 0.388379
R822 source.n256 source.n255 0.388379
R823 source.n222 source.n220 0.388379
R824 source source.n552 0.188
R825 source.n508 source.n503 0.155672
R826 source.n515 source.n503 0.155672
R827 source.n516 source.n515 0.155672
R828 source.n516 source.n499 0.155672
R829 source.n523 source.n499 0.155672
R830 source.n524 source.n523 0.155672
R831 source.n524 source.n495 0.155672
R832 source.n533 source.n495 0.155672
R833 source.n534 source.n533 0.155672
R834 source.n534 source.n491 0.155672
R835 source.n541 source.n491 0.155672
R836 source.n542 source.n541 0.155672
R837 source.n542 source.n487 0.155672
R838 source.n549 source.n487 0.155672
R839 source.n436 source.n431 0.155672
R840 source.n443 source.n431 0.155672
R841 source.n444 source.n443 0.155672
R842 source.n444 source.n427 0.155672
R843 source.n451 source.n427 0.155672
R844 source.n452 source.n451 0.155672
R845 source.n452 source.n423 0.155672
R846 source.n461 source.n423 0.155672
R847 source.n462 source.n461 0.155672
R848 source.n462 source.n419 0.155672
R849 source.n469 source.n419 0.155672
R850 source.n470 source.n469 0.155672
R851 source.n470 source.n415 0.155672
R852 source.n477 source.n415 0.155672
R853 source.n370 source.n365 0.155672
R854 source.n377 source.n365 0.155672
R855 source.n378 source.n377 0.155672
R856 source.n378 source.n361 0.155672
R857 source.n385 source.n361 0.155672
R858 source.n386 source.n385 0.155672
R859 source.n386 source.n357 0.155672
R860 source.n395 source.n357 0.155672
R861 source.n396 source.n395 0.155672
R862 source.n396 source.n353 0.155672
R863 source.n403 source.n353 0.155672
R864 source.n404 source.n403 0.155672
R865 source.n404 source.n349 0.155672
R866 source.n411 source.n349 0.155672
R867 source.n298 source.n293 0.155672
R868 source.n305 source.n293 0.155672
R869 source.n306 source.n305 0.155672
R870 source.n306 source.n289 0.155672
R871 source.n313 source.n289 0.155672
R872 source.n314 source.n313 0.155672
R873 source.n314 source.n285 0.155672
R874 source.n323 source.n285 0.155672
R875 source.n324 source.n323 0.155672
R876 source.n324 source.n281 0.155672
R877 source.n331 source.n281 0.155672
R878 source.n332 source.n331 0.155672
R879 source.n332 source.n277 0.155672
R880 source.n339 source.n277 0.155672
R881 source.n63 source.n1 0.155672
R882 source.n56 source.n1 0.155672
R883 source.n56 source.n55 0.155672
R884 source.n55 source.n5 0.155672
R885 source.n48 source.n5 0.155672
R886 source.n48 source.n47 0.155672
R887 source.n47 source.n9 0.155672
R888 source.n39 source.n9 0.155672
R889 source.n39 source.n38 0.155672
R890 source.n38 source.n14 0.155672
R891 source.n31 source.n14 0.155672
R892 source.n31 source.n30 0.155672
R893 source.n30 source.n18 0.155672
R894 source.n23 source.n18 0.155672
R895 source.n135 source.n73 0.155672
R896 source.n128 source.n73 0.155672
R897 source.n128 source.n127 0.155672
R898 source.n127 source.n77 0.155672
R899 source.n120 source.n77 0.155672
R900 source.n120 source.n119 0.155672
R901 source.n119 source.n81 0.155672
R902 source.n111 source.n81 0.155672
R903 source.n111 source.n110 0.155672
R904 source.n110 source.n86 0.155672
R905 source.n103 source.n86 0.155672
R906 source.n103 source.n102 0.155672
R907 source.n102 source.n90 0.155672
R908 source.n95 source.n90 0.155672
R909 source.n201 source.n139 0.155672
R910 source.n194 source.n139 0.155672
R911 source.n194 source.n193 0.155672
R912 source.n193 source.n143 0.155672
R913 source.n186 source.n143 0.155672
R914 source.n186 source.n185 0.155672
R915 source.n185 source.n147 0.155672
R916 source.n177 source.n147 0.155672
R917 source.n177 source.n176 0.155672
R918 source.n176 source.n152 0.155672
R919 source.n169 source.n152 0.155672
R920 source.n169 source.n168 0.155672
R921 source.n168 source.n156 0.155672
R922 source.n161 source.n156 0.155672
R923 source.n273 source.n211 0.155672
R924 source.n266 source.n211 0.155672
R925 source.n266 source.n265 0.155672
R926 source.n265 source.n215 0.155672
R927 source.n258 source.n215 0.155672
R928 source.n258 source.n257 0.155672
R929 source.n257 source.n219 0.155672
R930 source.n249 source.n219 0.155672
R931 source.n249 source.n248 0.155672
R932 source.n248 source.n224 0.155672
R933 source.n241 source.n224 0.155672
R934 source.n241 source.n240 0.155672
R935 source.n240 source.n228 0.155672
R936 source.n233 source.n228 0.155672
R937 drain_right.n5 drain_right.n3 60.3542
R938 drain_right.n2 drain_right.n0 60.3542
R939 drain_right.n9 drain_right.n7 60.3542
R940 drain_right.n9 drain_right.n8 59.5527
R941 drain_right.n11 drain_right.n10 59.5527
R942 drain_right.n13 drain_right.n12 59.5527
R943 drain_right.n5 drain_right.n4 59.5525
R944 drain_right.n2 drain_right.n1 59.5525
R945 drain_right drain_right.n6 32.0251
R946 drain_right drain_right.n13 6.45494
R947 drain_right.n3 drain_right.t6 1.6505
R948 drain_right.n3 drain_right.t1 1.6505
R949 drain_right.n4 drain_right.t14 1.6505
R950 drain_right.n4 drain_right.t15 1.6505
R951 drain_right.n1 drain_right.t8 1.6505
R952 drain_right.n1 drain_right.t0 1.6505
R953 drain_right.n0 drain_right.t4 1.6505
R954 drain_right.n0 drain_right.t13 1.6505
R955 drain_right.n7 drain_right.t3 1.6505
R956 drain_right.n7 drain_right.t2 1.6505
R957 drain_right.n8 drain_right.t7 1.6505
R958 drain_right.n8 drain_right.t5 1.6505
R959 drain_right.n10 drain_right.t9 1.6505
R960 drain_right.n10 drain_right.t11 1.6505
R961 drain_right.n12 drain_right.t12 1.6505
R962 drain_right.n12 drain_right.t10 1.6505
R963 drain_right.n13 drain_right.n11 0.802224
R964 drain_right.n11 drain_right.n9 0.802224
R965 drain_right.n6 drain_right.n5 0.346016
R966 drain_right.n6 drain_right.n2 0.346016
R967 plus.n6 plus.t12 568.453
R968 plus.n30 plus.t13 568.453
R969 plus.n22 plus.t1 547.472
R970 plus.n21 plus.t2 547.472
R971 plus.n1 plus.t4 547.472
R972 plus.n15 plus.t6 547.472
R973 plus.n3 plus.t7 547.472
R974 plus.n9 plus.t8 547.472
R975 plus.n5 plus.t11 547.472
R976 plus.n46 plus.t15 547.472
R977 plus.n45 plus.t10 547.472
R978 plus.n25 plus.t3 547.472
R979 plus.n39 plus.t0 547.472
R980 plus.n27 plus.t14 547.472
R981 plus.n33 plus.t9 547.472
R982 plus.n29 plus.t5 547.472
R983 plus.n8 plus.n7 161.3
R984 plus.n9 plus.n4 161.3
R985 plus.n11 plus.n10 161.3
R986 plus.n12 plus.n3 161.3
R987 plus.n14 plus.n13 161.3
R988 plus.n15 plus.n2 161.3
R989 plus.n17 plus.n16 161.3
R990 plus.n18 plus.n1 161.3
R991 plus.n20 plus.n19 161.3
R992 plus.n21 plus.n0 161.3
R993 plus.n23 plus.n22 161.3
R994 plus.n32 plus.n31 161.3
R995 plus.n33 plus.n28 161.3
R996 plus.n35 plus.n34 161.3
R997 plus.n36 plus.n27 161.3
R998 plus.n38 plus.n37 161.3
R999 plus.n39 plus.n26 161.3
R1000 plus.n41 plus.n40 161.3
R1001 plus.n42 plus.n25 161.3
R1002 plus.n44 plus.n43 161.3
R1003 plus.n45 plus.n24 161.3
R1004 plus.n47 plus.n46 161.3
R1005 plus.n7 plus.n6 70.4033
R1006 plus.n31 plus.n30 70.4033
R1007 plus.n22 plus.n21 48.2005
R1008 plus.n46 plus.n45 48.2005
R1009 plus.n20 plus.n1 44.549
R1010 plus.n9 plus.n8 44.549
R1011 plus.n44 plus.n25 44.549
R1012 plus.n33 plus.n32 44.549
R1013 plus.n16 plus.n15 34.3247
R1014 plus.n10 plus.n3 34.3247
R1015 plus.n40 plus.n39 34.3247
R1016 plus.n34 plus.n27 34.3247
R1017 plus plus.n47 32.2111
R1018 plus.n14 plus.n3 24.1005
R1019 plus.n15 plus.n14 24.1005
R1020 plus.n39 plus.n38 24.1005
R1021 plus.n38 plus.n27 24.1005
R1022 plus.n6 plus.n5 20.9576
R1023 plus.n30 plus.n29 20.9576
R1024 plus.n16 plus.n1 13.8763
R1025 plus.n10 plus.n9 13.8763
R1026 plus.n40 plus.n25 13.8763
R1027 plus.n34 plus.n33 13.8763
R1028 plus plus.n23 12.2997
R1029 plus.n21 plus.n20 3.65202
R1030 plus.n8 plus.n5 3.65202
R1031 plus.n45 plus.n44 3.65202
R1032 plus.n32 plus.n29 3.65202
R1033 plus.n7 plus.n4 0.189894
R1034 plus.n11 plus.n4 0.189894
R1035 plus.n12 plus.n11 0.189894
R1036 plus.n13 plus.n12 0.189894
R1037 plus.n13 plus.n2 0.189894
R1038 plus.n17 plus.n2 0.189894
R1039 plus.n18 plus.n17 0.189894
R1040 plus.n19 plus.n18 0.189894
R1041 plus.n19 plus.n0 0.189894
R1042 plus.n23 plus.n0 0.189894
R1043 plus.n47 plus.n24 0.189894
R1044 plus.n43 plus.n24 0.189894
R1045 plus.n43 plus.n42 0.189894
R1046 plus.n42 plus.n41 0.189894
R1047 plus.n41 plus.n26 0.189894
R1048 plus.n37 plus.n26 0.189894
R1049 plus.n37 plus.n36 0.189894
R1050 plus.n36 plus.n35 0.189894
R1051 plus.n35 plus.n28 0.189894
R1052 plus.n31 plus.n28 0.189894
R1053 drain_left.n9 drain_left.n7 60.3544
R1054 drain_left.n5 drain_left.n3 60.3542
R1055 drain_left.n2 drain_left.n0 60.3542
R1056 drain_left.n11 drain_left.n10 59.5527
R1057 drain_left.n9 drain_left.n8 59.5527
R1058 drain_left.n5 drain_left.n4 59.5525
R1059 drain_left.n2 drain_left.n1 59.5525
R1060 drain_left.n13 drain_left.n12 59.5525
R1061 drain_left drain_left.n6 32.5783
R1062 drain_left drain_left.n13 6.45494
R1063 drain_left.n3 drain_left.t10 1.6505
R1064 drain_left.n3 drain_left.t2 1.6505
R1065 drain_left.n4 drain_left.t1 1.6505
R1066 drain_left.n4 drain_left.t6 1.6505
R1067 drain_left.n1 drain_left.t12 1.6505
R1068 drain_left.n1 drain_left.t15 1.6505
R1069 drain_left.n0 drain_left.t0 1.6505
R1070 drain_left.n0 drain_left.t5 1.6505
R1071 drain_left.n12 drain_left.t13 1.6505
R1072 drain_left.n12 drain_left.t14 1.6505
R1073 drain_left.n10 drain_left.t9 1.6505
R1074 drain_left.n10 drain_left.t11 1.6505
R1075 drain_left.n8 drain_left.t7 1.6505
R1076 drain_left.n8 drain_left.t8 1.6505
R1077 drain_left.n7 drain_left.t3 1.6505
R1078 drain_left.n7 drain_left.t4 1.6505
R1079 drain_left.n11 drain_left.n9 0.802224
R1080 drain_left.n13 drain_left.n11 0.802224
R1081 drain_left.n6 drain_left.n5 0.346016
R1082 drain_left.n6 drain_left.n2 0.346016
C0 minus source 9.31807f
C1 drain_right source 21.41f
C2 plus source 9.33211f
C3 drain_left source 21.4083f
C4 drain_right minus 9.35956f
C5 minus plus 6.12424f
C6 drain_right plus 0.391974f
C7 minus drain_left 0.172752f
C8 drain_right drain_left 1.24373f
C9 drain_left plus 9.595469f
C10 drain_right a_n2390_n3288# 6.6733f
C11 drain_left a_n2390_n3288# 7.01416f
C12 source a_n2390_n3288# 9.14929f
C13 minus a_n2390_n3288# 9.483788f
C14 plus a_n2390_n3288# 11.29196f
C15 drain_left.t0 a_n2390_n3288# 0.266708f
C16 drain_left.t5 a_n2390_n3288# 0.266708f
C17 drain_left.n0 a_n2390_n3288# 2.37851f
C18 drain_left.t12 a_n2390_n3288# 0.266708f
C19 drain_left.t15 a_n2390_n3288# 0.266708f
C20 drain_left.n1 a_n2390_n3288# 2.37329f
C21 drain_left.n2 a_n2390_n3288# 0.729376f
C22 drain_left.t10 a_n2390_n3288# 0.266708f
C23 drain_left.t2 a_n2390_n3288# 0.266708f
C24 drain_left.n3 a_n2390_n3288# 2.37851f
C25 drain_left.t1 a_n2390_n3288# 0.266708f
C26 drain_left.t6 a_n2390_n3288# 0.266708f
C27 drain_left.n4 a_n2390_n3288# 2.37329f
C28 drain_left.n5 a_n2390_n3288# 0.729376f
C29 drain_left.n6 a_n2390_n3288# 1.55626f
C30 drain_left.t3 a_n2390_n3288# 0.266708f
C31 drain_left.t4 a_n2390_n3288# 0.266708f
C32 drain_left.n7 a_n2390_n3288# 2.37852f
C33 drain_left.t7 a_n2390_n3288# 0.266708f
C34 drain_left.t8 a_n2390_n3288# 0.266708f
C35 drain_left.n8 a_n2390_n3288# 2.3733f
C36 drain_left.n9 a_n2390_n3288# 0.768814f
C37 drain_left.t9 a_n2390_n3288# 0.266708f
C38 drain_left.t11 a_n2390_n3288# 0.266708f
C39 drain_left.n10 a_n2390_n3288# 2.3733f
C40 drain_left.n11 a_n2390_n3288# 0.381351f
C41 drain_left.t13 a_n2390_n3288# 0.266708f
C42 drain_left.t14 a_n2390_n3288# 0.266708f
C43 drain_left.n12 a_n2390_n3288# 2.37329f
C44 drain_left.n13 a_n2390_n3288# 0.626614f
C45 plus.n0 a_n2390_n3288# 0.043207f
C46 plus.t1 a_n2390_n3288# 0.88708f
C47 plus.t2 a_n2390_n3288# 0.88708f
C48 plus.t4 a_n2390_n3288# 0.88708f
C49 plus.n1 a_n2390_n3288# 0.357735f
C50 plus.n2 a_n2390_n3288# 0.043207f
C51 plus.t6 a_n2390_n3288# 0.88708f
C52 plus.t7 a_n2390_n3288# 0.88708f
C53 plus.n3 a_n2390_n3288# 0.357735f
C54 plus.n4 a_n2390_n3288# 0.043207f
C55 plus.t8 a_n2390_n3288# 0.88708f
C56 plus.t11 a_n2390_n3288# 0.88708f
C57 plus.n5 a_n2390_n3288# 0.356536f
C58 plus.t12 a_n2390_n3288# 0.900218f
C59 plus.n6 a_n2390_n3288# 0.343078f
C60 plus.n7 a_n2390_n3288# 0.145525f
C61 plus.n8 a_n2390_n3288# 0.009805f
C62 plus.n9 a_n2390_n3288# 0.357735f
C63 plus.n10 a_n2390_n3288# 0.009805f
C64 plus.n11 a_n2390_n3288# 0.043207f
C65 plus.n12 a_n2390_n3288# 0.043207f
C66 plus.n13 a_n2390_n3288# 0.043207f
C67 plus.n14 a_n2390_n3288# 0.009805f
C68 plus.n15 a_n2390_n3288# 0.357735f
C69 plus.n16 a_n2390_n3288# 0.009805f
C70 plus.n17 a_n2390_n3288# 0.043207f
C71 plus.n18 a_n2390_n3288# 0.043207f
C72 plus.n19 a_n2390_n3288# 0.043207f
C73 plus.n20 a_n2390_n3288# 0.009805f
C74 plus.n21 a_n2390_n3288# 0.356536f
C75 plus.n22 a_n2390_n3288# 0.35587f
C76 plus.n23 a_n2390_n3288# 0.499452f
C77 plus.n24 a_n2390_n3288# 0.043207f
C78 plus.t15 a_n2390_n3288# 0.88708f
C79 plus.t10 a_n2390_n3288# 0.88708f
C80 plus.t3 a_n2390_n3288# 0.88708f
C81 plus.n25 a_n2390_n3288# 0.357735f
C82 plus.n26 a_n2390_n3288# 0.043207f
C83 plus.t0 a_n2390_n3288# 0.88708f
C84 plus.t14 a_n2390_n3288# 0.88708f
C85 plus.n27 a_n2390_n3288# 0.357735f
C86 plus.n28 a_n2390_n3288# 0.043207f
C87 plus.t9 a_n2390_n3288# 0.88708f
C88 plus.t5 a_n2390_n3288# 0.88708f
C89 plus.n29 a_n2390_n3288# 0.356536f
C90 plus.t13 a_n2390_n3288# 0.900218f
C91 plus.n30 a_n2390_n3288# 0.343078f
C92 plus.n31 a_n2390_n3288# 0.145525f
C93 plus.n32 a_n2390_n3288# 0.009805f
C94 plus.n33 a_n2390_n3288# 0.357735f
C95 plus.n34 a_n2390_n3288# 0.009805f
C96 plus.n35 a_n2390_n3288# 0.043207f
C97 plus.n36 a_n2390_n3288# 0.043207f
C98 plus.n37 a_n2390_n3288# 0.043207f
C99 plus.n38 a_n2390_n3288# 0.009805f
C100 plus.n39 a_n2390_n3288# 0.357735f
C101 plus.n40 a_n2390_n3288# 0.009805f
C102 plus.n41 a_n2390_n3288# 0.043207f
C103 plus.n42 a_n2390_n3288# 0.043207f
C104 plus.n43 a_n2390_n3288# 0.043207f
C105 plus.n44 a_n2390_n3288# 0.009805f
C106 plus.n45 a_n2390_n3288# 0.356536f
C107 plus.n46 a_n2390_n3288# 0.35587f
C108 plus.n47 a_n2390_n3288# 1.42409f
C109 drain_right.t4 a_n2390_n3288# 0.265931f
C110 drain_right.t13 a_n2390_n3288# 0.265931f
C111 drain_right.n0 a_n2390_n3288# 2.37158f
C112 drain_right.t8 a_n2390_n3288# 0.265931f
C113 drain_right.t0 a_n2390_n3288# 0.265931f
C114 drain_right.n1 a_n2390_n3288# 2.36638f
C115 drain_right.n2 a_n2390_n3288# 0.727252f
C116 drain_right.t6 a_n2390_n3288# 0.265931f
C117 drain_right.t1 a_n2390_n3288# 0.265931f
C118 drain_right.n3 a_n2390_n3288# 2.37158f
C119 drain_right.t14 a_n2390_n3288# 0.265931f
C120 drain_right.t15 a_n2390_n3288# 0.265931f
C121 drain_right.n4 a_n2390_n3288# 2.36638f
C122 drain_right.n5 a_n2390_n3288# 0.727252f
C123 drain_right.n6 a_n2390_n3288# 1.49409f
C124 drain_right.t3 a_n2390_n3288# 0.265931f
C125 drain_right.t2 a_n2390_n3288# 0.265931f
C126 drain_right.n7 a_n2390_n3288# 2.37158f
C127 drain_right.t7 a_n2390_n3288# 0.265931f
C128 drain_right.t5 a_n2390_n3288# 0.265931f
C129 drain_right.n8 a_n2390_n3288# 2.36639f
C130 drain_right.n9 a_n2390_n3288# 0.766585f
C131 drain_right.t9 a_n2390_n3288# 0.265931f
C132 drain_right.t11 a_n2390_n3288# 0.265931f
C133 drain_right.n10 a_n2390_n3288# 2.36639f
C134 drain_right.n11 a_n2390_n3288# 0.38024f
C135 drain_right.t12 a_n2390_n3288# 0.265931f
C136 drain_right.t10 a_n2390_n3288# 0.265931f
C137 drain_right.n12 a_n2390_n3288# 2.36639f
C138 drain_right.n13 a_n2390_n3288# 0.624779f
C139 source.n0 a_n2390_n3288# 0.031634f
C140 source.n1 a_n2390_n3288# 0.023881f
C141 source.n2 a_n2390_n3288# 0.012833f
C142 source.n3 a_n2390_n3288# 0.030332f
C143 source.n4 a_n2390_n3288# 0.013587f
C144 source.n5 a_n2390_n3288# 0.023881f
C145 source.n6 a_n2390_n3288# 0.012833f
C146 source.n7 a_n2390_n3288# 0.030332f
C147 source.n8 a_n2390_n3288# 0.013587f
C148 source.n9 a_n2390_n3288# 0.023881f
C149 source.n10 a_n2390_n3288# 0.01321f
C150 source.n11 a_n2390_n3288# 0.030332f
C151 source.n12 a_n2390_n3288# 0.012833f
C152 source.n13 a_n2390_n3288# 0.013587f
C153 source.n14 a_n2390_n3288# 0.023881f
C154 source.n15 a_n2390_n3288# 0.012833f
C155 source.n16 a_n2390_n3288# 0.030332f
C156 source.n17 a_n2390_n3288# 0.013587f
C157 source.n18 a_n2390_n3288# 0.023881f
C158 source.n19 a_n2390_n3288# 0.012833f
C159 source.n20 a_n2390_n3288# 0.022749f
C160 source.n21 a_n2390_n3288# 0.021442f
C161 source.t6 a_n2390_n3288# 0.051228f
C162 source.n22 a_n2390_n3288# 0.17218f
C163 source.n23 a_n2390_n3288# 1.20476f
C164 source.n24 a_n2390_n3288# 0.012833f
C165 source.n25 a_n2390_n3288# 0.013587f
C166 source.n26 a_n2390_n3288# 0.030332f
C167 source.n27 a_n2390_n3288# 0.030332f
C168 source.n28 a_n2390_n3288# 0.013587f
C169 source.n29 a_n2390_n3288# 0.012833f
C170 source.n30 a_n2390_n3288# 0.023881f
C171 source.n31 a_n2390_n3288# 0.023881f
C172 source.n32 a_n2390_n3288# 0.012833f
C173 source.n33 a_n2390_n3288# 0.013587f
C174 source.n34 a_n2390_n3288# 0.030332f
C175 source.n35 a_n2390_n3288# 0.030332f
C176 source.n36 a_n2390_n3288# 0.013587f
C177 source.n37 a_n2390_n3288# 0.012833f
C178 source.n38 a_n2390_n3288# 0.023881f
C179 source.n39 a_n2390_n3288# 0.023881f
C180 source.n40 a_n2390_n3288# 0.012833f
C181 source.n41 a_n2390_n3288# 0.013587f
C182 source.n42 a_n2390_n3288# 0.030332f
C183 source.n43 a_n2390_n3288# 0.030332f
C184 source.n44 a_n2390_n3288# 0.030332f
C185 source.n45 a_n2390_n3288# 0.01321f
C186 source.n46 a_n2390_n3288# 0.012833f
C187 source.n47 a_n2390_n3288# 0.023881f
C188 source.n48 a_n2390_n3288# 0.023881f
C189 source.n49 a_n2390_n3288# 0.012833f
C190 source.n50 a_n2390_n3288# 0.013587f
C191 source.n51 a_n2390_n3288# 0.030332f
C192 source.n52 a_n2390_n3288# 0.030332f
C193 source.n53 a_n2390_n3288# 0.013587f
C194 source.n54 a_n2390_n3288# 0.012833f
C195 source.n55 a_n2390_n3288# 0.023881f
C196 source.n56 a_n2390_n3288# 0.023881f
C197 source.n57 a_n2390_n3288# 0.012833f
C198 source.n58 a_n2390_n3288# 0.013587f
C199 source.n59 a_n2390_n3288# 0.030332f
C200 source.n60 a_n2390_n3288# 0.062244f
C201 source.n61 a_n2390_n3288# 0.013587f
C202 source.n62 a_n2390_n3288# 0.012833f
C203 source.n63 a_n2390_n3288# 0.051285f
C204 source.n64 a_n2390_n3288# 0.034352f
C205 source.n65 a_n2390_n3288# 0.993725f
C206 source.t3 a_n2390_n3288# 0.226459f
C207 source.t14 a_n2390_n3288# 0.226459f
C208 source.n66 a_n2390_n3288# 1.93895f
C209 source.n67 a_n2390_n3288# 0.36754f
C210 source.t8 a_n2390_n3288# 0.226459f
C211 source.t4 a_n2390_n3288# 0.226459f
C212 source.n68 a_n2390_n3288# 1.93895f
C213 source.n69 a_n2390_n3288# 0.36754f
C214 source.t1 a_n2390_n3288# 0.226459f
C215 source.t11 a_n2390_n3288# 0.226459f
C216 source.n70 a_n2390_n3288# 1.93895f
C217 source.n71 a_n2390_n3288# 0.36754f
C218 source.n72 a_n2390_n3288# 0.031634f
C219 source.n73 a_n2390_n3288# 0.023881f
C220 source.n74 a_n2390_n3288# 0.012833f
C221 source.n75 a_n2390_n3288# 0.030332f
C222 source.n76 a_n2390_n3288# 0.013587f
C223 source.n77 a_n2390_n3288# 0.023881f
C224 source.n78 a_n2390_n3288# 0.012833f
C225 source.n79 a_n2390_n3288# 0.030332f
C226 source.n80 a_n2390_n3288# 0.013587f
C227 source.n81 a_n2390_n3288# 0.023881f
C228 source.n82 a_n2390_n3288# 0.01321f
C229 source.n83 a_n2390_n3288# 0.030332f
C230 source.n84 a_n2390_n3288# 0.012833f
C231 source.n85 a_n2390_n3288# 0.013587f
C232 source.n86 a_n2390_n3288# 0.023881f
C233 source.n87 a_n2390_n3288# 0.012833f
C234 source.n88 a_n2390_n3288# 0.030332f
C235 source.n89 a_n2390_n3288# 0.013587f
C236 source.n90 a_n2390_n3288# 0.023881f
C237 source.n91 a_n2390_n3288# 0.012833f
C238 source.n92 a_n2390_n3288# 0.022749f
C239 source.n93 a_n2390_n3288# 0.021442f
C240 source.t7 a_n2390_n3288# 0.051228f
C241 source.n94 a_n2390_n3288# 0.17218f
C242 source.n95 a_n2390_n3288# 1.20476f
C243 source.n96 a_n2390_n3288# 0.012833f
C244 source.n97 a_n2390_n3288# 0.013587f
C245 source.n98 a_n2390_n3288# 0.030332f
C246 source.n99 a_n2390_n3288# 0.030332f
C247 source.n100 a_n2390_n3288# 0.013587f
C248 source.n101 a_n2390_n3288# 0.012833f
C249 source.n102 a_n2390_n3288# 0.023881f
C250 source.n103 a_n2390_n3288# 0.023881f
C251 source.n104 a_n2390_n3288# 0.012833f
C252 source.n105 a_n2390_n3288# 0.013587f
C253 source.n106 a_n2390_n3288# 0.030332f
C254 source.n107 a_n2390_n3288# 0.030332f
C255 source.n108 a_n2390_n3288# 0.013587f
C256 source.n109 a_n2390_n3288# 0.012833f
C257 source.n110 a_n2390_n3288# 0.023881f
C258 source.n111 a_n2390_n3288# 0.023881f
C259 source.n112 a_n2390_n3288# 0.012833f
C260 source.n113 a_n2390_n3288# 0.013587f
C261 source.n114 a_n2390_n3288# 0.030332f
C262 source.n115 a_n2390_n3288# 0.030332f
C263 source.n116 a_n2390_n3288# 0.030332f
C264 source.n117 a_n2390_n3288# 0.01321f
C265 source.n118 a_n2390_n3288# 0.012833f
C266 source.n119 a_n2390_n3288# 0.023881f
C267 source.n120 a_n2390_n3288# 0.023881f
C268 source.n121 a_n2390_n3288# 0.012833f
C269 source.n122 a_n2390_n3288# 0.013587f
C270 source.n123 a_n2390_n3288# 0.030332f
C271 source.n124 a_n2390_n3288# 0.030332f
C272 source.n125 a_n2390_n3288# 0.013587f
C273 source.n126 a_n2390_n3288# 0.012833f
C274 source.n127 a_n2390_n3288# 0.023881f
C275 source.n128 a_n2390_n3288# 0.023881f
C276 source.n129 a_n2390_n3288# 0.012833f
C277 source.n130 a_n2390_n3288# 0.013587f
C278 source.n131 a_n2390_n3288# 0.030332f
C279 source.n132 a_n2390_n3288# 0.062244f
C280 source.n133 a_n2390_n3288# 0.013587f
C281 source.n134 a_n2390_n3288# 0.012833f
C282 source.n135 a_n2390_n3288# 0.051285f
C283 source.n136 a_n2390_n3288# 0.034352f
C284 source.n137 a_n2390_n3288# 0.116037f
C285 source.n138 a_n2390_n3288# 0.031634f
C286 source.n139 a_n2390_n3288# 0.023881f
C287 source.n140 a_n2390_n3288# 0.012833f
C288 source.n141 a_n2390_n3288# 0.030332f
C289 source.n142 a_n2390_n3288# 0.013587f
C290 source.n143 a_n2390_n3288# 0.023881f
C291 source.n144 a_n2390_n3288# 0.012833f
C292 source.n145 a_n2390_n3288# 0.030332f
C293 source.n146 a_n2390_n3288# 0.013587f
C294 source.n147 a_n2390_n3288# 0.023881f
C295 source.n148 a_n2390_n3288# 0.01321f
C296 source.n149 a_n2390_n3288# 0.030332f
C297 source.n150 a_n2390_n3288# 0.012833f
C298 source.n151 a_n2390_n3288# 0.013587f
C299 source.n152 a_n2390_n3288# 0.023881f
C300 source.n153 a_n2390_n3288# 0.012833f
C301 source.n154 a_n2390_n3288# 0.030332f
C302 source.n155 a_n2390_n3288# 0.013587f
C303 source.n156 a_n2390_n3288# 0.023881f
C304 source.n157 a_n2390_n3288# 0.012833f
C305 source.n158 a_n2390_n3288# 0.022749f
C306 source.n159 a_n2390_n3288# 0.021442f
C307 source.t19 a_n2390_n3288# 0.051228f
C308 source.n160 a_n2390_n3288# 0.17218f
C309 source.n161 a_n2390_n3288# 1.20476f
C310 source.n162 a_n2390_n3288# 0.012833f
C311 source.n163 a_n2390_n3288# 0.013587f
C312 source.n164 a_n2390_n3288# 0.030332f
C313 source.n165 a_n2390_n3288# 0.030332f
C314 source.n166 a_n2390_n3288# 0.013587f
C315 source.n167 a_n2390_n3288# 0.012833f
C316 source.n168 a_n2390_n3288# 0.023881f
C317 source.n169 a_n2390_n3288# 0.023881f
C318 source.n170 a_n2390_n3288# 0.012833f
C319 source.n171 a_n2390_n3288# 0.013587f
C320 source.n172 a_n2390_n3288# 0.030332f
C321 source.n173 a_n2390_n3288# 0.030332f
C322 source.n174 a_n2390_n3288# 0.013587f
C323 source.n175 a_n2390_n3288# 0.012833f
C324 source.n176 a_n2390_n3288# 0.023881f
C325 source.n177 a_n2390_n3288# 0.023881f
C326 source.n178 a_n2390_n3288# 0.012833f
C327 source.n179 a_n2390_n3288# 0.013587f
C328 source.n180 a_n2390_n3288# 0.030332f
C329 source.n181 a_n2390_n3288# 0.030332f
C330 source.n182 a_n2390_n3288# 0.030332f
C331 source.n183 a_n2390_n3288# 0.01321f
C332 source.n184 a_n2390_n3288# 0.012833f
C333 source.n185 a_n2390_n3288# 0.023881f
C334 source.n186 a_n2390_n3288# 0.023881f
C335 source.n187 a_n2390_n3288# 0.012833f
C336 source.n188 a_n2390_n3288# 0.013587f
C337 source.n189 a_n2390_n3288# 0.030332f
C338 source.n190 a_n2390_n3288# 0.030332f
C339 source.n191 a_n2390_n3288# 0.013587f
C340 source.n192 a_n2390_n3288# 0.012833f
C341 source.n193 a_n2390_n3288# 0.023881f
C342 source.n194 a_n2390_n3288# 0.023881f
C343 source.n195 a_n2390_n3288# 0.012833f
C344 source.n196 a_n2390_n3288# 0.013587f
C345 source.n197 a_n2390_n3288# 0.030332f
C346 source.n198 a_n2390_n3288# 0.062244f
C347 source.n199 a_n2390_n3288# 0.013587f
C348 source.n200 a_n2390_n3288# 0.012833f
C349 source.n201 a_n2390_n3288# 0.051285f
C350 source.n202 a_n2390_n3288# 0.034352f
C351 source.n203 a_n2390_n3288# 0.116037f
C352 source.t20 a_n2390_n3288# 0.226459f
C353 source.t23 a_n2390_n3288# 0.226459f
C354 source.n204 a_n2390_n3288# 1.93895f
C355 source.n205 a_n2390_n3288# 0.36754f
C356 source.t28 a_n2390_n3288# 0.226459f
C357 source.t31 a_n2390_n3288# 0.226459f
C358 source.n206 a_n2390_n3288# 1.93895f
C359 source.n207 a_n2390_n3288# 0.36754f
C360 source.t24 a_n2390_n3288# 0.226459f
C361 source.t29 a_n2390_n3288# 0.226459f
C362 source.n208 a_n2390_n3288# 1.93895f
C363 source.n209 a_n2390_n3288# 0.36754f
C364 source.n210 a_n2390_n3288# 0.031634f
C365 source.n211 a_n2390_n3288# 0.023881f
C366 source.n212 a_n2390_n3288# 0.012833f
C367 source.n213 a_n2390_n3288# 0.030332f
C368 source.n214 a_n2390_n3288# 0.013587f
C369 source.n215 a_n2390_n3288# 0.023881f
C370 source.n216 a_n2390_n3288# 0.012833f
C371 source.n217 a_n2390_n3288# 0.030332f
C372 source.n218 a_n2390_n3288# 0.013587f
C373 source.n219 a_n2390_n3288# 0.023881f
C374 source.n220 a_n2390_n3288# 0.01321f
C375 source.n221 a_n2390_n3288# 0.030332f
C376 source.n222 a_n2390_n3288# 0.012833f
C377 source.n223 a_n2390_n3288# 0.013587f
C378 source.n224 a_n2390_n3288# 0.023881f
C379 source.n225 a_n2390_n3288# 0.012833f
C380 source.n226 a_n2390_n3288# 0.030332f
C381 source.n227 a_n2390_n3288# 0.013587f
C382 source.n228 a_n2390_n3288# 0.023881f
C383 source.n229 a_n2390_n3288# 0.012833f
C384 source.n230 a_n2390_n3288# 0.022749f
C385 source.n231 a_n2390_n3288# 0.021442f
C386 source.t26 a_n2390_n3288# 0.051228f
C387 source.n232 a_n2390_n3288# 0.17218f
C388 source.n233 a_n2390_n3288# 1.20476f
C389 source.n234 a_n2390_n3288# 0.012833f
C390 source.n235 a_n2390_n3288# 0.013587f
C391 source.n236 a_n2390_n3288# 0.030332f
C392 source.n237 a_n2390_n3288# 0.030332f
C393 source.n238 a_n2390_n3288# 0.013587f
C394 source.n239 a_n2390_n3288# 0.012833f
C395 source.n240 a_n2390_n3288# 0.023881f
C396 source.n241 a_n2390_n3288# 0.023881f
C397 source.n242 a_n2390_n3288# 0.012833f
C398 source.n243 a_n2390_n3288# 0.013587f
C399 source.n244 a_n2390_n3288# 0.030332f
C400 source.n245 a_n2390_n3288# 0.030332f
C401 source.n246 a_n2390_n3288# 0.013587f
C402 source.n247 a_n2390_n3288# 0.012833f
C403 source.n248 a_n2390_n3288# 0.023881f
C404 source.n249 a_n2390_n3288# 0.023881f
C405 source.n250 a_n2390_n3288# 0.012833f
C406 source.n251 a_n2390_n3288# 0.013587f
C407 source.n252 a_n2390_n3288# 0.030332f
C408 source.n253 a_n2390_n3288# 0.030332f
C409 source.n254 a_n2390_n3288# 0.030332f
C410 source.n255 a_n2390_n3288# 0.01321f
C411 source.n256 a_n2390_n3288# 0.012833f
C412 source.n257 a_n2390_n3288# 0.023881f
C413 source.n258 a_n2390_n3288# 0.023881f
C414 source.n259 a_n2390_n3288# 0.012833f
C415 source.n260 a_n2390_n3288# 0.013587f
C416 source.n261 a_n2390_n3288# 0.030332f
C417 source.n262 a_n2390_n3288# 0.030332f
C418 source.n263 a_n2390_n3288# 0.013587f
C419 source.n264 a_n2390_n3288# 0.012833f
C420 source.n265 a_n2390_n3288# 0.023881f
C421 source.n266 a_n2390_n3288# 0.023881f
C422 source.n267 a_n2390_n3288# 0.012833f
C423 source.n268 a_n2390_n3288# 0.013587f
C424 source.n269 a_n2390_n3288# 0.030332f
C425 source.n270 a_n2390_n3288# 0.062244f
C426 source.n271 a_n2390_n3288# 0.013587f
C427 source.n272 a_n2390_n3288# 0.012833f
C428 source.n273 a_n2390_n3288# 0.051285f
C429 source.n274 a_n2390_n3288# 0.034352f
C430 source.n275 a_n2390_n3288# 1.37641f
C431 source.n276 a_n2390_n3288# 0.031634f
C432 source.n277 a_n2390_n3288# 0.023881f
C433 source.n278 a_n2390_n3288# 0.012833f
C434 source.n279 a_n2390_n3288# 0.030332f
C435 source.n280 a_n2390_n3288# 0.013587f
C436 source.n281 a_n2390_n3288# 0.023881f
C437 source.n282 a_n2390_n3288# 0.012833f
C438 source.n283 a_n2390_n3288# 0.030332f
C439 source.n284 a_n2390_n3288# 0.013587f
C440 source.n285 a_n2390_n3288# 0.023881f
C441 source.n286 a_n2390_n3288# 0.01321f
C442 source.n287 a_n2390_n3288# 0.030332f
C443 source.n288 a_n2390_n3288# 0.013587f
C444 source.n289 a_n2390_n3288# 0.023881f
C445 source.n290 a_n2390_n3288# 0.012833f
C446 source.n291 a_n2390_n3288# 0.030332f
C447 source.n292 a_n2390_n3288# 0.013587f
C448 source.n293 a_n2390_n3288# 0.023881f
C449 source.n294 a_n2390_n3288# 0.012833f
C450 source.n295 a_n2390_n3288# 0.022749f
C451 source.n296 a_n2390_n3288# 0.021442f
C452 source.t5 a_n2390_n3288# 0.051228f
C453 source.n297 a_n2390_n3288# 0.17218f
C454 source.n298 a_n2390_n3288# 1.20476f
C455 source.n299 a_n2390_n3288# 0.012833f
C456 source.n300 a_n2390_n3288# 0.013587f
C457 source.n301 a_n2390_n3288# 0.030332f
C458 source.n302 a_n2390_n3288# 0.030332f
C459 source.n303 a_n2390_n3288# 0.013587f
C460 source.n304 a_n2390_n3288# 0.012833f
C461 source.n305 a_n2390_n3288# 0.023881f
C462 source.n306 a_n2390_n3288# 0.023881f
C463 source.n307 a_n2390_n3288# 0.012833f
C464 source.n308 a_n2390_n3288# 0.013587f
C465 source.n309 a_n2390_n3288# 0.030332f
C466 source.n310 a_n2390_n3288# 0.030332f
C467 source.n311 a_n2390_n3288# 0.013587f
C468 source.n312 a_n2390_n3288# 0.012833f
C469 source.n313 a_n2390_n3288# 0.023881f
C470 source.n314 a_n2390_n3288# 0.023881f
C471 source.n315 a_n2390_n3288# 0.012833f
C472 source.n316 a_n2390_n3288# 0.012833f
C473 source.n317 a_n2390_n3288# 0.013587f
C474 source.n318 a_n2390_n3288# 0.030332f
C475 source.n319 a_n2390_n3288# 0.030332f
C476 source.n320 a_n2390_n3288# 0.030332f
C477 source.n321 a_n2390_n3288# 0.01321f
C478 source.n322 a_n2390_n3288# 0.012833f
C479 source.n323 a_n2390_n3288# 0.023881f
C480 source.n324 a_n2390_n3288# 0.023881f
C481 source.n325 a_n2390_n3288# 0.012833f
C482 source.n326 a_n2390_n3288# 0.013587f
C483 source.n327 a_n2390_n3288# 0.030332f
C484 source.n328 a_n2390_n3288# 0.030332f
C485 source.n329 a_n2390_n3288# 0.013587f
C486 source.n330 a_n2390_n3288# 0.012833f
C487 source.n331 a_n2390_n3288# 0.023881f
C488 source.n332 a_n2390_n3288# 0.023881f
C489 source.n333 a_n2390_n3288# 0.012833f
C490 source.n334 a_n2390_n3288# 0.013587f
C491 source.n335 a_n2390_n3288# 0.030332f
C492 source.n336 a_n2390_n3288# 0.062244f
C493 source.n337 a_n2390_n3288# 0.013587f
C494 source.n338 a_n2390_n3288# 0.012833f
C495 source.n339 a_n2390_n3288# 0.051285f
C496 source.n340 a_n2390_n3288# 0.034352f
C497 source.n341 a_n2390_n3288# 1.37641f
C498 source.t12 a_n2390_n3288# 0.226459f
C499 source.t15 a_n2390_n3288# 0.226459f
C500 source.n342 a_n2390_n3288# 1.93893f
C501 source.n343 a_n2390_n3288# 0.367552f
C502 source.t9 a_n2390_n3288# 0.226459f
C503 source.t13 a_n2390_n3288# 0.226459f
C504 source.n344 a_n2390_n3288# 1.93893f
C505 source.n345 a_n2390_n3288# 0.367552f
C506 source.t0 a_n2390_n3288# 0.226459f
C507 source.t10 a_n2390_n3288# 0.226459f
C508 source.n346 a_n2390_n3288# 1.93893f
C509 source.n347 a_n2390_n3288# 0.367552f
C510 source.n348 a_n2390_n3288# 0.031634f
C511 source.n349 a_n2390_n3288# 0.023881f
C512 source.n350 a_n2390_n3288# 0.012833f
C513 source.n351 a_n2390_n3288# 0.030332f
C514 source.n352 a_n2390_n3288# 0.013587f
C515 source.n353 a_n2390_n3288# 0.023881f
C516 source.n354 a_n2390_n3288# 0.012833f
C517 source.n355 a_n2390_n3288# 0.030332f
C518 source.n356 a_n2390_n3288# 0.013587f
C519 source.n357 a_n2390_n3288# 0.023881f
C520 source.n358 a_n2390_n3288# 0.01321f
C521 source.n359 a_n2390_n3288# 0.030332f
C522 source.n360 a_n2390_n3288# 0.013587f
C523 source.n361 a_n2390_n3288# 0.023881f
C524 source.n362 a_n2390_n3288# 0.012833f
C525 source.n363 a_n2390_n3288# 0.030332f
C526 source.n364 a_n2390_n3288# 0.013587f
C527 source.n365 a_n2390_n3288# 0.023881f
C528 source.n366 a_n2390_n3288# 0.012833f
C529 source.n367 a_n2390_n3288# 0.022749f
C530 source.n368 a_n2390_n3288# 0.021442f
C531 source.t2 a_n2390_n3288# 0.051228f
C532 source.n369 a_n2390_n3288# 0.17218f
C533 source.n370 a_n2390_n3288# 1.20476f
C534 source.n371 a_n2390_n3288# 0.012833f
C535 source.n372 a_n2390_n3288# 0.013587f
C536 source.n373 a_n2390_n3288# 0.030332f
C537 source.n374 a_n2390_n3288# 0.030332f
C538 source.n375 a_n2390_n3288# 0.013587f
C539 source.n376 a_n2390_n3288# 0.012833f
C540 source.n377 a_n2390_n3288# 0.023881f
C541 source.n378 a_n2390_n3288# 0.023881f
C542 source.n379 a_n2390_n3288# 0.012833f
C543 source.n380 a_n2390_n3288# 0.013587f
C544 source.n381 a_n2390_n3288# 0.030332f
C545 source.n382 a_n2390_n3288# 0.030332f
C546 source.n383 a_n2390_n3288# 0.013587f
C547 source.n384 a_n2390_n3288# 0.012833f
C548 source.n385 a_n2390_n3288# 0.023881f
C549 source.n386 a_n2390_n3288# 0.023881f
C550 source.n387 a_n2390_n3288# 0.012833f
C551 source.n388 a_n2390_n3288# 0.012833f
C552 source.n389 a_n2390_n3288# 0.013587f
C553 source.n390 a_n2390_n3288# 0.030332f
C554 source.n391 a_n2390_n3288# 0.030332f
C555 source.n392 a_n2390_n3288# 0.030332f
C556 source.n393 a_n2390_n3288# 0.01321f
C557 source.n394 a_n2390_n3288# 0.012833f
C558 source.n395 a_n2390_n3288# 0.023881f
C559 source.n396 a_n2390_n3288# 0.023881f
C560 source.n397 a_n2390_n3288# 0.012833f
C561 source.n398 a_n2390_n3288# 0.013587f
C562 source.n399 a_n2390_n3288# 0.030332f
C563 source.n400 a_n2390_n3288# 0.030332f
C564 source.n401 a_n2390_n3288# 0.013587f
C565 source.n402 a_n2390_n3288# 0.012833f
C566 source.n403 a_n2390_n3288# 0.023881f
C567 source.n404 a_n2390_n3288# 0.023881f
C568 source.n405 a_n2390_n3288# 0.012833f
C569 source.n406 a_n2390_n3288# 0.013587f
C570 source.n407 a_n2390_n3288# 0.030332f
C571 source.n408 a_n2390_n3288# 0.062244f
C572 source.n409 a_n2390_n3288# 0.013587f
C573 source.n410 a_n2390_n3288# 0.012833f
C574 source.n411 a_n2390_n3288# 0.051285f
C575 source.n412 a_n2390_n3288# 0.034352f
C576 source.n413 a_n2390_n3288# 0.116037f
C577 source.n414 a_n2390_n3288# 0.031634f
C578 source.n415 a_n2390_n3288# 0.023881f
C579 source.n416 a_n2390_n3288# 0.012833f
C580 source.n417 a_n2390_n3288# 0.030332f
C581 source.n418 a_n2390_n3288# 0.013587f
C582 source.n419 a_n2390_n3288# 0.023881f
C583 source.n420 a_n2390_n3288# 0.012833f
C584 source.n421 a_n2390_n3288# 0.030332f
C585 source.n422 a_n2390_n3288# 0.013587f
C586 source.n423 a_n2390_n3288# 0.023881f
C587 source.n424 a_n2390_n3288# 0.01321f
C588 source.n425 a_n2390_n3288# 0.030332f
C589 source.n426 a_n2390_n3288# 0.013587f
C590 source.n427 a_n2390_n3288# 0.023881f
C591 source.n428 a_n2390_n3288# 0.012833f
C592 source.n429 a_n2390_n3288# 0.030332f
C593 source.n430 a_n2390_n3288# 0.013587f
C594 source.n431 a_n2390_n3288# 0.023881f
C595 source.n432 a_n2390_n3288# 0.012833f
C596 source.n433 a_n2390_n3288# 0.022749f
C597 source.n434 a_n2390_n3288# 0.021442f
C598 source.t25 a_n2390_n3288# 0.051228f
C599 source.n435 a_n2390_n3288# 0.17218f
C600 source.n436 a_n2390_n3288# 1.20476f
C601 source.n437 a_n2390_n3288# 0.012833f
C602 source.n438 a_n2390_n3288# 0.013587f
C603 source.n439 a_n2390_n3288# 0.030332f
C604 source.n440 a_n2390_n3288# 0.030332f
C605 source.n441 a_n2390_n3288# 0.013587f
C606 source.n442 a_n2390_n3288# 0.012833f
C607 source.n443 a_n2390_n3288# 0.023881f
C608 source.n444 a_n2390_n3288# 0.023881f
C609 source.n445 a_n2390_n3288# 0.012833f
C610 source.n446 a_n2390_n3288# 0.013587f
C611 source.n447 a_n2390_n3288# 0.030332f
C612 source.n448 a_n2390_n3288# 0.030332f
C613 source.n449 a_n2390_n3288# 0.013587f
C614 source.n450 a_n2390_n3288# 0.012833f
C615 source.n451 a_n2390_n3288# 0.023881f
C616 source.n452 a_n2390_n3288# 0.023881f
C617 source.n453 a_n2390_n3288# 0.012833f
C618 source.n454 a_n2390_n3288# 0.012833f
C619 source.n455 a_n2390_n3288# 0.013587f
C620 source.n456 a_n2390_n3288# 0.030332f
C621 source.n457 a_n2390_n3288# 0.030332f
C622 source.n458 a_n2390_n3288# 0.030332f
C623 source.n459 a_n2390_n3288# 0.01321f
C624 source.n460 a_n2390_n3288# 0.012833f
C625 source.n461 a_n2390_n3288# 0.023881f
C626 source.n462 a_n2390_n3288# 0.023881f
C627 source.n463 a_n2390_n3288# 0.012833f
C628 source.n464 a_n2390_n3288# 0.013587f
C629 source.n465 a_n2390_n3288# 0.030332f
C630 source.n466 a_n2390_n3288# 0.030332f
C631 source.n467 a_n2390_n3288# 0.013587f
C632 source.n468 a_n2390_n3288# 0.012833f
C633 source.n469 a_n2390_n3288# 0.023881f
C634 source.n470 a_n2390_n3288# 0.023881f
C635 source.n471 a_n2390_n3288# 0.012833f
C636 source.n472 a_n2390_n3288# 0.013587f
C637 source.n473 a_n2390_n3288# 0.030332f
C638 source.n474 a_n2390_n3288# 0.062244f
C639 source.n475 a_n2390_n3288# 0.013587f
C640 source.n476 a_n2390_n3288# 0.012833f
C641 source.n477 a_n2390_n3288# 0.051285f
C642 source.n478 a_n2390_n3288# 0.034352f
C643 source.n479 a_n2390_n3288# 0.116037f
C644 source.t16 a_n2390_n3288# 0.226459f
C645 source.t22 a_n2390_n3288# 0.226459f
C646 source.n480 a_n2390_n3288# 1.93893f
C647 source.n481 a_n2390_n3288# 0.367552f
C648 source.t30 a_n2390_n3288# 0.226459f
C649 source.t27 a_n2390_n3288# 0.226459f
C650 source.n482 a_n2390_n3288# 1.93893f
C651 source.n483 a_n2390_n3288# 0.367552f
C652 source.t17 a_n2390_n3288# 0.226459f
C653 source.t21 a_n2390_n3288# 0.226459f
C654 source.n484 a_n2390_n3288# 1.93893f
C655 source.n485 a_n2390_n3288# 0.367552f
C656 source.n486 a_n2390_n3288# 0.031634f
C657 source.n487 a_n2390_n3288# 0.023881f
C658 source.n488 a_n2390_n3288# 0.012833f
C659 source.n489 a_n2390_n3288# 0.030332f
C660 source.n490 a_n2390_n3288# 0.013587f
C661 source.n491 a_n2390_n3288# 0.023881f
C662 source.n492 a_n2390_n3288# 0.012833f
C663 source.n493 a_n2390_n3288# 0.030332f
C664 source.n494 a_n2390_n3288# 0.013587f
C665 source.n495 a_n2390_n3288# 0.023881f
C666 source.n496 a_n2390_n3288# 0.01321f
C667 source.n497 a_n2390_n3288# 0.030332f
C668 source.n498 a_n2390_n3288# 0.013587f
C669 source.n499 a_n2390_n3288# 0.023881f
C670 source.n500 a_n2390_n3288# 0.012833f
C671 source.n501 a_n2390_n3288# 0.030332f
C672 source.n502 a_n2390_n3288# 0.013587f
C673 source.n503 a_n2390_n3288# 0.023881f
C674 source.n504 a_n2390_n3288# 0.012833f
C675 source.n505 a_n2390_n3288# 0.022749f
C676 source.n506 a_n2390_n3288# 0.021442f
C677 source.t18 a_n2390_n3288# 0.051228f
C678 source.n507 a_n2390_n3288# 0.17218f
C679 source.n508 a_n2390_n3288# 1.20476f
C680 source.n509 a_n2390_n3288# 0.012833f
C681 source.n510 a_n2390_n3288# 0.013587f
C682 source.n511 a_n2390_n3288# 0.030332f
C683 source.n512 a_n2390_n3288# 0.030332f
C684 source.n513 a_n2390_n3288# 0.013587f
C685 source.n514 a_n2390_n3288# 0.012833f
C686 source.n515 a_n2390_n3288# 0.023881f
C687 source.n516 a_n2390_n3288# 0.023881f
C688 source.n517 a_n2390_n3288# 0.012833f
C689 source.n518 a_n2390_n3288# 0.013587f
C690 source.n519 a_n2390_n3288# 0.030332f
C691 source.n520 a_n2390_n3288# 0.030332f
C692 source.n521 a_n2390_n3288# 0.013587f
C693 source.n522 a_n2390_n3288# 0.012833f
C694 source.n523 a_n2390_n3288# 0.023881f
C695 source.n524 a_n2390_n3288# 0.023881f
C696 source.n525 a_n2390_n3288# 0.012833f
C697 source.n526 a_n2390_n3288# 0.012833f
C698 source.n527 a_n2390_n3288# 0.013587f
C699 source.n528 a_n2390_n3288# 0.030332f
C700 source.n529 a_n2390_n3288# 0.030332f
C701 source.n530 a_n2390_n3288# 0.030332f
C702 source.n531 a_n2390_n3288# 0.01321f
C703 source.n532 a_n2390_n3288# 0.012833f
C704 source.n533 a_n2390_n3288# 0.023881f
C705 source.n534 a_n2390_n3288# 0.023881f
C706 source.n535 a_n2390_n3288# 0.012833f
C707 source.n536 a_n2390_n3288# 0.013587f
C708 source.n537 a_n2390_n3288# 0.030332f
C709 source.n538 a_n2390_n3288# 0.030332f
C710 source.n539 a_n2390_n3288# 0.013587f
C711 source.n540 a_n2390_n3288# 0.012833f
C712 source.n541 a_n2390_n3288# 0.023881f
C713 source.n542 a_n2390_n3288# 0.023881f
C714 source.n543 a_n2390_n3288# 0.012833f
C715 source.n544 a_n2390_n3288# 0.013587f
C716 source.n545 a_n2390_n3288# 0.030332f
C717 source.n546 a_n2390_n3288# 0.062244f
C718 source.n547 a_n2390_n3288# 0.013587f
C719 source.n548 a_n2390_n3288# 0.012833f
C720 source.n549 a_n2390_n3288# 0.051285f
C721 source.n550 a_n2390_n3288# 0.034352f
C722 source.n551 a_n2390_n3288# 0.266617f
C723 source.n552 a_n2390_n3288# 1.50946f
C724 minus.n0 a_n2390_n3288# 0.042712f
C725 minus.t6 a_n2390_n3288# 0.876919f
C726 minus.n1 a_n2390_n3288# 0.353637f
C727 minus.n2 a_n2390_n3288# 0.042712f
C728 minus.t8 a_n2390_n3288# 0.876919f
C729 minus.n3 a_n2390_n3288# 0.353637f
C730 minus.n4 a_n2390_n3288# 0.042712f
C731 minus.t12 a_n2390_n3288# 0.876919f
C732 minus.n5 a_n2390_n3288# 0.352452f
C733 minus.t13 a_n2390_n3288# 0.889906f
C734 minus.n6 a_n2390_n3288# 0.339148f
C735 minus.n7 a_n2390_n3288# 0.143858f
C736 minus.n8 a_n2390_n3288# 0.009692f
C737 minus.t10 a_n2390_n3288# 0.876919f
C738 minus.n9 a_n2390_n3288# 0.353637f
C739 minus.n10 a_n2390_n3288# 0.009692f
C740 minus.n11 a_n2390_n3288# 0.042712f
C741 minus.n12 a_n2390_n3288# 0.042712f
C742 minus.n13 a_n2390_n3288# 0.042712f
C743 minus.n14 a_n2390_n3288# 0.009692f
C744 minus.t4 a_n2390_n3288# 0.876919f
C745 minus.n15 a_n2390_n3288# 0.353637f
C746 minus.n16 a_n2390_n3288# 0.009692f
C747 minus.n17 a_n2390_n3288# 0.042712f
C748 minus.n18 a_n2390_n3288# 0.042712f
C749 minus.n19 a_n2390_n3288# 0.042712f
C750 minus.n20 a_n2390_n3288# 0.009692f
C751 minus.t5 a_n2390_n3288# 0.876919f
C752 minus.n21 a_n2390_n3288# 0.352452f
C753 minus.t3 a_n2390_n3288# 0.876919f
C754 minus.n22 a_n2390_n3288# 0.351793f
C755 minus.n23 a_n2390_n3288# 1.65416f
C756 minus.n24 a_n2390_n3288# 0.042712f
C757 minus.t0 a_n2390_n3288# 0.876919f
C758 minus.n25 a_n2390_n3288# 0.353637f
C759 minus.n26 a_n2390_n3288# 0.042712f
C760 minus.t15 a_n2390_n3288# 0.876919f
C761 minus.n27 a_n2390_n3288# 0.353637f
C762 minus.n28 a_n2390_n3288# 0.042712f
C763 minus.t2 a_n2390_n3288# 0.876919f
C764 minus.n29 a_n2390_n3288# 0.352452f
C765 minus.t11 a_n2390_n3288# 0.889906f
C766 minus.n30 a_n2390_n3288# 0.339148f
C767 minus.n31 a_n2390_n3288# 0.143858f
C768 minus.n32 a_n2390_n3288# 0.009692f
C769 minus.t7 a_n2390_n3288# 0.876919f
C770 minus.n33 a_n2390_n3288# 0.353637f
C771 minus.n34 a_n2390_n3288# 0.009692f
C772 minus.n35 a_n2390_n3288# 0.042712f
C773 minus.n36 a_n2390_n3288# 0.042712f
C774 minus.n37 a_n2390_n3288# 0.042712f
C775 minus.n38 a_n2390_n3288# 0.009692f
C776 minus.t1 a_n2390_n3288# 0.876919f
C777 minus.n39 a_n2390_n3288# 0.353637f
C778 minus.n40 a_n2390_n3288# 0.009692f
C779 minus.n41 a_n2390_n3288# 0.042712f
C780 minus.n42 a_n2390_n3288# 0.042712f
C781 minus.n43 a_n2390_n3288# 0.042712f
C782 minus.n44 a_n2390_n3288# 0.009692f
C783 minus.t9 a_n2390_n3288# 0.876919f
C784 minus.n45 a_n2390_n3288# 0.352452f
C785 minus.t14 a_n2390_n3288# 0.876919f
C786 minus.n46 a_n2390_n3288# 0.351793f
C787 minus.n47 a_n2390_n3288# 0.294806f
C788 minus.n48 a_n2390_n3288# 1.99207f
.ends

