* NGSPICE file created from diffpair608.ext - technology: sky130A

.subckt diffpair608 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t25 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t27 plus.t1 drain_left.t18 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 drain_right.t19 minus.t0 source.t9 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X3 a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X4 source.t36 plus.t2 drain_left.t17 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X5 source.t13 minus.t1 drain_right.t18 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t7 minus.t2 drain_right.t17 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X7 source.t38 plus.t3 drain_left.t16 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 source.t26 plus.t4 drain_left.t15 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X9 drain_left.t14 plus.t5 source.t34 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 source.t33 plus.t6 drain_left.t13 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X11 source.t8 minus.t3 drain_right.t16 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X12 drain_right.t15 minus.t4 source.t19 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X13 source.t10 minus.t5 drain_right.t14 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X14 drain_right.t13 minus.t6 source.t3 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 drain_right.t12 minus.t7 source.t5 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X16 source.t11 minus.t8 drain_right.t11 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X17 a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X18 drain_left.t12 plus.t7 source.t24 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 drain_left.t11 plus.t8 source.t29 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X20 drain_left.t10 plus.t9 source.t23 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X21 source.t32 plus.t10 drain_left.t9 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X22 source.t14 minus.t9 drain_right.t10 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 drain_right.t9 minus.t10 source.t0 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X24 source.t16 minus.t11 drain_right.t8 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X25 drain_left.t8 plus.t11 source.t22 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X26 source.t30 plus.t12 drain_left.t7 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X27 source.t35 plus.t13 drain_left.t6 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X28 drain_right.t7 minus.t12 source.t2 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X29 drain_left.t5 plus.t14 source.t28 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X30 drain_right.t6 minus.t13 source.t1 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X31 source.t18 minus.t14 drain_right.t5 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X32 drain_left.t4 plus.t15 source.t31 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X33 drain_right.t4 minus.t15 source.t4 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X34 a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X35 source.t17 minus.t16 drain_right.t3 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X36 drain_right.t2 minus.t17 source.t6 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X37 source.t12 minus.t18 drain_right.t1 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X38 source.t21 plus.t16 drain_left.t3 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X39 drain_right.t0 minus.t19 source.t15 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X40 drain_left.t2 plus.t17 source.t20 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X41 source.t37 plus.t18 drain_left.t1 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X42 a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X43 drain_left.t0 plus.t19 source.t39 a_n2542_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
R0 plus.n8 plus.t6 1063.55
R1 plus.n36 plus.t0 1063.55
R2 plus.n26 plus.t14 1042.57
R3 plus.n25 plus.t3 1042.57
R4 plus.n1 plus.t17 1042.57
R5 plus.n19 plus.t10 1042.57
R6 plus.n18 plus.t19 1042.57
R7 plus.n4 plus.t16 1042.57
R8 plus.n13 plus.t7 1042.57
R9 plus.n11 plus.t18 1042.57
R10 plus.n7 plus.t15 1042.57
R11 plus.n54 plus.t12 1042.57
R12 plus.n53 plus.t11 1042.57
R13 plus.n29 plus.t2 1042.57
R14 plus.n47 plus.t8 1042.57
R15 plus.n46 plus.t13 1042.57
R16 plus.n32 plus.t5 1042.57
R17 plus.n41 plus.t4 1042.57
R18 plus.n39 plus.t9 1042.57
R19 plus.n35 plus.t1 1042.57
R20 plus.n10 plus.n9 161.3
R21 plus.n11 plus.n6 161.3
R22 plus.n12 plus.n5 161.3
R23 plus.n14 plus.n13 161.3
R24 plus.n15 plus.n4 161.3
R25 plus.n17 plus.n16 161.3
R26 plus.n18 plus.n3 161.3
R27 plus.n19 plus.n2 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n22 plus.n1 161.3
R30 plus.n24 plus.n23 161.3
R31 plus.n25 plus.n0 161.3
R32 plus.n27 plus.n26 161.3
R33 plus.n38 plus.n37 161.3
R34 plus.n39 plus.n34 161.3
R35 plus.n40 plus.n33 161.3
R36 plus.n42 plus.n41 161.3
R37 plus.n43 plus.n32 161.3
R38 plus.n45 plus.n44 161.3
R39 plus.n46 plus.n31 161.3
R40 plus.n47 plus.n30 161.3
R41 plus.n49 plus.n48 161.3
R42 plus.n50 plus.n29 161.3
R43 plus.n52 plus.n51 161.3
R44 plus.n53 plus.n28 161.3
R45 plus.n55 plus.n54 161.3
R46 plus.n9 plus.n8 70.4033
R47 plus.n37 plus.n36 70.4033
R48 plus.n26 plus.n25 48.2005
R49 plus.n19 plus.n18 48.2005
R50 plus.n13 plus.n4 48.2005
R51 plus.n54 plus.n53 48.2005
R52 plus.n47 plus.n46 48.2005
R53 plus.n41 plus.n32 48.2005
R54 plus.n20 plus.n1 47.4702
R55 plus.n12 plus.n11 47.4702
R56 plus.n48 plus.n29 47.4702
R57 plus.n40 plus.n39 47.4702
R58 plus plus.n55 35.7528
R59 plus.n24 plus.n1 25.5611
R60 plus.n11 plus.n10 25.5611
R61 plus.n52 plus.n29 25.5611
R62 plus.n39 plus.n38 25.5611
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n25 plus.n24 22.6399
R68 plus.n10 plus.n7 22.6399
R69 plus.n53 plus.n52 22.6399
R70 plus.n38 plus.n35 22.6399
R71 plus.n8 plus.n7 20.9576
R72 plus.n36 plus.n35 20.9576
R73 plus plus.n27 15.2657
R74 plus.n20 plus.n19 0.730803
R75 plus.n13 plus.n12 0.730803
R76 plus.n48 plus.n47 0.730803
R77 plus.n41 plus.n40 0.730803
R78 plus.n9 plus.n6 0.189894
R79 plus.n6 plus.n5 0.189894
R80 plus.n14 plus.n5 0.189894
R81 plus.n15 plus.n14 0.189894
R82 plus.n16 plus.n15 0.189894
R83 plus.n16 plus.n3 0.189894
R84 plus.n3 plus.n2 0.189894
R85 plus.n21 plus.n2 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n23 plus.n22 0.189894
R88 plus.n23 plus.n0 0.189894
R89 plus.n27 plus.n0 0.189894
R90 plus.n55 plus.n28 0.189894
R91 plus.n51 plus.n28 0.189894
R92 plus.n51 plus.n50 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n30 0.189894
R95 plus.n31 plus.n30 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n34 plus.n33 0.189894
R101 plus.n37 plus.n34 0.189894
R102 source.n0 source.t28 44.1297
R103 source.n9 source.t33 44.1296
R104 source.n10 source.t1 44.1296
R105 source.n19 source.t8 44.1296
R106 source.n39 source.t15 44.1295
R107 source.n30 source.t10 44.1295
R108 source.n29 source.t25 44.1295
R109 source.n20 source.t30 44.1295
R110 source.n2 source.n1 43.1397
R111 source.n4 source.n3 43.1397
R112 source.n6 source.n5 43.1397
R113 source.n8 source.n7 43.1397
R114 source.n12 source.n11 43.1397
R115 source.n14 source.n13 43.1397
R116 source.n16 source.n15 43.1397
R117 source.n18 source.n17 43.1397
R118 source.n38 source.n37 43.1396
R119 source.n36 source.n35 43.1396
R120 source.n34 source.n33 43.1396
R121 source.n32 source.n31 43.1396
R122 source.n28 source.n27 43.1396
R123 source.n26 source.n25 43.1396
R124 source.n24 source.n23 43.1396
R125 source.n22 source.n21 43.1396
R126 source.n20 source.n19 28.0638
R127 source.n40 source.n0 22.4432
R128 source.n40 source.n39 5.62119
R129 source.n37 source.t0 0.9905
R130 source.n37 source.t7 0.9905
R131 source.n35 source.t6 0.9905
R132 source.n35 source.t17 0.9905
R133 source.n33 source.t2 0.9905
R134 source.n33 source.t11 0.9905
R135 source.n31 source.t19 0.9905
R136 source.n31 source.t18 0.9905
R137 source.n27 source.t23 0.9905
R138 source.n27 source.t27 0.9905
R139 source.n25 source.t34 0.9905
R140 source.n25 source.t26 0.9905
R141 source.n23 source.t29 0.9905
R142 source.n23 source.t35 0.9905
R143 source.n21 source.t22 0.9905
R144 source.n21 source.t36 0.9905
R145 source.n1 source.t20 0.9905
R146 source.n1 source.t38 0.9905
R147 source.n3 source.t39 0.9905
R148 source.n3 source.t32 0.9905
R149 source.n5 source.t24 0.9905
R150 source.n5 source.t21 0.9905
R151 source.n7 source.t31 0.9905
R152 source.n7 source.t37 0.9905
R153 source.n11 source.t5 0.9905
R154 source.n11 source.t13 0.9905
R155 source.n13 source.t3 0.9905
R156 source.n13 source.t12 0.9905
R157 source.n15 source.t9 0.9905
R158 source.n15 source.t14 0.9905
R159 source.n17 source.t4 0.9905
R160 source.n17 source.t16 0.9905
R161 source.n19 source.n18 0.716017
R162 source.n18 source.n16 0.716017
R163 source.n16 source.n14 0.716017
R164 source.n14 source.n12 0.716017
R165 source.n12 source.n10 0.716017
R166 source.n9 source.n8 0.716017
R167 source.n8 source.n6 0.716017
R168 source.n6 source.n4 0.716017
R169 source.n4 source.n2 0.716017
R170 source.n2 source.n0 0.716017
R171 source.n22 source.n20 0.716017
R172 source.n24 source.n22 0.716017
R173 source.n26 source.n24 0.716017
R174 source.n28 source.n26 0.716017
R175 source.n29 source.n28 0.716017
R176 source.n32 source.n30 0.716017
R177 source.n34 source.n32 0.716017
R178 source.n36 source.n34 0.716017
R179 source.n38 source.n36 0.716017
R180 source.n39 source.n38 0.716017
R181 source.n10 source.n9 0.470328
R182 source.n30 source.n29 0.470328
R183 source source.n40 0.188
R184 drain_left.n10 drain_left.n8 60.534
R185 drain_left.n6 drain_left.n4 60.5339
R186 drain_left.n2 drain_left.n0 60.5339
R187 drain_left.n16 drain_left.n15 59.8185
R188 drain_left.n14 drain_left.n13 59.8185
R189 drain_left.n12 drain_left.n11 59.8185
R190 drain_left.n10 drain_left.n9 59.8185
R191 drain_left.n7 drain_left.n3 59.8184
R192 drain_left.n6 drain_left.n5 59.8184
R193 drain_left.n2 drain_left.n1 59.8184
R194 drain_left drain_left.n7 39.1518
R195 drain_left drain_left.n16 6.36873
R196 drain_left.n3 drain_left.t6 0.9905
R197 drain_left.n3 drain_left.t14 0.9905
R198 drain_left.n4 drain_left.t18 0.9905
R199 drain_left.n4 drain_left.t19 0.9905
R200 drain_left.n5 drain_left.t15 0.9905
R201 drain_left.n5 drain_left.t10 0.9905
R202 drain_left.n1 drain_left.t17 0.9905
R203 drain_left.n1 drain_left.t11 0.9905
R204 drain_left.n0 drain_left.t7 0.9905
R205 drain_left.n0 drain_left.t8 0.9905
R206 drain_left.n15 drain_left.t16 0.9905
R207 drain_left.n15 drain_left.t5 0.9905
R208 drain_left.n13 drain_left.t9 0.9905
R209 drain_left.n13 drain_left.t2 0.9905
R210 drain_left.n11 drain_left.t3 0.9905
R211 drain_left.n11 drain_left.t0 0.9905
R212 drain_left.n9 drain_left.t1 0.9905
R213 drain_left.n9 drain_left.t12 0.9905
R214 drain_left.n8 drain_left.t13 0.9905
R215 drain_left.n8 drain_left.t4 0.9905
R216 drain_left.n12 drain_left.n10 0.716017
R217 drain_left.n14 drain_left.n12 0.716017
R218 drain_left.n16 drain_left.n14 0.716017
R219 drain_left.n7 drain_left.n6 0.660671
R220 drain_left.n7 drain_left.n2 0.660671
R221 minus.n6 minus.t13 1063.55
R222 minus.n34 minus.t5 1063.55
R223 minus.n7 minus.t1 1042.57
R224 minus.n5 minus.t7 1042.57
R225 minus.n13 minus.t18 1042.57
R226 minus.n14 minus.t6 1042.57
R227 minus.n18 minus.t9 1042.57
R228 minus.n19 minus.t0 1042.57
R229 minus.n1 minus.t11 1042.57
R230 minus.n25 minus.t15 1042.57
R231 minus.n26 minus.t3 1042.57
R232 minus.n35 minus.t4 1042.57
R233 minus.n33 minus.t14 1042.57
R234 minus.n41 minus.t12 1042.57
R235 minus.n42 minus.t8 1042.57
R236 minus.n46 minus.t17 1042.57
R237 minus.n47 minus.t16 1042.57
R238 minus.n29 minus.t10 1042.57
R239 minus.n53 minus.t2 1042.57
R240 minus.n54 minus.t19 1042.57
R241 minus.n27 minus.n26 161.3
R242 minus.n25 minus.n0 161.3
R243 minus.n24 minus.n23 161.3
R244 minus.n22 minus.n1 161.3
R245 minus.n21 minus.n20 161.3
R246 minus.n19 minus.n2 161.3
R247 minus.n18 minus.n17 161.3
R248 minus.n16 minus.n3 161.3
R249 minus.n15 minus.n14 161.3
R250 minus.n13 minus.n4 161.3
R251 minus.n12 minus.n11 161.3
R252 minus.n10 minus.n5 161.3
R253 minus.n9 minus.n8 161.3
R254 minus.n55 minus.n54 161.3
R255 minus.n53 minus.n28 161.3
R256 minus.n52 minus.n51 161.3
R257 minus.n50 minus.n29 161.3
R258 minus.n49 minus.n48 161.3
R259 minus.n47 minus.n30 161.3
R260 minus.n46 minus.n45 161.3
R261 minus.n44 minus.n31 161.3
R262 minus.n43 minus.n42 161.3
R263 minus.n41 minus.n32 161.3
R264 minus.n40 minus.n39 161.3
R265 minus.n38 minus.n33 161.3
R266 minus.n37 minus.n36 161.3
R267 minus.n9 minus.n6 70.4033
R268 minus.n37 minus.n34 70.4033
R269 minus.n14 minus.n13 48.2005
R270 minus.n19 minus.n18 48.2005
R271 minus.n26 minus.n25 48.2005
R272 minus.n42 minus.n41 48.2005
R273 minus.n47 minus.n46 48.2005
R274 minus.n54 minus.n53 48.2005
R275 minus.n12 minus.n5 47.4702
R276 minus.n20 minus.n1 47.4702
R277 minus.n40 minus.n33 47.4702
R278 minus.n48 minus.n29 47.4702
R279 minus.n56 minus.n27 44.902
R280 minus.n8 minus.n5 25.5611
R281 minus.n24 minus.n1 25.5611
R282 minus.n36 minus.n33 25.5611
R283 minus.n52 minus.n29 25.5611
R284 minus.n18 minus.n3 24.1005
R285 minus.n14 minus.n3 24.1005
R286 minus.n42 minus.n31 24.1005
R287 minus.n46 minus.n31 24.1005
R288 minus.n8 minus.n7 22.6399
R289 minus.n25 minus.n24 22.6399
R290 minus.n36 minus.n35 22.6399
R291 minus.n53 minus.n52 22.6399
R292 minus.n7 minus.n6 20.9576
R293 minus.n35 minus.n34 20.9576
R294 minus.n56 minus.n55 6.59141
R295 minus.n13 minus.n12 0.730803
R296 minus.n20 minus.n19 0.730803
R297 minus.n41 minus.n40 0.730803
R298 minus.n48 minus.n47 0.730803
R299 minus.n27 minus.n0 0.189894
R300 minus.n23 minus.n0 0.189894
R301 minus.n23 minus.n22 0.189894
R302 minus.n22 minus.n21 0.189894
R303 minus.n21 minus.n2 0.189894
R304 minus.n17 minus.n2 0.189894
R305 minus.n17 minus.n16 0.189894
R306 minus.n16 minus.n15 0.189894
R307 minus.n15 minus.n4 0.189894
R308 minus.n11 minus.n4 0.189894
R309 minus.n11 minus.n10 0.189894
R310 minus.n10 minus.n9 0.189894
R311 minus.n38 minus.n37 0.189894
R312 minus.n39 minus.n38 0.189894
R313 minus.n39 minus.n32 0.189894
R314 minus.n43 minus.n32 0.189894
R315 minus.n44 minus.n43 0.189894
R316 minus.n45 minus.n44 0.189894
R317 minus.n45 minus.n30 0.189894
R318 minus.n49 minus.n30 0.189894
R319 minus.n50 minus.n49 0.189894
R320 minus.n51 minus.n50 0.189894
R321 minus.n51 minus.n28 0.189894
R322 minus.n55 minus.n28 0.189894
R323 minus minus.n56 0.188
R324 drain_right.n10 drain_right.n8 60.534
R325 drain_right.n6 drain_right.n4 60.5339
R326 drain_right.n2 drain_right.n0 60.5339
R327 drain_right.n10 drain_right.n9 59.8185
R328 drain_right.n12 drain_right.n11 59.8185
R329 drain_right.n14 drain_right.n13 59.8185
R330 drain_right.n16 drain_right.n15 59.8185
R331 drain_right.n7 drain_right.n3 59.8184
R332 drain_right.n6 drain_right.n5 59.8184
R333 drain_right.n2 drain_right.n1 59.8184
R334 drain_right drain_right.n7 38.5986
R335 drain_right drain_right.n16 6.36873
R336 drain_right.n3 drain_right.t11 0.9905
R337 drain_right.n3 drain_right.t2 0.9905
R338 drain_right.n4 drain_right.t17 0.9905
R339 drain_right.n4 drain_right.t0 0.9905
R340 drain_right.n5 drain_right.t3 0.9905
R341 drain_right.n5 drain_right.t9 0.9905
R342 drain_right.n1 drain_right.t5 0.9905
R343 drain_right.n1 drain_right.t7 0.9905
R344 drain_right.n0 drain_right.t14 0.9905
R345 drain_right.n0 drain_right.t15 0.9905
R346 drain_right.n8 drain_right.t18 0.9905
R347 drain_right.n8 drain_right.t6 0.9905
R348 drain_right.n9 drain_right.t1 0.9905
R349 drain_right.n9 drain_right.t12 0.9905
R350 drain_right.n11 drain_right.t10 0.9905
R351 drain_right.n11 drain_right.t13 0.9905
R352 drain_right.n13 drain_right.t8 0.9905
R353 drain_right.n13 drain_right.t19 0.9905
R354 drain_right.n15 drain_right.t16 0.9905
R355 drain_right.n15 drain_right.t4 0.9905
R356 drain_right.n16 drain_right.n14 0.716017
R357 drain_right.n14 drain_right.n12 0.716017
R358 drain_right.n12 drain_right.n10 0.716017
R359 drain_right.n7 drain_right.n6 0.660671
R360 drain_right.n7 drain_right.n2 0.660671
C0 drain_left plus 16.899801f
C1 source drain_right 45.452698f
C2 minus plus 7.80147f
C3 drain_left minus 0.173163f
C4 drain_right plus 0.40825f
C5 source plus 16.325901f
C6 drain_left drain_right 1.35855f
C7 source drain_left 45.451397f
C8 drain_right minus 16.648f
C9 source minus 16.3119f
C10 drain_right a_n2542_n4888# 8.557309f
C11 drain_left a_n2542_n4888# 8.92526f
C12 source a_n2542_n4888# 13.521109f
C13 minus a_n2542_n4888# 10.658384f
C14 plus a_n2542_n4888# 13.01473f
C15 drain_right.t14 a_n2542_n4888# 0.465565f
C16 drain_right.t15 a_n2542_n4888# 0.465565f
C17 drain_right.n0 a_n2542_n4888# 4.26098f
C18 drain_right.t5 a_n2542_n4888# 0.465565f
C19 drain_right.t7 a_n2542_n4888# 0.465565f
C20 drain_right.n1 a_n2542_n4888# 4.2563f
C21 drain_right.n2 a_n2542_n4888# 0.771785f
C22 drain_right.t11 a_n2542_n4888# 0.465565f
C23 drain_right.t2 a_n2542_n4888# 0.465565f
C24 drain_right.n3 a_n2542_n4888# 4.2563f
C25 drain_right.t17 a_n2542_n4888# 0.465565f
C26 drain_right.t0 a_n2542_n4888# 0.465565f
C27 drain_right.n4 a_n2542_n4888# 4.26098f
C28 drain_right.t3 a_n2542_n4888# 0.465565f
C29 drain_right.t9 a_n2542_n4888# 0.465565f
C30 drain_right.n5 a_n2542_n4888# 4.2563f
C31 drain_right.n6 a_n2542_n4888# 0.771785f
C32 drain_right.n7 a_n2542_n4888# 2.50678f
C33 drain_right.t18 a_n2542_n4888# 0.465565f
C34 drain_right.t6 a_n2542_n4888# 0.465565f
C35 drain_right.n8 a_n2542_n4888# 4.26098f
C36 drain_right.t1 a_n2542_n4888# 0.465565f
C37 drain_right.t12 a_n2542_n4888# 0.465565f
C38 drain_right.n9 a_n2542_n4888# 4.25629f
C39 drain_right.n10 a_n2542_n4888# 0.776016f
C40 drain_right.t10 a_n2542_n4888# 0.465565f
C41 drain_right.t13 a_n2542_n4888# 0.465565f
C42 drain_right.n11 a_n2542_n4888# 4.25629f
C43 drain_right.n12 a_n2542_n4888# 0.384418f
C44 drain_right.t8 a_n2542_n4888# 0.465565f
C45 drain_right.t19 a_n2542_n4888# 0.465565f
C46 drain_right.n13 a_n2542_n4888# 4.25629f
C47 drain_right.n14 a_n2542_n4888# 0.384418f
C48 drain_right.t16 a_n2542_n4888# 0.465565f
C49 drain_right.t4 a_n2542_n4888# 0.465565f
C50 drain_right.n15 a_n2542_n4888# 4.25629f
C51 drain_right.n16 a_n2542_n4888# 0.637499f
C52 minus.n0 a_n2542_n4888# 0.043985f
C53 minus.t11 a_n2542_n4888# 1.2456f
C54 minus.n1 a_n2542_n4888# 0.472524f
C55 minus.n2 a_n2542_n4888# 0.043985f
C56 minus.n3 a_n2542_n4888# 0.009981f
C57 minus.t9 a_n2542_n4888# 1.2456f
C58 minus.n4 a_n2542_n4888# 0.043985f
C59 minus.t7 a_n2542_n4888# 1.2456f
C60 minus.n5 a_n2542_n4888# 0.472524f
C61 minus.t13 a_n2542_n4888# 1.25483f
C62 minus.n6 a_n2542_n4888# 0.459019f
C63 minus.t1 a_n2542_n4888# 1.2456f
C64 minus.n7 a_n2542_n4888# 0.472117f
C65 minus.n8 a_n2542_n4888# 0.009981f
C66 minus.n9 a_n2542_n4888# 0.144363f
C67 minus.n10 a_n2542_n4888# 0.043985f
C68 minus.n11 a_n2542_n4888# 0.043985f
C69 minus.n12 a_n2542_n4888# 0.009981f
C70 minus.t18 a_n2542_n4888# 1.2456f
C71 minus.n13 a_n2542_n4888# 0.468049f
C72 minus.t6 a_n2542_n4888# 1.2456f
C73 minus.n14 a_n2542_n4888# 0.472388f
C74 minus.n15 a_n2542_n4888# 0.043985f
C75 minus.n16 a_n2542_n4888# 0.043985f
C76 minus.n17 a_n2542_n4888# 0.043985f
C77 minus.n18 a_n2542_n4888# 0.472388f
C78 minus.t0 a_n2542_n4888# 1.2456f
C79 minus.n19 a_n2542_n4888# 0.468049f
C80 minus.n20 a_n2542_n4888# 0.009981f
C81 minus.n21 a_n2542_n4888# 0.043985f
C82 minus.n22 a_n2542_n4888# 0.043985f
C83 minus.n23 a_n2542_n4888# 0.043985f
C84 minus.n24 a_n2542_n4888# 0.009981f
C85 minus.t15 a_n2542_n4888# 1.2456f
C86 minus.n25 a_n2542_n4888# 0.472117f
C87 minus.t3 a_n2542_n4888# 1.2456f
C88 minus.n26 a_n2542_n4888# 0.467914f
C89 minus.n27 a_n2542_n4888# 2.14924f
C90 minus.n28 a_n2542_n4888# 0.043985f
C91 minus.t10 a_n2542_n4888# 1.2456f
C92 minus.n29 a_n2542_n4888# 0.472524f
C93 minus.n30 a_n2542_n4888# 0.043985f
C94 minus.n31 a_n2542_n4888# 0.009981f
C95 minus.n32 a_n2542_n4888# 0.043985f
C96 minus.t14 a_n2542_n4888# 1.2456f
C97 minus.n33 a_n2542_n4888# 0.472524f
C98 minus.t5 a_n2542_n4888# 1.25483f
C99 minus.n34 a_n2542_n4888# 0.459019f
C100 minus.t4 a_n2542_n4888# 1.2456f
C101 minus.n35 a_n2542_n4888# 0.472117f
C102 minus.n36 a_n2542_n4888# 0.009981f
C103 minus.n37 a_n2542_n4888# 0.144363f
C104 minus.n38 a_n2542_n4888# 0.043985f
C105 minus.n39 a_n2542_n4888# 0.043985f
C106 minus.n40 a_n2542_n4888# 0.009981f
C107 minus.t12 a_n2542_n4888# 1.2456f
C108 minus.n41 a_n2542_n4888# 0.468049f
C109 minus.t8 a_n2542_n4888# 1.2456f
C110 minus.n42 a_n2542_n4888# 0.472388f
C111 minus.n43 a_n2542_n4888# 0.043985f
C112 minus.n44 a_n2542_n4888# 0.043985f
C113 minus.n45 a_n2542_n4888# 0.043985f
C114 minus.t17 a_n2542_n4888# 1.2456f
C115 minus.n46 a_n2542_n4888# 0.472388f
C116 minus.t16 a_n2542_n4888# 1.2456f
C117 minus.n47 a_n2542_n4888# 0.468049f
C118 minus.n48 a_n2542_n4888# 0.009981f
C119 minus.n49 a_n2542_n4888# 0.043985f
C120 minus.n50 a_n2542_n4888# 0.043985f
C121 minus.n51 a_n2542_n4888# 0.043985f
C122 minus.n52 a_n2542_n4888# 0.009981f
C123 minus.t2 a_n2542_n4888# 1.2456f
C124 minus.n53 a_n2542_n4888# 0.472117f
C125 minus.t19 a_n2542_n4888# 1.2456f
C126 minus.n54 a_n2542_n4888# 0.467914f
C127 minus.n55 a_n2542_n4888# 0.296992f
C128 minus.n56 a_n2542_n4888# 2.54401f
C129 drain_left.t7 a_n2542_n4888# 0.466948f
C130 drain_left.t8 a_n2542_n4888# 0.466948f
C131 drain_left.n0 a_n2542_n4888# 4.27364f
C132 drain_left.t17 a_n2542_n4888# 0.466948f
C133 drain_left.t11 a_n2542_n4888# 0.466948f
C134 drain_left.n1 a_n2542_n4888# 4.26894f
C135 drain_left.n2 a_n2542_n4888# 0.774077f
C136 drain_left.t6 a_n2542_n4888# 0.466948f
C137 drain_left.t14 a_n2542_n4888# 0.466948f
C138 drain_left.n3 a_n2542_n4888# 4.26894f
C139 drain_left.t18 a_n2542_n4888# 0.466948f
C140 drain_left.t19 a_n2542_n4888# 0.466948f
C141 drain_left.n4 a_n2542_n4888# 4.27364f
C142 drain_left.t15 a_n2542_n4888# 0.466948f
C143 drain_left.t10 a_n2542_n4888# 0.466948f
C144 drain_left.n5 a_n2542_n4888# 4.26894f
C145 drain_left.n6 a_n2542_n4888# 0.774077f
C146 drain_left.n7 a_n2542_n4888# 2.57512f
C147 drain_left.t13 a_n2542_n4888# 0.466948f
C148 drain_left.t4 a_n2542_n4888# 0.466948f
C149 drain_left.n8 a_n2542_n4888# 4.27363f
C150 drain_left.t1 a_n2542_n4888# 0.466948f
C151 drain_left.t12 a_n2542_n4888# 0.466948f
C152 drain_left.n9 a_n2542_n4888# 4.26893f
C153 drain_left.n10 a_n2542_n4888# 0.778321f
C154 drain_left.t3 a_n2542_n4888# 0.466948f
C155 drain_left.t0 a_n2542_n4888# 0.466948f
C156 drain_left.n11 a_n2542_n4888# 4.26893f
C157 drain_left.n12 a_n2542_n4888# 0.385559f
C158 drain_left.t9 a_n2542_n4888# 0.466948f
C159 drain_left.t2 a_n2542_n4888# 0.466948f
C160 drain_left.n13 a_n2542_n4888# 4.26893f
C161 drain_left.n14 a_n2542_n4888# 0.385559f
C162 drain_left.t16 a_n2542_n4888# 0.466948f
C163 drain_left.t5 a_n2542_n4888# 0.466948f
C164 drain_left.n15 a_n2542_n4888# 4.26893f
C165 drain_left.n16 a_n2542_n4888# 0.639392f
C166 source.t28 a_n2542_n4888# 4.55041f
C167 source.n0 a_n2542_n4888# 1.9575f
C168 source.t20 a_n2542_n4888# 0.398168f
C169 source.t38 a_n2542_n4888# 0.398168f
C170 source.n1 a_n2542_n4888# 3.55979f
C171 source.n2 a_n2542_n4888# 0.374867f
C172 source.t39 a_n2542_n4888# 0.398168f
C173 source.t32 a_n2542_n4888# 0.398168f
C174 source.n3 a_n2542_n4888# 3.55979f
C175 source.n4 a_n2542_n4888# 0.374867f
C176 source.t24 a_n2542_n4888# 0.398168f
C177 source.t21 a_n2542_n4888# 0.398168f
C178 source.n5 a_n2542_n4888# 3.55979f
C179 source.n6 a_n2542_n4888# 0.374867f
C180 source.t31 a_n2542_n4888# 0.398168f
C181 source.t37 a_n2542_n4888# 0.398168f
C182 source.n7 a_n2542_n4888# 3.55979f
C183 source.n8 a_n2542_n4888# 0.374867f
C184 source.t33 a_n2542_n4888# 4.55042f
C185 source.n9 a_n2542_n4888# 0.450203f
C186 source.t1 a_n2542_n4888# 4.55042f
C187 source.n10 a_n2542_n4888# 0.450203f
C188 source.t5 a_n2542_n4888# 0.398168f
C189 source.t13 a_n2542_n4888# 0.398168f
C190 source.n11 a_n2542_n4888# 3.55979f
C191 source.n12 a_n2542_n4888# 0.374867f
C192 source.t3 a_n2542_n4888# 0.398168f
C193 source.t12 a_n2542_n4888# 0.398168f
C194 source.n13 a_n2542_n4888# 3.55979f
C195 source.n14 a_n2542_n4888# 0.374867f
C196 source.t9 a_n2542_n4888# 0.398168f
C197 source.t14 a_n2542_n4888# 0.398168f
C198 source.n15 a_n2542_n4888# 3.55979f
C199 source.n16 a_n2542_n4888# 0.374867f
C200 source.t4 a_n2542_n4888# 0.398168f
C201 source.t16 a_n2542_n4888# 0.398168f
C202 source.n17 a_n2542_n4888# 3.55979f
C203 source.n18 a_n2542_n4888# 0.374867f
C204 source.t8 a_n2542_n4888# 4.55042f
C205 source.n19 a_n2542_n4888# 2.40989f
C206 source.t30 a_n2542_n4888# 4.5504f
C207 source.n20 a_n2542_n4888# 2.40991f
C208 source.t22 a_n2542_n4888# 0.398168f
C209 source.t36 a_n2542_n4888# 0.398168f
C210 source.n21 a_n2542_n4888# 3.5598f
C211 source.n22 a_n2542_n4888# 0.37486f
C212 source.t29 a_n2542_n4888# 0.398168f
C213 source.t35 a_n2542_n4888# 0.398168f
C214 source.n23 a_n2542_n4888# 3.5598f
C215 source.n24 a_n2542_n4888# 0.37486f
C216 source.t34 a_n2542_n4888# 0.398168f
C217 source.t26 a_n2542_n4888# 0.398168f
C218 source.n25 a_n2542_n4888# 3.5598f
C219 source.n26 a_n2542_n4888# 0.37486f
C220 source.t23 a_n2542_n4888# 0.398168f
C221 source.t27 a_n2542_n4888# 0.398168f
C222 source.n27 a_n2542_n4888# 3.5598f
C223 source.n28 a_n2542_n4888# 0.37486f
C224 source.t25 a_n2542_n4888# 4.5504f
C225 source.n29 a_n2542_n4888# 0.450228f
C226 source.t10 a_n2542_n4888# 4.5504f
C227 source.n30 a_n2542_n4888# 0.450228f
C228 source.t19 a_n2542_n4888# 0.398168f
C229 source.t18 a_n2542_n4888# 0.398168f
C230 source.n31 a_n2542_n4888# 3.5598f
C231 source.n32 a_n2542_n4888# 0.37486f
C232 source.t2 a_n2542_n4888# 0.398168f
C233 source.t11 a_n2542_n4888# 0.398168f
C234 source.n33 a_n2542_n4888# 3.5598f
C235 source.n34 a_n2542_n4888# 0.37486f
C236 source.t6 a_n2542_n4888# 0.398168f
C237 source.t17 a_n2542_n4888# 0.398168f
C238 source.n35 a_n2542_n4888# 3.5598f
C239 source.n36 a_n2542_n4888# 0.37486f
C240 source.t0 a_n2542_n4888# 0.398168f
C241 source.t7 a_n2542_n4888# 0.398168f
C242 source.n37 a_n2542_n4888# 3.5598f
C243 source.n38 a_n2542_n4888# 0.37486f
C244 source.t15 a_n2542_n4888# 4.5504f
C245 source.n39 a_n2542_n4888# 0.603566f
C246 source.n40 a_n2542_n4888# 2.27666f
C247 plus.n0 a_n2542_n4888# 0.044406f
C248 plus.t14 a_n2542_n4888# 1.25753f
C249 plus.t3 a_n2542_n4888# 1.25753f
C250 plus.t17 a_n2542_n4888# 1.25753f
C251 plus.n1 a_n2542_n4888# 0.477049f
C252 plus.n2 a_n2542_n4888# 0.044406f
C253 plus.t10 a_n2542_n4888# 1.25753f
C254 plus.t19 a_n2542_n4888# 1.25753f
C255 plus.n3 a_n2542_n4888# 0.044406f
C256 plus.t16 a_n2542_n4888# 1.25753f
C257 plus.n4 a_n2542_n4888# 0.476912f
C258 plus.n5 a_n2542_n4888# 0.044406f
C259 plus.t7 a_n2542_n4888# 1.25753f
C260 plus.t18 a_n2542_n4888# 1.25753f
C261 plus.n6 a_n2542_n4888# 0.044406f
C262 plus.t15 a_n2542_n4888# 1.25753f
C263 plus.n7 a_n2542_n4888# 0.476639f
C264 plus.t6 a_n2542_n4888# 1.26685f
C265 plus.n8 a_n2542_n4888# 0.463415f
C266 plus.n9 a_n2542_n4888# 0.145745f
C267 plus.n10 a_n2542_n4888# 0.010077f
C268 plus.n11 a_n2542_n4888# 0.477049f
C269 plus.n12 a_n2542_n4888# 0.010077f
C270 plus.n13 a_n2542_n4888# 0.472532f
C271 plus.n14 a_n2542_n4888# 0.044406f
C272 plus.n15 a_n2542_n4888# 0.044406f
C273 plus.n16 a_n2542_n4888# 0.044406f
C274 plus.n17 a_n2542_n4888# 0.010077f
C275 plus.n18 a_n2542_n4888# 0.476912f
C276 plus.n19 a_n2542_n4888# 0.472532f
C277 plus.n20 a_n2542_n4888# 0.010077f
C278 plus.n21 a_n2542_n4888# 0.044406f
C279 plus.n22 a_n2542_n4888# 0.044406f
C280 plus.n23 a_n2542_n4888# 0.044406f
C281 plus.n24 a_n2542_n4888# 0.010077f
C282 plus.n25 a_n2542_n4888# 0.476639f
C283 plus.n26 a_n2542_n4888# 0.472395f
C284 plus.n27 a_n2542_n4888# 0.683596f
C285 plus.n28 a_n2542_n4888# 0.044406f
C286 plus.t12 a_n2542_n4888# 1.25753f
C287 plus.t11 a_n2542_n4888# 1.25753f
C288 plus.t2 a_n2542_n4888# 1.25753f
C289 plus.n29 a_n2542_n4888# 0.477049f
C290 plus.n30 a_n2542_n4888# 0.044406f
C291 plus.t8 a_n2542_n4888# 1.25753f
C292 plus.n31 a_n2542_n4888# 0.044406f
C293 plus.t13 a_n2542_n4888# 1.25753f
C294 plus.t5 a_n2542_n4888# 1.25753f
C295 plus.n32 a_n2542_n4888# 0.476912f
C296 plus.n33 a_n2542_n4888# 0.044406f
C297 plus.t4 a_n2542_n4888# 1.25753f
C298 plus.n34 a_n2542_n4888# 0.044406f
C299 plus.t9 a_n2542_n4888# 1.25753f
C300 plus.t1 a_n2542_n4888# 1.25753f
C301 plus.n35 a_n2542_n4888# 0.476639f
C302 plus.t0 a_n2542_n4888# 1.26685f
C303 plus.n36 a_n2542_n4888# 0.463415f
C304 plus.n37 a_n2542_n4888# 0.145745f
C305 plus.n38 a_n2542_n4888# 0.010077f
C306 plus.n39 a_n2542_n4888# 0.477049f
C307 plus.n40 a_n2542_n4888# 0.010077f
C308 plus.n41 a_n2542_n4888# 0.472532f
C309 plus.n42 a_n2542_n4888# 0.044406f
C310 plus.n43 a_n2542_n4888# 0.044406f
C311 plus.n44 a_n2542_n4888# 0.044406f
C312 plus.n45 a_n2542_n4888# 0.010077f
C313 plus.n46 a_n2542_n4888# 0.476912f
C314 plus.n47 a_n2542_n4888# 0.472532f
C315 plus.n48 a_n2542_n4888# 0.010077f
C316 plus.n49 a_n2542_n4888# 0.044406f
C317 plus.n50 a_n2542_n4888# 0.044406f
C318 plus.n51 a_n2542_n4888# 0.044406f
C319 plus.n52 a_n2542_n4888# 0.010077f
C320 plus.n53 a_n2542_n4888# 0.476639f
C321 plus.n54 a_n2542_n4888# 0.472395f
C322 plus.n55 a_n2542_n4888# 1.73578f
.ends

