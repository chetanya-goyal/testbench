* NGSPICE file created from diffpair133.ext - technology: sky130A

.subckt diffpair133 minus drain_right drain_left source plus
X0 a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X2 a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X3 source.t14 plus.t0 drain_left.t7 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X4 drain_right.t7 minus.t0 source.t15 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X5 source.t1 minus.t1 drain_right.t6 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_left.t6 plus.t1 source.t13 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 source.t12 plus.t2 drain_left.t0 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X8 source.t6 minus.t2 drain_right.t5 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_right.t4 minus.t3 source.t5 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X10 a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X11 drain_left.t1 plus.t3 source.t11 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X12 source.t4 minus.t4 drain_right.t3 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X13 source.t10 plus.t4 drain_left.t2 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 drain_right.t2 minus.t5 source.t0 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X15 source.t3 minus.t6 drain_right.t1 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 drain_left.t3 plus.t5 source.t9 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 source.t8 plus.t6 drain_left.t4 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X18 drain_right.t0 minus.t7 source.t2 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 drain_left.t5 plus.t7 source.t7 a_n1646_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
R0 plus.n1 plus.t6 172.626
R1 plus.n7 plus.t7 172.626
R2 plus.n5 plus.n4 161.3
R3 plus.n11 plus.n10 161.3
R4 plus.n4 plus.t3 145.805
R5 plus.n3 plus.t4 145.805
R6 plus.n2 plus.t5 145.805
R7 plus.n10 plus.t0 145.805
R8 plus.n9 plus.t1 145.805
R9 plus.n8 plus.t2 145.805
R10 plus.n3 plus.n0 80.6037
R11 plus.n9 plus.n6 80.6037
R12 plus.n4 plus.n3 48.2005
R13 plus.n3 plus.n2 48.2005
R14 plus.n10 plus.n9 48.2005
R15 plus.n9 plus.n8 48.2005
R16 plus.n1 plus.n0 45.2318
R17 plus.n7 plus.n6 45.2318
R18 plus plus.n11 25.5634
R19 plus.n2 plus.n1 13.3799
R20 plus.n8 plus.n7 13.3799
R21 plus plus.n5 8.4702
R22 plus.n5 plus.n0 0.285035
R23 plus.n11 plus.n6 0.285035
R24 drain_left.n5 drain_left.n3 101.597
R25 drain_left.n2 drain_left.n1 101.141
R26 drain_left.n2 drain_left.n0 101.141
R27 drain_left.n5 drain_left.n4 100.796
R28 drain_left drain_left.n2 22.5974
R29 drain_left.n1 drain_left.t0 9.9005
R30 drain_left.n1 drain_left.t5 9.9005
R31 drain_left.n0 drain_left.t7 9.9005
R32 drain_left.n0 drain_left.t6 9.9005
R33 drain_left.n4 drain_left.t2 9.9005
R34 drain_left.n4 drain_left.t1 9.9005
R35 drain_left.n3 drain_left.t4 9.9005
R36 drain_left.n3 drain_left.t3 9.9005
R37 drain_left drain_left.n5 6.45494
R38 source.n66 source.n64 289.615
R39 source.n56 source.n54 289.615
R40 source.n48 source.n46 289.615
R41 source.n38 source.n36 289.615
R42 source.n2 source.n0 289.615
R43 source.n12 source.n10 289.615
R44 source.n20 source.n18 289.615
R45 source.n30 source.n28 289.615
R46 source.n67 source.n66 185
R47 source.n57 source.n56 185
R48 source.n49 source.n48 185
R49 source.n39 source.n38 185
R50 source.n3 source.n2 185
R51 source.n13 source.n12 185
R52 source.n21 source.n20 185
R53 source.n31 source.n30 185
R54 source.t15 source.n65 167.117
R55 source.t1 source.n55 167.117
R56 source.t7 source.n47 167.117
R57 source.t14 source.n37 167.117
R58 source.t11 source.n1 167.117
R59 source.t8 source.n11 167.117
R60 source.t0 source.n19 167.117
R61 source.t6 source.n29 167.117
R62 source.n9 source.n8 84.1169
R63 source.n27 source.n26 84.1169
R64 source.n63 source.n62 84.1168
R65 source.n45 source.n44 84.1168
R66 source.n66 source.t15 52.3082
R67 source.n56 source.t1 52.3082
R68 source.n48 source.t7 52.3082
R69 source.n38 source.t14 52.3082
R70 source.n2 source.t11 52.3082
R71 source.n12 source.t8 52.3082
R72 source.n20 source.t0 52.3082
R73 source.n30 source.t6 52.3082
R74 source.n71 source.n70 31.4096
R75 source.n61 source.n60 31.4096
R76 source.n53 source.n52 31.4096
R77 source.n43 source.n42 31.4096
R78 source.n7 source.n6 31.4096
R79 source.n17 source.n16 31.4096
R80 source.n25 source.n24 31.4096
R81 source.n35 source.n34 31.4096
R82 source.n43 source.n35 14.5137
R83 source.n62 source.t2 9.9005
R84 source.n62 source.t3 9.9005
R85 source.n44 source.t13 9.9005
R86 source.n44 source.t12 9.9005
R87 source.n8 source.t9 9.9005
R88 source.n8 source.t10 9.9005
R89 source.n26 source.t5 9.9005
R90 source.n26 source.t4 9.9005
R91 source.n67 source.n65 9.71174
R92 source.n57 source.n55 9.71174
R93 source.n49 source.n47 9.71174
R94 source.n39 source.n37 9.71174
R95 source.n3 source.n1 9.71174
R96 source.n13 source.n11 9.71174
R97 source.n21 source.n19 9.71174
R98 source.n31 source.n29 9.71174
R99 source.n70 source.n69 9.45567
R100 source.n60 source.n59 9.45567
R101 source.n52 source.n51 9.45567
R102 source.n42 source.n41 9.45567
R103 source.n6 source.n5 9.45567
R104 source.n16 source.n15 9.45567
R105 source.n24 source.n23 9.45567
R106 source.n34 source.n33 9.45567
R107 source.n69 source.n68 9.3005
R108 source.n59 source.n58 9.3005
R109 source.n51 source.n50 9.3005
R110 source.n41 source.n40 9.3005
R111 source.n5 source.n4 9.3005
R112 source.n15 source.n14 9.3005
R113 source.n23 source.n22 9.3005
R114 source.n33 source.n32 9.3005
R115 source.n72 source.n7 8.8499
R116 source.n70 source.n64 8.14595
R117 source.n60 source.n54 8.14595
R118 source.n52 source.n46 8.14595
R119 source.n42 source.n36 8.14595
R120 source.n6 source.n0 8.14595
R121 source.n16 source.n10 8.14595
R122 source.n24 source.n18 8.14595
R123 source.n34 source.n28 8.14595
R124 source.n68 source.n67 7.3702
R125 source.n58 source.n57 7.3702
R126 source.n50 source.n49 7.3702
R127 source.n40 source.n39 7.3702
R128 source.n4 source.n3 7.3702
R129 source.n14 source.n13 7.3702
R130 source.n22 source.n21 7.3702
R131 source.n32 source.n31 7.3702
R132 source.n68 source.n64 5.81868
R133 source.n58 source.n54 5.81868
R134 source.n50 source.n46 5.81868
R135 source.n40 source.n36 5.81868
R136 source.n4 source.n0 5.81868
R137 source.n14 source.n10 5.81868
R138 source.n22 source.n18 5.81868
R139 source.n32 source.n28 5.81868
R140 source.n72 source.n71 5.66429
R141 source.n69 source.n65 3.44771
R142 source.n59 source.n55 3.44771
R143 source.n51 source.n47 3.44771
R144 source.n41 source.n37 3.44771
R145 source.n5 source.n1 3.44771
R146 source.n15 source.n11 3.44771
R147 source.n23 source.n19 3.44771
R148 source.n33 source.n29 3.44771
R149 source.n35 source.n27 0.802224
R150 source.n27 source.n25 0.802224
R151 source.n17 source.n9 0.802224
R152 source.n9 source.n7 0.802224
R153 source.n45 source.n43 0.802224
R154 source.n53 source.n45 0.802224
R155 source.n63 source.n61 0.802224
R156 source.n71 source.n63 0.802224
R157 source.n25 source.n17 0.470328
R158 source.n61 source.n53 0.470328
R159 source source.n72 0.188
R160 minus.n1 minus.t5 172.626
R161 minus.n7 minus.t1 172.626
R162 minus.n5 minus.n4 161.3
R163 minus.n11 minus.n10 161.3
R164 minus.n2 minus.t4 145.805
R165 minus.n3 minus.t3 145.805
R166 minus.n4 minus.t2 145.805
R167 minus.n8 minus.t7 145.805
R168 minus.n9 minus.t6 145.805
R169 minus.n10 minus.t0 145.805
R170 minus.n3 minus.n0 80.6037
R171 minus.n9 minus.n6 80.6037
R172 minus.n3 minus.n2 48.2005
R173 minus.n4 minus.n3 48.2005
R174 minus.n9 minus.n8 48.2005
R175 minus.n10 minus.n9 48.2005
R176 minus.n1 minus.n0 45.2318
R177 minus.n7 minus.n6 45.2318
R178 minus.n12 minus.n5 27.8944
R179 minus.n2 minus.n1 13.3799
R180 minus.n8 minus.n7 13.3799
R181 minus.n12 minus.n11 6.61414
R182 minus.n5 minus.n0 0.285035
R183 minus.n11 minus.n6 0.285035
R184 minus minus.n12 0.188
R185 drain_right.n5 drain_right.n3 101.597
R186 drain_right.n2 drain_right.n1 101.141
R187 drain_right.n2 drain_right.n0 101.141
R188 drain_right.n5 drain_right.n4 100.796
R189 drain_right drain_right.n2 22.0441
R190 drain_right.n1 drain_right.t1 9.9005
R191 drain_right.n1 drain_right.t7 9.9005
R192 drain_right.n0 drain_right.t6 9.9005
R193 drain_right.n0 drain_right.t0 9.9005
R194 drain_right.n3 drain_right.t3 9.9005
R195 drain_right.n3 drain_right.t2 9.9005
R196 drain_right.n4 drain_right.t5 9.9005
R197 drain_right.n4 drain_right.t4 9.9005
R198 drain_right drain_right.n5 6.45494
C0 drain_right drain_left 0.775958f
C1 drain_left minus 0.177176f
C2 drain_left plus 1.32097f
C3 drain_right source 3.73695f
C4 source minus 1.38867f
C5 source plus 1.40263f
C6 drain_left source 3.73581f
C7 drain_right minus 1.16259f
C8 drain_right plus 0.319354f
C9 plus minus 3.3513f
C10 drain_right a_n1646_n1288# 3.21806f
C11 drain_left a_n1646_n1288# 3.42317f
C12 source a_n1646_n1288# 3.023582f
C13 minus a_n1646_n1288# 5.549564f
C14 plus a_n1646_n1288# 6.143667f
C15 drain_right.t6 a_n1646_n1288# 0.031112f
C16 drain_right.t0 a_n1646_n1288# 0.031112f
C17 drain_right.n0 a_n1646_n1288# 0.196249f
C18 drain_right.t1 a_n1646_n1288# 0.031112f
C19 drain_right.t7 a_n1646_n1288# 0.031112f
C20 drain_right.n1 a_n1646_n1288# 0.196249f
C21 drain_right.n2 a_n1646_n1288# 0.962285f
C22 drain_right.t3 a_n1646_n1288# 0.031112f
C23 drain_right.t2 a_n1646_n1288# 0.031112f
C24 drain_right.n3 a_n1646_n1288# 0.197509f
C25 drain_right.t5 a_n1646_n1288# 0.031112f
C26 drain_right.t4 a_n1646_n1288# 0.031112f
C27 drain_right.n4 a_n1646_n1288# 0.195455f
C28 drain_right.n5 a_n1646_n1288# 0.68228f
C29 minus.n0 a_n1646_n1288# 0.137029f
C30 minus.t4 a_n1646_n1288# 0.104429f
C31 minus.t5 a_n1646_n1288# 0.115931f
C32 minus.n1 a_n1646_n1288# 0.063289f
C33 minus.n2 a_n1646_n1288# 0.080326f
C34 minus.t3 a_n1646_n1288# 0.104429f
C35 minus.n3 a_n1646_n1288# 0.080326f
C36 minus.t2 a_n1646_n1288# 0.104429f
C37 minus.n4 a_n1646_n1288# 0.073949f
C38 minus.n5 a_n1646_n1288# 0.656702f
C39 minus.n6 a_n1646_n1288# 0.137029f
C40 minus.t1 a_n1646_n1288# 0.115931f
C41 minus.n7 a_n1646_n1288# 0.063289f
C42 minus.t7 a_n1646_n1288# 0.104429f
C43 minus.n8 a_n1646_n1288# 0.080326f
C44 minus.t6 a_n1646_n1288# 0.104429f
C45 minus.n9 a_n1646_n1288# 0.080326f
C46 minus.t0 a_n1646_n1288# 0.104429f
C47 minus.n10 a_n1646_n1288# 0.073949f
C48 minus.n11 a_n1646_n1288# 0.200636f
C49 minus.n12 a_n1646_n1288# 0.795936f
C50 source.n0 a_n1646_n1288# 0.028251f
C51 source.n1 a_n1646_n1288# 0.062508f
C52 source.t11 a_n1646_n1288# 0.046909f
C53 source.n2 a_n1646_n1288# 0.048921f
C54 source.n3 a_n1646_n1288# 0.01577f
C55 source.n4 a_n1646_n1288# 0.010401f
C56 source.n5 a_n1646_n1288# 0.137783f
C57 source.n6 a_n1646_n1288# 0.030969f
C58 source.n7 a_n1646_n1288# 0.320836f
C59 source.t9 a_n1646_n1288# 0.030591f
C60 source.t10 a_n1646_n1288# 0.030591f
C61 source.n8 a_n1646_n1288# 0.163537f
C62 source.n9 a_n1646_n1288# 0.250484f
C63 source.n10 a_n1646_n1288# 0.028251f
C64 source.n11 a_n1646_n1288# 0.062508f
C65 source.t8 a_n1646_n1288# 0.046909f
C66 source.n12 a_n1646_n1288# 0.048921f
C67 source.n13 a_n1646_n1288# 0.01577f
C68 source.n14 a_n1646_n1288# 0.010401f
C69 source.n15 a_n1646_n1288# 0.137783f
C70 source.n16 a_n1646_n1288# 0.030969f
C71 source.n17 a_n1646_n1288# 0.095238f
C72 source.n18 a_n1646_n1288# 0.028251f
C73 source.n19 a_n1646_n1288# 0.062508f
C74 source.t0 a_n1646_n1288# 0.046909f
C75 source.n20 a_n1646_n1288# 0.048921f
C76 source.n21 a_n1646_n1288# 0.01577f
C77 source.n22 a_n1646_n1288# 0.010401f
C78 source.n23 a_n1646_n1288# 0.137783f
C79 source.n24 a_n1646_n1288# 0.030969f
C80 source.n25 a_n1646_n1288# 0.095238f
C81 source.t5 a_n1646_n1288# 0.030591f
C82 source.t4 a_n1646_n1288# 0.030591f
C83 source.n26 a_n1646_n1288# 0.163537f
C84 source.n27 a_n1646_n1288# 0.250484f
C85 source.n28 a_n1646_n1288# 0.028251f
C86 source.n29 a_n1646_n1288# 0.062508f
C87 source.t6 a_n1646_n1288# 0.046909f
C88 source.n30 a_n1646_n1288# 0.048921f
C89 source.n31 a_n1646_n1288# 0.01577f
C90 source.n32 a_n1646_n1288# 0.010401f
C91 source.n33 a_n1646_n1288# 0.137783f
C92 source.n34 a_n1646_n1288# 0.030969f
C93 source.n35 a_n1646_n1288# 0.504949f
C94 source.n36 a_n1646_n1288# 0.028251f
C95 source.n37 a_n1646_n1288# 0.062508f
C96 source.t14 a_n1646_n1288# 0.046909f
C97 source.n38 a_n1646_n1288# 0.048921f
C98 source.n39 a_n1646_n1288# 0.01577f
C99 source.n40 a_n1646_n1288# 0.010401f
C100 source.n41 a_n1646_n1288# 0.137783f
C101 source.n42 a_n1646_n1288# 0.030969f
C102 source.n43 a_n1646_n1288# 0.504949f
C103 source.t13 a_n1646_n1288# 0.030591f
C104 source.t12 a_n1646_n1288# 0.030591f
C105 source.n44 a_n1646_n1288# 0.163536f
C106 source.n45 a_n1646_n1288# 0.250485f
C107 source.n46 a_n1646_n1288# 0.028251f
C108 source.n47 a_n1646_n1288# 0.062508f
C109 source.t7 a_n1646_n1288# 0.046909f
C110 source.n48 a_n1646_n1288# 0.048921f
C111 source.n49 a_n1646_n1288# 0.01577f
C112 source.n50 a_n1646_n1288# 0.010401f
C113 source.n51 a_n1646_n1288# 0.137783f
C114 source.n52 a_n1646_n1288# 0.030969f
C115 source.n53 a_n1646_n1288# 0.095238f
C116 source.n54 a_n1646_n1288# 0.028251f
C117 source.n55 a_n1646_n1288# 0.062508f
C118 source.t1 a_n1646_n1288# 0.046909f
C119 source.n56 a_n1646_n1288# 0.048921f
C120 source.n57 a_n1646_n1288# 0.01577f
C121 source.n58 a_n1646_n1288# 0.010401f
C122 source.n59 a_n1646_n1288# 0.137783f
C123 source.n60 a_n1646_n1288# 0.030969f
C124 source.n61 a_n1646_n1288# 0.095238f
C125 source.t2 a_n1646_n1288# 0.030591f
C126 source.t3 a_n1646_n1288# 0.030591f
C127 source.n62 a_n1646_n1288# 0.163536f
C128 source.n63 a_n1646_n1288# 0.250485f
C129 source.n64 a_n1646_n1288# 0.028251f
C130 source.n65 a_n1646_n1288# 0.062508f
C131 source.t15 a_n1646_n1288# 0.046909f
C132 source.n66 a_n1646_n1288# 0.048921f
C133 source.n67 a_n1646_n1288# 0.01577f
C134 source.n68 a_n1646_n1288# 0.010401f
C135 source.n69 a_n1646_n1288# 0.137783f
C136 source.n70 a_n1646_n1288# 0.030969f
C137 source.n71 a_n1646_n1288# 0.217282f
C138 source.n72 a_n1646_n1288# 0.485546f
C139 drain_left.t7 a_n1646_n1288# 0.030477f
C140 drain_left.t6 a_n1646_n1288# 0.030477f
C141 drain_left.n0 a_n1646_n1288# 0.192248f
C142 drain_left.t0 a_n1646_n1288# 0.030477f
C143 drain_left.t5 a_n1646_n1288# 0.030477f
C144 drain_left.n1 a_n1646_n1288# 0.192248f
C145 drain_left.n2 a_n1646_n1288# 0.980526f
C146 drain_left.t4 a_n1646_n1288# 0.030477f
C147 drain_left.t3 a_n1646_n1288# 0.030477f
C148 drain_left.n3 a_n1646_n1288# 0.193482f
C149 drain_left.t2 a_n1646_n1288# 0.030477f
C150 drain_left.t1 a_n1646_n1288# 0.030477f
C151 drain_left.n4 a_n1646_n1288# 0.19147f
C152 drain_left.n5 a_n1646_n1288# 0.668369f
C153 plus.n0 a_n1646_n1288# 0.139358f
C154 plus.t3 a_n1646_n1288# 0.106204f
C155 plus.t4 a_n1646_n1288# 0.106204f
C156 plus.t5 a_n1646_n1288# 0.106204f
C157 plus.t6 a_n1646_n1288# 0.117901f
C158 plus.n1 a_n1646_n1288# 0.064365f
C159 plus.n2 a_n1646_n1288# 0.081691f
C160 plus.n3 a_n1646_n1288# 0.081691f
C161 plus.n4 a_n1646_n1288# 0.075206f
C162 plus.n5 a_n1646_n1288# 0.22193f
C163 plus.n6 a_n1646_n1288# 0.139358f
C164 plus.t0 a_n1646_n1288# 0.106204f
C165 plus.t1 a_n1646_n1288# 0.106204f
C166 plus.t7 a_n1646_n1288# 0.117901f
C167 plus.n7 a_n1646_n1288# 0.064365f
C168 plus.t2 a_n1646_n1288# 0.106204f
C169 plus.n8 a_n1646_n1288# 0.081691f
C170 plus.n9 a_n1646_n1288# 0.081691f
C171 plus.n10 a_n1646_n1288# 0.075206f
C172 plus.n11 a_n1646_n1288# 0.639522f
.ends

