* NGSPICE file created from diffpair649.ext - technology: sky130A

.subckt diffpair649 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t2 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 drain_right.t1 minus.t1 source.t46 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X2 source.t22 plus.t0 drain_left.t23 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X3 drain_right.t0 minus.t2 source.t45 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X4 source.t44 minus.t3 drain_right.t5 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X5 source.t6 plus.t1 drain_left.t22 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X6 drain_left.t21 plus.t2 source.t2 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X7 drain_left.t20 plus.t3 source.t5 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X8 source.t7 plus.t4 drain_left.t19 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X9 drain_left.t18 plus.t5 source.t10 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X10 a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X11 source.t14 plus.t6 drain_left.t17 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X12 a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X13 source.t43 minus.t4 drain_right.t4 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X14 drain_right.t3 minus.t5 source.t42 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X15 source.t0 plus.t7 drain_left.t16 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X16 drain_left.t15 plus.t8 source.t1 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 drain_right.t20 minus.t6 source.t41 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X18 drain_right.t19 minus.t7 source.t40 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 source.t39 minus.t8 drain_right.t18 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X20 a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X21 source.t38 minus.t9 drain_right.t11 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 drain_left.t14 plus.t9 source.t15 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X23 source.t37 minus.t10 drain_right.t10 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X24 drain_right.t9 minus.t11 source.t36 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X25 drain_left.t13 plus.t10 source.t17 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X26 drain_left.t12 plus.t11 source.t20 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X27 source.t11 plus.t12 drain_left.t11 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X28 drain_right.t8 minus.t12 source.t35 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X29 drain_right.t7 minus.t13 source.t34 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X30 drain_right.t6 minus.t14 source.t33 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X31 source.t16 plus.t13 drain_left.t10 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X32 source.t32 minus.t15 drain_right.t14 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X33 source.t31 minus.t16 drain_right.t13 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X34 drain_left.t9 plus.t14 source.t9 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X35 source.t30 minus.t17 drain_right.t12 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X36 drain_right.t23 minus.t18 source.t29 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X37 drain_right.t22 minus.t19 source.t28 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X38 drain_right.t21 minus.t20 source.t27 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X39 source.t19 plus.t15 drain_left.t8 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X40 drain_left.t7 plus.t16 source.t23 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X41 source.t12 plus.t17 drain_left.t6 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X42 source.t4 plus.t18 drain_left.t5 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X43 source.t26 minus.t21 drain_right.t17 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X44 source.t8 plus.t19 drain_left.t4 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X45 drain_left.t3 plus.t20 source.t13 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X46 drain_left.t2 plus.t21 source.t18 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X47 source.t25 minus.t22 drain_right.t16 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X48 a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X49 drain_left.t1 plus.t22 source.t21 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X50 source.t3 plus.t23 drain_left.t0 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X51 source.t24 minus.t23 drain_right.t15 a_n2406_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
R0 minus.n35 minus.t16 4273
R1 minus.n8 minus.t6 4273
R2 minus.n72 minus.t5 4273
R3 minus.n43 minus.t3 4273
R4 minus.n34 minus.t19 4225.53
R5 minus.n32 minus.t21 4225.53
R6 minus.n3 minus.t11 4225.53
R7 minus.n26 minus.t15 4225.53
R8 minus.n24 minus.t13 4225.53
R9 minus.n6 minus.t17 4225.53
R10 minus.n18 minus.t7 4225.53
R11 minus.n16 minus.t10 4225.53
R12 minus.n9 minus.t12 4225.53
R13 minus.n10 minus.t4 4225.53
R14 minus.n71 minus.t0 4225.53
R15 minus.n69 minus.t20 4225.53
R16 minus.n63 minus.t9 4225.53
R17 minus.n62 minus.t2 4225.53
R18 minus.n60 minus.t23 4225.53
R19 minus.n54 minus.t18 4225.53
R20 minus.n53 minus.t8 4225.53
R21 minus.n51 minus.t1 4225.53
R22 minus.n45 minus.t22 4225.53
R23 minus.n44 minus.t14 4225.53
R24 minus.n12 minus.n8 161.489
R25 minus.n47 minus.n43 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n31 minus.n30 161.3
R29 minus.n29 minus.n1 161.3
R30 minus.n28 minus.n27 161.3
R31 minus.n25 minus.n2 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n20 minus.n19 161.3
R35 minus.n17 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n7 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n68 minus.n67 161.3
R42 minus.n66 minus.n38 161.3
R43 minus.n65 minus.n64 161.3
R44 minus.n61 minus.n39 161.3
R45 minus.n59 minus.n58 161.3
R46 minus.n57 minus.n40 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n52 minus.n41 161.3
R49 minus.n50 minus.n49 161.3
R50 minus.n48 minus.n42 161.3
R51 minus.n47 minus.n46 161.3
R52 minus.n31 minus.n1 73.0308
R53 minus.n23 minus.n4 73.0308
R54 minus.n15 minus.n7 73.0308
R55 minus.n50 minus.n42 73.0308
R56 minus.n59 minus.n40 73.0308
R57 minus.n68 minus.n38 73.0308
R58 minus.n33 minus.n32 69.3793
R59 minus.n11 minus.n9 69.3793
R60 minus.n46 minus.n45 69.3793
R61 minus.n70 minus.n69 69.3793
R62 minus.n25 minus.n24 62.0763
R63 minus.n19 minus.n6 62.0763
R64 minus.n55 minus.n54 62.0763
R65 minus.n61 minus.n60 62.0763
R66 minus.n27 minus.n3 54.7732
R67 minus.n17 minus.n16 54.7732
R68 minus.n52 minus.n51 54.7732
R69 minus.n64 minus.n63 54.7732
R70 minus.n74 minus.n36 48.1066
R71 minus.n35 minus.n34 47.4702
R72 minus.n10 minus.n8 47.4702
R73 minus.n44 minus.n43 47.4702
R74 minus.n72 minus.n71 47.4702
R75 minus.n27 minus.n26 40.1672
R76 minus.n18 minus.n17 40.1672
R77 minus.n53 minus.n52 40.1672
R78 minus.n64 minus.n62 40.1672
R79 minus.n26 minus.n25 32.8641
R80 minus.n19 minus.n18 32.8641
R81 minus.n55 minus.n53 32.8641
R82 minus.n62 minus.n61 32.8641
R83 minus.n34 minus.n33 25.5611
R84 minus.n11 minus.n10 25.5611
R85 minus.n46 minus.n44 25.5611
R86 minus.n71 minus.n70 25.5611
R87 minus.n3 minus.n1 18.2581
R88 minus.n16 minus.n15 18.2581
R89 minus.n51 minus.n50 18.2581
R90 minus.n63 minus.n38 18.2581
R91 minus.n24 minus.n23 10.955
R92 minus.n6 minus.n4 10.955
R93 minus.n54 minus.n40 10.955
R94 minus.n60 minus.n59 10.955
R95 minus.n74 minus.n73 6.52323
R96 minus.n32 minus.n31 3.65202
R97 minus.n9 minus.n7 3.65202
R98 minus.n45 minus.n42 3.65202
R99 minus.n69 minus.n68 3.65202
R100 minus.n36 minus.n0 0.189894
R101 minus.n30 minus.n0 0.189894
R102 minus.n30 minus.n29 0.189894
R103 minus.n29 minus.n28 0.189894
R104 minus.n28 minus.n2 0.189894
R105 minus.n22 minus.n2 0.189894
R106 minus.n22 minus.n21 0.189894
R107 minus.n21 minus.n20 0.189894
R108 minus.n20 minus.n5 0.189894
R109 minus.n14 minus.n5 0.189894
R110 minus.n14 minus.n13 0.189894
R111 minus.n13 minus.n12 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n49 minus.n48 0.189894
R114 minus.n49 minus.n41 0.189894
R115 minus.n56 minus.n41 0.189894
R116 minus.n57 minus.n56 0.189894
R117 minus.n58 minus.n57 0.189894
R118 minus.n58 minus.n39 0.189894
R119 minus.n65 minus.n39 0.189894
R120 minus.n66 minus.n65 0.189894
R121 minus.n67 minus.n66 0.189894
R122 minus.n67 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 drain_right.n7 drain_right.n5 59.2758
R126 drain_right.n2 drain_right.n0 59.2758
R127 drain_right.n13 drain_right.n11 59.2756
R128 drain_right.n7 drain_right.n6 58.7154
R129 drain_right.n9 drain_right.n8 58.7154
R130 drain_right.n4 drain_right.n3 58.7154
R131 drain_right.n2 drain_right.n1 58.7154
R132 drain_right.n13 drain_right.n12 58.7154
R133 drain_right.n15 drain_right.n14 58.7154
R134 drain_right.n17 drain_right.n16 58.7154
R135 drain_right.n19 drain_right.n18 58.7154
R136 drain_right.n21 drain_right.n20 58.7154
R137 drain_right drain_right.n10 41.9856
R138 drain_right drain_right.n21 6.21356
R139 drain_right.n5 drain_right.t2 1.2005
R140 drain_right.n5 drain_right.t3 1.2005
R141 drain_right.n6 drain_right.t11 1.2005
R142 drain_right.n6 drain_right.t21 1.2005
R143 drain_right.n8 drain_right.t15 1.2005
R144 drain_right.n8 drain_right.t0 1.2005
R145 drain_right.n3 drain_right.t18 1.2005
R146 drain_right.n3 drain_right.t23 1.2005
R147 drain_right.n1 drain_right.t16 1.2005
R148 drain_right.n1 drain_right.t1 1.2005
R149 drain_right.n0 drain_right.t5 1.2005
R150 drain_right.n0 drain_right.t6 1.2005
R151 drain_right.n11 drain_right.t4 1.2005
R152 drain_right.n11 drain_right.t20 1.2005
R153 drain_right.n12 drain_right.t10 1.2005
R154 drain_right.n12 drain_right.t8 1.2005
R155 drain_right.n14 drain_right.t12 1.2005
R156 drain_right.n14 drain_right.t19 1.2005
R157 drain_right.n16 drain_right.t14 1.2005
R158 drain_right.n16 drain_right.t7 1.2005
R159 drain_right.n18 drain_right.t17 1.2005
R160 drain_right.n18 drain_right.t9 1.2005
R161 drain_right.n20 drain_right.t13 1.2005
R162 drain_right.n20 drain_right.t22 1.2005
R163 drain_right.n9 drain_right.n7 0.560845
R164 drain_right.n4 drain_right.n2 0.560845
R165 drain_right.n21 drain_right.n19 0.560845
R166 drain_right.n19 drain_right.n17 0.560845
R167 drain_right.n17 drain_right.n15 0.560845
R168 drain_right.n15 drain_right.n13 0.560845
R169 drain_right.n10 drain_right.n9 0.225326
R170 drain_right.n10 drain_right.n4 0.225326
R171 source.n11 source.t11 43.2366
R172 source.n12 source.t41 43.2366
R173 source.n23 source.t31 43.2366
R174 source.n47 source.t42 43.2365
R175 source.n36 source.t44 43.2365
R176 source.n35 source.t15 43.2365
R177 source.n24 source.t14 43.2365
R178 source.n0 source.t21 43.2365
R179 source.n46 source.n45 42.0366
R180 source.n44 source.n43 42.0366
R181 source.n42 source.n41 42.0366
R182 source.n40 source.n39 42.0366
R183 source.n38 source.n37 42.0366
R184 source.n34 source.n33 42.0366
R185 source.n32 source.n31 42.0366
R186 source.n30 source.n29 42.0366
R187 source.n28 source.n27 42.0366
R188 source.n26 source.n25 42.0366
R189 source.n2 source.n1 42.0366
R190 source.n4 source.n3 42.0366
R191 source.n6 source.n5 42.0366
R192 source.n8 source.n7 42.0366
R193 source.n10 source.n9 42.0366
R194 source.n14 source.n13 42.0366
R195 source.n16 source.n15 42.0366
R196 source.n18 source.n17 42.0366
R197 source.n20 source.n19 42.0366
R198 source.n22 source.n21 42.0366
R199 source.n24 source.n23 31.6966
R200 source.n48 source.n0 26.1535
R201 source.n48 source.n47 5.5436
R202 source.n45 source.t27 1.2005
R203 source.n45 source.t47 1.2005
R204 source.n43 source.t45 1.2005
R205 source.n43 source.t38 1.2005
R206 source.n41 source.t29 1.2005
R207 source.n41 source.t24 1.2005
R208 source.n39 source.t46 1.2005
R209 source.n39 source.t39 1.2005
R210 source.n37 source.t33 1.2005
R211 source.n37 source.t25 1.2005
R212 source.n33 source.t5 1.2005
R213 source.n33 source.t19 1.2005
R214 source.n31 source.t17 1.2005
R215 source.n31 source.t0 1.2005
R216 source.n29 source.t10 1.2005
R217 source.n29 source.t6 1.2005
R218 source.n27 source.t1 1.2005
R219 source.n27 source.t7 1.2005
R220 source.n25 source.t2 1.2005
R221 source.n25 source.t22 1.2005
R222 source.n1 source.t23 1.2005
R223 source.n1 source.t16 1.2005
R224 source.n3 source.t20 1.2005
R225 source.n3 source.t8 1.2005
R226 source.n5 source.t13 1.2005
R227 source.n5 source.t12 1.2005
R228 source.n7 source.t9 1.2005
R229 source.n7 source.t3 1.2005
R230 source.n9 source.t18 1.2005
R231 source.n9 source.t4 1.2005
R232 source.n13 source.t35 1.2005
R233 source.n13 source.t43 1.2005
R234 source.n15 source.t40 1.2005
R235 source.n15 source.t37 1.2005
R236 source.n17 source.t34 1.2005
R237 source.n17 source.t30 1.2005
R238 source.n19 source.t36 1.2005
R239 source.n19 source.t32 1.2005
R240 source.n21 source.t28 1.2005
R241 source.n21 source.t26 1.2005
R242 source.n23 source.n22 0.560845
R243 source.n22 source.n20 0.560845
R244 source.n20 source.n18 0.560845
R245 source.n18 source.n16 0.560845
R246 source.n16 source.n14 0.560845
R247 source.n14 source.n12 0.560845
R248 source.n11 source.n10 0.560845
R249 source.n10 source.n8 0.560845
R250 source.n8 source.n6 0.560845
R251 source.n6 source.n4 0.560845
R252 source.n4 source.n2 0.560845
R253 source.n2 source.n0 0.560845
R254 source.n26 source.n24 0.560845
R255 source.n28 source.n26 0.560845
R256 source.n30 source.n28 0.560845
R257 source.n32 source.n30 0.560845
R258 source.n34 source.n32 0.560845
R259 source.n35 source.n34 0.560845
R260 source.n38 source.n36 0.560845
R261 source.n40 source.n38 0.560845
R262 source.n42 source.n40 0.560845
R263 source.n44 source.n42 0.560845
R264 source.n46 source.n44 0.560845
R265 source.n47 source.n46 0.560845
R266 source.n12 source.n11 0.470328
R267 source.n36 source.n35 0.470328
R268 source source.n48 0.188
R269 plus.n6 plus.t12 4273
R270 plus.n35 plus.t22 4273
R271 plus.n45 plus.t9 4273
R272 plus.n72 plus.t6 4273
R273 plus.n7 plus.t21 4225.53
R274 plus.n8 plus.t18 4225.53
R275 plus.n14 plus.t14 4225.53
R276 plus.n16 plus.t23 4225.53
R277 plus.n17 plus.t20 4225.53
R278 plus.n23 plus.t17 4225.53
R279 plus.n25 plus.t11 4225.53
R280 plus.n26 plus.t19 4225.53
R281 plus.n32 plus.t16 4225.53
R282 plus.n34 plus.t13 4225.53
R283 plus.n47 plus.t15 4225.53
R284 plus.n46 plus.t3 4225.53
R285 plus.n53 plus.t7 4225.53
R286 plus.n55 plus.t10 4225.53
R287 plus.n43 plus.t1 4225.53
R288 plus.n61 plus.t5 4225.53
R289 plus.n63 plus.t4 4225.53
R290 plus.n40 plus.t8 4225.53
R291 plus.n69 plus.t0 4225.53
R292 plus.n71 plus.t2 4225.53
R293 plus.n10 plus.n6 161.489
R294 plus.n49 plus.n45 161.489
R295 plus.n10 plus.n9 161.3
R296 plus.n11 plus.n5 161.3
R297 plus.n13 plus.n12 161.3
R298 plus.n15 plus.n4 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n3 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n24 plus.n2 161.3
R303 plus.n28 plus.n27 161.3
R304 plus.n29 plus.n1 161.3
R305 plus.n31 plus.n30 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n49 plus.n48 161.3
R309 plus.n50 plus.n44 161.3
R310 plus.n52 plus.n51 161.3
R311 plus.n54 plus.n42 161.3
R312 plus.n57 plus.n56 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n39 161.3
R316 plus.n65 plus.n64 161.3
R317 plus.n66 plus.n38 161.3
R318 plus.n68 plus.n67 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n13 plus.n5 73.0308
R322 plus.n22 plus.n3 73.0308
R323 plus.n31 plus.n1 73.0308
R324 plus.n68 plus.n38 73.0308
R325 plus.n60 plus.n41 73.0308
R326 plus.n52 plus.n44 73.0308
R327 plus.n9 plus.n8 69.3793
R328 plus.n33 plus.n32 69.3793
R329 plus.n70 plus.n69 69.3793
R330 plus.n48 plus.n46 69.3793
R331 plus.n18 plus.n17 62.0763
R332 plus.n24 plus.n23 62.0763
R333 plus.n62 plus.n61 62.0763
R334 plus.n56 plus.n43 62.0763
R335 plus.n15 plus.n14 54.7732
R336 plus.n27 plus.n26 54.7732
R337 plus.n64 plus.n40 54.7732
R338 plus.n54 plus.n53 54.7732
R339 plus.n7 plus.n6 47.4702
R340 plus.n35 plus.n34 47.4702
R341 plus.n72 plus.n71 47.4702
R342 plus.n47 plus.n45 47.4702
R343 plus.n16 plus.n15 40.1672
R344 plus.n27 plus.n25 40.1672
R345 plus.n64 plus.n63 40.1672
R346 plus.n55 plus.n54 40.1672
R347 plus plus.n73 37.0634
R348 plus.n18 plus.n16 32.8641
R349 plus.n25 plus.n24 32.8641
R350 plus.n63 plus.n62 32.8641
R351 plus.n56 plus.n55 32.8641
R352 plus.n9 plus.n7 25.5611
R353 plus.n34 plus.n33 25.5611
R354 plus.n71 plus.n70 25.5611
R355 plus.n48 plus.n47 25.5611
R356 plus.n14 plus.n13 18.2581
R357 plus.n26 plus.n1 18.2581
R358 plus.n40 plus.n38 18.2581
R359 plus.n53 plus.n52 18.2581
R360 plus plus.n36 17.0914
R361 plus.n17 plus.n3 10.955
R362 plus.n23 plus.n22 10.955
R363 plus.n61 plus.n60 10.955
R364 plus.n43 plus.n41 10.955
R365 plus.n8 plus.n5 3.65202
R366 plus.n32 plus.n31 3.65202
R367 plus.n69 plus.n68 3.65202
R368 plus.n46 plus.n44 3.65202
R369 plus.n11 plus.n10 0.189894
R370 plus.n12 plus.n11 0.189894
R371 plus.n12 plus.n4 0.189894
R372 plus.n19 plus.n4 0.189894
R373 plus.n20 plus.n19 0.189894
R374 plus.n21 plus.n20 0.189894
R375 plus.n21 plus.n2 0.189894
R376 plus.n28 plus.n2 0.189894
R377 plus.n29 plus.n28 0.189894
R378 plus.n30 plus.n29 0.189894
R379 plus.n30 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n67 plus.n37 0.189894
R383 plus.n67 plus.n66 0.189894
R384 plus.n66 plus.n65 0.189894
R385 plus.n65 plus.n39 0.189894
R386 plus.n59 plus.n39 0.189894
R387 plus.n59 plus.n58 0.189894
R388 plus.n58 plus.n57 0.189894
R389 plus.n57 plus.n42 0.189894
R390 plus.n51 plus.n42 0.189894
R391 plus.n51 plus.n50 0.189894
R392 plus.n50 plus.n49 0.189894
R393 drain_left.n7 drain_left.n5 59.2758
R394 drain_left.n2 drain_left.n0 59.2758
R395 drain_left.n13 drain_left.n11 59.2758
R396 drain_left.n7 drain_left.n6 58.7154
R397 drain_left.n9 drain_left.n8 58.7154
R398 drain_left.n4 drain_left.n3 58.7154
R399 drain_left.n2 drain_left.n1 58.7154
R400 drain_left.n19 drain_left.n18 58.7154
R401 drain_left.n17 drain_left.n16 58.7154
R402 drain_left.n15 drain_left.n14 58.7154
R403 drain_left.n13 drain_left.n12 58.7154
R404 drain_left.n21 drain_left.n20 58.7153
R405 drain_left drain_left.n10 42.5388
R406 drain_left drain_left.n21 6.21356
R407 drain_left.n5 drain_left.t8 1.2005
R408 drain_left.n5 drain_left.t14 1.2005
R409 drain_left.n6 drain_left.t16 1.2005
R410 drain_left.n6 drain_left.t20 1.2005
R411 drain_left.n8 drain_left.t22 1.2005
R412 drain_left.n8 drain_left.t13 1.2005
R413 drain_left.n3 drain_left.t19 1.2005
R414 drain_left.n3 drain_left.t18 1.2005
R415 drain_left.n1 drain_left.t23 1.2005
R416 drain_left.n1 drain_left.t15 1.2005
R417 drain_left.n0 drain_left.t17 1.2005
R418 drain_left.n0 drain_left.t21 1.2005
R419 drain_left.n20 drain_left.t10 1.2005
R420 drain_left.n20 drain_left.t1 1.2005
R421 drain_left.n18 drain_left.t4 1.2005
R422 drain_left.n18 drain_left.t7 1.2005
R423 drain_left.n16 drain_left.t6 1.2005
R424 drain_left.n16 drain_left.t12 1.2005
R425 drain_left.n14 drain_left.t0 1.2005
R426 drain_left.n14 drain_left.t3 1.2005
R427 drain_left.n12 drain_left.t5 1.2005
R428 drain_left.n12 drain_left.t9 1.2005
R429 drain_left.n11 drain_left.t11 1.2005
R430 drain_left.n11 drain_left.t2 1.2005
R431 drain_left.n9 drain_left.n7 0.560845
R432 drain_left.n4 drain_left.n2 0.560845
R433 drain_left.n15 drain_left.n13 0.560845
R434 drain_left.n17 drain_left.n15 0.560845
R435 drain_left.n19 drain_left.n17 0.560845
R436 drain_left.n21 drain_left.n19 0.560845
R437 drain_left.n10 drain_left.n9 0.225326
R438 drain_left.n10 drain_left.n4 0.225326
C0 drain_left source 90.293106f
C1 minus drain_left 0.171476f
C2 plus drain_left 9.70437f
C3 drain_right drain_left 1.29455f
C4 minus source 8.42116f
C5 plus source 8.435201f
C6 drain_right source 90.29379f
C7 minus plus 8.54892f
C8 drain_right minus 9.46659f
C9 drain_right plus 0.392113f
C10 drain_right a_n2406_n5888# 9.20126f
C11 drain_left a_n2406_n5888# 9.546061f
C12 source a_n2406_n5888# 15.981501f
C13 minus a_n2406_n5888# 9.790675f
C14 plus a_n2406_n5888# 12.86996f
C15 drain_left.t17 a_n2406_n5888# 0.845245f
C16 drain_left.t21 a_n2406_n5888# 0.845245f
C17 drain_left.n0 a_n2406_n5888# 5.71939f
C18 drain_left.t23 a_n2406_n5888# 0.845245f
C19 drain_left.t15 a_n2406_n5888# 0.845245f
C20 drain_left.n1 a_n2406_n5888# 5.71607f
C21 drain_left.n2 a_n2406_n5888# 0.689372f
C22 drain_left.t19 a_n2406_n5888# 0.845245f
C23 drain_left.t18 a_n2406_n5888# 0.845245f
C24 drain_left.n3 a_n2406_n5888# 5.71607f
C25 drain_left.n4 a_n2406_n5888# 0.313046f
C26 drain_left.t8 a_n2406_n5888# 0.845245f
C27 drain_left.t14 a_n2406_n5888# 0.845245f
C28 drain_left.n5 a_n2406_n5888# 5.71939f
C29 drain_left.t16 a_n2406_n5888# 0.845245f
C30 drain_left.t20 a_n2406_n5888# 0.845245f
C31 drain_left.n6 a_n2406_n5888# 5.71607f
C32 drain_left.n7 a_n2406_n5888# 0.689372f
C33 drain_left.t22 a_n2406_n5888# 0.845245f
C34 drain_left.t13 a_n2406_n5888# 0.845245f
C35 drain_left.n8 a_n2406_n5888# 5.71607f
C36 drain_left.n9 a_n2406_n5888# 0.313046f
C37 drain_left.n10 a_n2406_n5888# 2.47327f
C38 drain_left.t11 a_n2406_n5888# 0.845245f
C39 drain_left.t2 a_n2406_n5888# 0.845245f
C40 drain_left.n11 a_n2406_n5888# 5.71939f
C41 drain_left.t5 a_n2406_n5888# 0.845245f
C42 drain_left.t9 a_n2406_n5888# 0.845245f
C43 drain_left.n12 a_n2406_n5888# 5.71607f
C44 drain_left.n13 a_n2406_n5888# 0.689369f
C45 drain_left.t0 a_n2406_n5888# 0.845245f
C46 drain_left.t3 a_n2406_n5888# 0.845245f
C47 drain_left.n14 a_n2406_n5888# 5.71607f
C48 drain_left.n15 a_n2406_n5888# 0.340662f
C49 drain_left.t6 a_n2406_n5888# 0.845245f
C50 drain_left.t12 a_n2406_n5888# 0.845245f
C51 drain_left.n16 a_n2406_n5888# 5.71607f
C52 drain_left.n17 a_n2406_n5888# 0.340662f
C53 drain_left.t4 a_n2406_n5888# 0.845245f
C54 drain_left.t7 a_n2406_n5888# 0.845245f
C55 drain_left.n18 a_n2406_n5888# 5.71607f
C56 drain_left.n19 a_n2406_n5888# 0.340662f
C57 drain_left.t10 a_n2406_n5888# 0.845245f
C58 drain_left.t1 a_n2406_n5888# 0.845245f
C59 drain_left.n20 a_n2406_n5888# 5.71605f
C60 drain_left.n21 a_n2406_n5888# 0.576491f
C61 plus.n0 a_n2406_n5888# 0.052259f
C62 plus.t13 a_n2406_n5888# 0.551398f
C63 plus.t16 a_n2406_n5888# 0.551398f
C64 plus.n1 a_n2406_n5888# 0.021363f
C65 plus.n2 a_n2406_n5888# 0.052259f
C66 plus.t11 a_n2406_n5888# 0.551398f
C67 plus.t17 a_n2406_n5888# 0.551398f
C68 plus.n3 a_n2406_n5888# 0.019753f
C69 plus.n4 a_n2406_n5888# 0.052259f
C70 plus.t23 a_n2406_n5888# 0.551398f
C71 plus.t14 a_n2406_n5888# 0.551398f
C72 plus.n5 a_n2406_n5888# 0.018142f
C73 plus.t12 a_n2406_n5888# 0.553707f
C74 plus.n6 a_n2406_n5888# 0.227823f
C75 plus.t21 a_n2406_n5888# 0.551398f
C76 plus.n7 a_n2406_n5888# 0.208696f
C77 plus.t18 a_n2406_n5888# 0.551398f
C78 plus.n8 a_n2406_n5888# 0.208696f
C79 plus.n9 a_n2406_n5888# 0.022169f
C80 plus.n10 a_n2406_n5888# 0.114111f
C81 plus.n11 a_n2406_n5888# 0.052259f
C82 plus.n12 a_n2406_n5888# 0.052259f
C83 plus.n13 a_n2406_n5888# 0.021363f
C84 plus.n14 a_n2406_n5888# 0.208696f
C85 plus.n15 a_n2406_n5888# 0.022169f
C86 plus.n16 a_n2406_n5888# 0.208696f
C87 plus.t20 a_n2406_n5888# 0.551398f
C88 plus.n17 a_n2406_n5888# 0.208696f
C89 plus.n18 a_n2406_n5888# 0.022169f
C90 plus.n19 a_n2406_n5888# 0.052259f
C91 plus.n20 a_n2406_n5888# 0.052259f
C92 plus.n21 a_n2406_n5888# 0.052259f
C93 plus.n22 a_n2406_n5888# 0.019753f
C94 plus.n23 a_n2406_n5888# 0.208696f
C95 plus.n24 a_n2406_n5888# 0.022169f
C96 plus.n25 a_n2406_n5888# 0.208696f
C97 plus.t19 a_n2406_n5888# 0.551398f
C98 plus.n26 a_n2406_n5888# 0.208696f
C99 plus.n27 a_n2406_n5888# 0.022169f
C100 plus.n28 a_n2406_n5888# 0.052259f
C101 plus.n29 a_n2406_n5888# 0.052259f
C102 plus.n30 a_n2406_n5888# 0.052259f
C103 plus.n31 a_n2406_n5888# 0.018142f
C104 plus.n32 a_n2406_n5888# 0.208696f
C105 plus.n33 a_n2406_n5888# 0.022169f
C106 plus.n34 a_n2406_n5888# 0.208696f
C107 plus.t22 a_n2406_n5888# 0.553707f
C108 plus.n35 a_n2406_n5888# 0.22775f
C109 plus.n36 a_n2406_n5888# 0.935581f
C110 plus.n37 a_n2406_n5888# 0.052259f
C111 plus.t6 a_n2406_n5888# 0.553707f
C112 plus.t2 a_n2406_n5888# 0.551398f
C113 plus.t0 a_n2406_n5888# 0.551398f
C114 plus.n38 a_n2406_n5888# 0.021363f
C115 plus.n39 a_n2406_n5888# 0.052259f
C116 plus.t8 a_n2406_n5888# 0.551398f
C117 plus.n40 a_n2406_n5888# 0.208696f
C118 plus.t4 a_n2406_n5888# 0.551398f
C119 plus.t5 a_n2406_n5888# 0.551398f
C120 plus.n41 a_n2406_n5888# 0.019753f
C121 plus.n42 a_n2406_n5888# 0.052259f
C122 plus.t1 a_n2406_n5888# 0.551398f
C123 plus.n43 a_n2406_n5888# 0.208696f
C124 plus.t10 a_n2406_n5888# 0.551398f
C125 plus.t7 a_n2406_n5888# 0.551398f
C126 plus.n44 a_n2406_n5888# 0.018142f
C127 plus.t9 a_n2406_n5888# 0.553707f
C128 plus.n45 a_n2406_n5888# 0.227823f
C129 plus.t3 a_n2406_n5888# 0.551398f
C130 plus.n46 a_n2406_n5888# 0.208696f
C131 plus.t15 a_n2406_n5888# 0.551398f
C132 plus.n47 a_n2406_n5888# 0.208696f
C133 plus.n48 a_n2406_n5888# 0.022169f
C134 plus.n49 a_n2406_n5888# 0.114111f
C135 plus.n50 a_n2406_n5888# 0.052259f
C136 plus.n51 a_n2406_n5888# 0.052259f
C137 plus.n52 a_n2406_n5888# 0.021363f
C138 plus.n53 a_n2406_n5888# 0.208696f
C139 plus.n54 a_n2406_n5888# 0.022169f
C140 plus.n55 a_n2406_n5888# 0.208696f
C141 plus.n56 a_n2406_n5888# 0.022169f
C142 plus.n57 a_n2406_n5888# 0.052259f
C143 plus.n58 a_n2406_n5888# 0.052259f
C144 plus.n59 a_n2406_n5888# 0.052259f
C145 plus.n60 a_n2406_n5888# 0.019753f
C146 plus.n61 a_n2406_n5888# 0.208696f
C147 plus.n62 a_n2406_n5888# 0.022169f
C148 plus.n63 a_n2406_n5888# 0.208696f
C149 plus.n64 a_n2406_n5888# 0.022169f
C150 plus.n65 a_n2406_n5888# 0.052259f
C151 plus.n66 a_n2406_n5888# 0.052259f
C152 plus.n67 a_n2406_n5888# 0.052259f
C153 plus.n68 a_n2406_n5888# 0.018142f
C154 plus.n69 a_n2406_n5888# 0.208696f
C155 plus.n70 a_n2406_n5888# 0.022169f
C156 plus.n71 a_n2406_n5888# 0.208696f
C157 plus.n72 a_n2406_n5888# 0.22775f
C158 plus.n73 a_n2406_n5888# 2.1738f
C159 source.t21 a_n2406_n5888# 6.114759f
C160 source.n0 a_n2406_n5888# 2.3398f
C161 source.t23 a_n2406_n5888# 0.741524f
C162 source.t16 a_n2406_n5888# 0.741524f
C163 source.n1 a_n2406_n5888# 4.93342f
C164 source.n2 a_n2406_n5888# 0.3464f
C165 source.t20 a_n2406_n5888# 0.741524f
C166 source.t8 a_n2406_n5888# 0.741524f
C167 source.n3 a_n2406_n5888# 4.93342f
C168 source.n4 a_n2406_n5888# 0.3464f
C169 source.t13 a_n2406_n5888# 0.741524f
C170 source.t12 a_n2406_n5888# 0.741524f
C171 source.n5 a_n2406_n5888# 4.93342f
C172 source.n6 a_n2406_n5888# 0.3464f
C173 source.t9 a_n2406_n5888# 0.741524f
C174 source.t3 a_n2406_n5888# 0.741524f
C175 source.n7 a_n2406_n5888# 4.93342f
C176 source.n8 a_n2406_n5888# 0.3464f
C177 source.t18 a_n2406_n5888# 0.741524f
C178 source.t4 a_n2406_n5888# 0.741524f
C179 source.n9 a_n2406_n5888# 4.93342f
C180 source.n10 a_n2406_n5888# 0.3464f
C181 source.t11 a_n2406_n5888# 6.11478f
C182 source.n11 a_n2406_n5888# 0.492565f
C183 source.t41 a_n2406_n5888# 6.11478f
C184 source.n12 a_n2406_n5888# 0.492565f
C185 source.t35 a_n2406_n5888# 0.741524f
C186 source.t43 a_n2406_n5888# 0.741524f
C187 source.n13 a_n2406_n5888# 4.93342f
C188 source.n14 a_n2406_n5888# 0.3464f
C189 source.t40 a_n2406_n5888# 0.741524f
C190 source.t37 a_n2406_n5888# 0.741524f
C191 source.n15 a_n2406_n5888# 4.93342f
C192 source.n16 a_n2406_n5888# 0.3464f
C193 source.t34 a_n2406_n5888# 0.741524f
C194 source.t30 a_n2406_n5888# 0.741524f
C195 source.n17 a_n2406_n5888# 4.93342f
C196 source.n18 a_n2406_n5888# 0.3464f
C197 source.t36 a_n2406_n5888# 0.741524f
C198 source.t32 a_n2406_n5888# 0.741524f
C199 source.n19 a_n2406_n5888# 4.93342f
C200 source.n20 a_n2406_n5888# 0.3464f
C201 source.t28 a_n2406_n5888# 0.741524f
C202 source.t26 a_n2406_n5888# 0.741524f
C203 source.n21 a_n2406_n5888# 4.93342f
C204 source.n22 a_n2406_n5888# 0.3464f
C205 source.t31 a_n2406_n5888# 6.11478f
C206 source.n23 a_n2406_n5888# 2.79869f
C207 source.t14 a_n2406_n5888# 6.114759f
C208 source.n24 a_n2406_n5888# 2.79871f
C209 source.t2 a_n2406_n5888# 0.741524f
C210 source.t22 a_n2406_n5888# 0.741524f
C211 source.n25 a_n2406_n5888# 4.93342f
C212 source.n26 a_n2406_n5888# 0.346402f
C213 source.t1 a_n2406_n5888# 0.741524f
C214 source.t7 a_n2406_n5888# 0.741524f
C215 source.n27 a_n2406_n5888# 4.93342f
C216 source.n28 a_n2406_n5888# 0.346402f
C217 source.t10 a_n2406_n5888# 0.741524f
C218 source.t6 a_n2406_n5888# 0.741524f
C219 source.n29 a_n2406_n5888# 4.93342f
C220 source.n30 a_n2406_n5888# 0.346402f
C221 source.t17 a_n2406_n5888# 0.741524f
C222 source.t0 a_n2406_n5888# 0.741524f
C223 source.n31 a_n2406_n5888# 4.93342f
C224 source.n32 a_n2406_n5888# 0.346402f
C225 source.t5 a_n2406_n5888# 0.741524f
C226 source.t19 a_n2406_n5888# 0.741524f
C227 source.n33 a_n2406_n5888# 4.93342f
C228 source.n34 a_n2406_n5888# 0.346402f
C229 source.t15 a_n2406_n5888# 6.114759f
C230 source.n35 a_n2406_n5888# 0.492581f
C231 source.t44 a_n2406_n5888# 6.114759f
C232 source.n36 a_n2406_n5888# 0.492581f
C233 source.t33 a_n2406_n5888# 0.741524f
C234 source.t25 a_n2406_n5888# 0.741524f
C235 source.n37 a_n2406_n5888# 4.93342f
C236 source.n38 a_n2406_n5888# 0.346402f
C237 source.t46 a_n2406_n5888# 0.741524f
C238 source.t39 a_n2406_n5888# 0.741524f
C239 source.n39 a_n2406_n5888# 4.93342f
C240 source.n40 a_n2406_n5888# 0.346402f
C241 source.t29 a_n2406_n5888# 0.741524f
C242 source.t24 a_n2406_n5888# 0.741524f
C243 source.n41 a_n2406_n5888# 4.93342f
C244 source.n42 a_n2406_n5888# 0.346402f
C245 source.t45 a_n2406_n5888# 0.741524f
C246 source.t38 a_n2406_n5888# 0.741524f
C247 source.n43 a_n2406_n5888# 4.93342f
C248 source.n44 a_n2406_n5888# 0.346402f
C249 source.t27 a_n2406_n5888# 0.741524f
C250 source.t47 a_n2406_n5888# 0.741524f
C251 source.n45 a_n2406_n5888# 4.93342f
C252 source.n46 a_n2406_n5888# 0.346402f
C253 source.t42 a_n2406_n5888# 6.114759f
C254 source.n47 a_n2406_n5888# 0.633522f
C255 source.n48 a_n2406_n5888# 2.64172f
C256 drain_right.t5 a_n2406_n5888# 0.844488f
C257 drain_right.t6 a_n2406_n5888# 0.844488f
C258 drain_right.n0 a_n2406_n5888# 5.71427f
C259 drain_right.t16 a_n2406_n5888# 0.844488f
C260 drain_right.t1 a_n2406_n5888# 0.844488f
C261 drain_right.n1 a_n2406_n5888# 5.71094f
C262 drain_right.n2 a_n2406_n5888# 0.688754f
C263 drain_right.t18 a_n2406_n5888# 0.844488f
C264 drain_right.t23 a_n2406_n5888# 0.844488f
C265 drain_right.n3 a_n2406_n5888# 5.71094f
C266 drain_right.n4 a_n2406_n5888# 0.312766f
C267 drain_right.t2 a_n2406_n5888# 0.844488f
C268 drain_right.t3 a_n2406_n5888# 0.844488f
C269 drain_right.n5 a_n2406_n5888# 5.71427f
C270 drain_right.t11 a_n2406_n5888# 0.844488f
C271 drain_right.t21 a_n2406_n5888# 0.844488f
C272 drain_right.n6 a_n2406_n5888# 5.71094f
C273 drain_right.n7 a_n2406_n5888# 0.688754f
C274 drain_right.t15 a_n2406_n5888# 0.844488f
C275 drain_right.t0 a_n2406_n5888# 0.844488f
C276 drain_right.n8 a_n2406_n5888# 5.71094f
C277 drain_right.n9 a_n2406_n5888# 0.312766f
C278 drain_right.n10 a_n2406_n5888# 2.41298f
C279 drain_right.t4 a_n2406_n5888# 0.844488f
C280 drain_right.t20 a_n2406_n5888# 0.844488f
C281 drain_right.n11 a_n2406_n5888# 5.71426f
C282 drain_right.t10 a_n2406_n5888# 0.844488f
C283 drain_right.t8 a_n2406_n5888# 0.844488f
C284 drain_right.n12 a_n2406_n5888# 5.71094f
C285 drain_right.n13 a_n2406_n5888# 0.688764f
C286 drain_right.t12 a_n2406_n5888# 0.844488f
C287 drain_right.t19 a_n2406_n5888# 0.844488f
C288 drain_right.n14 a_n2406_n5888# 5.71094f
C289 drain_right.n15 a_n2406_n5888# 0.340356f
C290 drain_right.t14 a_n2406_n5888# 0.844488f
C291 drain_right.t7 a_n2406_n5888# 0.844488f
C292 drain_right.n16 a_n2406_n5888# 5.71094f
C293 drain_right.n17 a_n2406_n5888# 0.340356f
C294 drain_right.t17 a_n2406_n5888# 0.844488f
C295 drain_right.t9 a_n2406_n5888# 0.844488f
C296 drain_right.n18 a_n2406_n5888# 5.71094f
C297 drain_right.n19 a_n2406_n5888# 0.340356f
C298 drain_right.t13 a_n2406_n5888# 0.844488f
C299 drain_right.t22 a_n2406_n5888# 0.844488f
C300 drain_right.n20 a_n2406_n5888# 5.71094f
C301 drain_right.n21 a_n2406_n5888# 0.575962f
C302 minus.n0 a_n2406_n5888# 0.051661f
C303 minus.t16 a_n2406_n5888# 0.54737f
C304 minus.t19 a_n2406_n5888# 0.545086f
C305 minus.t21 a_n2406_n5888# 0.545086f
C306 minus.n1 a_n2406_n5888# 0.021119f
C307 minus.n2 a_n2406_n5888# 0.051661f
C308 minus.t11 a_n2406_n5888# 0.545086f
C309 minus.n3 a_n2406_n5888# 0.206308f
C310 minus.t15 a_n2406_n5888# 0.545086f
C311 minus.t13 a_n2406_n5888# 0.545086f
C312 minus.n4 a_n2406_n5888# 0.019526f
C313 minus.n5 a_n2406_n5888# 0.051661f
C314 minus.t17 a_n2406_n5888# 0.545086f
C315 minus.n6 a_n2406_n5888# 0.206308f
C316 minus.t7 a_n2406_n5888# 0.545086f
C317 minus.t10 a_n2406_n5888# 0.545086f
C318 minus.n7 a_n2406_n5888# 0.017934f
C319 minus.t6 a_n2406_n5888# 0.54737f
C320 minus.n8 a_n2406_n5888# 0.225215f
C321 minus.t12 a_n2406_n5888# 0.545086f
C322 minus.n9 a_n2406_n5888# 0.206308f
C323 minus.t4 a_n2406_n5888# 0.545086f
C324 minus.n10 a_n2406_n5888# 0.206308f
C325 minus.n11 a_n2406_n5888# 0.021915f
C326 minus.n12 a_n2406_n5888# 0.112805f
C327 minus.n13 a_n2406_n5888# 0.051661f
C328 minus.n14 a_n2406_n5888# 0.051661f
C329 minus.n15 a_n2406_n5888# 0.021119f
C330 minus.n16 a_n2406_n5888# 0.206308f
C331 minus.n17 a_n2406_n5888# 0.021915f
C332 minus.n18 a_n2406_n5888# 0.206308f
C333 minus.n19 a_n2406_n5888# 0.021915f
C334 minus.n20 a_n2406_n5888# 0.051661f
C335 minus.n21 a_n2406_n5888# 0.051661f
C336 minus.n22 a_n2406_n5888# 0.051661f
C337 minus.n23 a_n2406_n5888# 0.019526f
C338 minus.n24 a_n2406_n5888# 0.206308f
C339 minus.n25 a_n2406_n5888# 0.021915f
C340 minus.n26 a_n2406_n5888# 0.206308f
C341 minus.n27 a_n2406_n5888# 0.021915f
C342 minus.n28 a_n2406_n5888# 0.051661f
C343 minus.n29 a_n2406_n5888# 0.051661f
C344 minus.n30 a_n2406_n5888# 0.051661f
C345 minus.n31 a_n2406_n5888# 0.017934f
C346 minus.n32 a_n2406_n5888# 0.206308f
C347 minus.n33 a_n2406_n5888# 0.021915f
C348 minus.n34 a_n2406_n5888# 0.206308f
C349 minus.n35 a_n2406_n5888# 0.225143f
C350 minus.n36 a_n2406_n5888# 2.78139f
C351 minus.n37 a_n2406_n5888# 0.051661f
C352 minus.t0 a_n2406_n5888# 0.545086f
C353 minus.t20 a_n2406_n5888# 0.545086f
C354 minus.n38 a_n2406_n5888# 0.021119f
C355 minus.n39 a_n2406_n5888# 0.051661f
C356 minus.t2 a_n2406_n5888# 0.545086f
C357 minus.t23 a_n2406_n5888# 0.545086f
C358 minus.n40 a_n2406_n5888# 0.019526f
C359 minus.n41 a_n2406_n5888# 0.051661f
C360 minus.t8 a_n2406_n5888# 0.545086f
C361 minus.t1 a_n2406_n5888# 0.545086f
C362 minus.n42 a_n2406_n5888# 0.017934f
C363 minus.t3 a_n2406_n5888# 0.54737f
C364 minus.n43 a_n2406_n5888# 0.225215f
C365 minus.t14 a_n2406_n5888# 0.545086f
C366 minus.n44 a_n2406_n5888# 0.206308f
C367 minus.t22 a_n2406_n5888# 0.545086f
C368 minus.n45 a_n2406_n5888# 0.206308f
C369 minus.n46 a_n2406_n5888# 0.021915f
C370 minus.n47 a_n2406_n5888# 0.112805f
C371 minus.n48 a_n2406_n5888# 0.051661f
C372 minus.n49 a_n2406_n5888# 0.051661f
C373 minus.n50 a_n2406_n5888# 0.021119f
C374 minus.n51 a_n2406_n5888# 0.206308f
C375 minus.n52 a_n2406_n5888# 0.021915f
C376 minus.n53 a_n2406_n5888# 0.206308f
C377 minus.t18 a_n2406_n5888# 0.545086f
C378 minus.n54 a_n2406_n5888# 0.206308f
C379 minus.n55 a_n2406_n5888# 0.021915f
C380 minus.n56 a_n2406_n5888# 0.051661f
C381 minus.n57 a_n2406_n5888# 0.051661f
C382 minus.n58 a_n2406_n5888# 0.051661f
C383 minus.n59 a_n2406_n5888# 0.019526f
C384 minus.n60 a_n2406_n5888# 0.206308f
C385 minus.n61 a_n2406_n5888# 0.021915f
C386 minus.n62 a_n2406_n5888# 0.206308f
C387 minus.t9 a_n2406_n5888# 0.545086f
C388 minus.n63 a_n2406_n5888# 0.206308f
C389 minus.n64 a_n2406_n5888# 0.021915f
C390 minus.n65 a_n2406_n5888# 0.051661f
C391 minus.n66 a_n2406_n5888# 0.051661f
C392 minus.n67 a_n2406_n5888# 0.051661f
C393 minus.n68 a_n2406_n5888# 0.017934f
C394 minus.n69 a_n2406_n5888# 0.206308f
C395 minus.n70 a_n2406_n5888# 0.021915f
C396 minus.n71 a_n2406_n5888# 0.206308f
C397 minus.t5 a_n2406_n5888# 0.54737f
C398 minus.n72 a_n2406_n5888# 0.225143f
C399 minus.n73 a_n2406_n5888# 0.340568f
C400 minus.n74 a_n2406_n5888# 3.2666f
.ends

