* NGSPICE file created from diffpair607.ext - technology: sky130A

.subckt diffpair607 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t23 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t18 plus.t1 drain_left.t14 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 drain_right.t15 minus.t0 source.t0 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X3 a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X4 source.t17 plus.t2 drain_left.t13 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X5 source.t9 minus.t1 drain_right.t14 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t16 plus.t3 drain_left.t12 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X7 drain_left.t11 plus.t4 source.t26 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 source.t21 plus.t5 drain_left.t10 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X9 drain_right.t13 minus.t2 source.t3 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 source.t10 minus.t3 drain_right.t12 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X11 drain_right.t11 minus.t4 source.t14 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X12 a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X13 drain_right.t10 minus.t5 source.t1 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X14 source.t13 minus.t6 drain_right.t9 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 drain_left.t9 plus.t6 source.t30 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X16 drain_left.t8 plus.t7 source.t29 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X17 drain_left.t7 plus.t8 source.t28 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X18 source.t20 plus.t9 drain_left.t6 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 source.t2 minus.t7 drain_right.t8 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X20 drain_right.t7 minus.t8 source.t6 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X21 source.t15 minus.t9 drain_right.t6 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X22 source.t31 plus.t10 drain_left.t5 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 drain_right.t5 minus.t10 source.t8 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X24 drain_right.t4 minus.t11 source.t12 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X25 source.t5 minus.t12 drain_right.t3 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X26 a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X27 drain_left.t4 plus.t11 source.t24 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X28 a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X29 source.t7 minus.t13 drain_right.t2 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X30 drain_right.t1 minus.t14 source.t11 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X31 source.t4 minus.t15 drain_right.t0 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X32 source.t25 plus.t12 drain_left.t3 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X33 drain_left.t2 plus.t13 source.t19 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X34 source.t27 plus.t14 drain_left.t1 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X35 drain_left.t0 plus.t15 source.t22 a_n2210_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
R0 plus.n5 plus.t5 1063.55
R1 plus.n27 plus.t0 1063.55
R2 plus.n20 plus.t13 1042.57
R3 plus.n19 plus.t9 1042.57
R4 plus.n1 plus.t15 1042.57
R5 plus.n13 plus.t12 1042.57
R6 plus.n12 plus.t6 1042.57
R7 plus.n4 plus.t14 1042.57
R8 plus.n6 plus.t11 1042.57
R9 plus.n42 plus.t2 1042.57
R10 plus.n41 plus.t7 1042.57
R11 plus.n23 plus.t10 1042.57
R12 plus.n35 plus.t4 1042.57
R13 plus.n34 plus.t3 1042.57
R14 plus.n26 plus.t8 1042.57
R15 plus.n28 plus.t1 1042.57
R16 plus.n8 plus.n7 161.3
R17 plus.n9 plus.n4 161.3
R18 plus.n11 plus.n10 161.3
R19 plus.n12 plus.n3 161.3
R20 plus.n13 plus.n2 161.3
R21 plus.n15 plus.n14 161.3
R22 plus.n16 plus.n1 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n21 plus.n20 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n31 plus.n26 161.3
R28 plus.n33 plus.n32 161.3
R29 plus.n34 plus.n25 161.3
R30 plus.n35 plus.n24 161.3
R31 plus.n37 plus.n36 161.3
R32 plus.n38 plus.n23 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n41 plus.n22 161.3
R35 plus.n43 plus.n42 161.3
R36 plus.n8 plus.n5 70.4033
R37 plus.n30 plus.n27 70.4033
R38 plus.n20 plus.n19 48.2005
R39 plus.n13 plus.n12 48.2005
R40 plus.n42 plus.n41 48.2005
R41 plus.n35 plus.n34 48.2005
R42 plus.n18 plus.n1 37.246
R43 plus.n7 plus.n4 37.246
R44 plus.n40 plus.n23 37.246
R45 plus.n29 plus.n26 37.246
R46 plus.n14 plus.n1 35.7853
R47 plus.n11 plus.n4 35.7853
R48 plus.n36 plus.n23 35.7853
R49 plus.n33 plus.n26 35.7853
R50 plus plus.n43 34.4649
R51 plus.n6 plus.n5 20.9576
R52 plus.n28 plus.n27 20.9576
R53 plus plus.n21 15.2353
R54 plus.n14 plus.n13 12.4157
R55 plus.n12 plus.n11 12.4157
R56 plus.n36 plus.n35 12.4157
R57 plus.n34 plus.n33 12.4157
R58 plus.n19 plus.n18 10.955
R59 plus.n7 plus.n6 10.955
R60 plus.n41 plus.n40 10.955
R61 plus.n29 plus.n28 10.955
R62 plus.n9 plus.n8 0.189894
R63 plus.n10 plus.n9 0.189894
R64 plus.n10 plus.n3 0.189894
R65 plus.n3 plus.n2 0.189894
R66 plus.n15 plus.n2 0.189894
R67 plus.n16 plus.n15 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n21 plus.n0 0.189894
R71 plus.n43 plus.n22 0.189894
R72 plus.n39 plus.n22 0.189894
R73 plus.n39 plus.n38 0.189894
R74 plus.n38 plus.n37 0.189894
R75 plus.n37 plus.n24 0.189894
R76 plus.n25 plus.n24 0.189894
R77 plus.n32 plus.n25 0.189894
R78 plus.n32 plus.n31 0.189894
R79 plus.n31 plus.n30 0.189894
R80 source.n0 source.t19 44.1297
R81 source.n7 source.t21 44.1296
R82 source.n8 source.t12 44.1296
R83 source.n15 source.t15 44.1296
R84 source.n31 source.t6 44.1295
R85 source.n24 source.t10 44.1295
R86 source.n23 source.t23 44.1295
R87 source.n16 source.t17 44.1295
R88 source.n2 source.n1 43.1397
R89 source.n4 source.n3 43.1397
R90 source.n6 source.n5 43.1397
R91 source.n10 source.n9 43.1397
R92 source.n12 source.n11 43.1397
R93 source.n14 source.n13 43.1397
R94 source.n30 source.n29 43.1396
R95 source.n28 source.n27 43.1396
R96 source.n26 source.n25 43.1396
R97 source.n22 source.n21 43.1396
R98 source.n20 source.n19 43.1396
R99 source.n18 source.n17 43.1396
R100 source.n16 source.n15 28.0638
R101 source.n32 source.n0 22.4432
R102 source.n32 source.n31 5.62119
R103 source.n29 source.t11 0.9905
R104 source.n29 source.t7 0.9905
R105 source.n27 source.t8 0.9905
R106 source.n27 source.t13 0.9905
R107 source.n25 source.t3 0.9905
R108 source.n25 source.t5 0.9905
R109 source.n21 source.t28 0.9905
R110 source.n21 source.t18 0.9905
R111 source.n19 source.t26 0.9905
R112 source.n19 source.t16 0.9905
R113 source.n17 source.t29 0.9905
R114 source.n17 source.t31 0.9905
R115 source.n1 source.t22 0.9905
R116 source.n1 source.t20 0.9905
R117 source.n3 source.t30 0.9905
R118 source.n3 source.t25 0.9905
R119 source.n5 source.t24 0.9905
R120 source.n5 source.t27 0.9905
R121 source.n9 source.t1 0.9905
R122 source.n9 source.t9 0.9905
R123 source.n11 source.t14 0.9905
R124 source.n11 source.t4 0.9905
R125 source.n13 source.t0 0.9905
R126 source.n13 source.t2 0.9905
R127 source.n15 source.n14 0.716017
R128 source.n14 source.n12 0.716017
R129 source.n12 source.n10 0.716017
R130 source.n10 source.n8 0.716017
R131 source.n7 source.n6 0.716017
R132 source.n6 source.n4 0.716017
R133 source.n4 source.n2 0.716017
R134 source.n2 source.n0 0.716017
R135 source.n18 source.n16 0.716017
R136 source.n20 source.n18 0.716017
R137 source.n22 source.n20 0.716017
R138 source.n23 source.n22 0.716017
R139 source.n26 source.n24 0.716017
R140 source.n28 source.n26 0.716017
R141 source.n30 source.n28 0.716017
R142 source.n31 source.n30 0.716017
R143 source.n8 source.n7 0.470328
R144 source.n24 source.n23 0.470328
R145 source source.n32 0.188
R146 drain_left.n9 drain_left.n7 60.534
R147 drain_left.n5 drain_left.n3 60.5339
R148 drain_left.n2 drain_left.n0 60.5339
R149 drain_left.n13 drain_left.n12 59.8185
R150 drain_left.n11 drain_left.n10 59.8185
R151 drain_left.n9 drain_left.n8 59.8185
R152 drain_left.n5 drain_left.n4 59.8184
R153 drain_left.n2 drain_left.n1 59.8184
R154 drain_left drain_left.n6 38.0785
R155 drain_left drain_left.n13 6.36873
R156 drain_left.n3 drain_left.t14 0.9905
R157 drain_left.n3 drain_left.t15 0.9905
R158 drain_left.n4 drain_left.t12 0.9905
R159 drain_left.n4 drain_left.t7 0.9905
R160 drain_left.n1 drain_left.t5 0.9905
R161 drain_left.n1 drain_left.t11 0.9905
R162 drain_left.n0 drain_left.t13 0.9905
R163 drain_left.n0 drain_left.t8 0.9905
R164 drain_left.n12 drain_left.t6 0.9905
R165 drain_left.n12 drain_left.t2 0.9905
R166 drain_left.n10 drain_left.t3 0.9905
R167 drain_left.n10 drain_left.t0 0.9905
R168 drain_left.n8 drain_left.t1 0.9905
R169 drain_left.n8 drain_left.t9 0.9905
R170 drain_left.n7 drain_left.t10 0.9905
R171 drain_left.n7 drain_left.t4 0.9905
R172 drain_left.n11 drain_left.n9 0.716017
R173 drain_left.n13 drain_left.n11 0.716017
R174 drain_left.n6 drain_left.n5 0.302913
R175 drain_left.n6 drain_left.n2 0.302913
R176 minus.n5 minus.t11 1063.55
R177 minus.n27 minus.t3 1063.55
R178 minus.n6 minus.t1 1042.57
R179 minus.n8 minus.t5 1042.57
R180 minus.n12 minus.t15 1042.57
R181 minus.n13 minus.t4 1042.57
R182 minus.n1 minus.t7 1042.57
R183 minus.n19 minus.t0 1042.57
R184 minus.n20 minus.t9 1042.57
R185 minus.n28 minus.t2 1042.57
R186 minus.n30 minus.t12 1042.57
R187 minus.n34 minus.t10 1042.57
R188 minus.n35 minus.t6 1042.57
R189 minus.n23 minus.t14 1042.57
R190 minus.n41 minus.t13 1042.57
R191 minus.n42 minus.t8 1042.57
R192 minus.n21 minus.n20 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n1 161.3
R196 minus.n15 minus.n14 161.3
R197 minus.n13 minus.n2 161.3
R198 minus.n12 minus.n11 161.3
R199 minus.n10 minus.n3 161.3
R200 minus.n9 minus.n8 161.3
R201 minus.n7 minus.n4 161.3
R202 minus.n43 minus.n42 161.3
R203 minus.n41 minus.n22 161.3
R204 minus.n40 minus.n39 161.3
R205 minus.n38 minus.n23 161.3
R206 minus.n37 minus.n36 161.3
R207 minus.n35 minus.n24 161.3
R208 minus.n34 minus.n33 161.3
R209 minus.n32 minus.n25 161.3
R210 minus.n31 minus.n30 161.3
R211 minus.n29 minus.n26 161.3
R212 minus.n5 minus.n4 70.4033
R213 minus.n27 minus.n26 70.4033
R214 minus.n13 minus.n12 48.2005
R215 minus.n20 minus.n19 48.2005
R216 minus.n35 minus.n34 48.2005
R217 minus.n42 minus.n41 48.2005
R218 minus.n44 minus.n21 43.6141
R219 minus.n8 minus.n7 37.246
R220 minus.n18 minus.n1 37.246
R221 minus.n30 minus.n29 37.246
R222 minus.n40 minus.n23 37.246
R223 minus.n8 minus.n3 35.7853
R224 minus.n14 minus.n1 35.7853
R225 minus.n30 minus.n25 35.7853
R226 minus.n36 minus.n23 35.7853
R227 minus.n6 minus.n5 20.9576
R228 minus.n28 minus.n27 20.9576
R229 minus.n12 minus.n3 12.4157
R230 minus.n14 minus.n13 12.4157
R231 minus.n34 minus.n25 12.4157
R232 minus.n36 minus.n35 12.4157
R233 minus.n7 minus.n6 10.955
R234 minus.n19 minus.n18 10.955
R235 minus.n29 minus.n28 10.955
R236 minus.n41 minus.n40 10.955
R237 minus.n44 minus.n43 6.56111
R238 minus.n21 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n15 0.189894
R242 minus.n15 minus.n2 0.189894
R243 minus.n11 minus.n2 0.189894
R244 minus.n11 minus.n10 0.189894
R245 minus.n10 minus.n9 0.189894
R246 minus.n9 minus.n4 0.189894
R247 minus.n31 minus.n26 0.189894
R248 minus.n32 minus.n31 0.189894
R249 minus.n33 minus.n32 0.189894
R250 minus.n33 minus.n24 0.189894
R251 minus.n37 minus.n24 0.189894
R252 minus.n38 minus.n37 0.189894
R253 minus.n39 minus.n38 0.189894
R254 minus.n39 minus.n22 0.189894
R255 minus.n43 minus.n22 0.189894
R256 minus minus.n44 0.188
R257 drain_right.n9 drain_right.n7 60.534
R258 drain_right.n5 drain_right.n3 60.5339
R259 drain_right.n2 drain_right.n0 60.5339
R260 drain_right.n9 drain_right.n8 59.8185
R261 drain_right.n11 drain_right.n10 59.8185
R262 drain_right.n13 drain_right.n12 59.8185
R263 drain_right.n5 drain_right.n4 59.8184
R264 drain_right.n2 drain_right.n1 59.8184
R265 drain_right drain_right.n6 37.5253
R266 drain_right drain_right.n13 6.36873
R267 drain_right.n3 drain_right.t2 0.9905
R268 drain_right.n3 drain_right.t7 0.9905
R269 drain_right.n4 drain_right.t9 0.9905
R270 drain_right.n4 drain_right.t1 0.9905
R271 drain_right.n1 drain_right.t3 0.9905
R272 drain_right.n1 drain_right.t5 0.9905
R273 drain_right.n0 drain_right.t12 0.9905
R274 drain_right.n0 drain_right.t13 0.9905
R275 drain_right.n7 drain_right.t14 0.9905
R276 drain_right.n7 drain_right.t4 0.9905
R277 drain_right.n8 drain_right.t0 0.9905
R278 drain_right.n8 drain_right.t10 0.9905
R279 drain_right.n10 drain_right.t8 0.9905
R280 drain_right.n10 drain_right.t11 0.9905
R281 drain_right.n12 drain_right.t6 0.9905
R282 drain_right.n12 drain_right.t15 0.9905
R283 drain_right.n13 drain_right.n11 0.716017
R284 drain_right.n11 drain_right.n9 0.716017
R285 drain_right.n6 drain_right.n5 0.302913
R286 drain_right.n6 drain_right.n2 0.302913
C0 drain_right source 37.1375f
C1 plus drain_left 13.7862f
C2 drain_right minus 13.569f
C3 minus source 13.133f
C4 drain_right plus 0.372806f
C5 plus source 13.147f
C6 plus minus 7.38812f
C7 drain_right drain_left 1.15071f
C8 drain_left source 37.1363f
C9 drain_left minus 0.172419f
C10 drain_right a_n2210_n4888# 8.10894f
C11 drain_left a_n2210_n4888# 8.42976f
C12 source a_n2210_n4888# 13.406878f
C13 minus a_n2210_n4888# 9.279306f
C14 plus a_n2210_n4888# 11.59166f
C15 drain_right.t12 a_n2210_n4888# 0.465083f
C16 drain_right.t13 a_n2210_n4888# 0.465083f
C17 drain_right.n0 a_n2210_n4888# 4.25657f
C18 drain_right.t3 a_n2210_n4888# 0.465083f
C19 drain_right.t5 a_n2210_n4888# 0.465083f
C20 drain_right.n1 a_n2210_n4888# 4.25189f
C21 drain_right.n2 a_n2210_n4888# 0.738285f
C22 drain_right.t2 a_n2210_n4888# 0.465083f
C23 drain_right.t7 a_n2210_n4888# 0.465083f
C24 drain_right.n3 a_n2210_n4888# 4.25657f
C25 drain_right.t9 a_n2210_n4888# 0.465083f
C26 drain_right.t1 a_n2210_n4888# 0.465083f
C27 drain_right.n4 a_n2210_n4888# 4.25189f
C28 drain_right.n5 a_n2210_n4888# 0.738285f
C29 drain_right.n6 a_n2210_n4888# 2.08382f
C30 drain_right.t14 a_n2210_n4888# 0.465083f
C31 drain_right.t4 a_n2210_n4888# 0.465083f
C32 drain_right.n7 a_n2210_n4888# 4.25656f
C33 drain_right.t0 a_n2210_n4888# 0.465083f
C34 drain_right.t10 a_n2210_n4888# 0.465083f
C35 drain_right.n8 a_n2210_n4888# 4.25188f
C36 drain_right.n9 a_n2210_n4888# 0.775212f
C37 drain_right.t8 a_n2210_n4888# 0.465083f
C38 drain_right.t11 a_n2210_n4888# 0.465083f
C39 drain_right.n10 a_n2210_n4888# 4.25188f
C40 drain_right.n11 a_n2210_n4888# 0.384019f
C41 drain_right.t6 a_n2210_n4888# 0.465083f
C42 drain_right.t15 a_n2210_n4888# 0.465083f
C43 drain_right.n12 a_n2210_n4888# 4.25188f
C44 drain_right.n13 a_n2210_n4888# 0.636839f
C45 minus.n0 a_n2210_n4888# 0.044978f
C46 minus.t7 a_n2210_n4888# 1.27374f
C47 minus.n1 a_n2210_n4888# 0.483197f
C48 minus.n2 a_n2210_n4888# 0.044978f
C49 minus.n3 a_n2210_n4888# 0.010207f
C50 minus.t15 a_n2210_n4888# 1.27374f
C51 minus.n4 a_n2210_n4888# 0.143204f
C52 minus.t1 a_n2210_n4888# 1.27374f
C53 minus.t11 a_n2210_n4888# 1.28318f
C54 minus.n5 a_n2210_n4888# 0.46937f
C55 minus.n6 a_n2210_n4888# 0.480563f
C56 minus.n7 a_n2210_n4888# 0.010207f
C57 minus.t5 a_n2210_n4888# 1.27374f
C58 minus.n8 a_n2210_n4888# 0.483197f
C59 minus.n9 a_n2210_n4888# 0.044978f
C60 minus.n10 a_n2210_n4888# 0.044978f
C61 minus.n11 a_n2210_n4888# 0.044978f
C62 minus.n12 a_n2210_n4888# 0.48084f
C63 minus.t4 a_n2210_n4888# 1.27374f
C64 minus.n13 a_n2210_n4888# 0.48084f
C65 minus.n14 a_n2210_n4888# 0.010207f
C66 minus.n15 a_n2210_n4888# 0.044978f
C67 minus.n16 a_n2210_n4888# 0.044978f
C68 minus.n17 a_n2210_n4888# 0.044978f
C69 minus.n18 a_n2210_n4888# 0.010207f
C70 minus.t0 a_n2210_n4888# 1.27374f
C71 minus.n19 a_n2210_n4888# 0.480563f
C72 minus.t9 a_n2210_n4888# 1.27374f
C73 minus.n20 a_n2210_n4888# 0.478483f
C74 minus.n21 a_n2210_n4888# 2.10662f
C75 minus.n22 a_n2210_n4888# 0.044978f
C76 minus.t14 a_n2210_n4888# 1.27374f
C77 minus.n23 a_n2210_n4888# 0.483197f
C78 minus.n24 a_n2210_n4888# 0.044978f
C79 minus.n25 a_n2210_n4888# 0.010207f
C80 minus.n26 a_n2210_n4888# 0.143204f
C81 minus.t3 a_n2210_n4888# 1.28318f
C82 minus.n27 a_n2210_n4888# 0.46937f
C83 minus.t2 a_n2210_n4888# 1.27374f
C84 minus.n28 a_n2210_n4888# 0.480563f
C85 minus.n29 a_n2210_n4888# 0.010207f
C86 minus.t12 a_n2210_n4888# 1.27374f
C87 minus.n30 a_n2210_n4888# 0.483197f
C88 minus.n31 a_n2210_n4888# 0.044978f
C89 minus.n32 a_n2210_n4888# 0.044978f
C90 minus.n33 a_n2210_n4888# 0.044978f
C91 minus.t10 a_n2210_n4888# 1.27374f
C92 minus.n34 a_n2210_n4888# 0.48084f
C93 minus.t6 a_n2210_n4888# 1.27374f
C94 minus.n35 a_n2210_n4888# 0.48084f
C95 minus.n36 a_n2210_n4888# 0.010207f
C96 minus.n37 a_n2210_n4888# 0.044978f
C97 minus.n38 a_n2210_n4888# 0.044978f
C98 minus.n39 a_n2210_n4888# 0.044978f
C99 minus.n40 a_n2210_n4888# 0.010207f
C100 minus.t13 a_n2210_n4888# 1.27374f
C101 minus.n41 a_n2210_n4888# 0.480563f
C102 minus.t8 a_n2210_n4888# 1.27374f
C103 minus.n42 a_n2210_n4888# 0.478483f
C104 minus.n43 a_n2210_n4888# 0.300513f
C105 minus.n44 a_n2210_n4888# 2.50283f
C106 drain_left.t13 a_n2210_n4888# 0.46586f
C107 drain_left.t8 a_n2210_n4888# 0.46586f
C108 drain_left.n0 a_n2210_n4888# 4.26368f
C109 drain_left.t5 a_n2210_n4888# 0.46586f
C110 drain_left.t11 a_n2210_n4888# 0.46586f
C111 drain_left.n1 a_n2210_n4888# 4.25899f
C112 drain_left.n2 a_n2210_n4888# 0.739519f
C113 drain_left.t14 a_n2210_n4888# 0.46586f
C114 drain_left.t15 a_n2210_n4888# 0.46586f
C115 drain_left.n3 a_n2210_n4888# 4.26368f
C116 drain_left.t12 a_n2210_n4888# 0.46586f
C117 drain_left.t7 a_n2210_n4888# 0.46586f
C118 drain_left.n4 a_n2210_n4888# 4.25899f
C119 drain_left.n5 a_n2210_n4888# 0.739519f
C120 drain_left.n6 a_n2210_n4888# 2.14833f
C121 drain_left.t10 a_n2210_n4888# 0.46586f
C122 drain_left.t4 a_n2210_n4888# 0.46586f
C123 drain_left.n7 a_n2210_n4888# 4.26367f
C124 drain_left.t1 a_n2210_n4888# 0.46586f
C125 drain_left.t9 a_n2210_n4888# 0.46586f
C126 drain_left.n8 a_n2210_n4888# 4.25899f
C127 drain_left.n9 a_n2210_n4888# 0.776507f
C128 drain_left.t3 a_n2210_n4888# 0.46586f
C129 drain_left.t0 a_n2210_n4888# 0.46586f
C130 drain_left.n10 a_n2210_n4888# 4.25899f
C131 drain_left.n11 a_n2210_n4888# 0.384661f
C132 drain_left.t6 a_n2210_n4888# 0.46586f
C133 drain_left.t2 a_n2210_n4888# 0.46586f
C134 drain_left.n12 a_n2210_n4888# 4.25899f
C135 drain_left.n13 a_n2210_n4888# 0.637903f
C136 source.t19 a_n2210_n4888# 4.36453f
C137 source.n0 a_n2210_n4888# 1.87754f
C138 source.t22 a_n2210_n4888# 0.381903f
C139 source.t20 a_n2210_n4888# 0.381903f
C140 source.n1 a_n2210_n4888# 3.41437f
C141 source.n2 a_n2210_n4888# 0.359554f
C142 source.t30 a_n2210_n4888# 0.381903f
C143 source.t25 a_n2210_n4888# 0.381903f
C144 source.n3 a_n2210_n4888# 3.41437f
C145 source.n4 a_n2210_n4888# 0.359554f
C146 source.t24 a_n2210_n4888# 0.381903f
C147 source.t27 a_n2210_n4888# 0.381903f
C148 source.n5 a_n2210_n4888# 3.41437f
C149 source.n6 a_n2210_n4888# 0.359554f
C150 source.t21 a_n2210_n4888# 4.36454f
C151 source.n7 a_n2210_n4888# 0.431812f
C152 source.t12 a_n2210_n4888# 4.36454f
C153 source.n8 a_n2210_n4888# 0.431812f
C154 source.t1 a_n2210_n4888# 0.381903f
C155 source.t9 a_n2210_n4888# 0.381903f
C156 source.n9 a_n2210_n4888# 3.41437f
C157 source.n10 a_n2210_n4888# 0.359554f
C158 source.t14 a_n2210_n4888# 0.381903f
C159 source.t4 a_n2210_n4888# 0.381903f
C160 source.n11 a_n2210_n4888# 3.41437f
C161 source.n12 a_n2210_n4888# 0.359554f
C162 source.t0 a_n2210_n4888# 0.381903f
C163 source.t2 a_n2210_n4888# 0.381903f
C164 source.n13 a_n2210_n4888# 3.41437f
C165 source.n14 a_n2210_n4888# 0.359554f
C166 source.t15 a_n2210_n4888# 4.36454f
C167 source.n15 a_n2210_n4888# 2.31144f
C168 source.t17 a_n2210_n4888# 4.36451f
C169 source.n16 a_n2210_n4888# 2.31147f
C170 source.t29 a_n2210_n4888# 0.381903f
C171 source.t31 a_n2210_n4888# 0.381903f
C172 source.n17 a_n2210_n4888# 3.41438f
C173 source.n18 a_n2210_n4888# 0.359547f
C174 source.t26 a_n2210_n4888# 0.381903f
C175 source.t16 a_n2210_n4888# 0.381903f
C176 source.n19 a_n2210_n4888# 3.41438f
C177 source.n20 a_n2210_n4888# 0.359547f
C178 source.t28 a_n2210_n4888# 0.381903f
C179 source.t18 a_n2210_n4888# 0.381903f
C180 source.n21 a_n2210_n4888# 3.41438f
C181 source.n22 a_n2210_n4888# 0.359547f
C182 source.t23 a_n2210_n4888# 4.36451f
C183 source.n23 a_n2210_n4888# 0.431836f
C184 source.t10 a_n2210_n4888# 4.36451f
C185 source.n24 a_n2210_n4888# 0.431836f
C186 source.t3 a_n2210_n4888# 0.381903f
C187 source.t5 a_n2210_n4888# 0.381903f
C188 source.n25 a_n2210_n4888# 3.41438f
C189 source.n26 a_n2210_n4888# 0.359547f
C190 source.t8 a_n2210_n4888# 0.381903f
C191 source.t13 a_n2210_n4888# 0.381903f
C192 source.n27 a_n2210_n4888# 3.41438f
C193 source.n28 a_n2210_n4888# 0.359547f
C194 source.t11 a_n2210_n4888# 0.381903f
C195 source.t7 a_n2210_n4888# 0.381903f
C196 source.n29 a_n2210_n4888# 3.41438f
C197 source.n30 a_n2210_n4888# 0.359547f
C198 source.t6 a_n2210_n4888# 4.36451f
C199 source.n31 a_n2210_n4888# 0.57891f
C200 source.n32 a_n2210_n4888# 2.18366f
C201 plus.n0 a_n2210_n4888# 0.045363f
C202 plus.t13 a_n2210_n4888# 1.28464f
C203 plus.t9 a_n2210_n4888# 1.28464f
C204 plus.t15 a_n2210_n4888# 1.28464f
C205 plus.n1 a_n2210_n4888# 0.487331f
C206 plus.n2 a_n2210_n4888# 0.045363f
C207 plus.t12 a_n2210_n4888# 1.28464f
C208 plus.t6 a_n2210_n4888# 1.28464f
C209 plus.n3 a_n2210_n4888# 0.045363f
C210 plus.t14 a_n2210_n4888# 1.28464f
C211 plus.n4 a_n2210_n4888# 0.487331f
C212 plus.t5 a_n2210_n4888# 1.29416f
C213 plus.n5 a_n2210_n4888# 0.473386f
C214 plus.t11 a_n2210_n4888# 1.28464f
C215 plus.n6 a_n2210_n4888# 0.484674f
C216 plus.n7 a_n2210_n4888# 0.010294f
C217 plus.n8 a_n2210_n4888# 0.144429f
C218 plus.n9 a_n2210_n4888# 0.045363f
C219 plus.n10 a_n2210_n4888# 0.045363f
C220 plus.n11 a_n2210_n4888# 0.010294f
C221 plus.n12 a_n2210_n4888# 0.484954f
C222 plus.n13 a_n2210_n4888# 0.484954f
C223 plus.n14 a_n2210_n4888# 0.010294f
C224 plus.n15 a_n2210_n4888# 0.045363f
C225 plus.n16 a_n2210_n4888# 0.045363f
C226 plus.n17 a_n2210_n4888# 0.045363f
C227 plus.n18 a_n2210_n4888# 0.010294f
C228 plus.n19 a_n2210_n4888# 0.484674f
C229 plus.n20 a_n2210_n4888# 0.482577f
C230 plus.n21 a_n2210_n4888# 0.695177f
C231 plus.n22 a_n2210_n4888# 0.045363f
C232 plus.t2 a_n2210_n4888# 1.28464f
C233 plus.t7 a_n2210_n4888# 1.28464f
C234 plus.t10 a_n2210_n4888# 1.28464f
C235 plus.n23 a_n2210_n4888# 0.487331f
C236 plus.n24 a_n2210_n4888# 0.045363f
C237 plus.t4 a_n2210_n4888# 1.28464f
C238 plus.n25 a_n2210_n4888# 0.045363f
C239 plus.t3 a_n2210_n4888# 1.28464f
C240 plus.t8 a_n2210_n4888# 1.28464f
C241 plus.n26 a_n2210_n4888# 0.487331f
C242 plus.t0 a_n2210_n4888# 1.29416f
C243 plus.n27 a_n2210_n4888# 0.473386f
C244 plus.t1 a_n2210_n4888# 1.28464f
C245 plus.n28 a_n2210_n4888# 0.484674f
C246 plus.n29 a_n2210_n4888# 0.010294f
C247 plus.n30 a_n2210_n4888# 0.144429f
C248 plus.n31 a_n2210_n4888# 0.045363f
C249 plus.n32 a_n2210_n4888# 0.045363f
C250 plus.n33 a_n2210_n4888# 0.010294f
C251 plus.n34 a_n2210_n4888# 0.484954f
C252 plus.n35 a_n2210_n4888# 0.484954f
C253 plus.n36 a_n2210_n4888# 0.010294f
C254 plus.n37 a_n2210_n4888# 0.045363f
C255 plus.n38 a_n2210_n4888# 0.045363f
C256 plus.n39 a_n2210_n4888# 0.045363f
C257 plus.n40 a_n2210_n4888# 0.010294f
C258 plus.n41 a_n2210_n4888# 0.484674f
C259 plus.n42 a_n2210_n4888# 0.482577f
C260 plus.n43 a_n2210_n4888# 1.69075f
.ends

