* NGSPICE file created from diffpair135.ext - technology: sky130A

.subckt diffpair135 minus drain_right drain_left source plus
X0 source.t20 minus.t0 drain_right.t3 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X1 drain_left.t11 plus.t0 source.t1 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X2 source.t22 plus.t1 drain_left.t10 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X3 drain_right.t7 minus.t1 source.t19 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X4 drain_right.t8 minus.t2 source.t18 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X5 a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X6 drain_right.t0 minus.t3 source.t17 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 source.t16 minus.t4 drain_right.t4 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X8 source.t15 minus.t5 drain_right.t11 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_left.t9 plus.t2 source.t8 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X10 source.t21 plus.t3 drain_left.t8 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X11 source.t7 plus.t4 drain_left.t7 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X12 source.t14 minus.t6 drain_right.t1 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X13 drain_right.t9 minus.t7 source.t13 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 drain_left.t6 plus.t5 source.t0 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 source.t12 minus.t8 drain_right.t6 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 source.t23 plus.t6 drain_left.t5 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 drain_right.t2 minus.t9 source.t11 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X18 source.t10 minus.t10 drain_right.t5 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X20 drain_left.t4 plus.t7 source.t4 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X21 source.t3 plus.t8 drain_left.t3 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X22 a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X23 source.t6 plus.t9 drain_left.t2 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X24 drain_right.t10 minus.t11 source.t9 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X25 a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X26 drain_left.t1 plus.t10 source.t5 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X27 drain_left.t0 plus.t11 source.t2 a_n2018_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
R0 minus.n2 minus.t9 170.865
R1 minus.n14 minus.t4 170.865
R2 minus.n11 minus.n10 161.3
R3 minus.n9 minus.n0 161.3
R4 minus.n8 minus.n7 161.3
R5 minus.n23 minus.n22 161.3
R6 minus.n21 minus.n12 161.3
R7 minus.n20 minus.n19 161.3
R8 minus.n3 minus.t8 145.805
R9 minus.n4 minus.t7 145.805
R10 minus.n1 minus.t6 145.805
R11 minus.n8 minus.t2 145.805
R12 minus.n10 minus.t5 145.805
R13 minus.n15 minus.t11 145.805
R14 minus.n16 minus.t10 145.805
R15 minus.n13 minus.t3 145.805
R16 minus.n20 minus.t0 145.805
R17 minus.n22 minus.t1 145.805
R18 minus.n6 minus.n1 80.6037
R19 minus.n5 minus.n4 80.6037
R20 minus.n18 minus.n13 80.6037
R21 minus.n17 minus.n16 80.6037
R22 minus.n4 minus.n3 48.2005
R23 minus.n4 minus.n1 48.2005
R24 minus.n8 minus.n1 48.2005
R25 minus.n16 minus.n15 48.2005
R26 minus.n16 minus.n13 48.2005
R27 minus.n20 minus.n13 48.2005
R28 minus.n5 minus.n2 45.0744
R29 minus.n17 minus.n14 45.0744
R30 minus.n10 minus.n9 40.1672
R31 minus.n22 minus.n21 40.1672
R32 minus.n24 minus.n11 29.277
R33 minus.n3 minus.n2 16.1124
R34 minus.n15 minus.n14 16.1124
R35 minus.n9 minus.n8 8.03383
R36 minus.n21 minus.n20 8.03383
R37 minus.n24 minus.n23 6.58762
R38 minus.n6 minus.n5 0.380177
R39 minus.n18 minus.n17 0.380177
R40 minus.n7 minus.n6 0.285035
R41 minus.n19 minus.n18 0.285035
R42 minus.n11 minus.n0 0.189894
R43 minus.n7 minus.n0 0.189894
R44 minus.n19 minus.n12 0.189894
R45 minus.n23 minus.n12 0.189894
R46 minus minus.n24 0.188
R47 drain_right.n6 drain_right.n4 101.597
R48 drain_right.n3 drain_right.n2 101.541
R49 drain_right.n3 drain_right.n0 101.541
R50 drain_right.n6 drain_right.n5 100.796
R51 drain_right.n8 drain_right.n7 100.796
R52 drain_right.n3 drain_right.n1 100.796
R53 drain_right drain_right.n3 23.2467
R54 drain_right.n1 drain_right.t5 9.9005
R55 drain_right.n1 drain_right.t0 9.9005
R56 drain_right.n2 drain_right.t3 9.9005
R57 drain_right.n2 drain_right.t7 9.9005
R58 drain_right.n0 drain_right.t4 9.9005
R59 drain_right.n0 drain_right.t10 9.9005
R60 drain_right.n4 drain_right.t6 9.9005
R61 drain_right.n4 drain_right.t2 9.9005
R62 drain_right.n5 drain_right.t1 9.9005
R63 drain_right.n5 drain_right.t9 9.9005
R64 drain_right.n7 drain_right.t11 9.9005
R65 drain_right.n7 drain_right.t8 9.9005
R66 drain_right drain_right.n8 6.45494
R67 drain_right.n8 drain_right.n6 0.802224
R68 source.n74 source.n72 289.615
R69 source.n62 source.n60 289.615
R70 source.n54 source.n52 289.615
R71 source.n42 source.n40 289.615
R72 source.n2 source.n0 289.615
R73 source.n14 source.n12 289.615
R74 source.n22 source.n20 289.615
R75 source.n34 source.n32 289.615
R76 source.n75 source.n74 185
R77 source.n63 source.n62 185
R78 source.n55 source.n54 185
R79 source.n43 source.n42 185
R80 source.n3 source.n2 185
R81 source.n15 source.n14 185
R82 source.n23 source.n22 185
R83 source.n35 source.n34 185
R84 source.t19 source.n73 167.117
R85 source.t16 source.n61 167.117
R86 source.t5 source.n53 167.117
R87 source.t6 source.n41 167.117
R88 source.t1 source.n1 167.117
R89 source.t3 source.n13 167.117
R90 source.t11 source.n21 167.117
R91 source.t15 source.n33 167.117
R92 source.n9 source.n8 84.1169
R93 source.n11 source.n10 84.1169
R94 source.n29 source.n28 84.1169
R95 source.n31 source.n30 84.1169
R96 source.n71 source.n70 84.1168
R97 source.n69 source.n68 84.1168
R98 source.n51 source.n50 84.1168
R99 source.n49 source.n48 84.1168
R100 source.n74 source.t19 52.3082
R101 source.n62 source.t16 52.3082
R102 source.n54 source.t5 52.3082
R103 source.n42 source.t6 52.3082
R104 source.n2 source.t1 52.3082
R105 source.n14 source.t3 52.3082
R106 source.n22 source.t11 52.3082
R107 source.n34 source.t15 52.3082
R108 source.n79 source.n78 31.4096
R109 source.n67 source.n66 31.4096
R110 source.n59 source.n58 31.4096
R111 source.n47 source.n46 31.4096
R112 source.n7 source.n6 31.4096
R113 source.n19 source.n18 31.4096
R114 source.n27 source.n26 31.4096
R115 source.n39 source.n38 31.4096
R116 source.n47 source.n39 14.5137
R117 source.n70 source.t17 9.9005
R118 source.n70 source.t20 9.9005
R119 source.n68 source.t9 9.9005
R120 source.n68 source.t10 9.9005
R121 source.n50 source.t8 9.9005
R122 source.n50 source.t7 9.9005
R123 source.n48 source.t2 9.9005
R124 source.n48 source.t22 9.9005
R125 source.n8 source.t0 9.9005
R126 source.n8 source.t21 9.9005
R127 source.n10 source.t4 9.9005
R128 source.n10 source.t23 9.9005
R129 source.n28 source.t13 9.9005
R130 source.n28 source.t12 9.9005
R131 source.n30 source.t18 9.9005
R132 source.n30 source.t14 9.9005
R133 source.n75 source.n73 9.71174
R134 source.n63 source.n61 9.71174
R135 source.n55 source.n53 9.71174
R136 source.n43 source.n41 9.71174
R137 source.n3 source.n1 9.71174
R138 source.n15 source.n13 9.71174
R139 source.n23 source.n21 9.71174
R140 source.n35 source.n33 9.71174
R141 source.n78 source.n77 9.45567
R142 source.n66 source.n65 9.45567
R143 source.n58 source.n57 9.45567
R144 source.n46 source.n45 9.45567
R145 source.n6 source.n5 9.45567
R146 source.n18 source.n17 9.45567
R147 source.n26 source.n25 9.45567
R148 source.n38 source.n37 9.45567
R149 source.n77 source.n76 9.3005
R150 source.n65 source.n64 9.3005
R151 source.n57 source.n56 9.3005
R152 source.n45 source.n44 9.3005
R153 source.n5 source.n4 9.3005
R154 source.n17 source.n16 9.3005
R155 source.n25 source.n24 9.3005
R156 source.n37 source.n36 9.3005
R157 source.n80 source.n7 8.8499
R158 source.n78 source.n72 8.14595
R159 source.n66 source.n60 8.14595
R160 source.n58 source.n52 8.14595
R161 source.n46 source.n40 8.14595
R162 source.n6 source.n0 8.14595
R163 source.n18 source.n12 8.14595
R164 source.n26 source.n20 8.14595
R165 source.n38 source.n32 8.14595
R166 source.n76 source.n75 7.3702
R167 source.n64 source.n63 7.3702
R168 source.n56 source.n55 7.3702
R169 source.n44 source.n43 7.3702
R170 source.n4 source.n3 7.3702
R171 source.n16 source.n15 7.3702
R172 source.n24 source.n23 7.3702
R173 source.n36 source.n35 7.3702
R174 source.n76 source.n72 5.81868
R175 source.n64 source.n60 5.81868
R176 source.n56 source.n52 5.81868
R177 source.n44 source.n40 5.81868
R178 source.n4 source.n0 5.81868
R179 source.n16 source.n12 5.81868
R180 source.n24 source.n20 5.81868
R181 source.n36 source.n32 5.81868
R182 source.n80 source.n79 5.66429
R183 source.n77 source.n73 3.44771
R184 source.n65 source.n61 3.44771
R185 source.n57 source.n53 3.44771
R186 source.n45 source.n41 3.44771
R187 source.n5 source.n1 3.44771
R188 source.n17 source.n13 3.44771
R189 source.n25 source.n21 3.44771
R190 source.n37 source.n33 3.44771
R191 source.n39 source.n31 0.802224
R192 source.n31 source.n29 0.802224
R193 source.n29 source.n27 0.802224
R194 source.n19 source.n11 0.802224
R195 source.n11 source.n9 0.802224
R196 source.n9 source.n7 0.802224
R197 source.n49 source.n47 0.802224
R198 source.n51 source.n49 0.802224
R199 source.n59 source.n51 0.802224
R200 source.n69 source.n67 0.802224
R201 source.n71 source.n69 0.802224
R202 source.n79 source.n71 0.802224
R203 source.n27 source.n19 0.470328
R204 source.n67 source.n59 0.470328
R205 source source.n80 0.188
R206 plus.n4 plus.t8 170.865
R207 plus.n16 plus.t10 170.865
R208 plus.n8 plus.n1 161.3
R209 plus.n9 plus.n0 161.3
R210 plus.n11 plus.n10 161.3
R211 plus.n20 plus.n13 161.3
R212 plus.n21 plus.n12 161.3
R213 plus.n23 plus.n22 161.3
R214 plus.n10 plus.t0 145.805
R215 plus.n8 plus.t3 145.805
R216 plus.n7 plus.t5 145.805
R217 plus.n6 plus.t6 145.805
R218 plus.n5 plus.t7 145.805
R219 plus.n22 plus.t9 145.805
R220 plus.n20 plus.t11 145.805
R221 plus.n19 plus.t1 145.805
R222 plus.n18 plus.t2 145.805
R223 plus.n17 plus.t4 145.805
R224 plus.n6 plus.n3 80.6037
R225 plus.n7 plus.n2 80.6037
R226 plus.n18 plus.n15 80.6037
R227 plus.n19 plus.n14 80.6037
R228 plus.n8 plus.n7 48.2005
R229 plus.n7 plus.n6 48.2005
R230 plus.n6 plus.n5 48.2005
R231 plus.n20 plus.n19 48.2005
R232 plus.n19 plus.n18 48.2005
R233 plus.n18 plus.n17 48.2005
R234 plus.n4 plus.n3 45.0744
R235 plus.n16 plus.n15 45.0744
R236 plus.n10 plus.n9 40.1672
R237 plus.n22 plus.n21 40.1672
R238 plus plus.n23 26.946
R239 plus.n5 plus.n4 16.1124
R240 plus.n17 plus.n16 16.1124
R241 plus plus.n11 8.44368
R242 plus.n9 plus.n8 8.03383
R243 plus.n21 plus.n20 8.03383
R244 plus.n3 plus.n2 0.380177
R245 plus.n15 plus.n14 0.380177
R246 plus.n2 plus.n1 0.285035
R247 plus.n14 plus.n13 0.285035
R248 plus.n1 plus.n0 0.189894
R249 plus.n11 plus.n0 0.189894
R250 plus.n23 plus.n12 0.189894
R251 plus.n13 plus.n12 0.189894
R252 drain_left.n6 drain_left.n4 101.597
R253 drain_left.n3 drain_left.n2 101.541
R254 drain_left.n3 drain_left.n0 101.541
R255 drain_left.n8 drain_left.n7 100.796
R256 drain_left.n6 drain_left.n5 100.796
R257 drain_left.n3 drain_left.n1 100.796
R258 drain_left drain_left.n3 23.7999
R259 drain_left.n1 drain_left.t10 9.9005
R260 drain_left.n1 drain_left.t9 9.9005
R261 drain_left.n2 drain_left.t7 9.9005
R262 drain_left.n2 drain_left.t1 9.9005
R263 drain_left.n0 drain_left.t2 9.9005
R264 drain_left.n0 drain_left.t0 9.9005
R265 drain_left.n7 drain_left.t8 9.9005
R266 drain_left.n7 drain_left.t11 9.9005
R267 drain_left.n5 drain_left.t5 9.9005
R268 drain_left.n5 drain_left.t6 9.9005
R269 drain_left.n4 drain_left.t3 9.9005
R270 drain_left.n4 drain_left.t4 9.9005
R271 drain_left drain_left.n8 6.45494
R272 drain_left.n8 drain_left.n6 0.802224
C0 drain_right minus 1.60036f
C1 source drain_right 5.01739f
C2 drain_right drain_left 1.01278f
C3 drain_right plus 0.359025f
C4 source minus 1.95743f
C5 minus drain_left 0.177888f
C6 plus minus 3.81991f
C7 source drain_left 5.01588f
C8 source plus 1.9714f
C9 plus drain_left 1.79744f
C10 drain_right a_n2018_n1288# 3.72189f
C11 drain_left a_n2018_n1288# 3.9778f
C12 source a_n2018_n1288# 3.163961f
C13 minus a_n2018_n1288# 7.111672f
C14 plus a_n2018_n1288# 7.638922f
C15 drain_left.t2 a_n2018_n1288# 0.031428f
C16 drain_left.t0 a_n2018_n1288# 0.031428f
C17 drain_left.n0 a_n2018_n1288# 0.199352f
C18 drain_left.t10 a_n2018_n1288# 0.031428f
C19 drain_left.t9 a_n2018_n1288# 0.031428f
C20 drain_left.n1 a_n2018_n1288# 0.197441f
C21 drain_left.t7 a_n2018_n1288# 0.031428f
C22 drain_left.t1 a_n2018_n1288# 0.031428f
C23 drain_left.n2 a_n2018_n1288# 0.199352f
C24 drain_left.n3 a_n2018_n1288# 1.33651f
C25 drain_left.t3 a_n2018_n1288# 0.031428f
C26 drain_left.t4 a_n2018_n1288# 0.031428f
C27 drain_left.n4 a_n2018_n1288# 0.199517f
C28 drain_left.t5 a_n2018_n1288# 0.031428f
C29 drain_left.t6 a_n2018_n1288# 0.031428f
C30 drain_left.n5 a_n2018_n1288# 0.197442f
C31 drain_left.n6 a_n2018_n1288# 0.515818f
C32 drain_left.t8 a_n2018_n1288# 0.031428f
C33 drain_left.t11 a_n2018_n1288# 0.031428f
C34 drain_left.n7 a_n2018_n1288# 0.197442f
C35 drain_left.n8 a_n2018_n1288# 0.428341f
C36 plus.n0 a_n2018_n1288# 0.024126f
C37 plus.t0 a_n2018_n1288# 0.089655f
C38 plus.t3 a_n2018_n1288# 0.089655f
C39 plus.n1 a_n2018_n1288# 0.032193f
C40 plus.t5 a_n2018_n1288# 0.089655f
C41 plus.n2 a_n2018_n1288# 0.040185f
C42 plus.t6 a_n2018_n1288# 0.089655f
C43 plus.n3 a_n2018_n1288# 0.12365f
C44 plus.t7 a_n2018_n1288# 0.089655f
C45 plus.t8 a_n2018_n1288# 0.098928f
C46 plus.n4 a_n2018_n1288# 0.055794f
C47 plus.n5 a_n2018_n1288# 0.06808f
C48 plus.n6 a_n2018_n1288# 0.068961f
C49 plus.n7 a_n2018_n1288# 0.068961f
C50 plus.n8 a_n2018_n1288# 0.064305f
C51 plus.n9 a_n2018_n1288# 0.005475f
C52 plus.n10 a_n2018_n1288# 0.062669f
C53 plus.n11 a_n2018_n1288# 0.177705f
C54 plus.n12 a_n2018_n1288# 0.024126f
C55 plus.t9 a_n2018_n1288# 0.089655f
C56 plus.n13 a_n2018_n1288# 0.032193f
C57 plus.t11 a_n2018_n1288# 0.089655f
C58 plus.n14 a_n2018_n1288# 0.040185f
C59 plus.t1 a_n2018_n1288# 0.089655f
C60 plus.n15 a_n2018_n1288# 0.12365f
C61 plus.t2 a_n2018_n1288# 0.089655f
C62 plus.t10 a_n2018_n1288# 0.098928f
C63 plus.n16 a_n2018_n1288# 0.055794f
C64 plus.t4 a_n2018_n1288# 0.089655f
C65 plus.n17 a_n2018_n1288# 0.06808f
C66 plus.n18 a_n2018_n1288# 0.068961f
C67 plus.n19 a_n2018_n1288# 0.068961f
C68 plus.n20 a_n2018_n1288# 0.064305f
C69 plus.n21 a_n2018_n1288# 0.005475f
C70 plus.n22 a_n2018_n1288# 0.062669f
C71 plus.n23 a_n2018_n1288# 0.575949f
C72 source.n0 a_n2018_n1288# 0.030374f
C73 source.n1 a_n2018_n1288# 0.067207f
C74 source.t1 a_n2018_n1288# 0.050435f
C75 source.n2 a_n2018_n1288# 0.052599f
C76 source.n3 a_n2018_n1288# 0.016956f
C77 source.n4 a_n2018_n1288# 0.011183f
C78 source.n5 a_n2018_n1288# 0.148141f
C79 source.n6 a_n2018_n1288# 0.033297f
C80 source.n7 a_n2018_n1288# 0.344955f
C81 source.t0 a_n2018_n1288# 0.03289f
C82 source.t21 a_n2018_n1288# 0.03289f
C83 source.n8 a_n2018_n1288# 0.175831f
C84 source.n9 a_n2018_n1288# 0.269314f
C85 source.t4 a_n2018_n1288# 0.03289f
C86 source.t23 a_n2018_n1288# 0.03289f
C87 source.n10 a_n2018_n1288# 0.175831f
C88 source.n11 a_n2018_n1288# 0.269314f
C89 source.n12 a_n2018_n1288# 0.030374f
C90 source.n13 a_n2018_n1288# 0.067207f
C91 source.t3 a_n2018_n1288# 0.050435f
C92 source.n14 a_n2018_n1288# 0.052599f
C93 source.n15 a_n2018_n1288# 0.016956f
C94 source.n16 a_n2018_n1288# 0.011183f
C95 source.n17 a_n2018_n1288# 0.148141f
C96 source.n18 a_n2018_n1288# 0.033297f
C97 source.n19 a_n2018_n1288# 0.102398f
C98 source.n20 a_n2018_n1288# 0.030374f
C99 source.n21 a_n2018_n1288# 0.067207f
C100 source.t11 a_n2018_n1288# 0.050435f
C101 source.n22 a_n2018_n1288# 0.052599f
C102 source.n23 a_n2018_n1288# 0.016956f
C103 source.n24 a_n2018_n1288# 0.011183f
C104 source.n25 a_n2018_n1288# 0.148141f
C105 source.n26 a_n2018_n1288# 0.033297f
C106 source.n27 a_n2018_n1288# 0.102398f
C107 source.t13 a_n2018_n1288# 0.03289f
C108 source.t12 a_n2018_n1288# 0.03289f
C109 source.n28 a_n2018_n1288# 0.175831f
C110 source.n29 a_n2018_n1288# 0.269314f
C111 source.t18 a_n2018_n1288# 0.03289f
C112 source.t14 a_n2018_n1288# 0.03289f
C113 source.n30 a_n2018_n1288# 0.175831f
C114 source.n31 a_n2018_n1288# 0.269314f
C115 source.n32 a_n2018_n1288# 0.030374f
C116 source.n33 a_n2018_n1288# 0.067207f
C117 source.t15 a_n2018_n1288# 0.050435f
C118 source.n34 a_n2018_n1288# 0.052599f
C119 source.n35 a_n2018_n1288# 0.016956f
C120 source.n36 a_n2018_n1288# 0.011183f
C121 source.n37 a_n2018_n1288# 0.148141f
C122 source.n38 a_n2018_n1288# 0.033297f
C123 source.n39 a_n2018_n1288# 0.542908f
C124 source.n40 a_n2018_n1288# 0.030374f
C125 source.n41 a_n2018_n1288# 0.067207f
C126 source.t6 a_n2018_n1288# 0.050435f
C127 source.n42 a_n2018_n1288# 0.052599f
C128 source.n43 a_n2018_n1288# 0.016956f
C129 source.n44 a_n2018_n1288# 0.011183f
C130 source.n45 a_n2018_n1288# 0.148141f
C131 source.n46 a_n2018_n1288# 0.033297f
C132 source.n47 a_n2018_n1288# 0.542908f
C133 source.t2 a_n2018_n1288# 0.03289f
C134 source.t22 a_n2018_n1288# 0.03289f
C135 source.n48 a_n2018_n1288# 0.17583f
C136 source.n49 a_n2018_n1288# 0.269315f
C137 source.t8 a_n2018_n1288# 0.03289f
C138 source.t7 a_n2018_n1288# 0.03289f
C139 source.n50 a_n2018_n1288# 0.17583f
C140 source.n51 a_n2018_n1288# 0.269315f
C141 source.n52 a_n2018_n1288# 0.030374f
C142 source.n53 a_n2018_n1288# 0.067207f
C143 source.t5 a_n2018_n1288# 0.050435f
C144 source.n54 a_n2018_n1288# 0.052599f
C145 source.n55 a_n2018_n1288# 0.016956f
C146 source.n56 a_n2018_n1288# 0.011183f
C147 source.n57 a_n2018_n1288# 0.148141f
C148 source.n58 a_n2018_n1288# 0.033297f
C149 source.n59 a_n2018_n1288# 0.102398f
C150 source.n60 a_n2018_n1288# 0.030374f
C151 source.n61 a_n2018_n1288# 0.067207f
C152 source.t16 a_n2018_n1288# 0.050435f
C153 source.n62 a_n2018_n1288# 0.052599f
C154 source.n63 a_n2018_n1288# 0.016956f
C155 source.n64 a_n2018_n1288# 0.011183f
C156 source.n65 a_n2018_n1288# 0.148141f
C157 source.n66 a_n2018_n1288# 0.033297f
C158 source.n67 a_n2018_n1288# 0.102398f
C159 source.t9 a_n2018_n1288# 0.03289f
C160 source.t10 a_n2018_n1288# 0.03289f
C161 source.n68 a_n2018_n1288# 0.17583f
C162 source.n69 a_n2018_n1288# 0.269315f
C163 source.t17 a_n2018_n1288# 0.03289f
C164 source.t20 a_n2018_n1288# 0.03289f
C165 source.n70 a_n2018_n1288# 0.17583f
C166 source.n71 a_n2018_n1288# 0.269315f
C167 source.n72 a_n2018_n1288# 0.030374f
C168 source.n73 a_n2018_n1288# 0.067207f
C169 source.t19 a_n2018_n1288# 0.050435f
C170 source.n74 a_n2018_n1288# 0.052599f
C171 source.n75 a_n2018_n1288# 0.016956f
C172 source.n76 a_n2018_n1288# 0.011183f
C173 source.n77 a_n2018_n1288# 0.148141f
C174 source.n78 a_n2018_n1288# 0.033297f
C175 source.n79 a_n2018_n1288# 0.233616f
C176 source.n80 a_n2018_n1288# 0.522048f
C177 drain_right.t4 a_n2018_n1288# 0.031925f
C178 drain_right.t10 a_n2018_n1288# 0.031925f
C179 drain_right.n0 a_n2018_n1288# 0.202503f
C180 drain_right.t5 a_n2018_n1288# 0.031925f
C181 drain_right.t0 a_n2018_n1288# 0.031925f
C182 drain_right.n1 a_n2018_n1288# 0.200561f
C183 drain_right.t3 a_n2018_n1288# 0.031925f
C184 drain_right.t7 a_n2018_n1288# 0.031925f
C185 drain_right.n2 a_n2018_n1288# 0.202503f
C186 drain_right.n3 a_n2018_n1288# 1.31812f
C187 drain_right.t6 a_n2018_n1288# 0.031925f
C188 drain_right.t2 a_n2018_n1288# 0.031925f
C189 drain_right.n4 a_n2018_n1288# 0.20267f
C190 drain_right.t1 a_n2018_n1288# 0.031925f
C191 drain_right.t9 a_n2018_n1288# 0.031925f
C192 drain_right.n5 a_n2018_n1288# 0.200562f
C193 drain_right.n6 a_n2018_n1288# 0.52397f
C194 drain_right.t11 a_n2018_n1288# 0.031925f
C195 drain_right.t8 a_n2018_n1288# 0.031925f
C196 drain_right.n7 a_n2018_n1288# 0.200562f
C197 drain_right.n8 a_n2018_n1288# 0.43511f
C198 minus.n0 a_n2018_n1288# 0.02382f
C199 minus.t6 a_n2018_n1288# 0.088518f
C200 minus.n1 a_n2018_n1288# 0.068087f
C201 minus.t2 a_n2018_n1288# 0.088518f
C202 minus.t9 a_n2018_n1288# 0.097674f
C203 minus.n2 a_n2018_n1288# 0.055087f
C204 minus.t8 a_n2018_n1288# 0.088518f
C205 minus.n3 a_n2018_n1288# 0.067217f
C206 minus.t7 a_n2018_n1288# 0.088518f
C207 minus.n4 a_n2018_n1288# 0.068087f
C208 minus.n5 a_n2018_n1288# 0.122083f
C209 minus.n6 a_n2018_n1288# 0.039676f
C210 minus.n7 a_n2018_n1288# 0.031785f
C211 minus.n8 a_n2018_n1288# 0.06349f
C212 minus.n9 a_n2018_n1288# 0.005405f
C213 minus.t5 a_n2018_n1288# 0.088518f
C214 minus.n10 a_n2018_n1288# 0.061874f
C215 minus.n11 a_n2018_n1288# 0.596221f
C216 minus.n12 a_n2018_n1288# 0.02382f
C217 minus.t3 a_n2018_n1288# 0.088518f
C218 minus.n13 a_n2018_n1288# 0.068087f
C219 minus.t4 a_n2018_n1288# 0.097674f
C220 minus.n14 a_n2018_n1288# 0.055087f
C221 minus.t11 a_n2018_n1288# 0.088518f
C222 minus.n15 a_n2018_n1288# 0.067217f
C223 minus.t10 a_n2018_n1288# 0.088518f
C224 minus.n16 a_n2018_n1288# 0.068087f
C225 minus.n17 a_n2018_n1288# 0.122083f
C226 minus.n18 a_n2018_n1288# 0.039676f
C227 minus.n19 a_n2018_n1288# 0.031785f
C228 minus.t0 a_n2018_n1288# 0.088518f
C229 minus.n20 a_n2018_n1288# 0.06349f
C230 minus.n21 a_n2018_n1288# 0.005405f
C231 minus.t1 a_n2018_n1288# 0.088518f
C232 minus.n22 a_n2018_n1288# 0.061874f
C233 minus.n23 a_n2018_n1288# 0.160628f
C234 minus.n24 a_n2018_n1288# 0.733755f
.ends

