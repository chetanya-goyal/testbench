* NGSPICE file created from diffpair506.ext - technology: sky130A

.subckt diffpair506 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t2 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X1 source.t26 plus.t1 drain_left.t11 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X2 source.t25 plus.t2 drain_left.t9 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X3 source.t11 minus.t0 drain_right.t13 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X4 drain_left.t8 plus.t3 source.t24 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X5 source.t1 minus.t1 drain_right.t12 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X6 source.t5 minus.t2 drain_right.t11 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X7 drain_right.t10 minus.t3 source.t7 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 source.t23 plus.t4 drain_left.t7 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X9 drain_left.t13 plus.t5 source.t22 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X10 a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X11 source.t0 minus.t4 drain_right.t9 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X12 source.t8 minus.t5 drain_right.t8 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X13 drain_left.t4 plus.t6 source.t21 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X14 drain_right.t7 minus.t6 source.t4 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X15 drain_left.t12 plus.t7 source.t20 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X16 drain_left.t6 plus.t8 source.t19 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X17 drain_left.t5 plus.t9 source.t18 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X18 drain_left.t1 plus.t10 source.t17 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X19 drain_right.t6 minus.t7 source.t6 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X20 drain_right.t5 minus.t8 source.t9 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X21 a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X22 a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X23 source.t3 minus.t9 drain_right.t4 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X24 drain_right.t3 minus.t10 source.t12 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X25 drain_right.t2 minus.t11 source.t13 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X26 drain_left.t3 plus.t11 source.t16 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X27 source.t15 plus.t12 drain_left.t0 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X28 source.t14 plus.t13 drain_left.t10 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X29 a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X30 drain_right.t1 minus.t12 source.t2 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X31 drain_right.t0 minus.t13 source.t10 a_n1644_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
R0 plus.n3 plus.t5 1606.37
R1 plus.n15 plus.t7 1606.37
R2 plus.n20 plus.t3 1606.37
R3 plus.n32 plus.t11 1606.37
R4 plus.n1 plus.t0 1571.32
R5 plus.n4 plus.t1 1571.32
R6 plus.n6 plus.t9 1571.32
R7 plus.n12 plus.t8 1571.32
R8 plus.n14 plus.t13 1571.32
R9 plus.n18 plus.t4 1571.32
R10 plus.n21 plus.t12 1571.32
R11 plus.n23 plus.t10 1571.32
R12 plus.n29 plus.t6 1571.32
R13 plus.n31 plus.t2 1571.32
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 30.3172
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus plus.n16 13.2316
R46 plus.n7 plus.n6 11.6853
R47 plus.n12 plus.n11 11.6853
R48 plus.n29 plus.n28 11.6853
R49 plus.n24 plus.n23 11.6853
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t13 62.6998
R61 drain_left.n1 drain_left.t3 62.6996
R62 drain_left.n4 drain_left.n2 61.3796
R63 drain_left.n9 drain_left.n8 60.8798
R64 drain_left.n7 drain_left.n6 60.8798
R65 drain_left.n11 drain_left.n10 60.8796
R66 drain_left.n4 drain_left.n3 60.8796
R67 drain_left.n1 drain_left.n0 60.8796
R68 drain_left drain_left.n5 32.5148
R69 drain_left drain_left.n11 6.15322
R70 drain_left.n2 drain_left.t0 1.3205
R71 drain_left.n2 drain_left.t8 1.3205
R72 drain_left.n3 drain_left.t7 1.3205
R73 drain_left.n3 drain_left.t1 1.3205
R74 drain_left.n0 drain_left.t9 1.3205
R75 drain_left.n0 drain_left.t4 1.3205
R76 drain_left.n10 drain_left.t10 1.3205
R77 drain_left.n10 drain_left.t12 1.3205
R78 drain_left.n8 drain_left.t2 1.3205
R79 drain_left.n8 drain_left.t6 1.3205
R80 drain_left.n6 drain_left.t11 1.3205
R81 drain_left.n6 drain_left.t5 1.3205
R82 drain_left.n9 drain_left.n7 0.5005
R83 drain_left.n11 drain_left.n9 0.5005
R84 drain_left.n5 drain_left.n1 0.320154
R85 drain_left.n5 drain_left.n4 0.070154
R86 source.n7 source.t9 45.521
R87 source.n27 source.t2 45.5208
R88 source.n20 source.t24 45.5208
R89 source.n0 source.t20 45.5208
R90 source.n2 source.n1 44.201
R91 source.n4 source.n3 44.201
R92 source.n6 source.n5 44.201
R93 source.n9 source.n8 44.201
R94 source.n11 source.n10 44.201
R95 source.n13 source.n12 44.201
R96 source.n26 source.n25 44.2008
R97 source.n24 source.n23 44.2008
R98 source.n22 source.n21 44.2008
R99 source.n19 source.n18 44.2008
R100 source.n17 source.n16 44.2008
R101 source.n15 source.n14 44.2008
R102 source.n15 source.n13 24.5605
R103 source.n28 source.n0 18.5475
R104 source.n28 source.n27 5.51343
R105 source.n25 source.t4 1.3205
R106 source.n25 source.t11 1.3205
R107 source.n23 source.t10 1.3205
R108 source.n23 source.t3 1.3205
R109 source.n21 source.t7 1.3205
R110 source.n21 source.t8 1.3205
R111 source.n18 source.t17 1.3205
R112 source.n18 source.t15 1.3205
R113 source.n16 source.t21 1.3205
R114 source.n16 source.t23 1.3205
R115 source.n14 source.t16 1.3205
R116 source.n14 source.t25 1.3205
R117 source.n1 source.t19 1.3205
R118 source.n1 source.t14 1.3205
R119 source.n3 source.t18 1.3205
R120 source.n3 source.t27 1.3205
R121 source.n5 source.t22 1.3205
R122 source.n5 source.t26 1.3205
R123 source.n8 source.t6 1.3205
R124 source.n8 source.t5 1.3205
R125 source.n10 source.t12 1.3205
R126 source.n10 source.t1 1.3205
R127 source.n12 source.t13 1.3205
R128 source.n12 source.t0 1.3205
R129 source.n7 source.n6 0.720328
R130 source.n22 source.n20 0.720328
R131 source.n13 source.n11 0.5005
R132 source.n11 source.n9 0.5005
R133 source.n9 source.n7 0.5005
R134 source.n6 source.n4 0.5005
R135 source.n4 source.n2 0.5005
R136 source.n2 source.n0 0.5005
R137 source.n17 source.n15 0.5005
R138 source.n19 source.n17 0.5005
R139 source.n20 source.n19 0.5005
R140 source.n24 source.n22 0.5005
R141 source.n26 source.n24 0.5005
R142 source.n27 source.n26 0.5005
R143 source source.n28 0.188
R144 minus.n15 minus.t11 1606.37
R145 minus.n3 minus.t8 1606.37
R146 minus.n32 minus.t12 1606.37
R147 minus.n20 minus.t3 1606.37
R148 minus.n1 minus.t1 1571.32
R149 minus.n14 minus.t4 1571.32
R150 minus.n12 minus.t10 1571.32
R151 minus.n6 minus.t7 1571.32
R152 minus.n4 minus.t2 1571.32
R153 minus.n18 minus.t9 1571.32
R154 minus.n31 minus.t0 1571.32
R155 minus.n29 minus.t6 1571.32
R156 minus.n23 minus.t13 1571.32
R157 minus.n21 minus.t5 1571.32
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 61.346
R177 minus.n6 minus.n5 61.346
R178 minus.n23 minus.n22 61.346
R179 minus.n30 minus.n29 61.346
R180 minus.n15 minus.n14 49.6611
R181 minus.n4 minus.n3 49.6611
R182 minus.n21 minus.n20 49.6611
R183 minus.n32 minus.n31 49.6611
R184 minus.n34 minus.n16 37.5725
R185 minus.n14 minus.n13 23.3702
R186 minus.n5 minus.n4 23.3702
R187 minus.n22 minus.n21 23.3702
R188 minus.n31 minus.n30 23.3702
R189 minus.n12 minus.n11 11.6853
R190 minus.n7 minus.n6 11.6853
R191 minus.n24 minus.n23 11.6853
R192 minus.n29 minus.n28 11.6853
R193 minus.n34 minus.n33 6.45126
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t10 62.6996
R206 drain_right.n11 drain_right.t2 62.1998
R207 drain_right.n8 drain_right.n6 61.3796
R208 drain_right.n4 drain_right.n2 61.3796
R209 drain_right.n8 drain_right.n7 60.8798
R210 drain_right.n10 drain_right.n9 60.8798
R211 drain_right.n4 drain_right.n3 60.8796
R212 drain_right.n1 drain_right.n0 60.8796
R213 drain_right drain_right.n5 31.9616
R214 drain_right drain_right.n11 5.90322
R215 drain_right.n2 drain_right.t13 1.3205
R216 drain_right.n2 drain_right.t1 1.3205
R217 drain_right.n3 drain_right.t4 1.3205
R218 drain_right.n3 drain_right.t7 1.3205
R219 drain_right.n0 drain_right.t8 1.3205
R220 drain_right.n0 drain_right.t0 1.3205
R221 drain_right.n6 drain_right.t11 1.3205
R222 drain_right.n6 drain_right.t5 1.3205
R223 drain_right.n7 drain_right.t12 1.3205
R224 drain_right.n7 drain_right.t6 1.3205
R225 drain_right.n9 drain_right.t9 1.3205
R226 drain_right.n9 drain_right.t3 1.3205
R227 drain_right.n11 drain_right.n10 0.5005
R228 drain_right.n10 drain_right.n8 0.5005
R229 drain_right.n5 drain_right.n1 0.320154
R230 drain_right.n5 drain_right.n4 0.070154
C0 source drain_left 37.373f
C1 drain_right minus 5.67871f
C2 drain_right plus 0.315543f
C3 plus minus 5.76176f
C4 drain_right drain_left 0.842315f
C5 drain_right source 37.3593f
C6 minus drain_left 0.171605f
C7 plus drain_left 5.83343f
C8 minus source 5.17001f
C9 plus source 5.1849f
C10 drain_right a_n1644_n3888# 8.36913f
C11 drain_left a_n1644_n3888# 8.635071f
C12 source a_n1644_n3888# 7.149228f
C13 minus a_n1644_n3888# 6.588956f
C14 plus a_n1644_n3888# 8.81657f
C15 drain_right.t10 a_n1644_n3888# 4.47532f
C16 drain_right.t8 a_n1644_n3888# 0.387597f
C17 drain_right.t0 a_n1644_n3888# 0.387597f
C18 drain_right.n0 a_n1644_n3888# 3.50342f
C19 drain_right.n1 a_n1644_n3888# 0.775427f
C20 drain_right.t13 a_n1644_n3888# 0.387597f
C21 drain_right.t1 a_n1644_n3888# 0.387597f
C22 drain_right.n2 a_n1644_n3888# 3.50657f
C23 drain_right.t4 a_n1644_n3888# 0.387597f
C24 drain_right.t7 a_n1644_n3888# 0.387597f
C25 drain_right.n3 a_n1644_n3888# 3.50342f
C26 drain_right.n4 a_n1644_n3888# 0.721942f
C27 drain_right.n5 a_n1644_n3888# 1.68779f
C28 drain_right.t11 a_n1644_n3888# 0.387597f
C29 drain_right.t5 a_n1644_n3888# 0.387597f
C30 drain_right.n6 a_n1644_n3888# 3.50656f
C31 drain_right.t12 a_n1644_n3888# 0.387597f
C32 drain_right.t6 a_n1644_n3888# 0.387597f
C33 drain_right.n7 a_n1644_n3888# 3.50343f
C34 drain_right.n8 a_n1644_n3888# 0.756408f
C35 drain_right.t9 a_n1644_n3888# 0.387597f
C36 drain_right.t3 a_n1644_n3888# 0.387597f
C37 drain_right.n9 a_n1644_n3888# 3.50343f
C38 drain_right.n10 a_n1644_n3888# 0.373186f
C39 drain_right.t2 a_n1644_n3888# 4.47195f
C40 drain_right.n11 a_n1644_n3888# 0.691518f
C41 minus.n0 a_n1644_n3888# 0.053353f
C42 minus.t11 a_n1644_n3888# 0.569223f
C43 minus.t4 a_n1644_n3888# 0.564439f
C44 minus.t10 a_n1644_n3888# 0.564439f
C45 minus.t1 a_n1644_n3888# 0.564439f
C46 minus.n1 a_n1644_n3888# 0.237245f
C47 minus.n2 a_n1644_n3888# 0.1142f
C48 minus.t7 a_n1644_n3888# 0.564439f
C49 minus.t2 a_n1644_n3888# 0.564439f
C50 minus.t8 a_n1644_n3888# 0.569223f
C51 minus.n3 a_n1644_n3888# 0.234835f
C52 minus.n4 a_n1644_n3888# 0.219546f
C53 minus.n5 a_n1644_n3888# 0.02033f
C54 minus.n6 a_n1644_n3888# 0.219546f
C55 minus.n7 a_n1644_n3888# 0.02033f
C56 minus.n8 a_n1644_n3888# 0.053353f
C57 minus.n9 a_n1644_n3888# 0.053353f
C58 minus.n10 a_n1644_n3888# 0.053353f
C59 minus.n11 a_n1644_n3888# 0.02033f
C60 minus.n12 a_n1644_n3888# 0.219546f
C61 minus.n13 a_n1644_n3888# 0.02033f
C62 minus.n14 a_n1644_n3888# 0.219546f
C63 minus.n15 a_n1644_n3888# 0.234763f
C64 minus.n16 a_n1644_n3888# 1.99619f
C65 minus.n17 a_n1644_n3888# 0.053353f
C66 minus.t0 a_n1644_n3888# 0.564439f
C67 minus.t6 a_n1644_n3888# 0.564439f
C68 minus.t9 a_n1644_n3888# 0.564439f
C69 minus.n18 a_n1644_n3888# 0.237245f
C70 minus.n19 a_n1644_n3888# 0.1142f
C71 minus.t13 a_n1644_n3888# 0.564439f
C72 minus.t5 a_n1644_n3888# 0.564439f
C73 minus.t3 a_n1644_n3888# 0.569223f
C74 minus.n20 a_n1644_n3888# 0.234835f
C75 minus.n21 a_n1644_n3888# 0.219546f
C76 minus.n22 a_n1644_n3888# 0.02033f
C77 minus.n23 a_n1644_n3888# 0.219546f
C78 minus.n24 a_n1644_n3888# 0.02033f
C79 minus.n25 a_n1644_n3888# 0.053353f
C80 minus.n26 a_n1644_n3888# 0.053353f
C81 minus.n27 a_n1644_n3888# 0.053353f
C82 minus.n28 a_n1644_n3888# 0.02033f
C83 minus.n29 a_n1644_n3888# 0.219546f
C84 minus.n30 a_n1644_n3888# 0.02033f
C85 minus.n31 a_n1644_n3888# 0.219546f
C86 minus.t12 a_n1644_n3888# 0.569223f
C87 minus.n32 a_n1644_n3888# 0.234763f
C88 minus.n33 a_n1644_n3888# 0.342668f
C89 minus.n34 a_n1644_n3888# 2.4169f
C90 source.t20 a_n1644_n3888# 4.45207f
C91 source.n0 a_n1644_n3888# 2.0546f
C92 source.t19 a_n1644_n3888# 0.397272f
C93 source.t14 a_n1644_n3888# 0.397272f
C94 source.n1 a_n1644_n3888# 3.4897f
C95 source.n2 a_n1644_n3888# 0.438123f
C96 source.t18 a_n1644_n3888# 0.397272f
C97 source.t27 a_n1644_n3888# 0.397272f
C98 source.n3 a_n1644_n3888# 3.4897f
C99 source.n4 a_n1644_n3888# 0.438123f
C100 source.t22 a_n1644_n3888# 0.397272f
C101 source.t26 a_n1644_n3888# 0.397272f
C102 source.n5 a_n1644_n3888# 3.4897f
C103 source.n6 a_n1644_n3888# 0.461863f
C104 source.t9 a_n1644_n3888# 4.45208f
C105 source.n7 a_n1644_n3888# 0.582956f
C106 source.t6 a_n1644_n3888# 0.397272f
C107 source.t5 a_n1644_n3888# 0.397272f
C108 source.n8 a_n1644_n3888# 3.4897f
C109 source.n9 a_n1644_n3888# 0.438123f
C110 source.t12 a_n1644_n3888# 0.397272f
C111 source.t1 a_n1644_n3888# 0.397272f
C112 source.n10 a_n1644_n3888# 3.4897f
C113 source.n11 a_n1644_n3888# 0.438123f
C114 source.t13 a_n1644_n3888# 0.397272f
C115 source.t0 a_n1644_n3888# 0.397272f
C116 source.n12 a_n1644_n3888# 3.4897f
C117 source.n13 a_n1644_n3888# 2.54293f
C118 source.t16 a_n1644_n3888# 0.397272f
C119 source.t25 a_n1644_n3888# 0.397272f
C120 source.n14 a_n1644_n3888# 3.48969f
C121 source.n15 a_n1644_n3888# 2.54293f
C122 source.t21 a_n1644_n3888# 0.397272f
C123 source.t23 a_n1644_n3888# 0.397272f
C124 source.n16 a_n1644_n3888# 3.48969f
C125 source.n17 a_n1644_n3888# 0.438128f
C126 source.t17 a_n1644_n3888# 0.397272f
C127 source.t15 a_n1644_n3888# 0.397272f
C128 source.n18 a_n1644_n3888# 3.48969f
C129 source.n19 a_n1644_n3888# 0.438128f
C130 source.t24 a_n1644_n3888# 4.45207f
C131 source.n20 a_n1644_n3888# 0.582961f
C132 source.t7 a_n1644_n3888# 0.397272f
C133 source.t8 a_n1644_n3888# 0.397272f
C134 source.n21 a_n1644_n3888# 3.48969f
C135 source.n22 a_n1644_n3888# 0.461868f
C136 source.t10 a_n1644_n3888# 0.397272f
C137 source.t3 a_n1644_n3888# 0.397272f
C138 source.n23 a_n1644_n3888# 3.48969f
C139 source.n24 a_n1644_n3888# 0.438128f
C140 source.t4 a_n1644_n3888# 0.397272f
C141 source.t11 a_n1644_n3888# 0.397272f
C142 source.n25 a_n1644_n3888# 3.48969f
C143 source.n26 a_n1644_n3888# 0.438128f
C144 source.t2 a_n1644_n3888# 4.45207f
C145 source.n27 a_n1644_n3888# 0.74143f
C146 source.n28 a_n1644_n3888# 2.44786f
C147 drain_left.t3 a_n1644_n3888# 4.47243f
C148 drain_left.t9 a_n1644_n3888# 0.387347f
C149 drain_left.t4 a_n1644_n3888# 0.387347f
C150 drain_left.n0 a_n1644_n3888# 3.50116f
C151 drain_left.n1 a_n1644_n3888# 0.774927f
C152 drain_left.t0 a_n1644_n3888# 0.387347f
C153 drain_left.t8 a_n1644_n3888# 0.387347f
C154 drain_left.n2 a_n1644_n3888# 3.50431f
C155 drain_left.t7 a_n1644_n3888# 0.387347f
C156 drain_left.t1 a_n1644_n3888# 0.387347f
C157 drain_left.n3 a_n1644_n3888# 3.50116f
C158 drain_left.n4 a_n1644_n3888# 0.721476f
C159 drain_left.n5 a_n1644_n3888# 1.75494f
C160 drain_left.t13 a_n1644_n3888# 4.47243f
C161 drain_left.t11 a_n1644_n3888# 0.387347f
C162 drain_left.t5 a_n1644_n3888# 0.387347f
C163 drain_left.n6 a_n1644_n3888# 3.50116f
C164 drain_left.n7 a_n1644_n3888# 0.79154f
C165 drain_left.t2 a_n1644_n3888# 0.387347f
C166 drain_left.t6 a_n1644_n3888# 0.387347f
C167 drain_left.n8 a_n1644_n3888# 3.50116f
C168 drain_left.n9 a_n1644_n3888# 0.372945f
C169 drain_left.t10 a_n1644_n3888# 0.387347f
C170 drain_left.t12 a_n1644_n3888# 0.387347f
C171 drain_left.n10 a_n1644_n3888# 3.50115f
C172 drain_left.n11 a_n1644_n3888# 0.642692f
C173 plus.n0 a_n1644_n3888# 0.054022f
C174 plus.t13 a_n1644_n3888# 0.571511f
C175 plus.t8 a_n1644_n3888# 0.571511f
C176 plus.t0 a_n1644_n3888# 0.571511f
C177 plus.n1 a_n1644_n3888# 0.240217f
C178 plus.n2 a_n1644_n3888# 0.115631f
C179 plus.t9 a_n1644_n3888# 0.571511f
C180 plus.t1 a_n1644_n3888# 0.571511f
C181 plus.t5 a_n1644_n3888# 0.576355f
C182 plus.n3 a_n1644_n3888# 0.237777f
C183 plus.n4 a_n1644_n3888# 0.222296f
C184 plus.n5 a_n1644_n3888# 0.020585f
C185 plus.n6 a_n1644_n3888# 0.222296f
C186 plus.n7 a_n1644_n3888# 0.020585f
C187 plus.n8 a_n1644_n3888# 0.054022f
C188 plus.n9 a_n1644_n3888# 0.054022f
C189 plus.n10 a_n1644_n3888# 0.054022f
C190 plus.n11 a_n1644_n3888# 0.020585f
C191 plus.n12 a_n1644_n3888# 0.222296f
C192 plus.n13 a_n1644_n3888# 0.020585f
C193 plus.n14 a_n1644_n3888# 0.222296f
C194 plus.t7 a_n1644_n3888# 0.576355f
C195 plus.n15 a_n1644_n3888# 0.237705f
C196 plus.n16 a_n1644_n3888# 0.676451f
C197 plus.n17 a_n1644_n3888# 0.054022f
C198 plus.t11 a_n1644_n3888# 0.576355f
C199 plus.t2 a_n1644_n3888# 0.571511f
C200 plus.t6 a_n1644_n3888# 0.571511f
C201 plus.t4 a_n1644_n3888# 0.571511f
C202 plus.n18 a_n1644_n3888# 0.240217f
C203 plus.n19 a_n1644_n3888# 0.115631f
C204 plus.t10 a_n1644_n3888# 0.571511f
C205 plus.t12 a_n1644_n3888# 0.571511f
C206 plus.t3 a_n1644_n3888# 0.576355f
C207 plus.n20 a_n1644_n3888# 0.237777f
C208 plus.n21 a_n1644_n3888# 0.222296f
C209 plus.n22 a_n1644_n3888# 0.020585f
C210 plus.n23 a_n1644_n3888# 0.222296f
C211 plus.n24 a_n1644_n3888# 0.020585f
C212 plus.n25 a_n1644_n3888# 0.054022f
C213 plus.n26 a_n1644_n3888# 0.054022f
C214 plus.n27 a_n1644_n3888# 0.054022f
C215 plus.n28 a_n1644_n3888# 0.020585f
C216 plus.n29 a_n1644_n3888# 0.222296f
C217 plus.n30 a_n1644_n3888# 0.020585f
C218 plus.n31 a_n1644_n3888# 0.222296f
C219 plus.n32 a_n1644_n3888# 0.237705f
C220 plus.n33 a_n1644_n3888# 1.65826f
.ends

