* NGSPICE file created from diffpair565.ext - technology: sky130A

.subckt diffpair565 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t22 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X1 a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X2 source.t23 minus.t1 drain_right.t10 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 source.t4 plus.t0 drain_left.t11 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X4 a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X5 a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X6 drain_left.t10 plus.t1 source.t10 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X7 source.t13 minus.t2 drain_right.t9 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X8 source.t9 plus.t2 drain_left.t9 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X9 drain_right.t8 minus.t3 source.t20 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X10 drain_right.t7 minus.t4 source.t19 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source.t18 minus.t5 drain_right.t6 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 source.t12 minus.t6 drain_right.t5 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X13 drain_left.t8 plus.t3 source.t1 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X14 source.t2 plus.t4 drain_left.t7 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X15 drain_right.t4 minus.t7 source.t17 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X16 drain_right.t3 minus.t8 source.t16 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_left.t6 plus.t5 source.t3 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X18 drain_left.t5 plus.t6 source.t6 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 source.t15 minus.t9 drain_right.t2 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X20 drain_right.t1 minus.t10 source.t14 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X21 source.t8 plus.t7 drain_left.t4 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 source.t0 plus.t8 drain_left.t3 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X23 drain_left.t2 plus.t9 source.t7 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X24 drain_left.t1 plus.t10 source.t5 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X25 a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X26 source.t21 minus.t11 drain_right.t0 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 source.t11 plus.t11 drain_left.t0 a_n1626_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n13 minus.t9 3476.97
R1 minus.n2 minus.t3 3476.97
R2 minus.n28 minus.t10 3476.97
R3 minus.n17 minus.t1 3476.97
R4 minus.n12 minus.t4 3422.2
R5 minus.n10 minus.t6 3422.2
R6 minus.n3 minus.t7 3422.2
R7 minus.n4 minus.t2 3422.2
R8 minus.n27 minus.t5 3422.2
R9 minus.n25 minus.t0 3422.2
R10 minus.n19 minus.t11 3422.2
R11 minus.n18 minus.t8 3422.2
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 62.0763
R27 minus.n5 minus.n3 62.0763
R28 minus.n20 minus.n19 62.0763
R29 minus.n26 minus.n25 62.0763
R30 minus.n30 minus.n14 41.3831
R31 minus.n13 minus.n12 40.1672
R32 minus.n4 minus.n2 40.1672
R33 minus.n18 minus.n17 40.1672
R34 minus.n28 minus.n27 40.1672
R35 minus.n12 minus.n11 32.8641
R36 minus.n5 minus.n4 32.8641
R37 minus.n20 minus.n18 32.8641
R38 minus.n27 minus.n26 32.8641
R39 minus.n10 minus.n9 10.955
R40 minus.n3 minus.n1 10.955
R41 minus.n19 minus.n16 10.955
R42 minus.n25 minus.n24 10.955
R43 minus.n30 minus.n29 6.54217
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 source.n0 source.t7 44.6397
R54 source.n5 source.t2 44.6396
R55 source.n6 source.t20 44.6396
R56 source.n11 source.t15 44.6396
R57 source.n23 source.t14 44.6395
R58 source.n18 source.t23 44.6395
R59 source.n17 source.t1 44.6395
R60 source.n12 source.t4 44.6395
R61 source.n2 source.n1 43.1397
R62 source.n4 source.n3 43.1397
R63 source.n8 source.n7 43.1397
R64 source.n10 source.n9 43.1397
R65 source.n22 source.n21 43.1396
R66 source.n20 source.n19 43.1396
R67 source.n16 source.n15 43.1396
R68 source.n14 source.n13 43.1396
R69 source.n12 source.n11 27.9087
R70 source.n24 source.n0 22.3656
R71 source.n24 source.n23 5.5436
R72 source.n21 source.t22 1.5005
R73 source.n21 source.t18 1.5005
R74 source.n19 source.t16 1.5005
R75 source.n19 source.t21 1.5005
R76 source.n15 source.t10 1.5005
R77 source.n15 source.t0 1.5005
R78 source.n13 source.t3 1.5005
R79 source.n13 source.t9 1.5005
R80 source.n1 source.t6 1.5005
R81 source.n1 source.t11 1.5005
R82 source.n3 source.t5 1.5005
R83 source.n3 source.t8 1.5005
R84 source.n7 source.t17 1.5005
R85 source.n7 source.t13 1.5005
R86 source.n9 source.t19 1.5005
R87 source.n9 source.t12 1.5005
R88 source.n11 source.n10 0.560845
R89 source.n10 source.n8 0.560845
R90 source.n8 source.n6 0.560845
R91 source.n5 source.n4 0.560845
R92 source.n4 source.n2 0.560845
R93 source.n2 source.n0 0.560845
R94 source.n14 source.n12 0.560845
R95 source.n16 source.n14 0.560845
R96 source.n17 source.n16 0.560845
R97 source.n20 source.n18 0.560845
R98 source.n22 source.n20 0.560845
R99 source.n23 source.n22 0.560845
R100 source.n6 source.n5 0.470328
R101 source.n18 source.n17 0.470328
R102 source source.n24 0.188
R103 drain_right.n6 drain_right.n4 60.3788
R104 drain_right.n3 drain_right.n2 60.3234
R105 drain_right.n3 drain_right.n0 60.3234
R106 drain_right.n6 drain_right.n5 59.8185
R107 drain_right.n8 drain_right.n7 59.8185
R108 drain_right.n3 drain_right.n1 59.8184
R109 drain_right drain_right.n3 35.6762
R110 drain_right drain_right.n8 6.21356
R111 drain_right.n1 drain_right.t0 1.5005
R112 drain_right.n1 drain_right.t11 1.5005
R113 drain_right.n2 drain_right.t6 1.5005
R114 drain_right.n2 drain_right.t1 1.5005
R115 drain_right.n0 drain_right.t10 1.5005
R116 drain_right.n0 drain_right.t3 1.5005
R117 drain_right.n4 drain_right.t9 1.5005
R118 drain_right.n4 drain_right.t8 1.5005
R119 drain_right.n5 drain_right.t5 1.5005
R120 drain_right.n5 drain_right.t4 1.5005
R121 drain_right.n7 drain_right.t2 1.5005
R122 drain_right.n7 drain_right.t7 1.5005
R123 drain_right.n8 drain_right.n6 0.560845
R124 plus.n2 plus.t4 3476.97
R125 plus.n13 plus.t9 3476.97
R126 plus.n17 plus.t3 3476.97
R127 plus.n28 plus.t0 3476.97
R128 plus.n3 plus.t10 3422.2
R129 plus.n4 plus.t7 3422.2
R130 plus.n10 plus.t6 3422.2
R131 plus.n12 plus.t11 3422.2
R132 plus.n19 plus.t8 3422.2
R133 plus.n18 plus.t1 3422.2
R134 plus.n25 plus.t2 3422.2
R135 plus.n27 plus.t5 3422.2
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 62.0763
R151 plus.n11 plus.n10 62.0763
R152 plus.n26 plus.n25 62.0763
R153 plus.n20 plus.n18 62.0763
R154 plus.n3 plus.n2 40.1672
R155 plus.n13 plus.n12 40.1672
R156 plus.n28 plus.n27 40.1672
R157 plus.n19 plus.n17 40.1672
R158 plus.n5 plus.n3 32.8641
R159 plus.n12 plus.n11 32.8641
R160 plus.n27 plus.n26 32.8641
R161 plus.n20 plus.n19 32.8641
R162 plus plus.n29 32.2339
R163 plus plus.n14 15.2164
R164 plus.n4 plus.n1 10.955
R165 plus.n10 plus.n9 10.955
R166 plus.n25 plus.n24 10.955
R167 plus.n18 plus.n16 10.955
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 60.3788
R177 drain_left.n3 drain_left.n2 60.3234
R178 drain_left.n3 drain_left.n0 60.3234
R179 drain_left.n8 drain_left.n7 59.8185
R180 drain_left.n6 drain_left.n5 59.8185
R181 drain_left.n3 drain_left.n1 59.8184
R182 drain_left drain_left.n3 36.2294
R183 drain_left drain_left.n8 6.21356
R184 drain_left.n1 drain_left.t9 1.5005
R185 drain_left.n1 drain_left.t10 1.5005
R186 drain_left.n2 drain_left.t3 1.5005
R187 drain_left.n2 drain_left.t8 1.5005
R188 drain_left.n0 drain_left.t11 1.5005
R189 drain_left.n0 drain_left.t6 1.5005
R190 drain_left.n7 drain_left.t0 1.5005
R191 drain_left.n7 drain_left.t2 1.5005
R192 drain_left.n5 drain_left.t4 1.5005
R193 drain_left.n5 drain_left.t5 1.5005
R194 drain_left.n4 drain_left.t7 1.5005
R195 drain_left.n4 drain_left.t1 1.5005
R196 drain_left.n8 drain_left.n6 0.560845
C0 minus plus 6.64522f
C1 source drain_right 38.4464f
C2 source minus 3.56719f
C3 source plus 3.58123f
C4 drain_right drain_left 0.801529f
C5 minus drain_left 0.170585f
C6 plus drain_left 4.63566f
C7 minus drain_right 4.47917f
C8 plus drain_right 0.309819f
C9 source drain_left 38.4465f
C10 drain_right a_n1626_n4888# 7.19558f
C11 drain_left a_n1626_n4888# 7.43771f
C12 source a_n1626_n4888# 13.029402f
C13 minus a_n1626_n4888# 6.520351f
C14 plus a_n1626_n4888# 9.277451f
C15 drain_left.t11 a_n1626_n4888# 0.674985f
C16 drain_left.t6 a_n1626_n4888# 0.674985f
C17 drain_left.n0 a_n1626_n4888# 4.53467f
C18 drain_left.t9 a_n1626_n4888# 0.674985f
C19 drain_left.t10 a_n1626_n4888# 0.674985f
C20 drain_left.n1 a_n1626_n4888# 4.53176f
C21 drain_left.t3 a_n1626_n4888# 0.674985f
C22 drain_left.t8 a_n1626_n4888# 0.674985f
C23 drain_left.n2 a_n1626_n4888# 4.53467f
C24 drain_left.n3 a_n1626_n4888# 2.8521f
C25 drain_left.t7 a_n1626_n4888# 0.674985f
C26 drain_left.t1 a_n1626_n4888# 0.674985f
C27 drain_left.n4 a_n1626_n4888# 4.53501f
C28 drain_left.t4 a_n1626_n4888# 0.674985f
C29 drain_left.t5 a_n1626_n4888# 0.674985f
C30 drain_left.n5 a_n1626_n4888# 4.53175f
C31 drain_left.n6 a_n1626_n4888# 0.687404f
C32 drain_left.t0 a_n1626_n4888# 0.674985f
C33 drain_left.t2 a_n1626_n4888# 0.674985f
C34 drain_left.n7 a_n1626_n4888# 4.53175f
C35 drain_left.n8 a_n1626_n4888# 0.575049f
C36 plus.n0 a_n1626_n4888# 0.057623f
C37 plus.t11 a_n1626_n4888# 0.486883f
C38 plus.t6 a_n1626_n4888# 0.486883f
C39 plus.n1 a_n1626_n4888# 0.02178f
C40 plus.t4 a_n1626_n4888# 0.489886f
C41 plus.n2 a_n1626_n4888# 0.212161f
C42 plus.t10 a_n1626_n4888# 0.486883f
C43 plus.n3 a_n1626_n4888# 0.189747f
C44 plus.t7 a_n1626_n4888# 0.486883f
C45 plus.n4 a_n1626_n4888# 0.189747f
C46 plus.n5 a_n1626_n4888# 0.024445f
C47 plus.n6 a_n1626_n4888# 0.129373f
C48 plus.n7 a_n1626_n4888# 0.057623f
C49 plus.n8 a_n1626_n4888# 0.057623f
C50 plus.n9 a_n1626_n4888# 0.02178f
C51 plus.n10 a_n1626_n4888# 0.189747f
C52 plus.n11 a_n1626_n4888# 0.024445f
C53 plus.n12 a_n1626_n4888# 0.189747f
C54 plus.t9 a_n1626_n4888# 0.489886f
C55 plus.n13 a_n1626_n4888# 0.212077f
C56 plus.n14 a_n1626_n4888# 0.880553f
C57 plus.n15 a_n1626_n4888# 0.057623f
C58 plus.t0 a_n1626_n4888# 0.489886f
C59 plus.t5 a_n1626_n4888# 0.486883f
C60 plus.t2 a_n1626_n4888# 0.486883f
C61 plus.n16 a_n1626_n4888# 0.02178f
C62 plus.t3 a_n1626_n4888# 0.489886f
C63 plus.n17 a_n1626_n4888# 0.212161f
C64 plus.t1 a_n1626_n4888# 0.486883f
C65 plus.n18 a_n1626_n4888# 0.189747f
C66 plus.t8 a_n1626_n4888# 0.486883f
C67 plus.n19 a_n1626_n4888# 0.189747f
C68 plus.n20 a_n1626_n4888# 0.024445f
C69 plus.n21 a_n1626_n4888# 0.129373f
C70 plus.n22 a_n1626_n4888# 0.057623f
C71 plus.n23 a_n1626_n4888# 0.057623f
C72 plus.n24 a_n1626_n4888# 0.02178f
C73 plus.n25 a_n1626_n4888# 0.189747f
C74 plus.n26 a_n1626_n4888# 0.024445f
C75 plus.n27 a_n1626_n4888# 0.189747f
C76 plus.n28 a_n1626_n4888# 0.212077f
C77 plus.n29 a_n1626_n4888# 1.971f
C78 drain_right.t10 a_n1626_n4888# 0.675146f
C79 drain_right.t3 a_n1626_n4888# 0.675146f
C80 drain_right.n0 a_n1626_n4888# 4.53575f
C81 drain_right.t0 a_n1626_n4888# 0.675146f
C82 drain_right.t11 a_n1626_n4888# 0.675146f
C83 drain_right.n1 a_n1626_n4888# 4.53284f
C84 drain_right.t6 a_n1626_n4888# 0.675146f
C85 drain_right.t1 a_n1626_n4888# 0.675146f
C86 drain_right.n2 a_n1626_n4888# 4.53575f
C87 drain_right.n3 a_n1626_n4888# 2.79391f
C88 drain_right.t9 a_n1626_n4888# 0.675146f
C89 drain_right.t8 a_n1626_n4888# 0.675146f
C90 drain_right.n4 a_n1626_n4888# 4.5361f
C91 drain_right.t5 a_n1626_n4888# 0.675146f
C92 drain_right.t4 a_n1626_n4888# 0.675146f
C93 drain_right.n5 a_n1626_n4888# 4.53284f
C94 drain_right.n6 a_n1626_n4888# 0.687569f
C95 drain_right.t2 a_n1626_n4888# 0.675146f
C96 drain_right.t7 a_n1626_n4888# 0.675146f
C97 drain_right.n7 a_n1626_n4888# 4.53284f
C98 drain_right.n8 a_n1626_n4888# 0.575186f
C99 source.t7 a_n1626_n4888# 4.32706f
C100 source.n0 a_n1626_n4888# 1.7568f
C101 source.t6 a_n1626_n4888# 0.532059f
C102 source.t11 a_n1626_n4888# 0.532059f
C103 source.n1 a_n1626_n4888# 3.50131f
C104 source.n2 a_n1626_n4888# 0.308391f
C105 source.t5 a_n1626_n4888# 0.532059f
C106 source.t8 a_n1626_n4888# 0.532059f
C107 source.n3 a_n1626_n4888# 3.50131f
C108 source.n4 a_n1626_n4888# 0.308391f
C109 source.t2 a_n1626_n4888# 4.32707f
C110 source.n5 a_n1626_n4888# 0.433858f
C111 source.t20 a_n1626_n4888# 4.32707f
C112 source.n6 a_n1626_n4888# 0.433858f
C113 source.t17 a_n1626_n4888# 0.532059f
C114 source.t13 a_n1626_n4888# 0.532059f
C115 source.n7 a_n1626_n4888# 3.50131f
C116 source.n8 a_n1626_n4888# 0.308391f
C117 source.t19 a_n1626_n4888# 0.532059f
C118 source.t12 a_n1626_n4888# 0.532059f
C119 source.n9 a_n1626_n4888# 3.50131f
C120 source.n10 a_n1626_n4888# 0.308391f
C121 source.t15 a_n1626_n4888# 4.32707f
C122 source.n11 a_n1626_n4888# 2.15107f
C123 source.t4 a_n1626_n4888# 4.32705f
C124 source.n12 a_n1626_n4888# 2.15109f
C125 source.t3 a_n1626_n4888# 0.532059f
C126 source.t9 a_n1626_n4888# 0.532059f
C127 source.n13 a_n1626_n4888# 3.50132f
C128 source.n14 a_n1626_n4888# 0.308384f
C129 source.t10 a_n1626_n4888# 0.532059f
C130 source.t0 a_n1626_n4888# 0.532059f
C131 source.n15 a_n1626_n4888# 3.50132f
C132 source.n16 a_n1626_n4888# 0.308384f
C133 source.t1 a_n1626_n4888# 4.32705f
C134 source.n17 a_n1626_n4888# 0.43388f
C135 source.t23 a_n1626_n4888# 4.32705f
C136 source.n18 a_n1626_n4888# 0.43388f
C137 source.t16 a_n1626_n4888# 0.532059f
C138 source.t21 a_n1626_n4888# 0.532059f
C139 source.n19 a_n1626_n4888# 3.50132f
C140 source.n20 a_n1626_n4888# 0.308384f
C141 source.t22 a_n1626_n4888# 0.532059f
C142 source.t18 a_n1626_n4888# 0.532059f
C143 source.n21 a_n1626_n4888# 3.50132f
C144 source.n22 a_n1626_n4888# 0.308384f
C145 source.t14 a_n1626_n4888# 4.32705f
C146 source.n23 a_n1626_n4888# 0.560291f
C147 source.n24 a_n1626_n4888# 2.00088f
C148 minus.n0 a_n1626_n4888# 0.056787f
C149 minus.t9 a_n1626_n4888# 0.482775f
C150 minus.t4 a_n1626_n4888# 0.479816f
C151 minus.t6 a_n1626_n4888# 0.479816f
C152 minus.n1 a_n1626_n4888# 0.021464f
C153 minus.t3 a_n1626_n4888# 0.482775f
C154 minus.n2 a_n1626_n4888# 0.209081f
C155 minus.t7 a_n1626_n4888# 0.479816f
C156 minus.n3 a_n1626_n4888# 0.186993f
C157 minus.t2 a_n1626_n4888# 0.479816f
C158 minus.n4 a_n1626_n4888# 0.186993f
C159 minus.n5 a_n1626_n4888# 0.02409f
C160 minus.n6 a_n1626_n4888# 0.127495f
C161 minus.n7 a_n1626_n4888# 0.056787f
C162 minus.n8 a_n1626_n4888# 0.056787f
C163 minus.n9 a_n1626_n4888# 0.021464f
C164 minus.n10 a_n1626_n4888# 0.186993f
C165 minus.n11 a_n1626_n4888# 0.02409f
C166 minus.n12 a_n1626_n4888# 0.186993f
C167 minus.n13 a_n1626_n4888# 0.208998f
C168 minus.n14 a_n1626_n4888# 2.46214f
C169 minus.n15 a_n1626_n4888# 0.056787f
C170 minus.t5 a_n1626_n4888# 0.479816f
C171 minus.t0 a_n1626_n4888# 0.479816f
C172 minus.n16 a_n1626_n4888# 0.021464f
C173 minus.t1 a_n1626_n4888# 0.482775f
C174 minus.n17 a_n1626_n4888# 0.209081f
C175 minus.t8 a_n1626_n4888# 0.479816f
C176 minus.n18 a_n1626_n4888# 0.186993f
C177 minus.t11 a_n1626_n4888# 0.479816f
C178 minus.n19 a_n1626_n4888# 0.186993f
C179 minus.n20 a_n1626_n4888# 0.02409f
C180 minus.n21 a_n1626_n4888# 0.127495f
C181 minus.n22 a_n1626_n4888# 0.056787f
C182 minus.n23 a_n1626_n4888# 0.056787f
C183 minus.n24 a_n1626_n4888# 0.021464f
C184 minus.n25 a_n1626_n4888# 0.186993f
C185 minus.n26 a_n1626_n4888# 0.02409f
C186 minus.n27 a_n1626_n4888# 0.186993f
C187 minus.t10 a_n1626_n4888# 0.482775f
C188 minus.n28 a_n1626_n4888# 0.208998f
C189 minus.n29 a_n1626_n4888# 0.376887f
C190 minus.n30 a_n1626_n4888# 2.94403f
.ends

