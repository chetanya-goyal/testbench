* NGSPICE file created from diffpair386.ext - technology: sky130A

.subckt diffpair386 minus drain_right drain_left source plus
X0 a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X1 drain_left.t13 plus.t0 source.t12 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X2 drain_left.t12 plus.t1 source.t19 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X3 source.t7 minus.t0 drain_right.t13 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X4 drain_left.t11 plus.t2 source.t13 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X5 drain_left.t10 plus.t3 source.t18 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X6 source.t14 plus.t4 drain_left.t9 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X7 drain_left.t8 plus.t5 source.t20 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X8 a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X9 drain_right.t12 minus.t1 source.t0 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X10 drain_right.t11 minus.t2 source.t1 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X11 drain_left.t7 plus.t6 source.t21 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X12 drain_right.t10 minus.t3 source.t2 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X13 source.t16 plus.t7 drain_left.t6 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X14 source.t24 plus.t8 drain_left.t5 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X15 source.t6 minus.t4 drain_right.t9 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X16 drain_right.t8 minus.t5 source.t9 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X17 a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X18 drain_right.t7 minus.t6 source.t27 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X19 source.t22 plus.t9 drain_left.t4 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X20 drain_left.t3 plus.t10 source.t17 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X21 drain_right.t6 minus.t7 source.t5 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X22 source.t15 plus.t11 drain_left.t2 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X23 source.t4 minus.t8 drain_right.t5 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X24 drain_right.t4 minus.t9 source.t11 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X25 source.t23 plus.t12 drain_left.t1 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X26 drain_left.t0 plus.t13 source.t25 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X27 source.t3 minus.t10 drain_right.t3 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X28 source.t8 minus.t11 drain_right.t2 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X29 source.t10 minus.t12 drain_right.t1 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X30 drain_right.t0 minus.t13 source.t26 a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X31 a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# a_n2364_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
R0 plus.n5 plus.t3 389.822
R1 plus.n27 plus.t10 389.822
R2 plus.n20 plus.t0 365.976
R3 plus.n18 plus.t8 365.976
R4 plus.n2 plus.t2 365.976
R5 plus.n12 plus.t7 365.976
R6 plus.n4 plus.t1 365.976
R7 plus.n6 plus.t9 365.976
R8 plus.n42 plus.t13 365.976
R9 plus.n40 plus.t12 365.976
R10 plus.n24 plus.t5 365.976
R11 plus.n34 plus.t4 365.976
R12 plus.n26 plus.t6 365.976
R13 plus.n28 plus.t11 365.976
R14 plus.n8 plus.n7 161.3
R15 plus.n9 plus.n4 161.3
R16 plus.n11 plus.n10 161.3
R17 plus.n12 plus.n3 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n15 plus.n2 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n18 plus.n1 161.3
R22 plus.n19 plus.n0 161.3
R23 plus.n21 plus.n20 161.3
R24 plus.n30 plus.n29 161.3
R25 plus.n31 plus.n26 161.3
R26 plus.n33 plus.n32 161.3
R27 plus.n34 plus.n25 161.3
R28 plus.n36 plus.n35 161.3
R29 plus.n37 plus.n24 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n40 plus.n23 161.3
R32 plus.n41 plus.n22 161.3
R33 plus.n43 plus.n42 161.3
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus plus.n43 30.9706
R39 plus.n18 plus.n17 30.6732
R40 plus.n7 plus.n6 30.6732
R41 plus.n40 plus.n39 30.6732
R42 plus.n29 plus.n28 30.6732
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus.n19 plus.n18 13.146
R58 plus.n41 plus.n40 13.146
R59 plus plus.n21 11.1577
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n7 source.t9 51.0588
R79 source.n27 source.t27 51.0586
R80 source.n20 source.t17 51.0586
R81 source.n0 source.t12 51.0586
R82 source.n2 source.n1 48.8588
R83 source.n4 source.n3 48.8588
R84 source.n6 source.n5 48.8588
R85 source.n9 source.n8 48.8588
R86 source.n11 source.n10 48.8588
R87 source.n13 source.n12 48.8588
R88 source.n26 source.n25 48.8586
R89 source.n24 source.n23 48.8586
R90 source.n22 source.n21 48.8586
R91 source.n19 source.n18 48.8586
R92 source.n17 source.n16 48.8586
R93 source.n15 source.n14 48.8586
R94 source.n15 source.n13 20.7909
R95 source.n28 source.n0 14.196
R96 source.n28 source.n27 5.7074
R97 source.n25 source.t11 2.2005
R98 source.n25 source.t6 2.2005
R99 source.n23 source.t5 2.2005
R100 source.n23 source.t4 2.2005
R101 source.n21 source.t26 2.2005
R102 source.n21 source.t10 2.2005
R103 source.n18 source.t21 2.2005
R104 source.n18 source.t15 2.2005
R105 source.n16 source.t20 2.2005
R106 source.n16 source.t14 2.2005
R107 source.n14 source.t25 2.2005
R108 source.n14 source.t23 2.2005
R109 source.n1 source.t13 2.2005
R110 source.n1 source.t24 2.2005
R111 source.n3 source.t19 2.2005
R112 source.n3 source.t16 2.2005
R113 source.n5 source.t18 2.2005
R114 source.n5 source.t22 2.2005
R115 source.n8 source.t2 2.2005
R116 source.n8 source.t7 2.2005
R117 source.n10 source.t1 2.2005
R118 source.n10 source.t3 2.2005
R119 source.n12 source.t0 2.2005
R120 source.n12 source.t8 2.2005
R121 source.n7 source.n6 0.914293
R122 source.n22 source.n20 0.914293
R123 source.n13 source.n11 0.888431
R124 source.n11 source.n9 0.888431
R125 source.n9 source.n7 0.888431
R126 source.n6 source.n4 0.888431
R127 source.n4 source.n2 0.888431
R128 source.n2 source.n0 0.888431
R129 source.n17 source.n15 0.888431
R130 source.n19 source.n17 0.888431
R131 source.n20 source.n19 0.888431
R132 source.n24 source.n22 0.888431
R133 source.n26 source.n24 0.888431
R134 source.n27 source.n26 0.888431
R135 source source.n28 0.188
R136 drain_left.n7 drain_left.t10 68.6255
R137 drain_left.n1 drain_left.t0 68.6253
R138 drain_left.n4 drain_left.n2 66.4253
R139 drain_left.n9 drain_left.n8 65.5376
R140 drain_left.n7 drain_left.n6 65.5376
R141 drain_left.n11 drain_left.n10 65.5374
R142 drain_left.n4 drain_left.n3 65.5373
R143 drain_left.n1 drain_left.n0 65.5373
R144 drain_left drain_left.n5 30.2
R145 drain_left drain_left.n11 6.54115
R146 drain_left.n2 drain_left.t2 2.2005
R147 drain_left.n2 drain_left.t3 2.2005
R148 drain_left.n3 drain_left.t9 2.2005
R149 drain_left.n3 drain_left.t7 2.2005
R150 drain_left.n0 drain_left.t1 2.2005
R151 drain_left.n0 drain_left.t8 2.2005
R152 drain_left.n10 drain_left.t5 2.2005
R153 drain_left.n10 drain_left.t13 2.2005
R154 drain_left.n8 drain_left.t6 2.2005
R155 drain_left.n8 drain_left.t11 2.2005
R156 drain_left.n6 drain_left.t4 2.2005
R157 drain_left.n6 drain_left.t12 2.2005
R158 drain_left.n9 drain_left.n7 0.888431
R159 drain_left.n11 drain_left.n9 0.888431
R160 drain_left.n5 drain_left.n1 0.611102
R161 drain_left.n5 drain_left.n4 0.167137
R162 minus.n5 minus.t5 389.822
R163 minus.n27 minus.t13 389.822
R164 minus.n6 minus.t0 365.976
R165 minus.n8 minus.t3 365.976
R166 minus.n12 minus.t10 365.976
R167 minus.n14 minus.t2 365.976
R168 minus.n18 minus.t11 365.976
R169 minus.n20 minus.t1 365.976
R170 minus.n28 minus.t12 365.976
R171 minus.n30 minus.t7 365.976
R172 minus.n34 minus.t8 365.976
R173 minus.n36 minus.t9 365.976
R174 minus.n40 minus.t4 365.976
R175 minus.n42 minus.t6 365.976
R176 minus.n21 minus.n20 161.3
R177 minus.n19 minus.n0 161.3
R178 minus.n18 minus.n17 161.3
R179 minus.n16 minus.n1 161.3
R180 minus.n15 minus.n14 161.3
R181 minus.n13 minus.n2 161.3
R182 minus.n12 minus.n11 161.3
R183 minus.n10 minus.n3 161.3
R184 minus.n9 minus.n8 161.3
R185 minus.n7 minus.n4 161.3
R186 minus.n43 minus.n42 161.3
R187 minus.n41 minus.n22 161.3
R188 minus.n40 minus.n39 161.3
R189 minus.n38 minus.n23 161.3
R190 minus.n37 minus.n36 161.3
R191 minus.n35 minus.n24 161.3
R192 minus.n34 minus.n33 161.3
R193 minus.n32 minus.n25 161.3
R194 minus.n31 minus.n30 161.3
R195 minus.n29 minus.n26 161.3
R196 minus.n5 minus.n4 44.9119
R197 minus.n27 minus.n26 44.9119
R198 minus.n44 minus.n21 35.9532
R199 minus.n20 minus.n19 35.055
R200 minus.n42 minus.n41 35.055
R201 minus.n7 minus.n6 30.6732
R202 minus.n18 minus.n1 30.6732
R203 minus.n29 minus.n28 30.6732
R204 minus.n40 minus.n23 30.6732
R205 minus.n8 minus.n3 26.2914
R206 minus.n14 minus.n13 26.2914
R207 minus.n30 minus.n25 26.2914
R208 minus.n36 minus.n35 26.2914
R209 minus.n12 minus.n3 21.9096
R210 minus.n13 minus.n12 21.9096
R211 minus.n34 minus.n25 21.9096
R212 minus.n35 minus.n34 21.9096
R213 minus.n6 minus.n5 17.739
R214 minus.n28 minus.n27 17.739
R215 minus.n8 minus.n7 17.5278
R216 minus.n14 minus.n1 17.5278
R217 minus.n30 minus.n29 17.5278
R218 minus.n36 minus.n23 17.5278
R219 minus.n19 minus.n18 13.146
R220 minus.n41 minus.n40 13.146
R221 minus.n44 minus.n43 6.65012
R222 minus.n21 minus.n0 0.189894
R223 minus.n17 minus.n0 0.189894
R224 minus.n17 minus.n16 0.189894
R225 minus.n16 minus.n15 0.189894
R226 minus.n15 minus.n2 0.189894
R227 minus.n11 minus.n2 0.189894
R228 minus.n11 minus.n10 0.189894
R229 minus.n10 minus.n9 0.189894
R230 minus.n9 minus.n4 0.189894
R231 minus.n31 minus.n26 0.189894
R232 minus.n32 minus.n31 0.189894
R233 minus.n33 minus.n32 0.189894
R234 minus.n33 minus.n24 0.189894
R235 minus.n37 minus.n24 0.189894
R236 minus.n38 minus.n37 0.189894
R237 minus.n39 minus.n38 0.189894
R238 minus.n39 minus.n22 0.189894
R239 minus.n43 minus.n22 0.189894
R240 minus minus.n44 0.188
R241 drain_right.n1 drain_right.t0 68.6253
R242 drain_right.n11 drain_right.t12 67.7376
R243 drain_right.n8 drain_right.n6 66.4254
R244 drain_right.n4 drain_right.n2 66.4253
R245 drain_right.n8 drain_right.n7 65.5376
R246 drain_right.n10 drain_right.n9 65.5376
R247 drain_right.n4 drain_right.n3 65.5373
R248 drain_right.n1 drain_right.n0 65.5373
R249 drain_right drain_right.n5 29.6467
R250 drain_right drain_right.n11 6.09718
R251 drain_right.n2 drain_right.t9 2.2005
R252 drain_right.n2 drain_right.t7 2.2005
R253 drain_right.n3 drain_right.t5 2.2005
R254 drain_right.n3 drain_right.t4 2.2005
R255 drain_right.n0 drain_right.t1 2.2005
R256 drain_right.n0 drain_right.t6 2.2005
R257 drain_right.n6 drain_right.t13 2.2005
R258 drain_right.n6 drain_right.t8 2.2005
R259 drain_right.n7 drain_right.t3 2.2005
R260 drain_right.n7 drain_right.t10 2.2005
R261 drain_right.n9 drain_right.t2 2.2005
R262 drain_right.n9 drain_right.t11 2.2005
R263 drain_right.n11 drain_right.n10 0.888431
R264 drain_right.n10 drain_right.n8 0.888431
R265 drain_right.n5 drain_right.n1 0.611102
R266 drain_right.n5 drain_right.n4 0.167137
C0 drain_left drain_right 1.23294f
C1 drain_left source 14.789001f
C2 plus minus 5.53692f
C3 drain_right source 14.784599f
C4 drain_left plus 7.16595f
C5 drain_left minus 0.172675f
C6 plus drain_right 0.390564f
C7 plus source 7.02972f
C8 minus drain_right 6.93453f
C9 minus source 7.0153f
C10 drain_right a_n2364_n2688# 6.71514f
C11 drain_left a_n2364_n2688# 7.07732f
C12 source a_n2364_n2688# 5.586095f
C13 minus a_n2364_n2688# 9.180644f
C14 plus a_n2364_n2688# 10.75873f
C15 drain_right.t0 a_n2364_n2688# 1.98039f
C16 drain_right.t1 a_n2364_n2688# 0.177476f
C17 drain_right.t6 a_n2364_n2688# 0.177476f
C18 drain_right.n0 a_n2364_n2688# 1.55232f
C19 drain_right.n1 a_n2364_n2688# 0.658611f
C20 drain_right.t9 a_n2364_n2688# 0.177476f
C21 drain_right.t7 a_n2364_n2688# 0.177476f
C22 drain_right.n2 a_n2364_n2688# 1.55703f
C23 drain_right.t5 a_n2364_n2688# 0.177476f
C24 drain_right.t4 a_n2364_n2688# 0.177476f
C25 drain_right.n3 a_n2364_n2688# 1.55232f
C26 drain_right.n4 a_n2364_n2688# 0.636167f
C27 drain_right.n5 a_n2364_n2688# 1.15794f
C28 drain_right.t13 a_n2364_n2688# 0.177476f
C29 drain_right.t8 a_n2364_n2688# 0.177476f
C30 drain_right.n6 a_n2364_n2688# 1.55703f
C31 drain_right.t3 a_n2364_n2688# 0.177476f
C32 drain_right.t10 a_n2364_n2688# 0.177476f
C33 drain_right.n7 a_n2364_n2688# 1.55232f
C34 drain_right.n8 a_n2364_n2688# 0.690693f
C35 drain_right.t2 a_n2364_n2688# 0.177476f
C36 drain_right.t11 a_n2364_n2688# 0.177476f
C37 drain_right.n9 a_n2364_n2688# 1.55232f
C38 drain_right.n10 a_n2364_n2688# 0.342675f
C39 drain_right.t12 a_n2364_n2688# 1.97597f
C40 drain_right.n11 a_n2364_n2688# 0.571045f
C41 minus.n0 a_n2364_n2688# 0.041151f
C42 minus.n1 a_n2364_n2688# 0.009338f
C43 minus.t11 a_n2364_n2688# 0.743497f
C44 minus.n2 a_n2364_n2688# 0.041151f
C45 minus.n3 a_n2364_n2688# 0.009338f
C46 minus.t10 a_n2364_n2688# 0.743497f
C47 minus.n4 a_n2364_n2688# 0.173387f
C48 minus.t5 a_n2364_n2688# 0.762609f
C49 minus.n5 a_n2364_n2688# 0.296845f
C50 minus.t0 a_n2364_n2688# 0.743497f
C51 minus.n6 a_n2364_n2688# 0.317478f
C52 minus.n7 a_n2364_n2688# 0.009338f
C53 minus.t3 a_n2364_n2688# 0.743497f
C54 minus.n8 a_n2364_n2688# 0.31238f
C55 minus.n9 a_n2364_n2688# 0.041151f
C56 minus.n10 a_n2364_n2688# 0.041151f
C57 minus.n11 a_n2364_n2688# 0.041151f
C58 minus.n12 a_n2364_n2688# 0.31238f
C59 minus.n13 a_n2364_n2688# 0.009338f
C60 minus.t2 a_n2364_n2688# 0.743497f
C61 minus.n14 a_n2364_n2688# 0.31238f
C62 minus.n15 a_n2364_n2688# 0.041151f
C63 minus.n16 a_n2364_n2688# 0.041151f
C64 minus.n17 a_n2364_n2688# 0.041151f
C65 minus.n18 a_n2364_n2688# 0.31238f
C66 minus.n19 a_n2364_n2688# 0.009338f
C67 minus.t1 a_n2364_n2688# 0.743497f
C68 minus.n20 a_n2364_n2688# 0.310858f
C69 minus.n21 a_n2364_n2688# 1.44401f
C70 minus.n22 a_n2364_n2688# 0.041151f
C71 minus.n23 a_n2364_n2688# 0.009338f
C72 minus.n24 a_n2364_n2688# 0.041151f
C73 minus.n25 a_n2364_n2688# 0.009338f
C74 minus.n26 a_n2364_n2688# 0.173387f
C75 minus.t13 a_n2364_n2688# 0.762609f
C76 minus.n27 a_n2364_n2688# 0.296845f
C77 minus.t12 a_n2364_n2688# 0.743497f
C78 minus.n28 a_n2364_n2688# 0.317478f
C79 minus.n29 a_n2364_n2688# 0.009338f
C80 minus.t7 a_n2364_n2688# 0.743497f
C81 minus.n30 a_n2364_n2688# 0.31238f
C82 minus.n31 a_n2364_n2688# 0.041151f
C83 minus.n32 a_n2364_n2688# 0.041151f
C84 minus.n33 a_n2364_n2688# 0.041151f
C85 minus.t8 a_n2364_n2688# 0.743497f
C86 minus.n34 a_n2364_n2688# 0.31238f
C87 minus.n35 a_n2364_n2688# 0.009338f
C88 minus.t9 a_n2364_n2688# 0.743497f
C89 minus.n36 a_n2364_n2688# 0.31238f
C90 minus.n37 a_n2364_n2688# 0.041151f
C91 minus.n38 a_n2364_n2688# 0.041151f
C92 minus.n39 a_n2364_n2688# 0.041151f
C93 minus.t4 a_n2364_n2688# 0.743497f
C94 minus.n40 a_n2364_n2688# 0.31238f
C95 minus.n41 a_n2364_n2688# 0.009338f
C96 minus.t6 a_n2364_n2688# 0.743497f
C97 minus.n42 a_n2364_n2688# 0.310858f
C98 minus.n43 a_n2364_n2688# 0.283487f
C99 minus.n44 a_n2364_n2688# 1.75032f
C100 drain_left.t0 a_n2364_n2688# 1.99878f
C101 drain_left.t1 a_n2364_n2688# 0.179123f
C102 drain_left.t8 a_n2364_n2688# 0.179123f
C103 drain_left.n0 a_n2364_n2688# 1.56673f
C104 drain_left.n1 a_n2364_n2688# 0.664726f
C105 drain_left.t2 a_n2364_n2688# 0.179123f
C106 drain_left.t3 a_n2364_n2688# 0.179123f
C107 drain_left.n2 a_n2364_n2688# 1.57149f
C108 drain_left.t9 a_n2364_n2688# 0.179123f
C109 drain_left.t7 a_n2364_n2688# 0.179123f
C110 drain_left.n3 a_n2364_n2688# 1.56673f
C111 drain_left.n4 a_n2364_n2688# 0.642073f
C112 drain_left.n5 a_n2364_n2688# 1.22009f
C113 drain_left.t10 a_n2364_n2688# 1.99878f
C114 drain_left.t4 a_n2364_n2688# 0.179123f
C115 drain_left.t12 a_n2364_n2688# 0.179123f
C116 drain_left.n6 a_n2364_n2688# 1.56673f
C117 drain_left.n7 a_n2364_n2688# 0.68627f
C118 drain_left.t6 a_n2364_n2688# 0.179123f
C119 drain_left.t11 a_n2364_n2688# 0.179123f
C120 drain_left.n8 a_n2364_n2688# 1.56673f
C121 drain_left.n9 a_n2364_n2688# 0.345857f
C122 drain_left.t5 a_n2364_n2688# 0.179123f
C123 drain_left.t13 a_n2364_n2688# 0.179123f
C124 drain_left.n10 a_n2364_n2688# 1.56673f
C125 drain_left.n11 a_n2364_n2688# 0.568633f
C126 source.t12 a_n2364_n2688# 2.04249f
C127 source.n0 a_n2364_n2688# 1.22452f
C128 source.t13 a_n2364_n2688# 0.191541f
C129 source.t24 a_n2364_n2688# 0.191541f
C130 source.n1 a_n2364_n2688# 1.60345f
C131 source.n2 a_n2364_n2688# 0.405119f
C132 source.t19 a_n2364_n2688# 0.191541f
C133 source.t16 a_n2364_n2688# 0.191541f
C134 source.n3 a_n2364_n2688# 1.60345f
C135 source.n4 a_n2364_n2688# 0.405119f
C136 source.t18 a_n2364_n2688# 0.191541f
C137 source.t22 a_n2364_n2688# 0.191541f
C138 source.n5 a_n2364_n2688# 1.60345f
C139 source.n6 a_n2364_n2688# 0.407363f
C140 source.t9 a_n2364_n2688# 2.04249f
C141 source.n7 a_n2364_n2688# 0.490708f
C142 source.t2 a_n2364_n2688# 0.191541f
C143 source.t7 a_n2364_n2688# 0.191541f
C144 source.n8 a_n2364_n2688# 1.60345f
C145 source.n9 a_n2364_n2688# 0.405119f
C146 source.t1 a_n2364_n2688# 0.191541f
C147 source.t3 a_n2364_n2688# 0.191541f
C148 source.n10 a_n2364_n2688# 1.60345f
C149 source.n11 a_n2364_n2688# 0.405119f
C150 source.t0 a_n2364_n2688# 0.191541f
C151 source.t8 a_n2364_n2688# 0.191541f
C152 source.n12 a_n2364_n2688# 1.60345f
C153 source.n13 a_n2364_n2688# 1.61936f
C154 source.t25 a_n2364_n2688# 0.191541f
C155 source.t23 a_n2364_n2688# 0.191541f
C156 source.n14 a_n2364_n2688# 1.60345f
C157 source.n15 a_n2364_n2688# 1.61936f
C158 source.t20 a_n2364_n2688# 0.191541f
C159 source.t14 a_n2364_n2688# 0.191541f
C160 source.n16 a_n2364_n2688# 1.60345f
C161 source.n17 a_n2364_n2688# 0.405123f
C162 source.t21 a_n2364_n2688# 0.191541f
C163 source.t15 a_n2364_n2688# 0.191541f
C164 source.n18 a_n2364_n2688# 1.60345f
C165 source.n19 a_n2364_n2688# 0.405123f
C166 source.t17 a_n2364_n2688# 2.04249f
C167 source.n20 a_n2364_n2688# 0.490713f
C168 source.t26 a_n2364_n2688# 0.191541f
C169 source.t10 a_n2364_n2688# 0.191541f
C170 source.n21 a_n2364_n2688# 1.60345f
C171 source.n22 a_n2364_n2688# 0.407368f
C172 source.t5 a_n2364_n2688# 0.191541f
C173 source.t4 a_n2364_n2688# 0.191541f
C174 source.n23 a_n2364_n2688# 1.60345f
C175 source.n24 a_n2364_n2688# 0.405123f
C176 source.t11 a_n2364_n2688# 0.191541f
C177 source.t6 a_n2364_n2688# 0.191541f
C178 source.n25 a_n2364_n2688# 1.60345f
C179 source.n26 a_n2364_n2688# 0.405123f
C180 source.t27 a_n2364_n2688# 2.04249f
C181 source.n27 a_n2364_n2688# 0.627862f
C182 source.n28 a_n2364_n2688# 1.41808f
C183 plus.n0 a_n2364_n2688# 0.041967f
C184 plus.t0 a_n2364_n2688# 0.758247f
C185 plus.t8 a_n2364_n2688# 0.758247f
C186 plus.n1 a_n2364_n2688# 0.041967f
C187 plus.t2 a_n2364_n2688# 0.758247f
C188 plus.n2 a_n2364_n2688# 0.318577f
C189 plus.n3 a_n2364_n2688# 0.041967f
C190 plus.t7 a_n2364_n2688# 0.758247f
C191 plus.t1 a_n2364_n2688# 0.758247f
C192 plus.n4 a_n2364_n2688# 0.318577f
C193 plus.t3 a_n2364_n2688# 0.777738f
C194 plus.n5 a_n2364_n2688# 0.302734f
C195 plus.t9 a_n2364_n2688# 0.758247f
C196 plus.n6 a_n2364_n2688# 0.323776f
C197 plus.n7 a_n2364_n2688# 0.009523f
C198 plus.n8 a_n2364_n2688# 0.176827f
C199 plus.n9 a_n2364_n2688# 0.041967f
C200 plus.n10 a_n2364_n2688# 0.041967f
C201 plus.n11 a_n2364_n2688# 0.009523f
C202 plus.n12 a_n2364_n2688# 0.318577f
C203 plus.n13 a_n2364_n2688# 0.009523f
C204 plus.n14 a_n2364_n2688# 0.041967f
C205 plus.n15 a_n2364_n2688# 0.041967f
C206 plus.n16 a_n2364_n2688# 0.041967f
C207 plus.n17 a_n2364_n2688# 0.009523f
C208 plus.n18 a_n2364_n2688# 0.318577f
C209 plus.n19 a_n2364_n2688# 0.009523f
C210 plus.n20 a_n2364_n2688# 0.317025f
C211 plus.n21 a_n2364_n2688# 0.42746f
C212 plus.n22 a_n2364_n2688# 0.041967f
C213 plus.t13 a_n2364_n2688# 0.758247f
C214 plus.n23 a_n2364_n2688# 0.041967f
C215 plus.t12 a_n2364_n2688# 0.758247f
C216 plus.t5 a_n2364_n2688# 0.758247f
C217 plus.n24 a_n2364_n2688# 0.318577f
C218 plus.n25 a_n2364_n2688# 0.041967f
C219 plus.t4 a_n2364_n2688# 0.758247f
C220 plus.t6 a_n2364_n2688# 0.758247f
C221 plus.n26 a_n2364_n2688# 0.318577f
C222 plus.t10 a_n2364_n2688# 0.777738f
C223 plus.n27 a_n2364_n2688# 0.302734f
C224 plus.t11 a_n2364_n2688# 0.758247f
C225 plus.n28 a_n2364_n2688# 0.323776f
C226 plus.n29 a_n2364_n2688# 0.009523f
C227 plus.n30 a_n2364_n2688# 0.176827f
C228 plus.n31 a_n2364_n2688# 0.041967f
C229 plus.n32 a_n2364_n2688# 0.041967f
C230 plus.n33 a_n2364_n2688# 0.009523f
C231 plus.n34 a_n2364_n2688# 0.318577f
C232 plus.n35 a_n2364_n2688# 0.009523f
C233 plus.n36 a_n2364_n2688# 0.041967f
C234 plus.n37 a_n2364_n2688# 0.041967f
C235 plus.n38 a_n2364_n2688# 0.041967f
C236 plus.n39 a_n2364_n2688# 0.009523f
C237 plus.n40 a_n2364_n2688# 0.318577f
C238 plus.n41 a_n2364_n2688# 0.009523f
C239 plus.n42 a_n2364_n2688# 0.317025f
C240 plus.n43 a_n2364_n2688# 1.28982f
.ends

