* NGSPICE file created from diffpair336.ext - technology: sky130A

.subckt diffpair336 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t23 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 drain_right.t12 minus.t1 source.t17 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X3 drain_right.t11 minus.t2 source.t15 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 drain_right.t10 minus.t3 source.t18 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X5 source.t27 minus.t4 drain_right.t9 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X6 source.t21 minus.t5 drain_right.t8 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X7 source.t19 minus.t6 drain_right.t7 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X8 drain_left.t13 plus.t0 source.t1 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X9 source.t0 plus.t1 drain_left.t12 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X10 drain_right.t6 minus.t7 source.t24 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X11 drain_right.t5 minus.t8 source.t22 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X12 source.t20 minus.t9 drain_right.t4 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X13 source.t25 minus.t10 drain_right.t3 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X14 a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X15 source.t13 plus.t2 drain_left.t11 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X16 drain_left.t10 plus.t3 source.t3 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X17 source.t12 plus.t4 drain_left.t9 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X18 source.t4 plus.t5 drain_left.t8 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X19 a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X20 drain_right.t2 minus.t11 source.t26 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X21 drain_right.t1 minus.t12 source.t16 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X22 drain_left.t7 plus.t6 source.t7 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X23 drain_left.t6 plus.t7 source.t9 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X24 drain_left.t5 plus.t8 source.t2 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X25 drain_left.t4 plus.t9 source.t10 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X26 a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X27 drain_left.t3 plus.t10 source.t6 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X28 source.t8 plus.t11 drain_left.t2 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X29 source.t11 plus.t12 drain_left.t1 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X30 source.t14 minus.t13 drain_right.t0 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X31 drain_left.t0 plus.t13 source.t5 a_n1564_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n14 minus.t3 1290.81
R1 minus.n3 minus.t11 1290.81
R2 minus.n30 minus.t7 1290.81
R3 minus.n19 minus.t1 1290.81
R4 minus.n13 minus.t9 1241.15
R5 minus.n11 minus.t12 1241.15
R6 minus.n1 minus.t13 1241.15
R7 minus.n6 minus.t2 1241.15
R8 minus.n4 minus.t10 1241.15
R9 minus.n29 minus.t6 1241.15
R10 minus.n27 minus.t8 1241.15
R11 minus.n17 minus.t4 1241.15
R12 minus.n22 minus.t0 1241.15
R13 minus.n20 minus.t5 1241.15
R14 minus.n3 minus.n2 161.489
R15 minus.n19 minus.n18 161.489
R16 minus.n15 minus.n14 161.3
R17 minus.n12 minus.n0 161.3
R18 minus.n10 minus.n9 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n5 minus.n2 161.3
R21 minus.n31 minus.n30 161.3
R22 minus.n28 minus.n16 161.3
R23 minus.n26 minus.n25 161.3
R24 minus.n24 minus.n23 161.3
R25 minus.n21 minus.n18 161.3
R26 minus.n13 minus.n12 45.2793
R27 minus.n5 minus.n4 45.2793
R28 minus.n21 minus.n20 45.2793
R29 minus.n29 minus.n28 45.2793
R30 minus.n11 minus.n10 40.8975
R31 minus.n7 minus.n6 40.8975
R32 minus.n23 minus.n22 40.8975
R33 minus.n27 minus.n26 40.8975
R34 minus.n10 minus.n1 36.5157
R35 minus.n7 minus.n1 36.5157
R36 minus.n23 minus.n17 36.5157
R37 minus.n26 minus.n17 36.5157
R38 minus.n32 minus.n15 32.7335
R39 minus.n12 minus.n11 32.1338
R40 minus.n6 minus.n5 32.1338
R41 minus.n22 minus.n21 32.1338
R42 minus.n28 minus.n27 32.1338
R43 minus.n14 minus.n13 27.752
R44 minus.n4 minus.n3 27.752
R45 minus.n20 minus.n19 27.752
R46 minus.n30 minus.n29 27.752
R47 minus.n32 minus.n31 6.46073
R48 minus.n15 minus.n0 0.189894
R49 minus.n9 minus.n0 0.189894
R50 minus.n9 minus.n8 0.189894
R51 minus.n8 minus.n2 0.189894
R52 minus.n24 minus.n18 0.189894
R53 minus.n25 minus.n24 0.189894
R54 minus.n25 minus.n16 0.189894
R55 minus.n31 minus.n16 0.189894
R56 minus minus.n32 0.188
R57 source.n7 source.t26 51.0588
R58 source.n27 source.t24 51.0586
R59 source.n20 source.t2 51.0586
R60 source.n0 source.t1 51.0586
R61 source.n2 source.n1 48.8588
R62 source.n4 source.n3 48.8588
R63 source.n6 source.n5 48.8588
R64 source.n9 source.n8 48.8588
R65 source.n11 source.n10 48.8588
R66 source.n13 source.n12 48.8588
R67 source.n26 source.n25 48.8586
R68 source.n24 source.n23 48.8586
R69 source.n22 source.n21 48.8586
R70 source.n19 source.n18 48.8586
R71 source.n17 source.n16 48.8586
R72 source.n15 source.n14 48.8586
R73 source.n15 source.n13 19.9288
R74 source.n28 source.n0 13.9805
R75 source.n28 source.n27 5.49188
R76 source.n25 source.t22 2.2005
R77 source.n25 source.t19 2.2005
R78 source.n23 source.t23 2.2005
R79 source.n23 source.t27 2.2005
R80 source.n21 source.t17 2.2005
R81 source.n21 source.t21 2.2005
R82 source.n18 source.t10 2.2005
R83 source.n18 source.t11 2.2005
R84 source.n16 source.t9 2.2005
R85 source.n16 source.t12 2.2005
R86 source.n14 source.t7 2.2005
R87 source.n14 source.t4 2.2005
R88 source.n1 source.t6 2.2005
R89 source.n1 source.t13 2.2005
R90 source.n3 source.t5 2.2005
R91 source.n3 source.t8 2.2005
R92 source.n5 source.t3 2.2005
R93 source.n5 source.t0 2.2005
R94 source.n8 source.t15 2.2005
R95 source.n8 source.t25 2.2005
R96 source.n10 source.t16 2.2005
R97 source.n10 source.t14 2.2005
R98 source.n12 source.t18 2.2005
R99 source.n12 source.t20 2.2005
R100 source.n7 source.n6 0.698776
R101 source.n22 source.n20 0.698776
R102 source.n13 source.n11 0.457397
R103 source.n11 source.n9 0.457397
R104 source.n9 source.n7 0.457397
R105 source.n6 source.n4 0.457397
R106 source.n4 source.n2 0.457397
R107 source.n2 source.n0 0.457397
R108 source.n17 source.n15 0.457397
R109 source.n19 source.n17 0.457397
R110 source.n20 source.n19 0.457397
R111 source.n24 source.n22 0.457397
R112 source.n26 source.n24 0.457397
R113 source.n27 source.n26 0.457397
R114 source source.n28 0.188
R115 drain_right.n1 drain_right.t12 68.1942
R116 drain_right.n11 drain_right.t10 67.7376
R117 drain_right.n8 drain_right.n6 65.9943
R118 drain_right.n4 drain_right.n2 65.9942
R119 drain_right.n8 drain_right.n7 65.5376
R120 drain_right.n10 drain_right.n9 65.5376
R121 drain_right.n4 drain_right.n3 65.5373
R122 drain_right.n1 drain_right.n0 65.5373
R123 drain_right drain_right.n5 27.1683
R124 drain_right drain_right.n11 5.88166
R125 drain_right.n2 drain_right.t7 2.2005
R126 drain_right.n2 drain_right.t6 2.2005
R127 drain_right.n3 drain_right.t9 2.2005
R128 drain_right.n3 drain_right.t5 2.2005
R129 drain_right.n0 drain_right.t8 2.2005
R130 drain_right.n0 drain_right.t13 2.2005
R131 drain_right.n6 drain_right.t3 2.2005
R132 drain_right.n6 drain_right.t2 2.2005
R133 drain_right.n7 drain_right.t0 2.2005
R134 drain_right.n7 drain_right.t11 2.2005
R135 drain_right.n9 drain_right.t4 2.2005
R136 drain_right.n9 drain_right.t1 2.2005
R137 drain_right.n11 drain_right.n10 0.457397
R138 drain_right.n10 drain_right.n8 0.457397
R139 drain_right.n5 drain_right.n1 0.287826
R140 drain_right.n5 drain_right.n4 0.0593781
R141 plus.n3 plus.t3 1290.81
R142 plus.n14 plus.t0 1290.81
R143 plus.n19 plus.t8 1290.81
R144 plus.n30 plus.t6 1290.81
R145 plus.n4 plus.t1 1241.15
R146 plus.n6 plus.t13 1241.15
R147 plus.n1 plus.t11 1241.15
R148 plus.n11 plus.t10 1241.15
R149 plus.n13 plus.t2 1241.15
R150 plus.n20 plus.t12 1241.15
R151 plus.n22 plus.t9 1241.15
R152 plus.n17 plus.t4 1241.15
R153 plus.n27 plus.t7 1241.15
R154 plus.n29 plus.t5 1241.15
R155 plus.n3 plus.n2 161.489
R156 plus.n19 plus.n18 161.489
R157 plus.n5 plus.n2 161.3
R158 plus.n8 plus.n7 161.3
R159 plus.n10 plus.n9 161.3
R160 plus.n12 plus.n0 161.3
R161 plus.n15 plus.n14 161.3
R162 plus.n21 plus.n18 161.3
R163 plus.n24 plus.n23 161.3
R164 plus.n26 plus.n25 161.3
R165 plus.n28 plus.n16 161.3
R166 plus.n31 plus.n30 161.3
R167 plus.n5 plus.n4 45.2793
R168 plus.n13 plus.n12 45.2793
R169 plus.n29 plus.n28 45.2793
R170 plus.n21 plus.n20 45.2793
R171 plus.n7 plus.n6 40.8975
R172 plus.n11 plus.n10 40.8975
R173 plus.n27 plus.n26 40.8975
R174 plus.n23 plus.n22 40.8975
R175 plus.n7 plus.n1 36.5157
R176 plus.n10 plus.n1 36.5157
R177 plus.n26 plus.n17 36.5157
R178 plus.n23 plus.n17 36.5157
R179 plus.n6 plus.n5 32.1338
R180 plus.n12 plus.n11 32.1338
R181 plus.n28 plus.n27 32.1338
R182 plus.n22 plus.n21 32.1338
R183 plus.n4 plus.n3 27.752
R184 plus.n14 plus.n13 27.752
R185 plus.n30 plus.n29 27.752
R186 plus.n20 plus.n19 27.752
R187 plus plus.n31 27.7509
R188 plus plus.n15 10.9683
R189 plus.n8 plus.n2 0.189894
R190 plus.n9 plus.n8 0.189894
R191 plus.n9 plus.n0 0.189894
R192 plus.n15 plus.n0 0.189894
R193 plus.n31 plus.n16 0.189894
R194 plus.n25 plus.n16 0.189894
R195 plus.n25 plus.n24 0.189894
R196 plus.n24 plus.n18 0.189894
R197 drain_left.n7 drain_left.t10 68.1945
R198 drain_left.n1 drain_left.t7 68.1942
R199 drain_left.n4 drain_left.n2 65.9942
R200 drain_left.n9 drain_left.n8 65.5376
R201 drain_left.n7 drain_left.n6 65.5376
R202 drain_left.n11 drain_left.n10 65.5374
R203 drain_left.n4 drain_left.n3 65.5373
R204 drain_left.n1 drain_left.n0 65.5373
R205 drain_left drain_left.n5 27.7215
R206 drain_left drain_left.n11 6.11011
R207 drain_left.n2 drain_left.t1 2.2005
R208 drain_left.n2 drain_left.t5 2.2005
R209 drain_left.n3 drain_left.t9 2.2005
R210 drain_left.n3 drain_left.t4 2.2005
R211 drain_left.n0 drain_left.t8 2.2005
R212 drain_left.n0 drain_left.t6 2.2005
R213 drain_left.n10 drain_left.t11 2.2005
R214 drain_left.n10 drain_left.t13 2.2005
R215 drain_left.n8 drain_left.t2 2.2005
R216 drain_left.n8 drain_left.t3 2.2005
R217 drain_left.n6 drain_left.t12 2.2005
R218 drain_left.n6 drain_left.t0 2.2005
R219 drain_left.n9 drain_left.n7 0.457397
R220 drain_left.n11 drain_left.n9 0.457397
R221 drain_left.n5 drain_left.n1 0.287826
R222 drain_left.n5 drain_left.n4 0.0593781
C0 drain_right drain_left 0.794104f
C1 drain_right minus 3.09484f
C2 drain_left minus 0.171065f
C3 drain_right source 25.706902f
C4 drain_left source 25.7161f
C5 source minus 2.80367f
C6 drain_right plus 0.305567f
C7 drain_left plus 3.24262f
C8 plus minus 4.54945f
C9 plus source 2.81823f
C10 drain_right a_n1564_n2688# 6.55369f
C11 drain_left a_n1564_n2688# 6.8133f
C12 source a_n1564_n2688# 5.018672f
C13 minus a_n1564_n2688# 5.850102f
C14 plus a_n1564_n2688# 7.67564f
C15 drain_left.t7 a_n1564_n2688# 2.73789f
C16 drain_left.t8 a_n1564_n2688# 0.245654f
C17 drain_left.t6 a_n1564_n2688# 0.245654f
C18 drain_left.n0 a_n1564_n2688# 2.14865f
C19 drain_left.n1 a_n1564_n2688# 0.784443f
C20 drain_left.t1 a_n1564_n2688# 0.245654f
C21 drain_left.t5 a_n1564_n2688# 0.245654f
C22 drain_left.n2 a_n1564_n2688# 2.15136f
C23 drain_left.t9 a_n1564_n2688# 0.245654f
C24 drain_left.t4 a_n1564_n2688# 0.245654f
C25 drain_left.n3 a_n1564_n2688# 2.14865f
C26 drain_left.n4 a_n1564_n2688# 0.737247f
C27 drain_left.n5 a_n1564_n2688# 1.3416f
C28 drain_left.t10 a_n1564_n2688# 2.7379f
C29 drain_left.t12 a_n1564_n2688# 0.245654f
C30 drain_left.t0 a_n1564_n2688# 0.245654f
C31 drain_left.n6 a_n1564_n2688# 2.14865f
C32 drain_left.n7 a_n1564_n2688# 0.80052f
C33 drain_left.t2 a_n1564_n2688# 0.245654f
C34 drain_left.t3 a_n1564_n2688# 0.245654f
C35 drain_left.n8 a_n1564_n2688# 2.14865f
C36 drain_left.n9 a_n1564_n2688# 0.37837f
C37 drain_left.t11 a_n1564_n2688# 0.245654f
C38 drain_left.t13 a_n1564_n2688# 0.245654f
C39 drain_left.n10 a_n1564_n2688# 2.14864f
C40 drain_left.n11 a_n1564_n2688# 0.66106f
C41 plus.n0 a_n1564_n2688# 0.055414f
C42 plus.t2 a_n1564_n2688# 0.282637f
C43 plus.t10 a_n1564_n2688# 0.282637f
C44 plus.t11 a_n1564_n2688# 0.282637f
C45 plus.n1 a_n1564_n2688# 0.123718f
C46 plus.n2 a_n1564_n2688# 0.12373f
C47 plus.t13 a_n1564_n2688# 0.282637f
C48 plus.t1 a_n1564_n2688# 0.282637f
C49 plus.t3 a_n1564_n2688# 0.287449f
C50 plus.n3 a_n1564_n2688# 0.13976f
C51 plus.n4 a_n1564_n2688# 0.123718f
C52 plus.n5 a_n1564_n2688# 0.019407f
C53 plus.n6 a_n1564_n2688# 0.123718f
C54 plus.n7 a_n1564_n2688# 0.019407f
C55 plus.n8 a_n1564_n2688# 0.055414f
C56 plus.n9 a_n1564_n2688# 0.055414f
C57 plus.n10 a_n1564_n2688# 0.019407f
C58 plus.n11 a_n1564_n2688# 0.123718f
C59 plus.n12 a_n1564_n2688# 0.019407f
C60 plus.n13 a_n1564_n2688# 0.123718f
C61 plus.t0 a_n1564_n2688# 0.287449f
C62 plus.n14 a_n1564_n2688# 0.13968f
C63 plus.n15 a_n1564_n2688# 0.539042f
C64 plus.n16 a_n1564_n2688# 0.055414f
C65 plus.t6 a_n1564_n2688# 0.287449f
C66 plus.t5 a_n1564_n2688# 0.282637f
C67 plus.t7 a_n1564_n2688# 0.282637f
C68 plus.t4 a_n1564_n2688# 0.282637f
C69 plus.n17 a_n1564_n2688# 0.123718f
C70 plus.n18 a_n1564_n2688# 0.12373f
C71 plus.t9 a_n1564_n2688# 0.282637f
C72 plus.t12 a_n1564_n2688# 0.282637f
C73 plus.t8 a_n1564_n2688# 0.287449f
C74 plus.n19 a_n1564_n2688# 0.13976f
C75 plus.n20 a_n1564_n2688# 0.123718f
C76 plus.n21 a_n1564_n2688# 0.019407f
C77 plus.n22 a_n1564_n2688# 0.123718f
C78 plus.n23 a_n1564_n2688# 0.019407f
C79 plus.n24 a_n1564_n2688# 0.055414f
C80 plus.n25 a_n1564_n2688# 0.055414f
C81 plus.n26 a_n1564_n2688# 0.019407f
C82 plus.n27 a_n1564_n2688# 0.123718f
C83 plus.n28 a_n1564_n2688# 0.019407f
C84 plus.n29 a_n1564_n2688# 0.123718f
C85 plus.n30 a_n1564_n2688# 0.13968f
C86 plus.n31 a_n1564_n2688# 1.45065f
C87 drain_right.t12 a_n1564_n2688# 2.74124f
C88 drain_right.t8 a_n1564_n2688# 0.245954f
C89 drain_right.t13 a_n1564_n2688# 0.245954f
C90 drain_right.n0 a_n1564_n2688# 2.15127f
C91 drain_right.n1 a_n1564_n2688# 0.785401f
C92 drain_right.t7 a_n1564_n2688# 0.245954f
C93 drain_right.t6 a_n1564_n2688# 0.245954f
C94 drain_right.n2 a_n1564_n2688# 2.15399f
C95 drain_right.t9 a_n1564_n2688# 0.245954f
C96 drain_right.t5 a_n1564_n2688# 0.245954f
C97 drain_right.n3 a_n1564_n2688# 2.15127f
C98 drain_right.n4 a_n1564_n2688# 0.738148f
C99 drain_right.n5 a_n1564_n2688# 1.27169f
C100 drain_right.t3 a_n1564_n2688# 0.245954f
C101 drain_right.t2 a_n1564_n2688# 0.245954f
C102 drain_right.n6 a_n1564_n2688# 2.15399f
C103 drain_right.t0 a_n1564_n2688# 0.245954f
C104 drain_right.t11 a_n1564_n2688# 0.245954f
C105 drain_right.n7 a_n1564_n2688# 2.15128f
C106 drain_right.n8 a_n1564_n2688# 0.768883f
C107 drain_right.t4 a_n1564_n2688# 0.245954f
C108 drain_right.t1 a_n1564_n2688# 0.245954f
C109 drain_right.n9 a_n1564_n2688# 2.15128f
C110 drain_right.n10 a_n1564_n2688# 0.378832f
C111 drain_right.t10 a_n1564_n2688# 2.73839f
C112 drain_right.n11 a_n1564_n2688# 0.706595f
C113 source.t1 a_n1564_n2688# 2.7456f
C114 source.n0 a_n1564_n2688# 1.56195f
C115 source.t6 a_n1564_n2688# 0.257477f
C116 source.t13 a_n1564_n2688# 0.257477f
C117 source.n1 a_n1564_n2688# 2.15543f
C118 source.n2 a_n1564_n2688# 0.444014f
C119 source.t5 a_n1564_n2688# 0.257477f
C120 source.t8 a_n1564_n2688# 0.257477f
C121 source.n3 a_n1564_n2688# 2.15543f
C122 source.n4 a_n1564_n2688# 0.444014f
C123 source.t3 a_n1564_n2688# 0.257477f
C124 source.t0 a_n1564_n2688# 0.257477f
C125 source.n5 a_n1564_n2688# 2.15543f
C126 source.n6 a_n1564_n2688# 0.472172f
C127 source.t26 a_n1564_n2688# 2.74561f
C128 source.n7 a_n1564_n2688# 0.584208f
C129 source.t15 a_n1564_n2688# 0.257477f
C130 source.t25 a_n1564_n2688# 0.257477f
C131 source.n8 a_n1564_n2688# 2.15543f
C132 source.n9 a_n1564_n2688# 0.444014f
C133 source.t16 a_n1564_n2688# 0.257477f
C134 source.t14 a_n1564_n2688# 0.257477f
C135 source.n10 a_n1564_n2688# 2.15543f
C136 source.n11 a_n1564_n2688# 0.444014f
C137 source.t18 a_n1564_n2688# 0.257477f
C138 source.t20 a_n1564_n2688# 0.257477f
C139 source.n12 a_n1564_n2688# 2.15543f
C140 source.n13 a_n1564_n2688# 2.02597f
C141 source.t7 a_n1564_n2688# 0.257477f
C142 source.t4 a_n1564_n2688# 0.257477f
C143 source.n14 a_n1564_n2688# 2.15543f
C144 source.n15 a_n1564_n2688# 2.02597f
C145 source.t9 a_n1564_n2688# 0.257477f
C146 source.t12 a_n1564_n2688# 0.257477f
C147 source.n16 a_n1564_n2688# 2.15543f
C148 source.n17 a_n1564_n2688# 0.444021f
C149 source.t10 a_n1564_n2688# 0.257477f
C150 source.t11 a_n1564_n2688# 0.257477f
C151 source.n18 a_n1564_n2688# 2.15543f
C152 source.n19 a_n1564_n2688# 0.444021f
C153 source.t2 a_n1564_n2688# 2.7456f
C154 source.n20 a_n1564_n2688# 0.584215f
C155 source.t17 a_n1564_n2688# 0.257477f
C156 source.t21 a_n1564_n2688# 0.257477f
C157 source.n21 a_n1564_n2688# 2.15543f
C158 source.n22 a_n1564_n2688# 0.472179f
C159 source.t23 a_n1564_n2688# 0.257477f
C160 source.t27 a_n1564_n2688# 0.257477f
C161 source.n23 a_n1564_n2688# 2.15543f
C162 source.n24 a_n1564_n2688# 0.444021f
C163 source.t22 a_n1564_n2688# 0.257477f
C164 source.t19 a_n1564_n2688# 0.257477f
C165 source.n25 a_n1564_n2688# 2.15543f
C166 source.n26 a_n1564_n2688# 0.444021f
C167 source.t24 a_n1564_n2688# 2.7456f
C168 source.n27 a_n1564_n2688# 0.753869f
C169 source.n28 a_n1564_n2688# 1.87935f
C170 minus.n0 a_n1564_n2688# 0.054306f
C171 minus.t3 a_n1564_n2688# 0.281705f
C172 minus.t9 a_n1564_n2688# 0.276989f
C173 minus.t12 a_n1564_n2688# 0.276989f
C174 minus.t13 a_n1564_n2688# 0.276989f
C175 minus.n1 a_n1564_n2688# 0.121246f
C176 minus.n2 a_n1564_n2688# 0.121257f
C177 minus.t2 a_n1564_n2688# 0.276989f
C178 minus.t10 a_n1564_n2688# 0.276989f
C179 minus.t11 a_n1564_n2688# 0.281705f
C180 minus.n3 a_n1564_n2688# 0.136968f
C181 minus.n4 a_n1564_n2688# 0.121246f
C182 minus.n5 a_n1564_n2688# 0.01902f
C183 minus.n6 a_n1564_n2688# 0.121246f
C184 minus.n7 a_n1564_n2688# 0.01902f
C185 minus.n8 a_n1564_n2688# 0.054306f
C186 minus.n9 a_n1564_n2688# 0.054306f
C187 minus.n10 a_n1564_n2688# 0.01902f
C188 minus.n11 a_n1564_n2688# 0.121246f
C189 minus.n12 a_n1564_n2688# 0.01902f
C190 minus.n13 a_n1564_n2688# 0.121246f
C191 minus.n14 a_n1564_n2688# 0.136889f
C192 minus.n15 a_n1564_n2688# 1.63254f
C193 minus.n16 a_n1564_n2688# 0.054306f
C194 minus.t6 a_n1564_n2688# 0.276989f
C195 minus.t8 a_n1564_n2688# 0.276989f
C196 minus.t4 a_n1564_n2688# 0.276989f
C197 minus.n17 a_n1564_n2688# 0.121246f
C198 minus.n18 a_n1564_n2688# 0.121257f
C199 minus.t0 a_n1564_n2688# 0.276989f
C200 minus.t5 a_n1564_n2688# 0.276989f
C201 minus.t1 a_n1564_n2688# 0.281705f
C202 minus.n19 a_n1564_n2688# 0.136968f
C203 minus.n20 a_n1564_n2688# 0.121246f
C204 minus.n21 a_n1564_n2688# 0.01902f
C205 minus.n22 a_n1564_n2688# 0.121246f
C206 minus.n23 a_n1564_n2688# 0.01902f
C207 minus.n24 a_n1564_n2688# 0.054306f
C208 minus.n25 a_n1564_n2688# 0.054306f
C209 minus.n26 a_n1564_n2688# 0.01902f
C210 minus.n27 a_n1564_n2688# 0.121246f
C211 minus.n28 a_n1564_n2688# 0.01902f
C212 minus.n29 a_n1564_n2688# 0.121246f
C213 minus.t7 a_n1564_n2688# 0.281705f
C214 minus.n30 a_n1564_n2688# 0.136889f
C215 minus.n31 a_n1564_n2688# 0.350007f
C216 minus.n32 a_n1564_n2688# 2.00439f
.ends

