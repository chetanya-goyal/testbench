* NGSPICE file created from diffpair141.ext - technology: sky130A

.subckt diffpair141 minus drain_right drain_left source plus
X0 a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X1 a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X2 source minus drain_right a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X3 source plus drain_left a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X4 a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X5 drain_right minus source a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X6 drain_right minus source a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X7 source minus drain_right a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X8 drain_left plus source a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X9 a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X10 source plus drain_left a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X11 drain_left plus source a_n1334_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
.ends

