* NGSPICE file created from diffpair561.ext - technology: sky130A

.subckt diffpair561 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t7 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X1 drain_left.t3 plus.t0 source.t0 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X2 source.t3 plus.t1 drain_left.t2 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 drain_right.t2 minus.t1 source.t6 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X4 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X5 source.t1 plus.t2 drain_left.t1 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X6 drain_left.t0 plus.t3 source.t2 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X7 source.t5 minus.t2 drain_right.t1 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X8 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X9 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X10 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X11 source.t4 minus.t3 drain_right.t0 a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
R0 minus.n0 minus.t3 3469.67
R1 minus.n0 minus.t0 3469.67
R2 minus.n1 minus.t1 3469.67
R3 minus.n1 minus.t2 3469.67
R4 minus.n2 minus.n0 200.709
R5 minus.n2 minus.n1 167.823
R6 minus minus.n2 0.188
R7 source.n0 source.t2 44.6397
R8 source.n1 source.t3 44.6396
R9 source.n2 source.t7 44.6396
R10 source.n3 source.t4 44.6396
R11 source.n7 source.t6 44.6395
R12 source.n6 source.t5 44.6395
R13 source.n5 source.t0 44.6395
R14 source.n4 source.t1 44.6395
R15 source.n4 source.n3 27.9238
R16 source.n8 source.n0 22.3807
R17 source.n8 source.n7 5.5436
R18 source.n3 source.n2 0.560845
R19 source.n1 source.n0 0.560845
R20 source.n5 source.n4 0.560845
R21 source.n7 source.n6 0.560845
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 93.8282
R26 drain_right drain_right.n1 66.0315
R27 drain_right.n0 drain_right.t1 1.5005
R28 drain_right.n0 drain_right.t2 1.5005
R29 drain_right.n1 drain_right.t0 1.5005
R30 drain_right.n1 drain_right.t3 1.5005
R31 plus.n0 plus.t1 3469.67
R32 plus.n0 plus.t3 3469.67
R33 plus.n1 plus.t0 3469.67
R34 plus.n1 plus.t2 3469.67
R35 plus plus.n1 191.56
R36 plus plus.n0 176.498
R37 drain_left drain_left.n0 94.3814
R38 drain_left drain_left.n1 66.0315
R39 drain_left.n0 drain_left.t1 1.5005
R40 drain_left.n0 drain_left.t3 1.5005
R41 drain_left.n1 drain_left.t2 1.5005
R42 drain_left.n1 drain_left.t0 1.5005
C0 plus source 1.33235f
C1 plus minus 5.99198f
C2 drain_left drain_right 0.481587f
C3 drain_left source 15.377601f
C4 drain_left minus 0.171192f
C5 source drain_right 15.376299f
C6 minus drain_right 2.32373f
C7 source minus 1.31831f
C8 plus drain_left 2.42602f
C9 plus drain_right 0.256158f
C10 drain_right a_n1106_n4892# 8.18471f
C11 drain_left a_n1106_n4892# 8.373321f
C12 source a_n1106_n4892# 13.060591f
C13 minus a_n1106_n4892# 4.575345f
C14 plus a_n1106_n4892# 9.612821f
C15 drain_left.t1 a_n1106_n4892# 0.681453f
C16 drain_left.t3 a_n1106_n4892# 0.681453f
C17 drain_left.n0 a_n1106_n4892# 5.25779f
C18 drain_left.t2 a_n1106_n4892# 0.681453f
C19 drain_left.t0 a_n1106_n4892# 0.681453f
C20 drain_left.n1 a_n1106_n4892# 4.63089f
C21 plus.t1 a_n1106_n4892# 0.50208f
C22 plus.t3 a_n1106_n4892# 0.50208f
C23 plus.n0 a_n1106_n4892# 0.485717f
C24 plus.t2 a_n1106_n4892# 0.50208f
C25 plus.t0 a_n1106_n4892# 0.50208f
C26 plus.n1 a_n1106_n4892# 0.703693f
C27 drain_right.t1 a_n1106_n4892# 0.68189f
C28 drain_right.t2 a_n1106_n4892# 0.68189f
C29 drain_right.n0 a_n1106_n4892# 5.23244f
C30 drain_right.t0 a_n1106_n4892# 0.68189f
C31 drain_right.t3 a_n1106_n4892# 0.68189f
C32 drain_right.n1 a_n1106_n4892# 4.63385f
C33 source.t2 a_n1106_n4892# 2.96064f
C34 source.n0 a_n1106_n4892# 1.20294f
C35 source.t3 a_n1106_n4892# 2.96065f
C36 source.n1 a_n1106_n4892# 0.296852f
C37 source.t7 a_n1106_n4892# 2.96065f
C38 source.n2 a_n1106_n4892# 0.296852f
C39 source.t4 a_n1106_n4892# 2.96065f
C40 source.n3 a_n1106_n4892# 1.47275f
C41 source.t1 a_n1106_n4892# 2.96063f
C42 source.n4 a_n1106_n4892# 1.47277f
C43 source.t0 a_n1106_n4892# 2.96063f
C44 source.n5 a_n1106_n4892# 0.296868f
C45 source.t5 a_n1106_n4892# 2.96063f
C46 source.n6 a_n1106_n4892# 0.296868f
C47 source.t6 a_n1106_n4892# 2.96063f
C48 source.n7 a_n1106_n4892# 0.38336f
C49 source.n8 a_n1106_n4892# 1.37005f
C50 minus.t3 a_n1106_n4892# 0.489142f
C51 minus.t0 a_n1106_n4892# 0.489142f
C52 minus.n0 a_n1106_n4892# 0.854352f
C53 minus.t2 a_n1106_n4892# 0.489142f
C54 minus.t1 a_n1106_n4892# 0.489142f
C55 minus.n1 a_n1106_n4892# 0.4119f
C56 minus.n2 a_n1106_n4892# 5.03936f
.ends

