* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t37 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X1 a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X2 source.t16 plus.t0 drain_left.t19 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X3 a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X4 source.t24 minus.t1 drain_right.t18 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X5 source.t27 minus.t2 drain_right.t17 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X6 drain_left.t18 plus.t1 source.t15 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X7 drain_left.t17 plus.t2 source.t17 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_left.t16 plus.t3 source.t19 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X9 source.t23 minus.t3 drain_right.t16 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X10 source.t38 minus.t4 drain_right.t15 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X11 source.t25 minus.t5 drain_right.t14 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X12 source.t35 minus.t6 drain_right.t13 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X13 drain_right.t12 minus.t7 source.t26 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X14 drain_left.t15 plus.t4 source.t18 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X15 drain_left.t14 plus.t5 source.t13 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X16 drain_left.t13 plus.t6 source.t12 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X17 source.t36 minus.t8 drain_right.t11 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_right.t10 minus.t9 source.t22 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X19 drain_right.t9 minus.t10 source.t20 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X20 source.t6 plus.t7 drain_left.t12 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 source.t34 minus.t11 drain_right.t8 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 drain_left.t11 plus.t8 source.t11 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X23 source.t33 minus.t12 drain_right.t7 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X24 drain_right.t6 minus.t13 source.t29 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X25 source.t3 plus.t9 drain_left.t10 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X26 drain_right.t5 minus.t14 source.t30 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X27 source.t5 plus.t10 drain_left.t9 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X28 drain_left.t8 plus.t11 source.t8 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X29 drain_left.t7 plus.t12 source.t10 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X30 source.t31 minus.t15 drain_right.t4 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X31 drain_right.t3 minus.t16 source.t28 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X32 drain_right.t2 minus.t17 source.t21 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X33 source.t1 plus.t13 drain_left.t6 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X34 a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X35 source.t2 plus.t14 drain_left.t5 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X36 drain_left.t4 plus.t15 source.t4 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X37 drain_right.t1 minus.t18 source.t32 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X38 a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X39 drain_right.t0 minus.t19 source.t39 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X40 source.t7 plus.t16 drain_left.t3 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X41 source.t9 plus.t17 drain_left.t2 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X42 source.t14 plus.t18 drain_left.t1 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X43 source.t0 plus.t19 drain_left.t0 a_n3202_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n29 minus.n28 161.3
R1 minus.n27 minus.n0 161.3
R2 minus.n26 minus.n25 161.3
R3 minus.n24 minus.n1 161.3
R4 minus.n20 minus.n19 161.3
R5 minus.n18 minus.n3 161.3
R6 minus.n17 minus.n16 161.3
R7 minus.n15 minus.n4 161.3
R8 minus.n14 minus.n13 161.3
R9 minus.n9 minus.n6 161.3
R10 minus.n59 minus.n58 161.3
R11 minus.n57 minus.n30 161.3
R12 minus.n56 minus.n55 161.3
R13 minus.n54 minus.n31 161.3
R14 minus.n50 minus.n49 161.3
R15 minus.n48 minus.n33 161.3
R16 minus.n47 minus.n46 161.3
R17 minus.n45 minus.n34 161.3
R18 minus.n44 minus.n43 161.3
R19 minus.n39 minus.n36 161.3
R20 minus.n7 minus.t10 101.019
R21 minus.n37 minus.t6 101.019
R22 minus.n23 minus.n22 80.6037
R23 minus.n21 minus.n2 80.6037
R24 minus.n12 minus.n5 80.6037
R25 minus.n11 minus.n10 80.6037
R26 minus.n53 minus.n52 80.6037
R27 minus.n51 minus.n32 80.6037
R28 minus.n42 minus.n35 80.6037
R29 minus.n41 minus.n40 80.6037
R30 minus.n8 minus.t8 79.2293
R31 minus.n10 minus.t7 79.2293
R32 minus.n5 minus.t12 79.2293
R33 minus.n15 minus.t14 79.2293
R34 minus.n3 minus.t11 79.2293
R35 minus.n21 minus.t9 79.2293
R36 minus.n22 minus.t15 79.2293
R37 minus.n26 minus.t13 79.2293
R38 minus.n28 minus.t4 79.2293
R39 minus.n38 minus.t17 79.2293
R40 minus.n40 minus.t5 79.2293
R41 minus.n35 minus.t16 79.2293
R42 minus.n45 minus.t2 79.2293
R43 minus.n33 minus.t18 79.2293
R44 minus.n51 minus.t1 79.2293
R45 minus.n52 minus.t19 79.2293
R46 minus.n56 minus.t3 79.2293
R47 minus.n58 minus.t0 79.2293
R48 minus.n10 minus.n5 48.2005
R49 minus.n22 minus.n21 48.2005
R50 minus.n40 minus.n35 48.2005
R51 minus.n52 minus.n51 48.2005
R52 minus.n7 minus.n6 44.8565
R53 minus.n37 minus.n36 44.8565
R54 minus.n14 minus.n5 43.0884
R55 minus.n21 minus.n20 43.0884
R56 minus.n44 minus.n35 43.0884
R57 minus.n51 minus.n50 43.0884
R58 minus.n10 minus.n9 40.1672
R59 minus.n22 minus.n1 40.1672
R60 minus.n40 minus.n39 40.1672
R61 minus.n52 minus.n31 40.1672
R62 minus.n60 minus.n29 33.1217
R63 minus.n28 minus.n27 27.0217
R64 minus.n58 minus.n57 27.0217
R65 minus.n16 minus.n3 24.1005
R66 minus.n16 minus.n15 24.1005
R67 minus.n46 minus.n45 24.1005
R68 minus.n46 minus.n33 24.1005
R69 minus.n27 minus.n26 21.1793
R70 minus.n57 minus.n56 21.1793
R71 minus.n8 minus.n7 20.1275
R72 minus.n38 minus.n37 20.1275
R73 minus.n9 minus.n8 8.03383
R74 minus.n26 minus.n1 8.03383
R75 minus.n39 minus.n38 8.03383
R76 minus.n56 minus.n31 8.03383
R77 minus.n60 minus.n59 6.70505
R78 minus.n15 minus.n14 5.11262
R79 minus.n20 minus.n3 5.11262
R80 minus.n45 minus.n44 5.11262
R81 minus.n50 minus.n33 5.11262
R82 minus.n23 minus.n2 0.380177
R83 minus.n12 minus.n11 0.380177
R84 minus.n42 minus.n41 0.380177
R85 minus.n53 minus.n32 0.380177
R86 minus.n24 minus.n23 0.285035
R87 minus.n19 minus.n2 0.285035
R88 minus.n13 minus.n12 0.285035
R89 minus.n11 minus.n6 0.285035
R90 minus.n41 minus.n36 0.285035
R91 minus.n43 minus.n42 0.285035
R92 minus.n49 minus.n32 0.285035
R93 minus.n54 minus.n53 0.285035
R94 minus.n29 minus.n0 0.189894
R95 minus.n25 minus.n0 0.189894
R96 minus.n25 minus.n24 0.189894
R97 minus.n19 minus.n18 0.189894
R98 minus.n18 minus.n17 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n13 minus.n4 0.189894
R101 minus.n43 minus.n34 0.189894
R102 minus.n47 minus.n34 0.189894
R103 minus.n48 minus.n47 0.189894
R104 minus.n49 minus.n48 0.189894
R105 minus.n55 minus.n54 0.189894
R106 minus.n55 minus.n30 0.189894
R107 minus.n59 minus.n30 0.189894
R108 minus minus.n60 0.188
R109 source.n0 source.t12 243.255
R110 source.n9 source.t9 243.255
R111 source.n10 source.t20 243.255
R112 source.n19 source.t38 243.255
R113 source.n39 source.t37 243.254
R114 source.n30 source.t35 243.254
R115 source.n29 source.t18 243.254
R116 source.n20 source.t16 243.254
R117 source.n2 source.n1 223.454
R118 source.n4 source.n3 223.454
R119 source.n6 source.n5 223.454
R120 source.n8 source.n7 223.454
R121 source.n12 source.n11 223.454
R122 source.n14 source.n13 223.454
R123 source.n16 source.n15 223.454
R124 source.n18 source.n17 223.454
R125 source.n38 source.n37 223.453
R126 source.n36 source.n35 223.453
R127 source.n34 source.n33 223.453
R128 source.n32 source.n31 223.453
R129 source.n28 source.n27 223.453
R130 source.n26 source.n25 223.453
R131 source.n24 source.n23 223.453
R132 source.n22 source.n21 223.453
R133 source.n37 source.t39 19.8005
R134 source.n37 source.t23 19.8005
R135 source.n35 source.t32 19.8005
R136 source.n35 source.t24 19.8005
R137 source.n33 source.t28 19.8005
R138 source.n33 source.t27 19.8005
R139 source.n31 source.t21 19.8005
R140 source.n31 source.t25 19.8005
R141 source.n27 source.t13 19.8005
R142 source.n27 source.t7 19.8005
R143 source.n25 source.t15 19.8005
R144 source.n25 source.t14 19.8005
R145 source.n23 source.t17 19.8005
R146 source.n23 source.t0 19.8005
R147 source.n21 source.t19 19.8005
R148 source.n21 source.t3 19.8005
R149 source.n1 source.t11 19.8005
R150 source.n1 source.t6 19.8005
R151 source.n3 source.t8 19.8005
R152 source.n3 source.t5 19.8005
R153 source.n5 source.t10 19.8005
R154 source.n5 source.t2 19.8005
R155 source.n7 source.t4 19.8005
R156 source.n7 source.t1 19.8005
R157 source.n11 source.t26 19.8005
R158 source.n11 source.t36 19.8005
R159 source.n13 source.t30 19.8005
R160 source.n13 source.t33 19.8005
R161 source.n15 source.t22 19.8005
R162 source.n15 source.t34 19.8005
R163 source.n17 source.t29 19.8005
R164 source.n17 source.t31 19.8005
R165 source.n20 source.n19 13.9285
R166 source.n40 source.n0 8.17853
R167 source.n40 source.n39 5.7505
R168 source.n19 source.n18 0.974638
R169 source.n18 source.n16 0.974638
R170 source.n16 source.n14 0.974638
R171 source.n14 source.n12 0.974638
R172 source.n12 source.n10 0.974638
R173 source.n9 source.n8 0.974638
R174 source.n8 source.n6 0.974638
R175 source.n6 source.n4 0.974638
R176 source.n4 source.n2 0.974638
R177 source.n2 source.n0 0.974638
R178 source.n22 source.n20 0.974638
R179 source.n24 source.n22 0.974638
R180 source.n26 source.n24 0.974638
R181 source.n28 source.n26 0.974638
R182 source.n29 source.n28 0.974638
R183 source.n32 source.n30 0.974638
R184 source.n34 source.n32 0.974638
R185 source.n36 source.n34 0.974638
R186 source.n38 source.n36 0.974638
R187 source.n39 source.n38 0.974638
R188 source.n10 source.n9 0.470328
R189 source.n30 source.n29 0.470328
R190 source source.n40 0.188
R191 drain_right.n10 drain_right.n8 241.107
R192 drain_right.n6 drain_right.n4 241.106
R193 drain_right.n2 drain_right.n0 241.106
R194 drain_right.n10 drain_right.n9 240.132
R195 drain_right.n12 drain_right.n11 240.132
R196 drain_right.n14 drain_right.n13 240.132
R197 drain_right.n16 drain_right.n15 240.132
R198 drain_right.n7 drain_right.n3 240.131
R199 drain_right.n6 drain_right.n5 240.131
R200 drain_right.n2 drain_right.n1 240.131
R201 drain_right drain_right.n7 26.2736
R202 drain_right.n3 drain_right.t17 19.8005
R203 drain_right.n3 drain_right.t1 19.8005
R204 drain_right.n4 drain_right.t16 19.8005
R205 drain_right.n4 drain_right.t19 19.8005
R206 drain_right.n5 drain_right.t18 19.8005
R207 drain_right.n5 drain_right.t0 19.8005
R208 drain_right.n1 drain_right.t14 19.8005
R209 drain_right.n1 drain_right.t3 19.8005
R210 drain_right.n0 drain_right.t13 19.8005
R211 drain_right.n0 drain_right.t2 19.8005
R212 drain_right.n8 drain_right.t11 19.8005
R213 drain_right.n8 drain_right.t9 19.8005
R214 drain_right.n9 drain_right.t7 19.8005
R215 drain_right.n9 drain_right.t12 19.8005
R216 drain_right.n11 drain_right.t8 19.8005
R217 drain_right.n11 drain_right.t5 19.8005
R218 drain_right.n13 drain_right.t4 19.8005
R219 drain_right.n13 drain_right.t10 19.8005
R220 drain_right.n15 drain_right.t15 19.8005
R221 drain_right.n15 drain_right.t6 19.8005
R222 drain_right drain_right.n16 6.62735
R223 drain_right.n16 drain_right.n14 0.974638
R224 drain_right.n14 drain_right.n12 0.974638
R225 drain_right.n12 drain_right.n10 0.974638
R226 drain_right.n7 drain_right.n6 0.919292
R227 drain_right.n7 drain_right.n2 0.919292
R228 plus.n11 plus.n10 161.3
R229 plus.n15 plus.n14 161.3
R230 plus.n16 plus.n5 161.3
R231 plus.n18 plus.n17 161.3
R232 plus.n19 plus.n4 161.3
R233 plus.n20 plus.n3 161.3
R234 plus.n25 plus.n24 161.3
R235 plus.n26 plus.n1 161.3
R236 plus.n27 plus.n0 161.3
R237 plus.n29 plus.n28 161.3
R238 plus.n41 plus.n40 161.3
R239 plus.n45 plus.n44 161.3
R240 plus.n46 plus.n35 161.3
R241 plus.n48 plus.n47 161.3
R242 plus.n49 plus.n34 161.3
R243 plus.n50 plus.n33 161.3
R244 plus.n55 plus.n54 161.3
R245 plus.n56 plus.n31 161.3
R246 plus.n57 plus.n30 161.3
R247 plus.n59 plus.n58 161.3
R248 plus.n9 plus.t17 101.019
R249 plus.n39 plus.t4 101.019
R250 plus.n12 plus.n7 80.6037
R251 plus.n13 plus.n6 80.6037
R252 plus.n22 plus.n21 80.6037
R253 plus.n23 plus.n2 80.6037
R254 plus.n42 plus.n37 80.6037
R255 plus.n43 plus.n36 80.6037
R256 plus.n52 plus.n51 80.6037
R257 plus.n53 plus.n32 80.6037
R258 plus.n28 plus.t6 79.2293
R259 plus.n26 plus.t7 79.2293
R260 plus.n2 plus.t8 79.2293
R261 plus.n21 plus.t10 79.2293
R262 plus.n19 plus.t11 79.2293
R263 plus.n5 plus.t14 79.2293
R264 plus.n13 plus.t12 79.2293
R265 plus.n12 plus.t13 79.2293
R266 plus.n8 plus.t15 79.2293
R267 plus.n58 plus.t0 79.2293
R268 plus.n56 plus.t3 79.2293
R269 plus.n32 plus.t9 79.2293
R270 plus.n51 plus.t2 79.2293
R271 plus.n49 plus.t19 79.2293
R272 plus.n35 plus.t1 79.2293
R273 plus.n43 plus.t18 79.2293
R274 plus.n42 plus.t5 79.2293
R275 plus.n38 plus.t16 79.2293
R276 plus.n21 plus.n2 48.2005
R277 plus.n13 plus.n12 48.2005
R278 plus.n51 plus.n32 48.2005
R279 plus.n43 plus.n42 48.2005
R280 plus.n40 plus.n39 44.8565
R281 plus.n10 plus.n9 44.8565
R282 plus.n21 plus.n20 43.0884
R283 plus.n14 plus.n13 43.0884
R284 plus.n51 plus.n50 43.0884
R285 plus.n44 plus.n43 43.0884
R286 plus.n25 plus.n2 40.1672
R287 plus.n12 plus.n11 40.1672
R288 plus.n55 plus.n32 40.1672
R289 plus.n42 plus.n41 40.1672
R290 plus plus.n59 31.1695
R291 plus.n28 plus.n27 27.0217
R292 plus.n58 plus.n57 27.0217
R293 plus.n18 plus.n5 24.1005
R294 plus.n19 plus.n18 24.1005
R295 plus.n49 plus.n48 24.1005
R296 plus.n48 plus.n35 24.1005
R297 plus.n27 plus.n26 21.1793
R298 plus.n57 plus.n56 21.1793
R299 plus.n39 plus.n38 20.1275
R300 plus.n9 plus.n8 20.1275
R301 plus plus.n29 8.18232
R302 plus.n26 plus.n25 8.03383
R303 plus.n11 plus.n8 8.03383
R304 plus.n56 plus.n55 8.03383
R305 plus.n41 plus.n38 8.03383
R306 plus.n20 plus.n19 5.11262
R307 plus.n14 plus.n5 5.11262
R308 plus.n50 plus.n49 5.11262
R309 plus.n44 plus.n35 5.11262
R310 plus.n7 plus.n6 0.380177
R311 plus.n23 plus.n22 0.380177
R312 plus.n53 plus.n52 0.380177
R313 plus.n37 plus.n36 0.380177
R314 plus.n10 plus.n7 0.285035
R315 plus.n15 plus.n6 0.285035
R316 plus.n22 plus.n3 0.285035
R317 plus.n24 plus.n23 0.285035
R318 plus.n54 plus.n53 0.285035
R319 plus.n52 plus.n33 0.285035
R320 plus.n45 plus.n36 0.285035
R321 plus.n40 plus.n37 0.285035
R322 plus.n16 plus.n15 0.189894
R323 plus.n17 plus.n16 0.189894
R324 plus.n17 plus.n4 0.189894
R325 plus.n4 plus.n3 0.189894
R326 plus.n24 plus.n1 0.189894
R327 plus.n1 plus.n0 0.189894
R328 plus.n29 plus.n0 0.189894
R329 plus.n59 plus.n30 0.189894
R330 plus.n31 plus.n30 0.189894
R331 plus.n54 plus.n31 0.189894
R332 plus.n34 plus.n33 0.189894
R333 plus.n47 plus.n34 0.189894
R334 plus.n47 plus.n46 0.189894
R335 plus.n46 plus.n45 0.189894
R336 drain_left.n10 drain_left.n8 241.107
R337 drain_left.n6 drain_left.n4 241.106
R338 drain_left.n2 drain_left.n0 241.106
R339 drain_left.n16 drain_left.n15 240.132
R340 drain_left.n14 drain_left.n13 240.132
R341 drain_left.n12 drain_left.n11 240.132
R342 drain_left.n10 drain_left.n9 240.132
R343 drain_left.n7 drain_left.n3 240.131
R344 drain_left.n6 drain_left.n5 240.131
R345 drain_left.n2 drain_left.n1 240.131
R346 drain_left drain_left.n7 26.8268
R347 drain_left.n3 drain_left.t0 19.8005
R348 drain_left.n3 drain_left.t18 19.8005
R349 drain_left.n4 drain_left.t3 19.8005
R350 drain_left.n4 drain_left.t15 19.8005
R351 drain_left.n5 drain_left.t1 19.8005
R352 drain_left.n5 drain_left.t14 19.8005
R353 drain_left.n1 drain_left.t10 19.8005
R354 drain_left.n1 drain_left.t17 19.8005
R355 drain_left.n0 drain_left.t19 19.8005
R356 drain_left.n0 drain_left.t16 19.8005
R357 drain_left.n15 drain_left.t12 19.8005
R358 drain_left.n15 drain_left.t13 19.8005
R359 drain_left.n13 drain_left.t9 19.8005
R360 drain_left.n13 drain_left.t11 19.8005
R361 drain_left.n11 drain_left.t5 19.8005
R362 drain_left.n11 drain_left.t8 19.8005
R363 drain_left.n9 drain_left.t6 19.8005
R364 drain_left.n9 drain_left.t7 19.8005
R365 drain_left.n8 drain_left.t2 19.8005
R366 drain_left.n8 drain_left.t4 19.8005
R367 drain_left drain_left.n16 6.62735
R368 drain_left.n12 drain_left.n10 0.974638
R369 drain_left.n14 drain_left.n12 0.974638
R370 drain_left.n16 drain_left.n14 0.974638
R371 drain_left.n7 drain_left.n6 0.919292
R372 drain_left.n7 drain_left.n2 0.919292
C0 plus drain_left 2.10013f
C1 drain_right minus 1.78f
C2 drain_right source 5.83903f
C3 drain_right plus 0.487177f
C4 minus source 2.72566f
C5 minus plus 5.11108f
C6 plus source 2.73952f
C7 drain_right drain_left 1.72967f
C8 minus drain_left 0.181407f
C9 drain_left source 5.83616f
C10 drain_right a_n3202_n1088# 5.01557f
C11 drain_left a_n3202_n1088# 5.890191f
C12 source a_n3202_n1088# 2.982263f
C13 minus a_n3202_n1088# 11.999421f
C14 plus a_n3202_n1088# 13.38209f
C15 drain_left.t19 a_n3202_n1088# 0.021247f
C16 drain_left.t16 a_n3202_n1088# 0.021247f
C17 drain_left.n0 a_n3202_n1088# 0.084045f
C18 drain_left.t10 a_n3202_n1088# 0.021247f
C19 drain_left.t17 a_n3202_n1088# 0.021247f
C20 drain_left.n1 a_n3202_n1088# 0.08256f
C21 drain_left.n2 a_n3202_n1088# 0.718862f
C22 drain_left.t0 a_n3202_n1088# 0.021247f
C23 drain_left.t18 a_n3202_n1088# 0.021247f
C24 drain_left.n3 a_n3202_n1088# 0.08256f
C25 drain_left.t3 a_n3202_n1088# 0.021247f
C26 drain_left.t15 a_n3202_n1088# 0.021247f
C27 drain_left.n4 a_n3202_n1088# 0.084045f
C28 drain_left.t1 a_n3202_n1088# 0.021247f
C29 drain_left.t14 a_n3202_n1088# 0.021247f
C30 drain_left.n5 a_n3202_n1088# 0.08256f
C31 drain_left.n6 a_n3202_n1088# 0.718862f
C32 drain_left.n7 a_n3202_n1088# 1.38629f
C33 drain_left.t2 a_n3202_n1088# 0.021247f
C34 drain_left.t4 a_n3202_n1088# 0.021247f
C35 drain_left.n8 a_n3202_n1088# 0.084045f
C36 drain_left.t6 a_n3202_n1088# 0.021247f
C37 drain_left.t7 a_n3202_n1088# 0.021247f
C38 drain_left.n9 a_n3202_n1088# 0.08256f
C39 drain_left.n10 a_n3202_n1088# 0.722978f
C40 drain_left.t5 a_n3202_n1088# 0.021247f
C41 drain_left.t8 a_n3202_n1088# 0.021247f
C42 drain_left.n11 a_n3202_n1088# 0.08256f
C43 drain_left.n12 a_n3202_n1088# 0.356817f
C44 drain_left.t9 a_n3202_n1088# 0.021247f
C45 drain_left.t11 a_n3202_n1088# 0.021247f
C46 drain_left.n13 a_n3202_n1088# 0.08256f
C47 drain_left.n14 a_n3202_n1088# 0.356817f
C48 drain_left.t12 a_n3202_n1088# 0.021247f
C49 drain_left.t13 a_n3202_n1088# 0.021247f
C50 drain_left.n15 a_n3202_n1088# 0.08256f
C51 drain_left.n16 a_n3202_n1088# 0.597913f
C52 plus.n0 a_n3202_n1088# 0.043722f
C53 plus.t6 a_n3202_n1088# 0.11861f
C54 plus.t7 a_n3202_n1088# 0.11861f
C55 plus.n1 a_n3202_n1088# 0.043722f
C56 plus.t8 a_n3202_n1088# 0.11861f
C57 plus.n2 a_n3202_n1088# 0.125861f
C58 plus.n3 a_n3202_n1088# 0.058342f
C59 plus.t10 a_n3202_n1088# 0.11861f
C60 plus.t11 a_n3202_n1088# 0.11861f
C61 plus.n4 a_n3202_n1088# 0.043722f
C62 plus.t14 a_n3202_n1088# 0.11861f
C63 plus.n5 a_n3202_n1088# 0.113917f
C64 plus.n6 a_n3202_n1088# 0.072825f
C65 plus.t12 a_n3202_n1088# 0.11861f
C66 plus.t13 a_n3202_n1088# 0.11861f
C67 plus.n7 a_n3202_n1088# 0.072825f
C68 plus.t15 a_n3202_n1088# 0.11861f
C69 plus.n8 a_n3202_n1088# 0.117592f
C70 plus.t17 a_n3202_n1088# 0.143709f
C71 plus.n9 a_n3202_n1088# 0.095586f
C72 plus.n10 a_n3202_n1088# 0.201253f
C73 plus.n11 a_n3202_n1088# 0.009922f
C74 plus.n12 a_n3202_n1088# 0.125861f
C75 plus.n13 a_n3202_n1088# 0.1264f
C76 plus.n14 a_n3202_n1088# 0.009922f
C77 plus.n15 a_n3202_n1088# 0.058342f
C78 plus.n16 a_n3202_n1088# 0.043722f
C79 plus.n17 a_n3202_n1088# 0.043722f
C80 plus.n18 a_n3202_n1088# 0.009922f
C81 plus.n19 a_n3202_n1088# 0.113917f
C82 plus.n20 a_n3202_n1088# 0.009922f
C83 plus.n21 a_n3202_n1088# 0.1264f
C84 plus.n22 a_n3202_n1088# 0.072825f
C85 plus.n23 a_n3202_n1088# 0.072825f
C86 plus.n24 a_n3202_n1088# 0.058342f
C87 plus.n25 a_n3202_n1088# 0.009922f
C88 plus.n26 a_n3202_n1088# 0.113917f
C89 plus.n27 a_n3202_n1088# 0.009922f
C90 plus.n28 a_n3202_n1088# 0.113513f
C91 plus.n29 a_n3202_n1088# 0.321825f
C92 plus.n30 a_n3202_n1088# 0.043722f
C93 plus.t0 a_n3202_n1088# 0.11861f
C94 plus.n31 a_n3202_n1088# 0.043722f
C95 plus.t3 a_n3202_n1088# 0.11861f
C96 plus.t9 a_n3202_n1088# 0.11861f
C97 plus.n32 a_n3202_n1088# 0.125861f
C98 plus.n33 a_n3202_n1088# 0.058342f
C99 plus.t2 a_n3202_n1088# 0.11861f
C100 plus.n34 a_n3202_n1088# 0.043722f
C101 plus.t19 a_n3202_n1088# 0.11861f
C102 plus.t1 a_n3202_n1088# 0.11861f
C103 plus.n35 a_n3202_n1088# 0.113917f
C104 plus.n36 a_n3202_n1088# 0.072825f
C105 plus.t18 a_n3202_n1088# 0.11861f
C106 plus.n37 a_n3202_n1088# 0.072825f
C107 plus.t5 a_n3202_n1088# 0.11861f
C108 plus.t16 a_n3202_n1088# 0.11861f
C109 plus.n38 a_n3202_n1088# 0.117592f
C110 plus.t4 a_n3202_n1088# 0.143709f
C111 plus.n39 a_n3202_n1088# 0.095586f
C112 plus.n40 a_n3202_n1088# 0.201253f
C113 plus.n41 a_n3202_n1088# 0.009922f
C114 plus.n42 a_n3202_n1088# 0.125861f
C115 plus.n43 a_n3202_n1088# 0.1264f
C116 plus.n44 a_n3202_n1088# 0.009922f
C117 plus.n45 a_n3202_n1088# 0.058342f
C118 plus.n46 a_n3202_n1088# 0.043722f
C119 plus.n47 a_n3202_n1088# 0.043722f
C120 plus.n48 a_n3202_n1088# 0.009922f
C121 plus.n49 a_n3202_n1088# 0.113917f
C122 plus.n50 a_n3202_n1088# 0.009922f
C123 plus.n51 a_n3202_n1088# 0.1264f
C124 plus.n52 a_n3202_n1088# 0.072825f
C125 plus.n53 a_n3202_n1088# 0.072825f
C126 plus.n54 a_n3202_n1088# 0.058342f
C127 plus.n55 a_n3202_n1088# 0.009922f
C128 plus.n56 a_n3202_n1088# 0.113917f
C129 plus.n57 a_n3202_n1088# 0.009922f
C130 plus.n58 a_n3202_n1088# 0.113513f
C131 plus.n59 a_n3202_n1088# 1.29862f
C132 drain_right.t13 a_n3202_n1088# 0.01581f
C133 drain_right.t2 a_n3202_n1088# 0.01581f
C134 drain_right.n0 a_n3202_n1088# 0.062537f
C135 drain_right.t14 a_n3202_n1088# 0.01581f
C136 drain_right.t3 a_n3202_n1088# 0.01581f
C137 drain_right.n1 a_n3202_n1088# 0.061432f
C138 drain_right.n2 a_n3202_n1088# 0.534893f
C139 drain_right.t17 a_n3202_n1088# 0.01581f
C140 drain_right.t1 a_n3202_n1088# 0.01581f
C141 drain_right.n3 a_n3202_n1088# 0.061432f
C142 drain_right.t16 a_n3202_n1088# 0.01581f
C143 drain_right.t19 a_n3202_n1088# 0.01581f
C144 drain_right.n4 a_n3202_n1088# 0.062537f
C145 drain_right.t18 a_n3202_n1088# 0.01581f
C146 drain_right.t0 a_n3202_n1088# 0.01581f
C147 drain_right.n5 a_n3202_n1088# 0.061432f
C148 drain_right.n6 a_n3202_n1088# 0.534893f
C149 drain_right.n7 a_n3202_n1088# 0.993206f
C150 drain_right.t11 a_n3202_n1088# 0.01581f
C151 drain_right.t9 a_n3202_n1088# 0.01581f
C152 drain_right.n8 a_n3202_n1088# 0.062537f
C153 drain_right.t7 a_n3202_n1088# 0.01581f
C154 drain_right.t12 a_n3202_n1088# 0.01581f
C155 drain_right.n9 a_n3202_n1088# 0.061432f
C156 drain_right.n10 a_n3202_n1088# 0.537956f
C157 drain_right.t8 a_n3202_n1088# 0.01581f
C158 drain_right.t5 a_n3202_n1088# 0.01581f
C159 drain_right.n11 a_n3202_n1088# 0.061432f
C160 drain_right.n12 a_n3202_n1088# 0.265502f
C161 drain_right.t4 a_n3202_n1088# 0.01581f
C162 drain_right.t10 a_n3202_n1088# 0.01581f
C163 drain_right.n13 a_n3202_n1088# 0.061432f
C164 drain_right.n14 a_n3202_n1088# 0.265502f
C165 drain_right.t15 a_n3202_n1088# 0.01581f
C166 drain_right.t6 a_n3202_n1088# 0.01581f
C167 drain_right.n15 a_n3202_n1088# 0.061432f
C168 drain_right.n16 a_n3202_n1088# 0.444897f
C169 source.t12 a_n3202_n1088# 0.16054f
C170 source.n0 a_n3202_n1088# 0.779789f
C171 source.t11 a_n3202_n1088# 0.028844f
C172 source.t6 a_n3202_n1088# 0.028844f
C173 source.n1 a_n3202_n1088# 0.093545f
C174 source.n2 a_n3202_n1088# 0.453316f
C175 source.t8 a_n3202_n1088# 0.028844f
C176 source.t5 a_n3202_n1088# 0.028844f
C177 source.n3 a_n3202_n1088# 0.093545f
C178 source.n4 a_n3202_n1088# 0.453316f
C179 source.t10 a_n3202_n1088# 0.028844f
C180 source.t2 a_n3202_n1088# 0.028844f
C181 source.n5 a_n3202_n1088# 0.093545f
C182 source.n6 a_n3202_n1088# 0.453316f
C183 source.t4 a_n3202_n1088# 0.028844f
C184 source.t1 a_n3202_n1088# 0.028844f
C185 source.n7 a_n3202_n1088# 0.093545f
C186 source.n8 a_n3202_n1088# 0.453316f
C187 source.t9 a_n3202_n1088# 0.16054f
C188 source.n9 a_n3202_n1088# 0.405672f
C189 source.t20 a_n3202_n1088# 0.16054f
C190 source.n10 a_n3202_n1088# 0.405672f
C191 source.t26 a_n3202_n1088# 0.028844f
C192 source.t36 a_n3202_n1088# 0.028844f
C193 source.n11 a_n3202_n1088# 0.093545f
C194 source.n12 a_n3202_n1088# 0.453316f
C195 source.t30 a_n3202_n1088# 0.028844f
C196 source.t33 a_n3202_n1088# 0.028844f
C197 source.n13 a_n3202_n1088# 0.093545f
C198 source.n14 a_n3202_n1088# 0.453316f
C199 source.t22 a_n3202_n1088# 0.028844f
C200 source.t34 a_n3202_n1088# 0.028844f
C201 source.n15 a_n3202_n1088# 0.093545f
C202 source.n16 a_n3202_n1088# 0.453316f
C203 source.t29 a_n3202_n1088# 0.028844f
C204 source.t31 a_n3202_n1088# 0.028844f
C205 source.n17 a_n3202_n1088# 0.093545f
C206 source.n18 a_n3202_n1088# 0.453316f
C207 source.t38 a_n3202_n1088# 0.16054f
C208 source.n19 a_n3202_n1088# 1.0832f
C209 source.t16 a_n3202_n1088# 0.16054f
C210 source.n20 a_n3202_n1088# 1.0832f
C211 source.t19 a_n3202_n1088# 0.028844f
C212 source.t3 a_n3202_n1088# 0.028844f
C213 source.n21 a_n3202_n1088# 0.093545f
C214 source.n22 a_n3202_n1088# 0.453316f
C215 source.t17 a_n3202_n1088# 0.028844f
C216 source.t0 a_n3202_n1088# 0.028844f
C217 source.n23 a_n3202_n1088# 0.093545f
C218 source.n24 a_n3202_n1088# 0.453316f
C219 source.t15 a_n3202_n1088# 0.028844f
C220 source.t14 a_n3202_n1088# 0.028844f
C221 source.n25 a_n3202_n1088# 0.093545f
C222 source.n26 a_n3202_n1088# 0.453316f
C223 source.t13 a_n3202_n1088# 0.028844f
C224 source.t7 a_n3202_n1088# 0.028844f
C225 source.n27 a_n3202_n1088# 0.093545f
C226 source.n28 a_n3202_n1088# 0.453316f
C227 source.t18 a_n3202_n1088# 0.16054f
C228 source.n29 a_n3202_n1088# 0.405672f
C229 source.t35 a_n3202_n1088# 0.16054f
C230 source.n30 a_n3202_n1088# 0.405672f
C231 source.t21 a_n3202_n1088# 0.028844f
C232 source.t25 a_n3202_n1088# 0.028844f
C233 source.n31 a_n3202_n1088# 0.093545f
C234 source.n32 a_n3202_n1088# 0.453316f
C235 source.t28 a_n3202_n1088# 0.028844f
C236 source.t27 a_n3202_n1088# 0.028844f
C237 source.n33 a_n3202_n1088# 0.093545f
C238 source.n34 a_n3202_n1088# 0.453316f
C239 source.t32 a_n3202_n1088# 0.028844f
C240 source.t24 a_n3202_n1088# 0.028844f
C241 source.n35 a_n3202_n1088# 0.093545f
C242 source.n36 a_n3202_n1088# 0.453316f
C243 source.t39 a_n3202_n1088# 0.028844f
C244 source.t23 a_n3202_n1088# 0.028844f
C245 source.n37 a_n3202_n1088# 0.093545f
C246 source.n38 a_n3202_n1088# 0.453316f
C247 source.t37 a_n3202_n1088# 0.16054f
C248 source.n39 a_n3202_n1088# 0.651668f
C249 source.n40 a_n3202_n1088# 0.760912f
C250 minus.n0 a_n3202_n1088# 0.034143f
C251 minus.n1 a_n3202_n1088# 0.007748f
C252 minus.t13 a_n3202_n1088# 0.092623f
C253 minus.n2 a_n3202_n1088# 0.056869f
C254 minus.t11 a_n3202_n1088# 0.092623f
C255 minus.n3 a_n3202_n1088# 0.088959f
C256 minus.n4 a_n3202_n1088# 0.034143f
C257 minus.t12 a_n3202_n1088# 0.092623f
C258 minus.n5 a_n3202_n1088# 0.098706f
C259 minus.n6 a_n3202_n1088# 0.157159f
C260 minus.t10 a_n3202_n1088# 0.112223f
C261 minus.n7 a_n3202_n1088# 0.074644f
C262 minus.t8 a_n3202_n1088# 0.092623f
C263 minus.n8 a_n3202_n1088# 0.091828f
C264 minus.n9 a_n3202_n1088# 0.007748f
C265 minus.t7 a_n3202_n1088# 0.092623f
C266 minus.n10 a_n3202_n1088# 0.098285f
C267 minus.n11 a_n3202_n1088# 0.056869f
C268 minus.n12 a_n3202_n1088# 0.056869f
C269 minus.n13 a_n3202_n1088# 0.04556f
C270 minus.n14 a_n3202_n1088# 0.007748f
C271 minus.t14 a_n3202_n1088# 0.092623f
C272 minus.n15 a_n3202_n1088# 0.088959f
C273 minus.n16 a_n3202_n1088# 0.007748f
C274 minus.n17 a_n3202_n1088# 0.034143f
C275 minus.n18 a_n3202_n1088# 0.034143f
C276 minus.n19 a_n3202_n1088# 0.04556f
C277 minus.n20 a_n3202_n1088# 0.007748f
C278 minus.t9 a_n3202_n1088# 0.092623f
C279 minus.n21 a_n3202_n1088# 0.098706f
C280 minus.t15 a_n3202_n1088# 0.092623f
C281 minus.n22 a_n3202_n1088# 0.098285f
C282 minus.n23 a_n3202_n1088# 0.056869f
C283 minus.n24 a_n3202_n1088# 0.04556f
C284 minus.n25 a_n3202_n1088# 0.034143f
C285 minus.n26 a_n3202_n1088# 0.088959f
C286 minus.n27 a_n3202_n1088# 0.007748f
C287 minus.t4 a_n3202_n1088# 0.092623f
C288 minus.n28 a_n3202_n1088# 0.088643f
C289 minus.n29 a_n3202_n1088# 1.0534f
C290 minus.n30 a_n3202_n1088# 0.034143f
C291 minus.n31 a_n3202_n1088# 0.007748f
C292 minus.n32 a_n3202_n1088# 0.056869f
C293 minus.t18 a_n3202_n1088# 0.092623f
C294 minus.n33 a_n3202_n1088# 0.088959f
C295 minus.n34 a_n3202_n1088# 0.034143f
C296 minus.t16 a_n3202_n1088# 0.092623f
C297 minus.n35 a_n3202_n1088# 0.098706f
C298 minus.n36 a_n3202_n1088# 0.157159f
C299 minus.t6 a_n3202_n1088# 0.112223f
C300 minus.n37 a_n3202_n1088# 0.074644f
C301 minus.t17 a_n3202_n1088# 0.092623f
C302 minus.n38 a_n3202_n1088# 0.091828f
C303 minus.n39 a_n3202_n1088# 0.007748f
C304 minus.t5 a_n3202_n1088# 0.092623f
C305 minus.n40 a_n3202_n1088# 0.098285f
C306 minus.n41 a_n3202_n1088# 0.056869f
C307 minus.n42 a_n3202_n1088# 0.056869f
C308 minus.n43 a_n3202_n1088# 0.04556f
C309 minus.n44 a_n3202_n1088# 0.007748f
C310 minus.t2 a_n3202_n1088# 0.092623f
C311 minus.n45 a_n3202_n1088# 0.088959f
C312 minus.n46 a_n3202_n1088# 0.007748f
C313 minus.n47 a_n3202_n1088# 0.034143f
C314 minus.n48 a_n3202_n1088# 0.034143f
C315 minus.n49 a_n3202_n1088# 0.04556f
C316 minus.n50 a_n3202_n1088# 0.007748f
C317 minus.t1 a_n3202_n1088# 0.092623f
C318 minus.n51 a_n3202_n1088# 0.098706f
C319 minus.t19 a_n3202_n1088# 0.092623f
C320 minus.n52 a_n3202_n1088# 0.098285f
C321 minus.n53 a_n3202_n1088# 0.056869f
C322 minus.n54 a_n3202_n1088# 0.04556f
C323 minus.n55 a_n3202_n1088# 0.034143f
C324 minus.t3 a_n3202_n1088# 0.092623f
C325 minus.n56 a_n3202_n1088# 0.088959f
C326 minus.n57 a_n3202_n1088# 0.007748f
C327 minus.t0 a_n3202_n1088# 0.092623f
C328 minus.n58 a_n3202_n1088# 0.088643f
C329 minus.n59 a_n3202_n1088# 0.239556f
C330 minus.n60 a_n3202_n1088# 1.28399f
.ends

