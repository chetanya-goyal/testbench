* NGSPICE file created from diffpair285.ext - technology: sky130A

.subckt diffpair285 minus drain_right drain_left source plus
X0 a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X1 source.t19 plus.t0 drain_left.t0 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X2 drain_right.t11 minus.t0 source.t22 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X3 source.t3 minus.t1 drain_right.t10 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X4 source.t2 minus.t2 drain_right.t9 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X5 a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X6 source.t18 plus.t1 drain_left.t4 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X7 drain_right.t8 minus.t3 source.t6 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X8 drain_right.t7 minus.t4 source.t1 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X9 drain_right.t6 minus.t5 source.t21 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X10 drain_left.t5 plus.t2 source.t17 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X11 source.t5 minus.t6 drain_right.t5 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X12 drain_left.t1 plus.t3 source.t16 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X13 source.t15 plus.t4 drain_left.t6 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X14 a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X15 drain_right.t4 minus.t7 source.t20 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X16 source.t14 plus.t5 drain_left.t2 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X17 drain_left.t3 plus.t6 source.t13 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X18 drain_left.t7 plus.t7 source.t12 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X19 drain_right.t3 minus.t8 source.t7 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X20 source.t0 minus.t9 drain_right.t2 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X21 source.t23 minus.t10 drain_right.t1 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X22 a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X23 source.t11 plus.t8 drain_left.t8 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X24 source.t4 minus.t11 drain_right.t0 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X25 source.t10 plus.t9 drain_left.t9 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X26 drain_left.t10 plus.t10 source.t9 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X27 drain_left.t11 plus.t11 source.t8 a_n1878_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
R0 plus.n5 plus.t1 394.435
R1 plus.n19 plus.t3 394.435
R2 plus.n12 plus.t11 367.767
R3 plus.n10 plus.t8 367.767
R4 plus.n9 plus.t2 367.767
R5 plus.n3 plus.t9 367.767
R6 plus.n4 plus.t7 367.767
R7 plus.n26 plus.t0 367.767
R8 plus.n24 plus.t6 367.767
R9 plus.n23 plus.t5 367.767
R10 plus.n17 plus.t10 367.767
R11 plus.n18 plus.t4 367.767
R12 plus.n6 plus.n3 161.3
R13 plus.n8 plus.n7 161.3
R14 plus.n9 plus.n2 161.3
R15 plus.n10 plus.n1 161.3
R16 plus.n11 plus.n0 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n20 plus.n17 161.3
R19 plus.n22 plus.n21 161.3
R20 plus.n23 plus.n16 161.3
R21 plus.n24 plus.n15 161.3
R22 plus.n25 plus.n14 161.3
R23 plus.n27 plus.n26 161.3
R24 plus.n10 plus.n9 48.2005
R25 plus.n4 plus.n3 48.2005
R26 plus.n24 plus.n23 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n12 plus.n11 47.4702
R29 plus.n26 plus.n25 47.4702
R30 plus.n6 plus.n5 45.1192
R31 plus.n20 plus.n19 45.1192
R32 plus plus.n27 27.874
R33 plus.n8 plus.n3 24.1005
R34 plus.n9 plus.n8 24.1005
R35 plus.n23 plus.n22 24.1005
R36 plus.n22 plus.n17 24.1005
R37 plus.n5 plus.n4 13.6377
R38 plus.n19 plus.n18 13.6377
R39 plus plus.n13 9.90202
R40 plus.n11 plus.n10 0.730803
R41 plus.n25 plus.n24 0.730803
R42 plus.n7 plus.n6 0.189894
R43 plus.n7 plus.n2 0.189894
R44 plus.n2 plus.n1 0.189894
R45 plus.n1 plus.n0 0.189894
R46 plus.n13 plus.n0 0.189894
R47 plus.n27 plus.n14 0.189894
R48 plus.n15 plus.n14 0.189894
R49 plus.n16 plus.n15 0.189894
R50 plus.n21 plus.n16 0.189894
R51 plus.n21 plus.n20 0.189894
R52 drain_left.n6 drain_left.n4 67.9063
R53 drain_left.n3 drain_left.n2 67.8508
R54 drain_left.n3 drain_left.n0 67.8508
R55 drain_left.n6 drain_left.n5 67.1908
R56 drain_left.n8 drain_left.n7 67.1907
R57 drain_left.n3 drain_left.n1 67.1907
R58 drain_left drain_left.n3 26.3992
R59 drain_left drain_left.n8 6.36873
R60 drain_left.n1 drain_left.t2 3.3005
R61 drain_left.n1 drain_left.t10 3.3005
R62 drain_left.n2 drain_left.t6 3.3005
R63 drain_left.n2 drain_left.t1 3.3005
R64 drain_left.n0 drain_left.t0 3.3005
R65 drain_left.n0 drain_left.t3 3.3005
R66 drain_left.n7 drain_left.t8 3.3005
R67 drain_left.n7 drain_left.t11 3.3005
R68 drain_left.n5 drain_left.t9 3.3005
R69 drain_left.n5 drain_left.t5 3.3005
R70 drain_left.n4 drain_left.t4 3.3005
R71 drain_left.n4 drain_left.t7 3.3005
R72 drain_left.n8 drain_left.n6 0.716017
R73 source.n266 source.n240 289.615
R74 source.n230 source.n204 289.615
R75 source.n198 source.n172 289.615
R76 source.n162 source.n136 289.615
R77 source.n26 source.n0 289.615
R78 source.n62 source.n36 289.615
R79 source.n94 source.n68 289.615
R80 source.n130 source.n104 289.615
R81 source.n251 source.n250 185
R82 source.n248 source.n247 185
R83 source.n257 source.n256 185
R84 source.n259 source.n258 185
R85 source.n244 source.n243 185
R86 source.n265 source.n264 185
R87 source.n267 source.n266 185
R88 source.n215 source.n214 185
R89 source.n212 source.n211 185
R90 source.n221 source.n220 185
R91 source.n223 source.n222 185
R92 source.n208 source.n207 185
R93 source.n229 source.n228 185
R94 source.n231 source.n230 185
R95 source.n183 source.n182 185
R96 source.n180 source.n179 185
R97 source.n189 source.n188 185
R98 source.n191 source.n190 185
R99 source.n176 source.n175 185
R100 source.n197 source.n196 185
R101 source.n199 source.n198 185
R102 source.n147 source.n146 185
R103 source.n144 source.n143 185
R104 source.n153 source.n152 185
R105 source.n155 source.n154 185
R106 source.n140 source.n139 185
R107 source.n161 source.n160 185
R108 source.n163 source.n162 185
R109 source.n27 source.n26 185
R110 source.n25 source.n24 185
R111 source.n4 source.n3 185
R112 source.n19 source.n18 185
R113 source.n17 source.n16 185
R114 source.n8 source.n7 185
R115 source.n11 source.n10 185
R116 source.n63 source.n62 185
R117 source.n61 source.n60 185
R118 source.n40 source.n39 185
R119 source.n55 source.n54 185
R120 source.n53 source.n52 185
R121 source.n44 source.n43 185
R122 source.n47 source.n46 185
R123 source.n95 source.n94 185
R124 source.n93 source.n92 185
R125 source.n72 source.n71 185
R126 source.n87 source.n86 185
R127 source.n85 source.n84 185
R128 source.n76 source.n75 185
R129 source.n79 source.n78 185
R130 source.n131 source.n130 185
R131 source.n129 source.n128 185
R132 source.n108 source.n107 185
R133 source.n123 source.n122 185
R134 source.n121 source.n120 185
R135 source.n112 source.n111 185
R136 source.n115 source.n114 185
R137 source.t6 source.n249 147.661
R138 source.t0 source.n213 147.661
R139 source.t16 source.n181 147.661
R140 source.t19 source.n145 147.661
R141 source.t8 source.n9 147.661
R142 source.t18 source.n45 147.661
R143 source.t20 source.n77 147.661
R144 source.t5 source.n113 147.661
R145 source.n250 source.n247 104.615
R146 source.n257 source.n247 104.615
R147 source.n258 source.n257 104.615
R148 source.n258 source.n243 104.615
R149 source.n265 source.n243 104.615
R150 source.n266 source.n265 104.615
R151 source.n214 source.n211 104.615
R152 source.n221 source.n211 104.615
R153 source.n222 source.n221 104.615
R154 source.n222 source.n207 104.615
R155 source.n229 source.n207 104.615
R156 source.n230 source.n229 104.615
R157 source.n182 source.n179 104.615
R158 source.n189 source.n179 104.615
R159 source.n190 source.n189 104.615
R160 source.n190 source.n175 104.615
R161 source.n197 source.n175 104.615
R162 source.n198 source.n197 104.615
R163 source.n146 source.n143 104.615
R164 source.n153 source.n143 104.615
R165 source.n154 source.n153 104.615
R166 source.n154 source.n139 104.615
R167 source.n161 source.n139 104.615
R168 source.n162 source.n161 104.615
R169 source.n26 source.n25 104.615
R170 source.n25 source.n3 104.615
R171 source.n18 source.n3 104.615
R172 source.n18 source.n17 104.615
R173 source.n17 source.n7 104.615
R174 source.n10 source.n7 104.615
R175 source.n62 source.n61 104.615
R176 source.n61 source.n39 104.615
R177 source.n54 source.n39 104.615
R178 source.n54 source.n53 104.615
R179 source.n53 source.n43 104.615
R180 source.n46 source.n43 104.615
R181 source.n94 source.n93 104.615
R182 source.n93 source.n71 104.615
R183 source.n86 source.n71 104.615
R184 source.n86 source.n85 104.615
R185 source.n85 source.n75 104.615
R186 source.n78 source.n75 104.615
R187 source.n130 source.n129 104.615
R188 source.n129 source.n107 104.615
R189 source.n122 source.n107 104.615
R190 source.n122 source.n121 104.615
R191 source.n121 source.n111 104.615
R192 source.n114 source.n111 104.615
R193 source.n250 source.t6 52.3082
R194 source.n214 source.t0 52.3082
R195 source.n182 source.t16 52.3082
R196 source.n146 source.t19 52.3082
R197 source.n10 source.t8 52.3082
R198 source.n46 source.t18 52.3082
R199 source.n78 source.t20 52.3082
R200 source.n114 source.t5 52.3082
R201 source.n33 source.n32 50.512
R202 source.n35 source.n34 50.512
R203 source.n101 source.n100 50.512
R204 source.n103 source.n102 50.512
R205 source.n239 source.n238 50.5119
R206 source.n237 source.n236 50.5119
R207 source.n171 source.n170 50.5119
R208 source.n169 source.n168 50.5119
R209 source.n271 source.n270 32.1853
R210 source.n235 source.n234 32.1853
R211 source.n203 source.n202 32.1853
R212 source.n167 source.n166 32.1853
R213 source.n31 source.n30 32.1853
R214 source.n67 source.n66 32.1853
R215 source.n99 source.n98 32.1853
R216 source.n135 source.n134 32.1853
R217 source.n167 source.n135 17.4578
R218 source.n251 source.n249 15.6674
R219 source.n215 source.n213 15.6674
R220 source.n183 source.n181 15.6674
R221 source.n147 source.n145 15.6674
R222 source.n11 source.n9 15.6674
R223 source.n47 source.n45 15.6674
R224 source.n79 source.n77 15.6674
R225 source.n115 source.n113 15.6674
R226 source.n252 source.n248 12.8005
R227 source.n216 source.n212 12.8005
R228 source.n184 source.n180 12.8005
R229 source.n148 source.n144 12.8005
R230 source.n12 source.n8 12.8005
R231 source.n48 source.n44 12.8005
R232 source.n80 source.n76 12.8005
R233 source.n116 source.n112 12.8005
R234 source.n256 source.n255 12.0247
R235 source.n220 source.n219 12.0247
R236 source.n188 source.n187 12.0247
R237 source.n152 source.n151 12.0247
R238 source.n16 source.n15 12.0247
R239 source.n52 source.n51 12.0247
R240 source.n84 source.n83 12.0247
R241 source.n120 source.n119 12.0247
R242 source.n272 source.n31 11.8371
R243 source.n259 source.n246 11.249
R244 source.n223 source.n210 11.249
R245 source.n191 source.n178 11.249
R246 source.n155 source.n142 11.249
R247 source.n19 source.n6 11.249
R248 source.n55 source.n42 11.249
R249 source.n87 source.n74 11.249
R250 source.n123 source.n110 11.249
R251 source.n260 source.n244 10.4732
R252 source.n224 source.n208 10.4732
R253 source.n192 source.n176 10.4732
R254 source.n156 source.n140 10.4732
R255 source.n20 source.n4 10.4732
R256 source.n56 source.n40 10.4732
R257 source.n88 source.n72 10.4732
R258 source.n124 source.n108 10.4732
R259 source.n264 source.n263 9.69747
R260 source.n228 source.n227 9.69747
R261 source.n196 source.n195 9.69747
R262 source.n160 source.n159 9.69747
R263 source.n24 source.n23 9.69747
R264 source.n60 source.n59 9.69747
R265 source.n92 source.n91 9.69747
R266 source.n128 source.n127 9.69747
R267 source.n270 source.n269 9.45567
R268 source.n234 source.n233 9.45567
R269 source.n202 source.n201 9.45567
R270 source.n166 source.n165 9.45567
R271 source.n30 source.n29 9.45567
R272 source.n66 source.n65 9.45567
R273 source.n98 source.n97 9.45567
R274 source.n134 source.n133 9.45567
R275 source.n269 source.n268 9.3005
R276 source.n242 source.n241 9.3005
R277 source.n263 source.n262 9.3005
R278 source.n261 source.n260 9.3005
R279 source.n246 source.n245 9.3005
R280 source.n255 source.n254 9.3005
R281 source.n253 source.n252 9.3005
R282 source.n233 source.n232 9.3005
R283 source.n206 source.n205 9.3005
R284 source.n227 source.n226 9.3005
R285 source.n225 source.n224 9.3005
R286 source.n210 source.n209 9.3005
R287 source.n219 source.n218 9.3005
R288 source.n217 source.n216 9.3005
R289 source.n201 source.n200 9.3005
R290 source.n174 source.n173 9.3005
R291 source.n195 source.n194 9.3005
R292 source.n193 source.n192 9.3005
R293 source.n178 source.n177 9.3005
R294 source.n187 source.n186 9.3005
R295 source.n185 source.n184 9.3005
R296 source.n165 source.n164 9.3005
R297 source.n138 source.n137 9.3005
R298 source.n159 source.n158 9.3005
R299 source.n157 source.n156 9.3005
R300 source.n142 source.n141 9.3005
R301 source.n151 source.n150 9.3005
R302 source.n149 source.n148 9.3005
R303 source.n29 source.n28 9.3005
R304 source.n2 source.n1 9.3005
R305 source.n23 source.n22 9.3005
R306 source.n21 source.n20 9.3005
R307 source.n6 source.n5 9.3005
R308 source.n15 source.n14 9.3005
R309 source.n13 source.n12 9.3005
R310 source.n65 source.n64 9.3005
R311 source.n38 source.n37 9.3005
R312 source.n59 source.n58 9.3005
R313 source.n57 source.n56 9.3005
R314 source.n42 source.n41 9.3005
R315 source.n51 source.n50 9.3005
R316 source.n49 source.n48 9.3005
R317 source.n97 source.n96 9.3005
R318 source.n70 source.n69 9.3005
R319 source.n91 source.n90 9.3005
R320 source.n89 source.n88 9.3005
R321 source.n74 source.n73 9.3005
R322 source.n83 source.n82 9.3005
R323 source.n81 source.n80 9.3005
R324 source.n133 source.n132 9.3005
R325 source.n106 source.n105 9.3005
R326 source.n127 source.n126 9.3005
R327 source.n125 source.n124 9.3005
R328 source.n110 source.n109 9.3005
R329 source.n119 source.n118 9.3005
R330 source.n117 source.n116 9.3005
R331 source.n267 source.n242 8.92171
R332 source.n231 source.n206 8.92171
R333 source.n199 source.n174 8.92171
R334 source.n163 source.n138 8.92171
R335 source.n27 source.n2 8.92171
R336 source.n63 source.n38 8.92171
R337 source.n95 source.n70 8.92171
R338 source.n131 source.n106 8.92171
R339 source.n268 source.n240 8.14595
R340 source.n232 source.n204 8.14595
R341 source.n200 source.n172 8.14595
R342 source.n164 source.n136 8.14595
R343 source.n28 source.n0 8.14595
R344 source.n64 source.n36 8.14595
R345 source.n96 source.n68 8.14595
R346 source.n132 source.n104 8.14595
R347 source.n270 source.n240 5.81868
R348 source.n234 source.n204 5.81868
R349 source.n202 source.n172 5.81868
R350 source.n166 source.n136 5.81868
R351 source.n30 source.n0 5.81868
R352 source.n66 source.n36 5.81868
R353 source.n98 source.n68 5.81868
R354 source.n134 source.n104 5.81868
R355 source.n272 source.n271 5.62119
R356 source.n268 source.n267 5.04292
R357 source.n232 source.n231 5.04292
R358 source.n200 source.n199 5.04292
R359 source.n164 source.n163 5.04292
R360 source.n28 source.n27 5.04292
R361 source.n64 source.n63 5.04292
R362 source.n96 source.n95 5.04292
R363 source.n132 source.n131 5.04292
R364 source.n253 source.n249 4.38594
R365 source.n217 source.n213 4.38594
R366 source.n185 source.n181 4.38594
R367 source.n149 source.n145 4.38594
R368 source.n13 source.n9 4.38594
R369 source.n49 source.n45 4.38594
R370 source.n81 source.n77 4.38594
R371 source.n117 source.n113 4.38594
R372 source.n264 source.n242 4.26717
R373 source.n228 source.n206 4.26717
R374 source.n196 source.n174 4.26717
R375 source.n160 source.n138 4.26717
R376 source.n24 source.n2 4.26717
R377 source.n60 source.n38 4.26717
R378 source.n92 source.n70 4.26717
R379 source.n128 source.n106 4.26717
R380 source.n263 source.n244 3.49141
R381 source.n227 source.n208 3.49141
R382 source.n195 source.n176 3.49141
R383 source.n159 source.n140 3.49141
R384 source.n23 source.n4 3.49141
R385 source.n59 source.n40 3.49141
R386 source.n91 source.n72 3.49141
R387 source.n127 source.n108 3.49141
R388 source.n238 source.t22 3.3005
R389 source.n238 source.t4 3.3005
R390 source.n236 source.t7 3.3005
R391 source.n236 source.t3 3.3005
R392 source.n170 source.t9 3.3005
R393 source.n170 source.t15 3.3005
R394 source.n168 source.t13 3.3005
R395 source.n168 source.t14 3.3005
R396 source.n32 source.t17 3.3005
R397 source.n32 source.t11 3.3005
R398 source.n34 source.t12 3.3005
R399 source.n34 source.t10 3.3005
R400 source.n100 source.t21 3.3005
R401 source.n100 source.t2 3.3005
R402 source.n102 source.t1 3.3005
R403 source.n102 source.t23 3.3005
R404 source.n260 source.n259 2.71565
R405 source.n224 source.n223 2.71565
R406 source.n192 source.n191 2.71565
R407 source.n156 source.n155 2.71565
R408 source.n20 source.n19 2.71565
R409 source.n56 source.n55 2.71565
R410 source.n88 source.n87 2.71565
R411 source.n124 source.n123 2.71565
R412 source.n256 source.n246 1.93989
R413 source.n220 source.n210 1.93989
R414 source.n188 source.n178 1.93989
R415 source.n152 source.n142 1.93989
R416 source.n16 source.n6 1.93989
R417 source.n52 source.n42 1.93989
R418 source.n84 source.n74 1.93989
R419 source.n120 source.n110 1.93989
R420 source.n255 source.n248 1.16414
R421 source.n219 source.n212 1.16414
R422 source.n187 source.n180 1.16414
R423 source.n151 source.n144 1.16414
R424 source.n15 source.n8 1.16414
R425 source.n51 source.n44 1.16414
R426 source.n83 source.n76 1.16414
R427 source.n119 source.n112 1.16414
R428 source.n135 source.n103 0.716017
R429 source.n103 source.n101 0.716017
R430 source.n101 source.n99 0.716017
R431 source.n67 source.n35 0.716017
R432 source.n35 source.n33 0.716017
R433 source.n33 source.n31 0.716017
R434 source.n169 source.n167 0.716017
R435 source.n171 source.n169 0.716017
R436 source.n203 source.n171 0.716017
R437 source.n237 source.n235 0.716017
R438 source.n239 source.n237 0.716017
R439 source.n271 source.n239 0.716017
R440 source.n99 source.n67 0.470328
R441 source.n235 source.n203 0.470328
R442 source.n252 source.n251 0.388379
R443 source.n216 source.n215 0.388379
R444 source.n184 source.n183 0.388379
R445 source.n148 source.n147 0.388379
R446 source.n12 source.n11 0.388379
R447 source.n48 source.n47 0.388379
R448 source.n80 source.n79 0.388379
R449 source.n116 source.n115 0.388379
R450 source source.n272 0.188
R451 source.n254 source.n253 0.155672
R452 source.n254 source.n245 0.155672
R453 source.n261 source.n245 0.155672
R454 source.n262 source.n261 0.155672
R455 source.n262 source.n241 0.155672
R456 source.n269 source.n241 0.155672
R457 source.n218 source.n217 0.155672
R458 source.n218 source.n209 0.155672
R459 source.n225 source.n209 0.155672
R460 source.n226 source.n225 0.155672
R461 source.n226 source.n205 0.155672
R462 source.n233 source.n205 0.155672
R463 source.n186 source.n185 0.155672
R464 source.n186 source.n177 0.155672
R465 source.n193 source.n177 0.155672
R466 source.n194 source.n193 0.155672
R467 source.n194 source.n173 0.155672
R468 source.n201 source.n173 0.155672
R469 source.n150 source.n149 0.155672
R470 source.n150 source.n141 0.155672
R471 source.n157 source.n141 0.155672
R472 source.n158 source.n157 0.155672
R473 source.n158 source.n137 0.155672
R474 source.n165 source.n137 0.155672
R475 source.n29 source.n1 0.155672
R476 source.n22 source.n1 0.155672
R477 source.n22 source.n21 0.155672
R478 source.n21 source.n5 0.155672
R479 source.n14 source.n5 0.155672
R480 source.n14 source.n13 0.155672
R481 source.n65 source.n37 0.155672
R482 source.n58 source.n37 0.155672
R483 source.n58 source.n57 0.155672
R484 source.n57 source.n41 0.155672
R485 source.n50 source.n41 0.155672
R486 source.n50 source.n49 0.155672
R487 source.n97 source.n69 0.155672
R488 source.n90 source.n69 0.155672
R489 source.n90 source.n89 0.155672
R490 source.n89 source.n73 0.155672
R491 source.n82 source.n73 0.155672
R492 source.n82 source.n81 0.155672
R493 source.n133 source.n105 0.155672
R494 source.n126 source.n105 0.155672
R495 source.n126 source.n125 0.155672
R496 source.n125 source.n109 0.155672
R497 source.n118 source.n109 0.155672
R498 source.n118 source.n117 0.155672
R499 minus.n3 minus.t7 394.435
R500 minus.n17 minus.t9 394.435
R501 minus.n4 minus.t2 367.767
R502 minus.n5 minus.t5 367.767
R503 minus.n1 minus.t10 367.767
R504 minus.n10 minus.t4 367.767
R505 minus.n12 minus.t6 367.767
R506 minus.n18 minus.t8 367.767
R507 minus.n19 minus.t1 367.767
R508 minus.n15 minus.t0 367.767
R509 minus.n24 minus.t11 367.767
R510 minus.n26 minus.t3 367.767
R511 minus.n13 minus.n12 161.3
R512 minus.n11 minus.n0 161.3
R513 minus.n10 minus.n9 161.3
R514 minus.n8 minus.n1 161.3
R515 minus.n7 minus.n6 161.3
R516 minus.n5 minus.n2 161.3
R517 minus.n27 minus.n26 161.3
R518 minus.n25 minus.n14 161.3
R519 minus.n24 minus.n23 161.3
R520 minus.n22 minus.n15 161.3
R521 minus.n21 minus.n20 161.3
R522 minus.n19 minus.n16 161.3
R523 minus.n5 minus.n4 48.2005
R524 minus.n10 minus.n1 48.2005
R525 minus.n19 minus.n18 48.2005
R526 minus.n24 minus.n15 48.2005
R527 minus.n12 minus.n11 47.4702
R528 minus.n26 minus.n25 47.4702
R529 minus.n3 minus.n2 45.1192
R530 minus.n17 minus.n16 45.1192
R531 minus.n28 minus.n13 31.7202
R532 minus.n6 minus.n1 24.1005
R533 minus.n6 minus.n5 24.1005
R534 minus.n20 minus.n19 24.1005
R535 minus.n20 minus.n15 24.1005
R536 minus.n4 minus.n3 13.6377
R537 minus.n18 minus.n17 13.6377
R538 minus.n28 minus.n27 6.5308
R539 minus.n11 minus.n10 0.730803
R540 minus.n25 minus.n24 0.730803
R541 minus.n13 minus.n0 0.189894
R542 minus.n9 minus.n0 0.189894
R543 minus.n9 minus.n8 0.189894
R544 minus.n8 minus.n7 0.189894
R545 minus.n7 minus.n2 0.189894
R546 minus.n21 minus.n16 0.189894
R547 minus.n22 minus.n21 0.189894
R548 minus.n23 minus.n22 0.189894
R549 minus.n23 minus.n14 0.189894
R550 minus.n27 minus.n14 0.189894
R551 minus minus.n28 0.188
R552 drain_right.n6 drain_right.n4 67.9062
R553 drain_right.n3 drain_right.n2 67.8508
R554 drain_right.n3 drain_right.n0 67.8508
R555 drain_right.n6 drain_right.n5 67.1908
R556 drain_right.n8 drain_right.n7 67.1908
R557 drain_right.n3 drain_right.n1 67.1907
R558 drain_right drain_right.n3 25.846
R559 drain_right drain_right.n8 6.36873
R560 drain_right.n1 drain_right.t10 3.3005
R561 drain_right.n1 drain_right.t11 3.3005
R562 drain_right.n2 drain_right.t0 3.3005
R563 drain_right.n2 drain_right.t8 3.3005
R564 drain_right.n0 drain_right.t2 3.3005
R565 drain_right.n0 drain_right.t3 3.3005
R566 drain_right.n4 drain_right.t9 3.3005
R567 drain_right.n4 drain_right.t4 3.3005
R568 drain_right.n5 drain_right.t1 3.3005
R569 drain_right.n5 drain_right.t6 3.3005
R570 drain_right.n7 drain_right.t5 3.3005
R571 drain_right.n7 drain_right.t7 3.3005
R572 drain_right.n8 drain_right.n6 0.716017
C0 source drain_left 10.4252f
C1 minus source 3.54459f
C2 source drain_right 10.426201f
C3 minus drain_left 0.171641f
C4 drain_left drain_right 0.936346f
C5 minus drain_right 3.47246f
C6 plus source 3.55861f
C7 plus drain_left 3.65505f
C8 plus minus 4.38212f
C9 plus drain_right 0.337327f
C10 drain_right a_n1878_n2088# 4.85409f
C11 drain_left a_n1878_n2088# 5.14037f
C12 source a_n1878_n2088# 5.403161f
C13 minus a_n1878_n2088# 6.877763f
C14 plus a_n1878_n2088# 8.373f
C15 drain_right.t2 a_n1878_n2088# 0.135938f
C16 drain_right.t3 a_n1878_n2088# 0.135938f
C17 drain_right.n0 a_n1878_n2088# 1.13735f
C18 drain_right.t10 a_n1878_n2088# 0.135938f
C19 drain_right.t11 a_n1878_n2088# 0.135938f
C20 drain_right.n1 a_n1878_n2088# 1.13372f
C21 drain_right.t0 a_n1878_n2088# 0.135938f
C22 drain_right.t8 a_n1878_n2088# 0.135938f
C23 drain_right.n2 a_n1878_n2088# 1.13735f
C24 drain_right.n3 a_n1878_n2088# 2.03395f
C25 drain_right.t9 a_n1878_n2088# 0.135938f
C26 drain_right.t4 a_n1878_n2088# 0.135938f
C27 drain_right.n4 a_n1878_n2088# 1.13769f
C28 drain_right.t1 a_n1878_n2088# 0.135938f
C29 drain_right.t6 a_n1878_n2088# 0.135938f
C30 drain_right.n5 a_n1878_n2088# 1.13373f
C31 drain_right.n6 a_n1878_n2088# 0.737382f
C32 drain_right.t5 a_n1878_n2088# 0.135938f
C33 drain_right.t7 a_n1878_n2088# 0.135938f
C34 drain_right.n7 a_n1878_n2088# 1.13373f
C35 drain_right.n8 a_n1878_n2088# 0.611218f
C36 minus.n0 a_n1878_n2088# 0.046998f
C37 minus.t10 a_n1878_n2088# 0.408961f
C38 minus.n1 a_n1878_n2088# 0.197426f
C39 minus.t4 a_n1878_n2088# 0.408961f
C40 minus.n2 a_n1878_n2088# 0.191406f
C41 minus.t7 a_n1878_n2088# 0.42199f
C42 minus.n3 a_n1878_n2088# 0.180768f
C43 minus.t2 a_n1878_n2088# 0.408961f
C44 minus.n4 a_n1878_n2088# 0.203091f
C45 minus.t5 a_n1878_n2088# 0.408961f
C46 minus.n5 a_n1878_n2088# 0.197426f
C47 minus.n6 a_n1878_n2088# 0.010665f
C48 minus.n7 a_n1878_n2088# 0.046998f
C49 minus.n8 a_n1878_n2088# 0.046998f
C50 minus.n9 a_n1878_n2088# 0.046998f
C51 minus.n10 a_n1878_n2088# 0.19279f
C52 minus.n11 a_n1878_n2088# 0.010665f
C53 minus.t6 a_n1878_n2088# 0.408961f
C54 minus.n12 a_n1878_n2088# 0.1925f
C55 minus.n13 a_n1878_n2088# 1.34424f
C56 minus.n14 a_n1878_n2088# 0.046998f
C57 minus.t0 a_n1878_n2088# 0.408961f
C58 minus.n15 a_n1878_n2088# 0.197426f
C59 minus.n16 a_n1878_n2088# 0.191406f
C60 minus.t9 a_n1878_n2088# 0.42199f
C61 minus.n17 a_n1878_n2088# 0.180768f
C62 minus.t8 a_n1878_n2088# 0.408961f
C63 minus.n18 a_n1878_n2088# 0.203091f
C64 minus.t1 a_n1878_n2088# 0.408961f
C65 minus.n19 a_n1878_n2088# 0.197426f
C66 minus.n20 a_n1878_n2088# 0.010665f
C67 minus.n21 a_n1878_n2088# 0.046998f
C68 minus.n22 a_n1878_n2088# 0.046998f
C69 minus.n23 a_n1878_n2088# 0.046998f
C70 minus.t11 a_n1878_n2088# 0.408961f
C71 minus.n24 a_n1878_n2088# 0.19279f
C72 minus.n25 a_n1878_n2088# 0.010665f
C73 minus.t3 a_n1878_n2088# 0.408961f
C74 minus.n26 a_n1878_n2088# 0.1925f
C75 minus.n27 a_n1878_n2088# 0.310667f
C76 minus.n28 a_n1878_n2088# 1.65118f
C77 source.n0 a_n1878_n2088# 0.034887f
C78 source.n1 a_n1878_n2088# 0.02482f
C79 source.n2 a_n1878_n2088# 0.013337f
C80 source.n3 a_n1878_n2088# 0.031524f
C81 source.n4 a_n1878_n2088# 0.014122f
C82 source.n5 a_n1878_n2088# 0.02482f
C83 source.n6 a_n1878_n2088# 0.013337f
C84 source.n7 a_n1878_n2088# 0.031524f
C85 source.n8 a_n1878_n2088# 0.014122f
C86 source.n9 a_n1878_n2088# 0.106213f
C87 source.t8 a_n1878_n2088# 0.051381f
C88 source.n10 a_n1878_n2088# 0.023643f
C89 source.n11 a_n1878_n2088# 0.018621f
C90 source.n12 a_n1878_n2088# 0.013337f
C91 source.n13 a_n1878_n2088# 0.590571f
C92 source.n14 a_n1878_n2088# 0.02482f
C93 source.n15 a_n1878_n2088# 0.013337f
C94 source.n16 a_n1878_n2088# 0.014122f
C95 source.n17 a_n1878_n2088# 0.031524f
C96 source.n18 a_n1878_n2088# 0.031524f
C97 source.n19 a_n1878_n2088# 0.014122f
C98 source.n20 a_n1878_n2088# 0.013337f
C99 source.n21 a_n1878_n2088# 0.02482f
C100 source.n22 a_n1878_n2088# 0.02482f
C101 source.n23 a_n1878_n2088# 0.013337f
C102 source.n24 a_n1878_n2088# 0.014122f
C103 source.n25 a_n1878_n2088# 0.031524f
C104 source.n26 a_n1878_n2088# 0.068245f
C105 source.n27 a_n1878_n2088# 0.014122f
C106 source.n28 a_n1878_n2088# 0.013337f
C107 source.n29 a_n1878_n2088# 0.057371f
C108 source.n30 a_n1878_n2088# 0.038186f
C109 source.n31 a_n1878_n2088# 0.624813f
C110 source.t17 a_n1878_n2088# 0.117682f
C111 source.t11 a_n1878_n2088# 0.117682f
C112 source.n32 a_n1878_n2088# 0.916514f
C113 source.n33 a_n1878_n2088# 0.347113f
C114 source.t12 a_n1878_n2088# 0.117682f
C115 source.t10 a_n1878_n2088# 0.117682f
C116 source.n34 a_n1878_n2088# 0.916514f
C117 source.n35 a_n1878_n2088# 0.347113f
C118 source.n36 a_n1878_n2088# 0.034887f
C119 source.n37 a_n1878_n2088# 0.02482f
C120 source.n38 a_n1878_n2088# 0.013337f
C121 source.n39 a_n1878_n2088# 0.031524f
C122 source.n40 a_n1878_n2088# 0.014122f
C123 source.n41 a_n1878_n2088# 0.02482f
C124 source.n42 a_n1878_n2088# 0.013337f
C125 source.n43 a_n1878_n2088# 0.031524f
C126 source.n44 a_n1878_n2088# 0.014122f
C127 source.n45 a_n1878_n2088# 0.106213f
C128 source.t18 a_n1878_n2088# 0.051381f
C129 source.n46 a_n1878_n2088# 0.023643f
C130 source.n47 a_n1878_n2088# 0.018621f
C131 source.n48 a_n1878_n2088# 0.013337f
C132 source.n49 a_n1878_n2088# 0.590571f
C133 source.n50 a_n1878_n2088# 0.02482f
C134 source.n51 a_n1878_n2088# 0.013337f
C135 source.n52 a_n1878_n2088# 0.014122f
C136 source.n53 a_n1878_n2088# 0.031524f
C137 source.n54 a_n1878_n2088# 0.031524f
C138 source.n55 a_n1878_n2088# 0.014122f
C139 source.n56 a_n1878_n2088# 0.013337f
C140 source.n57 a_n1878_n2088# 0.02482f
C141 source.n58 a_n1878_n2088# 0.02482f
C142 source.n59 a_n1878_n2088# 0.013337f
C143 source.n60 a_n1878_n2088# 0.014122f
C144 source.n61 a_n1878_n2088# 0.031524f
C145 source.n62 a_n1878_n2088# 0.068245f
C146 source.n63 a_n1878_n2088# 0.014122f
C147 source.n64 a_n1878_n2088# 0.013337f
C148 source.n65 a_n1878_n2088# 0.057371f
C149 source.n66 a_n1878_n2088# 0.038186f
C150 source.n67 a_n1878_n2088# 0.115997f
C151 source.n68 a_n1878_n2088# 0.034887f
C152 source.n69 a_n1878_n2088# 0.02482f
C153 source.n70 a_n1878_n2088# 0.013337f
C154 source.n71 a_n1878_n2088# 0.031524f
C155 source.n72 a_n1878_n2088# 0.014122f
C156 source.n73 a_n1878_n2088# 0.02482f
C157 source.n74 a_n1878_n2088# 0.013337f
C158 source.n75 a_n1878_n2088# 0.031524f
C159 source.n76 a_n1878_n2088# 0.014122f
C160 source.n77 a_n1878_n2088# 0.106213f
C161 source.t20 a_n1878_n2088# 0.051381f
C162 source.n78 a_n1878_n2088# 0.023643f
C163 source.n79 a_n1878_n2088# 0.018621f
C164 source.n80 a_n1878_n2088# 0.013337f
C165 source.n81 a_n1878_n2088# 0.590571f
C166 source.n82 a_n1878_n2088# 0.02482f
C167 source.n83 a_n1878_n2088# 0.013337f
C168 source.n84 a_n1878_n2088# 0.014122f
C169 source.n85 a_n1878_n2088# 0.031524f
C170 source.n86 a_n1878_n2088# 0.031524f
C171 source.n87 a_n1878_n2088# 0.014122f
C172 source.n88 a_n1878_n2088# 0.013337f
C173 source.n89 a_n1878_n2088# 0.02482f
C174 source.n90 a_n1878_n2088# 0.02482f
C175 source.n91 a_n1878_n2088# 0.013337f
C176 source.n92 a_n1878_n2088# 0.014122f
C177 source.n93 a_n1878_n2088# 0.031524f
C178 source.n94 a_n1878_n2088# 0.068245f
C179 source.n95 a_n1878_n2088# 0.014122f
C180 source.n96 a_n1878_n2088# 0.013337f
C181 source.n97 a_n1878_n2088# 0.057371f
C182 source.n98 a_n1878_n2088# 0.038186f
C183 source.n99 a_n1878_n2088# 0.115997f
C184 source.t21 a_n1878_n2088# 0.117682f
C185 source.t2 a_n1878_n2088# 0.117682f
C186 source.n100 a_n1878_n2088# 0.916514f
C187 source.n101 a_n1878_n2088# 0.347113f
C188 source.t1 a_n1878_n2088# 0.117682f
C189 source.t23 a_n1878_n2088# 0.117682f
C190 source.n102 a_n1878_n2088# 0.916514f
C191 source.n103 a_n1878_n2088# 0.347113f
C192 source.n104 a_n1878_n2088# 0.034887f
C193 source.n105 a_n1878_n2088# 0.02482f
C194 source.n106 a_n1878_n2088# 0.013337f
C195 source.n107 a_n1878_n2088# 0.031524f
C196 source.n108 a_n1878_n2088# 0.014122f
C197 source.n109 a_n1878_n2088# 0.02482f
C198 source.n110 a_n1878_n2088# 0.013337f
C199 source.n111 a_n1878_n2088# 0.031524f
C200 source.n112 a_n1878_n2088# 0.014122f
C201 source.n113 a_n1878_n2088# 0.106213f
C202 source.t5 a_n1878_n2088# 0.051381f
C203 source.n114 a_n1878_n2088# 0.023643f
C204 source.n115 a_n1878_n2088# 0.018621f
C205 source.n116 a_n1878_n2088# 0.013337f
C206 source.n117 a_n1878_n2088# 0.590571f
C207 source.n118 a_n1878_n2088# 0.02482f
C208 source.n119 a_n1878_n2088# 0.013337f
C209 source.n120 a_n1878_n2088# 0.014122f
C210 source.n121 a_n1878_n2088# 0.031524f
C211 source.n122 a_n1878_n2088# 0.031524f
C212 source.n123 a_n1878_n2088# 0.014122f
C213 source.n124 a_n1878_n2088# 0.013337f
C214 source.n125 a_n1878_n2088# 0.02482f
C215 source.n126 a_n1878_n2088# 0.02482f
C216 source.n127 a_n1878_n2088# 0.013337f
C217 source.n128 a_n1878_n2088# 0.014122f
C218 source.n129 a_n1878_n2088# 0.031524f
C219 source.n130 a_n1878_n2088# 0.068245f
C220 source.n131 a_n1878_n2088# 0.014122f
C221 source.n132 a_n1878_n2088# 0.013337f
C222 source.n133 a_n1878_n2088# 0.057371f
C223 source.n134 a_n1878_n2088# 0.038186f
C224 source.n135 a_n1878_n2088# 0.948304f
C225 source.n136 a_n1878_n2088# 0.034887f
C226 source.n137 a_n1878_n2088# 0.02482f
C227 source.n138 a_n1878_n2088# 0.013337f
C228 source.n139 a_n1878_n2088# 0.031524f
C229 source.n140 a_n1878_n2088# 0.014122f
C230 source.n141 a_n1878_n2088# 0.02482f
C231 source.n142 a_n1878_n2088# 0.013337f
C232 source.n143 a_n1878_n2088# 0.031524f
C233 source.n144 a_n1878_n2088# 0.014122f
C234 source.n145 a_n1878_n2088# 0.106213f
C235 source.t19 a_n1878_n2088# 0.051381f
C236 source.n146 a_n1878_n2088# 0.023643f
C237 source.n147 a_n1878_n2088# 0.018621f
C238 source.n148 a_n1878_n2088# 0.013337f
C239 source.n149 a_n1878_n2088# 0.590571f
C240 source.n150 a_n1878_n2088# 0.02482f
C241 source.n151 a_n1878_n2088# 0.013337f
C242 source.n152 a_n1878_n2088# 0.014122f
C243 source.n153 a_n1878_n2088# 0.031524f
C244 source.n154 a_n1878_n2088# 0.031524f
C245 source.n155 a_n1878_n2088# 0.014122f
C246 source.n156 a_n1878_n2088# 0.013337f
C247 source.n157 a_n1878_n2088# 0.02482f
C248 source.n158 a_n1878_n2088# 0.02482f
C249 source.n159 a_n1878_n2088# 0.013337f
C250 source.n160 a_n1878_n2088# 0.014122f
C251 source.n161 a_n1878_n2088# 0.031524f
C252 source.n162 a_n1878_n2088# 0.068245f
C253 source.n163 a_n1878_n2088# 0.014122f
C254 source.n164 a_n1878_n2088# 0.013337f
C255 source.n165 a_n1878_n2088# 0.057371f
C256 source.n166 a_n1878_n2088# 0.038186f
C257 source.n167 a_n1878_n2088# 0.948304f
C258 source.t13 a_n1878_n2088# 0.117682f
C259 source.t14 a_n1878_n2088# 0.117682f
C260 source.n168 a_n1878_n2088# 0.916508f
C261 source.n169 a_n1878_n2088# 0.347119f
C262 source.t9 a_n1878_n2088# 0.117682f
C263 source.t15 a_n1878_n2088# 0.117682f
C264 source.n170 a_n1878_n2088# 0.916508f
C265 source.n171 a_n1878_n2088# 0.347119f
C266 source.n172 a_n1878_n2088# 0.034887f
C267 source.n173 a_n1878_n2088# 0.02482f
C268 source.n174 a_n1878_n2088# 0.013337f
C269 source.n175 a_n1878_n2088# 0.031524f
C270 source.n176 a_n1878_n2088# 0.014122f
C271 source.n177 a_n1878_n2088# 0.02482f
C272 source.n178 a_n1878_n2088# 0.013337f
C273 source.n179 a_n1878_n2088# 0.031524f
C274 source.n180 a_n1878_n2088# 0.014122f
C275 source.n181 a_n1878_n2088# 0.106213f
C276 source.t16 a_n1878_n2088# 0.051381f
C277 source.n182 a_n1878_n2088# 0.023643f
C278 source.n183 a_n1878_n2088# 0.018621f
C279 source.n184 a_n1878_n2088# 0.013337f
C280 source.n185 a_n1878_n2088# 0.590571f
C281 source.n186 a_n1878_n2088# 0.02482f
C282 source.n187 a_n1878_n2088# 0.013337f
C283 source.n188 a_n1878_n2088# 0.014122f
C284 source.n189 a_n1878_n2088# 0.031524f
C285 source.n190 a_n1878_n2088# 0.031524f
C286 source.n191 a_n1878_n2088# 0.014122f
C287 source.n192 a_n1878_n2088# 0.013337f
C288 source.n193 a_n1878_n2088# 0.02482f
C289 source.n194 a_n1878_n2088# 0.02482f
C290 source.n195 a_n1878_n2088# 0.013337f
C291 source.n196 a_n1878_n2088# 0.014122f
C292 source.n197 a_n1878_n2088# 0.031524f
C293 source.n198 a_n1878_n2088# 0.068245f
C294 source.n199 a_n1878_n2088# 0.014122f
C295 source.n200 a_n1878_n2088# 0.013337f
C296 source.n201 a_n1878_n2088# 0.057371f
C297 source.n202 a_n1878_n2088# 0.038186f
C298 source.n203 a_n1878_n2088# 0.115997f
C299 source.n204 a_n1878_n2088# 0.034887f
C300 source.n205 a_n1878_n2088# 0.02482f
C301 source.n206 a_n1878_n2088# 0.013337f
C302 source.n207 a_n1878_n2088# 0.031524f
C303 source.n208 a_n1878_n2088# 0.014122f
C304 source.n209 a_n1878_n2088# 0.02482f
C305 source.n210 a_n1878_n2088# 0.013337f
C306 source.n211 a_n1878_n2088# 0.031524f
C307 source.n212 a_n1878_n2088# 0.014122f
C308 source.n213 a_n1878_n2088# 0.106213f
C309 source.t0 a_n1878_n2088# 0.051381f
C310 source.n214 a_n1878_n2088# 0.023643f
C311 source.n215 a_n1878_n2088# 0.018621f
C312 source.n216 a_n1878_n2088# 0.013337f
C313 source.n217 a_n1878_n2088# 0.590571f
C314 source.n218 a_n1878_n2088# 0.02482f
C315 source.n219 a_n1878_n2088# 0.013337f
C316 source.n220 a_n1878_n2088# 0.014122f
C317 source.n221 a_n1878_n2088# 0.031524f
C318 source.n222 a_n1878_n2088# 0.031524f
C319 source.n223 a_n1878_n2088# 0.014122f
C320 source.n224 a_n1878_n2088# 0.013337f
C321 source.n225 a_n1878_n2088# 0.02482f
C322 source.n226 a_n1878_n2088# 0.02482f
C323 source.n227 a_n1878_n2088# 0.013337f
C324 source.n228 a_n1878_n2088# 0.014122f
C325 source.n229 a_n1878_n2088# 0.031524f
C326 source.n230 a_n1878_n2088# 0.068245f
C327 source.n231 a_n1878_n2088# 0.014122f
C328 source.n232 a_n1878_n2088# 0.013337f
C329 source.n233 a_n1878_n2088# 0.057371f
C330 source.n234 a_n1878_n2088# 0.038186f
C331 source.n235 a_n1878_n2088# 0.115997f
C332 source.t7 a_n1878_n2088# 0.117682f
C333 source.t3 a_n1878_n2088# 0.117682f
C334 source.n236 a_n1878_n2088# 0.916508f
C335 source.n237 a_n1878_n2088# 0.347119f
C336 source.t22 a_n1878_n2088# 0.117682f
C337 source.t4 a_n1878_n2088# 0.117682f
C338 source.n238 a_n1878_n2088# 0.916508f
C339 source.n239 a_n1878_n2088# 0.347119f
C340 source.n240 a_n1878_n2088# 0.034887f
C341 source.n241 a_n1878_n2088# 0.02482f
C342 source.n242 a_n1878_n2088# 0.013337f
C343 source.n243 a_n1878_n2088# 0.031524f
C344 source.n244 a_n1878_n2088# 0.014122f
C345 source.n245 a_n1878_n2088# 0.02482f
C346 source.n246 a_n1878_n2088# 0.013337f
C347 source.n247 a_n1878_n2088# 0.031524f
C348 source.n248 a_n1878_n2088# 0.014122f
C349 source.n249 a_n1878_n2088# 0.106213f
C350 source.t6 a_n1878_n2088# 0.051381f
C351 source.n250 a_n1878_n2088# 0.023643f
C352 source.n251 a_n1878_n2088# 0.018621f
C353 source.n252 a_n1878_n2088# 0.013337f
C354 source.n253 a_n1878_n2088# 0.590571f
C355 source.n254 a_n1878_n2088# 0.02482f
C356 source.n255 a_n1878_n2088# 0.013337f
C357 source.n256 a_n1878_n2088# 0.014122f
C358 source.n257 a_n1878_n2088# 0.031524f
C359 source.n258 a_n1878_n2088# 0.031524f
C360 source.n259 a_n1878_n2088# 0.014122f
C361 source.n260 a_n1878_n2088# 0.013337f
C362 source.n261 a_n1878_n2088# 0.02482f
C363 source.n262 a_n1878_n2088# 0.02482f
C364 source.n263 a_n1878_n2088# 0.013337f
C365 source.n264 a_n1878_n2088# 0.014122f
C366 source.n265 a_n1878_n2088# 0.031524f
C367 source.n266 a_n1878_n2088# 0.068245f
C368 source.n267 a_n1878_n2088# 0.014122f
C369 source.n268 a_n1878_n2088# 0.013337f
C370 source.n269 a_n1878_n2088# 0.057371f
C371 source.n270 a_n1878_n2088# 0.038186f
C372 source.n271 a_n1878_n2088# 0.267065f
C373 source.n272 a_n1878_n2088# 1.02238f
C374 drain_left.t0 a_n1878_n2088# 0.13679f
C375 drain_left.t3 a_n1878_n2088# 0.13679f
C376 drain_left.n0 a_n1878_n2088# 1.14448f
C377 drain_left.t2 a_n1878_n2088# 0.13679f
C378 drain_left.t10 a_n1878_n2088# 0.13679f
C379 drain_left.n1 a_n1878_n2088# 1.14083f
C380 drain_left.t6 a_n1878_n2088# 0.13679f
C381 drain_left.t1 a_n1878_n2088# 0.13679f
C382 drain_left.n2 a_n1878_n2088# 1.14448f
C383 drain_left.n3 a_n1878_n2088# 2.10523f
C384 drain_left.t4 a_n1878_n2088# 0.13679f
C385 drain_left.t7 a_n1878_n2088# 0.13679f
C386 drain_left.n4 a_n1878_n2088# 1.14483f
C387 drain_left.t9 a_n1878_n2088# 0.13679f
C388 drain_left.t5 a_n1878_n2088# 0.13679f
C389 drain_left.n5 a_n1878_n2088# 1.14084f
C390 drain_left.n6 a_n1878_n2088# 0.742f
C391 drain_left.t8 a_n1878_n2088# 0.13679f
C392 drain_left.t11 a_n1878_n2088# 0.13679f
C393 drain_left.n7 a_n1878_n2088# 1.14083f
C394 drain_left.n8 a_n1878_n2088# 0.615055f
C395 plus.n0 a_n1878_n2088# 0.04864f
C396 plus.t11 a_n1878_n2088# 0.423252f
C397 plus.t8 a_n1878_n2088# 0.423252f
C398 plus.n1 a_n1878_n2088# 0.04864f
C399 plus.t2 a_n1878_n2088# 0.423252f
C400 plus.n2 a_n1878_n2088# 0.04864f
C401 plus.t9 a_n1878_n2088# 0.423252f
C402 plus.n3 a_n1878_n2088# 0.204325f
C403 plus.t7 a_n1878_n2088# 0.423252f
C404 plus.n4 a_n1878_n2088# 0.210188f
C405 plus.t1 a_n1878_n2088# 0.436736f
C406 plus.n5 a_n1878_n2088# 0.187084f
C407 plus.n6 a_n1878_n2088# 0.198094f
C408 plus.n7 a_n1878_n2088# 0.04864f
C409 plus.n8 a_n1878_n2088# 0.011038f
C410 plus.n9 a_n1878_n2088# 0.204325f
C411 plus.n10 a_n1878_n2088# 0.199527f
C412 plus.n11 a_n1878_n2088# 0.011038f
C413 plus.n12 a_n1878_n2088# 0.199227f
C414 plus.n13 a_n1878_n2088# 0.420474f
C415 plus.n14 a_n1878_n2088# 0.04864f
C416 plus.t0 a_n1878_n2088# 0.423252f
C417 plus.n15 a_n1878_n2088# 0.04864f
C418 plus.t6 a_n1878_n2088# 0.423252f
C419 plus.n16 a_n1878_n2088# 0.04864f
C420 plus.t5 a_n1878_n2088# 0.423252f
C421 plus.t10 a_n1878_n2088# 0.423252f
C422 plus.n17 a_n1878_n2088# 0.204325f
C423 plus.t3 a_n1878_n2088# 0.436736f
C424 plus.t4 a_n1878_n2088# 0.423252f
C425 plus.n18 a_n1878_n2088# 0.210188f
C426 plus.n19 a_n1878_n2088# 0.187084f
C427 plus.n20 a_n1878_n2088# 0.198094f
C428 plus.n21 a_n1878_n2088# 0.04864f
C429 plus.n22 a_n1878_n2088# 0.011038f
C430 plus.n23 a_n1878_n2088# 0.204325f
C431 plus.n24 a_n1878_n2088# 0.199527f
C432 plus.n25 a_n1878_n2088# 0.011038f
C433 plus.n26 a_n1878_n2088# 0.199227f
C434 plus.n27 a_n1878_n2088# 1.25705f
.ends

