* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X1 drain_left.t19 plus.t0 source.t19 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X2 drain_right.t19 minus.t0 source.t14 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X3 drain_right.t18 minus.t1 source.t1 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X4 source.t8 minus.t2 drain_right.t17 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X5 drain_right.t16 minus.t3 source.t10 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X6 source.t27 plus.t1 drain_left.t18 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X7 a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X8 source.t20 plus.t2 drain_left.t17 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X9 drain_left.t16 plus.t3 source.t24 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X10 source.t11 minus.t4 drain_right.t15 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X11 drain_left.t15 plus.t4 source.t33 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X12 source.t5 minus.t5 drain_right.t14 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X13 drain_right.t13 minus.t6 source.t4 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X14 source.t13 minus.t7 drain_right.t12 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X15 drain_left.t14 plus.t5 source.t30 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X16 drain_left.t13 plus.t6 source.t31 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X17 source.t12 minus.t8 drain_right.t11 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X18 drain_left.t12 plus.t7 source.t21 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X19 source.t15 minus.t9 drain_right.t10 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X20 drain_left.t11 plus.t8 source.t18 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X21 source.t23 plus.t9 drain_left.t10 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X22 drain_right.t9 minus.t10 source.t3 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X23 source.t36 plus.t10 drain_left.t9 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X24 source.t35 plus.t11 drain_left.t8 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X25 source.t28 plus.t12 drain_left.t7 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X26 drain_right.t8 minus.t11 source.t6 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X27 drain_right.t7 minus.t12 source.t2 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X28 drain_right.t6 minus.t13 source.t0 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X29 drain_right.t5 minus.t14 source.t17 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X30 source.t29 plus.t13 drain_left.t6 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X31 drain_left.t5 plus.t14 source.t32 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X32 a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X33 source.t26 plus.t15 drain_left.t4 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X34 drain_left.t3 plus.t16 source.t37 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X35 source.t16 minus.t15 drain_right.t4 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X36 source.t9 minus.t16 drain_right.t3 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X37 source.t7 minus.t17 drain_right.t2 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X38 drain_right.t1 minus.t18 source.t38 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X39 source.t34 plus.t17 drain_left.t2 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X40 drain_left.t1 plus.t18 source.t25 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X41 source.t22 plus.t19 drain_left.t0 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X42 a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X43 source.t39 minus.t19 drain_right.t0 a_n1882_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n5 plus.t9 574.384
R1 plus.n23 plus.t6 574.384
R2 plus.n30 plus.t4 574.384
R3 plus.n48 plus.t12 574.384
R4 plus.n6 plus.t3 518.15
R5 plus.n8 plus.t19 518.15
R6 plus.n3 plus.t16 518.15
R7 plus.n13 plus.t15 518.15
R8 plus.n15 plus.t8 518.15
R9 plus.n1 plus.t2 518.15
R10 plus.n20 plus.t18 518.15
R11 plus.n22 plus.t13 518.15
R12 plus.n31 plus.t11 518.15
R13 plus.n33 plus.t0 518.15
R14 plus.n28 plus.t10 518.15
R15 plus.n38 plus.t14 518.15
R16 plus.n40 plus.t1 518.15
R17 plus.n26 plus.t7 518.15
R18 plus.n45 plus.t17 518.15
R19 plus.n47 plus.t5 518.15
R20 plus.n5 plus.n4 161.489
R21 plus.n30 plus.n29 161.489
R22 plus.n7 plus.n4 161.3
R23 plus.n10 plus.n9 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n2 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n0 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n32 plus.n29 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n36 161.3
R33 plus.n39 plus.n27 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n25 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n7 plus.n6 51.852
R39 plus.n22 plus.n21 51.852
R40 plus.n47 plus.n46 51.852
R41 plus.n32 plus.n31 51.852
R42 plus.n9 plus.n8 47.4702
R43 plus.n20 plus.n19 47.4702
R44 plus.n45 plus.n44 47.4702
R45 plus.n34 plus.n33 47.4702
R46 plus.n12 plus.n3 43.0884
R47 plus.n16 plus.n1 43.0884
R48 plus.n41 plus.n26 43.0884
R49 plus.n37 plus.n28 43.0884
R50 plus.n14 plus.n13 38.7066
R51 plus.n15 plus.n14 38.7066
R52 plus.n40 plus.n39 38.7066
R53 plus.n39 plus.n38 38.7066
R54 plus.n13 plus.n12 34.3247
R55 plus.n16 plus.n15 34.3247
R56 plus.n41 plus.n40 34.3247
R57 plus.n38 plus.n37 34.3247
R58 plus.n9 plus.n3 29.9429
R59 plus.n19 plus.n1 29.9429
R60 plus.n44 plus.n26 29.9429
R61 plus.n34 plus.n28 29.9429
R62 plus plus.n49 26.6998
R63 plus.n8 plus.n7 25.5611
R64 plus.n21 plus.n20 25.5611
R65 plus.n46 plus.n45 25.5611
R66 plus.n33 plus.n32 25.5611
R67 plus.n6 plus.n5 21.1793
R68 plus.n23 plus.n22 21.1793
R69 plus.n48 plus.n47 21.1793
R70 plus.n31 plus.n30 21.1793
R71 plus plus.n24 8.71262
R72 plus.n10 plus.n4 0.189894
R73 plus.n11 plus.n10 0.189894
R74 plus.n11 plus.n2 0.189894
R75 plus.n17 plus.n2 0.189894
R76 plus.n18 plus.n17 0.189894
R77 plus.n18 plus.n0 0.189894
R78 plus.n24 plus.n0 0.189894
R79 plus.n49 plus.n25 0.189894
R80 plus.n43 plus.n25 0.189894
R81 plus.n43 plus.n42 0.189894
R82 plus.n42 plus.n27 0.189894
R83 plus.n36 plus.n27 0.189894
R84 plus.n36 plus.n35 0.189894
R85 plus.n35 plus.n29 0.189894
R86 source.n0 source.t31 69.6943
R87 source.n9 source.t23 69.6943
R88 source.n10 source.t0 69.6943
R89 source.n19 source.t15 69.6943
R90 source.n39 source.t4 69.6942
R91 source.n30 source.t11 69.6942
R92 source.n29 source.t33 69.6942
R93 source.n20 source.t28 69.6942
R94 source.n2 source.n1 63.0943
R95 source.n4 source.n3 63.0943
R96 source.n6 source.n5 63.0943
R97 source.n8 source.n7 63.0943
R98 source.n12 source.n11 63.0943
R99 source.n14 source.n13 63.0943
R100 source.n16 source.n15 63.0943
R101 source.n18 source.n17 63.0943
R102 source.n38 source.n37 63.0942
R103 source.n36 source.n35 63.0942
R104 source.n34 source.n33 63.0942
R105 source.n32 source.n31 63.0942
R106 source.n28 source.n27 63.0942
R107 source.n26 source.n25 63.0942
R108 source.n24 source.n23 63.0942
R109 source.n22 source.n21 63.0942
R110 source.n20 source.n19 14.9264
R111 source.n40 source.n0 9.43506
R112 source.n37 source.t2 6.6005
R113 source.n37 source.t7 6.6005
R114 source.n35 source.t38 6.6005
R115 source.n35 source.t8 6.6005
R116 source.n33 source.t10 6.6005
R117 source.n33 source.t12 6.6005
R118 source.n31 source.t3 6.6005
R119 source.n31 source.t39 6.6005
R120 source.n27 source.t19 6.6005
R121 source.n27 source.t35 6.6005
R122 source.n25 source.t32 6.6005
R123 source.n25 source.t36 6.6005
R124 source.n23 source.t21 6.6005
R125 source.n23 source.t27 6.6005
R126 source.n21 source.t30 6.6005
R127 source.n21 source.t34 6.6005
R128 source.n1 source.t25 6.6005
R129 source.n1 source.t29 6.6005
R130 source.n3 source.t18 6.6005
R131 source.n3 source.t20 6.6005
R132 source.n5 source.t37 6.6005
R133 source.n5 source.t26 6.6005
R134 source.n7 source.t24 6.6005
R135 source.n7 source.t22 6.6005
R136 source.n11 source.t14 6.6005
R137 source.n11 source.t13 6.6005
R138 source.n13 source.t17 6.6005
R139 source.n13 source.t16 6.6005
R140 source.n15 source.t1 6.6005
R141 source.n15 source.t5 6.6005
R142 source.n17 source.t6 6.6005
R143 source.n17 source.t9 6.6005
R144 source.n40 source.n39 5.49188
R145 source.n10 source.n9 0.470328
R146 source.n30 source.n29 0.470328
R147 source.n19 source.n18 0.457397
R148 source.n18 source.n16 0.457397
R149 source.n16 source.n14 0.457397
R150 source.n14 source.n12 0.457397
R151 source.n12 source.n10 0.457397
R152 source.n9 source.n8 0.457397
R153 source.n8 source.n6 0.457397
R154 source.n6 source.n4 0.457397
R155 source.n4 source.n2 0.457397
R156 source.n2 source.n0 0.457397
R157 source.n22 source.n20 0.457397
R158 source.n24 source.n22 0.457397
R159 source.n26 source.n24 0.457397
R160 source.n28 source.n26 0.457397
R161 source.n29 source.n28 0.457397
R162 source.n32 source.n30 0.457397
R163 source.n34 source.n32 0.457397
R164 source.n36 source.n34 0.457397
R165 source.n38 source.n36 0.457397
R166 source.n39 source.n38 0.457397
R167 source source.n40 0.188
R168 drain_left.n10 drain_left.n8 80.23
R169 drain_left.n6 drain_left.n4 80.2299
R170 drain_left.n2 drain_left.n0 80.2299
R171 drain_left.n16 drain_left.n15 79.7731
R172 drain_left.n14 drain_left.n13 79.7731
R173 drain_left.n12 drain_left.n11 79.7731
R174 drain_left.n10 drain_left.n9 79.7731
R175 drain_left.n7 drain_left.n3 79.773
R176 drain_left.n6 drain_left.n5 79.773
R177 drain_left.n2 drain_left.n1 79.773
R178 drain_left drain_left.n7 24.2041
R179 drain_left.n3 drain_left.t18 6.6005
R180 drain_left.n3 drain_left.t5 6.6005
R181 drain_left.n4 drain_left.t8 6.6005
R182 drain_left.n4 drain_left.t15 6.6005
R183 drain_left.n5 drain_left.t9 6.6005
R184 drain_left.n5 drain_left.t19 6.6005
R185 drain_left.n1 drain_left.t2 6.6005
R186 drain_left.n1 drain_left.t12 6.6005
R187 drain_left.n0 drain_left.t7 6.6005
R188 drain_left.n0 drain_left.t14 6.6005
R189 drain_left.n15 drain_left.t6 6.6005
R190 drain_left.n15 drain_left.t13 6.6005
R191 drain_left.n13 drain_left.t17 6.6005
R192 drain_left.n13 drain_left.t1 6.6005
R193 drain_left.n11 drain_left.t4 6.6005
R194 drain_left.n11 drain_left.t11 6.6005
R195 drain_left.n9 drain_left.t0 6.6005
R196 drain_left.n9 drain_left.t3 6.6005
R197 drain_left.n8 drain_left.t10 6.6005
R198 drain_left.n8 drain_left.t16 6.6005
R199 drain_left drain_left.n16 6.11011
R200 drain_left.n12 drain_left.n10 0.457397
R201 drain_left.n14 drain_left.n12 0.457397
R202 drain_left.n16 drain_left.n14 0.457397
R203 drain_left.n7 drain_left.n6 0.402051
R204 drain_left.n7 drain_left.n2 0.402051
R205 minus.n23 minus.t9 574.384
R206 minus.n5 minus.t13 574.384
R207 minus.n48 minus.t6 574.384
R208 minus.n30 minus.t4 574.384
R209 minus.n22 minus.t11 518.15
R210 minus.n20 minus.t16 518.15
R211 minus.n1 minus.t1 518.15
R212 minus.n15 minus.t5 518.15
R213 minus.n13 minus.t14 518.15
R214 minus.n3 minus.t15 518.15
R215 minus.n8 minus.t0 518.15
R216 minus.n6 minus.t7 518.15
R217 minus.n47 minus.t17 518.15
R218 minus.n45 minus.t12 518.15
R219 minus.n26 minus.t2 518.15
R220 minus.n40 minus.t18 518.15
R221 minus.n38 minus.t8 518.15
R222 minus.n28 minus.t3 518.15
R223 minus.n33 minus.t19 518.15
R224 minus.n31 minus.t10 518.15
R225 minus.n5 minus.n4 161.489
R226 minus.n30 minus.n29 161.489
R227 minus.n24 minus.n23 161.3
R228 minus.n21 minus.n0 161.3
R229 minus.n19 minus.n18 161.3
R230 minus.n17 minus.n16 161.3
R231 minus.n14 minus.n2 161.3
R232 minus.n12 minus.n11 161.3
R233 minus.n10 minus.n9 161.3
R234 minus.n7 minus.n4 161.3
R235 minus.n49 minus.n48 161.3
R236 minus.n46 minus.n25 161.3
R237 minus.n44 minus.n43 161.3
R238 minus.n42 minus.n41 161.3
R239 minus.n39 minus.n27 161.3
R240 minus.n37 minus.n36 161.3
R241 minus.n35 minus.n34 161.3
R242 minus.n32 minus.n29 161.3
R243 minus.n22 minus.n21 51.852
R244 minus.n7 minus.n6 51.852
R245 minus.n32 minus.n31 51.852
R246 minus.n47 minus.n46 51.852
R247 minus.n20 minus.n19 47.4702
R248 minus.n9 minus.n8 47.4702
R249 minus.n34 minus.n33 47.4702
R250 minus.n45 minus.n44 47.4702
R251 minus.n16 minus.n1 43.0884
R252 minus.n12 minus.n3 43.0884
R253 minus.n37 minus.n28 43.0884
R254 minus.n41 minus.n26 43.0884
R255 minus.n15 minus.n14 38.7066
R256 minus.n14 minus.n13 38.7066
R257 minus.n39 minus.n38 38.7066
R258 minus.n40 minus.n39 38.7066
R259 minus.n16 minus.n15 34.3247
R260 minus.n13 minus.n12 34.3247
R261 minus.n38 minus.n37 34.3247
R262 minus.n41 minus.n40 34.3247
R263 minus.n19 minus.n1 29.9429
R264 minus.n9 minus.n3 29.9429
R265 minus.n34 minus.n28 29.9429
R266 minus.n44 minus.n26 29.9429
R267 minus.n50 minus.n24 29.4096
R268 minus.n21 minus.n20 25.5611
R269 minus.n8 minus.n7 25.5611
R270 minus.n33 minus.n32 25.5611
R271 minus.n46 minus.n45 25.5611
R272 minus.n23 minus.n22 21.1793
R273 minus.n6 minus.n5 21.1793
R274 minus.n31 minus.n30 21.1793
R275 minus.n48 minus.n47 21.1793
R276 minus.n50 minus.n49 6.47777
R277 minus.n24 minus.n0 0.189894
R278 minus.n18 minus.n0 0.189894
R279 minus.n18 minus.n17 0.189894
R280 minus.n17 minus.n2 0.189894
R281 minus.n11 minus.n2 0.189894
R282 minus.n11 minus.n10 0.189894
R283 minus.n10 minus.n4 0.189894
R284 minus.n35 minus.n29 0.189894
R285 minus.n36 minus.n35 0.189894
R286 minus.n36 minus.n27 0.189894
R287 minus.n42 minus.n27 0.189894
R288 minus.n43 minus.n42 0.189894
R289 minus.n43 minus.n25 0.189894
R290 minus.n49 minus.n25 0.189894
R291 minus minus.n50 0.188
R292 drain_right.n10 drain_right.n8 80.23
R293 drain_right.n6 drain_right.n4 80.2299
R294 drain_right.n2 drain_right.n0 80.2299
R295 drain_right.n10 drain_right.n9 79.7731
R296 drain_right.n12 drain_right.n11 79.7731
R297 drain_right.n14 drain_right.n13 79.7731
R298 drain_right.n16 drain_right.n15 79.7731
R299 drain_right.n7 drain_right.n3 79.773
R300 drain_right.n6 drain_right.n5 79.773
R301 drain_right.n2 drain_right.n1 79.773
R302 drain_right drain_right.n7 23.6508
R303 drain_right.n3 drain_right.t11 6.6005
R304 drain_right.n3 drain_right.t1 6.6005
R305 drain_right.n4 drain_right.t2 6.6005
R306 drain_right.n4 drain_right.t13 6.6005
R307 drain_right.n5 drain_right.t17 6.6005
R308 drain_right.n5 drain_right.t7 6.6005
R309 drain_right.n1 drain_right.t0 6.6005
R310 drain_right.n1 drain_right.t16 6.6005
R311 drain_right.n0 drain_right.t15 6.6005
R312 drain_right.n0 drain_right.t9 6.6005
R313 drain_right.n8 drain_right.t12 6.6005
R314 drain_right.n8 drain_right.t6 6.6005
R315 drain_right.n9 drain_right.t4 6.6005
R316 drain_right.n9 drain_right.t19 6.6005
R317 drain_right.n11 drain_right.t14 6.6005
R318 drain_right.n11 drain_right.t5 6.6005
R319 drain_right.n13 drain_right.t3 6.6005
R320 drain_right.n13 drain_right.t18 6.6005
R321 drain_right.n15 drain_right.t10 6.6005
R322 drain_right.n15 drain_right.t8 6.6005
R323 drain_right drain_right.n16 6.11011
R324 drain_right.n16 drain_right.n14 0.457397
R325 drain_right.n14 drain_right.n12 0.457397
R326 drain_right.n12 drain_right.n10 0.457397
R327 drain_right.n7 drain_right.n6 0.402051
R328 drain_right.n7 drain_right.n2 0.402051
C0 drain_left minus 0.176325f
C1 drain_left plus 1.94529f
C2 drain_right minus 1.76222f
C3 drain_right plus 0.342781f
C4 source minus 1.86521f
C5 source plus 1.8792f
C6 drain_left drain_right 0.982057f
C7 source drain_left 13.6851f
C8 plus minus 3.84182f
C9 source drain_right 13.6851f
C10 drain_right a_n1882_n1488# 4.56526f
C11 drain_left a_n1882_n1488# 4.83651f
C12 source a_n1882_n1488# 3.695944f
C13 minus a_n1882_n1488# 6.586923f
C14 plus a_n1882_n1488# 7.216204f
C15 drain_right.t15 a_n1882_n1488# 0.076803f
C16 drain_right.t9 a_n1882_n1488# 0.076803f
C17 drain_right.n0 a_n1882_n1488# 0.555993f
C18 drain_right.t0 a_n1882_n1488# 0.076803f
C19 drain_right.t16 a_n1882_n1488# 0.076803f
C20 drain_right.n1 a_n1882_n1488# 0.553899f
C21 drain_right.n2 a_n1882_n1488# 0.716497f
C22 drain_right.t11 a_n1882_n1488# 0.076803f
C23 drain_right.t1 a_n1882_n1488# 0.076803f
C24 drain_right.n3 a_n1882_n1488# 0.553899f
C25 drain_right.t2 a_n1882_n1488# 0.076803f
C26 drain_right.t13 a_n1882_n1488# 0.076803f
C27 drain_right.n4 a_n1882_n1488# 0.555993f
C28 drain_right.t17 a_n1882_n1488# 0.076803f
C29 drain_right.t7 a_n1882_n1488# 0.076803f
C30 drain_right.n5 a_n1882_n1488# 0.553899f
C31 drain_right.n6 a_n1882_n1488# 0.716497f
C32 drain_right.n7 a_n1882_n1488# 1.23116f
C33 drain_right.t12 a_n1882_n1488# 0.076803f
C34 drain_right.t6 a_n1882_n1488# 0.076803f
C35 drain_right.n8 a_n1882_n1488# 0.555996f
C36 drain_right.t4 a_n1882_n1488# 0.076803f
C37 drain_right.t19 a_n1882_n1488# 0.076803f
C38 drain_right.n9 a_n1882_n1488# 0.553901f
C39 drain_right.n10 a_n1882_n1488# 0.720399f
C40 drain_right.t14 a_n1882_n1488# 0.076803f
C41 drain_right.t5 a_n1882_n1488# 0.076803f
C42 drain_right.n11 a_n1882_n1488# 0.553901f
C43 drain_right.n12 a_n1882_n1488# 0.354722f
C44 drain_right.t3 a_n1882_n1488# 0.076803f
C45 drain_right.t18 a_n1882_n1488# 0.076803f
C46 drain_right.n13 a_n1882_n1488# 0.553901f
C47 drain_right.n14 a_n1882_n1488# 0.354722f
C48 drain_right.t10 a_n1882_n1488# 0.076803f
C49 drain_right.t8 a_n1882_n1488# 0.076803f
C50 drain_right.n15 a_n1882_n1488# 0.553901f
C51 drain_right.n16 a_n1882_n1488# 0.619862f
C52 minus.n0 a_n1882_n1488# 0.026502f
C53 minus.t9 a_n1882_n1488# 0.049069f
C54 minus.t11 a_n1882_n1488# 0.046048f
C55 minus.t16 a_n1882_n1488# 0.046048f
C56 minus.t1 a_n1882_n1488# 0.046048f
C57 minus.n1 a_n1882_n1488# 0.029461f
C58 minus.n2 a_n1882_n1488# 0.026502f
C59 minus.t5 a_n1882_n1488# 0.046048f
C60 minus.t14 a_n1882_n1488# 0.046048f
C61 minus.t15 a_n1882_n1488# 0.046048f
C62 minus.n3 a_n1882_n1488# 0.029461f
C63 minus.n4 a_n1882_n1488# 0.060644f
C64 minus.t0 a_n1882_n1488# 0.046048f
C65 minus.t7 a_n1882_n1488# 0.046048f
C66 minus.t13 a_n1882_n1488# 0.049069f
C67 minus.n5 a_n1882_n1488# 0.037152f
C68 minus.n6 a_n1882_n1488# 0.029461f
C69 minus.n7 a_n1882_n1488# 0.009282f
C70 minus.n8 a_n1882_n1488# 0.029461f
C71 minus.n9 a_n1882_n1488# 0.009282f
C72 minus.n10 a_n1882_n1488# 0.026502f
C73 minus.n11 a_n1882_n1488# 0.026502f
C74 minus.n12 a_n1882_n1488# 0.009282f
C75 minus.n13 a_n1882_n1488# 0.029461f
C76 minus.n14 a_n1882_n1488# 0.009282f
C77 minus.n15 a_n1882_n1488# 0.029461f
C78 minus.n16 a_n1882_n1488# 0.009282f
C79 minus.n17 a_n1882_n1488# 0.026502f
C80 minus.n18 a_n1882_n1488# 0.026502f
C81 minus.n19 a_n1882_n1488# 0.009282f
C82 minus.n20 a_n1882_n1488# 0.029461f
C83 minus.n21 a_n1882_n1488# 0.009282f
C84 minus.n22 a_n1882_n1488# 0.029461f
C85 minus.n23 a_n1882_n1488# 0.037112f
C86 minus.n24 a_n1882_n1488# 0.665752f
C87 minus.n25 a_n1882_n1488# 0.026502f
C88 minus.t17 a_n1882_n1488# 0.046048f
C89 minus.t12 a_n1882_n1488# 0.046048f
C90 minus.t2 a_n1882_n1488# 0.046048f
C91 minus.n26 a_n1882_n1488# 0.029461f
C92 minus.n27 a_n1882_n1488# 0.026502f
C93 minus.t18 a_n1882_n1488# 0.046048f
C94 minus.t8 a_n1882_n1488# 0.046048f
C95 minus.t3 a_n1882_n1488# 0.046048f
C96 minus.n28 a_n1882_n1488# 0.029461f
C97 minus.n29 a_n1882_n1488# 0.060644f
C98 minus.t19 a_n1882_n1488# 0.046048f
C99 minus.t10 a_n1882_n1488# 0.046048f
C100 minus.t4 a_n1882_n1488# 0.049069f
C101 minus.n30 a_n1882_n1488# 0.037152f
C102 minus.n31 a_n1882_n1488# 0.029461f
C103 minus.n32 a_n1882_n1488# 0.009282f
C104 minus.n33 a_n1882_n1488# 0.029461f
C105 minus.n34 a_n1882_n1488# 0.009282f
C106 minus.n35 a_n1882_n1488# 0.026502f
C107 minus.n36 a_n1882_n1488# 0.026502f
C108 minus.n37 a_n1882_n1488# 0.009282f
C109 minus.n38 a_n1882_n1488# 0.029461f
C110 minus.n39 a_n1882_n1488# 0.009282f
C111 minus.n40 a_n1882_n1488# 0.029461f
C112 minus.n41 a_n1882_n1488# 0.009282f
C113 minus.n42 a_n1882_n1488# 0.026502f
C114 minus.n43 a_n1882_n1488# 0.026502f
C115 minus.n44 a_n1882_n1488# 0.009282f
C116 minus.n45 a_n1882_n1488# 0.029461f
C117 minus.n46 a_n1882_n1488# 0.009282f
C118 minus.n47 a_n1882_n1488# 0.029461f
C119 minus.t6 a_n1882_n1488# 0.049069f
C120 minus.n48 a_n1882_n1488# 0.037112f
C121 minus.n49 a_n1882_n1488# 0.171875f
C122 minus.n50 a_n1882_n1488# 0.822758f
C123 drain_left.t7 a_n1882_n1488# 0.0761f
C124 drain_left.t14 a_n1882_n1488# 0.0761f
C125 drain_left.n0 a_n1882_n1488# 0.550897f
C126 drain_left.t2 a_n1882_n1488# 0.0761f
C127 drain_left.t12 a_n1882_n1488# 0.0761f
C128 drain_left.n1 a_n1882_n1488# 0.548822f
C129 drain_left.n2 a_n1882_n1488# 0.70993f
C130 drain_left.t18 a_n1882_n1488# 0.0761f
C131 drain_left.t5 a_n1882_n1488# 0.0761f
C132 drain_left.n3 a_n1882_n1488# 0.548822f
C133 drain_left.t8 a_n1882_n1488# 0.0761f
C134 drain_left.t15 a_n1882_n1488# 0.0761f
C135 drain_left.n4 a_n1882_n1488# 0.550897f
C136 drain_left.t9 a_n1882_n1488# 0.0761f
C137 drain_left.t19 a_n1882_n1488# 0.0761f
C138 drain_left.n5 a_n1882_n1488# 0.548822f
C139 drain_left.n6 a_n1882_n1488# 0.70993f
C140 drain_left.n7 a_n1882_n1488# 1.28343f
C141 drain_left.t10 a_n1882_n1488# 0.0761f
C142 drain_left.t16 a_n1882_n1488# 0.0761f
C143 drain_left.n8 a_n1882_n1488# 0.5509f
C144 drain_left.t0 a_n1882_n1488# 0.0761f
C145 drain_left.t3 a_n1882_n1488# 0.0761f
C146 drain_left.n9 a_n1882_n1488# 0.548824f
C147 drain_left.n10 a_n1882_n1488# 0.713796f
C148 drain_left.t4 a_n1882_n1488# 0.0761f
C149 drain_left.t11 a_n1882_n1488# 0.0761f
C150 drain_left.n11 a_n1882_n1488# 0.548824f
C151 drain_left.n12 a_n1882_n1488# 0.351471f
C152 drain_left.t17 a_n1882_n1488# 0.0761f
C153 drain_left.t1 a_n1882_n1488# 0.0761f
C154 drain_left.n13 a_n1882_n1488# 0.548824f
C155 drain_left.n14 a_n1882_n1488# 0.351471f
C156 drain_left.t6 a_n1882_n1488# 0.0761f
C157 drain_left.t13 a_n1882_n1488# 0.0761f
C158 drain_left.n15 a_n1882_n1488# 0.548824f
C159 drain_left.n16 a_n1882_n1488# 0.61418f
C160 source.t31 a_n1882_n1488# 0.624527f
C161 source.n0 a_n1882_n1488# 0.836533f
C162 source.t25 a_n1882_n1488# 0.07521f
C163 source.t29 a_n1882_n1488# 0.07521f
C164 source.n1 a_n1882_n1488# 0.476872f
C165 source.n2 a_n1882_n1488# 0.369775f
C166 source.t18 a_n1882_n1488# 0.07521f
C167 source.t20 a_n1882_n1488# 0.07521f
C168 source.n3 a_n1882_n1488# 0.476872f
C169 source.n4 a_n1882_n1488# 0.369775f
C170 source.t37 a_n1882_n1488# 0.07521f
C171 source.t26 a_n1882_n1488# 0.07521f
C172 source.n5 a_n1882_n1488# 0.476872f
C173 source.n6 a_n1882_n1488# 0.369775f
C174 source.t24 a_n1882_n1488# 0.07521f
C175 source.t22 a_n1882_n1488# 0.07521f
C176 source.n7 a_n1882_n1488# 0.476872f
C177 source.n8 a_n1882_n1488# 0.369775f
C178 source.t23 a_n1882_n1488# 0.624527f
C179 source.n9 a_n1882_n1488# 0.428559f
C180 source.t0 a_n1882_n1488# 0.624527f
C181 source.n10 a_n1882_n1488# 0.428559f
C182 source.t14 a_n1882_n1488# 0.07521f
C183 source.t13 a_n1882_n1488# 0.07521f
C184 source.n11 a_n1882_n1488# 0.476872f
C185 source.n12 a_n1882_n1488# 0.369775f
C186 source.t17 a_n1882_n1488# 0.07521f
C187 source.t16 a_n1882_n1488# 0.07521f
C188 source.n13 a_n1882_n1488# 0.476872f
C189 source.n14 a_n1882_n1488# 0.369775f
C190 source.t1 a_n1882_n1488# 0.07521f
C191 source.t5 a_n1882_n1488# 0.07521f
C192 source.n15 a_n1882_n1488# 0.476872f
C193 source.n16 a_n1882_n1488# 0.369775f
C194 source.t6 a_n1882_n1488# 0.07521f
C195 source.t9 a_n1882_n1488# 0.07521f
C196 source.n17 a_n1882_n1488# 0.476872f
C197 source.n18 a_n1882_n1488# 0.369775f
C198 source.t15 a_n1882_n1488# 0.624527f
C199 source.n19 a_n1882_n1488# 1.16513f
C200 source.t28 a_n1882_n1488# 0.624524f
C201 source.n20 a_n1882_n1488# 1.16513f
C202 source.t30 a_n1882_n1488# 0.07521f
C203 source.t34 a_n1882_n1488# 0.07521f
C204 source.n21 a_n1882_n1488# 0.476869f
C205 source.n22 a_n1882_n1488# 0.369779f
C206 source.t21 a_n1882_n1488# 0.07521f
C207 source.t27 a_n1882_n1488# 0.07521f
C208 source.n23 a_n1882_n1488# 0.476869f
C209 source.n24 a_n1882_n1488# 0.369779f
C210 source.t32 a_n1882_n1488# 0.07521f
C211 source.t36 a_n1882_n1488# 0.07521f
C212 source.n25 a_n1882_n1488# 0.476869f
C213 source.n26 a_n1882_n1488# 0.369779f
C214 source.t19 a_n1882_n1488# 0.07521f
C215 source.t35 a_n1882_n1488# 0.07521f
C216 source.n27 a_n1882_n1488# 0.476869f
C217 source.n28 a_n1882_n1488# 0.369779f
C218 source.t33 a_n1882_n1488# 0.624524f
C219 source.n29 a_n1882_n1488# 0.428562f
C220 source.t11 a_n1882_n1488# 0.624524f
C221 source.n30 a_n1882_n1488# 0.428562f
C222 source.t3 a_n1882_n1488# 0.07521f
C223 source.t39 a_n1882_n1488# 0.07521f
C224 source.n31 a_n1882_n1488# 0.476869f
C225 source.n32 a_n1882_n1488# 0.369779f
C226 source.t10 a_n1882_n1488# 0.07521f
C227 source.t12 a_n1882_n1488# 0.07521f
C228 source.n33 a_n1882_n1488# 0.476869f
C229 source.n34 a_n1882_n1488# 0.369779f
C230 source.t38 a_n1882_n1488# 0.07521f
C231 source.t8 a_n1882_n1488# 0.07521f
C232 source.n35 a_n1882_n1488# 0.476869f
C233 source.n36 a_n1882_n1488# 0.369779f
C234 source.t2 a_n1882_n1488# 0.07521f
C235 source.t7 a_n1882_n1488# 0.07521f
C236 source.n37 a_n1882_n1488# 0.476869f
C237 source.n38 a_n1882_n1488# 0.369779f
C238 source.t4 a_n1882_n1488# 0.624524f
C239 source.n39 a_n1882_n1488# 0.600584f
C240 source.n40 a_n1882_n1488# 0.915705f
C241 plus.n0 a_n1882_n1488# 0.026881f
C242 plus.t13 a_n1882_n1488# 0.046707f
C243 plus.t18 a_n1882_n1488# 0.046707f
C244 plus.t2 a_n1882_n1488# 0.046707f
C245 plus.n1 a_n1882_n1488# 0.029882f
C246 plus.n2 a_n1882_n1488# 0.026881f
C247 plus.t8 a_n1882_n1488# 0.046707f
C248 plus.t15 a_n1882_n1488# 0.046707f
C249 plus.t16 a_n1882_n1488# 0.046707f
C250 plus.n3 a_n1882_n1488# 0.029882f
C251 plus.n4 a_n1882_n1488# 0.061511f
C252 plus.t19 a_n1882_n1488# 0.046707f
C253 plus.t3 a_n1882_n1488# 0.046707f
C254 plus.t9 a_n1882_n1488# 0.049771f
C255 plus.n5 a_n1882_n1488# 0.037683f
C256 plus.n6 a_n1882_n1488# 0.029882f
C257 plus.n7 a_n1882_n1488# 0.009415f
C258 plus.n8 a_n1882_n1488# 0.029882f
C259 plus.n9 a_n1882_n1488# 0.009415f
C260 plus.n10 a_n1882_n1488# 0.026881f
C261 plus.n11 a_n1882_n1488# 0.026881f
C262 plus.n12 a_n1882_n1488# 0.009415f
C263 plus.n13 a_n1882_n1488# 0.029882f
C264 plus.n14 a_n1882_n1488# 0.009415f
C265 plus.n15 a_n1882_n1488# 0.029882f
C266 plus.n16 a_n1882_n1488# 0.009415f
C267 plus.n17 a_n1882_n1488# 0.026881f
C268 plus.n18 a_n1882_n1488# 0.026881f
C269 plus.n19 a_n1882_n1488# 0.009415f
C270 plus.n20 a_n1882_n1488# 0.029882f
C271 plus.n21 a_n1882_n1488# 0.009415f
C272 plus.n22 a_n1882_n1488# 0.029882f
C273 plus.t6 a_n1882_n1488# 0.049771f
C274 plus.n23 a_n1882_n1488# 0.037642f
C275 plus.n24 a_n1882_n1488# 0.199318f
C276 plus.n25 a_n1882_n1488# 0.026881f
C277 plus.t12 a_n1882_n1488# 0.049771f
C278 plus.t5 a_n1882_n1488# 0.046707f
C279 plus.t17 a_n1882_n1488# 0.046707f
C280 plus.t7 a_n1882_n1488# 0.046707f
C281 plus.n26 a_n1882_n1488# 0.029882f
C282 plus.n27 a_n1882_n1488# 0.026881f
C283 plus.t1 a_n1882_n1488# 0.046707f
C284 plus.t14 a_n1882_n1488# 0.046707f
C285 plus.t10 a_n1882_n1488# 0.046707f
C286 plus.n28 a_n1882_n1488# 0.029882f
C287 plus.n29 a_n1882_n1488# 0.061511f
C288 plus.t0 a_n1882_n1488# 0.046707f
C289 plus.t11 a_n1882_n1488# 0.046707f
C290 plus.t4 a_n1882_n1488# 0.049771f
C291 plus.n30 a_n1882_n1488# 0.037683f
C292 plus.n31 a_n1882_n1488# 0.029882f
C293 plus.n32 a_n1882_n1488# 0.009415f
C294 plus.n33 a_n1882_n1488# 0.029882f
C295 plus.n34 a_n1882_n1488# 0.009415f
C296 plus.n35 a_n1882_n1488# 0.026881f
C297 plus.n36 a_n1882_n1488# 0.026881f
C298 plus.n37 a_n1882_n1488# 0.009415f
C299 plus.n38 a_n1882_n1488# 0.029882f
C300 plus.n39 a_n1882_n1488# 0.009415f
C301 plus.n40 a_n1882_n1488# 0.029882f
C302 plus.n41 a_n1882_n1488# 0.009415f
C303 plus.n42 a_n1882_n1488# 0.026881f
C304 plus.n43 a_n1882_n1488# 0.026881f
C305 plus.n44 a_n1882_n1488# 0.009415f
C306 plus.n45 a_n1882_n1488# 0.029882f
C307 plus.n46 a_n1882_n1488# 0.009415f
C308 plus.n47 a_n1882_n1488# 0.029882f
C309 plus.n48 a_n1882_n1488# 0.037642f
C310 plus.n49 a_n1882_n1488# 0.634978f
.ends

