* NGSPICE file created from diffpair349.ext - technology: sky130A

.subckt diffpair349 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t34 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 drain_left.t22 plus.t1 source.t31 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 drain_right.t23 minus.t0 source.t0 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_right.t22 minus.t1 source.t1 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 drain_left.t21 plus.t2 source.t43 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 drain_left.t20 plus.t3 source.t27 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X6 drain_left.t19 plus.t4 source.t46 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 source.t5 minus.t2 drain_right.t21 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 source.t9 minus.t3 drain_right.t20 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X9 drain_left.t18 plus.t5 source.t29 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X10 source.t13 minus.t4 drain_right.t19 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X11 drain_right.t18 minus.t5 source.t6 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X12 source.t39 plus.t6 drain_left.t17 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X13 drain_left.t16 plus.t7 source.t41 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X14 source.t36 plus.t8 drain_left.t15 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X15 source.t35 plus.t9 drain_left.t14 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X16 source.t15 minus.t6 drain_right.t17 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 source.t7 minus.t7 drain_right.t16 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X18 a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X19 source.t20 minus.t8 drain_right.t15 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X20 a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X21 source.t23 minus.t9 drain_right.t14 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X22 drain_left.t13 plus.t10 source.t32 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X23 source.t44 plus.t11 drain_left.t12 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X24 source.t37 plus.t12 drain_left.t11 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X25 source.t28 plus.t13 drain_left.t10 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X26 source.t47 plus.t14 drain_left.t9 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X27 drain_right.t13 minus.t10 source.t14 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X28 drain_right.t12 minus.t11 source.t2 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X29 drain_left.t8 plus.t15 source.t30 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X30 drain_right.t11 minus.t12 source.t4 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X31 source.t40 plus.t16 drain_left.t7 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X32 drain_left.t6 plus.t17 source.t42 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X33 source.t38 plus.t18 drain_left.t5 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X34 drain_right.t10 minus.t13 source.t10 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X35 source.t17 minus.t14 drain_right.t9 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X36 source.t22 minus.t15 drain_right.t8 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X37 source.t33 plus.t19 drain_left.t4 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X38 drain_right.t7 minus.t16 source.t3 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X39 source.t8 minus.t17 drain_right.t6 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X40 source.t11 minus.t18 drain_right.t5 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X41 a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X42 source.t45 plus.t20 drain_left.t3 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X43 drain_left.t2 plus.t21 source.t24 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X44 drain_right.t4 minus.t19 source.t16 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X45 source.t21 minus.t20 drain_right.t3 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X46 source.t26 plus.t22 drain_left.t1 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X47 a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X48 drain_right.t2 minus.t21 source.t12 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X49 drain_right.t1 minus.t22 source.t19 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X50 drain_right.t0 minus.t23 source.t18 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X51 drain_left.t0 plus.t23 source.t25 a_n2224_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
R0 plus.n6 plus.t8 1020.67
R1 plus.n33 plus.t3 1020.67
R2 plus.n42 plus.t21 1020.67
R3 plus.n68 plus.t9 1020.67
R4 plus.n7 plus.t1 992.92
R5 plus.n8 plus.t14 992.92
R6 plus.n14 plus.t0 992.92
R7 plus.n16 plus.t13 992.92
R8 plus.n3 plus.t23 992.92
R9 plus.n21 plus.t12 992.92
R10 plus.n23 plus.t5 992.92
R11 plus.n24 plus.t19 992.92
R12 plus.n30 plus.t4 992.92
R13 plus.n32 plus.t18 992.92
R14 plus.n44 plus.t16 992.92
R15 plus.n43 plus.t7 992.92
R16 plus.n50 plus.t22 992.92
R17 plus.n52 plus.t2 992.92
R18 plus.n39 plus.t20 992.92
R19 plus.n57 plus.t15 992.92
R20 plus.n59 plus.t6 992.92
R21 plus.n38 plus.t17 992.92
R22 plus.n65 plus.t11 992.92
R23 plus.n67 plus.t10 992.92
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus.n17 plus.n3 30.6732
R75 plus.n22 plus.n21 30.6732
R76 plus.n58 plus.n57 30.6732
R77 plus.n53 plus.n39 30.6732
R78 plus plus.n69 30.2225
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 10.9399
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n11 source.t36 51.0588
R119 source.n12 source.t3 51.0588
R120 source.n23 source.t11 51.0588
R121 source.n47 source.t2 51.0586
R122 source.n36 source.t21 51.0586
R123 source.n35 source.t24 51.0586
R124 source.n24 source.t35 51.0586
R125 source.n0 source.t27 51.0586
R126 source.n2 source.n1 48.8588
R127 source.n4 source.n3 48.8588
R128 source.n6 source.n5 48.8588
R129 source.n8 source.n7 48.8588
R130 source.n10 source.n9 48.8588
R131 source.n14 source.n13 48.8588
R132 source.n16 source.n15 48.8588
R133 source.n18 source.n17 48.8588
R134 source.n20 source.n19 48.8588
R135 source.n22 source.n21 48.8588
R136 source.n46 source.n45 48.8586
R137 source.n44 source.n43 48.8586
R138 source.n42 source.n41 48.8586
R139 source.n40 source.n39 48.8586
R140 source.n38 source.n37 48.8586
R141 source.n34 source.n33 48.8586
R142 source.n32 source.n31 48.8586
R143 source.n30 source.n29 48.8586
R144 source.n28 source.n27 48.8586
R145 source.n26 source.n25 48.8586
R146 source.n24 source.n23 19.515
R147 source.n48 source.n0 14.0021
R148 source.n48 source.n47 5.51343
R149 source.n45 source.t0 2.2005
R150 source.n45 source.t8 2.2005
R151 source.n43 source.t4 2.2005
R152 source.n43 source.t23 2.2005
R153 source.n41 source.t16 2.2005
R154 source.n41 source.t17 2.2005
R155 source.n39 source.t14 2.2005
R156 source.n39 source.t9 2.2005
R157 source.n37 source.t1 2.2005
R158 source.n37 source.t22 2.2005
R159 source.n33 source.t41 2.2005
R160 source.n33 source.t40 2.2005
R161 source.n31 source.t43 2.2005
R162 source.n31 source.t26 2.2005
R163 source.n29 source.t30 2.2005
R164 source.n29 source.t45 2.2005
R165 source.n27 source.t42 2.2005
R166 source.n27 source.t39 2.2005
R167 source.n25 source.t32 2.2005
R168 source.n25 source.t44 2.2005
R169 source.n1 source.t46 2.2005
R170 source.n1 source.t38 2.2005
R171 source.n3 source.t29 2.2005
R172 source.n3 source.t33 2.2005
R173 source.n5 source.t25 2.2005
R174 source.n5 source.t37 2.2005
R175 source.n7 source.t34 2.2005
R176 source.n7 source.t28 2.2005
R177 source.n9 source.t31 2.2005
R178 source.n9 source.t47 2.2005
R179 source.n13 source.t10 2.2005
R180 source.n13 source.t13 2.2005
R181 source.n15 source.t12 2.2005
R182 source.n15 source.t5 2.2005
R183 source.n17 source.t19 2.2005
R184 source.n17 source.t7 2.2005
R185 source.n19 source.t18 2.2005
R186 source.n19 source.t15 2.2005
R187 source.n21 source.t6 2.2005
R188 source.n21 source.t20 2.2005
R189 source.n23 source.n22 0.5005
R190 source.n22 source.n20 0.5005
R191 source.n20 source.n18 0.5005
R192 source.n18 source.n16 0.5005
R193 source.n16 source.n14 0.5005
R194 source.n14 source.n12 0.5005
R195 source.n11 source.n10 0.5005
R196 source.n10 source.n8 0.5005
R197 source.n8 source.n6 0.5005
R198 source.n6 source.n4 0.5005
R199 source.n4 source.n2 0.5005
R200 source.n2 source.n0 0.5005
R201 source.n26 source.n24 0.5005
R202 source.n28 source.n26 0.5005
R203 source.n30 source.n28 0.5005
R204 source.n32 source.n30 0.5005
R205 source.n34 source.n32 0.5005
R206 source.n35 source.n34 0.5005
R207 source.n38 source.n36 0.5005
R208 source.n40 source.n38 0.5005
R209 source.n42 source.n40 0.5005
R210 source.n44 source.n42 0.5005
R211 source.n46 source.n44 0.5005
R212 source.n47 source.n46 0.5005
R213 source.n12 source.n11 0.470328
R214 source.n36 source.n35 0.470328
R215 source source.n48 0.188
R216 drain_left.n13 drain_left.n11 66.0376
R217 drain_left.n7 drain_left.n5 66.0373
R218 drain_left.n2 drain_left.n0 66.0373
R219 drain_left.n19 drain_left.n18 65.5376
R220 drain_left.n17 drain_left.n16 65.5376
R221 drain_left.n15 drain_left.n14 65.5376
R222 drain_left.n13 drain_left.n12 65.5376
R223 drain_left.n21 drain_left.n20 65.5374
R224 drain_left.n7 drain_left.n6 65.5373
R225 drain_left.n9 drain_left.n8 65.5373
R226 drain_left.n4 drain_left.n3 65.5373
R227 drain_left.n2 drain_left.n1 65.5373
R228 drain_left drain_left.n10 29.8443
R229 drain_left drain_left.n21 6.15322
R230 drain_left.n5 drain_left.t7 2.2005
R231 drain_left.n5 drain_left.t2 2.2005
R232 drain_left.n6 drain_left.t1 2.2005
R233 drain_left.n6 drain_left.t16 2.2005
R234 drain_left.n8 drain_left.t3 2.2005
R235 drain_left.n8 drain_left.t21 2.2005
R236 drain_left.n3 drain_left.t17 2.2005
R237 drain_left.n3 drain_left.t8 2.2005
R238 drain_left.n1 drain_left.t12 2.2005
R239 drain_left.n1 drain_left.t6 2.2005
R240 drain_left.n0 drain_left.t14 2.2005
R241 drain_left.n0 drain_left.t13 2.2005
R242 drain_left.n20 drain_left.t5 2.2005
R243 drain_left.n20 drain_left.t20 2.2005
R244 drain_left.n18 drain_left.t4 2.2005
R245 drain_left.n18 drain_left.t19 2.2005
R246 drain_left.n16 drain_left.t11 2.2005
R247 drain_left.n16 drain_left.t18 2.2005
R248 drain_left.n14 drain_left.t10 2.2005
R249 drain_left.n14 drain_left.t0 2.2005
R250 drain_left.n12 drain_left.t9 2.2005
R251 drain_left.n12 drain_left.t23 2.2005
R252 drain_left.n11 drain_left.t15 2.2005
R253 drain_left.n11 drain_left.t22 2.2005
R254 drain_left.n9 drain_left.n7 0.5005
R255 drain_left.n4 drain_left.n2 0.5005
R256 drain_left.n15 drain_left.n13 0.5005
R257 drain_left.n17 drain_left.n15 0.5005
R258 drain_left.n19 drain_left.n17 0.5005
R259 drain_left.n21 drain_left.n19 0.5005
R260 drain_left.n10 drain_left.n9 0.195154
R261 drain_left.n10 drain_left.n4 0.195154
R262 minus.n33 minus.t18 1020.67
R263 minus.n7 minus.t16 1020.67
R264 minus.n68 minus.t11 1020.67
R265 minus.n41 minus.t20 1020.67
R266 minus.n32 minus.t5 992.92
R267 minus.n30 minus.t8 992.92
R268 minus.n3 minus.t23 992.92
R269 minus.n24 minus.t6 992.92
R270 minus.n22 minus.t22 992.92
R271 minus.n4 minus.t7 992.92
R272 minus.n17 minus.t21 992.92
R273 minus.n15 minus.t2 992.92
R274 minus.n8 minus.t13 992.92
R275 minus.n9 minus.t4 992.92
R276 minus.n67 minus.t17 992.92
R277 minus.n65 minus.t0 992.92
R278 minus.n59 minus.t9 992.92
R279 minus.n58 minus.t12 992.92
R280 minus.n56 minus.t14 992.92
R281 minus.n38 minus.t19 992.92
R282 minus.n51 minus.t3 992.92
R283 minus.n49 minus.t10 992.92
R284 minus.n43 minus.t15 992.92
R285 minus.n42 minus.t1 992.92
R286 minus.n11 minus.n7 161.489
R287 minus.n45 minus.n41 161.489
R288 minus.n34 minus.n33 161.3
R289 minus.n31 minus.n0 161.3
R290 minus.n29 minus.n28 161.3
R291 minus.n27 minus.n1 161.3
R292 minus.n26 minus.n25 161.3
R293 minus.n23 minus.n2 161.3
R294 minus.n21 minus.n20 161.3
R295 minus.n19 minus.n18 161.3
R296 minus.n16 minus.n5 161.3
R297 minus.n14 minus.n13 161.3
R298 minus.n12 minus.n6 161.3
R299 minus.n11 minus.n10 161.3
R300 minus.n69 minus.n68 161.3
R301 minus.n66 minus.n35 161.3
R302 minus.n64 minus.n63 161.3
R303 minus.n62 minus.n36 161.3
R304 minus.n61 minus.n60 161.3
R305 minus.n57 minus.n37 161.3
R306 minus.n55 minus.n54 161.3
R307 minus.n53 minus.n52 161.3
R308 minus.n50 minus.n39 161.3
R309 minus.n48 minus.n47 161.3
R310 minus.n46 minus.n40 161.3
R311 minus.n45 minus.n44 161.3
R312 minus.n29 minus.n1 73.0308
R313 minus.n14 minus.n6 73.0308
R314 minus.n48 minus.n40 73.0308
R315 minus.n64 minus.n36 73.0308
R316 minus.n31 minus.n30 68.649
R317 minus.n10 minus.n8 68.649
R318 minus.n44 minus.n43 68.649
R319 minus.n66 minus.n65 68.649
R320 minus.n25 minus.n3 65.7278
R321 minus.n16 minus.n15 65.7278
R322 minus.n50 minus.n49 65.7278
R323 minus.n60 minus.n59 65.7278
R324 minus.n33 minus.n32 56.9641
R325 minus.n9 minus.n7 56.9641
R326 minus.n42 minus.n41 56.9641
R327 minus.n68 minus.n67 56.9641
R328 minus.n24 minus.n23 54.0429
R329 minus.n18 minus.n17 54.0429
R330 minus.n52 minus.n51 54.0429
R331 minus.n58 minus.n57 54.0429
R332 minus.n22 minus.n21 42.3581
R333 minus.n21 minus.n4 42.3581
R334 minus.n55 minus.n38 42.3581
R335 minus.n56 minus.n55 42.3581
R336 minus.n70 minus.n34 35.205
R337 minus.n23 minus.n22 30.6732
R338 minus.n18 minus.n4 30.6732
R339 minus.n52 minus.n38 30.6732
R340 minus.n57 minus.n56 30.6732
R341 minus.n25 minus.n24 18.9884
R342 minus.n17 minus.n16 18.9884
R343 minus.n51 minus.n50 18.9884
R344 minus.n60 minus.n58 18.9884
R345 minus.n32 minus.n31 16.0672
R346 minus.n10 minus.n9 16.0672
R347 minus.n44 minus.n42 16.0672
R348 minus.n67 minus.n66 16.0672
R349 minus.n3 minus.n1 7.30353
R350 minus.n15 minus.n14 7.30353
R351 minus.n49 minus.n48 7.30353
R352 minus.n59 minus.n36 7.30353
R353 minus.n70 minus.n69 6.43232
R354 minus.n30 minus.n29 4.38232
R355 minus.n8 minus.n6 4.38232
R356 minus.n43 minus.n40 4.38232
R357 minus.n65 minus.n64 4.38232
R358 minus.n34 minus.n0 0.189894
R359 minus.n28 minus.n0 0.189894
R360 minus.n28 minus.n27 0.189894
R361 minus.n27 minus.n26 0.189894
R362 minus.n26 minus.n2 0.189894
R363 minus.n20 minus.n2 0.189894
R364 minus.n20 minus.n19 0.189894
R365 minus.n19 minus.n5 0.189894
R366 minus.n13 minus.n5 0.189894
R367 minus.n13 minus.n12 0.189894
R368 minus.n12 minus.n11 0.189894
R369 minus.n46 minus.n45 0.189894
R370 minus.n47 minus.n46 0.189894
R371 minus.n47 minus.n39 0.189894
R372 minus.n53 minus.n39 0.189894
R373 minus.n54 minus.n53 0.189894
R374 minus.n54 minus.n37 0.189894
R375 minus.n61 minus.n37 0.189894
R376 minus.n62 minus.n61 0.189894
R377 minus.n63 minus.n62 0.189894
R378 minus.n63 minus.n35 0.189894
R379 minus.n69 minus.n35 0.189894
R380 minus minus.n70 0.188
R381 drain_right.n13 drain_right.n11 66.0374
R382 drain_right.n7 drain_right.n5 66.0373
R383 drain_right.n2 drain_right.n0 66.0373
R384 drain_right.n13 drain_right.n12 65.5376
R385 drain_right.n15 drain_right.n14 65.5376
R386 drain_right.n17 drain_right.n16 65.5376
R387 drain_right.n19 drain_right.n18 65.5376
R388 drain_right.n21 drain_right.n20 65.5376
R389 drain_right.n7 drain_right.n6 65.5373
R390 drain_right.n9 drain_right.n8 65.5373
R391 drain_right.n4 drain_right.n3 65.5373
R392 drain_right.n2 drain_right.n1 65.5373
R393 drain_right drain_right.n10 29.2911
R394 drain_right drain_right.n21 6.15322
R395 drain_right.n5 drain_right.t6 2.2005
R396 drain_right.n5 drain_right.t12 2.2005
R397 drain_right.n6 drain_right.t14 2.2005
R398 drain_right.n6 drain_right.t23 2.2005
R399 drain_right.n8 drain_right.t9 2.2005
R400 drain_right.n8 drain_right.t11 2.2005
R401 drain_right.n3 drain_right.t20 2.2005
R402 drain_right.n3 drain_right.t4 2.2005
R403 drain_right.n1 drain_right.t8 2.2005
R404 drain_right.n1 drain_right.t13 2.2005
R405 drain_right.n0 drain_right.t3 2.2005
R406 drain_right.n0 drain_right.t22 2.2005
R407 drain_right.n11 drain_right.t19 2.2005
R408 drain_right.n11 drain_right.t7 2.2005
R409 drain_right.n12 drain_right.t21 2.2005
R410 drain_right.n12 drain_right.t10 2.2005
R411 drain_right.n14 drain_right.t16 2.2005
R412 drain_right.n14 drain_right.t2 2.2005
R413 drain_right.n16 drain_right.t17 2.2005
R414 drain_right.n16 drain_right.t1 2.2005
R415 drain_right.n18 drain_right.t15 2.2005
R416 drain_right.n18 drain_right.t0 2.2005
R417 drain_right.n20 drain_right.t5 2.2005
R418 drain_right.n20 drain_right.t18 2.2005
R419 drain_right.n9 drain_right.n7 0.5005
R420 drain_right.n4 drain_right.n2 0.5005
R421 drain_right.n21 drain_right.n19 0.5005
R422 drain_right.n19 drain_right.n17 0.5005
R423 drain_right.n17 drain_right.n15 0.5005
R424 drain_right.n15 drain_right.n13 0.5005
R425 drain_right.n10 drain_right.n9 0.195154
R426 drain_right.n10 drain_right.n4 0.195154
C0 minus plus 5.37859f
C1 drain_right drain_left 1.19771f
C2 source minus 5.55004f
C3 drain_right plus 0.374075f
C4 drain_right source 37.3453f
C5 drain_left plus 5.89868f
C6 drain_left source 37.3449f
C7 drain_right minus 5.68001f
C8 source plus 5.56408f
C9 drain_left minus 0.172313f
C10 drain_right a_n2224_n2688# 6.7013f
C11 drain_left a_n2224_n2688# 7.0406f
C12 source a_n2224_n2688# 7.236802f
C13 minus a_n2224_n2688# 8.519746f
C14 plus a_n2224_n2688# 10.40405f
C15 drain_right.t3 a_n2224_n2688# 0.256541f
C16 drain_right.t22 a_n2224_n2688# 0.256541f
C17 drain_right.n0 a_n2224_n2688# 2.24706f
C18 drain_right.t8 a_n2224_n2688# 0.256541f
C19 drain_right.t13 a_n2224_n2688# 0.256541f
C20 drain_right.n1 a_n2224_n2688# 2.24388f
C21 drain_right.n2 a_n2224_n2688# 0.82168f
C22 drain_right.t20 a_n2224_n2688# 0.256541f
C23 drain_right.t4 a_n2224_n2688# 0.256541f
C24 drain_right.n3 a_n2224_n2688# 2.24388f
C25 drain_right.n4 a_n2224_n2688# 0.37397f
C26 drain_right.t6 a_n2224_n2688# 0.256541f
C27 drain_right.t12 a_n2224_n2688# 0.256541f
C28 drain_right.n5 a_n2224_n2688# 2.24706f
C29 drain_right.t14 a_n2224_n2688# 0.256541f
C30 drain_right.t23 a_n2224_n2688# 0.256541f
C31 drain_right.n6 a_n2224_n2688# 2.24388f
C32 drain_right.n7 a_n2224_n2688# 0.82168f
C33 drain_right.t9 a_n2224_n2688# 0.256541f
C34 drain_right.t11 a_n2224_n2688# 0.256541f
C35 drain_right.n8 a_n2224_n2688# 2.24388f
C36 drain_right.n9 a_n2224_n2688# 0.37397f
C37 drain_right.n10 a_n2224_n2688# 1.58538f
C38 drain_right.t19 a_n2224_n2688# 0.256541f
C39 drain_right.t7 a_n2224_n2688# 0.256541f
C40 drain_right.n11 a_n2224_n2688# 2.24705f
C41 drain_right.t21 a_n2224_n2688# 0.256541f
C42 drain_right.t10 a_n2224_n2688# 0.256541f
C43 drain_right.n12 a_n2224_n2688# 2.24388f
C44 drain_right.n13 a_n2224_n2688# 0.82168f
C45 drain_right.t16 a_n2224_n2688# 0.256541f
C46 drain_right.t2 a_n2224_n2688# 0.256541f
C47 drain_right.n14 a_n2224_n2688# 2.24388f
C48 drain_right.n15 a_n2224_n2688# 0.40516f
C49 drain_right.t17 a_n2224_n2688# 0.256541f
C50 drain_right.t1 a_n2224_n2688# 0.256541f
C51 drain_right.n16 a_n2224_n2688# 2.24388f
C52 drain_right.n17 a_n2224_n2688# 0.40516f
C53 drain_right.t15 a_n2224_n2688# 0.256541f
C54 drain_right.t0 a_n2224_n2688# 0.256541f
C55 drain_right.n18 a_n2224_n2688# 2.24388f
C56 drain_right.n19 a_n2224_n2688# 0.40516f
C57 drain_right.t5 a_n2224_n2688# 0.256541f
C58 drain_right.t18 a_n2224_n2688# 0.256541f
C59 drain_right.n20 a_n2224_n2688# 2.24388f
C60 drain_right.n21 a_n2224_n2688# 0.702904f
C61 minus.n0 a_n2224_n2688# 0.050016f
C62 minus.t18 a_n2224_n2688# 0.322524f
C63 minus.t5 a_n2224_n2688# 0.318883f
C64 minus.t8 a_n2224_n2688# 0.318883f
C65 minus.n1 a_n2224_n2688# 0.018134f
C66 minus.n2 a_n2224_n2688# 0.050016f
C67 minus.t23 a_n2224_n2688# 0.318883f
C68 minus.n3 a_n2224_n2688# 0.13573f
C69 minus.t6 a_n2224_n2688# 0.318883f
C70 minus.t22 a_n2224_n2688# 0.318883f
C71 minus.t7 a_n2224_n2688# 0.318883f
C72 minus.n4 a_n2224_n2688# 0.13573f
C73 minus.n5 a_n2224_n2688# 0.050016f
C74 minus.t21 a_n2224_n2688# 0.318883f
C75 minus.t2 a_n2224_n2688# 0.318883f
C76 minus.n6 a_n2224_n2688# 0.017517f
C77 minus.t16 a_n2224_n2688# 0.322524f
C78 minus.n7 a_n2224_n2688# 0.149362f
C79 minus.t13 a_n2224_n2688# 0.318883f
C80 minus.n8 a_n2224_n2688# 0.13573f
C81 minus.t4 a_n2224_n2688# 0.318883f
C82 minus.n9 a_n2224_n2688# 0.13573f
C83 minus.n10 a_n2224_n2688# 0.019059f
C84 minus.n11 a_n2224_n2688# 0.103978f
C85 minus.n12 a_n2224_n2688# 0.050016f
C86 minus.n13 a_n2224_n2688# 0.050016f
C87 minus.n14 a_n2224_n2688# 0.018134f
C88 minus.n15 a_n2224_n2688# 0.13573f
C89 minus.n16 a_n2224_n2688# 0.019059f
C90 minus.n17 a_n2224_n2688# 0.13573f
C91 minus.n18 a_n2224_n2688# 0.019059f
C92 minus.n19 a_n2224_n2688# 0.050016f
C93 minus.n20 a_n2224_n2688# 0.050016f
C94 minus.n21 a_n2224_n2688# 0.019059f
C95 minus.n22 a_n2224_n2688# 0.13573f
C96 minus.n23 a_n2224_n2688# 0.019059f
C97 minus.n24 a_n2224_n2688# 0.13573f
C98 minus.n25 a_n2224_n2688# 0.019059f
C99 minus.n26 a_n2224_n2688# 0.050016f
C100 minus.n27 a_n2224_n2688# 0.050016f
C101 minus.n28 a_n2224_n2688# 0.050016f
C102 minus.n29 a_n2224_n2688# 0.017517f
C103 minus.n30 a_n2224_n2688# 0.13573f
C104 minus.n31 a_n2224_n2688# 0.019059f
C105 minus.n32 a_n2224_n2688# 0.13573f
C106 minus.n33 a_n2224_n2688# 0.149299f
C107 minus.n34 a_n2224_n2688# 1.68958f
C108 minus.n35 a_n2224_n2688# 0.050016f
C109 minus.t17 a_n2224_n2688# 0.318883f
C110 minus.t0 a_n2224_n2688# 0.318883f
C111 minus.n36 a_n2224_n2688# 0.018134f
C112 minus.n37 a_n2224_n2688# 0.050016f
C113 minus.t12 a_n2224_n2688# 0.318883f
C114 minus.t14 a_n2224_n2688# 0.318883f
C115 minus.t19 a_n2224_n2688# 0.318883f
C116 minus.n38 a_n2224_n2688# 0.13573f
C117 minus.n39 a_n2224_n2688# 0.050016f
C118 minus.t3 a_n2224_n2688# 0.318883f
C119 minus.t10 a_n2224_n2688# 0.318883f
C120 minus.n40 a_n2224_n2688# 0.017517f
C121 minus.t20 a_n2224_n2688# 0.322524f
C122 minus.n41 a_n2224_n2688# 0.149362f
C123 minus.t1 a_n2224_n2688# 0.318883f
C124 minus.n42 a_n2224_n2688# 0.13573f
C125 minus.t15 a_n2224_n2688# 0.318883f
C126 minus.n43 a_n2224_n2688# 0.13573f
C127 minus.n44 a_n2224_n2688# 0.019059f
C128 minus.n45 a_n2224_n2688# 0.103978f
C129 minus.n46 a_n2224_n2688# 0.050016f
C130 minus.n47 a_n2224_n2688# 0.050016f
C131 minus.n48 a_n2224_n2688# 0.018134f
C132 minus.n49 a_n2224_n2688# 0.13573f
C133 minus.n50 a_n2224_n2688# 0.019059f
C134 minus.n51 a_n2224_n2688# 0.13573f
C135 minus.n52 a_n2224_n2688# 0.019059f
C136 minus.n53 a_n2224_n2688# 0.050016f
C137 minus.n54 a_n2224_n2688# 0.050016f
C138 minus.n55 a_n2224_n2688# 0.019059f
C139 minus.n56 a_n2224_n2688# 0.13573f
C140 minus.n57 a_n2224_n2688# 0.019059f
C141 minus.n58 a_n2224_n2688# 0.13573f
C142 minus.t9 a_n2224_n2688# 0.318883f
C143 minus.n59 a_n2224_n2688# 0.13573f
C144 minus.n60 a_n2224_n2688# 0.019059f
C145 minus.n61 a_n2224_n2688# 0.050016f
C146 minus.n62 a_n2224_n2688# 0.050016f
C147 minus.n63 a_n2224_n2688# 0.050016f
C148 minus.n64 a_n2224_n2688# 0.017517f
C149 minus.n65 a_n2224_n2688# 0.13573f
C150 minus.n66 a_n2224_n2688# 0.019059f
C151 minus.n67 a_n2224_n2688# 0.13573f
C152 minus.t11 a_n2224_n2688# 0.322524f
C153 minus.n68 a_n2224_n2688# 0.149299f
C154 minus.n69 a_n2224_n2688# 0.318991f
C155 minus.n70 a_n2224_n2688# 2.06119f
C156 drain_left.t14 a_n2224_n2688# 0.256892f
C157 drain_left.t13 a_n2224_n2688# 0.256892f
C158 drain_left.n0 a_n2224_n2688# 2.25013f
C159 drain_left.t12 a_n2224_n2688# 0.256892f
C160 drain_left.t6 a_n2224_n2688# 0.256892f
C161 drain_left.n1 a_n2224_n2688# 2.24694f
C162 drain_left.n2 a_n2224_n2688# 0.822802f
C163 drain_left.t17 a_n2224_n2688# 0.256892f
C164 drain_left.t8 a_n2224_n2688# 0.256892f
C165 drain_left.n3 a_n2224_n2688# 2.24694f
C166 drain_left.n4 a_n2224_n2688# 0.374481f
C167 drain_left.t7 a_n2224_n2688# 0.256892f
C168 drain_left.t2 a_n2224_n2688# 0.256892f
C169 drain_left.n5 a_n2224_n2688# 2.25013f
C170 drain_left.t1 a_n2224_n2688# 0.256892f
C171 drain_left.t16 a_n2224_n2688# 0.256892f
C172 drain_left.n6 a_n2224_n2688# 2.24694f
C173 drain_left.n7 a_n2224_n2688# 0.822802f
C174 drain_left.t3 a_n2224_n2688# 0.256892f
C175 drain_left.t21 a_n2224_n2688# 0.256892f
C176 drain_left.n8 a_n2224_n2688# 2.24694f
C177 drain_left.n9 a_n2224_n2688# 0.374481f
C178 drain_left.n10 a_n2224_n2688# 1.66139f
C179 drain_left.t15 a_n2224_n2688# 0.256892f
C180 drain_left.t22 a_n2224_n2688# 0.256892f
C181 drain_left.n11 a_n2224_n2688# 2.25013f
C182 drain_left.t9 a_n2224_n2688# 0.256892f
C183 drain_left.t23 a_n2224_n2688# 0.256892f
C184 drain_left.n12 a_n2224_n2688# 2.24695f
C185 drain_left.n13 a_n2224_n2688# 0.822793f
C186 drain_left.t10 a_n2224_n2688# 0.256892f
C187 drain_left.t0 a_n2224_n2688# 0.256892f
C188 drain_left.n14 a_n2224_n2688# 2.24695f
C189 drain_left.n15 a_n2224_n2688# 0.405713f
C190 drain_left.t11 a_n2224_n2688# 0.256892f
C191 drain_left.t18 a_n2224_n2688# 0.256892f
C192 drain_left.n16 a_n2224_n2688# 2.24695f
C193 drain_left.n17 a_n2224_n2688# 0.405713f
C194 drain_left.t4 a_n2224_n2688# 0.256892f
C195 drain_left.t19 a_n2224_n2688# 0.256892f
C196 drain_left.n18 a_n2224_n2688# 2.24695f
C197 drain_left.n19 a_n2224_n2688# 0.405713f
C198 drain_left.t5 a_n2224_n2688# 0.256892f
C199 drain_left.t20 a_n2224_n2688# 0.256892f
C200 drain_left.n20 a_n2224_n2688# 2.24694f
C201 drain_left.n21 a_n2224_n2688# 0.703873f
C202 source.t27 a_n2224_n2688# 2.47528f
C203 source.n0 a_n2224_n2688# 1.41576f
C204 source.t46 a_n2224_n2688# 0.232127f
C205 source.t38 a_n2224_n2688# 0.232127f
C206 source.n1 a_n2224_n2688# 1.94322f
C207 source.n2 a_n2224_n2688# 0.409364f
C208 source.t29 a_n2224_n2688# 0.232127f
C209 source.t33 a_n2224_n2688# 0.232127f
C210 source.n3 a_n2224_n2688# 1.94322f
C211 source.n4 a_n2224_n2688# 0.409364f
C212 source.t25 a_n2224_n2688# 0.232127f
C213 source.t37 a_n2224_n2688# 0.232127f
C214 source.n5 a_n2224_n2688# 1.94322f
C215 source.n6 a_n2224_n2688# 0.409364f
C216 source.t34 a_n2224_n2688# 0.232127f
C217 source.t28 a_n2224_n2688# 0.232127f
C218 source.n7 a_n2224_n2688# 1.94322f
C219 source.n8 a_n2224_n2688# 0.409364f
C220 source.t31 a_n2224_n2688# 0.232127f
C221 source.t47 a_n2224_n2688# 0.232127f
C222 source.n9 a_n2224_n2688# 1.94322f
C223 source.n10 a_n2224_n2688# 0.409364f
C224 source.t36 a_n2224_n2688# 2.47528f
C225 source.n11 a_n2224_n2688# 0.507197f
C226 source.t3 a_n2224_n2688# 2.47528f
C227 source.n12 a_n2224_n2688# 0.507197f
C228 source.t10 a_n2224_n2688# 0.232127f
C229 source.t13 a_n2224_n2688# 0.232127f
C230 source.n13 a_n2224_n2688# 1.94322f
C231 source.n14 a_n2224_n2688# 0.409364f
C232 source.t12 a_n2224_n2688# 0.232127f
C233 source.t5 a_n2224_n2688# 0.232127f
C234 source.n15 a_n2224_n2688# 1.94322f
C235 source.n16 a_n2224_n2688# 0.409364f
C236 source.t19 a_n2224_n2688# 0.232127f
C237 source.t7 a_n2224_n2688# 0.232127f
C238 source.n17 a_n2224_n2688# 1.94322f
C239 source.n18 a_n2224_n2688# 0.409364f
C240 source.t18 a_n2224_n2688# 0.232127f
C241 source.t15 a_n2224_n2688# 0.232127f
C242 source.n19 a_n2224_n2688# 1.94322f
C243 source.n20 a_n2224_n2688# 0.409364f
C244 source.t6 a_n2224_n2688# 0.232127f
C245 source.t20 a_n2224_n2688# 0.232127f
C246 source.n21 a_n2224_n2688# 1.94322f
C247 source.n22 a_n2224_n2688# 0.409364f
C248 source.t11 a_n2224_n2688# 2.47528f
C249 source.n23 a_n2224_n2688# 1.88852f
C250 source.t35 a_n2224_n2688# 2.47528f
C251 source.n24 a_n2224_n2688# 1.88852f
C252 source.t32 a_n2224_n2688# 0.232127f
C253 source.t44 a_n2224_n2688# 0.232127f
C254 source.n25 a_n2224_n2688# 1.94321f
C255 source.n26 a_n2224_n2688# 0.40937f
C256 source.t42 a_n2224_n2688# 0.232127f
C257 source.t39 a_n2224_n2688# 0.232127f
C258 source.n27 a_n2224_n2688# 1.94321f
C259 source.n28 a_n2224_n2688# 0.40937f
C260 source.t30 a_n2224_n2688# 0.232127f
C261 source.t45 a_n2224_n2688# 0.232127f
C262 source.n29 a_n2224_n2688# 1.94321f
C263 source.n30 a_n2224_n2688# 0.40937f
C264 source.t43 a_n2224_n2688# 0.232127f
C265 source.t26 a_n2224_n2688# 0.232127f
C266 source.n31 a_n2224_n2688# 1.94321f
C267 source.n32 a_n2224_n2688# 0.40937f
C268 source.t41 a_n2224_n2688# 0.232127f
C269 source.t40 a_n2224_n2688# 0.232127f
C270 source.n33 a_n2224_n2688# 1.94321f
C271 source.n34 a_n2224_n2688# 0.40937f
C272 source.t24 a_n2224_n2688# 2.47528f
C273 source.n35 a_n2224_n2688# 0.507203f
C274 source.t21 a_n2224_n2688# 2.47528f
C275 source.n36 a_n2224_n2688# 0.507203f
C276 source.t1 a_n2224_n2688# 0.232127f
C277 source.t22 a_n2224_n2688# 0.232127f
C278 source.n37 a_n2224_n2688# 1.94321f
C279 source.n38 a_n2224_n2688# 0.40937f
C280 source.t14 a_n2224_n2688# 0.232127f
C281 source.t9 a_n2224_n2688# 0.232127f
C282 source.n39 a_n2224_n2688# 1.94321f
C283 source.n40 a_n2224_n2688# 0.40937f
C284 source.t16 a_n2224_n2688# 0.232127f
C285 source.t17 a_n2224_n2688# 0.232127f
C286 source.n41 a_n2224_n2688# 1.94321f
C287 source.n42 a_n2224_n2688# 0.40937f
C288 source.t4 a_n2224_n2688# 0.232127f
C289 source.t23 a_n2224_n2688# 0.232127f
C290 source.n43 a_n2224_n2688# 1.94321f
C291 source.n44 a_n2224_n2688# 0.40937f
C292 source.t0 a_n2224_n2688# 0.232127f
C293 source.t8 a_n2224_n2688# 0.232127f
C294 source.n45 a_n2224_n2688# 1.94321f
C295 source.n46 a_n2224_n2688# 0.40937f
C296 source.t2 a_n2224_n2688# 2.47528f
C297 source.n47 a_n2224_n2688# 0.687818f
C298 source.n48 a_n2224_n2688# 1.69668f
C299 plus.n0 a_n2224_n2688# 0.050924f
C300 plus.t18 a_n2224_n2688# 0.324669f
C301 plus.t4 a_n2224_n2688# 0.324669f
C302 plus.n1 a_n2224_n2688# 0.018463f
C303 plus.n2 a_n2224_n2688# 0.050924f
C304 plus.t5 a_n2224_n2688# 0.324669f
C305 plus.t12 a_n2224_n2688# 0.324669f
C306 plus.t23 a_n2224_n2688# 0.324669f
C307 plus.n3 a_n2224_n2688# 0.138192f
C308 plus.n4 a_n2224_n2688# 0.050924f
C309 plus.t13 a_n2224_n2688# 0.324669f
C310 plus.t0 a_n2224_n2688# 0.324669f
C311 plus.n5 a_n2224_n2688# 0.017835f
C312 plus.t8 a_n2224_n2688# 0.328375f
C313 plus.n6 a_n2224_n2688# 0.152072f
C314 plus.t1 a_n2224_n2688# 0.324669f
C315 plus.n7 a_n2224_n2688# 0.138192f
C316 plus.t14 a_n2224_n2688# 0.324669f
C317 plus.n8 a_n2224_n2688# 0.138192f
C318 plus.n9 a_n2224_n2688# 0.019405f
C319 plus.n10 a_n2224_n2688# 0.105864f
C320 plus.n11 a_n2224_n2688# 0.050924f
C321 plus.n12 a_n2224_n2688# 0.050924f
C322 plus.n13 a_n2224_n2688# 0.018463f
C323 plus.n14 a_n2224_n2688# 0.138192f
C324 plus.n15 a_n2224_n2688# 0.019405f
C325 plus.n16 a_n2224_n2688# 0.138192f
C326 plus.n17 a_n2224_n2688# 0.019405f
C327 plus.n18 a_n2224_n2688# 0.050924f
C328 plus.n19 a_n2224_n2688# 0.050924f
C329 plus.n20 a_n2224_n2688# 0.019405f
C330 plus.n21 a_n2224_n2688# 0.138192f
C331 plus.n22 a_n2224_n2688# 0.019405f
C332 plus.n23 a_n2224_n2688# 0.138192f
C333 plus.t19 a_n2224_n2688# 0.324669f
C334 plus.n24 a_n2224_n2688# 0.138192f
C335 plus.n25 a_n2224_n2688# 0.019405f
C336 plus.n26 a_n2224_n2688# 0.050924f
C337 plus.n27 a_n2224_n2688# 0.050924f
C338 plus.n28 a_n2224_n2688# 0.050924f
C339 plus.n29 a_n2224_n2688# 0.017835f
C340 plus.n30 a_n2224_n2688# 0.138192f
C341 plus.n31 a_n2224_n2688# 0.019405f
C342 plus.n32 a_n2224_n2688# 0.138192f
C343 plus.t3 a_n2224_n2688# 0.328375f
C344 plus.n33 a_n2224_n2688# 0.152007f
C345 plus.n34 a_n2224_n2688# 0.491843f
C346 plus.n35 a_n2224_n2688# 0.050924f
C347 plus.t9 a_n2224_n2688# 0.328375f
C348 plus.t10 a_n2224_n2688# 0.324669f
C349 plus.t11 a_n2224_n2688# 0.324669f
C350 plus.n36 a_n2224_n2688# 0.018463f
C351 plus.n37 a_n2224_n2688# 0.050924f
C352 plus.t17 a_n2224_n2688# 0.324669f
C353 plus.n38 a_n2224_n2688# 0.138192f
C354 plus.t6 a_n2224_n2688# 0.324669f
C355 plus.t15 a_n2224_n2688# 0.324669f
C356 plus.t20 a_n2224_n2688# 0.324669f
C357 plus.n39 a_n2224_n2688# 0.138192f
C358 plus.n40 a_n2224_n2688# 0.050924f
C359 plus.t2 a_n2224_n2688# 0.324669f
C360 plus.t22 a_n2224_n2688# 0.324669f
C361 plus.n41 a_n2224_n2688# 0.017835f
C362 plus.t21 a_n2224_n2688# 0.328375f
C363 plus.n42 a_n2224_n2688# 0.152072f
C364 plus.t7 a_n2224_n2688# 0.324669f
C365 plus.n43 a_n2224_n2688# 0.138192f
C366 plus.t16 a_n2224_n2688# 0.324669f
C367 plus.n44 a_n2224_n2688# 0.138192f
C368 plus.n45 a_n2224_n2688# 0.019405f
C369 plus.n46 a_n2224_n2688# 0.105864f
C370 plus.n47 a_n2224_n2688# 0.050924f
C371 plus.n48 a_n2224_n2688# 0.050924f
C372 plus.n49 a_n2224_n2688# 0.018463f
C373 plus.n50 a_n2224_n2688# 0.138192f
C374 plus.n51 a_n2224_n2688# 0.019405f
C375 plus.n52 a_n2224_n2688# 0.138192f
C376 plus.n53 a_n2224_n2688# 0.019405f
C377 plus.n54 a_n2224_n2688# 0.050924f
C378 plus.n55 a_n2224_n2688# 0.050924f
C379 plus.n56 a_n2224_n2688# 0.019405f
C380 plus.n57 a_n2224_n2688# 0.138192f
C381 plus.n58 a_n2224_n2688# 0.019405f
C382 plus.n59 a_n2224_n2688# 0.138192f
C383 plus.n60 a_n2224_n2688# 0.019405f
C384 plus.n61 a_n2224_n2688# 0.050924f
C385 plus.n62 a_n2224_n2688# 0.050924f
C386 plus.n63 a_n2224_n2688# 0.050924f
C387 plus.n64 a_n2224_n2688# 0.017835f
C388 plus.n65 a_n2224_n2688# 0.138192f
C389 plus.n66 a_n2224_n2688# 0.019405f
C390 plus.n67 a_n2224_n2688# 0.138192f
C391 plus.n68 a_n2224_n2688# 0.152007f
C392 plus.n69 a_n2224_n2688# 1.50234f
.ends

