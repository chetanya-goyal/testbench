* NGSPICE file created from diffpair306.ext - technology: sky130A

.subckt diffpair306 minus drain_right drain_left source plus
X0 a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X1 drain_left.t13 plus.t0 source.t26 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X2 source.t18 plus.t1 drain_left.t12 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 drain_left.t11 plus.t2 source.t20 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 source.t6 minus.t0 drain_right.t13 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X5 drain_left.t10 plus.t3 source.t22 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X6 a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X7 drain_left.t9 plus.t4 source.t24 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X8 drain_left.t8 plus.t5 source.t14 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X9 drain_left.t7 plus.t6 source.t16 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X10 drain_right.t12 minus.t1 source.t7 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X11 source.t9 minus.t2 drain_right.t11 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 drain_right.t10 minus.t3 source.t5 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 drain_right.t9 minus.t4 source.t13 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X14 drain_left.t6 plus.t7 source.t15 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X15 drain_right.t8 minus.t5 source.t2 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X16 drain_right.t7 minus.t6 source.t1 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X17 source.t27 plus.t8 drain_left.t5 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X18 source.t17 plus.t9 drain_left.t4 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X19 source.t3 minus.t7 drain_right.t6 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X20 source.t19 plus.t10 drain_left.t3 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X21 drain_right.t5 minus.t8 source.t4 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X22 a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X23 drain_right.t4 minus.t9 source.t8 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X24 source.t21 plus.t11 drain_left.t2 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X25 source.t23 plus.t12 drain_left.t1 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X26 drain_left.t0 plus.t13 source.t25 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X27 drain_right.t3 minus.t10 source.t10 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X28 source.t0 minus.t11 drain_right.t2 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X29 a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X30 source.t12 minus.t12 drain_right.t1 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X31 source.t11 minus.t13 drain_right.t0 a_n2364_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n5 plus.t5 286.536
R1 plus.n27 plus.t7 286.536
R2 plus.n20 plus.t0 262.69
R3 plus.n18 plus.t10 262.69
R4 plus.n2 plus.t4 262.69
R5 plus.n12 plus.t9 262.69
R6 plus.n4 plus.t2 262.69
R7 plus.n6 plus.t11 262.69
R8 plus.n42 plus.t13 262.69
R9 plus.n40 plus.t12 262.69
R10 plus.n24 plus.t3 262.69
R11 plus.n34 plus.t1 262.69
R12 plus.n26 plus.t6 262.69
R13 plus.n28 plus.t8 262.69
R14 plus.n8 plus.n7 161.3
R15 plus.n9 plus.n4 161.3
R16 plus.n11 plus.n10 161.3
R17 plus.n12 plus.n3 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n15 plus.n2 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n18 plus.n1 161.3
R22 plus.n19 plus.n0 161.3
R23 plus.n21 plus.n20 161.3
R24 plus.n30 plus.n29 161.3
R25 plus.n31 plus.n26 161.3
R26 plus.n33 plus.n32 161.3
R27 plus.n34 plus.n25 161.3
R28 plus.n36 plus.n35 161.3
R29 plus.n37 plus.n24 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n40 plus.n23 161.3
R32 plus.n41 plus.n22 161.3
R33 plus.n43 plus.n42 161.3
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus.n18 plus.n17 30.6732
R39 plus.n7 plus.n6 30.6732
R40 plus.n40 plus.n39 30.6732
R41 plus.n29 plus.n28 30.6732
R42 plus plus.n43 29.8342
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus.n19 plus.n18 13.146
R58 plus.n41 plus.n40 13.146
R59 plus plus.n21 10.0213
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n146 source.n120 289.615
R79 source.n108 source.n82 289.615
R80 source.n26 source.n0 289.615
R81 source.n64 source.n38 289.615
R82 source.n131 source.n130 185
R83 source.n128 source.n127 185
R84 source.n137 source.n136 185
R85 source.n139 source.n138 185
R86 source.n124 source.n123 185
R87 source.n145 source.n144 185
R88 source.n147 source.n146 185
R89 source.n93 source.n92 185
R90 source.n90 source.n89 185
R91 source.n99 source.n98 185
R92 source.n101 source.n100 185
R93 source.n86 source.n85 185
R94 source.n107 source.n106 185
R95 source.n109 source.n108 185
R96 source.n27 source.n26 185
R97 source.n25 source.n24 185
R98 source.n4 source.n3 185
R99 source.n19 source.n18 185
R100 source.n17 source.n16 185
R101 source.n8 source.n7 185
R102 source.n11 source.n10 185
R103 source.n65 source.n64 185
R104 source.n63 source.n62 185
R105 source.n42 source.n41 185
R106 source.n57 source.n56 185
R107 source.n55 source.n54 185
R108 source.n46 source.n45 185
R109 source.n49 source.n48 185
R110 source.t13 source.n129 147.661
R111 source.t15 source.n91 147.661
R112 source.t26 source.n9 147.661
R113 source.t4 source.n47 147.661
R114 source.n130 source.n127 104.615
R115 source.n137 source.n127 104.615
R116 source.n138 source.n137 104.615
R117 source.n138 source.n123 104.615
R118 source.n145 source.n123 104.615
R119 source.n146 source.n145 104.615
R120 source.n92 source.n89 104.615
R121 source.n99 source.n89 104.615
R122 source.n100 source.n99 104.615
R123 source.n100 source.n85 104.615
R124 source.n107 source.n85 104.615
R125 source.n108 source.n107 104.615
R126 source.n26 source.n25 104.615
R127 source.n25 source.n3 104.615
R128 source.n18 source.n3 104.615
R129 source.n18 source.n17 104.615
R130 source.n17 source.n7 104.615
R131 source.n10 source.n7 104.615
R132 source.n64 source.n63 104.615
R133 source.n63 source.n41 104.615
R134 source.n56 source.n41 104.615
R135 source.n56 source.n55 104.615
R136 source.n55 source.n45 104.615
R137 source.n48 source.n45 104.615
R138 source.n130 source.t13 52.3082
R139 source.n92 source.t15 52.3082
R140 source.n10 source.t26 52.3082
R141 source.n48 source.t4 52.3082
R142 source.n33 source.n32 50.512
R143 source.n35 source.n34 50.512
R144 source.n37 source.n36 50.512
R145 source.n71 source.n70 50.512
R146 source.n73 source.n72 50.512
R147 source.n75 source.n74 50.512
R148 source.n119 source.n118 50.5119
R149 source.n117 source.n116 50.5119
R150 source.n115 source.n114 50.5119
R151 source.n81 source.n80 50.5119
R152 source.n79 source.n78 50.5119
R153 source.n77 source.n76 50.5119
R154 source.n151 source.n150 32.1853
R155 source.n113 source.n112 32.1853
R156 source.n31 source.n30 32.1853
R157 source.n69 source.n68 32.1853
R158 source.n77 source.n75 18.5181
R159 source.n131 source.n129 15.6674
R160 source.n93 source.n91 15.6674
R161 source.n11 source.n9 15.6674
R162 source.n49 source.n47 15.6674
R163 source.n132 source.n128 12.8005
R164 source.n94 source.n90 12.8005
R165 source.n12 source.n8 12.8005
R166 source.n50 source.n46 12.8005
R167 source.n136 source.n135 12.0247
R168 source.n98 source.n97 12.0247
R169 source.n16 source.n15 12.0247
R170 source.n54 source.n53 12.0247
R171 source.n152 source.n31 11.9233
R172 source.n139 source.n126 11.249
R173 source.n101 source.n88 11.249
R174 source.n19 source.n6 11.249
R175 source.n57 source.n44 11.249
R176 source.n140 source.n124 10.4732
R177 source.n102 source.n86 10.4732
R178 source.n20 source.n4 10.4732
R179 source.n58 source.n42 10.4732
R180 source.n144 source.n143 9.69747
R181 source.n106 source.n105 9.69747
R182 source.n24 source.n23 9.69747
R183 source.n62 source.n61 9.69747
R184 source.n150 source.n149 9.45567
R185 source.n112 source.n111 9.45567
R186 source.n30 source.n29 9.45567
R187 source.n68 source.n67 9.45567
R188 source.n149 source.n148 9.3005
R189 source.n122 source.n121 9.3005
R190 source.n143 source.n142 9.3005
R191 source.n141 source.n140 9.3005
R192 source.n126 source.n125 9.3005
R193 source.n135 source.n134 9.3005
R194 source.n133 source.n132 9.3005
R195 source.n111 source.n110 9.3005
R196 source.n84 source.n83 9.3005
R197 source.n105 source.n104 9.3005
R198 source.n103 source.n102 9.3005
R199 source.n88 source.n87 9.3005
R200 source.n97 source.n96 9.3005
R201 source.n95 source.n94 9.3005
R202 source.n29 source.n28 9.3005
R203 source.n2 source.n1 9.3005
R204 source.n23 source.n22 9.3005
R205 source.n21 source.n20 9.3005
R206 source.n6 source.n5 9.3005
R207 source.n15 source.n14 9.3005
R208 source.n13 source.n12 9.3005
R209 source.n67 source.n66 9.3005
R210 source.n40 source.n39 9.3005
R211 source.n61 source.n60 9.3005
R212 source.n59 source.n58 9.3005
R213 source.n44 source.n43 9.3005
R214 source.n53 source.n52 9.3005
R215 source.n51 source.n50 9.3005
R216 source.n147 source.n122 8.92171
R217 source.n109 source.n84 8.92171
R218 source.n27 source.n2 8.92171
R219 source.n65 source.n40 8.92171
R220 source.n148 source.n120 8.14595
R221 source.n110 source.n82 8.14595
R222 source.n28 source.n0 8.14595
R223 source.n66 source.n38 8.14595
R224 source.n150 source.n120 5.81868
R225 source.n112 source.n82 5.81868
R226 source.n30 source.n0 5.81868
R227 source.n68 source.n38 5.81868
R228 source.n152 source.n151 5.7074
R229 source.n148 source.n147 5.04292
R230 source.n110 source.n109 5.04292
R231 source.n28 source.n27 5.04292
R232 source.n66 source.n65 5.04292
R233 source.n133 source.n129 4.38594
R234 source.n95 source.n91 4.38594
R235 source.n13 source.n9 4.38594
R236 source.n51 source.n47 4.38594
R237 source.n144 source.n122 4.26717
R238 source.n106 source.n84 4.26717
R239 source.n24 source.n2 4.26717
R240 source.n62 source.n40 4.26717
R241 source.n143 source.n124 3.49141
R242 source.n105 source.n86 3.49141
R243 source.n23 source.n4 3.49141
R244 source.n61 source.n42 3.49141
R245 source.n118 source.t8 3.3005
R246 source.n118 source.t9 3.3005
R247 source.n116 source.t1 3.3005
R248 source.n116 source.t3 3.3005
R249 source.n114 source.t10 3.3005
R250 source.n114 source.t0 3.3005
R251 source.n80 source.t16 3.3005
R252 source.n80 source.t27 3.3005
R253 source.n78 source.t22 3.3005
R254 source.n78 source.t18 3.3005
R255 source.n76 source.t25 3.3005
R256 source.n76 source.t23 3.3005
R257 source.n32 source.t24 3.3005
R258 source.n32 source.t19 3.3005
R259 source.n34 source.t20 3.3005
R260 source.n34 source.t17 3.3005
R261 source.n36 source.t14 3.3005
R262 source.n36 source.t21 3.3005
R263 source.n70 source.t2 3.3005
R264 source.n70 source.t6 3.3005
R265 source.n72 source.t5 3.3005
R266 source.n72 source.t12 3.3005
R267 source.n74 source.t7 3.3005
R268 source.n74 source.t11 3.3005
R269 source.n140 source.n139 2.71565
R270 source.n102 source.n101 2.71565
R271 source.n20 source.n19 2.71565
R272 source.n58 source.n57 2.71565
R273 source.n136 source.n126 1.93989
R274 source.n98 source.n88 1.93989
R275 source.n16 source.n6 1.93989
R276 source.n54 source.n44 1.93989
R277 source.n135 source.n128 1.16414
R278 source.n97 source.n90 1.16414
R279 source.n15 source.n8 1.16414
R280 source.n53 source.n46 1.16414
R281 source.n69 source.n37 0.914293
R282 source.n115 source.n113 0.914293
R283 source.n75 source.n73 0.888431
R284 source.n73 source.n71 0.888431
R285 source.n71 source.n69 0.888431
R286 source.n37 source.n35 0.888431
R287 source.n35 source.n33 0.888431
R288 source.n33 source.n31 0.888431
R289 source.n79 source.n77 0.888431
R290 source.n81 source.n79 0.888431
R291 source.n113 source.n81 0.888431
R292 source.n117 source.n115 0.888431
R293 source.n119 source.n117 0.888431
R294 source.n151 source.n119 0.888431
R295 source.n132 source.n131 0.388379
R296 source.n94 source.n93 0.388379
R297 source.n12 source.n11 0.388379
R298 source.n50 source.n49 0.388379
R299 source source.n152 0.188
R300 source.n134 source.n133 0.155672
R301 source.n134 source.n125 0.155672
R302 source.n141 source.n125 0.155672
R303 source.n142 source.n141 0.155672
R304 source.n142 source.n121 0.155672
R305 source.n149 source.n121 0.155672
R306 source.n96 source.n95 0.155672
R307 source.n96 source.n87 0.155672
R308 source.n103 source.n87 0.155672
R309 source.n104 source.n103 0.155672
R310 source.n104 source.n83 0.155672
R311 source.n111 source.n83 0.155672
R312 source.n29 source.n1 0.155672
R313 source.n22 source.n1 0.155672
R314 source.n22 source.n21 0.155672
R315 source.n21 source.n5 0.155672
R316 source.n14 source.n5 0.155672
R317 source.n14 source.n13 0.155672
R318 source.n67 source.n39 0.155672
R319 source.n60 source.n39 0.155672
R320 source.n60 source.n59 0.155672
R321 source.n59 source.n43 0.155672
R322 source.n52 source.n43 0.155672
R323 source.n52 source.n51 0.155672
R324 drain_left.n26 drain_left.n0 289.615
R325 drain_left.n63 drain_left.n37 289.615
R326 drain_left.n11 drain_left.n10 185
R327 drain_left.n8 drain_left.n7 185
R328 drain_left.n17 drain_left.n16 185
R329 drain_left.n19 drain_left.n18 185
R330 drain_left.n4 drain_left.n3 185
R331 drain_left.n25 drain_left.n24 185
R332 drain_left.n27 drain_left.n26 185
R333 drain_left.n64 drain_left.n63 185
R334 drain_left.n62 drain_left.n61 185
R335 drain_left.n41 drain_left.n40 185
R336 drain_left.n56 drain_left.n55 185
R337 drain_left.n54 drain_left.n53 185
R338 drain_left.n45 drain_left.n44 185
R339 drain_left.n48 drain_left.n47 185
R340 drain_left.t0 drain_left.n9 147.661
R341 drain_left.t8 drain_left.n46 147.661
R342 drain_left.n10 drain_left.n7 104.615
R343 drain_left.n17 drain_left.n7 104.615
R344 drain_left.n18 drain_left.n17 104.615
R345 drain_left.n18 drain_left.n3 104.615
R346 drain_left.n25 drain_left.n3 104.615
R347 drain_left.n26 drain_left.n25 104.615
R348 drain_left.n63 drain_left.n62 104.615
R349 drain_left.n62 drain_left.n40 104.615
R350 drain_left.n55 drain_left.n40 104.615
R351 drain_left.n55 drain_left.n54 104.615
R352 drain_left.n54 drain_left.n44 104.615
R353 drain_left.n47 drain_left.n44 104.615
R354 drain_left.n35 drain_left.n33 68.0786
R355 drain_left.n71 drain_left.n70 67.1908
R356 drain_left.n69 drain_left.n68 67.1908
R357 drain_left.n73 drain_left.n72 67.1907
R358 drain_left.n35 drain_left.n34 67.1907
R359 drain_left.n32 drain_left.n31 67.1907
R360 drain_left.n10 drain_left.t0 52.3082
R361 drain_left.n47 drain_left.t8 52.3082
R362 drain_left.n32 drain_left.n30 49.7521
R363 drain_left.n69 drain_left.n67 49.7521
R364 drain_left drain_left.n36 27.9272
R365 drain_left.n11 drain_left.n9 15.6674
R366 drain_left.n48 drain_left.n46 15.6674
R367 drain_left.n12 drain_left.n8 12.8005
R368 drain_left.n49 drain_left.n45 12.8005
R369 drain_left.n16 drain_left.n15 12.0247
R370 drain_left.n53 drain_left.n52 12.0247
R371 drain_left.n19 drain_left.n6 11.249
R372 drain_left.n56 drain_left.n43 11.249
R373 drain_left.n20 drain_left.n4 10.4732
R374 drain_left.n57 drain_left.n41 10.4732
R375 drain_left.n24 drain_left.n23 9.69747
R376 drain_left.n61 drain_left.n60 9.69747
R377 drain_left.n30 drain_left.n29 9.45567
R378 drain_left.n67 drain_left.n66 9.45567
R379 drain_left.n29 drain_left.n28 9.3005
R380 drain_left.n2 drain_left.n1 9.3005
R381 drain_left.n23 drain_left.n22 9.3005
R382 drain_left.n21 drain_left.n20 9.3005
R383 drain_left.n6 drain_left.n5 9.3005
R384 drain_left.n15 drain_left.n14 9.3005
R385 drain_left.n13 drain_left.n12 9.3005
R386 drain_left.n66 drain_left.n65 9.3005
R387 drain_left.n39 drain_left.n38 9.3005
R388 drain_left.n60 drain_left.n59 9.3005
R389 drain_left.n58 drain_left.n57 9.3005
R390 drain_left.n43 drain_left.n42 9.3005
R391 drain_left.n52 drain_left.n51 9.3005
R392 drain_left.n50 drain_left.n49 9.3005
R393 drain_left.n27 drain_left.n2 8.92171
R394 drain_left.n64 drain_left.n39 8.92171
R395 drain_left.n28 drain_left.n0 8.14595
R396 drain_left.n65 drain_left.n37 8.14595
R397 drain_left drain_left.n73 6.54115
R398 drain_left.n30 drain_left.n0 5.81868
R399 drain_left.n67 drain_left.n37 5.81868
R400 drain_left.n28 drain_left.n27 5.04292
R401 drain_left.n65 drain_left.n64 5.04292
R402 drain_left.n13 drain_left.n9 4.38594
R403 drain_left.n50 drain_left.n46 4.38594
R404 drain_left.n24 drain_left.n2 4.26717
R405 drain_left.n61 drain_left.n39 4.26717
R406 drain_left.n23 drain_left.n4 3.49141
R407 drain_left.n60 drain_left.n41 3.49141
R408 drain_left.n33 drain_left.t5 3.3005
R409 drain_left.n33 drain_left.t6 3.3005
R410 drain_left.n34 drain_left.t12 3.3005
R411 drain_left.n34 drain_left.t7 3.3005
R412 drain_left.n31 drain_left.t1 3.3005
R413 drain_left.n31 drain_left.t10 3.3005
R414 drain_left.n72 drain_left.t3 3.3005
R415 drain_left.n72 drain_left.t13 3.3005
R416 drain_left.n70 drain_left.t4 3.3005
R417 drain_left.n70 drain_left.t9 3.3005
R418 drain_left.n68 drain_left.t2 3.3005
R419 drain_left.n68 drain_left.t11 3.3005
R420 drain_left.n20 drain_left.n19 2.71565
R421 drain_left.n57 drain_left.n56 2.71565
R422 drain_left.n16 drain_left.n6 1.93989
R423 drain_left.n53 drain_left.n43 1.93989
R424 drain_left.n15 drain_left.n8 1.16414
R425 drain_left.n52 drain_left.n45 1.16414
R426 drain_left.n71 drain_left.n69 0.888431
R427 drain_left.n73 drain_left.n71 0.888431
R428 drain_left.n36 drain_left.n32 0.611102
R429 drain_left.n12 drain_left.n11 0.388379
R430 drain_left.n49 drain_left.n48 0.388379
R431 drain_left.n36 drain_left.n35 0.167137
R432 drain_left.n14 drain_left.n13 0.155672
R433 drain_left.n14 drain_left.n5 0.155672
R434 drain_left.n21 drain_left.n5 0.155672
R435 drain_left.n22 drain_left.n21 0.155672
R436 drain_left.n22 drain_left.n1 0.155672
R437 drain_left.n29 drain_left.n1 0.155672
R438 drain_left.n66 drain_left.n38 0.155672
R439 drain_left.n59 drain_left.n38 0.155672
R440 drain_left.n59 drain_left.n58 0.155672
R441 drain_left.n58 drain_left.n42 0.155672
R442 drain_left.n51 drain_left.n42 0.155672
R443 drain_left.n51 drain_left.n50 0.155672
R444 minus.n5 minus.t8 286.536
R445 minus.n27 minus.t10 286.536
R446 minus.n6 minus.t0 262.69
R447 minus.n8 minus.t5 262.69
R448 minus.n12 minus.t12 262.69
R449 minus.n14 minus.t3 262.69
R450 minus.n18 minus.t13 262.69
R451 minus.n20 minus.t1 262.69
R452 minus.n28 minus.t11 262.69
R453 minus.n30 minus.t6 262.69
R454 minus.n34 minus.t7 262.69
R455 minus.n36 minus.t9 262.69
R456 minus.n40 minus.t2 262.69
R457 minus.n42 minus.t4 262.69
R458 minus.n21 minus.n20 161.3
R459 minus.n19 minus.n0 161.3
R460 minus.n18 minus.n17 161.3
R461 minus.n16 minus.n1 161.3
R462 minus.n15 minus.n14 161.3
R463 minus.n13 minus.n2 161.3
R464 minus.n12 minus.n11 161.3
R465 minus.n10 minus.n3 161.3
R466 minus.n9 minus.n8 161.3
R467 minus.n7 minus.n4 161.3
R468 minus.n43 minus.n42 161.3
R469 minus.n41 minus.n22 161.3
R470 minus.n40 minus.n39 161.3
R471 minus.n38 minus.n23 161.3
R472 minus.n37 minus.n36 161.3
R473 minus.n35 minus.n24 161.3
R474 minus.n34 minus.n33 161.3
R475 minus.n32 minus.n25 161.3
R476 minus.n31 minus.n30 161.3
R477 minus.n29 minus.n26 161.3
R478 minus.n5 minus.n4 44.9119
R479 minus.n27 minus.n26 44.9119
R480 minus.n20 minus.n19 35.055
R481 minus.n42 minus.n41 35.055
R482 minus.n44 minus.n21 33.6804
R483 minus.n7 minus.n6 30.6732
R484 minus.n18 minus.n1 30.6732
R485 minus.n29 minus.n28 30.6732
R486 minus.n40 minus.n23 30.6732
R487 minus.n8 minus.n3 26.2914
R488 minus.n14 minus.n13 26.2914
R489 minus.n30 minus.n25 26.2914
R490 minus.n36 minus.n35 26.2914
R491 minus.n12 minus.n3 21.9096
R492 minus.n13 minus.n12 21.9096
R493 minus.n34 minus.n25 21.9096
R494 minus.n35 minus.n34 21.9096
R495 minus.n6 minus.n5 17.739
R496 minus.n28 minus.n27 17.739
R497 minus.n8 minus.n7 17.5278
R498 minus.n14 minus.n1 17.5278
R499 minus.n30 minus.n29 17.5278
R500 minus.n36 minus.n23 17.5278
R501 minus.n19 minus.n18 13.146
R502 minus.n41 minus.n40 13.146
R503 minus.n44 minus.n43 6.65012
R504 minus.n21 minus.n0 0.189894
R505 minus.n17 minus.n0 0.189894
R506 minus.n17 minus.n16 0.189894
R507 minus.n16 minus.n15 0.189894
R508 minus.n15 minus.n2 0.189894
R509 minus.n11 minus.n2 0.189894
R510 minus.n11 minus.n10 0.189894
R511 minus.n10 minus.n9 0.189894
R512 minus.n9 minus.n4 0.189894
R513 minus.n31 minus.n26 0.189894
R514 minus.n32 minus.n31 0.189894
R515 minus.n33 minus.n32 0.189894
R516 minus.n33 minus.n24 0.189894
R517 minus.n37 minus.n24 0.189894
R518 minus.n38 minus.n37 0.189894
R519 minus.n39 minus.n38 0.189894
R520 minus.n39 minus.n22 0.189894
R521 minus.n43 minus.n22 0.189894
R522 minus minus.n44 0.188
R523 drain_right.n26 drain_right.n0 289.615
R524 drain_right.n68 drain_right.n42 289.615
R525 drain_right.n11 drain_right.n10 185
R526 drain_right.n8 drain_right.n7 185
R527 drain_right.n17 drain_right.n16 185
R528 drain_right.n19 drain_right.n18 185
R529 drain_right.n4 drain_right.n3 185
R530 drain_right.n25 drain_right.n24 185
R531 drain_right.n27 drain_right.n26 185
R532 drain_right.n69 drain_right.n68 185
R533 drain_right.n67 drain_right.n66 185
R534 drain_right.n46 drain_right.n45 185
R535 drain_right.n61 drain_right.n60 185
R536 drain_right.n59 drain_right.n58 185
R537 drain_right.n50 drain_right.n49 185
R538 drain_right.n53 drain_right.n52 185
R539 drain_right.t3 drain_right.n9 147.661
R540 drain_right.t12 drain_right.n51 147.661
R541 drain_right.n10 drain_right.n7 104.615
R542 drain_right.n17 drain_right.n7 104.615
R543 drain_right.n18 drain_right.n17 104.615
R544 drain_right.n18 drain_right.n3 104.615
R545 drain_right.n25 drain_right.n3 104.615
R546 drain_right.n26 drain_right.n25 104.615
R547 drain_right.n68 drain_right.n67 104.615
R548 drain_right.n67 drain_right.n45 104.615
R549 drain_right.n60 drain_right.n45 104.615
R550 drain_right.n60 drain_right.n59 104.615
R551 drain_right.n59 drain_right.n49 104.615
R552 drain_right.n52 drain_right.n49 104.615
R553 drain_right.n39 drain_right.n37 68.0786
R554 drain_right.n35 drain_right.n33 68.0786
R555 drain_right.n39 drain_right.n38 67.1908
R556 drain_right.n41 drain_right.n40 67.1908
R557 drain_right.n35 drain_right.n34 67.1907
R558 drain_right.n32 drain_right.n31 67.1907
R559 drain_right.n10 drain_right.t3 52.3082
R560 drain_right.n52 drain_right.t12 52.3082
R561 drain_right.n32 drain_right.n30 49.7521
R562 drain_right.n73 drain_right.n72 48.8641
R563 drain_right drain_right.n36 27.374
R564 drain_right.n11 drain_right.n9 15.6674
R565 drain_right.n53 drain_right.n51 15.6674
R566 drain_right.n12 drain_right.n8 12.8005
R567 drain_right.n54 drain_right.n50 12.8005
R568 drain_right.n16 drain_right.n15 12.0247
R569 drain_right.n58 drain_right.n57 12.0247
R570 drain_right.n19 drain_right.n6 11.249
R571 drain_right.n61 drain_right.n48 11.249
R572 drain_right.n20 drain_right.n4 10.4732
R573 drain_right.n62 drain_right.n46 10.4732
R574 drain_right.n24 drain_right.n23 9.69747
R575 drain_right.n66 drain_right.n65 9.69747
R576 drain_right.n30 drain_right.n29 9.45567
R577 drain_right.n72 drain_right.n71 9.45567
R578 drain_right.n29 drain_right.n28 9.3005
R579 drain_right.n2 drain_right.n1 9.3005
R580 drain_right.n23 drain_right.n22 9.3005
R581 drain_right.n21 drain_right.n20 9.3005
R582 drain_right.n6 drain_right.n5 9.3005
R583 drain_right.n15 drain_right.n14 9.3005
R584 drain_right.n13 drain_right.n12 9.3005
R585 drain_right.n71 drain_right.n70 9.3005
R586 drain_right.n44 drain_right.n43 9.3005
R587 drain_right.n65 drain_right.n64 9.3005
R588 drain_right.n63 drain_right.n62 9.3005
R589 drain_right.n48 drain_right.n47 9.3005
R590 drain_right.n57 drain_right.n56 9.3005
R591 drain_right.n55 drain_right.n54 9.3005
R592 drain_right.n27 drain_right.n2 8.92171
R593 drain_right.n69 drain_right.n44 8.92171
R594 drain_right.n28 drain_right.n0 8.14595
R595 drain_right.n70 drain_right.n42 8.14595
R596 drain_right drain_right.n73 6.09718
R597 drain_right.n30 drain_right.n0 5.81868
R598 drain_right.n72 drain_right.n42 5.81868
R599 drain_right.n28 drain_right.n27 5.04292
R600 drain_right.n70 drain_right.n69 5.04292
R601 drain_right.n13 drain_right.n9 4.38594
R602 drain_right.n55 drain_right.n51 4.38594
R603 drain_right.n24 drain_right.n2 4.26717
R604 drain_right.n66 drain_right.n44 4.26717
R605 drain_right.n23 drain_right.n4 3.49141
R606 drain_right.n65 drain_right.n46 3.49141
R607 drain_right.n33 drain_right.t11 3.3005
R608 drain_right.n33 drain_right.t9 3.3005
R609 drain_right.n34 drain_right.t6 3.3005
R610 drain_right.n34 drain_right.t4 3.3005
R611 drain_right.n31 drain_right.t2 3.3005
R612 drain_right.n31 drain_right.t7 3.3005
R613 drain_right.n37 drain_right.t13 3.3005
R614 drain_right.n37 drain_right.t5 3.3005
R615 drain_right.n38 drain_right.t1 3.3005
R616 drain_right.n38 drain_right.t8 3.3005
R617 drain_right.n40 drain_right.t0 3.3005
R618 drain_right.n40 drain_right.t10 3.3005
R619 drain_right.n20 drain_right.n19 2.71565
R620 drain_right.n62 drain_right.n61 2.71565
R621 drain_right.n16 drain_right.n6 1.93989
R622 drain_right.n58 drain_right.n48 1.93989
R623 drain_right.n15 drain_right.n8 1.16414
R624 drain_right.n57 drain_right.n50 1.16414
R625 drain_right.n73 drain_right.n41 0.888431
R626 drain_right.n41 drain_right.n39 0.888431
R627 drain_right.n36 drain_right.n32 0.611102
R628 drain_right.n12 drain_right.n11 0.388379
R629 drain_right.n54 drain_right.n53 0.388379
R630 drain_right.n36 drain_right.n35 0.167137
R631 drain_right.n14 drain_right.n13 0.155672
R632 drain_right.n14 drain_right.n5 0.155672
R633 drain_right.n21 drain_right.n5 0.155672
R634 drain_right.n22 drain_right.n21 0.155672
R635 drain_right.n22 drain_right.n1 0.155672
R636 drain_right.n29 drain_right.n1 0.155672
R637 drain_right.n71 drain_right.n43 0.155672
R638 drain_right.n64 drain_right.n43 0.155672
R639 drain_right.n64 drain_right.n63 0.155672
R640 drain_right.n63 drain_right.n47 0.155672
R641 drain_right.n56 drain_right.n47 0.155672
R642 drain_right.n56 drain_right.n55 0.155672
C0 drain_left plus 5.03919f
C1 source drain_left 10.932099f
C2 source plus 5.10992f
C3 drain_right drain_left 1.23199f
C4 drain_right plus 0.390107f
C5 minus drain_left 0.172675f
C6 minus plus 4.98137f
C7 source drain_right 10.9296f
C8 minus source 5.09565f
C9 minus drain_right 4.80719f
C10 drain_right a_n2364_n2088# 5.86045f
C11 drain_left a_n2364_n2088# 6.21486f
C12 source a_n2364_n2088# 4.292094f
C13 minus a_n2364_n2088# 8.873696f
C14 plus a_n2364_n2088# 10.31577f
C15 drain_right.n0 a_n2364_n2088# 0.035096f
C16 drain_right.n1 a_n2364_n2088# 0.024969f
C17 drain_right.n2 a_n2364_n2088# 0.013417f
C18 drain_right.n3 a_n2364_n2088# 0.031713f
C19 drain_right.n4 a_n2364_n2088# 0.014206f
C20 drain_right.n5 a_n2364_n2088# 0.024969f
C21 drain_right.n6 a_n2364_n2088# 0.013417f
C22 drain_right.n7 a_n2364_n2088# 0.031713f
C23 drain_right.n8 a_n2364_n2088# 0.014206f
C24 drain_right.n9 a_n2364_n2088# 0.106848f
C25 drain_right.t3 a_n2364_n2088# 0.051688f
C26 drain_right.n10 a_n2364_n2088# 0.023785f
C27 drain_right.n11 a_n2364_n2088# 0.018733f
C28 drain_right.n12 a_n2364_n2088# 0.013417f
C29 drain_right.n13 a_n2364_n2088# 0.594103f
C30 drain_right.n14 a_n2364_n2088# 0.024969f
C31 drain_right.n15 a_n2364_n2088# 0.013417f
C32 drain_right.n16 a_n2364_n2088# 0.014206f
C33 drain_right.n17 a_n2364_n2088# 0.031713f
C34 drain_right.n18 a_n2364_n2088# 0.031713f
C35 drain_right.n19 a_n2364_n2088# 0.014206f
C36 drain_right.n20 a_n2364_n2088# 0.013417f
C37 drain_right.n21 a_n2364_n2088# 0.024969f
C38 drain_right.n22 a_n2364_n2088# 0.024969f
C39 drain_right.n23 a_n2364_n2088# 0.013417f
C40 drain_right.n24 a_n2364_n2088# 0.014206f
C41 drain_right.n25 a_n2364_n2088# 0.031713f
C42 drain_right.n26 a_n2364_n2088# 0.068653f
C43 drain_right.n27 a_n2364_n2088# 0.014206f
C44 drain_right.n28 a_n2364_n2088# 0.013417f
C45 drain_right.n29 a_n2364_n2088# 0.057714f
C46 drain_right.n30 a_n2364_n2088# 0.057787f
C47 drain_right.t2 a_n2364_n2088# 0.118385f
C48 drain_right.t7 a_n2364_n2088# 0.118385f
C49 drain_right.n31 a_n2364_n2088# 0.987335f
C50 drain_right.n32 a_n2364_n2088# 0.441549f
C51 drain_right.t11 a_n2364_n2088# 0.118385f
C52 drain_right.t9 a_n2364_n2088# 0.118385f
C53 drain_right.n33 a_n2364_n2088# 0.991973f
C54 drain_right.t6 a_n2364_n2088# 0.118385f
C55 drain_right.t4 a_n2364_n2088# 0.118385f
C56 drain_right.n34 a_n2364_n2088# 0.987335f
C57 drain_right.n35 a_n2364_n2088# 0.64192f
C58 drain_right.n36 a_n2364_n2088# 1.00084f
C59 drain_right.t13 a_n2364_n2088# 0.118385f
C60 drain_right.t5 a_n2364_n2088# 0.118385f
C61 drain_right.n37 a_n2364_n2088# 0.991973f
C62 drain_right.t1 a_n2364_n2088# 0.118385f
C63 drain_right.t8 a_n2364_n2088# 0.118385f
C64 drain_right.n38 a_n2364_n2088# 0.98734f
C65 drain_right.n39 a_n2364_n2088# 0.696473f
C66 drain_right.t0 a_n2364_n2088# 0.118385f
C67 drain_right.t10 a_n2364_n2088# 0.118385f
C68 drain_right.n40 a_n2364_n2088# 0.98734f
C69 drain_right.n41 a_n2364_n2088# 0.345525f
C70 drain_right.n42 a_n2364_n2088# 0.035096f
C71 drain_right.n43 a_n2364_n2088# 0.024969f
C72 drain_right.n44 a_n2364_n2088# 0.013417f
C73 drain_right.n45 a_n2364_n2088# 0.031713f
C74 drain_right.n46 a_n2364_n2088# 0.014206f
C75 drain_right.n47 a_n2364_n2088# 0.024969f
C76 drain_right.n48 a_n2364_n2088# 0.013417f
C77 drain_right.n49 a_n2364_n2088# 0.031713f
C78 drain_right.n50 a_n2364_n2088# 0.014206f
C79 drain_right.n51 a_n2364_n2088# 0.106848f
C80 drain_right.t12 a_n2364_n2088# 0.051688f
C81 drain_right.n52 a_n2364_n2088# 0.023785f
C82 drain_right.n53 a_n2364_n2088# 0.018733f
C83 drain_right.n54 a_n2364_n2088# 0.013417f
C84 drain_right.n55 a_n2364_n2088# 0.594103f
C85 drain_right.n56 a_n2364_n2088# 0.024969f
C86 drain_right.n57 a_n2364_n2088# 0.013417f
C87 drain_right.n58 a_n2364_n2088# 0.014206f
C88 drain_right.n59 a_n2364_n2088# 0.031713f
C89 drain_right.n60 a_n2364_n2088# 0.031713f
C90 drain_right.n61 a_n2364_n2088# 0.014206f
C91 drain_right.n62 a_n2364_n2088# 0.013417f
C92 drain_right.n63 a_n2364_n2088# 0.024969f
C93 drain_right.n64 a_n2364_n2088# 0.024969f
C94 drain_right.n65 a_n2364_n2088# 0.013417f
C95 drain_right.n66 a_n2364_n2088# 0.014206f
C96 drain_right.n67 a_n2364_n2088# 0.031713f
C97 drain_right.n68 a_n2364_n2088# 0.068653f
C98 drain_right.n69 a_n2364_n2088# 0.014206f
C99 drain_right.n70 a_n2364_n2088# 0.013417f
C100 drain_right.n71 a_n2364_n2088# 0.057714f
C101 drain_right.n72 a_n2364_n2088# 0.055654f
C102 drain_right.n73 a_n2364_n2088# 0.348992f
C103 minus.n0 a_n2364_n2088# 0.042069f
C104 minus.n1 a_n2364_n2088# 0.009546f
C105 minus.t13 a_n2364_n2088# 0.512501f
C106 minus.n2 a_n2364_n2088# 0.042069f
C107 minus.n3 a_n2364_n2088# 0.009546f
C108 minus.t12 a_n2364_n2088# 0.512501f
C109 minus.n4 a_n2364_n2088# 0.177256f
C110 minus.t8 a_n2364_n2088# 0.532213f
C111 minus.n5 a_n2364_n2088# 0.220765f
C112 minus.t0 a_n2364_n2088# 0.512501f
C113 minus.n6 a_n2364_n2088# 0.242033f
C114 minus.n7 a_n2364_n2088# 0.009546f
C115 minus.t5 a_n2364_n2088# 0.512501f
C116 minus.n8 a_n2364_n2088# 0.236821f
C117 minus.n9 a_n2364_n2088# 0.042069f
C118 minus.n10 a_n2364_n2088# 0.042069f
C119 minus.n11 a_n2364_n2088# 0.042069f
C120 minus.n12 a_n2364_n2088# 0.236821f
C121 minus.n13 a_n2364_n2088# 0.009546f
C122 minus.t3 a_n2364_n2088# 0.512501f
C123 minus.n14 a_n2364_n2088# 0.236821f
C124 minus.n15 a_n2364_n2088# 0.042069f
C125 minus.n16 a_n2364_n2088# 0.042069f
C126 minus.n17 a_n2364_n2088# 0.042069f
C127 minus.n18 a_n2364_n2088# 0.236821f
C128 minus.n19 a_n2364_n2088# 0.009546f
C129 minus.t1 a_n2364_n2088# 0.512501f
C130 minus.n20 a_n2364_n2088# 0.235265f
C131 minus.n21 a_n2364_n2088# 1.33138f
C132 minus.n22 a_n2364_n2088# 0.042069f
C133 minus.n23 a_n2364_n2088# 0.009546f
C134 minus.n24 a_n2364_n2088# 0.042069f
C135 minus.n25 a_n2364_n2088# 0.009546f
C136 minus.n26 a_n2364_n2088# 0.177256f
C137 minus.t10 a_n2364_n2088# 0.532213f
C138 minus.n27 a_n2364_n2088# 0.220765f
C139 minus.t11 a_n2364_n2088# 0.512501f
C140 minus.n28 a_n2364_n2088# 0.242033f
C141 minus.n29 a_n2364_n2088# 0.009546f
C142 minus.t6 a_n2364_n2088# 0.512501f
C143 minus.n30 a_n2364_n2088# 0.236821f
C144 minus.n31 a_n2364_n2088# 0.042069f
C145 minus.n32 a_n2364_n2088# 0.042069f
C146 minus.n33 a_n2364_n2088# 0.042069f
C147 minus.t7 a_n2364_n2088# 0.512501f
C148 minus.n34 a_n2364_n2088# 0.236821f
C149 minus.n35 a_n2364_n2088# 0.009546f
C150 minus.t9 a_n2364_n2088# 0.512501f
C151 minus.n36 a_n2364_n2088# 0.236821f
C152 minus.n37 a_n2364_n2088# 0.042069f
C153 minus.n38 a_n2364_n2088# 0.042069f
C154 minus.n39 a_n2364_n2088# 0.042069f
C155 minus.t2 a_n2364_n2088# 0.512501f
C156 minus.n40 a_n2364_n2088# 0.236821f
C157 minus.n41 a_n2364_n2088# 0.009546f
C158 minus.t4 a_n2364_n2088# 0.512501f
C159 minus.n42 a_n2364_n2088# 0.235265f
C160 minus.n43 a_n2364_n2088# 0.289812f
C161 minus.n44 a_n2364_n2088# 1.62297f
C162 drain_left.n0 a_n2364_n2088# 0.035323f
C163 drain_left.n1 a_n2364_n2088# 0.02513f
C164 drain_left.n2 a_n2364_n2088# 0.013504f
C165 drain_left.n3 a_n2364_n2088# 0.031918f
C166 drain_left.n4 a_n2364_n2088# 0.014298f
C167 drain_left.n5 a_n2364_n2088# 0.02513f
C168 drain_left.n6 a_n2364_n2088# 0.013504f
C169 drain_left.n7 a_n2364_n2088# 0.031918f
C170 drain_left.n8 a_n2364_n2088# 0.014298f
C171 drain_left.n9 a_n2364_n2088# 0.10754f
C172 drain_left.t0 a_n2364_n2088# 0.052023f
C173 drain_left.n10 a_n2364_n2088# 0.023939f
C174 drain_left.n11 a_n2364_n2088# 0.018854f
C175 drain_left.n12 a_n2364_n2088# 0.013504f
C176 drain_left.n13 a_n2364_n2088# 0.597951f
C177 drain_left.n14 a_n2364_n2088# 0.02513f
C178 drain_left.n15 a_n2364_n2088# 0.013504f
C179 drain_left.n16 a_n2364_n2088# 0.014298f
C180 drain_left.n17 a_n2364_n2088# 0.031918f
C181 drain_left.n18 a_n2364_n2088# 0.031918f
C182 drain_left.n19 a_n2364_n2088# 0.014298f
C183 drain_left.n20 a_n2364_n2088# 0.013504f
C184 drain_left.n21 a_n2364_n2088# 0.02513f
C185 drain_left.n22 a_n2364_n2088# 0.02513f
C186 drain_left.n23 a_n2364_n2088# 0.013504f
C187 drain_left.n24 a_n2364_n2088# 0.014298f
C188 drain_left.n25 a_n2364_n2088# 0.031918f
C189 drain_left.n26 a_n2364_n2088# 0.069098f
C190 drain_left.n27 a_n2364_n2088# 0.014298f
C191 drain_left.n28 a_n2364_n2088# 0.013504f
C192 drain_left.n29 a_n2364_n2088# 0.058088f
C193 drain_left.n30 a_n2364_n2088# 0.058162f
C194 drain_left.t1 a_n2364_n2088# 0.119152f
C195 drain_left.t10 a_n2364_n2088# 0.119152f
C196 drain_left.n31 a_n2364_n2088# 0.993731f
C197 drain_left.n32 a_n2364_n2088# 0.444409f
C198 drain_left.t5 a_n2364_n2088# 0.119152f
C199 drain_left.t6 a_n2364_n2088# 0.119152f
C200 drain_left.n33 a_n2364_n2088# 0.998398f
C201 drain_left.t12 a_n2364_n2088# 0.119152f
C202 drain_left.t7 a_n2364_n2088# 0.119152f
C203 drain_left.n34 a_n2364_n2088# 0.993731f
C204 drain_left.n35 a_n2364_n2088# 0.646078f
C205 drain_left.n36 a_n2364_n2088# 1.05793f
C206 drain_left.n37 a_n2364_n2088# 0.035323f
C207 drain_left.n38 a_n2364_n2088# 0.02513f
C208 drain_left.n39 a_n2364_n2088# 0.013504f
C209 drain_left.n40 a_n2364_n2088# 0.031918f
C210 drain_left.n41 a_n2364_n2088# 0.014298f
C211 drain_left.n42 a_n2364_n2088# 0.02513f
C212 drain_left.n43 a_n2364_n2088# 0.013504f
C213 drain_left.n44 a_n2364_n2088# 0.031918f
C214 drain_left.n45 a_n2364_n2088# 0.014298f
C215 drain_left.n46 a_n2364_n2088# 0.10754f
C216 drain_left.t8 a_n2364_n2088# 0.052023f
C217 drain_left.n47 a_n2364_n2088# 0.023939f
C218 drain_left.n48 a_n2364_n2088# 0.018854f
C219 drain_left.n49 a_n2364_n2088# 0.013504f
C220 drain_left.n50 a_n2364_n2088# 0.597951f
C221 drain_left.n51 a_n2364_n2088# 0.02513f
C222 drain_left.n52 a_n2364_n2088# 0.013504f
C223 drain_left.n53 a_n2364_n2088# 0.014298f
C224 drain_left.n54 a_n2364_n2088# 0.031918f
C225 drain_left.n55 a_n2364_n2088# 0.031918f
C226 drain_left.n56 a_n2364_n2088# 0.014298f
C227 drain_left.n57 a_n2364_n2088# 0.013504f
C228 drain_left.n58 a_n2364_n2088# 0.02513f
C229 drain_left.n59 a_n2364_n2088# 0.02513f
C230 drain_left.n60 a_n2364_n2088# 0.013504f
C231 drain_left.n61 a_n2364_n2088# 0.014298f
C232 drain_left.n62 a_n2364_n2088# 0.031918f
C233 drain_left.n63 a_n2364_n2088# 0.069098f
C234 drain_left.n64 a_n2364_n2088# 0.014298f
C235 drain_left.n65 a_n2364_n2088# 0.013504f
C236 drain_left.n66 a_n2364_n2088# 0.058088f
C237 drain_left.n67 a_n2364_n2088# 0.058162f
C238 drain_left.t2 a_n2364_n2088# 0.119152f
C239 drain_left.t11 a_n2364_n2088# 0.119152f
C240 drain_left.n68 a_n2364_n2088# 0.993735f
C241 drain_left.n69 a_n2364_n2088# 0.465906f
C242 drain_left.t4 a_n2364_n2088# 0.119152f
C243 drain_left.t9 a_n2364_n2088# 0.119152f
C244 drain_left.n70 a_n2364_n2088# 0.993735f
C245 drain_left.n71 a_n2364_n2088# 0.347763f
C246 drain_left.t3 a_n2364_n2088# 0.119152f
C247 drain_left.t13 a_n2364_n2088# 0.119152f
C248 drain_left.n72 a_n2364_n2088# 0.993731f
C249 drain_left.n73 a_n2364_n2088# 0.570046f
C250 source.n0 a_n2364_n2088# 0.039549f
C251 source.n1 a_n2364_n2088# 0.028137f
C252 source.n2 a_n2364_n2088# 0.01512f
C253 source.n3 a_n2364_n2088# 0.035737f
C254 source.n4 a_n2364_n2088# 0.016009f
C255 source.n5 a_n2364_n2088# 0.028137f
C256 source.n6 a_n2364_n2088# 0.01512f
C257 source.n7 a_n2364_n2088# 0.035737f
C258 source.n8 a_n2364_n2088# 0.016009f
C259 source.n9 a_n2364_n2088# 0.120406f
C260 source.t26 a_n2364_n2088# 0.058247f
C261 source.n10 a_n2364_n2088# 0.026803f
C262 source.n11 a_n2364_n2088# 0.02111f
C263 source.n12 a_n2364_n2088# 0.01512f
C264 source.n13 a_n2364_n2088# 0.669491f
C265 source.n14 a_n2364_n2088# 0.028137f
C266 source.n15 a_n2364_n2088# 0.01512f
C267 source.n16 a_n2364_n2088# 0.016009f
C268 source.n17 a_n2364_n2088# 0.035737f
C269 source.n18 a_n2364_n2088# 0.035737f
C270 source.n19 a_n2364_n2088# 0.016009f
C271 source.n20 a_n2364_n2088# 0.01512f
C272 source.n21 a_n2364_n2088# 0.028137f
C273 source.n22 a_n2364_n2088# 0.028137f
C274 source.n23 a_n2364_n2088# 0.01512f
C275 source.n24 a_n2364_n2088# 0.016009f
C276 source.n25 a_n2364_n2088# 0.035737f
C277 source.n26 a_n2364_n2088# 0.077365f
C278 source.n27 a_n2364_n2088# 0.016009f
C279 source.n28 a_n2364_n2088# 0.01512f
C280 source.n29 a_n2364_n2088# 0.065037f
C281 source.n30 a_n2364_n2088# 0.043289f
C282 source.n31 a_n2364_n2088# 0.735037f
C283 source.t24 a_n2364_n2088# 0.133408f
C284 source.t19 a_n2364_n2088# 0.133408f
C285 source.n32 a_n2364_n2088# 1.03899f
C286 source.n33 a_n2364_n2088# 0.424763f
C287 source.t20 a_n2364_n2088# 0.133408f
C288 source.t17 a_n2364_n2088# 0.133408f
C289 source.n34 a_n2364_n2088# 1.03899f
C290 source.n35 a_n2364_n2088# 0.424763f
C291 source.t14 a_n2364_n2088# 0.133408f
C292 source.t21 a_n2364_n2088# 0.133408f
C293 source.n36 a_n2364_n2088# 1.03899f
C294 source.n37 a_n2364_n2088# 0.427107f
C295 source.n38 a_n2364_n2088# 0.039549f
C296 source.n39 a_n2364_n2088# 0.028137f
C297 source.n40 a_n2364_n2088# 0.01512f
C298 source.n41 a_n2364_n2088# 0.035737f
C299 source.n42 a_n2364_n2088# 0.016009f
C300 source.n43 a_n2364_n2088# 0.028137f
C301 source.n44 a_n2364_n2088# 0.01512f
C302 source.n45 a_n2364_n2088# 0.035737f
C303 source.n46 a_n2364_n2088# 0.016009f
C304 source.n47 a_n2364_n2088# 0.120406f
C305 source.t4 a_n2364_n2088# 0.058247f
C306 source.n48 a_n2364_n2088# 0.026803f
C307 source.n49 a_n2364_n2088# 0.02111f
C308 source.n50 a_n2364_n2088# 0.01512f
C309 source.n51 a_n2364_n2088# 0.669491f
C310 source.n52 a_n2364_n2088# 0.028137f
C311 source.n53 a_n2364_n2088# 0.01512f
C312 source.n54 a_n2364_n2088# 0.016009f
C313 source.n55 a_n2364_n2088# 0.035737f
C314 source.n56 a_n2364_n2088# 0.035737f
C315 source.n57 a_n2364_n2088# 0.016009f
C316 source.n58 a_n2364_n2088# 0.01512f
C317 source.n59 a_n2364_n2088# 0.028137f
C318 source.n60 a_n2364_n2088# 0.028137f
C319 source.n61 a_n2364_n2088# 0.01512f
C320 source.n62 a_n2364_n2088# 0.016009f
C321 source.n63 a_n2364_n2088# 0.035737f
C322 source.n64 a_n2364_n2088# 0.077365f
C323 source.n65 a_n2364_n2088# 0.016009f
C324 source.n66 a_n2364_n2088# 0.01512f
C325 source.n67 a_n2364_n2088# 0.065037f
C326 source.n68 a_n2364_n2088# 0.043289f
C327 source.n69 a_n2364_n2088# 0.187382f
C328 source.t2 a_n2364_n2088# 0.133408f
C329 source.t6 a_n2364_n2088# 0.133408f
C330 source.n70 a_n2364_n2088# 1.03899f
C331 source.n71 a_n2364_n2088# 0.424763f
C332 source.t5 a_n2364_n2088# 0.133408f
C333 source.t12 a_n2364_n2088# 0.133408f
C334 source.n72 a_n2364_n2088# 1.03899f
C335 source.n73 a_n2364_n2088# 0.424763f
C336 source.t7 a_n2364_n2088# 0.133408f
C337 source.t11 a_n2364_n2088# 0.133408f
C338 source.n74 a_n2364_n2088# 1.03899f
C339 source.n75 a_n2364_n2088# 1.42652f
C340 source.t25 a_n2364_n2088# 0.133408f
C341 source.t23 a_n2364_n2088# 0.133408f
C342 source.n76 a_n2364_n2088# 1.03898f
C343 source.n77 a_n2364_n2088# 1.42653f
C344 source.t22 a_n2364_n2088# 0.133408f
C345 source.t18 a_n2364_n2088# 0.133408f
C346 source.n78 a_n2364_n2088# 1.03898f
C347 source.n79 a_n2364_n2088# 0.42477f
C348 source.t16 a_n2364_n2088# 0.133408f
C349 source.t27 a_n2364_n2088# 0.133408f
C350 source.n80 a_n2364_n2088# 1.03898f
C351 source.n81 a_n2364_n2088# 0.42477f
C352 source.n82 a_n2364_n2088# 0.039549f
C353 source.n83 a_n2364_n2088# 0.028137f
C354 source.n84 a_n2364_n2088# 0.01512f
C355 source.n85 a_n2364_n2088# 0.035737f
C356 source.n86 a_n2364_n2088# 0.016009f
C357 source.n87 a_n2364_n2088# 0.028137f
C358 source.n88 a_n2364_n2088# 0.01512f
C359 source.n89 a_n2364_n2088# 0.035737f
C360 source.n90 a_n2364_n2088# 0.016009f
C361 source.n91 a_n2364_n2088# 0.120406f
C362 source.t15 a_n2364_n2088# 0.058247f
C363 source.n92 a_n2364_n2088# 0.026803f
C364 source.n93 a_n2364_n2088# 0.02111f
C365 source.n94 a_n2364_n2088# 0.01512f
C366 source.n95 a_n2364_n2088# 0.669491f
C367 source.n96 a_n2364_n2088# 0.028137f
C368 source.n97 a_n2364_n2088# 0.01512f
C369 source.n98 a_n2364_n2088# 0.016009f
C370 source.n99 a_n2364_n2088# 0.035737f
C371 source.n100 a_n2364_n2088# 0.035737f
C372 source.n101 a_n2364_n2088# 0.016009f
C373 source.n102 a_n2364_n2088# 0.01512f
C374 source.n103 a_n2364_n2088# 0.028137f
C375 source.n104 a_n2364_n2088# 0.028137f
C376 source.n105 a_n2364_n2088# 0.01512f
C377 source.n106 a_n2364_n2088# 0.016009f
C378 source.n107 a_n2364_n2088# 0.035737f
C379 source.n108 a_n2364_n2088# 0.077365f
C380 source.n109 a_n2364_n2088# 0.016009f
C381 source.n110 a_n2364_n2088# 0.01512f
C382 source.n111 a_n2364_n2088# 0.065037f
C383 source.n112 a_n2364_n2088# 0.043289f
C384 source.n113 a_n2364_n2088# 0.187382f
C385 source.t10 a_n2364_n2088# 0.133408f
C386 source.t0 a_n2364_n2088# 0.133408f
C387 source.n114 a_n2364_n2088# 1.03898f
C388 source.n115 a_n2364_n2088# 0.427114f
C389 source.t1 a_n2364_n2088# 0.133408f
C390 source.t3 a_n2364_n2088# 0.133408f
C391 source.n116 a_n2364_n2088# 1.03898f
C392 source.n117 a_n2364_n2088# 0.42477f
C393 source.t8 a_n2364_n2088# 0.133408f
C394 source.t9 a_n2364_n2088# 0.133408f
C395 source.n118 a_n2364_n2088# 1.03898f
C396 source.n119 a_n2364_n2088# 0.42477f
C397 source.n120 a_n2364_n2088# 0.039549f
C398 source.n121 a_n2364_n2088# 0.028137f
C399 source.n122 a_n2364_n2088# 0.01512f
C400 source.n123 a_n2364_n2088# 0.035737f
C401 source.n124 a_n2364_n2088# 0.016009f
C402 source.n125 a_n2364_n2088# 0.028137f
C403 source.n126 a_n2364_n2088# 0.01512f
C404 source.n127 a_n2364_n2088# 0.035737f
C405 source.n128 a_n2364_n2088# 0.016009f
C406 source.n129 a_n2364_n2088# 0.120406f
C407 source.t13 a_n2364_n2088# 0.058247f
C408 source.n130 a_n2364_n2088# 0.026803f
C409 source.n131 a_n2364_n2088# 0.02111f
C410 source.n132 a_n2364_n2088# 0.01512f
C411 source.n133 a_n2364_n2088# 0.669491f
C412 source.n134 a_n2364_n2088# 0.028137f
C413 source.n135 a_n2364_n2088# 0.01512f
C414 source.n136 a_n2364_n2088# 0.016009f
C415 source.n137 a_n2364_n2088# 0.035737f
C416 source.n138 a_n2364_n2088# 0.035737f
C417 source.n139 a_n2364_n2088# 0.016009f
C418 source.n140 a_n2364_n2088# 0.01512f
C419 source.n141 a_n2364_n2088# 0.028137f
C420 source.n142 a_n2364_n2088# 0.028137f
C421 source.n143 a_n2364_n2088# 0.01512f
C422 source.n144 a_n2364_n2088# 0.016009f
C423 source.n145 a_n2364_n2088# 0.035737f
C424 source.n146 a_n2364_n2088# 0.077365f
C425 source.n147 a_n2364_n2088# 0.016009f
C426 source.n148 a_n2364_n2088# 0.01512f
C427 source.n149 a_n2364_n2088# 0.065037f
C428 source.n150 a_n2364_n2088# 0.043289f
C429 source.n151 a_n2364_n2088# 0.330668f
C430 source.n152 a_n2364_n2088# 1.16689f
C431 plus.n0 a_n2364_n2088# 0.042879f
C432 plus.t0 a_n2364_n2088# 0.522362f
C433 plus.t10 a_n2364_n2088# 0.522362f
C434 plus.n1 a_n2364_n2088# 0.042879f
C435 plus.t4 a_n2364_n2088# 0.522362f
C436 plus.n2 a_n2364_n2088# 0.241378f
C437 plus.n3 a_n2364_n2088# 0.042879f
C438 plus.t9 a_n2364_n2088# 0.522362f
C439 plus.t2 a_n2364_n2088# 0.522362f
C440 plus.n4 a_n2364_n2088# 0.241378f
C441 plus.t5 a_n2364_n2088# 0.542454f
C442 plus.n5 a_n2364_n2088# 0.225013f
C443 plus.t11 a_n2364_n2088# 0.522362f
C444 plus.n6 a_n2364_n2088# 0.24669f
C445 plus.n7 a_n2364_n2088# 0.00973f
C446 plus.n8 a_n2364_n2088# 0.180667f
C447 plus.n9 a_n2364_n2088# 0.042879f
C448 plus.n10 a_n2364_n2088# 0.042879f
C449 plus.n11 a_n2364_n2088# 0.00973f
C450 plus.n12 a_n2364_n2088# 0.241378f
C451 plus.n13 a_n2364_n2088# 0.00973f
C452 plus.n14 a_n2364_n2088# 0.042879f
C453 plus.n15 a_n2364_n2088# 0.042879f
C454 plus.n16 a_n2364_n2088# 0.042879f
C455 plus.n17 a_n2364_n2088# 0.00973f
C456 plus.n18 a_n2364_n2088# 0.241378f
C457 plus.n19 a_n2364_n2088# 0.00973f
C458 plus.n20 a_n2364_n2088# 0.239792f
C459 plus.n21 a_n2364_n2088# 0.383163f
C460 plus.n22 a_n2364_n2088# 0.042879f
C461 plus.t13 a_n2364_n2088# 0.522362f
C462 plus.n23 a_n2364_n2088# 0.042879f
C463 plus.t12 a_n2364_n2088# 0.522362f
C464 plus.t3 a_n2364_n2088# 0.522362f
C465 plus.n24 a_n2364_n2088# 0.241378f
C466 plus.n25 a_n2364_n2088# 0.042879f
C467 plus.t1 a_n2364_n2088# 0.522362f
C468 plus.t6 a_n2364_n2088# 0.522362f
C469 plus.n26 a_n2364_n2088# 0.241378f
C470 plus.t7 a_n2364_n2088# 0.542454f
C471 plus.n27 a_n2364_n2088# 0.225013f
C472 plus.t8 a_n2364_n2088# 0.522362f
C473 plus.n28 a_n2364_n2088# 0.24669f
C474 plus.n29 a_n2364_n2088# 0.00973f
C475 plus.n30 a_n2364_n2088# 0.180667f
C476 plus.n31 a_n2364_n2088# 0.042879f
C477 plus.n32 a_n2364_n2088# 0.042879f
C478 plus.n33 a_n2364_n2088# 0.00973f
C479 plus.n34 a_n2364_n2088# 0.241378f
C480 plus.n35 a_n2364_n2088# 0.00973f
C481 plus.n36 a_n2364_n2088# 0.042879f
C482 plus.n37 a_n2364_n2088# 0.042879f
C483 plus.n38 a_n2364_n2088# 0.042879f
C484 plus.n39 a_n2364_n2088# 0.00973f
C485 plus.n40 a_n2364_n2088# 0.241378f
C486 plus.n41 a_n2364_n2088# 0.00973f
C487 plus.n42 a_n2364_n2088# 0.239792f
C488 plus.n43 a_n2364_n2088# 1.22805f
.ends

