* NGSPICE file created from diffpair137.ext - technology: sky130A

.subckt diffpair137 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t26 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X1 source.t27 plus.t1 drain_left.t14 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X2 source.t6 minus.t0 drain_right.t15 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X3 drain_left.t13 plus.t2 source.t19 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X4 source.t7 minus.t1 drain_right.t14 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t28 plus.t3 drain_left.t12 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right.t13 minus.t2 source.t9 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 drain_right.t12 minus.t3 source.t5 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X8 drain_right.t11 minus.t4 source.t15 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_right.t10 minus.t5 source.t2 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X10 source.t1 minus.t6 drain_right.t9 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X11 source.t31 plus.t4 drain_left.t11 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X12 a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X13 source.t3 minus.t7 drain_right.t8 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 drain_left.t10 plus.t5 source.t24 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 drain_left.t9 plus.t6 source.t21 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 source.t16 plus.t7 drain_left.t8 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 source.t22 plus.t8 drain_left.t7 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X18 source.t4 minus.t8 drain_right.t7 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 drain_right.t6 minus.t9 source.t8 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X20 a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X21 drain_left.t6 plus.t9 source.t18 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X22 source.t10 minus.t10 drain_right.t5 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X23 source.t17 plus.t10 drain_left.t5 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X24 drain_right.t4 minus.t11 source.t0 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X25 a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X26 drain_right.t3 minus.t12 source.t13 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X27 source.t11 minus.t13 drain_right.t2 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X28 drain_left.t4 plus.t11 source.t20 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X29 source.t23 plus.t12 drain_left.t3 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X30 a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X31 source.t12 minus.t14 drain_right.t1 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X32 source.t30 plus.t13 drain_left.t2 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X33 drain_right.t0 minus.t15 source.t14 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X34 drain_left.t1 plus.t14 source.t29 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X35 drain_left.t0 plus.t15 source.t25 a_n2390_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
R0 plus.n6 plus.t12 166.787
R1 plus.n30 plus.t14 166.787
R2 plus.n8 plus.n7 161.3
R3 plus.n9 plus.n4 161.3
R4 plus.n11 plus.n10 161.3
R5 plus.n12 plus.n3 161.3
R6 plus.n14 plus.n13 161.3
R7 plus.n15 plus.n2 161.3
R8 plus.n17 plus.n16 161.3
R9 plus.n18 plus.n1 161.3
R10 plus.n20 plus.n19 161.3
R11 plus.n21 plus.n0 161.3
R12 plus.n23 plus.n22 161.3
R13 plus.n32 plus.n31 161.3
R14 plus.n33 plus.n28 161.3
R15 plus.n35 plus.n34 161.3
R16 plus.n36 plus.n27 161.3
R17 plus.n38 plus.n37 161.3
R18 plus.n39 plus.n26 161.3
R19 plus.n41 plus.n40 161.3
R20 plus.n42 plus.n25 161.3
R21 plus.n44 plus.n43 161.3
R22 plus.n45 plus.n24 161.3
R23 plus.n47 plus.n46 161.3
R24 plus.n22 plus.t0 145.805
R25 plus.n21 plus.t1 145.805
R26 plus.n1 plus.t2 145.805
R27 plus.n15 plus.t7 145.805
R28 plus.n3 plus.t9 145.805
R29 plus.n9 plus.t10 145.805
R30 plus.n5 plus.t11 145.805
R31 plus.n46 plus.t4 145.805
R32 plus.n45 plus.t6 145.805
R33 plus.n25 plus.t13 145.805
R34 plus.n39 plus.t15 145.805
R35 plus.n27 plus.t3 145.805
R36 plus.n33 plus.t5 145.805
R37 plus.n29 plus.t8 145.805
R38 plus.n7 plus.n6 70.4033
R39 plus.n31 plus.n30 70.4033
R40 plus.n22 plus.n21 48.2005
R41 plus.n46 plus.n45 48.2005
R42 plus.n20 plus.n1 44.549
R43 plus.n9 plus.n8 44.549
R44 plus.n44 plus.n25 44.549
R45 plus.n33 plus.n32 44.549
R46 plus.n16 plus.n15 34.3247
R47 plus.n10 plus.n3 34.3247
R48 plus.n40 plus.n39 34.3247
R49 plus.n34 plus.n27 34.3247
R50 plus plus.n47 28.4233
R51 plus.n14 plus.n3 24.1005
R52 plus.n15 plus.n14 24.1005
R53 plus.n39 plus.n38 24.1005
R54 plus.n38 plus.n27 24.1005
R55 plus.n6 plus.n5 20.9576
R56 plus.n30 plus.n29 20.9576
R57 plus.n16 plus.n1 13.8763
R58 plus.n10 plus.n9 13.8763
R59 plus.n40 plus.n25 13.8763
R60 plus.n34 plus.n33 13.8763
R61 plus plus.n23 8.51186
R62 plus.n21 plus.n20 3.65202
R63 plus.n8 plus.n5 3.65202
R64 plus.n45 plus.n44 3.65202
R65 plus.n32 plus.n29 3.65202
R66 plus.n7 plus.n4 0.189894
R67 plus.n11 plus.n4 0.189894
R68 plus.n12 plus.n11 0.189894
R69 plus.n13 plus.n12 0.189894
R70 plus.n13 plus.n2 0.189894
R71 plus.n17 plus.n2 0.189894
R72 plus.n18 plus.n17 0.189894
R73 plus.n19 plus.n18 0.189894
R74 plus.n19 plus.n0 0.189894
R75 plus.n23 plus.n0 0.189894
R76 plus.n47 plus.n24 0.189894
R77 plus.n43 plus.n24 0.189894
R78 plus.n43 plus.n42 0.189894
R79 plus.n42 plus.n41 0.189894
R80 plus.n41 plus.n26 0.189894
R81 plus.n37 plus.n26 0.189894
R82 plus.n37 plus.n36 0.189894
R83 plus.n36 plus.n35 0.189894
R84 plus.n35 plus.n28 0.189894
R85 plus.n31 plus.n28 0.189894
R86 source.n82 source.n80 289.615
R87 source.n68 source.n66 289.615
R88 source.n60 source.n58 289.615
R89 source.n46 source.n44 289.615
R90 source.n2 source.n0 289.615
R91 source.n16 source.n14 289.615
R92 source.n24 source.n22 289.615
R93 source.n38 source.n36 289.615
R94 source.n83 source.n82 185
R95 source.n69 source.n68 185
R96 source.n61 source.n60 185
R97 source.n47 source.n46 185
R98 source.n3 source.n2 185
R99 source.n17 source.n16 185
R100 source.n25 source.n24 185
R101 source.n39 source.n38 185
R102 source.t13 source.n81 167.117
R103 source.t1 source.n67 167.117
R104 source.t29 source.n59 167.117
R105 source.t31 source.n45 167.117
R106 source.t26 source.n1 167.117
R107 source.t23 source.n15 167.117
R108 source.t0 source.n23 167.117
R109 source.t7 source.n37 167.117
R110 source.n9 source.n8 84.1169
R111 source.n11 source.n10 84.1169
R112 source.n13 source.n12 84.1169
R113 source.n31 source.n30 84.1169
R114 source.n33 source.n32 84.1169
R115 source.n35 source.n34 84.1169
R116 source.n79 source.n78 84.1168
R117 source.n77 source.n76 84.1168
R118 source.n75 source.n74 84.1168
R119 source.n57 source.n56 84.1168
R120 source.n55 source.n54 84.1168
R121 source.n53 source.n52 84.1168
R122 source.n82 source.t13 52.3082
R123 source.n68 source.t1 52.3082
R124 source.n60 source.t29 52.3082
R125 source.n46 source.t31 52.3082
R126 source.n2 source.t26 52.3082
R127 source.n16 source.t23 52.3082
R128 source.n24 source.t0 52.3082
R129 source.n38 source.t7 52.3082
R130 source.n87 source.n86 31.4096
R131 source.n73 source.n72 31.4096
R132 source.n65 source.n64 31.4096
R133 source.n51 source.n50 31.4096
R134 source.n7 source.n6 31.4096
R135 source.n21 source.n20 31.4096
R136 source.n29 source.n28 31.4096
R137 source.n43 source.n42 31.4096
R138 source.n51 source.n43 14.5137
R139 source.n78 source.t9 9.9005
R140 source.n78 source.t12 9.9005
R141 source.n76 source.t2 9.9005
R142 source.n76 source.t6 9.9005
R143 source.n74 source.t14 9.9005
R144 source.n74 source.t11 9.9005
R145 source.n56 source.t24 9.9005
R146 source.n56 source.t22 9.9005
R147 source.n54 source.t25 9.9005
R148 source.n54 source.t28 9.9005
R149 source.n52 source.t21 9.9005
R150 source.n52 source.t30 9.9005
R151 source.n8 source.t19 9.9005
R152 source.n8 source.t27 9.9005
R153 source.n10 source.t18 9.9005
R154 source.n10 source.t16 9.9005
R155 source.n12 source.t20 9.9005
R156 source.n12 source.t17 9.9005
R157 source.n30 source.t8 9.9005
R158 source.n30 source.t10 9.9005
R159 source.n32 source.t5 9.9005
R160 source.n32 source.t4 9.9005
R161 source.n34 source.t15 9.9005
R162 source.n34 source.t3 9.9005
R163 source.n83 source.n81 9.71174
R164 source.n69 source.n67 9.71174
R165 source.n61 source.n59 9.71174
R166 source.n47 source.n45 9.71174
R167 source.n3 source.n1 9.71174
R168 source.n17 source.n15 9.71174
R169 source.n25 source.n23 9.71174
R170 source.n39 source.n37 9.71174
R171 source.n86 source.n85 9.45567
R172 source.n72 source.n71 9.45567
R173 source.n64 source.n63 9.45567
R174 source.n50 source.n49 9.45567
R175 source.n6 source.n5 9.45567
R176 source.n20 source.n19 9.45567
R177 source.n28 source.n27 9.45567
R178 source.n42 source.n41 9.45567
R179 source.n85 source.n84 9.3005
R180 source.n71 source.n70 9.3005
R181 source.n63 source.n62 9.3005
R182 source.n49 source.n48 9.3005
R183 source.n5 source.n4 9.3005
R184 source.n19 source.n18 9.3005
R185 source.n27 source.n26 9.3005
R186 source.n41 source.n40 9.3005
R187 source.n88 source.n7 8.8499
R188 source.n86 source.n80 8.14595
R189 source.n72 source.n66 8.14595
R190 source.n64 source.n58 8.14595
R191 source.n50 source.n44 8.14595
R192 source.n6 source.n0 8.14595
R193 source.n20 source.n14 8.14595
R194 source.n28 source.n22 8.14595
R195 source.n42 source.n36 8.14595
R196 source.n84 source.n83 7.3702
R197 source.n70 source.n69 7.3702
R198 source.n62 source.n61 7.3702
R199 source.n48 source.n47 7.3702
R200 source.n4 source.n3 7.3702
R201 source.n18 source.n17 7.3702
R202 source.n26 source.n25 7.3702
R203 source.n40 source.n39 7.3702
R204 source.n84 source.n80 5.81868
R205 source.n70 source.n66 5.81868
R206 source.n62 source.n58 5.81868
R207 source.n48 source.n44 5.81868
R208 source.n4 source.n0 5.81868
R209 source.n18 source.n14 5.81868
R210 source.n26 source.n22 5.81868
R211 source.n40 source.n36 5.81868
R212 source.n88 source.n87 5.66429
R213 source.n85 source.n81 3.44771
R214 source.n71 source.n67 3.44771
R215 source.n63 source.n59 3.44771
R216 source.n49 source.n45 3.44771
R217 source.n5 source.n1 3.44771
R218 source.n19 source.n15 3.44771
R219 source.n27 source.n23 3.44771
R220 source.n41 source.n37 3.44771
R221 source.n43 source.n35 0.802224
R222 source.n35 source.n33 0.802224
R223 source.n33 source.n31 0.802224
R224 source.n31 source.n29 0.802224
R225 source.n21 source.n13 0.802224
R226 source.n13 source.n11 0.802224
R227 source.n11 source.n9 0.802224
R228 source.n9 source.n7 0.802224
R229 source.n53 source.n51 0.802224
R230 source.n55 source.n53 0.802224
R231 source.n57 source.n55 0.802224
R232 source.n65 source.n57 0.802224
R233 source.n75 source.n73 0.802224
R234 source.n77 source.n75 0.802224
R235 source.n79 source.n77 0.802224
R236 source.n87 source.n79 0.802224
R237 source.n29 source.n21 0.470328
R238 source.n73 source.n65 0.470328
R239 source source.n88 0.188
R240 drain_left.n9 drain_left.n7 101.597
R241 drain_left.n5 drain_left.n3 101.597
R242 drain_left.n2 drain_left.n0 101.597
R243 drain_left.n13 drain_left.n12 100.796
R244 drain_left.n11 drain_left.n10 100.796
R245 drain_left.n9 drain_left.n8 100.796
R246 drain_left.n5 drain_left.n4 100.796
R247 drain_left.n2 drain_left.n1 100.796
R248 drain_left drain_left.n6 25.0025
R249 drain_left.n3 drain_left.t7 9.9005
R250 drain_left.n3 drain_left.t1 9.9005
R251 drain_left.n4 drain_left.t12 9.9005
R252 drain_left.n4 drain_left.t10 9.9005
R253 drain_left.n1 drain_left.t2 9.9005
R254 drain_left.n1 drain_left.t0 9.9005
R255 drain_left.n0 drain_left.t11 9.9005
R256 drain_left.n0 drain_left.t9 9.9005
R257 drain_left.n12 drain_left.t14 9.9005
R258 drain_left.n12 drain_left.t15 9.9005
R259 drain_left.n10 drain_left.t8 9.9005
R260 drain_left.n10 drain_left.t13 9.9005
R261 drain_left.n8 drain_left.t5 9.9005
R262 drain_left.n8 drain_left.t6 9.9005
R263 drain_left.n7 drain_left.t3 9.9005
R264 drain_left.n7 drain_left.t4 9.9005
R265 drain_left drain_left.n13 6.45494
R266 drain_left.n11 drain_left.n9 0.802224
R267 drain_left.n13 drain_left.n11 0.802224
R268 drain_left.n6 drain_left.n5 0.346016
R269 drain_left.n6 drain_left.n2 0.346016
R270 minus.n6 minus.t11 166.787
R271 minus.n30 minus.t6 166.787
R272 minus.n23 minus.n22 161.3
R273 minus.n21 minus.n0 161.3
R274 minus.n20 minus.n19 161.3
R275 minus.n18 minus.n1 161.3
R276 minus.n17 minus.n16 161.3
R277 minus.n15 minus.n2 161.3
R278 minus.n14 minus.n13 161.3
R279 minus.n12 minus.n3 161.3
R280 minus.n11 minus.n10 161.3
R281 minus.n9 minus.n4 161.3
R282 minus.n8 minus.n7 161.3
R283 minus.n47 minus.n46 161.3
R284 minus.n45 minus.n24 161.3
R285 minus.n44 minus.n43 161.3
R286 minus.n42 minus.n25 161.3
R287 minus.n41 minus.n40 161.3
R288 minus.n39 minus.n26 161.3
R289 minus.n38 minus.n37 161.3
R290 minus.n36 minus.n27 161.3
R291 minus.n35 minus.n34 161.3
R292 minus.n33 minus.n28 161.3
R293 minus.n32 minus.n31 161.3
R294 minus.n5 minus.t10 145.805
R295 minus.n9 minus.t9 145.805
R296 minus.n3 minus.t8 145.805
R297 minus.n15 minus.t3 145.805
R298 minus.n1 minus.t7 145.805
R299 minus.n21 minus.t4 145.805
R300 minus.n22 minus.t1 145.805
R301 minus.n29 minus.t15 145.805
R302 minus.n33 minus.t13 145.805
R303 minus.n27 minus.t5 145.805
R304 minus.n39 minus.t0 145.805
R305 minus.n25 minus.t2 145.805
R306 minus.n45 minus.t14 145.805
R307 minus.n46 minus.t12 145.805
R308 minus.n7 minus.n6 70.4033
R309 minus.n31 minus.n30 70.4033
R310 minus.n22 minus.n21 48.2005
R311 minus.n46 minus.n45 48.2005
R312 minus.n9 minus.n8 44.549
R313 minus.n20 minus.n1 44.549
R314 minus.n33 minus.n32 44.549
R315 minus.n44 minus.n25 44.549
R316 minus.n10 minus.n3 34.3247
R317 minus.n16 minus.n15 34.3247
R318 minus.n34 minus.n27 34.3247
R319 minus.n40 minus.n39 34.3247
R320 minus.n48 minus.n23 30.7543
R321 minus.n15 minus.n14 24.1005
R322 minus.n14 minus.n3 24.1005
R323 minus.n38 minus.n27 24.1005
R324 minus.n39 minus.n38 24.1005
R325 minus.n6 minus.n5 20.9576
R326 minus.n30 minus.n29 20.9576
R327 minus.n10 minus.n9 13.8763
R328 minus.n16 minus.n1 13.8763
R329 minus.n34 minus.n33 13.8763
R330 minus.n40 minus.n25 13.8763
R331 minus.n48 minus.n47 6.6558
R332 minus.n8 minus.n5 3.65202
R333 minus.n21 minus.n20 3.65202
R334 minus.n32 minus.n29 3.65202
R335 minus.n45 minus.n44 3.65202
R336 minus.n23 minus.n0 0.189894
R337 minus.n19 minus.n0 0.189894
R338 minus.n19 minus.n18 0.189894
R339 minus.n18 minus.n17 0.189894
R340 minus.n17 minus.n2 0.189894
R341 minus.n13 minus.n2 0.189894
R342 minus.n13 minus.n12 0.189894
R343 minus.n12 minus.n11 0.189894
R344 minus.n11 minus.n4 0.189894
R345 minus.n7 minus.n4 0.189894
R346 minus.n31 minus.n28 0.189894
R347 minus.n35 minus.n28 0.189894
R348 minus.n36 minus.n35 0.189894
R349 minus.n37 minus.n36 0.189894
R350 minus.n37 minus.n26 0.189894
R351 minus.n41 minus.n26 0.189894
R352 minus.n42 minus.n41 0.189894
R353 minus.n43 minus.n42 0.189894
R354 minus.n43 minus.n24 0.189894
R355 minus.n47 minus.n24 0.189894
R356 minus minus.n48 0.188
R357 drain_right.n9 drain_right.n7 101.597
R358 drain_right.n5 drain_right.n3 101.597
R359 drain_right.n2 drain_right.n0 101.597
R360 drain_right.n9 drain_right.n8 100.796
R361 drain_right.n11 drain_right.n10 100.796
R362 drain_right.n13 drain_right.n12 100.796
R363 drain_right.n5 drain_right.n4 100.796
R364 drain_right.n2 drain_right.n1 100.796
R365 drain_right drain_right.n6 24.4493
R366 drain_right.n3 drain_right.t1 9.9005
R367 drain_right.n3 drain_right.t3 9.9005
R368 drain_right.n4 drain_right.t15 9.9005
R369 drain_right.n4 drain_right.t13 9.9005
R370 drain_right.n1 drain_right.t2 9.9005
R371 drain_right.n1 drain_right.t10 9.9005
R372 drain_right.n0 drain_right.t9 9.9005
R373 drain_right.n0 drain_right.t0 9.9005
R374 drain_right.n7 drain_right.t5 9.9005
R375 drain_right.n7 drain_right.t4 9.9005
R376 drain_right.n8 drain_right.t7 9.9005
R377 drain_right.n8 drain_right.t6 9.9005
R378 drain_right.n10 drain_right.t8 9.9005
R379 drain_right.n10 drain_right.t12 9.9005
R380 drain_right.n12 drain_right.t14 9.9005
R381 drain_right.n12 drain_right.t11 9.9005
R382 drain_right drain_right.n13 6.45494
R383 drain_right.n13 drain_right.n11 0.802224
R384 drain_right.n11 drain_right.n9 0.802224
R385 drain_right.n6 drain_right.n5 0.346016
R386 drain_right.n6 drain_right.n2 0.346016
C0 drain_right drain_left 1.24373f
C1 drain_right source 6.3097f
C2 drain_right minus 2.03603f
C3 drain_right plus 0.398723f
C4 source drain_left 6.30798f
C5 minus drain_left 0.178671f
C6 minus source 2.53086f
C7 plus drain_left 2.27185f
C8 plus source 2.54483f
C9 plus minus 4.28028f
C10 drain_right a_n2390_n1288# 4.63672f
C11 drain_left a_n2390_n1288# 5.00929f
C12 source a_n2390_n1288# 3.311003f
C13 minus a_n2390_n1288# 8.664556f
C14 plus a_n2390_n1288# 9.96924f
C15 drain_right.t9 a_n2390_n1288# 0.042715f
C16 drain_right.t0 a_n2390_n1288# 0.042715f
C17 drain_right.n0 a_n2390_n1288# 0.27117f
C18 drain_right.t2 a_n2390_n1288# 0.042715f
C19 drain_right.t10 a_n2390_n1288# 0.042715f
C20 drain_right.n1 a_n2390_n1288# 0.26835f
C21 drain_right.n2 a_n2390_n1288# 0.663154f
C22 drain_right.t1 a_n2390_n1288# 0.042715f
C23 drain_right.t3 a_n2390_n1288# 0.042715f
C24 drain_right.n3 a_n2390_n1288# 0.27117f
C25 drain_right.t15 a_n2390_n1288# 0.042715f
C26 drain_right.t13 a_n2390_n1288# 0.042715f
C27 drain_right.n4 a_n2390_n1288# 0.26835f
C28 drain_right.n5 a_n2390_n1288# 0.663155f
C29 drain_right.n6 a_n2390_n1288# 0.882924f
C30 drain_right.t5 a_n2390_n1288# 0.042715f
C31 drain_right.t4 a_n2390_n1288# 0.042715f
C32 drain_right.n7 a_n2390_n1288# 0.271171f
C33 drain_right.t7 a_n2390_n1288# 0.042715f
C34 drain_right.t6 a_n2390_n1288# 0.042715f
C35 drain_right.n8 a_n2390_n1288# 0.268351f
C36 drain_right.n9 a_n2390_n1288# 0.701069f
C37 drain_right.t8 a_n2390_n1288# 0.042715f
C38 drain_right.t12 a_n2390_n1288# 0.042715f
C39 drain_right.n10 a_n2390_n1288# 0.268351f
C40 drain_right.n11 a_n2390_n1288# 0.346501f
C41 drain_right.t14 a_n2390_n1288# 0.042715f
C42 drain_right.t11 a_n2390_n1288# 0.042715f
C43 drain_right.n12 a_n2390_n1288# 0.268351f
C44 drain_right.n13 a_n2390_n1288# 0.582175f
C45 minus.n0 a_n2390_n1288# 0.044613f
C46 minus.t7 a_n2390_n1288# 0.165784f
C47 minus.n1 a_n2390_n1288# 0.119321f
C48 minus.n2 a_n2390_n1288# 0.044613f
C49 minus.t8 a_n2390_n1288# 0.165784f
C50 minus.n3 a_n2390_n1288# 0.119321f
C51 minus.n4 a_n2390_n1288# 0.044613f
C52 minus.t10 a_n2390_n1288# 0.165784f
C53 minus.n5 a_n2390_n1288# 0.118083f
C54 minus.t11 a_n2390_n1288# 0.180562f
C55 minus.n6 a_n2390_n1288# 0.102975f
C56 minus.n7 a_n2390_n1288# 0.15026f
C57 minus.n8 a_n2390_n1288# 0.010124f
C58 minus.t9 a_n2390_n1288# 0.165784f
C59 minus.n9 a_n2390_n1288# 0.119321f
C60 minus.n10 a_n2390_n1288# 0.010124f
C61 minus.n11 a_n2390_n1288# 0.044613f
C62 minus.n12 a_n2390_n1288# 0.044613f
C63 minus.n13 a_n2390_n1288# 0.044613f
C64 minus.n14 a_n2390_n1288# 0.010124f
C65 minus.t3 a_n2390_n1288# 0.165784f
C66 minus.n15 a_n2390_n1288# 0.119321f
C67 minus.n16 a_n2390_n1288# 0.010124f
C68 minus.n17 a_n2390_n1288# 0.044613f
C69 minus.n18 a_n2390_n1288# 0.044613f
C70 minus.n19 a_n2390_n1288# 0.044613f
C71 minus.n20 a_n2390_n1288# 0.010124f
C72 minus.t4 a_n2390_n1288# 0.165784f
C73 minus.n21 a_n2390_n1288# 0.118083f
C74 minus.t1 a_n2390_n1288# 0.165784f
C75 minus.n22 a_n2390_n1288# 0.117396f
C76 minus.n23 a_n2390_n1288# 1.21682f
C77 minus.n24 a_n2390_n1288# 0.044613f
C78 minus.t2 a_n2390_n1288# 0.165784f
C79 minus.n25 a_n2390_n1288# 0.119321f
C80 minus.n26 a_n2390_n1288# 0.044613f
C81 minus.t5 a_n2390_n1288# 0.165784f
C82 minus.n27 a_n2390_n1288# 0.119321f
C83 minus.n28 a_n2390_n1288# 0.044613f
C84 minus.t15 a_n2390_n1288# 0.165784f
C85 minus.n29 a_n2390_n1288# 0.118083f
C86 minus.t6 a_n2390_n1288# 0.180562f
C87 minus.n30 a_n2390_n1288# 0.102975f
C88 minus.n31 a_n2390_n1288# 0.15026f
C89 minus.n32 a_n2390_n1288# 0.010124f
C90 minus.t13 a_n2390_n1288# 0.165784f
C91 minus.n33 a_n2390_n1288# 0.119321f
C92 minus.n34 a_n2390_n1288# 0.010124f
C93 minus.n35 a_n2390_n1288# 0.044613f
C94 minus.n36 a_n2390_n1288# 0.044613f
C95 minus.n37 a_n2390_n1288# 0.044613f
C96 minus.n38 a_n2390_n1288# 0.010124f
C97 minus.t0 a_n2390_n1288# 0.165784f
C98 minus.n39 a_n2390_n1288# 0.119321f
C99 minus.n40 a_n2390_n1288# 0.010124f
C100 minus.n41 a_n2390_n1288# 0.044613f
C101 minus.n42 a_n2390_n1288# 0.044613f
C102 minus.n43 a_n2390_n1288# 0.044613f
C103 minus.n44 a_n2390_n1288# 0.010124f
C104 minus.t14 a_n2390_n1288# 0.165784f
C105 minus.n45 a_n2390_n1288# 0.118083f
C106 minus.t12 a_n2390_n1288# 0.165784f
C107 minus.n46 a_n2390_n1288# 0.117396f
C108 minus.n47 a_n2390_n1288# 0.307924f
C109 minus.n48 a_n2390_n1288# 1.49143f
C110 drain_left.t11 a_n2390_n1288# 0.043702f
C111 drain_left.t9 a_n2390_n1288# 0.043702f
C112 drain_left.n0 a_n2390_n1288# 0.277438f
C113 drain_left.t2 a_n2390_n1288# 0.043702f
C114 drain_left.t0 a_n2390_n1288# 0.043702f
C115 drain_left.n1 a_n2390_n1288# 0.274552f
C116 drain_left.n2 a_n2390_n1288# 0.678481f
C117 drain_left.t7 a_n2390_n1288# 0.043702f
C118 drain_left.t1 a_n2390_n1288# 0.043702f
C119 drain_left.n3 a_n2390_n1288# 0.277438f
C120 drain_left.t12 a_n2390_n1288# 0.043702f
C121 drain_left.t10 a_n2390_n1288# 0.043702f
C122 drain_left.n4 a_n2390_n1288# 0.274552f
C123 drain_left.n5 a_n2390_n1288# 0.678481f
C124 drain_left.n6 a_n2390_n1288# 0.957218f
C125 drain_left.t3 a_n2390_n1288# 0.043702f
C126 drain_left.t4 a_n2390_n1288# 0.043702f
C127 drain_left.n7 a_n2390_n1288# 0.277439f
C128 drain_left.t5 a_n2390_n1288# 0.043702f
C129 drain_left.t6 a_n2390_n1288# 0.043702f
C130 drain_left.n8 a_n2390_n1288# 0.274553f
C131 drain_left.n9 a_n2390_n1288# 0.717272f
C132 drain_left.t8 a_n2390_n1288# 0.043702f
C133 drain_left.t13 a_n2390_n1288# 0.043702f
C134 drain_left.n10 a_n2390_n1288# 0.274553f
C135 drain_left.n11 a_n2390_n1288# 0.35451f
C136 drain_left.t14 a_n2390_n1288# 0.043702f
C137 drain_left.t15 a_n2390_n1288# 0.043702f
C138 drain_left.n12 a_n2390_n1288# 0.274553f
C139 drain_left.n13 a_n2390_n1288# 0.59563f
C140 source.n0 a_n2390_n1288# 0.044387f
C141 source.n1 a_n2390_n1288# 0.098213f
C142 source.t26 a_n2390_n1288# 0.073703f
C143 source.n2 a_n2390_n1288# 0.076865f
C144 source.n3 a_n2390_n1288# 0.024778f
C145 source.n4 a_n2390_n1288# 0.016342f
C146 source.n5 a_n2390_n1288# 0.216484f
C147 source.n6 a_n2390_n1288# 0.048659f
C148 source.n7 a_n2390_n1288# 0.504098f
C149 source.t19 a_n2390_n1288# 0.048064f
C150 source.t27 a_n2390_n1288# 0.048064f
C151 source.n8 a_n2390_n1288# 0.256949f
C152 source.n9 a_n2390_n1288# 0.393561f
C153 source.t18 a_n2390_n1288# 0.048064f
C154 source.t16 a_n2390_n1288# 0.048064f
C155 source.n10 a_n2390_n1288# 0.256949f
C156 source.n11 a_n2390_n1288# 0.393561f
C157 source.t20 a_n2390_n1288# 0.048064f
C158 source.t17 a_n2390_n1288# 0.048064f
C159 source.n12 a_n2390_n1288# 0.256949f
C160 source.n13 a_n2390_n1288# 0.393561f
C161 source.n14 a_n2390_n1288# 0.044387f
C162 source.n15 a_n2390_n1288# 0.098213f
C163 source.t23 a_n2390_n1288# 0.073703f
C164 source.n16 a_n2390_n1288# 0.076865f
C165 source.n17 a_n2390_n1288# 0.024778f
C166 source.n18 a_n2390_n1288# 0.016342f
C167 source.n19 a_n2390_n1288# 0.216484f
C168 source.n20 a_n2390_n1288# 0.048659f
C169 source.n21 a_n2390_n1288# 0.149638f
C170 source.n22 a_n2390_n1288# 0.044387f
C171 source.n23 a_n2390_n1288# 0.098213f
C172 source.t0 a_n2390_n1288# 0.073703f
C173 source.n24 a_n2390_n1288# 0.076865f
C174 source.n25 a_n2390_n1288# 0.024778f
C175 source.n26 a_n2390_n1288# 0.016342f
C176 source.n27 a_n2390_n1288# 0.216484f
C177 source.n28 a_n2390_n1288# 0.048659f
C178 source.n29 a_n2390_n1288# 0.149638f
C179 source.t8 a_n2390_n1288# 0.048064f
C180 source.t10 a_n2390_n1288# 0.048064f
C181 source.n30 a_n2390_n1288# 0.256949f
C182 source.n31 a_n2390_n1288# 0.393561f
C183 source.t5 a_n2390_n1288# 0.048064f
C184 source.t4 a_n2390_n1288# 0.048064f
C185 source.n32 a_n2390_n1288# 0.256949f
C186 source.n33 a_n2390_n1288# 0.393561f
C187 source.t15 a_n2390_n1288# 0.048064f
C188 source.t3 a_n2390_n1288# 0.048064f
C189 source.n34 a_n2390_n1288# 0.256949f
C190 source.n35 a_n2390_n1288# 0.393561f
C191 source.n36 a_n2390_n1288# 0.044387f
C192 source.n37 a_n2390_n1288# 0.098213f
C193 source.t7 a_n2390_n1288# 0.073703f
C194 source.n38 a_n2390_n1288# 0.076865f
C195 source.n39 a_n2390_n1288# 0.024778f
C196 source.n40 a_n2390_n1288# 0.016342f
C197 source.n41 a_n2390_n1288# 0.216484f
C198 source.n42 a_n2390_n1288# 0.048659f
C199 source.n43 a_n2390_n1288# 0.793376f
C200 source.n44 a_n2390_n1288# 0.044387f
C201 source.n45 a_n2390_n1288# 0.098213f
C202 source.t31 a_n2390_n1288# 0.073703f
C203 source.n46 a_n2390_n1288# 0.076865f
C204 source.n47 a_n2390_n1288# 0.024778f
C205 source.n48 a_n2390_n1288# 0.016342f
C206 source.n49 a_n2390_n1288# 0.216484f
C207 source.n50 a_n2390_n1288# 0.048659f
C208 source.n51 a_n2390_n1288# 0.793376f
C209 source.t21 a_n2390_n1288# 0.048064f
C210 source.t30 a_n2390_n1288# 0.048064f
C211 source.n52 a_n2390_n1288# 0.256948f
C212 source.n53 a_n2390_n1288# 0.393562f
C213 source.t25 a_n2390_n1288# 0.048064f
C214 source.t28 a_n2390_n1288# 0.048064f
C215 source.n54 a_n2390_n1288# 0.256948f
C216 source.n55 a_n2390_n1288# 0.393562f
C217 source.t24 a_n2390_n1288# 0.048064f
C218 source.t22 a_n2390_n1288# 0.048064f
C219 source.n56 a_n2390_n1288# 0.256948f
C220 source.n57 a_n2390_n1288# 0.393562f
C221 source.n58 a_n2390_n1288# 0.044387f
C222 source.n59 a_n2390_n1288# 0.098213f
C223 source.t29 a_n2390_n1288# 0.073703f
C224 source.n60 a_n2390_n1288# 0.076865f
C225 source.n61 a_n2390_n1288# 0.024778f
C226 source.n62 a_n2390_n1288# 0.016342f
C227 source.n63 a_n2390_n1288# 0.216484f
C228 source.n64 a_n2390_n1288# 0.048659f
C229 source.n65 a_n2390_n1288# 0.149638f
C230 source.n66 a_n2390_n1288# 0.044387f
C231 source.n67 a_n2390_n1288# 0.098213f
C232 source.t1 a_n2390_n1288# 0.073703f
C233 source.n68 a_n2390_n1288# 0.076865f
C234 source.n69 a_n2390_n1288# 0.024778f
C235 source.n70 a_n2390_n1288# 0.016342f
C236 source.n71 a_n2390_n1288# 0.216484f
C237 source.n72 a_n2390_n1288# 0.048659f
C238 source.n73 a_n2390_n1288# 0.149638f
C239 source.t14 a_n2390_n1288# 0.048064f
C240 source.t11 a_n2390_n1288# 0.048064f
C241 source.n74 a_n2390_n1288# 0.256948f
C242 source.n75 a_n2390_n1288# 0.393562f
C243 source.t2 a_n2390_n1288# 0.048064f
C244 source.t6 a_n2390_n1288# 0.048064f
C245 source.n76 a_n2390_n1288# 0.256948f
C246 source.n77 a_n2390_n1288# 0.393562f
C247 source.t9 a_n2390_n1288# 0.048064f
C248 source.t12 a_n2390_n1288# 0.048064f
C249 source.n78 a_n2390_n1288# 0.256948f
C250 source.n79 a_n2390_n1288# 0.393562f
C251 source.n80 a_n2390_n1288# 0.044387f
C252 source.n81 a_n2390_n1288# 0.098213f
C253 source.t13 a_n2390_n1288# 0.073703f
C254 source.n82 a_n2390_n1288# 0.076865f
C255 source.n83 a_n2390_n1288# 0.024778f
C256 source.n84 a_n2390_n1288# 0.016342f
C257 source.n85 a_n2390_n1288# 0.216484f
C258 source.n86 a_n2390_n1288# 0.048659f
C259 source.n87 a_n2390_n1288# 0.341394f
C260 source.n88 a_n2390_n1288# 0.762891f
C261 plus.n0 a_n2390_n1288# 0.046611f
C262 plus.t0 a_n2390_n1288# 0.173212f
C263 plus.t1 a_n2390_n1288# 0.173212f
C264 plus.t2 a_n2390_n1288# 0.173212f
C265 plus.n1 a_n2390_n1288# 0.124667f
C266 plus.n2 a_n2390_n1288# 0.046611f
C267 plus.t7 a_n2390_n1288# 0.173212f
C268 plus.t9 a_n2390_n1288# 0.173212f
C269 plus.n3 a_n2390_n1288# 0.124667f
C270 plus.n4 a_n2390_n1288# 0.046611f
C271 plus.t10 a_n2390_n1288# 0.173212f
C272 plus.t11 a_n2390_n1288# 0.173212f
C273 plus.n5 a_n2390_n1288# 0.123374f
C274 plus.t12 a_n2390_n1288# 0.188651f
C275 plus.n6 a_n2390_n1288# 0.107589f
C276 plus.n7 a_n2390_n1288# 0.156992f
C277 plus.n8 a_n2390_n1288# 0.010577f
C278 plus.n9 a_n2390_n1288# 0.124667f
C279 plus.n10 a_n2390_n1288# 0.010577f
C280 plus.n11 a_n2390_n1288# 0.046611f
C281 plus.n12 a_n2390_n1288# 0.046611f
C282 plus.n13 a_n2390_n1288# 0.046611f
C283 plus.n14 a_n2390_n1288# 0.010577f
C284 plus.n15 a_n2390_n1288# 0.124667f
C285 plus.n16 a_n2390_n1288# 0.010577f
C286 plus.n17 a_n2390_n1288# 0.046611f
C287 plus.n18 a_n2390_n1288# 0.046611f
C288 plus.n19 a_n2390_n1288# 0.046611f
C289 plus.n20 a_n2390_n1288# 0.010577f
C290 plus.n21 a_n2390_n1288# 0.123374f
C291 plus.n22 a_n2390_n1288# 0.122655f
C292 plus.n23 a_n2390_n1288# 0.351136f
C293 plus.n24 a_n2390_n1288# 0.046611f
C294 plus.t4 a_n2390_n1288# 0.173212f
C295 plus.t6 a_n2390_n1288# 0.173212f
C296 plus.t13 a_n2390_n1288# 0.173212f
C297 plus.n25 a_n2390_n1288# 0.124667f
C298 plus.n26 a_n2390_n1288# 0.046611f
C299 plus.t15 a_n2390_n1288# 0.173212f
C300 plus.t3 a_n2390_n1288# 0.173212f
C301 plus.n27 a_n2390_n1288# 0.124667f
C302 plus.n28 a_n2390_n1288# 0.046611f
C303 plus.t5 a_n2390_n1288# 0.173212f
C304 plus.t8 a_n2390_n1288# 0.173212f
C305 plus.n29 a_n2390_n1288# 0.123374f
C306 plus.t14 a_n2390_n1288# 0.188651f
C307 plus.n30 a_n2390_n1288# 0.107589f
C308 plus.n31 a_n2390_n1288# 0.156992f
C309 plus.n32 a_n2390_n1288# 0.010577f
C310 plus.n33 a_n2390_n1288# 0.124667f
C311 plus.n34 a_n2390_n1288# 0.010577f
C312 plus.n35 a_n2390_n1288# 0.046611f
C313 plus.n36 a_n2390_n1288# 0.046611f
C314 plus.n37 a_n2390_n1288# 0.046611f
C315 plus.n38 a_n2390_n1288# 0.010577f
C316 plus.n39 a_n2390_n1288# 0.124667f
C317 plus.n40 a_n2390_n1288# 0.010577f
C318 plus.n41 a_n2390_n1288# 0.046611f
C319 plus.n42 a_n2390_n1288# 0.046611f
C320 plus.n43 a_n2390_n1288# 0.046611f
C321 plus.n44 a_n2390_n1288# 0.010577f
C322 plus.n45 a_n2390_n1288# 0.123374f
C323 plus.n46 a_n2390_n1288# 0.122655f
C324 plus.n47 a_n2390_n1288# 1.21039f
.ends

