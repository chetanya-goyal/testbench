* NGSPICE file created from diffpair171.ext - technology: sky130A

.subckt diffpair171 minus drain_right drain_left source plus
X0 drain_right minus source a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X1 a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X2 source minus drain_right a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X3 a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X4 drain_right minus source a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X5 a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X6 drain_left plus source a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X7 a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X8 drain_left plus source a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X9 source minus drain_right a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X10 source plus drain_left a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X11 source plus drain_left a_n1034_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
.ends

