* NGSPICE file created from diffpair41.ext - technology: sky130A

.subckt diffpair41 minus drain_right drain_left source plus
X0 source.t7 minus.t0 drain_right.t0 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X1 source.t3 plus.t0 drain_left.t3 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 source.t6 minus.t1 drain_right.t3 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_left.t2 plus.t1 source.t2 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X5 drain_right.t2 minus.t2 source.t5 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X6 drain_right.t1 minus.t3 source.t4 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X7 drain_left.t1 plus.t2 source.t1 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X8 source.t0 plus.t3 drain_left.t0 a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X9 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X10 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X11 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
R0 minus.n0 minus.t2 147.749
R1 minus.n1 minus.t1 147.749
R2 minus.n0 minus.t0 147.724
R3 minus.n1 minus.t3 147.724
R4 minus.n2 minus.n0 95.6647
R5 minus.n2 minus.n1 76.7783
R6 minus minus.n2 0.188
R7 drain_right drain_right.n0 260.043
R8 drain_right drain_right.n1 246.501
R9 drain_right.n0 drain_right.t3 19.8005
R10 drain_right.n0 drain_right.t1 19.8005
R11 drain_right.n1 drain_right.t0 19.8005
R12 drain_right.n1 drain_right.t2 19.8005
R13 source.n0 source.t1 243.255
R14 source.n1 source.t3 243.255
R15 source.n2 source.t5 243.255
R16 source.n3 source.t7 243.255
R17 source.n7 source.t4 243.254
R18 source.n6 source.t6 243.254
R19 source.n5 source.t2 243.254
R20 source.n4 source.t0 243.254
R21 source.n4 source.n3 13.6699
R22 source.n8 source.n0 8.04922
R23 source.n8 source.n7 5.62119
R24 source.n3 source.n2 0.716017
R25 source.n1 source.n0 0.716017
R26 source.n5 source.n4 0.716017
R27 source.n7 source.n6 0.716017
R28 source.n2 source.n1 0.470328
R29 source.n6 source.n5 0.470328
R30 source source.n8 0.188
R31 plus.n0 plus.t0 147.749
R32 plus.n1 plus.t1 147.749
R33 plus.n0 plus.t2 147.724
R34 plus.n1 plus.t3 147.724
R35 plus plus.n1 93.7124
R36 plus plus.n0 78.2556
R37 drain_left drain_left.n0 260.596
R38 drain_left drain_left.n1 246.501
R39 drain_left.n0 drain_left.t0 19.8005
R40 drain_left.n0 drain_left.t2 19.8005
R41 drain_left.n1 drain_left.t3 19.8005
R42 drain_left.n1 drain_left.t1 19.8005
C0 plus drain_right 0.274688f
C1 plus source 0.642999f
C2 plus minus 2.6303f
C3 drain_left drain_right 0.522929f
C4 drain_left source 1.9499f
C5 drain_left minus 0.177386f
C6 source drain_right 1.94964f
C7 minus drain_right 0.485446f
C8 source minus 0.629135f
C9 plus drain_left 0.598857f
C10 drain_right a_n1214_n1088# 1.6441f
C11 drain_left a_n1214_n1088# 1.76467f
C12 source a_n1214_n1088# 2.19687f
C13 minus a_n1214_n1088# 3.687742f
C14 plus a_n1214_n1088# 5.31956f
C15 plus.t2 a_n1214_n1088# 0.077916f
C16 plus.t0 a_n1214_n1088# 0.077934f
C17 plus.n0 a_n1214_n1088# 0.155069f
C18 plus.t3 a_n1214_n1088# 0.077916f
C19 plus.t1 a_n1214_n1088# 0.077934f
C20 plus.n1 a_n1214_n1088# 0.324826f
C21 minus.t2 a_n1214_n1088# 0.07558f
C22 minus.t0 a_n1214_n1088# 0.075562f
C23 minus.n0 a_n1214_n1088# 0.331165f
C24 minus.t1 a_n1214_n1088# 0.07558f
C25 minus.t3 a_n1214_n1088# 0.075562f
C26 minus.n1 a_n1214_n1088# 0.143791f
C27 minus.n2 a_n1214_n1088# 1.79726f
.ends

