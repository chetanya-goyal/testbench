* NGSPICE file created from diffpair121.ext - technology: sky130A

.subckt diffpair121 minus drain_right drain_left source plus
X0 drain_right minus source a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X1 source plus drain_left a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X2 source minus drain_right a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X3 a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X4 source plus drain_left a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X5 a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X6 a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X7 drain_right minus source a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X8 drain_left plus source a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X9 source minus drain_right a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X10 a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X11 drain_left plus source a_n1214_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
.ends

