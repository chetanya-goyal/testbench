* NGSPICE file created from diffpair704.ext - technology: sky130A

.subckt diffpair704 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t19 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X1 source.t1 plus.t0 drain_left.t9 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X2 source.t18 minus.t1 drain_right.t8 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X3 a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.7
X4 drain_left.t8 plus.t1 source.t8 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X5 source.t17 minus.t2 drain_right.t7 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X6 a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X7 drain_right.t6 minus.t3 source.t16 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X8 a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X9 drain_left.t7 plus.t2 source.t5 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X10 drain_left.t6 plus.t3 source.t0 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X11 source.t11 minus.t4 drain_right.t5 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X12 drain_right.t4 minus.t5 source.t13 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X13 drain_right.t3 minus.t6 source.t12 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X14 a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X15 drain_right.t2 minus.t7 source.t14 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X16 source.t9 plus.t4 drain_left.t5 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X17 source.t2 plus.t5 drain_left.t4 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X18 drain_left.t3 plus.t6 source.t3 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X19 drain_right.t1 minus.t8 source.t15 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X20 source.t7 plus.t7 drain_left.t2 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X21 drain_left.t1 plus.t8 source.t4 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X22 source.t10 minus.t9 drain_right.t0 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X23 drain_left.t0 plus.t9 source.t6 a_n1952_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
R0 minus.n3 minus.t8 939.582
R1 minus.n17 minus.t5 939.582
R2 minus.n4 minus.t2 916.833
R3 minus.n6 minus.t7 916.833
R4 minus.n10 minus.t9 916.833
R5 minus.n12 minus.t6 916.833
R6 minus.n18 minus.t4 916.833
R7 minus.n20 minus.t0 916.833
R8 minus.n24 minus.t1 916.833
R9 minus.n26 minus.t3 916.833
R10 minus.n13 minus.n12 161.3
R11 minus.n11 minus.n0 161.3
R12 minus.n10 minus.n9 161.3
R13 minus.n8 minus.n1 161.3
R14 minus.n7 minus.n6 161.3
R15 minus.n5 minus.n2 161.3
R16 minus.n27 minus.n26 161.3
R17 minus.n25 minus.n14 161.3
R18 minus.n24 minus.n23 161.3
R19 minus.n22 minus.n15 161.3
R20 minus.n21 minus.n20 161.3
R21 minus.n19 minus.n16 161.3
R22 minus.n28 minus.n13 46.5024
R23 minus.n3 minus.n2 44.8741
R24 minus.n17 minus.n16 44.8741
R25 minus.n12 minus.n11 30.6732
R26 minus.n26 minus.n25 30.6732
R27 minus.n5 minus.n4 26.2914
R28 minus.n10 minus.n1 26.2914
R29 minus.n19 minus.n18 26.2914
R30 minus.n24 minus.n15 26.2914
R31 minus.n6 minus.n5 21.9096
R32 minus.n6 minus.n1 21.9096
R33 minus.n20 minus.n19 21.9096
R34 minus.n20 minus.n15 21.9096
R35 minus.n4 minus.n3 19.0667
R36 minus.n18 minus.n17 19.0667
R37 minus.n11 minus.n10 17.5278
R38 minus.n25 minus.n24 17.5278
R39 minus.n28 minus.n27 6.63876
R40 minus.n13 minus.n0 0.189894
R41 minus.n9 minus.n0 0.189894
R42 minus.n9 minus.n8 0.189894
R43 minus.n8 minus.n7 0.189894
R44 minus.n7 minus.n2 0.189894
R45 minus.n21 minus.n16 0.189894
R46 minus.n22 minus.n21 0.189894
R47 minus.n23 minus.n22 0.189894
R48 minus.n23 minus.n14 0.189894
R49 minus.n27 minus.n14 0.189894
R50 minus minus.n28 0.188
R51 source.n570 source.n436 289.615
R52 source.n426 source.n292 289.615
R53 source.n134 source.n0 289.615
R54 source.n278 source.n144 289.615
R55 source.n480 source.n479 185
R56 source.n485 source.n484 185
R57 source.n487 source.n486 185
R58 source.n476 source.n475 185
R59 source.n493 source.n492 185
R60 source.n495 source.n494 185
R61 source.n472 source.n471 185
R62 source.n502 source.n501 185
R63 source.n503 source.n470 185
R64 source.n505 source.n504 185
R65 source.n468 source.n467 185
R66 source.n511 source.n510 185
R67 source.n513 source.n512 185
R68 source.n464 source.n463 185
R69 source.n519 source.n518 185
R70 source.n521 source.n520 185
R71 source.n460 source.n459 185
R72 source.n527 source.n526 185
R73 source.n529 source.n528 185
R74 source.n456 source.n455 185
R75 source.n535 source.n534 185
R76 source.n537 source.n536 185
R77 source.n452 source.n451 185
R78 source.n543 source.n542 185
R79 source.n546 source.n545 185
R80 source.n544 source.n448 185
R81 source.n551 source.n447 185
R82 source.n553 source.n552 185
R83 source.n555 source.n554 185
R84 source.n444 source.n443 185
R85 source.n561 source.n560 185
R86 source.n563 source.n562 185
R87 source.n440 source.n439 185
R88 source.n569 source.n568 185
R89 source.n571 source.n570 185
R90 source.n336 source.n335 185
R91 source.n341 source.n340 185
R92 source.n343 source.n342 185
R93 source.n332 source.n331 185
R94 source.n349 source.n348 185
R95 source.n351 source.n350 185
R96 source.n328 source.n327 185
R97 source.n358 source.n357 185
R98 source.n359 source.n326 185
R99 source.n361 source.n360 185
R100 source.n324 source.n323 185
R101 source.n367 source.n366 185
R102 source.n369 source.n368 185
R103 source.n320 source.n319 185
R104 source.n375 source.n374 185
R105 source.n377 source.n376 185
R106 source.n316 source.n315 185
R107 source.n383 source.n382 185
R108 source.n385 source.n384 185
R109 source.n312 source.n311 185
R110 source.n391 source.n390 185
R111 source.n393 source.n392 185
R112 source.n308 source.n307 185
R113 source.n399 source.n398 185
R114 source.n402 source.n401 185
R115 source.n400 source.n304 185
R116 source.n407 source.n303 185
R117 source.n409 source.n408 185
R118 source.n411 source.n410 185
R119 source.n300 source.n299 185
R120 source.n417 source.n416 185
R121 source.n419 source.n418 185
R122 source.n296 source.n295 185
R123 source.n425 source.n424 185
R124 source.n427 source.n426 185
R125 source.n135 source.n134 185
R126 source.n133 source.n132 185
R127 source.n4 source.n3 185
R128 source.n127 source.n126 185
R129 source.n125 source.n124 185
R130 source.n8 source.n7 185
R131 source.n119 source.n118 185
R132 source.n117 source.n116 185
R133 source.n115 source.n11 185
R134 source.n15 source.n12 185
R135 source.n110 source.n109 185
R136 source.n108 source.n107 185
R137 source.n17 source.n16 185
R138 source.n102 source.n101 185
R139 source.n100 source.n99 185
R140 source.n21 source.n20 185
R141 source.n94 source.n93 185
R142 source.n92 source.n91 185
R143 source.n25 source.n24 185
R144 source.n86 source.n85 185
R145 source.n84 source.n83 185
R146 source.n29 source.n28 185
R147 source.n78 source.n77 185
R148 source.n76 source.n75 185
R149 source.n33 source.n32 185
R150 source.n70 source.n69 185
R151 source.n68 source.n35 185
R152 source.n67 source.n66 185
R153 source.n38 source.n36 185
R154 source.n61 source.n60 185
R155 source.n59 source.n58 185
R156 source.n42 source.n41 185
R157 source.n53 source.n52 185
R158 source.n51 source.n50 185
R159 source.n46 source.n45 185
R160 source.n279 source.n278 185
R161 source.n277 source.n276 185
R162 source.n148 source.n147 185
R163 source.n271 source.n270 185
R164 source.n269 source.n268 185
R165 source.n152 source.n151 185
R166 source.n263 source.n262 185
R167 source.n261 source.n260 185
R168 source.n259 source.n155 185
R169 source.n159 source.n156 185
R170 source.n254 source.n253 185
R171 source.n252 source.n251 185
R172 source.n161 source.n160 185
R173 source.n246 source.n245 185
R174 source.n244 source.n243 185
R175 source.n165 source.n164 185
R176 source.n238 source.n237 185
R177 source.n236 source.n235 185
R178 source.n169 source.n168 185
R179 source.n230 source.n229 185
R180 source.n228 source.n227 185
R181 source.n173 source.n172 185
R182 source.n222 source.n221 185
R183 source.n220 source.n219 185
R184 source.n177 source.n176 185
R185 source.n214 source.n213 185
R186 source.n212 source.n179 185
R187 source.n211 source.n210 185
R188 source.n182 source.n180 185
R189 source.n205 source.n204 185
R190 source.n203 source.n202 185
R191 source.n186 source.n185 185
R192 source.n197 source.n196 185
R193 source.n195 source.n194 185
R194 source.n190 source.n189 185
R195 source.n481 source.t16 149.524
R196 source.n337 source.t6 149.524
R197 source.n47 source.t5 149.524
R198 source.n191 source.t15 149.524
R199 source.n485 source.n479 104.615
R200 source.n486 source.n485 104.615
R201 source.n486 source.n475 104.615
R202 source.n493 source.n475 104.615
R203 source.n494 source.n493 104.615
R204 source.n494 source.n471 104.615
R205 source.n502 source.n471 104.615
R206 source.n503 source.n502 104.615
R207 source.n504 source.n503 104.615
R208 source.n504 source.n467 104.615
R209 source.n511 source.n467 104.615
R210 source.n512 source.n511 104.615
R211 source.n512 source.n463 104.615
R212 source.n519 source.n463 104.615
R213 source.n520 source.n519 104.615
R214 source.n520 source.n459 104.615
R215 source.n527 source.n459 104.615
R216 source.n528 source.n527 104.615
R217 source.n528 source.n455 104.615
R218 source.n535 source.n455 104.615
R219 source.n536 source.n535 104.615
R220 source.n536 source.n451 104.615
R221 source.n543 source.n451 104.615
R222 source.n545 source.n543 104.615
R223 source.n545 source.n544 104.615
R224 source.n544 source.n447 104.615
R225 source.n553 source.n447 104.615
R226 source.n554 source.n553 104.615
R227 source.n554 source.n443 104.615
R228 source.n561 source.n443 104.615
R229 source.n562 source.n561 104.615
R230 source.n562 source.n439 104.615
R231 source.n569 source.n439 104.615
R232 source.n570 source.n569 104.615
R233 source.n341 source.n335 104.615
R234 source.n342 source.n341 104.615
R235 source.n342 source.n331 104.615
R236 source.n349 source.n331 104.615
R237 source.n350 source.n349 104.615
R238 source.n350 source.n327 104.615
R239 source.n358 source.n327 104.615
R240 source.n359 source.n358 104.615
R241 source.n360 source.n359 104.615
R242 source.n360 source.n323 104.615
R243 source.n367 source.n323 104.615
R244 source.n368 source.n367 104.615
R245 source.n368 source.n319 104.615
R246 source.n375 source.n319 104.615
R247 source.n376 source.n375 104.615
R248 source.n376 source.n315 104.615
R249 source.n383 source.n315 104.615
R250 source.n384 source.n383 104.615
R251 source.n384 source.n311 104.615
R252 source.n391 source.n311 104.615
R253 source.n392 source.n391 104.615
R254 source.n392 source.n307 104.615
R255 source.n399 source.n307 104.615
R256 source.n401 source.n399 104.615
R257 source.n401 source.n400 104.615
R258 source.n400 source.n303 104.615
R259 source.n409 source.n303 104.615
R260 source.n410 source.n409 104.615
R261 source.n410 source.n299 104.615
R262 source.n417 source.n299 104.615
R263 source.n418 source.n417 104.615
R264 source.n418 source.n295 104.615
R265 source.n425 source.n295 104.615
R266 source.n426 source.n425 104.615
R267 source.n134 source.n133 104.615
R268 source.n133 source.n3 104.615
R269 source.n126 source.n3 104.615
R270 source.n126 source.n125 104.615
R271 source.n125 source.n7 104.615
R272 source.n118 source.n7 104.615
R273 source.n118 source.n117 104.615
R274 source.n117 source.n11 104.615
R275 source.n15 source.n11 104.615
R276 source.n109 source.n15 104.615
R277 source.n109 source.n108 104.615
R278 source.n108 source.n16 104.615
R279 source.n101 source.n16 104.615
R280 source.n101 source.n100 104.615
R281 source.n100 source.n20 104.615
R282 source.n93 source.n20 104.615
R283 source.n93 source.n92 104.615
R284 source.n92 source.n24 104.615
R285 source.n85 source.n24 104.615
R286 source.n85 source.n84 104.615
R287 source.n84 source.n28 104.615
R288 source.n77 source.n28 104.615
R289 source.n77 source.n76 104.615
R290 source.n76 source.n32 104.615
R291 source.n69 source.n32 104.615
R292 source.n69 source.n68 104.615
R293 source.n68 source.n67 104.615
R294 source.n67 source.n36 104.615
R295 source.n60 source.n36 104.615
R296 source.n60 source.n59 104.615
R297 source.n59 source.n41 104.615
R298 source.n52 source.n41 104.615
R299 source.n52 source.n51 104.615
R300 source.n51 source.n45 104.615
R301 source.n278 source.n277 104.615
R302 source.n277 source.n147 104.615
R303 source.n270 source.n147 104.615
R304 source.n270 source.n269 104.615
R305 source.n269 source.n151 104.615
R306 source.n262 source.n151 104.615
R307 source.n262 source.n261 104.615
R308 source.n261 source.n155 104.615
R309 source.n159 source.n155 104.615
R310 source.n253 source.n159 104.615
R311 source.n253 source.n252 104.615
R312 source.n252 source.n160 104.615
R313 source.n245 source.n160 104.615
R314 source.n245 source.n244 104.615
R315 source.n244 source.n164 104.615
R316 source.n237 source.n164 104.615
R317 source.n237 source.n236 104.615
R318 source.n236 source.n168 104.615
R319 source.n229 source.n168 104.615
R320 source.n229 source.n228 104.615
R321 source.n228 source.n172 104.615
R322 source.n221 source.n172 104.615
R323 source.n221 source.n220 104.615
R324 source.n220 source.n176 104.615
R325 source.n213 source.n176 104.615
R326 source.n213 source.n212 104.615
R327 source.n212 source.n211 104.615
R328 source.n211 source.n180 104.615
R329 source.n204 source.n180 104.615
R330 source.n204 source.n203 104.615
R331 source.n203 source.n185 104.615
R332 source.n196 source.n185 104.615
R333 source.n196 source.n195 104.615
R334 source.n195 source.n189 104.615
R335 source.t16 source.n479 52.3082
R336 source.t6 source.n335 52.3082
R337 source.t5 source.n45 52.3082
R338 source.t15 source.n189 52.3082
R339 source.n435 source.n434 42.0366
R340 source.n433 source.n432 42.0366
R341 source.n291 source.n290 42.0366
R342 source.n289 source.n288 42.0366
R343 source.n141 source.n140 42.0366
R344 source.n143 source.n142 42.0366
R345 source.n285 source.n284 42.0366
R346 source.n287 source.n286 42.0366
R347 source.n289 source.n287 32.9121
R348 source.n575 source.n574 30.6338
R349 source.n431 source.n430 30.6338
R350 source.n139 source.n138 30.6338
R351 source.n283 source.n282 30.6338
R352 source.n576 source.n139 26.3172
R353 source.n505 source.n470 13.1884
R354 source.n552 source.n551 13.1884
R355 source.n361 source.n326 13.1884
R356 source.n408 source.n407 13.1884
R357 source.n116 source.n115 13.1884
R358 source.n70 source.n35 13.1884
R359 source.n260 source.n259 13.1884
R360 source.n214 source.n179 13.1884
R361 source.n501 source.n500 12.8005
R362 source.n506 source.n468 12.8005
R363 source.n550 source.n448 12.8005
R364 source.n555 source.n446 12.8005
R365 source.n357 source.n356 12.8005
R366 source.n362 source.n324 12.8005
R367 source.n406 source.n304 12.8005
R368 source.n411 source.n302 12.8005
R369 source.n119 source.n10 12.8005
R370 source.n114 source.n12 12.8005
R371 source.n71 source.n33 12.8005
R372 source.n66 source.n37 12.8005
R373 source.n263 source.n154 12.8005
R374 source.n258 source.n156 12.8005
R375 source.n215 source.n177 12.8005
R376 source.n210 source.n181 12.8005
R377 source.n499 source.n472 12.0247
R378 source.n510 source.n509 12.0247
R379 source.n547 source.n546 12.0247
R380 source.n556 source.n444 12.0247
R381 source.n355 source.n328 12.0247
R382 source.n366 source.n365 12.0247
R383 source.n403 source.n402 12.0247
R384 source.n412 source.n300 12.0247
R385 source.n120 source.n8 12.0247
R386 source.n111 source.n110 12.0247
R387 source.n75 source.n74 12.0247
R388 source.n65 source.n38 12.0247
R389 source.n264 source.n152 12.0247
R390 source.n255 source.n254 12.0247
R391 source.n219 source.n218 12.0247
R392 source.n209 source.n182 12.0247
R393 source.n496 source.n495 11.249
R394 source.n513 source.n466 11.249
R395 source.n542 source.n450 11.249
R396 source.n560 source.n559 11.249
R397 source.n352 source.n351 11.249
R398 source.n369 source.n322 11.249
R399 source.n398 source.n306 11.249
R400 source.n416 source.n415 11.249
R401 source.n124 source.n123 11.249
R402 source.n107 source.n14 11.249
R403 source.n78 source.n31 11.249
R404 source.n62 source.n61 11.249
R405 source.n268 source.n267 11.249
R406 source.n251 source.n158 11.249
R407 source.n222 source.n175 11.249
R408 source.n206 source.n205 11.249
R409 source.n492 source.n474 10.4732
R410 source.n514 source.n464 10.4732
R411 source.n541 source.n452 10.4732
R412 source.n563 source.n442 10.4732
R413 source.n348 source.n330 10.4732
R414 source.n370 source.n320 10.4732
R415 source.n397 source.n308 10.4732
R416 source.n419 source.n298 10.4732
R417 source.n127 source.n6 10.4732
R418 source.n106 source.n17 10.4732
R419 source.n79 source.n29 10.4732
R420 source.n58 source.n40 10.4732
R421 source.n271 source.n150 10.4732
R422 source.n250 source.n161 10.4732
R423 source.n223 source.n173 10.4732
R424 source.n202 source.n184 10.4732
R425 source.n481 source.n480 10.2747
R426 source.n337 source.n336 10.2747
R427 source.n47 source.n46 10.2747
R428 source.n191 source.n190 10.2747
R429 source.n491 source.n476 9.69747
R430 source.n518 source.n517 9.69747
R431 source.n538 source.n537 9.69747
R432 source.n564 source.n440 9.69747
R433 source.n347 source.n332 9.69747
R434 source.n374 source.n373 9.69747
R435 source.n394 source.n393 9.69747
R436 source.n420 source.n296 9.69747
R437 source.n128 source.n4 9.69747
R438 source.n103 source.n102 9.69747
R439 source.n83 source.n82 9.69747
R440 source.n57 source.n42 9.69747
R441 source.n272 source.n148 9.69747
R442 source.n247 source.n246 9.69747
R443 source.n227 source.n226 9.69747
R444 source.n201 source.n186 9.69747
R445 source.n574 source.n573 9.45567
R446 source.n430 source.n429 9.45567
R447 source.n138 source.n137 9.45567
R448 source.n282 source.n281 9.45567
R449 source.n438 source.n437 9.3005
R450 source.n567 source.n566 9.3005
R451 source.n565 source.n564 9.3005
R452 source.n442 source.n441 9.3005
R453 source.n559 source.n558 9.3005
R454 source.n557 source.n556 9.3005
R455 source.n446 source.n445 9.3005
R456 source.n525 source.n524 9.3005
R457 source.n523 source.n522 9.3005
R458 source.n462 source.n461 9.3005
R459 source.n517 source.n516 9.3005
R460 source.n515 source.n514 9.3005
R461 source.n466 source.n465 9.3005
R462 source.n509 source.n508 9.3005
R463 source.n507 source.n506 9.3005
R464 source.n483 source.n482 9.3005
R465 source.n478 source.n477 9.3005
R466 source.n489 source.n488 9.3005
R467 source.n491 source.n490 9.3005
R468 source.n474 source.n473 9.3005
R469 source.n497 source.n496 9.3005
R470 source.n499 source.n498 9.3005
R471 source.n500 source.n469 9.3005
R472 source.n458 source.n457 9.3005
R473 source.n531 source.n530 9.3005
R474 source.n533 source.n532 9.3005
R475 source.n454 source.n453 9.3005
R476 source.n539 source.n538 9.3005
R477 source.n541 source.n540 9.3005
R478 source.n450 source.n449 9.3005
R479 source.n548 source.n547 9.3005
R480 source.n550 source.n549 9.3005
R481 source.n573 source.n572 9.3005
R482 source.n294 source.n293 9.3005
R483 source.n423 source.n422 9.3005
R484 source.n421 source.n420 9.3005
R485 source.n298 source.n297 9.3005
R486 source.n415 source.n414 9.3005
R487 source.n413 source.n412 9.3005
R488 source.n302 source.n301 9.3005
R489 source.n381 source.n380 9.3005
R490 source.n379 source.n378 9.3005
R491 source.n318 source.n317 9.3005
R492 source.n373 source.n372 9.3005
R493 source.n371 source.n370 9.3005
R494 source.n322 source.n321 9.3005
R495 source.n365 source.n364 9.3005
R496 source.n363 source.n362 9.3005
R497 source.n339 source.n338 9.3005
R498 source.n334 source.n333 9.3005
R499 source.n345 source.n344 9.3005
R500 source.n347 source.n346 9.3005
R501 source.n330 source.n329 9.3005
R502 source.n353 source.n352 9.3005
R503 source.n355 source.n354 9.3005
R504 source.n356 source.n325 9.3005
R505 source.n314 source.n313 9.3005
R506 source.n387 source.n386 9.3005
R507 source.n389 source.n388 9.3005
R508 source.n310 source.n309 9.3005
R509 source.n395 source.n394 9.3005
R510 source.n397 source.n396 9.3005
R511 source.n306 source.n305 9.3005
R512 source.n404 source.n403 9.3005
R513 source.n406 source.n405 9.3005
R514 source.n429 source.n428 9.3005
R515 source.n49 source.n48 9.3005
R516 source.n44 source.n43 9.3005
R517 source.n55 source.n54 9.3005
R518 source.n57 source.n56 9.3005
R519 source.n40 source.n39 9.3005
R520 source.n63 source.n62 9.3005
R521 source.n65 source.n64 9.3005
R522 source.n37 source.n34 9.3005
R523 source.n96 source.n95 9.3005
R524 source.n98 source.n97 9.3005
R525 source.n19 source.n18 9.3005
R526 source.n104 source.n103 9.3005
R527 source.n106 source.n105 9.3005
R528 source.n14 source.n13 9.3005
R529 source.n112 source.n111 9.3005
R530 source.n114 source.n113 9.3005
R531 source.n137 source.n136 9.3005
R532 source.n2 source.n1 9.3005
R533 source.n131 source.n130 9.3005
R534 source.n129 source.n128 9.3005
R535 source.n6 source.n5 9.3005
R536 source.n123 source.n122 9.3005
R537 source.n121 source.n120 9.3005
R538 source.n10 source.n9 9.3005
R539 source.n23 source.n22 9.3005
R540 source.n90 source.n89 9.3005
R541 source.n88 source.n87 9.3005
R542 source.n27 source.n26 9.3005
R543 source.n82 source.n81 9.3005
R544 source.n80 source.n79 9.3005
R545 source.n31 source.n30 9.3005
R546 source.n74 source.n73 9.3005
R547 source.n72 source.n71 9.3005
R548 source.n193 source.n192 9.3005
R549 source.n188 source.n187 9.3005
R550 source.n199 source.n198 9.3005
R551 source.n201 source.n200 9.3005
R552 source.n184 source.n183 9.3005
R553 source.n207 source.n206 9.3005
R554 source.n209 source.n208 9.3005
R555 source.n181 source.n178 9.3005
R556 source.n240 source.n239 9.3005
R557 source.n242 source.n241 9.3005
R558 source.n163 source.n162 9.3005
R559 source.n248 source.n247 9.3005
R560 source.n250 source.n249 9.3005
R561 source.n158 source.n157 9.3005
R562 source.n256 source.n255 9.3005
R563 source.n258 source.n257 9.3005
R564 source.n281 source.n280 9.3005
R565 source.n146 source.n145 9.3005
R566 source.n275 source.n274 9.3005
R567 source.n273 source.n272 9.3005
R568 source.n150 source.n149 9.3005
R569 source.n267 source.n266 9.3005
R570 source.n265 source.n264 9.3005
R571 source.n154 source.n153 9.3005
R572 source.n167 source.n166 9.3005
R573 source.n234 source.n233 9.3005
R574 source.n232 source.n231 9.3005
R575 source.n171 source.n170 9.3005
R576 source.n226 source.n225 9.3005
R577 source.n224 source.n223 9.3005
R578 source.n175 source.n174 9.3005
R579 source.n218 source.n217 9.3005
R580 source.n216 source.n215 9.3005
R581 source.n488 source.n487 8.92171
R582 source.n521 source.n462 8.92171
R583 source.n534 source.n454 8.92171
R584 source.n568 source.n567 8.92171
R585 source.n344 source.n343 8.92171
R586 source.n377 source.n318 8.92171
R587 source.n390 source.n310 8.92171
R588 source.n424 source.n423 8.92171
R589 source.n132 source.n131 8.92171
R590 source.n99 source.n19 8.92171
R591 source.n86 source.n27 8.92171
R592 source.n54 source.n53 8.92171
R593 source.n276 source.n275 8.92171
R594 source.n243 source.n163 8.92171
R595 source.n230 source.n171 8.92171
R596 source.n198 source.n197 8.92171
R597 source.n484 source.n478 8.14595
R598 source.n522 source.n460 8.14595
R599 source.n533 source.n456 8.14595
R600 source.n571 source.n438 8.14595
R601 source.n340 source.n334 8.14595
R602 source.n378 source.n316 8.14595
R603 source.n389 source.n312 8.14595
R604 source.n427 source.n294 8.14595
R605 source.n135 source.n2 8.14595
R606 source.n98 source.n21 8.14595
R607 source.n87 source.n25 8.14595
R608 source.n50 source.n44 8.14595
R609 source.n279 source.n146 8.14595
R610 source.n242 source.n165 8.14595
R611 source.n231 source.n169 8.14595
R612 source.n194 source.n188 8.14595
R613 source.n483 source.n480 7.3702
R614 source.n526 source.n525 7.3702
R615 source.n530 source.n529 7.3702
R616 source.n572 source.n436 7.3702
R617 source.n339 source.n336 7.3702
R618 source.n382 source.n381 7.3702
R619 source.n386 source.n385 7.3702
R620 source.n428 source.n292 7.3702
R621 source.n136 source.n0 7.3702
R622 source.n95 source.n94 7.3702
R623 source.n91 source.n90 7.3702
R624 source.n49 source.n46 7.3702
R625 source.n280 source.n144 7.3702
R626 source.n239 source.n238 7.3702
R627 source.n235 source.n234 7.3702
R628 source.n193 source.n190 7.3702
R629 source.n526 source.n458 6.59444
R630 source.n529 source.n458 6.59444
R631 source.n574 source.n436 6.59444
R632 source.n382 source.n314 6.59444
R633 source.n385 source.n314 6.59444
R634 source.n430 source.n292 6.59444
R635 source.n138 source.n0 6.59444
R636 source.n94 source.n23 6.59444
R637 source.n91 source.n23 6.59444
R638 source.n282 source.n144 6.59444
R639 source.n238 source.n167 6.59444
R640 source.n235 source.n167 6.59444
R641 source.n484 source.n483 5.81868
R642 source.n525 source.n460 5.81868
R643 source.n530 source.n456 5.81868
R644 source.n572 source.n571 5.81868
R645 source.n340 source.n339 5.81868
R646 source.n381 source.n316 5.81868
R647 source.n386 source.n312 5.81868
R648 source.n428 source.n427 5.81868
R649 source.n136 source.n135 5.81868
R650 source.n95 source.n21 5.81868
R651 source.n90 source.n25 5.81868
R652 source.n50 source.n49 5.81868
R653 source.n280 source.n279 5.81868
R654 source.n239 source.n165 5.81868
R655 source.n234 source.n169 5.81868
R656 source.n194 source.n193 5.81868
R657 source.n576 source.n575 5.7074
R658 source.n487 source.n478 5.04292
R659 source.n522 source.n521 5.04292
R660 source.n534 source.n533 5.04292
R661 source.n568 source.n438 5.04292
R662 source.n343 source.n334 5.04292
R663 source.n378 source.n377 5.04292
R664 source.n390 source.n389 5.04292
R665 source.n424 source.n294 5.04292
R666 source.n132 source.n2 5.04292
R667 source.n99 source.n98 5.04292
R668 source.n87 source.n86 5.04292
R669 source.n53 source.n44 5.04292
R670 source.n276 source.n146 5.04292
R671 source.n243 source.n242 5.04292
R672 source.n231 source.n230 5.04292
R673 source.n197 source.n188 5.04292
R674 source.n488 source.n476 4.26717
R675 source.n518 source.n462 4.26717
R676 source.n537 source.n454 4.26717
R677 source.n567 source.n440 4.26717
R678 source.n344 source.n332 4.26717
R679 source.n374 source.n318 4.26717
R680 source.n393 source.n310 4.26717
R681 source.n423 source.n296 4.26717
R682 source.n131 source.n4 4.26717
R683 source.n102 source.n19 4.26717
R684 source.n83 source.n27 4.26717
R685 source.n54 source.n42 4.26717
R686 source.n275 source.n148 4.26717
R687 source.n246 source.n163 4.26717
R688 source.n227 source.n171 4.26717
R689 source.n198 source.n186 4.26717
R690 source.n492 source.n491 3.49141
R691 source.n517 source.n464 3.49141
R692 source.n538 source.n452 3.49141
R693 source.n564 source.n563 3.49141
R694 source.n348 source.n347 3.49141
R695 source.n373 source.n320 3.49141
R696 source.n394 source.n308 3.49141
R697 source.n420 source.n419 3.49141
R698 source.n128 source.n127 3.49141
R699 source.n103 source.n17 3.49141
R700 source.n82 source.n29 3.49141
R701 source.n58 source.n57 3.49141
R702 source.n272 source.n271 3.49141
R703 source.n247 source.n161 3.49141
R704 source.n226 source.n173 3.49141
R705 source.n202 source.n201 3.49141
R706 source.n48 source.n47 2.84303
R707 source.n192 source.n191 2.84303
R708 source.n482 source.n481 2.84303
R709 source.n338 source.n337 2.84303
R710 source.n495 source.n474 2.71565
R711 source.n514 source.n513 2.71565
R712 source.n542 source.n541 2.71565
R713 source.n560 source.n442 2.71565
R714 source.n351 source.n330 2.71565
R715 source.n370 source.n369 2.71565
R716 source.n398 source.n397 2.71565
R717 source.n416 source.n298 2.71565
R718 source.n124 source.n6 2.71565
R719 source.n107 source.n106 2.71565
R720 source.n79 source.n78 2.71565
R721 source.n61 source.n40 2.71565
R722 source.n268 source.n150 2.71565
R723 source.n251 source.n250 2.71565
R724 source.n223 source.n222 2.71565
R725 source.n205 source.n184 2.71565
R726 source.n496 source.n472 1.93989
R727 source.n510 source.n466 1.93989
R728 source.n546 source.n450 1.93989
R729 source.n559 source.n444 1.93989
R730 source.n352 source.n328 1.93989
R731 source.n366 source.n322 1.93989
R732 source.n402 source.n306 1.93989
R733 source.n415 source.n300 1.93989
R734 source.n123 source.n8 1.93989
R735 source.n110 source.n14 1.93989
R736 source.n75 source.n31 1.93989
R737 source.n62 source.n38 1.93989
R738 source.n267 source.n152 1.93989
R739 source.n254 source.n158 1.93989
R740 source.n219 source.n175 1.93989
R741 source.n206 source.n182 1.93989
R742 source.n501 source.n499 1.16414
R743 source.n509 source.n468 1.16414
R744 source.n547 source.n448 1.16414
R745 source.n556 source.n555 1.16414
R746 source.n357 source.n355 1.16414
R747 source.n365 source.n324 1.16414
R748 source.n403 source.n304 1.16414
R749 source.n412 source.n411 1.16414
R750 source.n120 source.n119 1.16414
R751 source.n111 source.n12 1.16414
R752 source.n74 source.n33 1.16414
R753 source.n66 source.n65 1.16414
R754 source.n264 source.n263 1.16414
R755 source.n255 source.n156 1.16414
R756 source.n218 source.n177 1.16414
R757 source.n210 source.n209 1.16414
R758 source.n283 source.n143 0.914293
R759 source.n433 source.n431 0.914293
R760 source.n287 source.n285 0.888431
R761 source.n285 source.n283 0.888431
R762 source.n143 source.n141 0.888431
R763 source.n141 source.n139 0.888431
R764 source.n291 source.n289 0.888431
R765 source.n431 source.n291 0.888431
R766 source.n435 source.n433 0.888431
R767 source.n575 source.n435 0.888431
R768 source.n434 source.t19 0.7925
R769 source.n434 source.t18 0.7925
R770 source.n432 source.t13 0.7925
R771 source.n432 source.t11 0.7925
R772 source.n290 source.t4 0.7925
R773 source.n290 source.t1 0.7925
R774 source.n288 source.t3 0.7925
R775 source.n288 source.t9 0.7925
R776 source.n140 source.t8 0.7925
R777 source.n140 source.t2 0.7925
R778 source.n142 source.t0 0.7925
R779 source.n142 source.t7 0.7925
R780 source.n284 source.t14 0.7925
R781 source.n284 source.t17 0.7925
R782 source.n286 source.t12 0.7925
R783 source.n286 source.t10 0.7925
R784 source.n500 source.n470 0.388379
R785 source.n506 source.n505 0.388379
R786 source.n551 source.n550 0.388379
R787 source.n552 source.n446 0.388379
R788 source.n356 source.n326 0.388379
R789 source.n362 source.n361 0.388379
R790 source.n407 source.n406 0.388379
R791 source.n408 source.n302 0.388379
R792 source.n116 source.n10 0.388379
R793 source.n115 source.n114 0.388379
R794 source.n71 source.n70 0.388379
R795 source.n37 source.n35 0.388379
R796 source.n260 source.n154 0.388379
R797 source.n259 source.n258 0.388379
R798 source.n215 source.n214 0.388379
R799 source.n181 source.n179 0.388379
R800 source source.n576 0.188
R801 source.n482 source.n477 0.155672
R802 source.n489 source.n477 0.155672
R803 source.n490 source.n489 0.155672
R804 source.n490 source.n473 0.155672
R805 source.n497 source.n473 0.155672
R806 source.n498 source.n497 0.155672
R807 source.n498 source.n469 0.155672
R808 source.n507 source.n469 0.155672
R809 source.n508 source.n507 0.155672
R810 source.n508 source.n465 0.155672
R811 source.n515 source.n465 0.155672
R812 source.n516 source.n515 0.155672
R813 source.n516 source.n461 0.155672
R814 source.n523 source.n461 0.155672
R815 source.n524 source.n523 0.155672
R816 source.n524 source.n457 0.155672
R817 source.n531 source.n457 0.155672
R818 source.n532 source.n531 0.155672
R819 source.n532 source.n453 0.155672
R820 source.n539 source.n453 0.155672
R821 source.n540 source.n539 0.155672
R822 source.n540 source.n449 0.155672
R823 source.n548 source.n449 0.155672
R824 source.n549 source.n548 0.155672
R825 source.n549 source.n445 0.155672
R826 source.n557 source.n445 0.155672
R827 source.n558 source.n557 0.155672
R828 source.n558 source.n441 0.155672
R829 source.n565 source.n441 0.155672
R830 source.n566 source.n565 0.155672
R831 source.n566 source.n437 0.155672
R832 source.n573 source.n437 0.155672
R833 source.n338 source.n333 0.155672
R834 source.n345 source.n333 0.155672
R835 source.n346 source.n345 0.155672
R836 source.n346 source.n329 0.155672
R837 source.n353 source.n329 0.155672
R838 source.n354 source.n353 0.155672
R839 source.n354 source.n325 0.155672
R840 source.n363 source.n325 0.155672
R841 source.n364 source.n363 0.155672
R842 source.n364 source.n321 0.155672
R843 source.n371 source.n321 0.155672
R844 source.n372 source.n371 0.155672
R845 source.n372 source.n317 0.155672
R846 source.n379 source.n317 0.155672
R847 source.n380 source.n379 0.155672
R848 source.n380 source.n313 0.155672
R849 source.n387 source.n313 0.155672
R850 source.n388 source.n387 0.155672
R851 source.n388 source.n309 0.155672
R852 source.n395 source.n309 0.155672
R853 source.n396 source.n395 0.155672
R854 source.n396 source.n305 0.155672
R855 source.n404 source.n305 0.155672
R856 source.n405 source.n404 0.155672
R857 source.n405 source.n301 0.155672
R858 source.n413 source.n301 0.155672
R859 source.n414 source.n413 0.155672
R860 source.n414 source.n297 0.155672
R861 source.n421 source.n297 0.155672
R862 source.n422 source.n421 0.155672
R863 source.n422 source.n293 0.155672
R864 source.n429 source.n293 0.155672
R865 source.n137 source.n1 0.155672
R866 source.n130 source.n1 0.155672
R867 source.n130 source.n129 0.155672
R868 source.n129 source.n5 0.155672
R869 source.n122 source.n5 0.155672
R870 source.n122 source.n121 0.155672
R871 source.n121 source.n9 0.155672
R872 source.n113 source.n9 0.155672
R873 source.n113 source.n112 0.155672
R874 source.n112 source.n13 0.155672
R875 source.n105 source.n13 0.155672
R876 source.n105 source.n104 0.155672
R877 source.n104 source.n18 0.155672
R878 source.n97 source.n18 0.155672
R879 source.n97 source.n96 0.155672
R880 source.n96 source.n22 0.155672
R881 source.n89 source.n22 0.155672
R882 source.n89 source.n88 0.155672
R883 source.n88 source.n26 0.155672
R884 source.n81 source.n26 0.155672
R885 source.n81 source.n80 0.155672
R886 source.n80 source.n30 0.155672
R887 source.n73 source.n30 0.155672
R888 source.n73 source.n72 0.155672
R889 source.n72 source.n34 0.155672
R890 source.n64 source.n34 0.155672
R891 source.n64 source.n63 0.155672
R892 source.n63 source.n39 0.155672
R893 source.n56 source.n39 0.155672
R894 source.n56 source.n55 0.155672
R895 source.n55 source.n43 0.155672
R896 source.n48 source.n43 0.155672
R897 source.n281 source.n145 0.155672
R898 source.n274 source.n145 0.155672
R899 source.n274 source.n273 0.155672
R900 source.n273 source.n149 0.155672
R901 source.n266 source.n149 0.155672
R902 source.n266 source.n265 0.155672
R903 source.n265 source.n153 0.155672
R904 source.n257 source.n153 0.155672
R905 source.n257 source.n256 0.155672
R906 source.n256 source.n157 0.155672
R907 source.n249 source.n157 0.155672
R908 source.n249 source.n248 0.155672
R909 source.n248 source.n162 0.155672
R910 source.n241 source.n162 0.155672
R911 source.n241 source.n240 0.155672
R912 source.n240 source.n166 0.155672
R913 source.n233 source.n166 0.155672
R914 source.n233 source.n232 0.155672
R915 source.n232 source.n170 0.155672
R916 source.n225 source.n170 0.155672
R917 source.n225 source.n224 0.155672
R918 source.n224 source.n174 0.155672
R919 source.n217 source.n174 0.155672
R920 source.n217 source.n216 0.155672
R921 source.n216 source.n178 0.155672
R922 source.n208 source.n178 0.155672
R923 source.n208 source.n207 0.155672
R924 source.n207 source.n183 0.155672
R925 source.n200 source.n183 0.155672
R926 source.n200 source.n199 0.155672
R927 source.n199 source.n187 0.155672
R928 source.n192 source.n187 0.155672
R929 drain_right.n134 drain_right.n0 289.615
R930 drain_right.n280 drain_right.n146 289.615
R931 drain_right.n44 drain_right.n43 185
R932 drain_right.n49 drain_right.n48 185
R933 drain_right.n51 drain_right.n50 185
R934 drain_right.n40 drain_right.n39 185
R935 drain_right.n57 drain_right.n56 185
R936 drain_right.n59 drain_right.n58 185
R937 drain_right.n36 drain_right.n35 185
R938 drain_right.n66 drain_right.n65 185
R939 drain_right.n67 drain_right.n34 185
R940 drain_right.n69 drain_right.n68 185
R941 drain_right.n32 drain_right.n31 185
R942 drain_right.n75 drain_right.n74 185
R943 drain_right.n77 drain_right.n76 185
R944 drain_right.n28 drain_right.n27 185
R945 drain_right.n83 drain_right.n82 185
R946 drain_right.n85 drain_right.n84 185
R947 drain_right.n24 drain_right.n23 185
R948 drain_right.n91 drain_right.n90 185
R949 drain_right.n93 drain_right.n92 185
R950 drain_right.n20 drain_right.n19 185
R951 drain_right.n99 drain_right.n98 185
R952 drain_right.n101 drain_right.n100 185
R953 drain_right.n16 drain_right.n15 185
R954 drain_right.n107 drain_right.n106 185
R955 drain_right.n110 drain_right.n109 185
R956 drain_right.n108 drain_right.n12 185
R957 drain_right.n115 drain_right.n11 185
R958 drain_right.n117 drain_right.n116 185
R959 drain_right.n119 drain_right.n118 185
R960 drain_right.n8 drain_right.n7 185
R961 drain_right.n125 drain_right.n124 185
R962 drain_right.n127 drain_right.n126 185
R963 drain_right.n4 drain_right.n3 185
R964 drain_right.n133 drain_right.n132 185
R965 drain_right.n135 drain_right.n134 185
R966 drain_right.n281 drain_right.n280 185
R967 drain_right.n279 drain_right.n278 185
R968 drain_right.n150 drain_right.n149 185
R969 drain_right.n273 drain_right.n272 185
R970 drain_right.n271 drain_right.n270 185
R971 drain_right.n154 drain_right.n153 185
R972 drain_right.n265 drain_right.n264 185
R973 drain_right.n263 drain_right.n262 185
R974 drain_right.n261 drain_right.n157 185
R975 drain_right.n161 drain_right.n158 185
R976 drain_right.n256 drain_right.n255 185
R977 drain_right.n254 drain_right.n253 185
R978 drain_right.n163 drain_right.n162 185
R979 drain_right.n248 drain_right.n247 185
R980 drain_right.n246 drain_right.n245 185
R981 drain_right.n167 drain_right.n166 185
R982 drain_right.n240 drain_right.n239 185
R983 drain_right.n238 drain_right.n237 185
R984 drain_right.n171 drain_right.n170 185
R985 drain_right.n232 drain_right.n231 185
R986 drain_right.n230 drain_right.n229 185
R987 drain_right.n175 drain_right.n174 185
R988 drain_right.n224 drain_right.n223 185
R989 drain_right.n222 drain_right.n221 185
R990 drain_right.n179 drain_right.n178 185
R991 drain_right.n216 drain_right.n215 185
R992 drain_right.n214 drain_right.n181 185
R993 drain_right.n213 drain_right.n212 185
R994 drain_right.n184 drain_right.n182 185
R995 drain_right.n207 drain_right.n206 185
R996 drain_right.n205 drain_right.n204 185
R997 drain_right.n188 drain_right.n187 185
R998 drain_right.n199 drain_right.n198 185
R999 drain_right.n197 drain_right.n196 185
R1000 drain_right.n192 drain_right.n191 185
R1001 drain_right.n45 drain_right.t4 149.524
R1002 drain_right.n193 drain_right.t3 149.524
R1003 drain_right.n49 drain_right.n43 104.615
R1004 drain_right.n50 drain_right.n49 104.615
R1005 drain_right.n50 drain_right.n39 104.615
R1006 drain_right.n57 drain_right.n39 104.615
R1007 drain_right.n58 drain_right.n57 104.615
R1008 drain_right.n58 drain_right.n35 104.615
R1009 drain_right.n66 drain_right.n35 104.615
R1010 drain_right.n67 drain_right.n66 104.615
R1011 drain_right.n68 drain_right.n67 104.615
R1012 drain_right.n68 drain_right.n31 104.615
R1013 drain_right.n75 drain_right.n31 104.615
R1014 drain_right.n76 drain_right.n75 104.615
R1015 drain_right.n76 drain_right.n27 104.615
R1016 drain_right.n83 drain_right.n27 104.615
R1017 drain_right.n84 drain_right.n83 104.615
R1018 drain_right.n84 drain_right.n23 104.615
R1019 drain_right.n91 drain_right.n23 104.615
R1020 drain_right.n92 drain_right.n91 104.615
R1021 drain_right.n92 drain_right.n19 104.615
R1022 drain_right.n99 drain_right.n19 104.615
R1023 drain_right.n100 drain_right.n99 104.615
R1024 drain_right.n100 drain_right.n15 104.615
R1025 drain_right.n107 drain_right.n15 104.615
R1026 drain_right.n109 drain_right.n107 104.615
R1027 drain_right.n109 drain_right.n108 104.615
R1028 drain_right.n108 drain_right.n11 104.615
R1029 drain_right.n117 drain_right.n11 104.615
R1030 drain_right.n118 drain_right.n117 104.615
R1031 drain_right.n118 drain_right.n7 104.615
R1032 drain_right.n125 drain_right.n7 104.615
R1033 drain_right.n126 drain_right.n125 104.615
R1034 drain_right.n126 drain_right.n3 104.615
R1035 drain_right.n133 drain_right.n3 104.615
R1036 drain_right.n134 drain_right.n133 104.615
R1037 drain_right.n280 drain_right.n279 104.615
R1038 drain_right.n279 drain_right.n149 104.615
R1039 drain_right.n272 drain_right.n149 104.615
R1040 drain_right.n272 drain_right.n271 104.615
R1041 drain_right.n271 drain_right.n153 104.615
R1042 drain_right.n264 drain_right.n153 104.615
R1043 drain_right.n264 drain_right.n263 104.615
R1044 drain_right.n263 drain_right.n157 104.615
R1045 drain_right.n161 drain_right.n157 104.615
R1046 drain_right.n255 drain_right.n161 104.615
R1047 drain_right.n255 drain_right.n254 104.615
R1048 drain_right.n254 drain_right.n162 104.615
R1049 drain_right.n247 drain_right.n162 104.615
R1050 drain_right.n247 drain_right.n246 104.615
R1051 drain_right.n246 drain_right.n166 104.615
R1052 drain_right.n239 drain_right.n166 104.615
R1053 drain_right.n239 drain_right.n238 104.615
R1054 drain_right.n238 drain_right.n170 104.615
R1055 drain_right.n231 drain_right.n170 104.615
R1056 drain_right.n231 drain_right.n230 104.615
R1057 drain_right.n230 drain_right.n174 104.615
R1058 drain_right.n223 drain_right.n174 104.615
R1059 drain_right.n223 drain_right.n222 104.615
R1060 drain_right.n222 drain_right.n178 104.615
R1061 drain_right.n215 drain_right.n178 104.615
R1062 drain_right.n215 drain_right.n214 104.615
R1063 drain_right.n214 drain_right.n213 104.615
R1064 drain_right.n213 drain_right.n182 104.615
R1065 drain_right.n206 drain_right.n182 104.615
R1066 drain_right.n206 drain_right.n205 104.615
R1067 drain_right.n205 drain_right.n187 104.615
R1068 drain_right.n198 drain_right.n187 104.615
R1069 drain_right.n198 drain_right.n197 104.615
R1070 drain_right.n197 drain_right.n191 104.615
R1071 drain_right.n145 drain_right.n143 59.6032
R1072 drain_right.n142 drain_right.n141 59.326
R1073 drain_right.n140 drain_right.n139 58.7154
R1074 drain_right.n145 drain_right.n144 58.7154
R1075 drain_right.t4 drain_right.n43 52.3082
R1076 drain_right.t3 drain_right.n191 52.3082
R1077 drain_right.n140 drain_right.n138 48.2006
R1078 drain_right.n285 drain_right.n284 47.3126
R1079 drain_right drain_right.n142 40.436
R1080 drain_right.n69 drain_right.n34 13.1884
R1081 drain_right.n116 drain_right.n115 13.1884
R1082 drain_right.n262 drain_right.n261 13.1884
R1083 drain_right.n216 drain_right.n181 13.1884
R1084 drain_right.n65 drain_right.n64 12.8005
R1085 drain_right.n70 drain_right.n32 12.8005
R1086 drain_right.n114 drain_right.n12 12.8005
R1087 drain_right.n119 drain_right.n10 12.8005
R1088 drain_right.n265 drain_right.n156 12.8005
R1089 drain_right.n260 drain_right.n158 12.8005
R1090 drain_right.n217 drain_right.n179 12.8005
R1091 drain_right.n212 drain_right.n183 12.8005
R1092 drain_right.n63 drain_right.n36 12.0247
R1093 drain_right.n74 drain_right.n73 12.0247
R1094 drain_right.n111 drain_right.n110 12.0247
R1095 drain_right.n120 drain_right.n8 12.0247
R1096 drain_right.n266 drain_right.n154 12.0247
R1097 drain_right.n257 drain_right.n256 12.0247
R1098 drain_right.n221 drain_right.n220 12.0247
R1099 drain_right.n211 drain_right.n184 12.0247
R1100 drain_right.n60 drain_right.n59 11.249
R1101 drain_right.n77 drain_right.n30 11.249
R1102 drain_right.n106 drain_right.n14 11.249
R1103 drain_right.n124 drain_right.n123 11.249
R1104 drain_right.n270 drain_right.n269 11.249
R1105 drain_right.n253 drain_right.n160 11.249
R1106 drain_right.n224 drain_right.n177 11.249
R1107 drain_right.n208 drain_right.n207 11.249
R1108 drain_right.n56 drain_right.n38 10.4732
R1109 drain_right.n78 drain_right.n28 10.4732
R1110 drain_right.n105 drain_right.n16 10.4732
R1111 drain_right.n127 drain_right.n6 10.4732
R1112 drain_right.n273 drain_right.n152 10.4732
R1113 drain_right.n252 drain_right.n163 10.4732
R1114 drain_right.n225 drain_right.n175 10.4732
R1115 drain_right.n204 drain_right.n186 10.4732
R1116 drain_right.n45 drain_right.n44 10.2747
R1117 drain_right.n193 drain_right.n192 10.2747
R1118 drain_right.n55 drain_right.n40 9.69747
R1119 drain_right.n82 drain_right.n81 9.69747
R1120 drain_right.n102 drain_right.n101 9.69747
R1121 drain_right.n128 drain_right.n4 9.69747
R1122 drain_right.n274 drain_right.n150 9.69747
R1123 drain_right.n249 drain_right.n248 9.69747
R1124 drain_right.n229 drain_right.n228 9.69747
R1125 drain_right.n203 drain_right.n188 9.69747
R1126 drain_right.n138 drain_right.n137 9.45567
R1127 drain_right.n284 drain_right.n283 9.45567
R1128 drain_right.n2 drain_right.n1 9.3005
R1129 drain_right.n131 drain_right.n130 9.3005
R1130 drain_right.n129 drain_right.n128 9.3005
R1131 drain_right.n6 drain_right.n5 9.3005
R1132 drain_right.n123 drain_right.n122 9.3005
R1133 drain_right.n121 drain_right.n120 9.3005
R1134 drain_right.n10 drain_right.n9 9.3005
R1135 drain_right.n89 drain_right.n88 9.3005
R1136 drain_right.n87 drain_right.n86 9.3005
R1137 drain_right.n26 drain_right.n25 9.3005
R1138 drain_right.n81 drain_right.n80 9.3005
R1139 drain_right.n79 drain_right.n78 9.3005
R1140 drain_right.n30 drain_right.n29 9.3005
R1141 drain_right.n73 drain_right.n72 9.3005
R1142 drain_right.n71 drain_right.n70 9.3005
R1143 drain_right.n47 drain_right.n46 9.3005
R1144 drain_right.n42 drain_right.n41 9.3005
R1145 drain_right.n53 drain_right.n52 9.3005
R1146 drain_right.n55 drain_right.n54 9.3005
R1147 drain_right.n38 drain_right.n37 9.3005
R1148 drain_right.n61 drain_right.n60 9.3005
R1149 drain_right.n63 drain_right.n62 9.3005
R1150 drain_right.n64 drain_right.n33 9.3005
R1151 drain_right.n22 drain_right.n21 9.3005
R1152 drain_right.n95 drain_right.n94 9.3005
R1153 drain_right.n97 drain_right.n96 9.3005
R1154 drain_right.n18 drain_right.n17 9.3005
R1155 drain_right.n103 drain_right.n102 9.3005
R1156 drain_right.n105 drain_right.n104 9.3005
R1157 drain_right.n14 drain_right.n13 9.3005
R1158 drain_right.n112 drain_right.n111 9.3005
R1159 drain_right.n114 drain_right.n113 9.3005
R1160 drain_right.n137 drain_right.n136 9.3005
R1161 drain_right.n195 drain_right.n194 9.3005
R1162 drain_right.n190 drain_right.n189 9.3005
R1163 drain_right.n201 drain_right.n200 9.3005
R1164 drain_right.n203 drain_right.n202 9.3005
R1165 drain_right.n186 drain_right.n185 9.3005
R1166 drain_right.n209 drain_right.n208 9.3005
R1167 drain_right.n211 drain_right.n210 9.3005
R1168 drain_right.n183 drain_right.n180 9.3005
R1169 drain_right.n242 drain_right.n241 9.3005
R1170 drain_right.n244 drain_right.n243 9.3005
R1171 drain_right.n165 drain_right.n164 9.3005
R1172 drain_right.n250 drain_right.n249 9.3005
R1173 drain_right.n252 drain_right.n251 9.3005
R1174 drain_right.n160 drain_right.n159 9.3005
R1175 drain_right.n258 drain_right.n257 9.3005
R1176 drain_right.n260 drain_right.n259 9.3005
R1177 drain_right.n283 drain_right.n282 9.3005
R1178 drain_right.n148 drain_right.n147 9.3005
R1179 drain_right.n277 drain_right.n276 9.3005
R1180 drain_right.n275 drain_right.n274 9.3005
R1181 drain_right.n152 drain_right.n151 9.3005
R1182 drain_right.n269 drain_right.n268 9.3005
R1183 drain_right.n267 drain_right.n266 9.3005
R1184 drain_right.n156 drain_right.n155 9.3005
R1185 drain_right.n169 drain_right.n168 9.3005
R1186 drain_right.n236 drain_right.n235 9.3005
R1187 drain_right.n234 drain_right.n233 9.3005
R1188 drain_right.n173 drain_right.n172 9.3005
R1189 drain_right.n228 drain_right.n227 9.3005
R1190 drain_right.n226 drain_right.n225 9.3005
R1191 drain_right.n177 drain_right.n176 9.3005
R1192 drain_right.n220 drain_right.n219 9.3005
R1193 drain_right.n218 drain_right.n217 9.3005
R1194 drain_right.n52 drain_right.n51 8.92171
R1195 drain_right.n85 drain_right.n26 8.92171
R1196 drain_right.n98 drain_right.n18 8.92171
R1197 drain_right.n132 drain_right.n131 8.92171
R1198 drain_right.n278 drain_right.n277 8.92171
R1199 drain_right.n245 drain_right.n165 8.92171
R1200 drain_right.n232 drain_right.n173 8.92171
R1201 drain_right.n200 drain_right.n199 8.92171
R1202 drain_right.n48 drain_right.n42 8.14595
R1203 drain_right.n86 drain_right.n24 8.14595
R1204 drain_right.n97 drain_right.n20 8.14595
R1205 drain_right.n135 drain_right.n2 8.14595
R1206 drain_right.n281 drain_right.n148 8.14595
R1207 drain_right.n244 drain_right.n167 8.14595
R1208 drain_right.n233 drain_right.n171 8.14595
R1209 drain_right.n196 drain_right.n190 8.14595
R1210 drain_right.n47 drain_right.n44 7.3702
R1211 drain_right.n90 drain_right.n89 7.3702
R1212 drain_right.n94 drain_right.n93 7.3702
R1213 drain_right.n136 drain_right.n0 7.3702
R1214 drain_right.n282 drain_right.n146 7.3702
R1215 drain_right.n241 drain_right.n240 7.3702
R1216 drain_right.n237 drain_right.n236 7.3702
R1217 drain_right.n195 drain_right.n192 7.3702
R1218 drain_right.n90 drain_right.n22 6.59444
R1219 drain_right.n93 drain_right.n22 6.59444
R1220 drain_right.n138 drain_right.n0 6.59444
R1221 drain_right.n284 drain_right.n146 6.59444
R1222 drain_right.n240 drain_right.n169 6.59444
R1223 drain_right.n237 drain_right.n169 6.59444
R1224 drain_right drain_right.n285 6.09718
R1225 drain_right.n48 drain_right.n47 5.81868
R1226 drain_right.n89 drain_right.n24 5.81868
R1227 drain_right.n94 drain_right.n20 5.81868
R1228 drain_right.n136 drain_right.n135 5.81868
R1229 drain_right.n282 drain_right.n281 5.81868
R1230 drain_right.n241 drain_right.n167 5.81868
R1231 drain_right.n236 drain_right.n171 5.81868
R1232 drain_right.n196 drain_right.n195 5.81868
R1233 drain_right.n51 drain_right.n42 5.04292
R1234 drain_right.n86 drain_right.n85 5.04292
R1235 drain_right.n98 drain_right.n97 5.04292
R1236 drain_right.n132 drain_right.n2 5.04292
R1237 drain_right.n278 drain_right.n148 5.04292
R1238 drain_right.n245 drain_right.n244 5.04292
R1239 drain_right.n233 drain_right.n232 5.04292
R1240 drain_right.n199 drain_right.n190 5.04292
R1241 drain_right.n52 drain_right.n40 4.26717
R1242 drain_right.n82 drain_right.n26 4.26717
R1243 drain_right.n101 drain_right.n18 4.26717
R1244 drain_right.n131 drain_right.n4 4.26717
R1245 drain_right.n277 drain_right.n150 4.26717
R1246 drain_right.n248 drain_right.n165 4.26717
R1247 drain_right.n229 drain_right.n173 4.26717
R1248 drain_right.n200 drain_right.n188 4.26717
R1249 drain_right.n56 drain_right.n55 3.49141
R1250 drain_right.n81 drain_right.n28 3.49141
R1251 drain_right.n102 drain_right.n16 3.49141
R1252 drain_right.n128 drain_right.n127 3.49141
R1253 drain_right.n274 drain_right.n273 3.49141
R1254 drain_right.n249 drain_right.n163 3.49141
R1255 drain_right.n228 drain_right.n175 3.49141
R1256 drain_right.n204 drain_right.n203 3.49141
R1257 drain_right.n194 drain_right.n193 2.84303
R1258 drain_right.n46 drain_right.n45 2.84303
R1259 drain_right.n59 drain_right.n38 2.71565
R1260 drain_right.n78 drain_right.n77 2.71565
R1261 drain_right.n106 drain_right.n105 2.71565
R1262 drain_right.n124 drain_right.n6 2.71565
R1263 drain_right.n270 drain_right.n152 2.71565
R1264 drain_right.n253 drain_right.n252 2.71565
R1265 drain_right.n225 drain_right.n224 2.71565
R1266 drain_right.n207 drain_right.n186 2.71565
R1267 drain_right.n60 drain_right.n36 1.93989
R1268 drain_right.n74 drain_right.n30 1.93989
R1269 drain_right.n110 drain_right.n14 1.93989
R1270 drain_right.n123 drain_right.n8 1.93989
R1271 drain_right.n269 drain_right.n154 1.93989
R1272 drain_right.n256 drain_right.n160 1.93989
R1273 drain_right.n221 drain_right.n177 1.93989
R1274 drain_right.n208 drain_right.n184 1.93989
R1275 drain_right.n65 drain_right.n63 1.16414
R1276 drain_right.n73 drain_right.n32 1.16414
R1277 drain_right.n111 drain_right.n12 1.16414
R1278 drain_right.n120 drain_right.n119 1.16414
R1279 drain_right.n266 drain_right.n265 1.16414
R1280 drain_right.n257 drain_right.n158 1.16414
R1281 drain_right.n220 drain_right.n179 1.16414
R1282 drain_right.n212 drain_right.n211 1.16414
R1283 drain_right.n285 drain_right.n145 0.888431
R1284 drain_right.n141 drain_right.t8 0.7925
R1285 drain_right.n141 drain_right.t6 0.7925
R1286 drain_right.n139 drain_right.t5 0.7925
R1287 drain_right.n139 drain_right.t9 0.7925
R1288 drain_right.n143 drain_right.t7 0.7925
R1289 drain_right.n143 drain_right.t1 0.7925
R1290 drain_right.n144 drain_right.t0 0.7925
R1291 drain_right.n144 drain_right.t2 0.7925
R1292 drain_right.n64 drain_right.n34 0.388379
R1293 drain_right.n70 drain_right.n69 0.388379
R1294 drain_right.n115 drain_right.n114 0.388379
R1295 drain_right.n116 drain_right.n10 0.388379
R1296 drain_right.n262 drain_right.n156 0.388379
R1297 drain_right.n261 drain_right.n260 0.388379
R1298 drain_right.n217 drain_right.n216 0.388379
R1299 drain_right.n183 drain_right.n181 0.388379
R1300 drain_right.n142 drain_right.n140 0.167137
R1301 drain_right.n46 drain_right.n41 0.155672
R1302 drain_right.n53 drain_right.n41 0.155672
R1303 drain_right.n54 drain_right.n53 0.155672
R1304 drain_right.n54 drain_right.n37 0.155672
R1305 drain_right.n61 drain_right.n37 0.155672
R1306 drain_right.n62 drain_right.n61 0.155672
R1307 drain_right.n62 drain_right.n33 0.155672
R1308 drain_right.n71 drain_right.n33 0.155672
R1309 drain_right.n72 drain_right.n71 0.155672
R1310 drain_right.n72 drain_right.n29 0.155672
R1311 drain_right.n79 drain_right.n29 0.155672
R1312 drain_right.n80 drain_right.n79 0.155672
R1313 drain_right.n80 drain_right.n25 0.155672
R1314 drain_right.n87 drain_right.n25 0.155672
R1315 drain_right.n88 drain_right.n87 0.155672
R1316 drain_right.n88 drain_right.n21 0.155672
R1317 drain_right.n95 drain_right.n21 0.155672
R1318 drain_right.n96 drain_right.n95 0.155672
R1319 drain_right.n96 drain_right.n17 0.155672
R1320 drain_right.n103 drain_right.n17 0.155672
R1321 drain_right.n104 drain_right.n103 0.155672
R1322 drain_right.n104 drain_right.n13 0.155672
R1323 drain_right.n112 drain_right.n13 0.155672
R1324 drain_right.n113 drain_right.n112 0.155672
R1325 drain_right.n113 drain_right.n9 0.155672
R1326 drain_right.n121 drain_right.n9 0.155672
R1327 drain_right.n122 drain_right.n121 0.155672
R1328 drain_right.n122 drain_right.n5 0.155672
R1329 drain_right.n129 drain_right.n5 0.155672
R1330 drain_right.n130 drain_right.n129 0.155672
R1331 drain_right.n130 drain_right.n1 0.155672
R1332 drain_right.n137 drain_right.n1 0.155672
R1333 drain_right.n283 drain_right.n147 0.155672
R1334 drain_right.n276 drain_right.n147 0.155672
R1335 drain_right.n276 drain_right.n275 0.155672
R1336 drain_right.n275 drain_right.n151 0.155672
R1337 drain_right.n268 drain_right.n151 0.155672
R1338 drain_right.n268 drain_right.n267 0.155672
R1339 drain_right.n267 drain_right.n155 0.155672
R1340 drain_right.n259 drain_right.n155 0.155672
R1341 drain_right.n259 drain_right.n258 0.155672
R1342 drain_right.n258 drain_right.n159 0.155672
R1343 drain_right.n251 drain_right.n159 0.155672
R1344 drain_right.n251 drain_right.n250 0.155672
R1345 drain_right.n250 drain_right.n164 0.155672
R1346 drain_right.n243 drain_right.n164 0.155672
R1347 drain_right.n243 drain_right.n242 0.155672
R1348 drain_right.n242 drain_right.n168 0.155672
R1349 drain_right.n235 drain_right.n168 0.155672
R1350 drain_right.n235 drain_right.n234 0.155672
R1351 drain_right.n234 drain_right.n172 0.155672
R1352 drain_right.n227 drain_right.n172 0.155672
R1353 drain_right.n227 drain_right.n226 0.155672
R1354 drain_right.n226 drain_right.n176 0.155672
R1355 drain_right.n219 drain_right.n176 0.155672
R1356 drain_right.n219 drain_right.n218 0.155672
R1357 drain_right.n218 drain_right.n180 0.155672
R1358 drain_right.n210 drain_right.n180 0.155672
R1359 drain_right.n210 drain_right.n209 0.155672
R1360 drain_right.n209 drain_right.n185 0.155672
R1361 drain_right.n202 drain_right.n185 0.155672
R1362 drain_right.n202 drain_right.n201 0.155672
R1363 drain_right.n201 drain_right.n189 0.155672
R1364 drain_right.n194 drain_right.n189 0.155672
R1365 plus.n3 plus.t3 939.582
R1366 plus.n17 plus.t9 939.582
R1367 plus.n12 plus.t2 916.833
R1368 plus.n10 plus.t5 916.833
R1369 plus.n2 plus.t1 916.833
R1370 plus.n4 plus.t7 916.833
R1371 plus.n26 plus.t6 916.833
R1372 plus.n24 plus.t4 916.833
R1373 plus.n16 plus.t8 916.833
R1374 plus.n18 plus.t0 916.833
R1375 plus.n6 plus.n5 161.3
R1376 plus.n7 plus.n2 161.3
R1377 plus.n9 plus.n8 161.3
R1378 plus.n10 plus.n1 161.3
R1379 plus.n11 plus.n0 161.3
R1380 plus.n13 plus.n12 161.3
R1381 plus.n20 plus.n19 161.3
R1382 plus.n21 plus.n16 161.3
R1383 plus.n23 plus.n22 161.3
R1384 plus.n24 plus.n15 161.3
R1385 plus.n25 plus.n14 161.3
R1386 plus.n27 plus.n26 161.3
R1387 plus.n6 plus.n3 44.8741
R1388 plus.n20 plus.n17 44.8741
R1389 plus plus.n27 35.4593
R1390 plus.n12 plus.n11 30.6732
R1391 plus.n26 plus.n25 30.6732
R1392 plus.n10 plus.n9 26.2914
R1393 plus.n5 plus.n4 26.2914
R1394 plus.n24 plus.n23 26.2914
R1395 plus.n19 plus.n18 26.2914
R1396 plus.n9 plus.n2 21.9096
R1397 plus.n5 plus.n2 21.9096
R1398 plus.n23 plus.n16 21.9096
R1399 plus.n19 plus.n16 21.9096
R1400 plus.n4 plus.n3 19.0667
R1401 plus.n18 plus.n17 19.0667
R1402 plus.n11 plus.n10 17.5278
R1403 plus.n25 plus.n24 17.5278
R1404 plus plus.n13 17.2069
R1405 plus.n7 plus.n6 0.189894
R1406 plus.n8 plus.n7 0.189894
R1407 plus.n8 plus.n1 0.189894
R1408 plus.n1 plus.n0 0.189894
R1409 plus.n13 plus.n0 0.189894
R1410 plus.n27 plus.n14 0.189894
R1411 plus.n15 plus.n14 0.189894
R1412 plus.n22 plus.n15 0.189894
R1413 plus.n22 plus.n21 0.189894
R1414 plus.n21 plus.n20 0.189894
R1415 drain_left.n134 drain_left.n0 289.615
R1416 drain_left.n277 drain_left.n143 289.615
R1417 drain_left.n44 drain_left.n43 185
R1418 drain_left.n49 drain_left.n48 185
R1419 drain_left.n51 drain_left.n50 185
R1420 drain_left.n40 drain_left.n39 185
R1421 drain_left.n57 drain_left.n56 185
R1422 drain_left.n59 drain_left.n58 185
R1423 drain_left.n36 drain_left.n35 185
R1424 drain_left.n66 drain_left.n65 185
R1425 drain_left.n67 drain_left.n34 185
R1426 drain_left.n69 drain_left.n68 185
R1427 drain_left.n32 drain_left.n31 185
R1428 drain_left.n75 drain_left.n74 185
R1429 drain_left.n77 drain_left.n76 185
R1430 drain_left.n28 drain_left.n27 185
R1431 drain_left.n83 drain_left.n82 185
R1432 drain_left.n85 drain_left.n84 185
R1433 drain_left.n24 drain_left.n23 185
R1434 drain_left.n91 drain_left.n90 185
R1435 drain_left.n93 drain_left.n92 185
R1436 drain_left.n20 drain_left.n19 185
R1437 drain_left.n99 drain_left.n98 185
R1438 drain_left.n101 drain_left.n100 185
R1439 drain_left.n16 drain_left.n15 185
R1440 drain_left.n107 drain_left.n106 185
R1441 drain_left.n110 drain_left.n109 185
R1442 drain_left.n108 drain_left.n12 185
R1443 drain_left.n115 drain_left.n11 185
R1444 drain_left.n117 drain_left.n116 185
R1445 drain_left.n119 drain_left.n118 185
R1446 drain_left.n8 drain_left.n7 185
R1447 drain_left.n125 drain_left.n124 185
R1448 drain_left.n127 drain_left.n126 185
R1449 drain_left.n4 drain_left.n3 185
R1450 drain_left.n133 drain_left.n132 185
R1451 drain_left.n135 drain_left.n134 185
R1452 drain_left.n278 drain_left.n277 185
R1453 drain_left.n276 drain_left.n275 185
R1454 drain_left.n147 drain_left.n146 185
R1455 drain_left.n270 drain_left.n269 185
R1456 drain_left.n268 drain_left.n267 185
R1457 drain_left.n151 drain_left.n150 185
R1458 drain_left.n262 drain_left.n261 185
R1459 drain_left.n260 drain_left.n259 185
R1460 drain_left.n258 drain_left.n154 185
R1461 drain_left.n158 drain_left.n155 185
R1462 drain_left.n253 drain_left.n252 185
R1463 drain_left.n251 drain_left.n250 185
R1464 drain_left.n160 drain_left.n159 185
R1465 drain_left.n245 drain_left.n244 185
R1466 drain_left.n243 drain_left.n242 185
R1467 drain_left.n164 drain_left.n163 185
R1468 drain_left.n237 drain_left.n236 185
R1469 drain_left.n235 drain_left.n234 185
R1470 drain_left.n168 drain_left.n167 185
R1471 drain_left.n229 drain_left.n228 185
R1472 drain_left.n227 drain_left.n226 185
R1473 drain_left.n172 drain_left.n171 185
R1474 drain_left.n221 drain_left.n220 185
R1475 drain_left.n219 drain_left.n218 185
R1476 drain_left.n176 drain_left.n175 185
R1477 drain_left.n213 drain_left.n212 185
R1478 drain_left.n211 drain_left.n178 185
R1479 drain_left.n210 drain_left.n209 185
R1480 drain_left.n181 drain_left.n179 185
R1481 drain_left.n204 drain_left.n203 185
R1482 drain_left.n202 drain_left.n201 185
R1483 drain_left.n185 drain_left.n184 185
R1484 drain_left.n196 drain_left.n195 185
R1485 drain_left.n194 drain_left.n193 185
R1486 drain_left.n189 drain_left.n188 185
R1487 drain_left.n45 drain_left.t3 149.524
R1488 drain_left.n190 drain_left.t6 149.524
R1489 drain_left.n49 drain_left.n43 104.615
R1490 drain_left.n50 drain_left.n49 104.615
R1491 drain_left.n50 drain_left.n39 104.615
R1492 drain_left.n57 drain_left.n39 104.615
R1493 drain_left.n58 drain_left.n57 104.615
R1494 drain_left.n58 drain_left.n35 104.615
R1495 drain_left.n66 drain_left.n35 104.615
R1496 drain_left.n67 drain_left.n66 104.615
R1497 drain_left.n68 drain_left.n67 104.615
R1498 drain_left.n68 drain_left.n31 104.615
R1499 drain_left.n75 drain_left.n31 104.615
R1500 drain_left.n76 drain_left.n75 104.615
R1501 drain_left.n76 drain_left.n27 104.615
R1502 drain_left.n83 drain_left.n27 104.615
R1503 drain_left.n84 drain_left.n83 104.615
R1504 drain_left.n84 drain_left.n23 104.615
R1505 drain_left.n91 drain_left.n23 104.615
R1506 drain_left.n92 drain_left.n91 104.615
R1507 drain_left.n92 drain_left.n19 104.615
R1508 drain_left.n99 drain_left.n19 104.615
R1509 drain_left.n100 drain_left.n99 104.615
R1510 drain_left.n100 drain_left.n15 104.615
R1511 drain_left.n107 drain_left.n15 104.615
R1512 drain_left.n109 drain_left.n107 104.615
R1513 drain_left.n109 drain_left.n108 104.615
R1514 drain_left.n108 drain_left.n11 104.615
R1515 drain_left.n117 drain_left.n11 104.615
R1516 drain_left.n118 drain_left.n117 104.615
R1517 drain_left.n118 drain_left.n7 104.615
R1518 drain_left.n125 drain_left.n7 104.615
R1519 drain_left.n126 drain_left.n125 104.615
R1520 drain_left.n126 drain_left.n3 104.615
R1521 drain_left.n133 drain_left.n3 104.615
R1522 drain_left.n134 drain_left.n133 104.615
R1523 drain_left.n277 drain_left.n276 104.615
R1524 drain_left.n276 drain_left.n146 104.615
R1525 drain_left.n269 drain_left.n146 104.615
R1526 drain_left.n269 drain_left.n268 104.615
R1527 drain_left.n268 drain_left.n150 104.615
R1528 drain_left.n261 drain_left.n150 104.615
R1529 drain_left.n261 drain_left.n260 104.615
R1530 drain_left.n260 drain_left.n154 104.615
R1531 drain_left.n158 drain_left.n154 104.615
R1532 drain_left.n252 drain_left.n158 104.615
R1533 drain_left.n252 drain_left.n251 104.615
R1534 drain_left.n251 drain_left.n159 104.615
R1535 drain_left.n244 drain_left.n159 104.615
R1536 drain_left.n244 drain_left.n243 104.615
R1537 drain_left.n243 drain_left.n163 104.615
R1538 drain_left.n236 drain_left.n163 104.615
R1539 drain_left.n236 drain_left.n235 104.615
R1540 drain_left.n235 drain_left.n167 104.615
R1541 drain_left.n228 drain_left.n167 104.615
R1542 drain_left.n228 drain_left.n227 104.615
R1543 drain_left.n227 drain_left.n171 104.615
R1544 drain_left.n220 drain_left.n171 104.615
R1545 drain_left.n220 drain_left.n219 104.615
R1546 drain_left.n219 drain_left.n175 104.615
R1547 drain_left.n212 drain_left.n175 104.615
R1548 drain_left.n212 drain_left.n211 104.615
R1549 drain_left.n211 drain_left.n210 104.615
R1550 drain_left.n210 drain_left.n179 104.615
R1551 drain_left.n203 drain_left.n179 104.615
R1552 drain_left.n203 drain_left.n202 104.615
R1553 drain_left.n202 drain_left.n184 104.615
R1554 drain_left.n195 drain_left.n184 104.615
R1555 drain_left.n195 drain_left.n194 104.615
R1556 drain_left.n194 drain_left.n188 104.615
R1557 drain_left.n142 drain_left.n141 59.326
R1558 drain_left.n140 drain_left.n139 58.7154
R1559 drain_left.n283 drain_left.n282 58.7154
R1560 drain_left.n285 drain_left.n284 58.7153
R1561 drain_left.t3 drain_left.n43 52.3082
R1562 drain_left.t6 drain_left.n188 52.3082
R1563 drain_left.n140 drain_left.n138 48.2006
R1564 drain_left.n283 drain_left.n281 48.2006
R1565 drain_left drain_left.n142 40.9893
R1566 drain_left.n69 drain_left.n34 13.1884
R1567 drain_left.n116 drain_left.n115 13.1884
R1568 drain_left.n259 drain_left.n258 13.1884
R1569 drain_left.n213 drain_left.n178 13.1884
R1570 drain_left.n65 drain_left.n64 12.8005
R1571 drain_left.n70 drain_left.n32 12.8005
R1572 drain_left.n114 drain_left.n12 12.8005
R1573 drain_left.n119 drain_left.n10 12.8005
R1574 drain_left.n262 drain_left.n153 12.8005
R1575 drain_left.n257 drain_left.n155 12.8005
R1576 drain_left.n214 drain_left.n176 12.8005
R1577 drain_left.n209 drain_left.n180 12.8005
R1578 drain_left.n63 drain_left.n36 12.0247
R1579 drain_left.n74 drain_left.n73 12.0247
R1580 drain_left.n111 drain_left.n110 12.0247
R1581 drain_left.n120 drain_left.n8 12.0247
R1582 drain_left.n263 drain_left.n151 12.0247
R1583 drain_left.n254 drain_left.n253 12.0247
R1584 drain_left.n218 drain_left.n217 12.0247
R1585 drain_left.n208 drain_left.n181 12.0247
R1586 drain_left.n60 drain_left.n59 11.249
R1587 drain_left.n77 drain_left.n30 11.249
R1588 drain_left.n106 drain_left.n14 11.249
R1589 drain_left.n124 drain_left.n123 11.249
R1590 drain_left.n267 drain_left.n266 11.249
R1591 drain_left.n250 drain_left.n157 11.249
R1592 drain_left.n221 drain_left.n174 11.249
R1593 drain_left.n205 drain_left.n204 11.249
R1594 drain_left.n56 drain_left.n38 10.4732
R1595 drain_left.n78 drain_left.n28 10.4732
R1596 drain_left.n105 drain_left.n16 10.4732
R1597 drain_left.n127 drain_left.n6 10.4732
R1598 drain_left.n270 drain_left.n149 10.4732
R1599 drain_left.n249 drain_left.n160 10.4732
R1600 drain_left.n222 drain_left.n172 10.4732
R1601 drain_left.n201 drain_left.n183 10.4732
R1602 drain_left.n45 drain_left.n44 10.2747
R1603 drain_left.n190 drain_left.n189 10.2747
R1604 drain_left.n55 drain_left.n40 9.69747
R1605 drain_left.n82 drain_left.n81 9.69747
R1606 drain_left.n102 drain_left.n101 9.69747
R1607 drain_left.n128 drain_left.n4 9.69747
R1608 drain_left.n271 drain_left.n147 9.69747
R1609 drain_left.n246 drain_left.n245 9.69747
R1610 drain_left.n226 drain_left.n225 9.69747
R1611 drain_left.n200 drain_left.n185 9.69747
R1612 drain_left.n138 drain_left.n137 9.45567
R1613 drain_left.n281 drain_left.n280 9.45567
R1614 drain_left.n2 drain_left.n1 9.3005
R1615 drain_left.n131 drain_left.n130 9.3005
R1616 drain_left.n129 drain_left.n128 9.3005
R1617 drain_left.n6 drain_left.n5 9.3005
R1618 drain_left.n123 drain_left.n122 9.3005
R1619 drain_left.n121 drain_left.n120 9.3005
R1620 drain_left.n10 drain_left.n9 9.3005
R1621 drain_left.n89 drain_left.n88 9.3005
R1622 drain_left.n87 drain_left.n86 9.3005
R1623 drain_left.n26 drain_left.n25 9.3005
R1624 drain_left.n81 drain_left.n80 9.3005
R1625 drain_left.n79 drain_left.n78 9.3005
R1626 drain_left.n30 drain_left.n29 9.3005
R1627 drain_left.n73 drain_left.n72 9.3005
R1628 drain_left.n71 drain_left.n70 9.3005
R1629 drain_left.n47 drain_left.n46 9.3005
R1630 drain_left.n42 drain_left.n41 9.3005
R1631 drain_left.n53 drain_left.n52 9.3005
R1632 drain_left.n55 drain_left.n54 9.3005
R1633 drain_left.n38 drain_left.n37 9.3005
R1634 drain_left.n61 drain_left.n60 9.3005
R1635 drain_left.n63 drain_left.n62 9.3005
R1636 drain_left.n64 drain_left.n33 9.3005
R1637 drain_left.n22 drain_left.n21 9.3005
R1638 drain_left.n95 drain_left.n94 9.3005
R1639 drain_left.n97 drain_left.n96 9.3005
R1640 drain_left.n18 drain_left.n17 9.3005
R1641 drain_left.n103 drain_left.n102 9.3005
R1642 drain_left.n105 drain_left.n104 9.3005
R1643 drain_left.n14 drain_left.n13 9.3005
R1644 drain_left.n112 drain_left.n111 9.3005
R1645 drain_left.n114 drain_left.n113 9.3005
R1646 drain_left.n137 drain_left.n136 9.3005
R1647 drain_left.n192 drain_left.n191 9.3005
R1648 drain_left.n187 drain_left.n186 9.3005
R1649 drain_left.n198 drain_left.n197 9.3005
R1650 drain_left.n200 drain_left.n199 9.3005
R1651 drain_left.n183 drain_left.n182 9.3005
R1652 drain_left.n206 drain_left.n205 9.3005
R1653 drain_left.n208 drain_left.n207 9.3005
R1654 drain_left.n180 drain_left.n177 9.3005
R1655 drain_left.n239 drain_left.n238 9.3005
R1656 drain_left.n241 drain_left.n240 9.3005
R1657 drain_left.n162 drain_left.n161 9.3005
R1658 drain_left.n247 drain_left.n246 9.3005
R1659 drain_left.n249 drain_left.n248 9.3005
R1660 drain_left.n157 drain_left.n156 9.3005
R1661 drain_left.n255 drain_left.n254 9.3005
R1662 drain_left.n257 drain_left.n256 9.3005
R1663 drain_left.n280 drain_left.n279 9.3005
R1664 drain_left.n145 drain_left.n144 9.3005
R1665 drain_left.n274 drain_left.n273 9.3005
R1666 drain_left.n272 drain_left.n271 9.3005
R1667 drain_left.n149 drain_left.n148 9.3005
R1668 drain_left.n266 drain_left.n265 9.3005
R1669 drain_left.n264 drain_left.n263 9.3005
R1670 drain_left.n153 drain_left.n152 9.3005
R1671 drain_left.n166 drain_left.n165 9.3005
R1672 drain_left.n233 drain_left.n232 9.3005
R1673 drain_left.n231 drain_left.n230 9.3005
R1674 drain_left.n170 drain_left.n169 9.3005
R1675 drain_left.n225 drain_left.n224 9.3005
R1676 drain_left.n223 drain_left.n222 9.3005
R1677 drain_left.n174 drain_left.n173 9.3005
R1678 drain_left.n217 drain_left.n216 9.3005
R1679 drain_left.n215 drain_left.n214 9.3005
R1680 drain_left.n52 drain_left.n51 8.92171
R1681 drain_left.n85 drain_left.n26 8.92171
R1682 drain_left.n98 drain_left.n18 8.92171
R1683 drain_left.n132 drain_left.n131 8.92171
R1684 drain_left.n275 drain_left.n274 8.92171
R1685 drain_left.n242 drain_left.n162 8.92171
R1686 drain_left.n229 drain_left.n170 8.92171
R1687 drain_left.n197 drain_left.n196 8.92171
R1688 drain_left.n48 drain_left.n42 8.14595
R1689 drain_left.n86 drain_left.n24 8.14595
R1690 drain_left.n97 drain_left.n20 8.14595
R1691 drain_left.n135 drain_left.n2 8.14595
R1692 drain_left.n278 drain_left.n145 8.14595
R1693 drain_left.n241 drain_left.n164 8.14595
R1694 drain_left.n230 drain_left.n168 8.14595
R1695 drain_left.n193 drain_left.n187 8.14595
R1696 drain_left.n47 drain_left.n44 7.3702
R1697 drain_left.n90 drain_left.n89 7.3702
R1698 drain_left.n94 drain_left.n93 7.3702
R1699 drain_left.n136 drain_left.n0 7.3702
R1700 drain_left.n279 drain_left.n143 7.3702
R1701 drain_left.n238 drain_left.n237 7.3702
R1702 drain_left.n234 drain_left.n233 7.3702
R1703 drain_left.n192 drain_left.n189 7.3702
R1704 drain_left.n90 drain_left.n22 6.59444
R1705 drain_left.n93 drain_left.n22 6.59444
R1706 drain_left.n138 drain_left.n0 6.59444
R1707 drain_left.n281 drain_left.n143 6.59444
R1708 drain_left.n237 drain_left.n166 6.59444
R1709 drain_left.n234 drain_left.n166 6.59444
R1710 drain_left drain_left.n285 6.54115
R1711 drain_left.n48 drain_left.n47 5.81868
R1712 drain_left.n89 drain_left.n24 5.81868
R1713 drain_left.n94 drain_left.n20 5.81868
R1714 drain_left.n136 drain_left.n135 5.81868
R1715 drain_left.n279 drain_left.n278 5.81868
R1716 drain_left.n238 drain_left.n164 5.81868
R1717 drain_left.n233 drain_left.n168 5.81868
R1718 drain_left.n193 drain_left.n192 5.81868
R1719 drain_left.n51 drain_left.n42 5.04292
R1720 drain_left.n86 drain_left.n85 5.04292
R1721 drain_left.n98 drain_left.n97 5.04292
R1722 drain_left.n132 drain_left.n2 5.04292
R1723 drain_left.n275 drain_left.n145 5.04292
R1724 drain_left.n242 drain_left.n241 5.04292
R1725 drain_left.n230 drain_left.n229 5.04292
R1726 drain_left.n196 drain_left.n187 5.04292
R1727 drain_left.n52 drain_left.n40 4.26717
R1728 drain_left.n82 drain_left.n26 4.26717
R1729 drain_left.n101 drain_left.n18 4.26717
R1730 drain_left.n131 drain_left.n4 4.26717
R1731 drain_left.n274 drain_left.n147 4.26717
R1732 drain_left.n245 drain_left.n162 4.26717
R1733 drain_left.n226 drain_left.n170 4.26717
R1734 drain_left.n197 drain_left.n185 4.26717
R1735 drain_left.n56 drain_left.n55 3.49141
R1736 drain_left.n81 drain_left.n28 3.49141
R1737 drain_left.n102 drain_left.n16 3.49141
R1738 drain_left.n128 drain_left.n127 3.49141
R1739 drain_left.n271 drain_left.n270 3.49141
R1740 drain_left.n246 drain_left.n160 3.49141
R1741 drain_left.n225 drain_left.n172 3.49141
R1742 drain_left.n201 drain_left.n200 3.49141
R1743 drain_left.n191 drain_left.n190 2.84303
R1744 drain_left.n46 drain_left.n45 2.84303
R1745 drain_left.n59 drain_left.n38 2.71565
R1746 drain_left.n78 drain_left.n77 2.71565
R1747 drain_left.n106 drain_left.n105 2.71565
R1748 drain_left.n124 drain_left.n6 2.71565
R1749 drain_left.n267 drain_left.n149 2.71565
R1750 drain_left.n250 drain_left.n249 2.71565
R1751 drain_left.n222 drain_left.n221 2.71565
R1752 drain_left.n204 drain_left.n183 2.71565
R1753 drain_left.n60 drain_left.n36 1.93989
R1754 drain_left.n74 drain_left.n30 1.93989
R1755 drain_left.n110 drain_left.n14 1.93989
R1756 drain_left.n123 drain_left.n8 1.93989
R1757 drain_left.n266 drain_left.n151 1.93989
R1758 drain_left.n253 drain_left.n157 1.93989
R1759 drain_left.n218 drain_left.n174 1.93989
R1760 drain_left.n205 drain_left.n181 1.93989
R1761 drain_left.n65 drain_left.n63 1.16414
R1762 drain_left.n73 drain_left.n32 1.16414
R1763 drain_left.n111 drain_left.n12 1.16414
R1764 drain_left.n120 drain_left.n119 1.16414
R1765 drain_left.n263 drain_left.n262 1.16414
R1766 drain_left.n254 drain_left.n155 1.16414
R1767 drain_left.n217 drain_left.n176 1.16414
R1768 drain_left.n209 drain_left.n208 1.16414
R1769 drain_left.n285 drain_left.n283 0.888431
R1770 drain_left.n141 drain_left.t9 0.7925
R1771 drain_left.n141 drain_left.t0 0.7925
R1772 drain_left.n139 drain_left.t5 0.7925
R1773 drain_left.n139 drain_left.t1 0.7925
R1774 drain_left.n284 drain_left.t4 0.7925
R1775 drain_left.n284 drain_left.t7 0.7925
R1776 drain_left.n282 drain_left.t2 0.7925
R1777 drain_left.n282 drain_left.t8 0.7925
R1778 drain_left.n64 drain_left.n34 0.388379
R1779 drain_left.n70 drain_left.n69 0.388379
R1780 drain_left.n115 drain_left.n114 0.388379
R1781 drain_left.n116 drain_left.n10 0.388379
R1782 drain_left.n259 drain_left.n153 0.388379
R1783 drain_left.n258 drain_left.n257 0.388379
R1784 drain_left.n214 drain_left.n213 0.388379
R1785 drain_left.n180 drain_left.n178 0.388379
R1786 drain_left.n142 drain_left.n140 0.167137
R1787 drain_left.n46 drain_left.n41 0.155672
R1788 drain_left.n53 drain_left.n41 0.155672
R1789 drain_left.n54 drain_left.n53 0.155672
R1790 drain_left.n54 drain_left.n37 0.155672
R1791 drain_left.n61 drain_left.n37 0.155672
R1792 drain_left.n62 drain_left.n61 0.155672
R1793 drain_left.n62 drain_left.n33 0.155672
R1794 drain_left.n71 drain_left.n33 0.155672
R1795 drain_left.n72 drain_left.n71 0.155672
R1796 drain_left.n72 drain_left.n29 0.155672
R1797 drain_left.n79 drain_left.n29 0.155672
R1798 drain_left.n80 drain_left.n79 0.155672
R1799 drain_left.n80 drain_left.n25 0.155672
R1800 drain_left.n87 drain_left.n25 0.155672
R1801 drain_left.n88 drain_left.n87 0.155672
R1802 drain_left.n88 drain_left.n21 0.155672
R1803 drain_left.n95 drain_left.n21 0.155672
R1804 drain_left.n96 drain_left.n95 0.155672
R1805 drain_left.n96 drain_left.n17 0.155672
R1806 drain_left.n103 drain_left.n17 0.155672
R1807 drain_left.n104 drain_left.n103 0.155672
R1808 drain_left.n104 drain_left.n13 0.155672
R1809 drain_left.n112 drain_left.n13 0.155672
R1810 drain_left.n113 drain_left.n112 0.155672
R1811 drain_left.n113 drain_left.n9 0.155672
R1812 drain_left.n121 drain_left.n9 0.155672
R1813 drain_left.n122 drain_left.n121 0.155672
R1814 drain_left.n122 drain_left.n5 0.155672
R1815 drain_left.n129 drain_left.n5 0.155672
R1816 drain_left.n130 drain_left.n129 0.155672
R1817 drain_left.n130 drain_left.n1 0.155672
R1818 drain_left.n137 drain_left.n1 0.155672
R1819 drain_left.n280 drain_left.n144 0.155672
R1820 drain_left.n273 drain_left.n144 0.155672
R1821 drain_left.n273 drain_left.n272 0.155672
R1822 drain_left.n272 drain_left.n148 0.155672
R1823 drain_left.n265 drain_left.n148 0.155672
R1824 drain_left.n265 drain_left.n264 0.155672
R1825 drain_left.n264 drain_left.n152 0.155672
R1826 drain_left.n256 drain_left.n152 0.155672
R1827 drain_left.n256 drain_left.n255 0.155672
R1828 drain_left.n255 drain_left.n156 0.155672
R1829 drain_left.n248 drain_left.n156 0.155672
R1830 drain_left.n248 drain_left.n247 0.155672
R1831 drain_left.n247 drain_left.n161 0.155672
R1832 drain_left.n240 drain_left.n161 0.155672
R1833 drain_left.n240 drain_left.n239 0.155672
R1834 drain_left.n239 drain_left.n165 0.155672
R1835 drain_left.n232 drain_left.n165 0.155672
R1836 drain_left.n232 drain_left.n231 0.155672
R1837 drain_left.n231 drain_left.n169 0.155672
R1838 drain_left.n224 drain_left.n169 0.155672
R1839 drain_left.n224 drain_left.n223 0.155672
R1840 drain_left.n223 drain_left.n173 0.155672
R1841 drain_left.n216 drain_left.n173 0.155672
R1842 drain_left.n216 drain_left.n215 0.155672
R1843 drain_left.n215 drain_left.n177 0.155672
R1844 drain_left.n207 drain_left.n177 0.155672
R1845 drain_left.n207 drain_left.n206 0.155672
R1846 drain_left.n206 drain_left.n182 0.155672
R1847 drain_left.n199 drain_left.n182 0.155672
R1848 drain_left.n199 drain_left.n198 0.155672
R1849 drain_left.n198 drain_left.n186 0.155672
R1850 drain_left.n191 drain_left.n186 0.155672
C0 source drain_left 27.138699f
C1 drain_right drain_left 0.973273f
C2 plus minus 7.984509f
C3 drain_right source 27.123901f
C4 plus drain_left 13.6936f
C5 plus source 12.8445f
C6 drain_right plus 0.349144f
C7 minus drain_left 0.171897f
C8 minus source 12.829401f
C9 drain_right minus 13.508201f
C10 drain_right a_n1952_n5888# 10.48311f
C11 drain_left a_n1952_n5888# 10.77967f
C12 source a_n1952_n5888# 11.260633f
C13 minus a_n1952_n5888# 8.512239f
C14 plus a_n1952_n5888# 10.87721f
C15 drain_left.n0 a_n1952_n5888# 0.033526f
C16 drain_left.n1 a_n1952_n5888# 0.024319f
C17 drain_left.n2 a_n1952_n5888# 0.013068f
C18 drain_left.n3 a_n1952_n5888# 0.030888f
C19 drain_left.n4 a_n1952_n5888# 0.013837f
C20 drain_left.n5 a_n1952_n5888# 0.024319f
C21 drain_left.n6 a_n1952_n5888# 0.013068f
C22 drain_left.n7 a_n1952_n5888# 0.030888f
C23 drain_left.n8 a_n1952_n5888# 0.013837f
C24 drain_left.n9 a_n1952_n5888# 0.024319f
C25 drain_left.n10 a_n1952_n5888# 0.013068f
C26 drain_left.n11 a_n1952_n5888# 0.030888f
C27 drain_left.n12 a_n1952_n5888# 0.013837f
C28 drain_left.n13 a_n1952_n5888# 0.024319f
C29 drain_left.n14 a_n1952_n5888# 0.013068f
C30 drain_left.n15 a_n1952_n5888# 0.030888f
C31 drain_left.n16 a_n1952_n5888# 0.013837f
C32 drain_left.n17 a_n1952_n5888# 0.024319f
C33 drain_left.n18 a_n1952_n5888# 0.013068f
C34 drain_left.n19 a_n1952_n5888# 0.030888f
C35 drain_left.n20 a_n1952_n5888# 0.013837f
C36 drain_left.n21 a_n1952_n5888# 0.024319f
C37 drain_left.n22 a_n1952_n5888# 0.013068f
C38 drain_left.n23 a_n1952_n5888# 0.030888f
C39 drain_left.n24 a_n1952_n5888# 0.013837f
C40 drain_left.n25 a_n1952_n5888# 0.024319f
C41 drain_left.n26 a_n1952_n5888# 0.013068f
C42 drain_left.n27 a_n1952_n5888# 0.030888f
C43 drain_left.n28 a_n1952_n5888# 0.013837f
C44 drain_left.n29 a_n1952_n5888# 0.024319f
C45 drain_left.n30 a_n1952_n5888# 0.013068f
C46 drain_left.n31 a_n1952_n5888# 0.030888f
C47 drain_left.n32 a_n1952_n5888# 0.013837f
C48 drain_left.n33 a_n1952_n5888# 0.024319f
C49 drain_left.n34 a_n1952_n5888# 0.013452f
C50 drain_left.n35 a_n1952_n5888# 0.030888f
C51 drain_left.n36 a_n1952_n5888# 0.013837f
C52 drain_left.n37 a_n1952_n5888# 0.024319f
C53 drain_left.n38 a_n1952_n5888# 0.013068f
C54 drain_left.n39 a_n1952_n5888# 0.030888f
C55 drain_left.n40 a_n1952_n5888# 0.013837f
C56 drain_left.n41 a_n1952_n5888# 0.024319f
C57 drain_left.n42 a_n1952_n5888# 0.013068f
C58 drain_left.n43 a_n1952_n5888# 0.023166f
C59 drain_left.n44 a_n1952_n5888# 0.021835f
C60 drain_left.t3 a_n1952_n5888# 0.05387f
C61 drain_left.n45 a_n1952_n5888# 0.296712f
C62 drain_left.n46 a_n1952_n5888# 2.63303f
C63 drain_left.n47 a_n1952_n5888# 0.013068f
C64 drain_left.n48 a_n1952_n5888# 0.013837f
C65 drain_left.n49 a_n1952_n5888# 0.030888f
C66 drain_left.n50 a_n1952_n5888# 0.030888f
C67 drain_left.n51 a_n1952_n5888# 0.013837f
C68 drain_left.n52 a_n1952_n5888# 0.013068f
C69 drain_left.n53 a_n1952_n5888# 0.024319f
C70 drain_left.n54 a_n1952_n5888# 0.024319f
C71 drain_left.n55 a_n1952_n5888# 0.013068f
C72 drain_left.n56 a_n1952_n5888# 0.013837f
C73 drain_left.n57 a_n1952_n5888# 0.030888f
C74 drain_left.n58 a_n1952_n5888# 0.030888f
C75 drain_left.n59 a_n1952_n5888# 0.013837f
C76 drain_left.n60 a_n1952_n5888# 0.013068f
C77 drain_left.n61 a_n1952_n5888# 0.024319f
C78 drain_left.n62 a_n1952_n5888# 0.024319f
C79 drain_left.n63 a_n1952_n5888# 0.013068f
C80 drain_left.n64 a_n1952_n5888# 0.013068f
C81 drain_left.n65 a_n1952_n5888# 0.013837f
C82 drain_left.n66 a_n1952_n5888# 0.030888f
C83 drain_left.n67 a_n1952_n5888# 0.030888f
C84 drain_left.n68 a_n1952_n5888# 0.030888f
C85 drain_left.n69 a_n1952_n5888# 0.013452f
C86 drain_left.n70 a_n1952_n5888# 0.013068f
C87 drain_left.n71 a_n1952_n5888# 0.024319f
C88 drain_left.n72 a_n1952_n5888# 0.024319f
C89 drain_left.n73 a_n1952_n5888# 0.013068f
C90 drain_left.n74 a_n1952_n5888# 0.013837f
C91 drain_left.n75 a_n1952_n5888# 0.030888f
C92 drain_left.n76 a_n1952_n5888# 0.030888f
C93 drain_left.n77 a_n1952_n5888# 0.013837f
C94 drain_left.n78 a_n1952_n5888# 0.013068f
C95 drain_left.n79 a_n1952_n5888# 0.024319f
C96 drain_left.n80 a_n1952_n5888# 0.024319f
C97 drain_left.n81 a_n1952_n5888# 0.013068f
C98 drain_left.n82 a_n1952_n5888# 0.013837f
C99 drain_left.n83 a_n1952_n5888# 0.030888f
C100 drain_left.n84 a_n1952_n5888# 0.030888f
C101 drain_left.n85 a_n1952_n5888# 0.013837f
C102 drain_left.n86 a_n1952_n5888# 0.013068f
C103 drain_left.n87 a_n1952_n5888# 0.024319f
C104 drain_left.n88 a_n1952_n5888# 0.024319f
C105 drain_left.n89 a_n1952_n5888# 0.013068f
C106 drain_left.n90 a_n1952_n5888# 0.013837f
C107 drain_left.n91 a_n1952_n5888# 0.030888f
C108 drain_left.n92 a_n1952_n5888# 0.030888f
C109 drain_left.n93 a_n1952_n5888# 0.013837f
C110 drain_left.n94 a_n1952_n5888# 0.013068f
C111 drain_left.n95 a_n1952_n5888# 0.024319f
C112 drain_left.n96 a_n1952_n5888# 0.024319f
C113 drain_left.n97 a_n1952_n5888# 0.013068f
C114 drain_left.n98 a_n1952_n5888# 0.013837f
C115 drain_left.n99 a_n1952_n5888# 0.030888f
C116 drain_left.n100 a_n1952_n5888# 0.030888f
C117 drain_left.n101 a_n1952_n5888# 0.013837f
C118 drain_left.n102 a_n1952_n5888# 0.013068f
C119 drain_left.n103 a_n1952_n5888# 0.024319f
C120 drain_left.n104 a_n1952_n5888# 0.024319f
C121 drain_left.n105 a_n1952_n5888# 0.013068f
C122 drain_left.n106 a_n1952_n5888# 0.013837f
C123 drain_left.n107 a_n1952_n5888# 0.030888f
C124 drain_left.n108 a_n1952_n5888# 0.030888f
C125 drain_left.n109 a_n1952_n5888# 0.030888f
C126 drain_left.n110 a_n1952_n5888# 0.013837f
C127 drain_left.n111 a_n1952_n5888# 0.013068f
C128 drain_left.n112 a_n1952_n5888# 0.024319f
C129 drain_left.n113 a_n1952_n5888# 0.024319f
C130 drain_left.n114 a_n1952_n5888# 0.013068f
C131 drain_left.n115 a_n1952_n5888# 0.013452f
C132 drain_left.n116 a_n1952_n5888# 0.013452f
C133 drain_left.n117 a_n1952_n5888# 0.030888f
C134 drain_left.n118 a_n1952_n5888# 0.030888f
C135 drain_left.n119 a_n1952_n5888# 0.013837f
C136 drain_left.n120 a_n1952_n5888# 0.013068f
C137 drain_left.n121 a_n1952_n5888# 0.024319f
C138 drain_left.n122 a_n1952_n5888# 0.024319f
C139 drain_left.n123 a_n1952_n5888# 0.013068f
C140 drain_left.n124 a_n1952_n5888# 0.013837f
C141 drain_left.n125 a_n1952_n5888# 0.030888f
C142 drain_left.n126 a_n1952_n5888# 0.030888f
C143 drain_left.n127 a_n1952_n5888# 0.013837f
C144 drain_left.n128 a_n1952_n5888# 0.013068f
C145 drain_left.n129 a_n1952_n5888# 0.024319f
C146 drain_left.n130 a_n1952_n5888# 0.024319f
C147 drain_left.n131 a_n1952_n5888# 0.013068f
C148 drain_left.n132 a_n1952_n5888# 0.013837f
C149 drain_left.n133 a_n1952_n5888# 0.030888f
C150 drain_left.n134 a_n1952_n5888# 0.065706f
C151 drain_left.n135 a_n1952_n5888# 0.013837f
C152 drain_left.n136 a_n1952_n5888# 0.013068f
C153 drain_left.n137 a_n1952_n5888# 0.053554f
C154 drain_left.n138 a_n1952_n5888# 0.055493f
C155 drain_left.t5 a_n1952_n5888# 0.48044f
C156 drain_left.t1 a_n1952_n5888# 0.48044f
C157 drain_left.n139 a_n1952_n5888# 4.42777f
C158 drain_left.n140 a_n1952_n5888# 0.404357f
C159 drain_left.t9 a_n1952_n5888# 0.48044f
C160 drain_left.t0 a_n1952_n5888# 0.48044f
C161 drain_left.n141 a_n1952_n5888# 4.43121f
C162 drain_left.n142 a_n1952_n5888# 2.36641f
C163 drain_left.n143 a_n1952_n5888# 0.033526f
C164 drain_left.n144 a_n1952_n5888# 0.024319f
C165 drain_left.n145 a_n1952_n5888# 0.013068f
C166 drain_left.n146 a_n1952_n5888# 0.030888f
C167 drain_left.n147 a_n1952_n5888# 0.013837f
C168 drain_left.n148 a_n1952_n5888# 0.024319f
C169 drain_left.n149 a_n1952_n5888# 0.013068f
C170 drain_left.n150 a_n1952_n5888# 0.030888f
C171 drain_left.n151 a_n1952_n5888# 0.013837f
C172 drain_left.n152 a_n1952_n5888# 0.024319f
C173 drain_left.n153 a_n1952_n5888# 0.013068f
C174 drain_left.n154 a_n1952_n5888# 0.030888f
C175 drain_left.n155 a_n1952_n5888# 0.013837f
C176 drain_left.n156 a_n1952_n5888# 0.024319f
C177 drain_left.n157 a_n1952_n5888# 0.013068f
C178 drain_left.n158 a_n1952_n5888# 0.030888f
C179 drain_left.n159 a_n1952_n5888# 0.030888f
C180 drain_left.n160 a_n1952_n5888# 0.013837f
C181 drain_left.n161 a_n1952_n5888# 0.024319f
C182 drain_left.n162 a_n1952_n5888# 0.013068f
C183 drain_left.n163 a_n1952_n5888# 0.030888f
C184 drain_left.n164 a_n1952_n5888# 0.013837f
C185 drain_left.n165 a_n1952_n5888# 0.024319f
C186 drain_left.n166 a_n1952_n5888# 0.013068f
C187 drain_left.n167 a_n1952_n5888# 0.030888f
C188 drain_left.n168 a_n1952_n5888# 0.013837f
C189 drain_left.n169 a_n1952_n5888# 0.024319f
C190 drain_left.n170 a_n1952_n5888# 0.013068f
C191 drain_left.n171 a_n1952_n5888# 0.030888f
C192 drain_left.n172 a_n1952_n5888# 0.013837f
C193 drain_left.n173 a_n1952_n5888# 0.024319f
C194 drain_left.n174 a_n1952_n5888# 0.013068f
C195 drain_left.n175 a_n1952_n5888# 0.030888f
C196 drain_left.n176 a_n1952_n5888# 0.013837f
C197 drain_left.n177 a_n1952_n5888# 0.024319f
C198 drain_left.n178 a_n1952_n5888# 0.013452f
C199 drain_left.n179 a_n1952_n5888# 0.030888f
C200 drain_left.n180 a_n1952_n5888# 0.013068f
C201 drain_left.n181 a_n1952_n5888# 0.013837f
C202 drain_left.n182 a_n1952_n5888# 0.024319f
C203 drain_left.n183 a_n1952_n5888# 0.013068f
C204 drain_left.n184 a_n1952_n5888# 0.030888f
C205 drain_left.n185 a_n1952_n5888# 0.013837f
C206 drain_left.n186 a_n1952_n5888# 0.024319f
C207 drain_left.n187 a_n1952_n5888# 0.013068f
C208 drain_left.n188 a_n1952_n5888# 0.023166f
C209 drain_left.n189 a_n1952_n5888# 0.021835f
C210 drain_left.t6 a_n1952_n5888# 0.05387f
C211 drain_left.n190 a_n1952_n5888# 0.296712f
C212 drain_left.n191 a_n1952_n5888# 2.63303f
C213 drain_left.n192 a_n1952_n5888# 0.013068f
C214 drain_left.n193 a_n1952_n5888# 0.013837f
C215 drain_left.n194 a_n1952_n5888# 0.030888f
C216 drain_left.n195 a_n1952_n5888# 0.030888f
C217 drain_left.n196 a_n1952_n5888# 0.013837f
C218 drain_left.n197 a_n1952_n5888# 0.013068f
C219 drain_left.n198 a_n1952_n5888# 0.024319f
C220 drain_left.n199 a_n1952_n5888# 0.024319f
C221 drain_left.n200 a_n1952_n5888# 0.013068f
C222 drain_left.n201 a_n1952_n5888# 0.013837f
C223 drain_left.n202 a_n1952_n5888# 0.030888f
C224 drain_left.n203 a_n1952_n5888# 0.030888f
C225 drain_left.n204 a_n1952_n5888# 0.013837f
C226 drain_left.n205 a_n1952_n5888# 0.013068f
C227 drain_left.n206 a_n1952_n5888# 0.024319f
C228 drain_left.n207 a_n1952_n5888# 0.024319f
C229 drain_left.n208 a_n1952_n5888# 0.013068f
C230 drain_left.n209 a_n1952_n5888# 0.013837f
C231 drain_left.n210 a_n1952_n5888# 0.030888f
C232 drain_left.n211 a_n1952_n5888# 0.030888f
C233 drain_left.n212 a_n1952_n5888# 0.030888f
C234 drain_left.n213 a_n1952_n5888# 0.013452f
C235 drain_left.n214 a_n1952_n5888# 0.013068f
C236 drain_left.n215 a_n1952_n5888# 0.024319f
C237 drain_left.n216 a_n1952_n5888# 0.024319f
C238 drain_left.n217 a_n1952_n5888# 0.013068f
C239 drain_left.n218 a_n1952_n5888# 0.013837f
C240 drain_left.n219 a_n1952_n5888# 0.030888f
C241 drain_left.n220 a_n1952_n5888# 0.030888f
C242 drain_left.n221 a_n1952_n5888# 0.013837f
C243 drain_left.n222 a_n1952_n5888# 0.013068f
C244 drain_left.n223 a_n1952_n5888# 0.024319f
C245 drain_left.n224 a_n1952_n5888# 0.024319f
C246 drain_left.n225 a_n1952_n5888# 0.013068f
C247 drain_left.n226 a_n1952_n5888# 0.013837f
C248 drain_left.n227 a_n1952_n5888# 0.030888f
C249 drain_left.n228 a_n1952_n5888# 0.030888f
C250 drain_left.n229 a_n1952_n5888# 0.013837f
C251 drain_left.n230 a_n1952_n5888# 0.013068f
C252 drain_left.n231 a_n1952_n5888# 0.024319f
C253 drain_left.n232 a_n1952_n5888# 0.024319f
C254 drain_left.n233 a_n1952_n5888# 0.013068f
C255 drain_left.n234 a_n1952_n5888# 0.013837f
C256 drain_left.n235 a_n1952_n5888# 0.030888f
C257 drain_left.n236 a_n1952_n5888# 0.030888f
C258 drain_left.n237 a_n1952_n5888# 0.013837f
C259 drain_left.n238 a_n1952_n5888# 0.013068f
C260 drain_left.n239 a_n1952_n5888# 0.024319f
C261 drain_left.n240 a_n1952_n5888# 0.024319f
C262 drain_left.n241 a_n1952_n5888# 0.013068f
C263 drain_left.n242 a_n1952_n5888# 0.013837f
C264 drain_left.n243 a_n1952_n5888# 0.030888f
C265 drain_left.n244 a_n1952_n5888# 0.030888f
C266 drain_left.n245 a_n1952_n5888# 0.013837f
C267 drain_left.n246 a_n1952_n5888# 0.013068f
C268 drain_left.n247 a_n1952_n5888# 0.024319f
C269 drain_left.n248 a_n1952_n5888# 0.024319f
C270 drain_left.n249 a_n1952_n5888# 0.013068f
C271 drain_left.n250 a_n1952_n5888# 0.013837f
C272 drain_left.n251 a_n1952_n5888# 0.030888f
C273 drain_left.n252 a_n1952_n5888# 0.030888f
C274 drain_left.n253 a_n1952_n5888# 0.013837f
C275 drain_left.n254 a_n1952_n5888# 0.013068f
C276 drain_left.n255 a_n1952_n5888# 0.024319f
C277 drain_left.n256 a_n1952_n5888# 0.024319f
C278 drain_left.n257 a_n1952_n5888# 0.013068f
C279 drain_left.n258 a_n1952_n5888# 0.013452f
C280 drain_left.n259 a_n1952_n5888# 0.013452f
C281 drain_left.n260 a_n1952_n5888# 0.030888f
C282 drain_left.n261 a_n1952_n5888# 0.030888f
C283 drain_left.n262 a_n1952_n5888# 0.013837f
C284 drain_left.n263 a_n1952_n5888# 0.013068f
C285 drain_left.n264 a_n1952_n5888# 0.024319f
C286 drain_left.n265 a_n1952_n5888# 0.024319f
C287 drain_left.n266 a_n1952_n5888# 0.013068f
C288 drain_left.n267 a_n1952_n5888# 0.013837f
C289 drain_left.n268 a_n1952_n5888# 0.030888f
C290 drain_left.n269 a_n1952_n5888# 0.030888f
C291 drain_left.n270 a_n1952_n5888# 0.013837f
C292 drain_left.n271 a_n1952_n5888# 0.013068f
C293 drain_left.n272 a_n1952_n5888# 0.024319f
C294 drain_left.n273 a_n1952_n5888# 0.024319f
C295 drain_left.n274 a_n1952_n5888# 0.013068f
C296 drain_left.n275 a_n1952_n5888# 0.013837f
C297 drain_left.n276 a_n1952_n5888# 0.030888f
C298 drain_left.n277 a_n1952_n5888# 0.065706f
C299 drain_left.n278 a_n1952_n5888# 0.013837f
C300 drain_left.n279 a_n1952_n5888# 0.013068f
C301 drain_left.n280 a_n1952_n5888# 0.053554f
C302 drain_left.n281 a_n1952_n5888# 0.055493f
C303 drain_left.t2 a_n1952_n5888# 0.48044f
C304 drain_left.t8 a_n1952_n5888# 0.48044f
C305 drain_left.n282 a_n1952_n5888# 4.42777f
C306 drain_left.n283 a_n1952_n5888# 0.457494f
C307 drain_left.t4 a_n1952_n5888# 0.48044f
C308 drain_left.t7 a_n1952_n5888# 0.48044f
C309 drain_left.n284 a_n1952_n5888# 4.42776f
C310 drain_left.n285 a_n1952_n5888# 0.559837f
C311 plus.n0 a_n1952_n5888# 0.042565f
C312 plus.t2 a_n1952_n5888# 2.10505f
C313 plus.t5 a_n1952_n5888# 2.10505f
C314 plus.n1 a_n1952_n5888# 0.042565f
C315 plus.t1 a_n1952_n5888# 2.10505f
C316 plus.n2 a_n1952_n5888# 0.768449f
C317 plus.t3 a_n1952_n5888# 2.12365f
C318 plus.n3 a_n1952_n5888# 0.753729f
C319 plus.t7 a_n1952_n5888# 2.10505f
C320 plus.n4 a_n1952_n5888# 0.772738f
C321 plus.n5 a_n1952_n5888# 0.009659f
C322 plus.n6 a_n1952_n5888# 0.177785f
C323 plus.n7 a_n1952_n5888# 0.042565f
C324 plus.n8 a_n1952_n5888# 0.042565f
C325 plus.n9 a_n1952_n5888# 0.009659f
C326 plus.n10 a_n1952_n5888# 0.768449f
C327 plus.n11 a_n1952_n5888# 0.009659f
C328 plus.n12 a_n1952_n5888# 0.766087f
C329 plus.n13 a_n1952_n5888# 0.773067f
C330 plus.n14 a_n1952_n5888# 0.042565f
C331 plus.t6 a_n1952_n5888# 2.10505f
C332 plus.n15 a_n1952_n5888# 0.042565f
C333 plus.t4 a_n1952_n5888# 2.10505f
C334 plus.t8 a_n1952_n5888# 2.10505f
C335 plus.n16 a_n1952_n5888# 0.768449f
C336 plus.t9 a_n1952_n5888# 2.12365f
C337 plus.n17 a_n1952_n5888# 0.753729f
C338 plus.t0 a_n1952_n5888# 2.10505f
C339 plus.n18 a_n1952_n5888# 0.772738f
C340 plus.n19 a_n1952_n5888# 0.009659f
C341 plus.n20 a_n1952_n5888# 0.177785f
C342 plus.n21 a_n1952_n5888# 0.042565f
C343 plus.n22 a_n1952_n5888# 0.042565f
C344 plus.n23 a_n1952_n5888# 0.009659f
C345 plus.n24 a_n1952_n5888# 0.768449f
C346 plus.n25 a_n1952_n5888# 0.009659f
C347 plus.n26 a_n1952_n5888# 0.766087f
C348 plus.n27 a_n1952_n5888# 1.67965f
C349 drain_right.n0 a_n1952_n5888# 0.03344f
C350 drain_right.n1 a_n1952_n5888# 0.024256f
C351 drain_right.n2 a_n1952_n5888# 0.013034f
C352 drain_right.n3 a_n1952_n5888# 0.030808f
C353 drain_right.n4 a_n1952_n5888# 0.013801f
C354 drain_right.n5 a_n1952_n5888# 0.024256f
C355 drain_right.n6 a_n1952_n5888# 0.013034f
C356 drain_right.n7 a_n1952_n5888# 0.030808f
C357 drain_right.n8 a_n1952_n5888# 0.013801f
C358 drain_right.n9 a_n1952_n5888# 0.024256f
C359 drain_right.n10 a_n1952_n5888# 0.013034f
C360 drain_right.n11 a_n1952_n5888# 0.030808f
C361 drain_right.n12 a_n1952_n5888# 0.013801f
C362 drain_right.n13 a_n1952_n5888# 0.024256f
C363 drain_right.n14 a_n1952_n5888# 0.013034f
C364 drain_right.n15 a_n1952_n5888# 0.030808f
C365 drain_right.n16 a_n1952_n5888# 0.013801f
C366 drain_right.n17 a_n1952_n5888# 0.024256f
C367 drain_right.n18 a_n1952_n5888# 0.013034f
C368 drain_right.n19 a_n1952_n5888# 0.030808f
C369 drain_right.n20 a_n1952_n5888# 0.013801f
C370 drain_right.n21 a_n1952_n5888# 0.024256f
C371 drain_right.n22 a_n1952_n5888# 0.013034f
C372 drain_right.n23 a_n1952_n5888# 0.030808f
C373 drain_right.n24 a_n1952_n5888# 0.013801f
C374 drain_right.n25 a_n1952_n5888# 0.024256f
C375 drain_right.n26 a_n1952_n5888# 0.013034f
C376 drain_right.n27 a_n1952_n5888# 0.030808f
C377 drain_right.n28 a_n1952_n5888# 0.013801f
C378 drain_right.n29 a_n1952_n5888# 0.024256f
C379 drain_right.n30 a_n1952_n5888# 0.013034f
C380 drain_right.n31 a_n1952_n5888# 0.030808f
C381 drain_right.n32 a_n1952_n5888# 0.013801f
C382 drain_right.n33 a_n1952_n5888# 0.024256f
C383 drain_right.n34 a_n1952_n5888# 0.013418f
C384 drain_right.n35 a_n1952_n5888# 0.030808f
C385 drain_right.n36 a_n1952_n5888# 0.013801f
C386 drain_right.n37 a_n1952_n5888# 0.024256f
C387 drain_right.n38 a_n1952_n5888# 0.013034f
C388 drain_right.n39 a_n1952_n5888# 0.030808f
C389 drain_right.n40 a_n1952_n5888# 0.013801f
C390 drain_right.n41 a_n1952_n5888# 0.024256f
C391 drain_right.n42 a_n1952_n5888# 0.013034f
C392 drain_right.n43 a_n1952_n5888# 0.023106f
C393 drain_right.n44 a_n1952_n5888# 0.021779f
C394 drain_right.t4 a_n1952_n5888# 0.053732f
C395 drain_right.n45 a_n1952_n5888# 0.295948f
C396 drain_right.n46 a_n1952_n5888# 2.62625f
C397 drain_right.n47 a_n1952_n5888# 0.013034f
C398 drain_right.n48 a_n1952_n5888# 0.013801f
C399 drain_right.n49 a_n1952_n5888# 0.030808f
C400 drain_right.n50 a_n1952_n5888# 0.030808f
C401 drain_right.n51 a_n1952_n5888# 0.013801f
C402 drain_right.n52 a_n1952_n5888# 0.013034f
C403 drain_right.n53 a_n1952_n5888# 0.024256f
C404 drain_right.n54 a_n1952_n5888# 0.024256f
C405 drain_right.n55 a_n1952_n5888# 0.013034f
C406 drain_right.n56 a_n1952_n5888# 0.013801f
C407 drain_right.n57 a_n1952_n5888# 0.030808f
C408 drain_right.n58 a_n1952_n5888# 0.030808f
C409 drain_right.n59 a_n1952_n5888# 0.013801f
C410 drain_right.n60 a_n1952_n5888# 0.013034f
C411 drain_right.n61 a_n1952_n5888# 0.024256f
C412 drain_right.n62 a_n1952_n5888# 0.024256f
C413 drain_right.n63 a_n1952_n5888# 0.013034f
C414 drain_right.n64 a_n1952_n5888# 0.013034f
C415 drain_right.n65 a_n1952_n5888# 0.013801f
C416 drain_right.n66 a_n1952_n5888# 0.030808f
C417 drain_right.n67 a_n1952_n5888# 0.030808f
C418 drain_right.n68 a_n1952_n5888# 0.030808f
C419 drain_right.n69 a_n1952_n5888# 0.013418f
C420 drain_right.n70 a_n1952_n5888# 0.013034f
C421 drain_right.n71 a_n1952_n5888# 0.024256f
C422 drain_right.n72 a_n1952_n5888# 0.024256f
C423 drain_right.n73 a_n1952_n5888# 0.013034f
C424 drain_right.n74 a_n1952_n5888# 0.013801f
C425 drain_right.n75 a_n1952_n5888# 0.030808f
C426 drain_right.n76 a_n1952_n5888# 0.030808f
C427 drain_right.n77 a_n1952_n5888# 0.013801f
C428 drain_right.n78 a_n1952_n5888# 0.013034f
C429 drain_right.n79 a_n1952_n5888# 0.024256f
C430 drain_right.n80 a_n1952_n5888# 0.024256f
C431 drain_right.n81 a_n1952_n5888# 0.013034f
C432 drain_right.n82 a_n1952_n5888# 0.013801f
C433 drain_right.n83 a_n1952_n5888# 0.030808f
C434 drain_right.n84 a_n1952_n5888# 0.030808f
C435 drain_right.n85 a_n1952_n5888# 0.013801f
C436 drain_right.n86 a_n1952_n5888# 0.013034f
C437 drain_right.n87 a_n1952_n5888# 0.024256f
C438 drain_right.n88 a_n1952_n5888# 0.024256f
C439 drain_right.n89 a_n1952_n5888# 0.013034f
C440 drain_right.n90 a_n1952_n5888# 0.013801f
C441 drain_right.n91 a_n1952_n5888# 0.030808f
C442 drain_right.n92 a_n1952_n5888# 0.030808f
C443 drain_right.n93 a_n1952_n5888# 0.013801f
C444 drain_right.n94 a_n1952_n5888# 0.013034f
C445 drain_right.n95 a_n1952_n5888# 0.024256f
C446 drain_right.n96 a_n1952_n5888# 0.024256f
C447 drain_right.n97 a_n1952_n5888# 0.013034f
C448 drain_right.n98 a_n1952_n5888# 0.013801f
C449 drain_right.n99 a_n1952_n5888# 0.030808f
C450 drain_right.n100 a_n1952_n5888# 0.030808f
C451 drain_right.n101 a_n1952_n5888# 0.013801f
C452 drain_right.n102 a_n1952_n5888# 0.013034f
C453 drain_right.n103 a_n1952_n5888# 0.024256f
C454 drain_right.n104 a_n1952_n5888# 0.024256f
C455 drain_right.n105 a_n1952_n5888# 0.013034f
C456 drain_right.n106 a_n1952_n5888# 0.013801f
C457 drain_right.n107 a_n1952_n5888# 0.030808f
C458 drain_right.n108 a_n1952_n5888# 0.030808f
C459 drain_right.n109 a_n1952_n5888# 0.030808f
C460 drain_right.n110 a_n1952_n5888# 0.013801f
C461 drain_right.n111 a_n1952_n5888# 0.013034f
C462 drain_right.n112 a_n1952_n5888# 0.024256f
C463 drain_right.n113 a_n1952_n5888# 0.024256f
C464 drain_right.n114 a_n1952_n5888# 0.013034f
C465 drain_right.n115 a_n1952_n5888# 0.013418f
C466 drain_right.n116 a_n1952_n5888# 0.013418f
C467 drain_right.n117 a_n1952_n5888# 0.030808f
C468 drain_right.n118 a_n1952_n5888# 0.030808f
C469 drain_right.n119 a_n1952_n5888# 0.013801f
C470 drain_right.n120 a_n1952_n5888# 0.013034f
C471 drain_right.n121 a_n1952_n5888# 0.024256f
C472 drain_right.n122 a_n1952_n5888# 0.024256f
C473 drain_right.n123 a_n1952_n5888# 0.013034f
C474 drain_right.n124 a_n1952_n5888# 0.013801f
C475 drain_right.n125 a_n1952_n5888# 0.030808f
C476 drain_right.n126 a_n1952_n5888# 0.030808f
C477 drain_right.n127 a_n1952_n5888# 0.013801f
C478 drain_right.n128 a_n1952_n5888# 0.013034f
C479 drain_right.n129 a_n1952_n5888# 0.024256f
C480 drain_right.n130 a_n1952_n5888# 0.024256f
C481 drain_right.n131 a_n1952_n5888# 0.013034f
C482 drain_right.n132 a_n1952_n5888# 0.013801f
C483 drain_right.n133 a_n1952_n5888# 0.030808f
C484 drain_right.n134 a_n1952_n5888# 0.065537f
C485 drain_right.n135 a_n1952_n5888# 0.013801f
C486 drain_right.n136 a_n1952_n5888# 0.013034f
C487 drain_right.n137 a_n1952_n5888# 0.053417f
C488 drain_right.n138 a_n1952_n5888# 0.05535f
C489 drain_right.t5 a_n1952_n5888# 0.479202f
C490 drain_right.t9 a_n1952_n5888# 0.479202f
C491 drain_right.n139 a_n1952_n5888# 4.41637f
C492 drain_right.n140 a_n1952_n5888# 0.403315f
C493 drain_right.t8 a_n1952_n5888# 0.479202f
C494 drain_right.t6 a_n1952_n5888# 0.479202f
C495 drain_right.n141 a_n1952_n5888# 4.41979f
C496 drain_right.n142 a_n1952_n5888# 2.31008f
C497 drain_right.t7 a_n1952_n5888# 0.479202f
C498 drain_right.t1 a_n1952_n5888# 0.479202f
C499 drain_right.n143 a_n1952_n5888# 4.42162f
C500 drain_right.t0 a_n1952_n5888# 0.479202f
C501 drain_right.t2 a_n1952_n5888# 0.479202f
C502 drain_right.n144 a_n1952_n5888# 4.41637f
C503 drain_right.n145 a_n1952_n5888# 0.692184f
C504 drain_right.n146 a_n1952_n5888# 0.03344f
C505 drain_right.n147 a_n1952_n5888# 0.024256f
C506 drain_right.n148 a_n1952_n5888# 0.013034f
C507 drain_right.n149 a_n1952_n5888# 0.030808f
C508 drain_right.n150 a_n1952_n5888# 0.013801f
C509 drain_right.n151 a_n1952_n5888# 0.024256f
C510 drain_right.n152 a_n1952_n5888# 0.013034f
C511 drain_right.n153 a_n1952_n5888# 0.030808f
C512 drain_right.n154 a_n1952_n5888# 0.013801f
C513 drain_right.n155 a_n1952_n5888# 0.024256f
C514 drain_right.n156 a_n1952_n5888# 0.013034f
C515 drain_right.n157 a_n1952_n5888# 0.030808f
C516 drain_right.n158 a_n1952_n5888# 0.013801f
C517 drain_right.n159 a_n1952_n5888# 0.024256f
C518 drain_right.n160 a_n1952_n5888# 0.013034f
C519 drain_right.n161 a_n1952_n5888# 0.030808f
C520 drain_right.n162 a_n1952_n5888# 0.030808f
C521 drain_right.n163 a_n1952_n5888# 0.013801f
C522 drain_right.n164 a_n1952_n5888# 0.024256f
C523 drain_right.n165 a_n1952_n5888# 0.013034f
C524 drain_right.n166 a_n1952_n5888# 0.030808f
C525 drain_right.n167 a_n1952_n5888# 0.013801f
C526 drain_right.n168 a_n1952_n5888# 0.024256f
C527 drain_right.n169 a_n1952_n5888# 0.013034f
C528 drain_right.n170 a_n1952_n5888# 0.030808f
C529 drain_right.n171 a_n1952_n5888# 0.013801f
C530 drain_right.n172 a_n1952_n5888# 0.024256f
C531 drain_right.n173 a_n1952_n5888# 0.013034f
C532 drain_right.n174 a_n1952_n5888# 0.030808f
C533 drain_right.n175 a_n1952_n5888# 0.013801f
C534 drain_right.n176 a_n1952_n5888# 0.024256f
C535 drain_right.n177 a_n1952_n5888# 0.013034f
C536 drain_right.n178 a_n1952_n5888# 0.030808f
C537 drain_right.n179 a_n1952_n5888# 0.013801f
C538 drain_right.n180 a_n1952_n5888# 0.024256f
C539 drain_right.n181 a_n1952_n5888# 0.013418f
C540 drain_right.n182 a_n1952_n5888# 0.030808f
C541 drain_right.n183 a_n1952_n5888# 0.013034f
C542 drain_right.n184 a_n1952_n5888# 0.013801f
C543 drain_right.n185 a_n1952_n5888# 0.024256f
C544 drain_right.n186 a_n1952_n5888# 0.013034f
C545 drain_right.n187 a_n1952_n5888# 0.030808f
C546 drain_right.n188 a_n1952_n5888# 0.013801f
C547 drain_right.n189 a_n1952_n5888# 0.024256f
C548 drain_right.n190 a_n1952_n5888# 0.013034f
C549 drain_right.n191 a_n1952_n5888# 0.023106f
C550 drain_right.n192 a_n1952_n5888# 0.021779f
C551 drain_right.t3 a_n1952_n5888# 0.053732f
C552 drain_right.n193 a_n1952_n5888# 0.295948f
C553 drain_right.n194 a_n1952_n5888# 2.62625f
C554 drain_right.n195 a_n1952_n5888# 0.013034f
C555 drain_right.n196 a_n1952_n5888# 0.013801f
C556 drain_right.n197 a_n1952_n5888# 0.030808f
C557 drain_right.n198 a_n1952_n5888# 0.030808f
C558 drain_right.n199 a_n1952_n5888# 0.013801f
C559 drain_right.n200 a_n1952_n5888# 0.013034f
C560 drain_right.n201 a_n1952_n5888# 0.024256f
C561 drain_right.n202 a_n1952_n5888# 0.024256f
C562 drain_right.n203 a_n1952_n5888# 0.013034f
C563 drain_right.n204 a_n1952_n5888# 0.013801f
C564 drain_right.n205 a_n1952_n5888# 0.030808f
C565 drain_right.n206 a_n1952_n5888# 0.030808f
C566 drain_right.n207 a_n1952_n5888# 0.013801f
C567 drain_right.n208 a_n1952_n5888# 0.013034f
C568 drain_right.n209 a_n1952_n5888# 0.024256f
C569 drain_right.n210 a_n1952_n5888# 0.024256f
C570 drain_right.n211 a_n1952_n5888# 0.013034f
C571 drain_right.n212 a_n1952_n5888# 0.013801f
C572 drain_right.n213 a_n1952_n5888# 0.030808f
C573 drain_right.n214 a_n1952_n5888# 0.030808f
C574 drain_right.n215 a_n1952_n5888# 0.030808f
C575 drain_right.n216 a_n1952_n5888# 0.013418f
C576 drain_right.n217 a_n1952_n5888# 0.013034f
C577 drain_right.n218 a_n1952_n5888# 0.024256f
C578 drain_right.n219 a_n1952_n5888# 0.024256f
C579 drain_right.n220 a_n1952_n5888# 0.013034f
C580 drain_right.n221 a_n1952_n5888# 0.013801f
C581 drain_right.n222 a_n1952_n5888# 0.030808f
C582 drain_right.n223 a_n1952_n5888# 0.030808f
C583 drain_right.n224 a_n1952_n5888# 0.013801f
C584 drain_right.n225 a_n1952_n5888# 0.013034f
C585 drain_right.n226 a_n1952_n5888# 0.024256f
C586 drain_right.n227 a_n1952_n5888# 0.024256f
C587 drain_right.n228 a_n1952_n5888# 0.013034f
C588 drain_right.n229 a_n1952_n5888# 0.013801f
C589 drain_right.n230 a_n1952_n5888# 0.030808f
C590 drain_right.n231 a_n1952_n5888# 0.030808f
C591 drain_right.n232 a_n1952_n5888# 0.013801f
C592 drain_right.n233 a_n1952_n5888# 0.013034f
C593 drain_right.n234 a_n1952_n5888# 0.024256f
C594 drain_right.n235 a_n1952_n5888# 0.024256f
C595 drain_right.n236 a_n1952_n5888# 0.013034f
C596 drain_right.n237 a_n1952_n5888# 0.013801f
C597 drain_right.n238 a_n1952_n5888# 0.030808f
C598 drain_right.n239 a_n1952_n5888# 0.030808f
C599 drain_right.n240 a_n1952_n5888# 0.013801f
C600 drain_right.n241 a_n1952_n5888# 0.013034f
C601 drain_right.n242 a_n1952_n5888# 0.024256f
C602 drain_right.n243 a_n1952_n5888# 0.024256f
C603 drain_right.n244 a_n1952_n5888# 0.013034f
C604 drain_right.n245 a_n1952_n5888# 0.013801f
C605 drain_right.n246 a_n1952_n5888# 0.030808f
C606 drain_right.n247 a_n1952_n5888# 0.030808f
C607 drain_right.n248 a_n1952_n5888# 0.013801f
C608 drain_right.n249 a_n1952_n5888# 0.013034f
C609 drain_right.n250 a_n1952_n5888# 0.024256f
C610 drain_right.n251 a_n1952_n5888# 0.024256f
C611 drain_right.n252 a_n1952_n5888# 0.013034f
C612 drain_right.n253 a_n1952_n5888# 0.013801f
C613 drain_right.n254 a_n1952_n5888# 0.030808f
C614 drain_right.n255 a_n1952_n5888# 0.030808f
C615 drain_right.n256 a_n1952_n5888# 0.013801f
C616 drain_right.n257 a_n1952_n5888# 0.013034f
C617 drain_right.n258 a_n1952_n5888# 0.024256f
C618 drain_right.n259 a_n1952_n5888# 0.024256f
C619 drain_right.n260 a_n1952_n5888# 0.013034f
C620 drain_right.n261 a_n1952_n5888# 0.013418f
C621 drain_right.n262 a_n1952_n5888# 0.013418f
C622 drain_right.n263 a_n1952_n5888# 0.030808f
C623 drain_right.n264 a_n1952_n5888# 0.030808f
C624 drain_right.n265 a_n1952_n5888# 0.013801f
C625 drain_right.n266 a_n1952_n5888# 0.013034f
C626 drain_right.n267 a_n1952_n5888# 0.024256f
C627 drain_right.n268 a_n1952_n5888# 0.024256f
C628 drain_right.n269 a_n1952_n5888# 0.013034f
C629 drain_right.n270 a_n1952_n5888# 0.013801f
C630 drain_right.n271 a_n1952_n5888# 0.030808f
C631 drain_right.n272 a_n1952_n5888# 0.030808f
C632 drain_right.n273 a_n1952_n5888# 0.013801f
C633 drain_right.n274 a_n1952_n5888# 0.013034f
C634 drain_right.n275 a_n1952_n5888# 0.024256f
C635 drain_right.n276 a_n1952_n5888# 0.024256f
C636 drain_right.n277 a_n1952_n5888# 0.013034f
C637 drain_right.n278 a_n1952_n5888# 0.013801f
C638 drain_right.n279 a_n1952_n5888# 0.030808f
C639 drain_right.n280 a_n1952_n5888# 0.065537f
C640 drain_right.n281 a_n1952_n5888# 0.013801f
C641 drain_right.n282 a_n1952_n5888# 0.013034f
C642 drain_right.n283 a_n1952_n5888# 0.053417f
C643 drain_right.n284 a_n1952_n5888# 0.053239f
C644 drain_right.n285 a_n1952_n5888# 0.33752f
C645 source.n0 a_n1952_n5888# 0.033851f
C646 source.n1 a_n1952_n5888# 0.024555f
C647 source.n2 a_n1952_n5888# 0.013195f
C648 source.n3 a_n1952_n5888# 0.031187f
C649 source.n4 a_n1952_n5888# 0.013971f
C650 source.n5 a_n1952_n5888# 0.024555f
C651 source.n6 a_n1952_n5888# 0.013195f
C652 source.n7 a_n1952_n5888# 0.031187f
C653 source.n8 a_n1952_n5888# 0.013971f
C654 source.n9 a_n1952_n5888# 0.024555f
C655 source.n10 a_n1952_n5888# 0.013195f
C656 source.n11 a_n1952_n5888# 0.031187f
C657 source.n12 a_n1952_n5888# 0.013971f
C658 source.n13 a_n1952_n5888# 0.024555f
C659 source.n14 a_n1952_n5888# 0.013195f
C660 source.n15 a_n1952_n5888# 0.031187f
C661 source.n16 a_n1952_n5888# 0.031187f
C662 source.n17 a_n1952_n5888# 0.013971f
C663 source.n18 a_n1952_n5888# 0.024555f
C664 source.n19 a_n1952_n5888# 0.013195f
C665 source.n20 a_n1952_n5888# 0.031187f
C666 source.n21 a_n1952_n5888# 0.013971f
C667 source.n22 a_n1952_n5888# 0.024555f
C668 source.n23 a_n1952_n5888# 0.013195f
C669 source.n24 a_n1952_n5888# 0.031187f
C670 source.n25 a_n1952_n5888# 0.013971f
C671 source.n26 a_n1952_n5888# 0.024555f
C672 source.n27 a_n1952_n5888# 0.013195f
C673 source.n28 a_n1952_n5888# 0.031187f
C674 source.n29 a_n1952_n5888# 0.013971f
C675 source.n30 a_n1952_n5888# 0.024555f
C676 source.n31 a_n1952_n5888# 0.013195f
C677 source.n32 a_n1952_n5888# 0.031187f
C678 source.n33 a_n1952_n5888# 0.013971f
C679 source.n34 a_n1952_n5888# 0.024555f
C680 source.n35 a_n1952_n5888# 0.013583f
C681 source.n36 a_n1952_n5888# 0.031187f
C682 source.n37 a_n1952_n5888# 0.013195f
C683 source.n38 a_n1952_n5888# 0.013971f
C684 source.n39 a_n1952_n5888# 0.024555f
C685 source.n40 a_n1952_n5888# 0.013195f
C686 source.n41 a_n1952_n5888# 0.031187f
C687 source.n42 a_n1952_n5888# 0.013971f
C688 source.n43 a_n1952_n5888# 0.024555f
C689 source.n44 a_n1952_n5888# 0.013195f
C690 source.n45 a_n1952_n5888# 0.02339f
C691 source.n46 a_n1952_n5888# 0.022047f
C692 source.t5 a_n1952_n5888# 0.054392f
C693 source.n47 a_n1952_n5888# 0.299587f
C694 source.n48 a_n1952_n5888# 2.65854f
C695 source.n49 a_n1952_n5888# 0.013195f
C696 source.n50 a_n1952_n5888# 0.013971f
C697 source.n51 a_n1952_n5888# 0.031187f
C698 source.n52 a_n1952_n5888# 0.031187f
C699 source.n53 a_n1952_n5888# 0.013971f
C700 source.n54 a_n1952_n5888# 0.013195f
C701 source.n55 a_n1952_n5888# 0.024555f
C702 source.n56 a_n1952_n5888# 0.024555f
C703 source.n57 a_n1952_n5888# 0.013195f
C704 source.n58 a_n1952_n5888# 0.013971f
C705 source.n59 a_n1952_n5888# 0.031187f
C706 source.n60 a_n1952_n5888# 0.031187f
C707 source.n61 a_n1952_n5888# 0.013971f
C708 source.n62 a_n1952_n5888# 0.013195f
C709 source.n63 a_n1952_n5888# 0.024555f
C710 source.n64 a_n1952_n5888# 0.024555f
C711 source.n65 a_n1952_n5888# 0.013195f
C712 source.n66 a_n1952_n5888# 0.013971f
C713 source.n67 a_n1952_n5888# 0.031187f
C714 source.n68 a_n1952_n5888# 0.031187f
C715 source.n69 a_n1952_n5888# 0.031187f
C716 source.n70 a_n1952_n5888# 0.013583f
C717 source.n71 a_n1952_n5888# 0.013195f
C718 source.n72 a_n1952_n5888# 0.024555f
C719 source.n73 a_n1952_n5888# 0.024555f
C720 source.n74 a_n1952_n5888# 0.013195f
C721 source.n75 a_n1952_n5888# 0.013971f
C722 source.n76 a_n1952_n5888# 0.031187f
C723 source.n77 a_n1952_n5888# 0.031187f
C724 source.n78 a_n1952_n5888# 0.013971f
C725 source.n79 a_n1952_n5888# 0.013195f
C726 source.n80 a_n1952_n5888# 0.024555f
C727 source.n81 a_n1952_n5888# 0.024555f
C728 source.n82 a_n1952_n5888# 0.013195f
C729 source.n83 a_n1952_n5888# 0.013971f
C730 source.n84 a_n1952_n5888# 0.031187f
C731 source.n85 a_n1952_n5888# 0.031187f
C732 source.n86 a_n1952_n5888# 0.013971f
C733 source.n87 a_n1952_n5888# 0.013195f
C734 source.n88 a_n1952_n5888# 0.024555f
C735 source.n89 a_n1952_n5888# 0.024555f
C736 source.n90 a_n1952_n5888# 0.013195f
C737 source.n91 a_n1952_n5888# 0.013971f
C738 source.n92 a_n1952_n5888# 0.031187f
C739 source.n93 a_n1952_n5888# 0.031187f
C740 source.n94 a_n1952_n5888# 0.013971f
C741 source.n95 a_n1952_n5888# 0.013195f
C742 source.n96 a_n1952_n5888# 0.024555f
C743 source.n97 a_n1952_n5888# 0.024555f
C744 source.n98 a_n1952_n5888# 0.013195f
C745 source.n99 a_n1952_n5888# 0.013971f
C746 source.n100 a_n1952_n5888# 0.031187f
C747 source.n101 a_n1952_n5888# 0.031187f
C748 source.n102 a_n1952_n5888# 0.013971f
C749 source.n103 a_n1952_n5888# 0.013195f
C750 source.n104 a_n1952_n5888# 0.024555f
C751 source.n105 a_n1952_n5888# 0.024555f
C752 source.n106 a_n1952_n5888# 0.013195f
C753 source.n107 a_n1952_n5888# 0.013971f
C754 source.n108 a_n1952_n5888# 0.031187f
C755 source.n109 a_n1952_n5888# 0.031187f
C756 source.n110 a_n1952_n5888# 0.013971f
C757 source.n111 a_n1952_n5888# 0.013195f
C758 source.n112 a_n1952_n5888# 0.024555f
C759 source.n113 a_n1952_n5888# 0.024555f
C760 source.n114 a_n1952_n5888# 0.013195f
C761 source.n115 a_n1952_n5888# 0.013583f
C762 source.n116 a_n1952_n5888# 0.013583f
C763 source.n117 a_n1952_n5888# 0.031187f
C764 source.n118 a_n1952_n5888# 0.031187f
C765 source.n119 a_n1952_n5888# 0.013971f
C766 source.n120 a_n1952_n5888# 0.013195f
C767 source.n121 a_n1952_n5888# 0.024555f
C768 source.n122 a_n1952_n5888# 0.024555f
C769 source.n123 a_n1952_n5888# 0.013195f
C770 source.n124 a_n1952_n5888# 0.013971f
C771 source.n125 a_n1952_n5888# 0.031187f
C772 source.n126 a_n1952_n5888# 0.031187f
C773 source.n127 a_n1952_n5888# 0.013971f
C774 source.n128 a_n1952_n5888# 0.013195f
C775 source.n129 a_n1952_n5888# 0.024555f
C776 source.n130 a_n1952_n5888# 0.024555f
C777 source.n131 a_n1952_n5888# 0.013195f
C778 source.n132 a_n1952_n5888# 0.013971f
C779 source.n133 a_n1952_n5888# 0.031187f
C780 source.n134 a_n1952_n5888# 0.066343f
C781 source.n135 a_n1952_n5888# 0.013971f
C782 source.n136 a_n1952_n5888# 0.013195f
C783 source.n137 a_n1952_n5888# 0.054073f
C784 source.n138 a_n1952_n5888# 0.036917f
C785 source.n139 a_n1952_n5888# 1.97204f
C786 source.t8 a_n1952_n5888# 0.485095f
C787 source.t2 a_n1952_n5888# 0.485095f
C788 source.n140 a_n1952_n5888# 4.39018f
C789 source.n141 a_n1952_n5888# 0.395187f
C790 source.t0 a_n1952_n5888# 0.485095f
C791 source.t7 a_n1952_n5888# 0.485095f
C792 source.n142 a_n1952_n5888# 4.39018f
C793 source.n143 a_n1952_n5888# 0.397233f
C794 source.n144 a_n1952_n5888# 0.033851f
C795 source.n145 a_n1952_n5888# 0.024555f
C796 source.n146 a_n1952_n5888# 0.013195f
C797 source.n147 a_n1952_n5888# 0.031187f
C798 source.n148 a_n1952_n5888# 0.013971f
C799 source.n149 a_n1952_n5888# 0.024555f
C800 source.n150 a_n1952_n5888# 0.013195f
C801 source.n151 a_n1952_n5888# 0.031187f
C802 source.n152 a_n1952_n5888# 0.013971f
C803 source.n153 a_n1952_n5888# 0.024555f
C804 source.n154 a_n1952_n5888# 0.013195f
C805 source.n155 a_n1952_n5888# 0.031187f
C806 source.n156 a_n1952_n5888# 0.013971f
C807 source.n157 a_n1952_n5888# 0.024555f
C808 source.n158 a_n1952_n5888# 0.013195f
C809 source.n159 a_n1952_n5888# 0.031187f
C810 source.n160 a_n1952_n5888# 0.031187f
C811 source.n161 a_n1952_n5888# 0.013971f
C812 source.n162 a_n1952_n5888# 0.024555f
C813 source.n163 a_n1952_n5888# 0.013195f
C814 source.n164 a_n1952_n5888# 0.031187f
C815 source.n165 a_n1952_n5888# 0.013971f
C816 source.n166 a_n1952_n5888# 0.024555f
C817 source.n167 a_n1952_n5888# 0.013195f
C818 source.n168 a_n1952_n5888# 0.031187f
C819 source.n169 a_n1952_n5888# 0.013971f
C820 source.n170 a_n1952_n5888# 0.024555f
C821 source.n171 a_n1952_n5888# 0.013195f
C822 source.n172 a_n1952_n5888# 0.031187f
C823 source.n173 a_n1952_n5888# 0.013971f
C824 source.n174 a_n1952_n5888# 0.024555f
C825 source.n175 a_n1952_n5888# 0.013195f
C826 source.n176 a_n1952_n5888# 0.031187f
C827 source.n177 a_n1952_n5888# 0.013971f
C828 source.n178 a_n1952_n5888# 0.024555f
C829 source.n179 a_n1952_n5888# 0.013583f
C830 source.n180 a_n1952_n5888# 0.031187f
C831 source.n181 a_n1952_n5888# 0.013195f
C832 source.n182 a_n1952_n5888# 0.013971f
C833 source.n183 a_n1952_n5888# 0.024555f
C834 source.n184 a_n1952_n5888# 0.013195f
C835 source.n185 a_n1952_n5888# 0.031187f
C836 source.n186 a_n1952_n5888# 0.013971f
C837 source.n187 a_n1952_n5888# 0.024555f
C838 source.n188 a_n1952_n5888# 0.013195f
C839 source.n189 a_n1952_n5888# 0.02339f
C840 source.n190 a_n1952_n5888# 0.022047f
C841 source.t15 a_n1952_n5888# 0.054392f
C842 source.n191 a_n1952_n5888# 0.299587f
C843 source.n192 a_n1952_n5888# 2.65854f
C844 source.n193 a_n1952_n5888# 0.013195f
C845 source.n194 a_n1952_n5888# 0.013971f
C846 source.n195 a_n1952_n5888# 0.031187f
C847 source.n196 a_n1952_n5888# 0.031187f
C848 source.n197 a_n1952_n5888# 0.013971f
C849 source.n198 a_n1952_n5888# 0.013195f
C850 source.n199 a_n1952_n5888# 0.024555f
C851 source.n200 a_n1952_n5888# 0.024555f
C852 source.n201 a_n1952_n5888# 0.013195f
C853 source.n202 a_n1952_n5888# 0.013971f
C854 source.n203 a_n1952_n5888# 0.031187f
C855 source.n204 a_n1952_n5888# 0.031187f
C856 source.n205 a_n1952_n5888# 0.013971f
C857 source.n206 a_n1952_n5888# 0.013195f
C858 source.n207 a_n1952_n5888# 0.024555f
C859 source.n208 a_n1952_n5888# 0.024555f
C860 source.n209 a_n1952_n5888# 0.013195f
C861 source.n210 a_n1952_n5888# 0.013971f
C862 source.n211 a_n1952_n5888# 0.031187f
C863 source.n212 a_n1952_n5888# 0.031187f
C864 source.n213 a_n1952_n5888# 0.031187f
C865 source.n214 a_n1952_n5888# 0.013583f
C866 source.n215 a_n1952_n5888# 0.013195f
C867 source.n216 a_n1952_n5888# 0.024555f
C868 source.n217 a_n1952_n5888# 0.024555f
C869 source.n218 a_n1952_n5888# 0.013195f
C870 source.n219 a_n1952_n5888# 0.013971f
C871 source.n220 a_n1952_n5888# 0.031187f
C872 source.n221 a_n1952_n5888# 0.031187f
C873 source.n222 a_n1952_n5888# 0.013971f
C874 source.n223 a_n1952_n5888# 0.013195f
C875 source.n224 a_n1952_n5888# 0.024555f
C876 source.n225 a_n1952_n5888# 0.024555f
C877 source.n226 a_n1952_n5888# 0.013195f
C878 source.n227 a_n1952_n5888# 0.013971f
C879 source.n228 a_n1952_n5888# 0.031187f
C880 source.n229 a_n1952_n5888# 0.031187f
C881 source.n230 a_n1952_n5888# 0.013971f
C882 source.n231 a_n1952_n5888# 0.013195f
C883 source.n232 a_n1952_n5888# 0.024555f
C884 source.n233 a_n1952_n5888# 0.024555f
C885 source.n234 a_n1952_n5888# 0.013195f
C886 source.n235 a_n1952_n5888# 0.013971f
C887 source.n236 a_n1952_n5888# 0.031187f
C888 source.n237 a_n1952_n5888# 0.031187f
C889 source.n238 a_n1952_n5888# 0.013971f
C890 source.n239 a_n1952_n5888# 0.013195f
C891 source.n240 a_n1952_n5888# 0.024555f
C892 source.n241 a_n1952_n5888# 0.024555f
C893 source.n242 a_n1952_n5888# 0.013195f
C894 source.n243 a_n1952_n5888# 0.013971f
C895 source.n244 a_n1952_n5888# 0.031187f
C896 source.n245 a_n1952_n5888# 0.031187f
C897 source.n246 a_n1952_n5888# 0.013971f
C898 source.n247 a_n1952_n5888# 0.013195f
C899 source.n248 a_n1952_n5888# 0.024555f
C900 source.n249 a_n1952_n5888# 0.024555f
C901 source.n250 a_n1952_n5888# 0.013195f
C902 source.n251 a_n1952_n5888# 0.013971f
C903 source.n252 a_n1952_n5888# 0.031187f
C904 source.n253 a_n1952_n5888# 0.031187f
C905 source.n254 a_n1952_n5888# 0.013971f
C906 source.n255 a_n1952_n5888# 0.013195f
C907 source.n256 a_n1952_n5888# 0.024555f
C908 source.n257 a_n1952_n5888# 0.024555f
C909 source.n258 a_n1952_n5888# 0.013195f
C910 source.n259 a_n1952_n5888# 0.013583f
C911 source.n260 a_n1952_n5888# 0.013583f
C912 source.n261 a_n1952_n5888# 0.031187f
C913 source.n262 a_n1952_n5888# 0.031187f
C914 source.n263 a_n1952_n5888# 0.013971f
C915 source.n264 a_n1952_n5888# 0.013195f
C916 source.n265 a_n1952_n5888# 0.024555f
C917 source.n266 a_n1952_n5888# 0.024555f
C918 source.n267 a_n1952_n5888# 0.013195f
C919 source.n268 a_n1952_n5888# 0.013971f
C920 source.n269 a_n1952_n5888# 0.031187f
C921 source.n270 a_n1952_n5888# 0.031187f
C922 source.n271 a_n1952_n5888# 0.013971f
C923 source.n272 a_n1952_n5888# 0.013195f
C924 source.n273 a_n1952_n5888# 0.024555f
C925 source.n274 a_n1952_n5888# 0.024555f
C926 source.n275 a_n1952_n5888# 0.013195f
C927 source.n276 a_n1952_n5888# 0.013971f
C928 source.n277 a_n1952_n5888# 0.031187f
C929 source.n278 a_n1952_n5888# 0.066343f
C930 source.n279 a_n1952_n5888# 0.013971f
C931 source.n280 a_n1952_n5888# 0.013195f
C932 source.n281 a_n1952_n5888# 0.054073f
C933 source.n282 a_n1952_n5888# 0.036917f
C934 source.n283 a_n1952_n5888# 0.162012f
C935 source.t14 a_n1952_n5888# 0.485095f
C936 source.t17 a_n1952_n5888# 0.485095f
C937 source.n284 a_n1952_n5888# 4.39018f
C938 source.n285 a_n1952_n5888# 0.395187f
C939 source.t12 a_n1952_n5888# 0.485095f
C940 source.t10 a_n1952_n5888# 0.485095f
C941 source.n286 a_n1952_n5888# 4.39018f
C942 source.n287 a_n1952_n5888# 2.7441f
C943 source.t3 a_n1952_n5888# 0.485095f
C944 source.t9 a_n1952_n5888# 0.485095f
C945 source.n288 a_n1952_n5888# 4.39018f
C946 source.n289 a_n1952_n5888# 2.7441f
C947 source.t4 a_n1952_n5888# 0.485095f
C948 source.t1 a_n1952_n5888# 0.485095f
C949 source.n290 a_n1952_n5888# 4.39018f
C950 source.n291 a_n1952_n5888# 0.395189f
C951 source.n292 a_n1952_n5888# 0.033851f
C952 source.n293 a_n1952_n5888# 0.024555f
C953 source.n294 a_n1952_n5888# 0.013195f
C954 source.n295 a_n1952_n5888# 0.031187f
C955 source.n296 a_n1952_n5888# 0.013971f
C956 source.n297 a_n1952_n5888# 0.024555f
C957 source.n298 a_n1952_n5888# 0.013195f
C958 source.n299 a_n1952_n5888# 0.031187f
C959 source.n300 a_n1952_n5888# 0.013971f
C960 source.n301 a_n1952_n5888# 0.024555f
C961 source.n302 a_n1952_n5888# 0.013195f
C962 source.n303 a_n1952_n5888# 0.031187f
C963 source.n304 a_n1952_n5888# 0.013971f
C964 source.n305 a_n1952_n5888# 0.024555f
C965 source.n306 a_n1952_n5888# 0.013195f
C966 source.n307 a_n1952_n5888# 0.031187f
C967 source.n308 a_n1952_n5888# 0.013971f
C968 source.n309 a_n1952_n5888# 0.024555f
C969 source.n310 a_n1952_n5888# 0.013195f
C970 source.n311 a_n1952_n5888# 0.031187f
C971 source.n312 a_n1952_n5888# 0.013971f
C972 source.n313 a_n1952_n5888# 0.024555f
C973 source.n314 a_n1952_n5888# 0.013195f
C974 source.n315 a_n1952_n5888# 0.031187f
C975 source.n316 a_n1952_n5888# 0.013971f
C976 source.n317 a_n1952_n5888# 0.024555f
C977 source.n318 a_n1952_n5888# 0.013195f
C978 source.n319 a_n1952_n5888# 0.031187f
C979 source.n320 a_n1952_n5888# 0.013971f
C980 source.n321 a_n1952_n5888# 0.024555f
C981 source.n322 a_n1952_n5888# 0.013195f
C982 source.n323 a_n1952_n5888# 0.031187f
C983 source.n324 a_n1952_n5888# 0.013971f
C984 source.n325 a_n1952_n5888# 0.024555f
C985 source.n326 a_n1952_n5888# 0.013583f
C986 source.n327 a_n1952_n5888# 0.031187f
C987 source.n328 a_n1952_n5888# 0.013971f
C988 source.n329 a_n1952_n5888# 0.024555f
C989 source.n330 a_n1952_n5888# 0.013195f
C990 source.n331 a_n1952_n5888# 0.031187f
C991 source.n332 a_n1952_n5888# 0.013971f
C992 source.n333 a_n1952_n5888# 0.024555f
C993 source.n334 a_n1952_n5888# 0.013195f
C994 source.n335 a_n1952_n5888# 0.02339f
C995 source.n336 a_n1952_n5888# 0.022047f
C996 source.t6 a_n1952_n5888# 0.054392f
C997 source.n337 a_n1952_n5888# 0.299587f
C998 source.n338 a_n1952_n5888# 2.65854f
C999 source.n339 a_n1952_n5888# 0.013195f
C1000 source.n340 a_n1952_n5888# 0.013971f
C1001 source.n341 a_n1952_n5888# 0.031187f
C1002 source.n342 a_n1952_n5888# 0.031187f
C1003 source.n343 a_n1952_n5888# 0.013971f
C1004 source.n344 a_n1952_n5888# 0.013195f
C1005 source.n345 a_n1952_n5888# 0.024555f
C1006 source.n346 a_n1952_n5888# 0.024555f
C1007 source.n347 a_n1952_n5888# 0.013195f
C1008 source.n348 a_n1952_n5888# 0.013971f
C1009 source.n349 a_n1952_n5888# 0.031187f
C1010 source.n350 a_n1952_n5888# 0.031187f
C1011 source.n351 a_n1952_n5888# 0.013971f
C1012 source.n352 a_n1952_n5888# 0.013195f
C1013 source.n353 a_n1952_n5888# 0.024555f
C1014 source.n354 a_n1952_n5888# 0.024555f
C1015 source.n355 a_n1952_n5888# 0.013195f
C1016 source.n356 a_n1952_n5888# 0.013195f
C1017 source.n357 a_n1952_n5888# 0.013971f
C1018 source.n358 a_n1952_n5888# 0.031187f
C1019 source.n359 a_n1952_n5888# 0.031187f
C1020 source.n360 a_n1952_n5888# 0.031187f
C1021 source.n361 a_n1952_n5888# 0.013583f
C1022 source.n362 a_n1952_n5888# 0.013195f
C1023 source.n363 a_n1952_n5888# 0.024555f
C1024 source.n364 a_n1952_n5888# 0.024555f
C1025 source.n365 a_n1952_n5888# 0.013195f
C1026 source.n366 a_n1952_n5888# 0.013971f
C1027 source.n367 a_n1952_n5888# 0.031187f
C1028 source.n368 a_n1952_n5888# 0.031187f
C1029 source.n369 a_n1952_n5888# 0.013971f
C1030 source.n370 a_n1952_n5888# 0.013195f
C1031 source.n371 a_n1952_n5888# 0.024555f
C1032 source.n372 a_n1952_n5888# 0.024555f
C1033 source.n373 a_n1952_n5888# 0.013195f
C1034 source.n374 a_n1952_n5888# 0.013971f
C1035 source.n375 a_n1952_n5888# 0.031187f
C1036 source.n376 a_n1952_n5888# 0.031187f
C1037 source.n377 a_n1952_n5888# 0.013971f
C1038 source.n378 a_n1952_n5888# 0.013195f
C1039 source.n379 a_n1952_n5888# 0.024555f
C1040 source.n380 a_n1952_n5888# 0.024555f
C1041 source.n381 a_n1952_n5888# 0.013195f
C1042 source.n382 a_n1952_n5888# 0.013971f
C1043 source.n383 a_n1952_n5888# 0.031187f
C1044 source.n384 a_n1952_n5888# 0.031187f
C1045 source.n385 a_n1952_n5888# 0.013971f
C1046 source.n386 a_n1952_n5888# 0.013195f
C1047 source.n387 a_n1952_n5888# 0.024555f
C1048 source.n388 a_n1952_n5888# 0.024555f
C1049 source.n389 a_n1952_n5888# 0.013195f
C1050 source.n390 a_n1952_n5888# 0.013971f
C1051 source.n391 a_n1952_n5888# 0.031187f
C1052 source.n392 a_n1952_n5888# 0.031187f
C1053 source.n393 a_n1952_n5888# 0.013971f
C1054 source.n394 a_n1952_n5888# 0.013195f
C1055 source.n395 a_n1952_n5888# 0.024555f
C1056 source.n396 a_n1952_n5888# 0.024555f
C1057 source.n397 a_n1952_n5888# 0.013195f
C1058 source.n398 a_n1952_n5888# 0.013971f
C1059 source.n399 a_n1952_n5888# 0.031187f
C1060 source.n400 a_n1952_n5888# 0.031187f
C1061 source.n401 a_n1952_n5888# 0.031187f
C1062 source.n402 a_n1952_n5888# 0.013971f
C1063 source.n403 a_n1952_n5888# 0.013195f
C1064 source.n404 a_n1952_n5888# 0.024555f
C1065 source.n405 a_n1952_n5888# 0.024555f
C1066 source.n406 a_n1952_n5888# 0.013195f
C1067 source.n407 a_n1952_n5888# 0.013583f
C1068 source.n408 a_n1952_n5888# 0.013583f
C1069 source.n409 a_n1952_n5888# 0.031187f
C1070 source.n410 a_n1952_n5888# 0.031187f
C1071 source.n411 a_n1952_n5888# 0.013971f
C1072 source.n412 a_n1952_n5888# 0.013195f
C1073 source.n413 a_n1952_n5888# 0.024555f
C1074 source.n414 a_n1952_n5888# 0.024555f
C1075 source.n415 a_n1952_n5888# 0.013195f
C1076 source.n416 a_n1952_n5888# 0.013971f
C1077 source.n417 a_n1952_n5888# 0.031187f
C1078 source.n418 a_n1952_n5888# 0.031187f
C1079 source.n419 a_n1952_n5888# 0.013971f
C1080 source.n420 a_n1952_n5888# 0.013195f
C1081 source.n421 a_n1952_n5888# 0.024555f
C1082 source.n422 a_n1952_n5888# 0.024555f
C1083 source.n423 a_n1952_n5888# 0.013195f
C1084 source.n424 a_n1952_n5888# 0.013971f
C1085 source.n425 a_n1952_n5888# 0.031187f
C1086 source.n426 a_n1952_n5888# 0.066343f
C1087 source.n427 a_n1952_n5888# 0.013971f
C1088 source.n428 a_n1952_n5888# 0.013195f
C1089 source.n429 a_n1952_n5888# 0.054073f
C1090 source.n430 a_n1952_n5888# 0.036917f
C1091 source.n431 a_n1952_n5888# 0.162012f
C1092 source.t13 a_n1952_n5888# 0.485095f
C1093 source.t11 a_n1952_n5888# 0.485095f
C1094 source.n432 a_n1952_n5888# 4.39018f
C1095 source.n433 a_n1952_n5888# 0.397235f
C1096 source.t19 a_n1952_n5888# 0.485095f
C1097 source.t18 a_n1952_n5888# 0.485095f
C1098 source.n434 a_n1952_n5888# 4.39018f
C1099 source.n435 a_n1952_n5888# 0.395189f
C1100 source.n436 a_n1952_n5888# 0.033851f
C1101 source.n437 a_n1952_n5888# 0.024555f
C1102 source.n438 a_n1952_n5888# 0.013195f
C1103 source.n439 a_n1952_n5888# 0.031187f
C1104 source.n440 a_n1952_n5888# 0.013971f
C1105 source.n441 a_n1952_n5888# 0.024555f
C1106 source.n442 a_n1952_n5888# 0.013195f
C1107 source.n443 a_n1952_n5888# 0.031187f
C1108 source.n444 a_n1952_n5888# 0.013971f
C1109 source.n445 a_n1952_n5888# 0.024555f
C1110 source.n446 a_n1952_n5888# 0.013195f
C1111 source.n447 a_n1952_n5888# 0.031187f
C1112 source.n448 a_n1952_n5888# 0.013971f
C1113 source.n449 a_n1952_n5888# 0.024555f
C1114 source.n450 a_n1952_n5888# 0.013195f
C1115 source.n451 a_n1952_n5888# 0.031187f
C1116 source.n452 a_n1952_n5888# 0.013971f
C1117 source.n453 a_n1952_n5888# 0.024555f
C1118 source.n454 a_n1952_n5888# 0.013195f
C1119 source.n455 a_n1952_n5888# 0.031187f
C1120 source.n456 a_n1952_n5888# 0.013971f
C1121 source.n457 a_n1952_n5888# 0.024555f
C1122 source.n458 a_n1952_n5888# 0.013195f
C1123 source.n459 a_n1952_n5888# 0.031187f
C1124 source.n460 a_n1952_n5888# 0.013971f
C1125 source.n461 a_n1952_n5888# 0.024555f
C1126 source.n462 a_n1952_n5888# 0.013195f
C1127 source.n463 a_n1952_n5888# 0.031187f
C1128 source.n464 a_n1952_n5888# 0.013971f
C1129 source.n465 a_n1952_n5888# 0.024555f
C1130 source.n466 a_n1952_n5888# 0.013195f
C1131 source.n467 a_n1952_n5888# 0.031187f
C1132 source.n468 a_n1952_n5888# 0.013971f
C1133 source.n469 a_n1952_n5888# 0.024555f
C1134 source.n470 a_n1952_n5888# 0.013583f
C1135 source.n471 a_n1952_n5888# 0.031187f
C1136 source.n472 a_n1952_n5888# 0.013971f
C1137 source.n473 a_n1952_n5888# 0.024555f
C1138 source.n474 a_n1952_n5888# 0.013195f
C1139 source.n475 a_n1952_n5888# 0.031187f
C1140 source.n476 a_n1952_n5888# 0.013971f
C1141 source.n477 a_n1952_n5888# 0.024555f
C1142 source.n478 a_n1952_n5888# 0.013195f
C1143 source.n479 a_n1952_n5888# 0.02339f
C1144 source.n480 a_n1952_n5888# 0.022047f
C1145 source.t16 a_n1952_n5888# 0.054392f
C1146 source.n481 a_n1952_n5888# 0.299587f
C1147 source.n482 a_n1952_n5888# 2.65854f
C1148 source.n483 a_n1952_n5888# 0.013195f
C1149 source.n484 a_n1952_n5888# 0.013971f
C1150 source.n485 a_n1952_n5888# 0.031187f
C1151 source.n486 a_n1952_n5888# 0.031187f
C1152 source.n487 a_n1952_n5888# 0.013971f
C1153 source.n488 a_n1952_n5888# 0.013195f
C1154 source.n489 a_n1952_n5888# 0.024555f
C1155 source.n490 a_n1952_n5888# 0.024555f
C1156 source.n491 a_n1952_n5888# 0.013195f
C1157 source.n492 a_n1952_n5888# 0.013971f
C1158 source.n493 a_n1952_n5888# 0.031187f
C1159 source.n494 a_n1952_n5888# 0.031187f
C1160 source.n495 a_n1952_n5888# 0.013971f
C1161 source.n496 a_n1952_n5888# 0.013195f
C1162 source.n497 a_n1952_n5888# 0.024555f
C1163 source.n498 a_n1952_n5888# 0.024555f
C1164 source.n499 a_n1952_n5888# 0.013195f
C1165 source.n500 a_n1952_n5888# 0.013195f
C1166 source.n501 a_n1952_n5888# 0.013971f
C1167 source.n502 a_n1952_n5888# 0.031187f
C1168 source.n503 a_n1952_n5888# 0.031187f
C1169 source.n504 a_n1952_n5888# 0.031187f
C1170 source.n505 a_n1952_n5888# 0.013583f
C1171 source.n506 a_n1952_n5888# 0.013195f
C1172 source.n507 a_n1952_n5888# 0.024555f
C1173 source.n508 a_n1952_n5888# 0.024555f
C1174 source.n509 a_n1952_n5888# 0.013195f
C1175 source.n510 a_n1952_n5888# 0.013971f
C1176 source.n511 a_n1952_n5888# 0.031187f
C1177 source.n512 a_n1952_n5888# 0.031187f
C1178 source.n513 a_n1952_n5888# 0.013971f
C1179 source.n514 a_n1952_n5888# 0.013195f
C1180 source.n515 a_n1952_n5888# 0.024555f
C1181 source.n516 a_n1952_n5888# 0.024555f
C1182 source.n517 a_n1952_n5888# 0.013195f
C1183 source.n518 a_n1952_n5888# 0.013971f
C1184 source.n519 a_n1952_n5888# 0.031187f
C1185 source.n520 a_n1952_n5888# 0.031187f
C1186 source.n521 a_n1952_n5888# 0.013971f
C1187 source.n522 a_n1952_n5888# 0.013195f
C1188 source.n523 a_n1952_n5888# 0.024555f
C1189 source.n524 a_n1952_n5888# 0.024555f
C1190 source.n525 a_n1952_n5888# 0.013195f
C1191 source.n526 a_n1952_n5888# 0.013971f
C1192 source.n527 a_n1952_n5888# 0.031187f
C1193 source.n528 a_n1952_n5888# 0.031187f
C1194 source.n529 a_n1952_n5888# 0.013971f
C1195 source.n530 a_n1952_n5888# 0.013195f
C1196 source.n531 a_n1952_n5888# 0.024555f
C1197 source.n532 a_n1952_n5888# 0.024555f
C1198 source.n533 a_n1952_n5888# 0.013195f
C1199 source.n534 a_n1952_n5888# 0.013971f
C1200 source.n535 a_n1952_n5888# 0.031187f
C1201 source.n536 a_n1952_n5888# 0.031187f
C1202 source.n537 a_n1952_n5888# 0.013971f
C1203 source.n538 a_n1952_n5888# 0.013195f
C1204 source.n539 a_n1952_n5888# 0.024555f
C1205 source.n540 a_n1952_n5888# 0.024555f
C1206 source.n541 a_n1952_n5888# 0.013195f
C1207 source.n542 a_n1952_n5888# 0.013971f
C1208 source.n543 a_n1952_n5888# 0.031187f
C1209 source.n544 a_n1952_n5888# 0.031187f
C1210 source.n545 a_n1952_n5888# 0.031187f
C1211 source.n546 a_n1952_n5888# 0.013971f
C1212 source.n547 a_n1952_n5888# 0.013195f
C1213 source.n548 a_n1952_n5888# 0.024555f
C1214 source.n549 a_n1952_n5888# 0.024555f
C1215 source.n550 a_n1952_n5888# 0.013195f
C1216 source.n551 a_n1952_n5888# 0.013583f
C1217 source.n552 a_n1952_n5888# 0.013583f
C1218 source.n553 a_n1952_n5888# 0.031187f
C1219 source.n554 a_n1952_n5888# 0.031187f
C1220 source.n555 a_n1952_n5888# 0.013971f
C1221 source.n556 a_n1952_n5888# 0.013195f
C1222 source.n557 a_n1952_n5888# 0.024555f
C1223 source.n558 a_n1952_n5888# 0.024555f
C1224 source.n559 a_n1952_n5888# 0.013195f
C1225 source.n560 a_n1952_n5888# 0.013971f
C1226 source.n561 a_n1952_n5888# 0.031187f
C1227 source.n562 a_n1952_n5888# 0.031187f
C1228 source.n563 a_n1952_n5888# 0.013971f
C1229 source.n564 a_n1952_n5888# 0.013195f
C1230 source.n565 a_n1952_n5888# 0.024555f
C1231 source.n566 a_n1952_n5888# 0.024555f
C1232 source.n567 a_n1952_n5888# 0.013195f
C1233 source.n568 a_n1952_n5888# 0.013971f
C1234 source.n569 a_n1952_n5888# 0.031187f
C1235 source.n570 a_n1952_n5888# 0.066343f
C1236 source.n571 a_n1952_n5888# 0.013971f
C1237 source.n572 a_n1952_n5888# 0.013195f
C1238 source.n573 a_n1952_n5888# 0.054073f
C1239 source.n574 a_n1952_n5888# 0.036917f
C1240 source.n575 a_n1952_n5888# 0.287056f
C1241 source.n576 a_n1952_n5888# 2.63561f
C1242 minus.n0 a_n1952_n5888# 0.042213f
C1243 minus.n1 a_n1952_n5888# 0.009579f
C1244 minus.t9 a_n1952_n5888# 2.08764f
C1245 minus.n2 a_n1952_n5888# 0.176314f
C1246 minus.t8 a_n1952_n5888# 2.10609f
C1247 minus.n3 a_n1952_n5888# 0.747494f
C1248 minus.t2 a_n1952_n5888# 2.08764f
C1249 minus.n4 a_n1952_n5888# 0.766346f
C1250 minus.n5 a_n1952_n5888# 0.009579f
C1251 minus.t7 a_n1952_n5888# 2.08764f
C1252 minus.n6 a_n1952_n5888# 0.762093f
C1253 minus.n7 a_n1952_n5888# 0.042213f
C1254 minus.n8 a_n1952_n5888# 0.042213f
C1255 minus.n9 a_n1952_n5888# 0.042213f
C1256 minus.n10 a_n1952_n5888# 0.762093f
C1257 minus.n11 a_n1952_n5888# 0.009579f
C1258 minus.t6 a_n1952_n5888# 2.08764f
C1259 minus.n12 a_n1952_n5888# 0.759751f
C1260 minus.n13 a_n1952_n5888# 2.16945f
C1261 minus.n14 a_n1952_n5888# 0.042213f
C1262 minus.n15 a_n1952_n5888# 0.009579f
C1263 minus.n16 a_n1952_n5888# 0.176314f
C1264 minus.t5 a_n1952_n5888# 2.10609f
C1265 minus.n17 a_n1952_n5888# 0.747494f
C1266 minus.t4 a_n1952_n5888# 2.08764f
C1267 minus.n18 a_n1952_n5888# 0.766346f
C1268 minus.n19 a_n1952_n5888# 0.009579f
C1269 minus.t0 a_n1952_n5888# 2.08764f
C1270 minus.n20 a_n1952_n5888# 0.762093f
C1271 minus.n21 a_n1952_n5888# 0.042213f
C1272 minus.n22 a_n1952_n5888# 0.042213f
C1273 minus.n23 a_n1952_n5888# 0.042213f
C1274 minus.t1 a_n1952_n5888# 2.08764f
C1275 minus.n24 a_n1952_n5888# 0.762093f
C1276 minus.n25 a_n1952_n5888# 0.009579f
C1277 minus.t3 a_n1952_n5888# 2.08764f
C1278 minus.n26 a_n1952_n5888# 0.759751f
C1279 minus.n27 a_n1952_n5888# 0.289686f
C1280 minus.n28 a_n1952_n5888# 2.5565f
.ends

