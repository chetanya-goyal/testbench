* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right minus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X1 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X2 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X3 source plus drain_left a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5 source minus drain_right a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7 drain_left plus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X8 source minus drain_right a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X9 drain_right minus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X10 drain_right minus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X11 drain_left plus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X12 drain_right minus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X13 drain_left plus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X14 source plus drain_left a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X15 drain_left plus source a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
.ends

