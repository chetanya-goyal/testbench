* NGSPICE file created from diffpair79.ext - technology: sky130A

.subckt diffpair79 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t31 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X1 drain_right.t22 minus.t1 source.t33 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X2 source.t10 plus.t0 drain_left.t23 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X3 a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X4 a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X5 source.t32 minus.t2 drain_right.t21 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X6 source.t24 minus.t3 drain_right.t20 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X7 drain_left.t22 plus.t1 source.t23 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_left.t21 plus.t2 source.t19 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X9 drain_left.t20 plus.t3 source.t8 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X10 source.t43 minus.t4 drain_right.t19 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X11 source.t47 minus.t5 drain_right.t18 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X12 source.t30 minus.t6 drain_right.t17 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X13 source.t45 minus.t7 drain_right.t16 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X14 drain_left.t19 plus.t4 source.t18 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X15 drain_left.t18 plus.t5 source.t22 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X16 source.t5 plus.t6 drain_left.t17 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X17 drain_right.t15 minus.t8 source.t41 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_left.t16 plus.t7 source.t21 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X19 drain_left.t15 plus.t8 source.t7 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X20 drain_left.t14 plus.t9 source.t14 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 source.t28 minus.t9 drain_right.t14 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 source.t46 minus.t10 drain_right.t13 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X23 drain_right.t12 minus.t11 source.t37 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X24 drain_right.t11 minus.t12 source.t29 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X25 drain_right.t10 minus.t13 source.t40 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X26 source.t17 plus.t10 drain_left.t13 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X27 source.t38 minus.t14 drain_right.t9 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X28 source.t36 minus.t15 drain_right.t8 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X29 drain_left.t12 plus.t11 source.t4 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X30 source.t25 minus.t16 drain_right.t7 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X31 drain_right.t6 minus.t17 source.t44 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X32 source.t1 plus.t12 drain_left.t11 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X33 drain_right.t5 minus.t18 source.t26 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X34 source.t3 plus.t13 drain_left.t10 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X35 a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X36 drain_left.t9 plus.t14 source.t6 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X37 drain_left.t8 plus.t15 source.t13 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X38 source.t39 minus.t19 drain_right.t4 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X39 drain_right.t3 minus.t20 source.t27 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X40 drain_right.t2 minus.t21 source.t34 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X41 source.t16 plus.t16 drain_left.t7 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X42 source.t0 plus.t17 drain_left.t6 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X43 source.t20 plus.t18 drain_left.t5 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X44 drain_left.t4 plus.t19 source.t2 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X45 drain_right.t1 minus.t22 source.t35 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X46 a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X47 drain_right.t0 minus.t23 source.t42 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X48 source.t12 plus.t20 drain_left.t3 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X49 source.t15 plus.t21 drain_left.t2 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X50 source.t9 plus.t22 drain_left.t1 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X51 source.t11 plus.t23 drain_left.t0 a_n3654_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n35 minus.n34 161.3
R1 minus.n33 minus.n0 161.3
R2 minus.n29 minus.n28 161.3
R3 minus.n27 minus.n2 161.3
R4 minus.n26 minus.n25 161.3
R5 minus.n24 minus.n3 161.3
R6 minus.n23 minus.n22 161.3
R7 minus.n18 minus.n5 161.3
R8 minus.n17 minus.n16 161.3
R9 minus.n15 minus.n6 161.3
R10 minus.n14 minus.n13 161.3
R11 minus.n12 minus.n7 161.3
R12 minus.n71 minus.n70 161.3
R13 minus.n69 minus.n36 161.3
R14 minus.n65 minus.n64 161.3
R15 minus.n63 minus.n38 161.3
R16 minus.n62 minus.n61 161.3
R17 minus.n60 minus.n39 161.3
R18 minus.n59 minus.n58 161.3
R19 minus.n54 minus.n41 161.3
R20 minus.n53 minus.n52 161.3
R21 minus.n51 minus.n42 161.3
R22 minus.n50 minus.n49 161.3
R23 minus.n48 minus.n43 161.3
R24 minus.n8 minus.t13 100.665
R25 minus.n44 minus.t7 100.665
R26 minus.n32 minus.n31 80.6037
R27 minus.n30 minus.n1 80.6037
R28 minus.n21 minus.n4 80.6037
R29 minus.n20 minus.n19 80.6037
R30 minus.n11 minus.n10 80.6037
R31 minus.n68 minus.n67 80.6037
R32 minus.n66 minus.n37 80.6037
R33 minus.n57 minus.n40 80.6037
R34 minus.n56 minus.n55 80.6037
R35 minus.n47 minus.n46 80.6037
R36 minus.n9 minus.t9 79.2293
R37 minus.n10 minus.t8 79.2293
R38 minus.n14 minus.t16 79.2293
R39 minus.n16 minus.t18 79.2293
R40 minus.n20 minus.t14 79.2293
R41 minus.n21 minus.t11 79.2293
R42 minus.n3 minus.t19 79.2293
R43 minus.n27 minus.t17 79.2293
R44 minus.n1 minus.t5 79.2293
R45 minus.n32 minus.t12 79.2293
R46 minus.n34 minus.t10 79.2293
R47 minus.n45 minus.t21 79.2293
R48 minus.n46 minus.t6 79.2293
R49 minus.n50 minus.t20 79.2293
R50 minus.n52 minus.t3 79.2293
R51 minus.n56 minus.t22 79.2293
R52 minus.n57 minus.t2 79.2293
R53 minus.n39 minus.t23 79.2293
R54 minus.n63 minus.t4 79.2293
R55 minus.n37 minus.t0 79.2293
R56 minus.n68 minus.t15 79.2293
R57 minus.n70 minus.t1 79.2293
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n20 minus.n5 41.6278
R69 minus.n22 minus.n21 41.6278
R70 minus.n56 minus.n41 41.6278
R71 minus.n58 minus.n57 41.6278
R72 minus.n33 minus.n32 38.7066
R73 minus.n69 minus.n68 38.7066
R74 minus.n72 minus.n35 34.7884
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 source.n0 source.t18 243.255
R132 source.n11 source.t15 243.255
R133 source.n12 source.t40 243.255
R134 source.n23 source.t46 243.255
R135 source.n47 source.t33 243.254
R136 source.n36 source.t45 243.254
R137 source.n35 source.t21 243.254
R138 source.n24 source.t0 243.254
R139 source.n2 source.n1 223.454
R140 source.n4 source.n3 223.454
R141 source.n6 source.n5 223.454
R142 source.n8 source.n7 223.454
R143 source.n10 source.n9 223.454
R144 source.n14 source.n13 223.454
R145 source.n16 source.n15 223.454
R146 source.n18 source.n17 223.454
R147 source.n20 source.n19 223.454
R148 source.n22 source.n21 223.454
R149 source.n46 source.n45 223.453
R150 source.n44 source.n43 223.453
R151 source.n42 source.n41 223.453
R152 source.n40 source.n39 223.453
R153 source.n38 source.n37 223.453
R154 source.n34 source.n33 223.453
R155 source.n32 source.n31 223.453
R156 source.n30 source.n29 223.453
R157 source.n28 source.n27 223.453
R158 source.n26 source.n25 223.453
R159 source.n45 source.t31 19.8005
R160 source.n45 source.t36 19.8005
R161 source.n43 source.t42 19.8005
R162 source.n43 source.t43 19.8005
R163 source.n41 source.t35 19.8005
R164 source.n41 source.t32 19.8005
R165 source.n39 source.t27 19.8005
R166 source.n39 source.t24 19.8005
R167 source.n37 source.t34 19.8005
R168 source.n37 source.t30 19.8005
R169 source.n33 source.t7 19.8005
R170 source.n33 source.t12 19.8005
R171 source.n31 source.t23 19.8005
R172 source.n31 source.t9 19.8005
R173 source.n29 source.t19 19.8005
R174 source.n29 source.t11 19.8005
R175 source.n27 source.t8 19.8005
R176 source.n27 source.t1 19.8005
R177 source.n25 source.t22 19.8005
R178 source.n25 source.t10 19.8005
R179 source.n1 source.t14 19.8005
R180 source.n1 source.t5 19.8005
R181 source.n3 source.t4 19.8005
R182 source.n3 source.t17 19.8005
R183 source.n5 source.t6 19.8005
R184 source.n5 source.t3 19.8005
R185 source.n7 source.t13 19.8005
R186 source.n7 source.t20 19.8005
R187 source.n9 source.t2 19.8005
R188 source.n9 source.t16 19.8005
R189 source.n13 source.t41 19.8005
R190 source.n13 source.t28 19.8005
R191 source.n15 source.t26 19.8005
R192 source.n15 source.t25 19.8005
R193 source.n17 source.t37 19.8005
R194 source.n17 source.t38 19.8005
R195 source.n19 source.t44 19.8005
R196 source.n19 source.t39 19.8005
R197 source.n21 source.t29 19.8005
R198 source.n21 source.t47 19.8005
R199 source.n24 source.n23 13.9285
R200 source.n48 source.n0 8.17853
R201 source.n48 source.n47 5.7505
R202 source.n23 source.n22 0.974638
R203 source.n22 source.n20 0.974638
R204 source.n20 source.n18 0.974638
R205 source.n18 source.n16 0.974638
R206 source.n16 source.n14 0.974638
R207 source.n14 source.n12 0.974638
R208 source.n11 source.n10 0.974638
R209 source.n10 source.n8 0.974638
R210 source.n8 source.n6 0.974638
R211 source.n6 source.n4 0.974638
R212 source.n4 source.n2 0.974638
R213 source.n2 source.n0 0.974638
R214 source.n26 source.n24 0.974638
R215 source.n28 source.n26 0.974638
R216 source.n30 source.n28 0.974638
R217 source.n32 source.n30 0.974638
R218 source.n34 source.n32 0.974638
R219 source.n35 source.n34 0.974638
R220 source.n38 source.n36 0.974638
R221 source.n40 source.n38 0.974638
R222 source.n42 source.n40 0.974638
R223 source.n44 source.n42 0.974638
R224 source.n46 source.n44 0.974638
R225 source.n47 source.n46 0.974638
R226 source.n12 source.n11 0.470328
R227 source.n36 source.n35 0.470328
R228 source source.n48 0.188
R229 drain_right.n13 drain_right.n11 241.107
R230 drain_right.n7 drain_right.n5 241.106
R231 drain_right.n2 drain_right.n0 241.106
R232 drain_right.n13 drain_right.n12 240.132
R233 drain_right.n15 drain_right.n14 240.132
R234 drain_right.n17 drain_right.n16 240.132
R235 drain_right.n19 drain_right.n18 240.132
R236 drain_right.n21 drain_right.n20 240.132
R237 drain_right.n7 drain_right.n6 240.131
R238 drain_right.n9 drain_right.n8 240.131
R239 drain_right.n4 drain_right.n3 240.131
R240 drain_right.n2 drain_right.n1 240.131
R241 drain_right drain_right.n10 27.7348
R242 drain_right.n5 drain_right.t8 19.8005
R243 drain_right.n5 drain_right.t22 19.8005
R244 drain_right.n6 drain_right.t19 19.8005
R245 drain_right.n6 drain_right.t23 19.8005
R246 drain_right.n8 drain_right.t21 19.8005
R247 drain_right.n8 drain_right.t0 19.8005
R248 drain_right.n3 drain_right.t20 19.8005
R249 drain_right.n3 drain_right.t1 19.8005
R250 drain_right.n1 drain_right.t17 19.8005
R251 drain_right.n1 drain_right.t3 19.8005
R252 drain_right.n0 drain_right.t16 19.8005
R253 drain_right.n0 drain_right.t2 19.8005
R254 drain_right.n11 drain_right.t14 19.8005
R255 drain_right.n11 drain_right.t10 19.8005
R256 drain_right.n12 drain_right.t7 19.8005
R257 drain_right.n12 drain_right.t15 19.8005
R258 drain_right.n14 drain_right.t9 19.8005
R259 drain_right.n14 drain_right.t5 19.8005
R260 drain_right.n16 drain_right.t4 19.8005
R261 drain_right.n16 drain_right.t12 19.8005
R262 drain_right.n18 drain_right.t18 19.8005
R263 drain_right.n18 drain_right.t6 19.8005
R264 drain_right.n20 drain_right.t13 19.8005
R265 drain_right.n20 drain_right.t11 19.8005
R266 drain_right drain_right.n21 6.62735
R267 drain_right.n9 drain_right.n7 0.974638
R268 drain_right.n4 drain_right.n2 0.974638
R269 drain_right.n21 drain_right.n19 0.974638
R270 drain_right.n19 drain_right.n17 0.974638
R271 drain_right.n17 drain_right.n15 0.974638
R272 drain_right.n15 drain_right.n13 0.974638
R273 drain_right.n10 drain_right.n9 0.432223
R274 drain_right.n10 drain_right.n4 0.432223
R275 plus.n14 plus.n13 161.3
R276 plus.n15 plus.n8 161.3
R277 plus.n17 plus.n16 161.3
R278 plus.n18 plus.n7 161.3
R279 plus.n19 plus.n6 161.3
R280 plus.n24 plus.n23 161.3
R281 plus.n25 plus.n4 161.3
R282 plus.n27 plus.n26 161.3
R283 plus.n28 plus.n3 161.3
R284 plus.n30 plus.n29 161.3
R285 plus.n33 plus.n0 161.3
R286 plus.n35 plus.n34 161.3
R287 plus.n50 plus.n49 161.3
R288 plus.n51 plus.n44 161.3
R289 plus.n53 plus.n52 161.3
R290 plus.n54 plus.n43 161.3
R291 plus.n55 plus.n42 161.3
R292 plus.n60 plus.n59 161.3
R293 plus.n61 plus.n40 161.3
R294 plus.n63 plus.n62 161.3
R295 plus.n64 plus.n39 161.3
R296 plus.n66 plus.n65 161.3
R297 plus.n69 plus.n36 161.3
R298 plus.n71 plus.n70 161.3
R299 plus.n10 plus.t21 100.665
R300 plus.n46 plus.t7 100.665
R301 plus.n12 plus.n9 80.6037
R302 plus.n21 plus.n20 80.6037
R303 plus.n22 plus.n5 80.6037
R304 plus.n31 plus.n2 80.6037
R305 plus.n32 plus.n1 80.6037
R306 plus.n48 plus.n45 80.6037
R307 plus.n57 plus.n56 80.6037
R308 plus.n58 plus.n41 80.6037
R309 plus.n67 plus.n38 80.6037
R310 plus.n68 plus.n37 80.6037
R311 plus.n34 plus.t4 79.2293
R312 plus.n32 plus.t6 79.2293
R313 plus.n31 plus.t9 79.2293
R314 plus.n3 plus.t10 79.2293
R315 plus.n25 plus.t11 79.2293
R316 plus.n5 plus.t13 79.2293
R317 plus.n20 plus.t14 79.2293
R318 plus.n18 plus.t18 79.2293
R319 plus.n8 plus.t15 79.2293
R320 plus.n12 plus.t16 79.2293
R321 plus.n11 plus.t19 79.2293
R322 plus.n70 plus.t17 79.2293
R323 plus.n68 plus.t5 79.2293
R324 plus.n67 plus.t0 79.2293
R325 plus.n39 plus.t3 79.2293
R326 plus.n61 plus.t12 79.2293
R327 plus.n41 plus.t2 79.2293
R328 plus.n56 plus.t23 79.2293
R329 plus.n54 plus.t1 79.2293
R330 plus.n44 plus.t22 79.2293
R331 plus.n48 plus.t8 79.2293
R332 plus.n47 plus.t20 79.2293
R333 plus.n32 plus.n31 48.2005
R334 plus.n20 plus.n5 48.2005
R335 plus.n12 plus.n11 48.2005
R336 plus.n68 plus.n67 48.2005
R337 plus.n56 plus.n41 48.2005
R338 plus.n48 plus.n47 48.2005
R339 plus.n31 plus.n30 44.549
R340 plus.n13 plus.n12 44.549
R341 plus.n67 plus.n66 44.549
R342 plus.n49 plus.n48 44.549
R343 plus.n24 plus.n5 41.6278
R344 plus.n20 plus.n19 41.6278
R345 plus.n60 plus.n41 41.6278
R346 plus.n56 plus.n55 41.6278
R347 plus.n33 plus.n32 38.7066
R348 plus.n69 plus.n68 38.7066
R349 plus plus.n71 32.8361
R350 plus.n10 plus.n9 31.6825
R351 plus.n46 plus.n45 31.6825
R352 plus.n26 plus.n3 25.5611
R353 plus.n17 plus.n8 25.5611
R354 plus.n62 plus.n39 25.5611
R355 plus.n53 plus.n44 25.5611
R356 plus.n26 plus.n25 22.6399
R357 plus.n18 plus.n17 22.6399
R358 plus.n62 plus.n61 22.6399
R359 plus.n54 plus.n53 22.6399
R360 plus.n11 plus.n10 17.2341
R361 plus.n47 plus.n46 17.2341
R362 plus.n34 plus.n33 9.49444
R363 plus.n70 plus.n69 9.49444
R364 plus plus.n35 8.13686
R365 plus.n25 plus.n24 6.57323
R366 plus.n19 plus.n18 6.57323
R367 plus.n61 plus.n60 6.57323
R368 plus.n55 plus.n54 6.57323
R369 plus.n30 plus.n3 3.65202
R370 plus.n13 plus.n8 3.65202
R371 plus.n66 plus.n39 3.65202
R372 plus.n49 plus.n44 3.65202
R373 plus.n22 plus.n21 0.380177
R374 plus.n2 plus.n1 0.380177
R375 plus.n38 plus.n37 0.380177
R376 plus.n58 plus.n57 0.380177
R377 plus.n14 plus.n9 0.285035
R378 plus.n21 plus.n6 0.285035
R379 plus.n23 plus.n22 0.285035
R380 plus.n29 plus.n2 0.285035
R381 plus.n1 plus.n0 0.285035
R382 plus.n37 plus.n36 0.285035
R383 plus.n65 plus.n38 0.285035
R384 plus.n59 plus.n58 0.285035
R385 plus.n57 plus.n42 0.285035
R386 plus.n50 plus.n45 0.285035
R387 plus.n15 plus.n14 0.189894
R388 plus.n16 plus.n15 0.189894
R389 plus.n16 plus.n7 0.189894
R390 plus.n7 plus.n6 0.189894
R391 plus.n23 plus.n4 0.189894
R392 plus.n27 plus.n4 0.189894
R393 plus.n28 plus.n27 0.189894
R394 plus.n29 plus.n28 0.189894
R395 plus.n35 plus.n0 0.189894
R396 plus.n71 plus.n36 0.189894
R397 plus.n65 plus.n64 0.189894
R398 plus.n64 plus.n63 0.189894
R399 plus.n63 plus.n40 0.189894
R400 plus.n59 plus.n40 0.189894
R401 plus.n43 plus.n42 0.189894
R402 plus.n52 plus.n43 0.189894
R403 plus.n52 plus.n51 0.189894
R404 plus.n51 plus.n50 0.189894
R405 drain_left.n13 drain_left.n11 241.107
R406 drain_left.n7 drain_left.n5 241.106
R407 drain_left.n2 drain_left.n0 241.106
R408 drain_left.n21 drain_left.n20 240.132
R409 drain_left.n19 drain_left.n18 240.132
R410 drain_left.n17 drain_left.n16 240.132
R411 drain_left.n15 drain_left.n14 240.132
R412 drain_left.n13 drain_left.n12 240.132
R413 drain_left.n7 drain_left.n6 240.131
R414 drain_left.n9 drain_left.n8 240.131
R415 drain_left.n4 drain_left.n3 240.131
R416 drain_left.n2 drain_left.n1 240.131
R417 drain_left drain_left.n10 28.288
R418 drain_left.n5 drain_left.t3 19.8005
R419 drain_left.n5 drain_left.t16 19.8005
R420 drain_left.n6 drain_left.t1 19.8005
R421 drain_left.n6 drain_left.t15 19.8005
R422 drain_left.n8 drain_left.t0 19.8005
R423 drain_left.n8 drain_left.t22 19.8005
R424 drain_left.n3 drain_left.t11 19.8005
R425 drain_left.n3 drain_left.t21 19.8005
R426 drain_left.n1 drain_left.t23 19.8005
R427 drain_left.n1 drain_left.t20 19.8005
R428 drain_left.n0 drain_left.t6 19.8005
R429 drain_left.n0 drain_left.t18 19.8005
R430 drain_left.n20 drain_left.t17 19.8005
R431 drain_left.n20 drain_left.t19 19.8005
R432 drain_left.n18 drain_left.t13 19.8005
R433 drain_left.n18 drain_left.t14 19.8005
R434 drain_left.n16 drain_left.t10 19.8005
R435 drain_left.n16 drain_left.t12 19.8005
R436 drain_left.n14 drain_left.t5 19.8005
R437 drain_left.n14 drain_left.t9 19.8005
R438 drain_left.n12 drain_left.t7 19.8005
R439 drain_left.n12 drain_left.t8 19.8005
R440 drain_left.n11 drain_left.t2 19.8005
R441 drain_left.n11 drain_left.t4 19.8005
R442 drain_left drain_left.n21 6.62735
R443 drain_left.n9 drain_left.n7 0.974638
R444 drain_left.n4 drain_left.n2 0.974638
R445 drain_left.n15 drain_left.n13 0.974638
R446 drain_left.n17 drain_left.n15 0.974638
R447 drain_left.n19 drain_left.n17 0.974638
R448 drain_left.n21 drain_left.n19 0.974638
R449 drain_left.n10 drain_left.n9 0.432223
R450 drain_left.n10 drain_left.n4 0.432223
C0 drain_right source 6.80487f
C1 minus plus 5.68179f
C2 drain_left source 6.80179f
C3 source plus 3.22889f
C4 drain_left drain_right 2.02893f
C5 minus source 3.21503f
C6 drain_right plus 0.536075f
C7 drain_right minus 2.07518f
C8 drain_left plus 2.44224f
C9 drain_left minus 0.182851f
C10 drain_right a_n3654_n1088# 6.46608f
C11 drain_left a_n3654_n1088# 7.00121f
C12 source a_n3654_n1088# 3.140654f
C13 minus a_n3654_n1088# 13.941257f
C14 plus a_n3654_n1088# 15.400749f
C15 drain_left.t6 a_n3654_n1088# 0.026102f
C16 drain_left.t18 a_n3654_n1088# 0.026102f
C17 drain_left.n0 a_n3654_n1088# 0.103248f
C18 drain_left.t23 a_n3654_n1088# 0.026102f
C19 drain_left.t20 a_n3654_n1088# 0.026102f
C20 drain_left.n1 a_n3654_n1088# 0.101423f
C21 drain_left.n2 a_n3654_n1088# 0.888167f
C22 drain_left.t11 a_n3654_n1088# 0.026102f
C23 drain_left.t21 a_n3654_n1088# 0.026102f
C24 drain_left.n3 a_n3654_n1088# 0.101423f
C25 drain_left.n4 a_n3654_n1088# 0.382387f
C26 drain_left.t3 a_n3654_n1088# 0.026102f
C27 drain_left.t16 a_n3654_n1088# 0.026102f
C28 drain_left.n5 a_n3654_n1088# 0.103248f
C29 drain_left.t1 a_n3654_n1088# 0.026102f
C30 drain_left.t15 a_n3654_n1088# 0.026102f
C31 drain_left.n6 a_n3654_n1088# 0.101423f
C32 drain_left.n7 a_n3654_n1088# 0.888167f
C33 drain_left.t0 a_n3654_n1088# 0.026102f
C34 drain_left.t22 a_n3654_n1088# 0.026102f
C35 drain_left.n8 a_n3654_n1088# 0.101423f
C36 drain_left.n9 a_n3654_n1088# 0.382387f
C37 drain_left.n10 a_n3654_n1088# 1.51478f
C38 drain_left.t2 a_n3654_n1088# 0.026102f
C39 drain_left.t4 a_n3654_n1088# 0.026102f
C40 drain_left.n11 a_n3654_n1088# 0.103248f
C41 drain_left.t7 a_n3654_n1088# 0.026102f
C42 drain_left.t8 a_n3654_n1088# 0.026102f
C43 drain_left.n12 a_n3654_n1088# 0.101424f
C44 drain_left.n13 a_n3654_n1088# 0.888167f
C45 drain_left.t5 a_n3654_n1088# 0.026102f
C46 drain_left.t9 a_n3654_n1088# 0.026102f
C47 drain_left.n14 a_n3654_n1088# 0.101424f
C48 drain_left.n15 a_n3654_n1088# 0.438344f
C49 drain_left.t10 a_n3654_n1088# 0.026102f
C50 drain_left.t12 a_n3654_n1088# 0.026102f
C51 drain_left.n16 a_n3654_n1088# 0.101424f
C52 drain_left.n17 a_n3654_n1088# 0.438344f
C53 drain_left.t13 a_n3654_n1088# 0.026102f
C54 drain_left.t14 a_n3654_n1088# 0.026102f
C55 drain_left.n18 a_n3654_n1088# 0.101424f
C56 drain_left.n19 a_n3654_n1088# 0.438344f
C57 drain_left.t17 a_n3654_n1088# 0.026102f
C58 drain_left.t19 a_n3654_n1088# 0.026102f
C59 drain_left.n20 a_n3654_n1088# 0.101424f
C60 drain_left.n21 a_n3654_n1088# 0.734526f
C61 plus.n0 a_n3654_n1088# 0.057124f
C62 plus.t4 a_n3654_n1088# 0.116134f
C63 plus.t6 a_n3654_n1088# 0.116134f
C64 plus.n1 a_n3654_n1088# 0.071305f
C65 plus.t9 a_n3654_n1088# 0.116134f
C66 plus.n2 a_n3654_n1088# 0.071305f
C67 plus.t10 a_n3654_n1088# 0.116134f
C68 plus.n3 a_n3654_n1088# 0.111539f
C69 plus.n4 a_n3654_n1088# 0.04281f
C70 plus.t11 a_n3654_n1088# 0.116134f
C71 plus.t13 a_n3654_n1088# 0.116134f
C72 plus.n5 a_n3654_n1088# 0.123497f
C73 plus.n6 a_n3654_n1088# 0.057124f
C74 plus.t14 a_n3654_n1088# 0.116134f
C75 plus.t18 a_n3654_n1088# 0.116134f
C76 plus.n7 a_n3654_n1088# 0.04281f
C77 plus.t15 a_n3654_n1088# 0.116134f
C78 plus.n8 a_n3654_n1088# 0.111539f
C79 plus.n9 a_n3654_n1088# 0.246055f
C80 plus.t16 a_n3654_n1088# 0.116134f
C81 plus.t19 a_n3654_n1088# 0.116134f
C82 plus.t21 a_n3654_n1088# 0.140654f
C83 plus.n10 a_n3654_n1088# 0.094697f
C84 plus.n11 a_n3654_n1088# 0.124003f
C85 plus.n12 a_n3654_n1088# 0.124025f
C86 plus.n13 a_n3654_n1088# 0.009714f
C87 plus.n14 a_n3654_n1088# 0.057124f
C88 plus.n15 a_n3654_n1088# 0.04281f
C89 plus.n16 a_n3654_n1088# 0.04281f
C90 plus.n17 a_n3654_n1088# 0.009714f
C91 plus.n18 a_n3654_n1088# 0.111539f
C92 plus.n19 a_n3654_n1088# 0.009714f
C93 plus.n20 a_n3654_n1088# 0.123497f
C94 plus.n21 a_n3654_n1088# 0.071305f
C95 plus.n22 a_n3654_n1088# 0.071305f
C96 plus.n23 a_n3654_n1088# 0.057124f
C97 plus.n24 a_n3654_n1088# 0.009714f
C98 plus.n25 a_n3654_n1088# 0.111539f
C99 plus.n26 a_n3654_n1088# 0.009714f
C100 plus.n27 a_n3654_n1088# 0.04281f
C101 plus.n28 a_n3654_n1088# 0.04281f
C102 plus.n29 a_n3654_n1088# 0.057124f
C103 plus.n30 a_n3654_n1088# 0.009714f
C104 plus.n31 a_n3654_n1088# 0.124025f
C105 plus.n32 a_n3654_n1088# 0.12297f
C106 plus.n33 a_n3654_n1088# 0.009714f
C107 plus.n34 a_n3654_n1088# 0.107976f
C108 plus.n35 a_n3654_n1088# 0.31035f
C109 plus.n36 a_n3654_n1088# 0.057124f
C110 plus.t17 a_n3654_n1088# 0.116134f
C111 plus.n37 a_n3654_n1088# 0.071305f
C112 plus.t5 a_n3654_n1088# 0.116134f
C113 plus.n38 a_n3654_n1088# 0.071305f
C114 plus.t0 a_n3654_n1088# 0.116134f
C115 plus.t3 a_n3654_n1088# 0.116134f
C116 plus.n39 a_n3654_n1088# 0.111539f
C117 plus.n40 a_n3654_n1088# 0.04281f
C118 plus.t12 a_n3654_n1088# 0.116134f
C119 plus.t2 a_n3654_n1088# 0.116134f
C120 plus.n41 a_n3654_n1088# 0.123497f
C121 plus.n42 a_n3654_n1088# 0.057124f
C122 plus.t23 a_n3654_n1088# 0.116134f
C123 plus.n43 a_n3654_n1088# 0.04281f
C124 plus.t1 a_n3654_n1088# 0.116134f
C125 plus.t22 a_n3654_n1088# 0.116134f
C126 plus.n44 a_n3654_n1088# 0.111539f
C127 plus.n45 a_n3654_n1088# 0.246055f
C128 plus.t8 a_n3654_n1088# 0.116134f
C129 plus.t7 a_n3654_n1088# 0.140654f
C130 plus.n46 a_n3654_n1088# 0.094697f
C131 plus.t20 a_n3654_n1088# 0.116134f
C132 plus.n47 a_n3654_n1088# 0.124003f
C133 plus.n48 a_n3654_n1088# 0.124025f
C134 plus.n49 a_n3654_n1088# 0.009714f
C135 plus.n50 a_n3654_n1088# 0.057124f
C136 plus.n51 a_n3654_n1088# 0.04281f
C137 plus.n52 a_n3654_n1088# 0.04281f
C138 plus.n53 a_n3654_n1088# 0.009714f
C139 plus.n54 a_n3654_n1088# 0.111539f
C140 plus.n55 a_n3654_n1088# 0.009714f
C141 plus.n56 a_n3654_n1088# 0.123497f
C142 plus.n57 a_n3654_n1088# 0.071305f
C143 plus.n58 a_n3654_n1088# 0.071305f
C144 plus.n59 a_n3654_n1088# 0.057124f
C145 plus.n60 a_n3654_n1088# 0.009714f
C146 plus.n61 a_n3654_n1088# 0.111539f
C147 plus.n62 a_n3654_n1088# 0.009714f
C148 plus.n63 a_n3654_n1088# 0.04281f
C149 plus.n64 a_n3654_n1088# 0.04281f
C150 plus.n65 a_n3654_n1088# 0.057124f
C151 plus.n66 a_n3654_n1088# 0.009714f
C152 plus.n67 a_n3654_n1088# 0.124025f
C153 plus.n68 a_n3654_n1088# 0.12297f
C154 plus.n69 a_n3654_n1088# 0.009714f
C155 plus.n70 a_n3654_n1088# 0.107976f
C156 plus.n71 a_n3654_n1088# 1.37254f
C157 drain_right.t16 a_n3654_n1088# 0.025699f
C158 drain_right.t2 a_n3654_n1088# 0.025699f
C159 drain_right.n0 a_n3654_n1088# 0.101655f
C160 drain_right.t17 a_n3654_n1088# 0.025699f
C161 drain_right.t3 a_n3654_n1088# 0.025699f
C162 drain_right.n1 a_n3654_n1088# 0.099859f
C163 drain_right.n2 a_n3654_n1088# 0.874465f
C164 drain_right.t20 a_n3654_n1088# 0.025699f
C165 drain_right.t1 a_n3654_n1088# 0.025699f
C166 drain_right.n3 a_n3654_n1088# 0.099859f
C167 drain_right.n4 a_n3654_n1088# 0.376488f
C168 drain_right.t8 a_n3654_n1088# 0.025699f
C169 drain_right.t22 a_n3654_n1088# 0.025699f
C170 drain_right.n5 a_n3654_n1088# 0.101655f
C171 drain_right.t19 a_n3654_n1088# 0.025699f
C172 drain_right.t23 a_n3654_n1088# 0.025699f
C173 drain_right.n6 a_n3654_n1088# 0.099859f
C174 drain_right.n7 a_n3654_n1088# 0.874465f
C175 drain_right.t21 a_n3654_n1088# 0.025699f
C176 drain_right.t0 a_n3654_n1088# 0.025699f
C177 drain_right.n8 a_n3654_n1088# 0.099859f
C178 drain_right.n9 a_n3654_n1088# 0.376488f
C179 drain_right.n10 a_n3654_n1088# 1.42933f
C180 drain_right.t14 a_n3654_n1088# 0.025699f
C181 drain_right.t10 a_n3654_n1088# 0.025699f
C182 drain_right.n11 a_n3654_n1088# 0.101656f
C183 drain_right.t7 a_n3654_n1088# 0.025699f
C184 drain_right.t15 a_n3654_n1088# 0.025699f
C185 drain_right.n12 a_n3654_n1088# 0.099859f
C186 drain_right.n13 a_n3654_n1088# 0.874465f
C187 drain_right.t9 a_n3654_n1088# 0.025699f
C188 drain_right.t5 a_n3654_n1088# 0.025699f
C189 drain_right.n14 a_n3654_n1088# 0.099859f
C190 drain_right.n15 a_n3654_n1088# 0.431581f
C191 drain_right.t4 a_n3654_n1088# 0.025699f
C192 drain_right.t12 a_n3654_n1088# 0.025699f
C193 drain_right.n16 a_n3654_n1088# 0.099859f
C194 drain_right.n17 a_n3654_n1088# 0.431581f
C195 drain_right.t18 a_n3654_n1088# 0.025699f
C196 drain_right.t6 a_n3654_n1088# 0.025699f
C197 drain_right.n18 a_n3654_n1088# 0.099859f
C198 drain_right.n19 a_n3654_n1088# 0.431581f
C199 drain_right.t13 a_n3654_n1088# 0.025699f
C200 drain_right.t11 a_n3654_n1088# 0.025699f
C201 drain_right.n20 a_n3654_n1088# 0.099859f
C202 drain_right.n21 a_n3654_n1088# 0.723195f
C203 source.t18 a_n3654_n1088# 0.16535f
C204 source.n0 a_n3654_n1088# 0.803153f
C205 source.t14 a_n3654_n1088# 0.029708f
C206 source.t5 a_n3654_n1088# 0.029708f
C207 source.n1 a_n3654_n1088# 0.096348f
C208 source.n2 a_n3654_n1088# 0.466898f
C209 source.t4 a_n3654_n1088# 0.029708f
C210 source.t17 a_n3654_n1088# 0.029708f
C211 source.n3 a_n3654_n1088# 0.096348f
C212 source.n4 a_n3654_n1088# 0.466898f
C213 source.t6 a_n3654_n1088# 0.029708f
C214 source.t3 a_n3654_n1088# 0.029708f
C215 source.n5 a_n3654_n1088# 0.096348f
C216 source.n6 a_n3654_n1088# 0.466898f
C217 source.t13 a_n3654_n1088# 0.029708f
C218 source.t20 a_n3654_n1088# 0.029708f
C219 source.n7 a_n3654_n1088# 0.096348f
C220 source.n8 a_n3654_n1088# 0.466898f
C221 source.t2 a_n3654_n1088# 0.029708f
C222 source.t16 a_n3654_n1088# 0.029708f
C223 source.n9 a_n3654_n1088# 0.096348f
C224 source.n10 a_n3654_n1088# 0.466898f
C225 source.t15 a_n3654_n1088# 0.16535f
C226 source.n11 a_n3654_n1088# 0.417827f
C227 source.t40 a_n3654_n1088# 0.16535f
C228 source.n12 a_n3654_n1088# 0.417827f
C229 source.t41 a_n3654_n1088# 0.029708f
C230 source.t28 a_n3654_n1088# 0.029708f
C231 source.n13 a_n3654_n1088# 0.096348f
C232 source.n14 a_n3654_n1088# 0.466898f
C233 source.t26 a_n3654_n1088# 0.029708f
C234 source.t25 a_n3654_n1088# 0.029708f
C235 source.n15 a_n3654_n1088# 0.096348f
C236 source.n16 a_n3654_n1088# 0.466898f
C237 source.t37 a_n3654_n1088# 0.029708f
C238 source.t38 a_n3654_n1088# 0.029708f
C239 source.n17 a_n3654_n1088# 0.096348f
C240 source.n18 a_n3654_n1088# 0.466898f
C241 source.t44 a_n3654_n1088# 0.029708f
C242 source.t39 a_n3654_n1088# 0.029708f
C243 source.n19 a_n3654_n1088# 0.096348f
C244 source.n20 a_n3654_n1088# 0.466898f
C245 source.t29 a_n3654_n1088# 0.029708f
C246 source.t47 a_n3654_n1088# 0.029708f
C247 source.n21 a_n3654_n1088# 0.096348f
C248 source.n22 a_n3654_n1088# 0.466898f
C249 source.t46 a_n3654_n1088# 0.16535f
C250 source.n23 a_n3654_n1088# 1.11566f
C251 source.t0 a_n3654_n1088# 0.16535f
C252 source.n24 a_n3654_n1088# 1.11566f
C253 source.t22 a_n3654_n1088# 0.029708f
C254 source.t10 a_n3654_n1088# 0.029708f
C255 source.n25 a_n3654_n1088# 0.096348f
C256 source.n26 a_n3654_n1088# 0.466898f
C257 source.t8 a_n3654_n1088# 0.029708f
C258 source.t1 a_n3654_n1088# 0.029708f
C259 source.n27 a_n3654_n1088# 0.096348f
C260 source.n28 a_n3654_n1088# 0.466898f
C261 source.t19 a_n3654_n1088# 0.029708f
C262 source.t11 a_n3654_n1088# 0.029708f
C263 source.n29 a_n3654_n1088# 0.096348f
C264 source.n30 a_n3654_n1088# 0.466898f
C265 source.t23 a_n3654_n1088# 0.029708f
C266 source.t9 a_n3654_n1088# 0.029708f
C267 source.n31 a_n3654_n1088# 0.096348f
C268 source.n32 a_n3654_n1088# 0.466898f
C269 source.t7 a_n3654_n1088# 0.029708f
C270 source.t12 a_n3654_n1088# 0.029708f
C271 source.n33 a_n3654_n1088# 0.096348f
C272 source.n34 a_n3654_n1088# 0.466898f
C273 source.t21 a_n3654_n1088# 0.16535f
C274 source.n35 a_n3654_n1088# 0.417827f
C275 source.t45 a_n3654_n1088# 0.16535f
C276 source.n36 a_n3654_n1088# 0.417827f
C277 source.t34 a_n3654_n1088# 0.029708f
C278 source.t30 a_n3654_n1088# 0.029708f
C279 source.n37 a_n3654_n1088# 0.096348f
C280 source.n38 a_n3654_n1088# 0.466898f
C281 source.t27 a_n3654_n1088# 0.029708f
C282 source.t24 a_n3654_n1088# 0.029708f
C283 source.n39 a_n3654_n1088# 0.096348f
C284 source.n40 a_n3654_n1088# 0.466898f
C285 source.t35 a_n3654_n1088# 0.029708f
C286 source.t32 a_n3654_n1088# 0.029708f
C287 source.n41 a_n3654_n1088# 0.096348f
C288 source.n42 a_n3654_n1088# 0.466898f
C289 source.t42 a_n3654_n1088# 0.029708f
C290 source.t43 a_n3654_n1088# 0.029708f
C291 source.n43 a_n3654_n1088# 0.096348f
C292 source.n44 a_n3654_n1088# 0.466898f
C293 source.t31 a_n3654_n1088# 0.029708f
C294 source.t36 a_n3654_n1088# 0.029708f
C295 source.n45 a_n3654_n1088# 0.096348f
C296 source.n46 a_n3654_n1088# 0.466898f
C297 source.t33 a_n3654_n1088# 0.16535f
C298 source.n47 a_n3654_n1088# 0.671193f
C299 source.n48 a_n3654_n1088# 0.783711f
C300 minus.n0 a_n3654_n1088# 0.055185f
C301 minus.t5 a_n3654_n1088# 0.112191f
C302 minus.n1 a_n3654_n1088# 0.119815f
C303 minus.t12 a_n3654_n1088# 0.112191f
C304 minus.n2 a_n3654_n1088# 0.041356f
C305 minus.t19 a_n3654_n1088# 0.112191f
C306 minus.n3 a_n3654_n1088# 0.107753f
C307 minus.n4 a_n3654_n1088# 0.068884f
C308 minus.n5 a_n3654_n1088# 0.009385f
C309 minus.t14 a_n3654_n1088# 0.112191f
C310 minus.n6 a_n3654_n1088# 0.041356f
C311 minus.n7 a_n3654_n1088# 0.009385f
C312 minus.t16 a_n3654_n1088# 0.112191f
C313 minus.t13 a_n3654_n1088# 0.135879f
C314 minus.n8 a_n3654_n1088# 0.091482f
C315 minus.t9 a_n3654_n1088# 0.112191f
C316 minus.n9 a_n3654_n1088# 0.119793f
C317 minus.t8 a_n3654_n1088# 0.112191f
C318 minus.n10 a_n3654_n1088# 0.119815f
C319 minus.n11 a_n3654_n1088# 0.237701f
C320 minus.n12 a_n3654_n1088# 0.055185f
C321 minus.n13 a_n3654_n1088# 0.041356f
C322 minus.n14 a_n3654_n1088# 0.107753f
C323 minus.n15 a_n3654_n1088# 0.009385f
C324 minus.t18 a_n3654_n1088# 0.112191f
C325 minus.n16 a_n3654_n1088# 0.107753f
C326 minus.n17 a_n3654_n1088# 0.041356f
C327 minus.n18 a_n3654_n1088# 0.055185f
C328 minus.n19 a_n3654_n1088# 0.068884f
C329 minus.n20 a_n3654_n1088# 0.119305f
C330 minus.t11 a_n3654_n1088# 0.112191f
C331 minus.n21 a_n3654_n1088# 0.119305f
C332 minus.n22 a_n3654_n1088# 0.009385f
C333 minus.n23 a_n3654_n1088# 0.055185f
C334 minus.n24 a_n3654_n1088# 0.041356f
C335 minus.n25 a_n3654_n1088# 0.041356f
C336 minus.n26 a_n3654_n1088# 0.009385f
C337 minus.t17 a_n3654_n1088# 0.112191f
C338 minus.n27 a_n3654_n1088# 0.107753f
C339 minus.n28 a_n3654_n1088# 0.009385f
C340 minus.n29 a_n3654_n1088# 0.055185f
C341 minus.n30 a_n3654_n1088# 0.068884f
C342 minus.n31 a_n3654_n1088# 0.068884f
C343 minus.n32 a_n3654_n1088# 0.118795f
C344 minus.n33 a_n3654_n1088# 0.009385f
C345 minus.t10 a_n3654_n1088# 0.112191f
C346 minus.n34 a_n3654_n1088# 0.104311f
C347 minus.n35 a_n3654_n1088# 1.37838f
C348 minus.n36 a_n3654_n1088# 0.055185f
C349 minus.t0 a_n3654_n1088# 0.112191f
C350 minus.n37 a_n3654_n1088# 0.119815f
C351 minus.n38 a_n3654_n1088# 0.041356f
C352 minus.t23 a_n3654_n1088# 0.112191f
C353 minus.n39 a_n3654_n1088# 0.107753f
C354 minus.n40 a_n3654_n1088# 0.068884f
C355 minus.n41 a_n3654_n1088# 0.009385f
C356 minus.n42 a_n3654_n1088# 0.041356f
C357 minus.n43 a_n3654_n1088# 0.009385f
C358 minus.t7 a_n3654_n1088# 0.135879f
C359 minus.n44 a_n3654_n1088# 0.091482f
C360 minus.t21 a_n3654_n1088# 0.112191f
C361 minus.n45 a_n3654_n1088# 0.119793f
C362 minus.t6 a_n3654_n1088# 0.112191f
C363 minus.n46 a_n3654_n1088# 0.119815f
C364 minus.n47 a_n3654_n1088# 0.237701f
C365 minus.n48 a_n3654_n1088# 0.055185f
C366 minus.n49 a_n3654_n1088# 0.041356f
C367 minus.t20 a_n3654_n1088# 0.112191f
C368 minus.n50 a_n3654_n1088# 0.107753f
C369 minus.n51 a_n3654_n1088# 0.009385f
C370 minus.t3 a_n3654_n1088# 0.112191f
C371 minus.n52 a_n3654_n1088# 0.107753f
C372 minus.n53 a_n3654_n1088# 0.041356f
C373 minus.n54 a_n3654_n1088# 0.055185f
C374 minus.n55 a_n3654_n1088# 0.068884f
C375 minus.t22 a_n3654_n1088# 0.112191f
C376 minus.n56 a_n3654_n1088# 0.119305f
C377 minus.t2 a_n3654_n1088# 0.112191f
C378 minus.n57 a_n3654_n1088# 0.119305f
C379 minus.n58 a_n3654_n1088# 0.009385f
C380 minus.n59 a_n3654_n1088# 0.055185f
C381 minus.n60 a_n3654_n1088# 0.041356f
C382 minus.n61 a_n3654_n1088# 0.041356f
C383 minus.n62 a_n3654_n1088# 0.009385f
C384 minus.t4 a_n3654_n1088# 0.112191f
C385 minus.n63 a_n3654_n1088# 0.107753f
C386 minus.n64 a_n3654_n1088# 0.009385f
C387 minus.n65 a_n3654_n1088# 0.055185f
C388 minus.n66 a_n3654_n1088# 0.068884f
C389 minus.n67 a_n3654_n1088# 0.068884f
C390 minus.t15 a_n3654_n1088# 0.112191f
C391 minus.n68 a_n3654_n1088# 0.118795f
C392 minus.n69 a_n3654_n1088# 0.009385f
C393 minus.t1 a_n3654_n1088# 0.112191f
C394 minus.n70 a_n3654_n1088# 0.104311f
C395 minus.n71 a_n3654_n1088# 0.285811f
C396 minus.n72 a_n3654_n1088# 1.67544f
.ends

