* NGSPICE file created from diffpair421.ext - technology: sky130A

.subckt diffpair421 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t7 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X1 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X2 source.t0 plus.t0 drain_left.t3 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X3 drain_left.t2 plus.t1 source.t1 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X4 source.t4 minus.t1 drain_right.t2 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X5 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X6 drain_left.t1 plus.t2 source.t3 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X7 source.t5 minus.t2 drain_right.t1 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X8 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X9 drain_right.t0 minus.t3 source.t6 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X10 source.t2 plus.t3 drain_left.t0 a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X11 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
R0 minus.n0 minus.t2 1324.48
R1 minus.n0 minus.t0 1324.48
R2 minus.n1 minus.t3 1324.48
R3 minus.n1 minus.t1 1324.48
R4 minus.n2 minus.n0 194.436
R5 minus.n2 minus.n1 167.77
R6 minus minus.n2 0.188
R7 source.n522 source.n462 289.615
R8 source.n456 source.n396 289.615
R9 source.n390 source.n330 289.615
R10 source.n324 source.n264 289.615
R11 source.n60 source.n0 289.615
R12 source.n126 source.n66 289.615
R13 source.n192 source.n132 289.615
R14 source.n258 source.n198 289.615
R15 source.n482 source.n481 185
R16 source.n487 source.n486 185
R17 source.n489 source.n488 185
R18 source.n478 source.n477 185
R19 source.n495 source.n494 185
R20 source.n497 source.n496 185
R21 source.n474 source.n473 185
R22 source.n504 source.n503 185
R23 source.n505 source.n472 185
R24 source.n507 source.n506 185
R25 source.n470 source.n469 185
R26 source.n513 source.n512 185
R27 source.n515 source.n514 185
R28 source.n466 source.n465 185
R29 source.n521 source.n520 185
R30 source.n523 source.n522 185
R31 source.n416 source.n415 185
R32 source.n421 source.n420 185
R33 source.n423 source.n422 185
R34 source.n412 source.n411 185
R35 source.n429 source.n428 185
R36 source.n431 source.n430 185
R37 source.n408 source.n407 185
R38 source.n438 source.n437 185
R39 source.n439 source.n406 185
R40 source.n441 source.n440 185
R41 source.n404 source.n403 185
R42 source.n447 source.n446 185
R43 source.n449 source.n448 185
R44 source.n400 source.n399 185
R45 source.n455 source.n454 185
R46 source.n457 source.n456 185
R47 source.n350 source.n349 185
R48 source.n355 source.n354 185
R49 source.n357 source.n356 185
R50 source.n346 source.n345 185
R51 source.n363 source.n362 185
R52 source.n365 source.n364 185
R53 source.n342 source.n341 185
R54 source.n372 source.n371 185
R55 source.n373 source.n340 185
R56 source.n375 source.n374 185
R57 source.n338 source.n337 185
R58 source.n381 source.n380 185
R59 source.n383 source.n382 185
R60 source.n334 source.n333 185
R61 source.n389 source.n388 185
R62 source.n391 source.n390 185
R63 source.n284 source.n283 185
R64 source.n289 source.n288 185
R65 source.n291 source.n290 185
R66 source.n280 source.n279 185
R67 source.n297 source.n296 185
R68 source.n299 source.n298 185
R69 source.n276 source.n275 185
R70 source.n306 source.n305 185
R71 source.n307 source.n274 185
R72 source.n309 source.n308 185
R73 source.n272 source.n271 185
R74 source.n315 source.n314 185
R75 source.n317 source.n316 185
R76 source.n268 source.n267 185
R77 source.n323 source.n322 185
R78 source.n325 source.n324 185
R79 source.n61 source.n60 185
R80 source.n59 source.n58 185
R81 source.n4 source.n3 185
R82 source.n53 source.n52 185
R83 source.n51 source.n50 185
R84 source.n8 source.n7 185
R85 source.n45 source.n44 185
R86 source.n43 source.n10 185
R87 source.n42 source.n41 185
R88 source.n13 source.n11 185
R89 source.n36 source.n35 185
R90 source.n34 source.n33 185
R91 source.n17 source.n16 185
R92 source.n28 source.n27 185
R93 source.n26 source.n25 185
R94 source.n21 source.n20 185
R95 source.n127 source.n126 185
R96 source.n125 source.n124 185
R97 source.n70 source.n69 185
R98 source.n119 source.n118 185
R99 source.n117 source.n116 185
R100 source.n74 source.n73 185
R101 source.n111 source.n110 185
R102 source.n109 source.n76 185
R103 source.n108 source.n107 185
R104 source.n79 source.n77 185
R105 source.n102 source.n101 185
R106 source.n100 source.n99 185
R107 source.n83 source.n82 185
R108 source.n94 source.n93 185
R109 source.n92 source.n91 185
R110 source.n87 source.n86 185
R111 source.n193 source.n192 185
R112 source.n191 source.n190 185
R113 source.n136 source.n135 185
R114 source.n185 source.n184 185
R115 source.n183 source.n182 185
R116 source.n140 source.n139 185
R117 source.n177 source.n176 185
R118 source.n175 source.n142 185
R119 source.n174 source.n173 185
R120 source.n145 source.n143 185
R121 source.n168 source.n167 185
R122 source.n166 source.n165 185
R123 source.n149 source.n148 185
R124 source.n160 source.n159 185
R125 source.n158 source.n157 185
R126 source.n153 source.n152 185
R127 source.n259 source.n258 185
R128 source.n257 source.n256 185
R129 source.n202 source.n201 185
R130 source.n251 source.n250 185
R131 source.n249 source.n248 185
R132 source.n206 source.n205 185
R133 source.n243 source.n242 185
R134 source.n241 source.n208 185
R135 source.n240 source.n239 185
R136 source.n211 source.n209 185
R137 source.n234 source.n233 185
R138 source.n232 source.n231 185
R139 source.n215 source.n214 185
R140 source.n226 source.n225 185
R141 source.n224 source.n223 185
R142 source.n219 source.n218 185
R143 source.n483 source.t6 149.524
R144 source.n417 source.t4 149.524
R145 source.n351 source.t1 149.524
R146 source.n285 source.t0 149.524
R147 source.n22 source.t3 149.524
R148 source.n88 source.t2 149.524
R149 source.n154 source.t7 149.524
R150 source.n220 source.t5 149.524
R151 source.n487 source.n481 104.615
R152 source.n488 source.n487 104.615
R153 source.n488 source.n477 104.615
R154 source.n495 source.n477 104.615
R155 source.n496 source.n495 104.615
R156 source.n496 source.n473 104.615
R157 source.n504 source.n473 104.615
R158 source.n505 source.n504 104.615
R159 source.n506 source.n505 104.615
R160 source.n506 source.n469 104.615
R161 source.n513 source.n469 104.615
R162 source.n514 source.n513 104.615
R163 source.n514 source.n465 104.615
R164 source.n521 source.n465 104.615
R165 source.n522 source.n521 104.615
R166 source.n421 source.n415 104.615
R167 source.n422 source.n421 104.615
R168 source.n422 source.n411 104.615
R169 source.n429 source.n411 104.615
R170 source.n430 source.n429 104.615
R171 source.n430 source.n407 104.615
R172 source.n438 source.n407 104.615
R173 source.n439 source.n438 104.615
R174 source.n440 source.n439 104.615
R175 source.n440 source.n403 104.615
R176 source.n447 source.n403 104.615
R177 source.n448 source.n447 104.615
R178 source.n448 source.n399 104.615
R179 source.n455 source.n399 104.615
R180 source.n456 source.n455 104.615
R181 source.n355 source.n349 104.615
R182 source.n356 source.n355 104.615
R183 source.n356 source.n345 104.615
R184 source.n363 source.n345 104.615
R185 source.n364 source.n363 104.615
R186 source.n364 source.n341 104.615
R187 source.n372 source.n341 104.615
R188 source.n373 source.n372 104.615
R189 source.n374 source.n373 104.615
R190 source.n374 source.n337 104.615
R191 source.n381 source.n337 104.615
R192 source.n382 source.n381 104.615
R193 source.n382 source.n333 104.615
R194 source.n389 source.n333 104.615
R195 source.n390 source.n389 104.615
R196 source.n289 source.n283 104.615
R197 source.n290 source.n289 104.615
R198 source.n290 source.n279 104.615
R199 source.n297 source.n279 104.615
R200 source.n298 source.n297 104.615
R201 source.n298 source.n275 104.615
R202 source.n306 source.n275 104.615
R203 source.n307 source.n306 104.615
R204 source.n308 source.n307 104.615
R205 source.n308 source.n271 104.615
R206 source.n315 source.n271 104.615
R207 source.n316 source.n315 104.615
R208 source.n316 source.n267 104.615
R209 source.n323 source.n267 104.615
R210 source.n324 source.n323 104.615
R211 source.n60 source.n59 104.615
R212 source.n59 source.n3 104.615
R213 source.n52 source.n3 104.615
R214 source.n52 source.n51 104.615
R215 source.n51 source.n7 104.615
R216 source.n44 source.n7 104.615
R217 source.n44 source.n43 104.615
R218 source.n43 source.n42 104.615
R219 source.n42 source.n11 104.615
R220 source.n35 source.n11 104.615
R221 source.n35 source.n34 104.615
R222 source.n34 source.n16 104.615
R223 source.n27 source.n16 104.615
R224 source.n27 source.n26 104.615
R225 source.n26 source.n20 104.615
R226 source.n126 source.n125 104.615
R227 source.n125 source.n69 104.615
R228 source.n118 source.n69 104.615
R229 source.n118 source.n117 104.615
R230 source.n117 source.n73 104.615
R231 source.n110 source.n73 104.615
R232 source.n110 source.n109 104.615
R233 source.n109 source.n108 104.615
R234 source.n108 source.n77 104.615
R235 source.n101 source.n77 104.615
R236 source.n101 source.n100 104.615
R237 source.n100 source.n82 104.615
R238 source.n93 source.n82 104.615
R239 source.n93 source.n92 104.615
R240 source.n92 source.n86 104.615
R241 source.n192 source.n191 104.615
R242 source.n191 source.n135 104.615
R243 source.n184 source.n135 104.615
R244 source.n184 source.n183 104.615
R245 source.n183 source.n139 104.615
R246 source.n176 source.n139 104.615
R247 source.n176 source.n175 104.615
R248 source.n175 source.n174 104.615
R249 source.n174 source.n143 104.615
R250 source.n167 source.n143 104.615
R251 source.n167 source.n166 104.615
R252 source.n166 source.n148 104.615
R253 source.n159 source.n148 104.615
R254 source.n159 source.n158 104.615
R255 source.n158 source.n152 104.615
R256 source.n258 source.n257 104.615
R257 source.n257 source.n201 104.615
R258 source.n250 source.n201 104.615
R259 source.n250 source.n249 104.615
R260 source.n249 source.n205 104.615
R261 source.n242 source.n205 104.615
R262 source.n242 source.n241 104.615
R263 source.n241 source.n240 104.615
R264 source.n240 source.n209 104.615
R265 source.n233 source.n209 104.615
R266 source.n233 source.n232 104.615
R267 source.n232 source.n214 104.615
R268 source.n225 source.n214 104.615
R269 source.n225 source.n224 104.615
R270 source.n224 source.n218 104.615
R271 source.t6 source.n481 52.3082
R272 source.t4 source.n415 52.3082
R273 source.t1 source.n349 52.3082
R274 source.t0 source.n283 52.3082
R275 source.t3 source.n20 52.3082
R276 source.t2 source.n86 52.3082
R277 source.t7 source.n152 52.3082
R278 source.t5 source.n218 52.3082
R279 source.n527 source.n526 29.8581
R280 source.n461 source.n460 29.8581
R281 source.n395 source.n394 29.8581
R282 source.n329 source.n328 29.8581
R283 source.n65 source.n64 29.8581
R284 source.n131 source.n130 29.8581
R285 source.n197 source.n196 29.8581
R286 source.n263 source.n262 29.8581
R287 source.n329 source.n263 21.8029
R288 source.n528 source.n65 16.2899
R289 source.n507 source.n472 13.1884
R290 source.n441 source.n406 13.1884
R291 source.n375 source.n340 13.1884
R292 source.n309 source.n274 13.1884
R293 source.n45 source.n10 13.1884
R294 source.n111 source.n76 13.1884
R295 source.n177 source.n142 13.1884
R296 source.n243 source.n208 13.1884
R297 source.n503 source.n502 12.8005
R298 source.n508 source.n470 12.8005
R299 source.n437 source.n436 12.8005
R300 source.n442 source.n404 12.8005
R301 source.n371 source.n370 12.8005
R302 source.n376 source.n338 12.8005
R303 source.n305 source.n304 12.8005
R304 source.n310 source.n272 12.8005
R305 source.n46 source.n8 12.8005
R306 source.n41 source.n12 12.8005
R307 source.n112 source.n74 12.8005
R308 source.n107 source.n78 12.8005
R309 source.n178 source.n140 12.8005
R310 source.n173 source.n144 12.8005
R311 source.n244 source.n206 12.8005
R312 source.n239 source.n210 12.8005
R313 source.n501 source.n474 12.0247
R314 source.n512 source.n511 12.0247
R315 source.n435 source.n408 12.0247
R316 source.n446 source.n445 12.0247
R317 source.n369 source.n342 12.0247
R318 source.n380 source.n379 12.0247
R319 source.n303 source.n276 12.0247
R320 source.n314 source.n313 12.0247
R321 source.n50 source.n49 12.0247
R322 source.n40 source.n13 12.0247
R323 source.n116 source.n115 12.0247
R324 source.n106 source.n79 12.0247
R325 source.n182 source.n181 12.0247
R326 source.n172 source.n145 12.0247
R327 source.n248 source.n247 12.0247
R328 source.n238 source.n211 12.0247
R329 source.n498 source.n497 11.249
R330 source.n515 source.n468 11.249
R331 source.n432 source.n431 11.249
R332 source.n449 source.n402 11.249
R333 source.n366 source.n365 11.249
R334 source.n383 source.n336 11.249
R335 source.n300 source.n299 11.249
R336 source.n317 source.n270 11.249
R337 source.n53 source.n6 11.249
R338 source.n37 source.n36 11.249
R339 source.n119 source.n72 11.249
R340 source.n103 source.n102 11.249
R341 source.n185 source.n138 11.249
R342 source.n169 source.n168 11.249
R343 source.n251 source.n204 11.249
R344 source.n235 source.n234 11.249
R345 source.n494 source.n476 10.4732
R346 source.n516 source.n466 10.4732
R347 source.n428 source.n410 10.4732
R348 source.n450 source.n400 10.4732
R349 source.n362 source.n344 10.4732
R350 source.n384 source.n334 10.4732
R351 source.n296 source.n278 10.4732
R352 source.n318 source.n268 10.4732
R353 source.n54 source.n4 10.4732
R354 source.n33 source.n15 10.4732
R355 source.n120 source.n70 10.4732
R356 source.n99 source.n81 10.4732
R357 source.n186 source.n136 10.4732
R358 source.n165 source.n147 10.4732
R359 source.n252 source.n202 10.4732
R360 source.n231 source.n213 10.4732
R361 source.n483 source.n482 10.2747
R362 source.n417 source.n416 10.2747
R363 source.n351 source.n350 10.2747
R364 source.n285 source.n284 10.2747
R365 source.n22 source.n21 10.2747
R366 source.n88 source.n87 10.2747
R367 source.n154 source.n153 10.2747
R368 source.n220 source.n219 10.2747
R369 source.n493 source.n478 9.69747
R370 source.n520 source.n519 9.69747
R371 source.n427 source.n412 9.69747
R372 source.n454 source.n453 9.69747
R373 source.n361 source.n346 9.69747
R374 source.n388 source.n387 9.69747
R375 source.n295 source.n280 9.69747
R376 source.n322 source.n321 9.69747
R377 source.n58 source.n57 9.69747
R378 source.n32 source.n17 9.69747
R379 source.n124 source.n123 9.69747
R380 source.n98 source.n83 9.69747
R381 source.n190 source.n189 9.69747
R382 source.n164 source.n149 9.69747
R383 source.n256 source.n255 9.69747
R384 source.n230 source.n215 9.69747
R385 source.n526 source.n525 9.45567
R386 source.n460 source.n459 9.45567
R387 source.n394 source.n393 9.45567
R388 source.n328 source.n327 9.45567
R389 source.n64 source.n63 9.45567
R390 source.n130 source.n129 9.45567
R391 source.n196 source.n195 9.45567
R392 source.n262 source.n261 9.45567
R393 source.n525 source.n524 9.3005
R394 source.n464 source.n463 9.3005
R395 source.n519 source.n518 9.3005
R396 source.n517 source.n516 9.3005
R397 source.n468 source.n467 9.3005
R398 source.n511 source.n510 9.3005
R399 source.n509 source.n508 9.3005
R400 source.n485 source.n484 9.3005
R401 source.n480 source.n479 9.3005
R402 source.n491 source.n490 9.3005
R403 source.n493 source.n492 9.3005
R404 source.n476 source.n475 9.3005
R405 source.n499 source.n498 9.3005
R406 source.n501 source.n500 9.3005
R407 source.n502 source.n471 9.3005
R408 source.n459 source.n458 9.3005
R409 source.n398 source.n397 9.3005
R410 source.n453 source.n452 9.3005
R411 source.n451 source.n450 9.3005
R412 source.n402 source.n401 9.3005
R413 source.n445 source.n444 9.3005
R414 source.n443 source.n442 9.3005
R415 source.n419 source.n418 9.3005
R416 source.n414 source.n413 9.3005
R417 source.n425 source.n424 9.3005
R418 source.n427 source.n426 9.3005
R419 source.n410 source.n409 9.3005
R420 source.n433 source.n432 9.3005
R421 source.n435 source.n434 9.3005
R422 source.n436 source.n405 9.3005
R423 source.n393 source.n392 9.3005
R424 source.n332 source.n331 9.3005
R425 source.n387 source.n386 9.3005
R426 source.n385 source.n384 9.3005
R427 source.n336 source.n335 9.3005
R428 source.n379 source.n378 9.3005
R429 source.n377 source.n376 9.3005
R430 source.n353 source.n352 9.3005
R431 source.n348 source.n347 9.3005
R432 source.n359 source.n358 9.3005
R433 source.n361 source.n360 9.3005
R434 source.n344 source.n343 9.3005
R435 source.n367 source.n366 9.3005
R436 source.n369 source.n368 9.3005
R437 source.n370 source.n339 9.3005
R438 source.n327 source.n326 9.3005
R439 source.n266 source.n265 9.3005
R440 source.n321 source.n320 9.3005
R441 source.n319 source.n318 9.3005
R442 source.n270 source.n269 9.3005
R443 source.n313 source.n312 9.3005
R444 source.n311 source.n310 9.3005
R445 source.n287 source.n286 9.3005
R446 source.n282 source.n281 9.3005
R447 source.n293 source.n292 9.3005
R448 source.n295 source.n294 9.3005
R449 source.n278 source.n277 9.3005
R450 source.n301 source.n300 9.3005
R451 source.n303 source.n302 9.3005
R452 source.n304 source.n273 9.3005
R453 source.n24 source.n23 9.3005
R454 source.n19 source.n18 9.3005
R455 source.n30 source.n29 9.3005
R456 source.n32 source.n31 9.3005
R457 source.n15 source.n14 9.3005
R458 source.n38 source.n37 9.3005
R459 source.n40 source.n39 9.3005
R460 source.n12 source.n9 9.3005
R461 source.n63 source.n62 9.3005
R462 source.n2 source.n1 9.3005
R463 source.n57 source.n56 9.3005
R464 source.n55 source.n54 9.3005
R465 source.n6 source.n5 9.3005
R466 source.n49 source.n48 9.3005
R467 source.n47 source.n46 9.3005
R468 source.n90 source.n89 9.3005
R469 source.n85 source.n84 9.3005
R470 source.n96 source.n95 9.3005
R471 source.n98 source.n97 9.3005
R472 source.n81 source.n80 9.3005
R473 source.n104 source.n103 9.3005
R474 source.n106 source.n105 9.3005
R475 source.n78 source.n75 9.3005
R476 source.n129 source.n128 9.3005
R477 source.n68 source.n67 9.3005
R478 source.n123 source.n122 9.3005
R479 source.n121 source.n120 9.3005
R480 source.n72 source.n71 9.3005
R481 source.n115 source.n114 9.3005
R482 source.n113 source.n112 9.3005
R483 source.n156 source.n155 9.3005
R484 source.n151 source.n150 9.3005
R485 source.n162 source.n161 9.3005
R486 source.n164 source.n163 9.3005
R487 source.n147 source.n146 9.3005
R488 source.n170 source.n169 9.3005
R489 source.n172 source.n171 9.3005
R490 source.n144 source.n141 9.3005
R491 source.n195 source.n194 9.3005
R492 source.n134 source.n133 9.3005
R493 source.n189 source.n188 9.3005
R494 source.n187 source.n186 9.3005
R495 source.n138 source.n137 9.3005
R496 source.n181 source.n180 9.3005
R497 source.n179 source.n178 9.3005
R498 source.n222 source.n221 9.3005
R499 source.n217 source.n216 9.3005
R500 source.n228 source.n227 9.3005
R501 source.n230 source.n229 9.3005
R502 source.n213 source.n212 9.3005
R503 source.n236 source.n235 9.3005
R504 source.n238 source.n237 9.3005
R505 source.n210 source.n207 9.3005
R506 source.n261 source.n260 9.3005
R507 source.n200 source.n199 9.3005
R508 source.n255 source.n254 9.3005
R509 source.n253 source.n252 9.3005
R510 source.n204 source.n203 9.3005
R511 source.n247 source.n246 9.3005
R512 source.n245 source.n244 9.3005
R513 source.n490 source.n489 8.92171
R514 source.n523 source.n464 8.92171
R515 source.n424 source.n423 8.92171
R516 source.n457 source.n398 8.92171
R517 source.n358 source.n357 8.92171
R518 source.n391 source.n332 8.92171
R519 source.n292 source.n291 8.92171
R520 source.n325 source.n266 8.92171
R521 source.n61 source.n2 8.92171
R522 source.n29 source.n28 8.92171
R523 source.n127 source.n68 8.92171
R524 source.n95 source.n94 8.92171
R525 source.n193 source.n134 8.92171
R526 source.n161 source.n160 8.92171
R527 source.n259 source.n200 8.92171
R528 source.n227 source.n226 8.92171
R529 source.n486 source.n480 8.14595
R530 source.n524 source.n462 8.14595
R531 source.n420 source.n414 8.14595
R532 source.n458 source.n396 8.14595
R533 source.n354 source.n348 8.14595
R534 source.n392 source.n330 8.14595
R535 source.n288 source.n282 8.14595
R536 source.n326 source.n264 8.14595
R537 source.n62 source.n0 8.14595
R538 source.n25 source.n19 8.14595
R539 source.n128 source.n66 8.14595
R540 source.n91 source.n85 8.14595
R541 source.n194 source.n132 8.14595
R542 source.n157 source.n151 8.14595
R543 source.n260 source.n198 8.14595
R544 source.n223 source.n217 8.14595
R545 source.n485 source.n482 7.3702
R546 source.n419 source.n416 7.3702
R547 source.n353 source.n350 7.3702
R548 source.n287 source.n284 7.3702
R549 source.n24 source.n21 7.3702
R550 source.n90 source.n87 7.3702
R551 source.n156 source.n153 7.3702
R552 source.n222 source.n219 7.3702
R553 source.n486 source.n485 5.81868
R554 source.n526 source.n462 5.81868
R555 source.n420 source.n419 5.81868
R556 source.n460 source.n396 5.81868
R557 source.n354 source.n353 5.81868
R558 source.n394 source.n330 5.81868
R559 source.n288 source.n287 5.81868
R560 source.n328 source.n264 5.81868
R561 source.n64 source.n0 5.81868
R562 source.n25 source.n24 5.81868
R563 source.n130 source.n66 5.81868
R564 source.n91 source.n90 5.81868
R565 source.n196 source.n132 5.81868
R566 source.n157 source.n156 5.81868
R567 source.n262 source.n198 5.81868
R568 source.n223 source.n222 5.81868
R569 source.n528 source.n527 5.51343
R570 source.n489 source.n480 5.04292
R571 source.n524 source.n523 5.04292
R572 source.n423 source.n414 5.04292
R573 source.n458 source.n457 5.04292
R574 source.n357 source.n348 5.04292
R575 source.n392 source.n391 5.04292
R576 source.n291 source.n282 5.04292
R577 source.n326 source.n325 5.04292
R578 source.n62 source.n61 5.04292
R579 source.n28 source.n19 5.04292
R580 source.n128 source.n127 5.04292
R581 source.n94 source.n85 5.04292
R582 source.n194 source.n193 5.04292
R583 source.n160 source.n151 5.04292
R584 source.n260 source.n259 5.04292
R585 source.n226 source.n217 5.04292
R586 source.n490 source.n478 4.26717
R587 source.n520 source.n464 4.26717
R588 source.n424 source.n412 4.26717
R589 source.n454 source.n398 4.26717
R590 source.n358 source.n346 4.26717
R591 source.n388 source.n332 4.26717
R592 source.n292 source.n280 4.26717
R593 source.n322 source.n266 4.26717
R594 source.n58 source.n2 4.26717
R595 source.n29 source.n17 4.26717
R596 source.n124 source.n68 4.26717
R597 source.n95 source.n83 4.26717
R598 source.n190 source.n134 4.26717
R599 source.n161 source.n149 4.26717
R600 source.n256 source.n200 4.26717
R601 source.n227 source.n215 4.26717
R602 source.n494 source.n493 3.49141
R603 source.n519 source.n466 3.49141
R604 source.n428 source.n427 3.49141
R605 source.n453 source.n400 3.49141
R606 source.n362 source.n361 3.49141
R607 source.n387 source.n334 3.49141
R608 source.n296 source.n295 3.49141
R609 source.n321 source.n268 3.49141
R610 source.n57 source.n4 3.49141
R611 source.n33 source.n32 3.49141
R612 source.n123 source.n70 3.49141
R613 source.n99 source.n98 3.49141
R614 source.n189 source.n136 3.49141
R615 source.n165 source.n164 3.49141
R616 source.n255 source.n202 3.49141
R617 source.n231 source.n230 3.49141
R618 source.n484 source.n483 2.84303
R619 source.n418 source.n417 2.84303
R620 source.n352 source.n351 2.84303
R621 source.n286 source.n285 2.84303
R622 source.n23 source.n22 2.84303
R623 source.n89 source.n88 2.84303
R624 source.n155 source.n154 2.84303
R625 source.n221 source.n220 2.84303
R626 source.n497 source.n476 2.71565
R627 source.n516 source.n515 2.71565
R628 source.n431 source.n410 2.71565
R629 source.n450 source.n449 2.71565
R630 source.n365 source.n344 2.71565
R631 source.n384 source.n383 2.71565
R632 source.n299 source.n278 2.71565
R633 source.n318 source.n317 2.71565
R634 source.n54 source.n53 2.71565
R635 source.n36 source.n15 2.71565
R636 source.n120 source.n119 2.71565
R637 source.n102 source.n81 2.71565
R638 source.n186 source.n185 2.71565
R639 source.n168 source.n147 2.71565
R640 source.n252 source.n251 2.71565
R641 source.n234 source.n213 2.71565
R642 source.n498 source.n474 1.93989
R643 source.n512 source.n468 1.93989
R644 source.n432 source.n408 1.93989
R645 source.n446 source.n402 1.93989
R646 source.n366 source.n342 1.93989
R647 source.n380 source.n336 1.93989
R648 source.n300 source.n276 1.93989
R649 source.n314 source.n270 1.93989
R650 source.n50 source.n6 1.93989
R651 source.n37 source.n13 1.93989
R652 source.n116 source.n72 1.93989
R653 source.n103 source.n79 1.93989
R654 source.n182 source.n138 1.93989
R655 source.n169 source.n145 1.93989
R656 source.n248 source.n204 1.93989
R657 source.n235 source.n211 1.93989
R658 source.n503 source.n501 1.16414
R659 source.n511 source.n470 1.16414
R660 source.n437 source.n435 1.16414
R661 source.n445 source.n404 1.16414
R662 source.n371 source.n369 1.16414
R663 source.n379 source.n338 1.16414
R664 source.n305 source.n303 1.16414
R665 source.n313 source.n272 1.16414
R666 source.n49 source.n8 1.16414
R667 source.n41 source.n40 1.16414
R668 source.n115 source.n74 1.16414
R669 source.n107 source.n106 1.16414
R670 source.n181 source.n140 1.16414
R671 source.n173 source.n172 1.16414
R672 source.n247 source.n206 1.16414
R673 source.n239 source.n238 1.16414
R674 source.n263 source.n197 0.5005
R675 source.n131 source.n65 0.5005
R676 source.n395 source.n329 0.5005
R677 source.n527 source.n461 0.5005
R678 source.n197 source.n131 0.470328
R679 source.n461 source.n395 0.470328
R680 source.n502 source.n472 0.388379
R681 source.n508 source.n507 0.388379
R682 source.n436 source.n406 0.388379
R683 source.n442 source.n441 0.388379
R684 source.n370 source.n340 0.388379
R685 source.n376 source.n375 0.388379
R686 source.n304 source.n274 0.388379
R687 source.n310 source.n309 0.388379
R688 source.n46 source.n45 0.388379
R689 source.n12 source.n10 0.388379
R690 source.n112 source.n111 0.388379
R691 source.n78 source.n76 0.388379
R692 source.n178 source.n177 0.388379
R693 source.n144 source.n142 0.388379
R694 source.n244 source.n243 0.388379
R695 source.n210 source.n208 0.388379
R696 source source.n528 0.188
R697 source.n484 source.n479 0.155672
R698 source.n491 source.n479 0.155672
R699 source.n492 source.n491 0.155672
R700 source.n492 source.n475 0.155672
R701 source.n499 source.n475 0.155672
R702 source.n500 source.n499 0.155672
R703 source.n500 source.n471 0.155672
R704 source.n509 source.n471 0.155672
R705 source.n510 source.n509 0.155672
R706 source.n510 source.n467 0.155672
R707 source.n517 source.n467 0.155672
R708 source.n518 source.n517 0.155672
R709 source.n518 source.n463 0.155672
R710 source.n525 source.n463 0.155672
R711 source.n418 source.n413 0.155672
R712 source.n425 source.n413 0.155672
R713 source.n426 source.n425 0.155672
R714 source.n426 source.n409 0.155672
R715 source.n433 source.n409 0.155672
R716 source.n434 source.n433 0.155672
R717 source.n434 source.n405 0.155672
R718 source.n443 source.n405 0.155672
R719 source.n444 source.n443 0.155672
R720 source.n444 source.n401 0.155672
R721 source.n451 source.n401 0.155672
R722 source.n452 source.n451 0.155672
R723 source.n452 source.n397 0.155672
R724 source.n459 source.n397 0.155672
R725 source.n352 source.n347 0.155672
R726 source.n359 source.n347 0.155672
R727 source.n360 source.n359 0.155672
R728 source.n360 source.n343 0.155672
R729 source.n367 source.n343 0.155672
R730 source.n368 source.n367 0.155672
R731 source.n368 source.n339 0.155672
R732 source.n377 source.n339 0.155672
R733 source.n378 source.n377 0.155672
R734 source.n378 source.n335 0.155672
R735 source.n385 source.n335 0.155672
R736 source.n386 source.n385 0.155672
R737 source.n386 source.n331 0.155672
R738 source.n393 source.n331 0.155672
R739 source.n286 source.n281 0.155672
R740 source.n293 source.n281 0.155672
R741 source.n294 source.n293 0.155672
R742 source.n294 source.n277 0.155672
R743 source.n301 source.n277 0.155672
R744 source.n302 source.n301 0.155672
R745 source.n302 source.n273 0.155672
R746 source.n311 source.n273 0.155672
R747 source.n312 source.n311 0.155672
R748 source.n312 source.n269 0.155672
R749 source.n319 source.n269 0.155672
R750 source.n320 source.n319 0.155672
R751 source.n320 source.n265 0.155672
R752 source.n327 source.n265 0.155672
R753 source.n63 source.n1 0.155672
R754 source.n56 source.n1 0.155672
R755 source.n56 source.n55 0.155672
R756 source.n55 source.n5 0.155672
R757 source.n48 source.n5 0.155672
R758 source.n48 source.n47 0.155672
R759 source.n47 source.n9 0.155672
R760 source.n39 source.n9 0.155672
R761 source.n39 source.n38 0.155672
R762 source.n38 source.n14 0.155672
R763 source.n31 source.n14 0.155672
R764 source.n31 source.n30 0.155672
R765 source.n30 source.n18 0.155672
R766 source.n23 source.n18 0.155672
R767 source.n129 source.n67 0.155672
R768 source.n122 source.n67 0.155672
R769 source.n122 source.n121 0.155672
R770 source.n121 source.n71 0.155672
R771 source.n114 source.n71 0.155672
R772 source.n114 source.n113 0.155672
R773 source.n113 source.n75 0.155672
R774 source.n105 source.n75 0.155672
R775 source.n105 source.n104 0.155672
R776 source.n104 source.n80 0.155672
R777 source.n97 source.n80 0.155672
R778 source.n97 source.n96 0.155672
R779 source.n96 source.n84 0.155672
R780 source.n89 source.n84 0.155672
R781 source.n195 source.n133 0.155672
R782 source.n188 source.n133 0.155672
R783 source.n188 source.n187 0.155672
R784 source.n187 source.n137 0.155672
R785 source.n180 source.n137 0.155672
R786 source.n180 source.n179 0.155672
R787 source.n179 source.n141 0.155672
R788 source.n171 source.n141 0.155672
R789 source.n171 source.n170 0.155672
R790 source.n170 source.n146 0.155672
R791 source.n163 source.n146 0.155672
R792 source.n163 source.n162 0.155672
R793 source.n162 source.n150 0.155672
R794 source.n155 source.n150 0.155672
R795 source.n261 source.n199 0.155672
R796 source.n254 source.n199 0.155672
R797 source.n254 source.n253 0.155672
R798 source.n253 source.n203 0.155672
R799 source.n246 source.n203 0.155672
R800 source.n246 source.n245 0.155672
R801 source.n245 source.n207 0.155672
R802 source.n237 source.n207 0.155672
R803 source.n237 source.n236 0.155672
R804 source.n236 source.n212 0.155672
R805 source.n229 source.n212 0.155672
R806 source.n229 source.n228 0.155672
R807 source.n228 source.n216 0.155672
R808 source.n221 source.n216 0.155672
R809 drain_right drain_right.n0 87.381
R810 drain_right drain_right.n1 65.7052
R811 drain_right.n0 drain_right.t2 1.6505
R812 drain_right.n0 drain_right.t0 1.6505
R813 drain_right.n1 drain_right.t1 1.6505
R814 drain_right.n1 drain_right.t3 1.6505
R815 plus.n0 plus.t3 1324.48
R816 plus.n0 plus.t2 1324.48
R817 plus.n1 plus.t1 1324.48
R818 plus.n1 plus.t0 1324.48
R819 plus plus.n1 188.317
R820 plus plus.n0 173.415
R821 drain_left drain_left.n0 87.9342
R822 drain_left drain_left.n1 65.7052
R823 drain_left.n0 drain_left.t3 1.6505
R824 drain_left.n0 drain_left.t2 1.6505
R825 drain_left.n1 drain_left.t0 1.6505
R826 drain_left.n1 drain_left.t1 1.6505
C0 drain_right drain_left 0.467153f
C1 source plus 1.37602f
C2 source drain_left 10.267799f
C3 drain_right minus 1.91541f
C4 drain_left plus 2.01324f
C5 source minus 1.36198f
C6 drain_right source 10.2661f
C7 plus minus 4.47425f
C8 drain_left minus 0.171285f
C9 drain_right plus 0.251889f
C10 drain_right a_n1064_n3292# 6.32156f
C11 drain_left a_n1064_n3292# 7.240781f
C12 source a_n1064_n3292# 8.05946f
C13 minus a_n1064_n3292# 4.042283f
C14 plus a_n1064_n3292# 7.57701f
C15 drain_left.t3 a_n1064_n3292# 0.321123f
C16 drain_left.t2 a_n1064_n3292# 0.321123f
C17 drain_left.n0 a_n1064_n3292# 3.35802f
C18 drain_left.t0 a_n1064_n3292# 0.321123f
C19 drain_left.t1 a_n1064_n3292# 0.321123f
C20 drain_left.n1 a_n1064_n3292# 2.92178f
C21 plus.t3 a_n1064_n3292# 0.45667f
C22 plus.t2 a_n1064_n3292# 0.45667f
C23 plus.n0 a_n1064_n3292# 0.416384f
C24 plus.t0 a_n1064_n3292# 0.45667f
C25 plus.t1 a_n1064_n3292# 0.45667f
C26 plus.n1 a_n1064_n3292# 0.572827f
C27 drain_right.t2 a_n1064_n3292# 0.271835f
C28 drain_right.t0 a_n1064_n3292# 0.271835f
C29 drain_right.n0 a_n1064_n3292# 2.81777f
C30 drain_right.t1 a_n1064_n3292# 0.271835f
C31 drain_right.t3 a_n1064_n3292# 0.271835f
C32 drain_right.n1 a_n1064_n3292# 2.47333f
C33 source.n0 a_n1064_n3292# 0.023261f
C34 source.n1 a_n1064_n3292# 0.01756f
C35 source.n2 a_n1064_n3292# 0.009436f
C36 source.n3 a_n1064_n3292# 0.022304f
C37 source.n4 a_n1064_n3292# 0.009991f
C38 source.n5 a_n1064_n3292# 0.01756f
C39 source.n6 a_n1064_n3292# 0.009436f
C40 source.n7 a_n1064_n3292# 0.022304f
C41 source.n8 a_n1064_n3292# 0.009991f
C42 source.n9 a_n1064_n3292# 0.01756f
C43 source.n10 a_n1064_n3292# 0.009714f
C44 source.n11 a_n1064_n3292# 0.022304f
C45 source.n12 a_n1064_n3292# 0.009436f
C46 source.n13 a_n1064_n3292# 0.009991f
C47 source.n14 a_n1064_n3292# 0.01756f
C48 source.n15 a_n1064_n3292# 0.009436f
C49 source.n16 a_n1064_n3292# 0.022304f
C50 source.n17 a_n1064_n3292# 0.009991f
C51 source.n18 a_n1064_n3292# 0.01756f
C52 source.n19 a_n1064_n3292# 0.009436f
C53 source.n20 a_n1064_n3292# 0.016728f
C54 source.n21 a_n1064_n3292# 0.015767f
C55 source.t3 a_n1064_n3292# 0.03767f
C56 source.n22 a_n1064_n3292# 0.126609f
C57 source.n23 a_n1064_n3292# 0.885899f
C58 source.n24 a_n1064_n3292# 0.009436f
C59 source.n25 a_n1064_n3292# 0.009991f
C60 source.n26 a_n1064_n3292# 0.022304f
C61 source.n27 a_n1064_n3292# 0.022304f
C62 source.n28 a_n1064_n3292# 0.009991f
C63 source.n29 a_n1064_n3292# 0.009436f
C64 source.n30 a_n1064_n3292# 0.01756f
C65 source.n31 a_n1064_n3292# 0.01756f
C66 source.n32 a_n1064_n3292# 0.009436f
C67 source.n33 a_n1064_n3292# 0.009991f
C68 source.n34 a_n1064_n3292# 0.022304f
C69 source.n35 a_n1064_n3292# 0.022304f
C70 source.n36 a_n1064_n3292# 0.009991f
C71 source.n37 a_n1064_n3292# 0.009436f
C72 source.n38 a_n1064_n3292# 0.01756f
C73 source.n39 a_n1064_n3292# 0.01756f
C74 source.n40 a_n1064_n3292# 0.009436f
C75 source.n41 a_n1064_n3292# 0.009991f
C76 source.n42 a_n1064_n3292# 0.022304f
C77 source.n43 a_n1064_n3292# 0.022304f
C78 source.n44 a_n1064_n3292# 0.022304f
C79 source.n45 a_n1064_n3292# 0.009714f
C80 source.n46 a_n1064_n3292# 0.009436f
C81 source.n47 a_n1064_n3292# 0.01756f
C82 source.n48 a_n1064_n3292# 0.01756f
C83 source.n49 a_n1064_n3292# 0.009436f
C84 source.n50 a_n1064_n3292# 0.009991f
C85 source.n51 a_n1064_n3292# 0.022304f
C86 source.n52 a_n1064_n3292# 0.022304f
C87 source.n53 a_n1064_n3292# 0.009991f
C88 source.n54 a_n1064_n3292# 0.009436f
C89 source.n55 a_n1064_n3292# 0.01756f
C90 source.n56 a_n1064_n3292# 0.01756f
C91 source.n57 a_n1064_n3292# 0.009436f
C92 source.n58 a_n1064_n3292# 0.009991f
C93 source.n59 a_n1064_n3292# 0.022304f
C94 source.n60 a_n1064_n3292# 0.04577f
C95 source.n61 a_n1064_n3292# 0.009991f
C96 source.n62 a_n1064_n3292# 0.009436f
C97 source.n63 a_n1064_n3292# 0.037712f
C98 source.n64 a_n1064_n3292# 0.02526f
C99 source.n65 a_n1064_n3292# 0.703712f
C100 source.n66 a_n1064_n3292# 0.023261f
C101 source.n67 a_n1064_n3292# 0.01756f
C102 source.n68 a_n1064_n3292# 0.009436f
C103 source.n69 a_n1064_n3292# 0.022304f
C104 source.n70 a_n1064_n3292# 0.009991f
C105 source.n71 a_n1064_n3292# 0.01756f
C106 source.n72 a_n1064_n3292# 0.009436f
C107 source.n73 a_n1064_n3292# 0.022304f
C108 source.n74 a_n1064_n3292# 0.009991f
C109 source.n75 a_n1064_n3292# 0.01756f
C110 source.n76 a_n1064_n3292# 0.009714f
C111 source.n77 a_n1064_n3292# 0.022304f
C112 source.n78 a_n1064_n3292# 0.009436f
C113 source.n79 a_n1064_n3292# 0.009991f
C114 source.n80 a_n1064_n3292# 0.01756f
C115 source.n81 a_n1064_n3292# 0.009436f
C116 source.n82 a_n1064_n3292# 0.022304f
C117 source.n83 a_n1064_n3292# 0.009991f
C118 source.n84 a_n1064_n3292# 0.01756f
C119 source.n85 a_n1064_n3292# 0.009436f
C120 source.n86 a_n1064_n3292# 0.016728f
C121 source.n87 a_n1064_n3292# 0.015767f
C122 source.t2 a_n1064_n3292# 0.03767f
C123 source.n88 a_n1064_n3292# 0.126609f
C124 source.n89 a_n1064_n3292# 0.885899f
C125 source.n90 a_n1064_n3292# 0.009436f
C126 source.n91 a_n1064_n3292# 0.009991f
C127 source.n92 a_n1064_n3292# 0.022304f
C128 source.n93 a_n1064_n3292# 0.022304f
C129 source.n94 a_n1064_n3292# 0.009991f
C130 source.n95 a_n1064_n3292# 0.009436f
C131 source.n96 a_n1064_n3292# 0.01756f
C132 source.n97 a_n1064_n3292# 0.01756f
C133 source.n98 a_n1064_n3292# 0.009436f
C134 source.n99 a_n1064_n3292# 0.009991f
C135 source.n100 a_n1064_n3292# 0.022304f
C136 source.n101 a_n1064_n3292# 0.022304f
C137 source.n102 a_n1064_n3292# 0.009991f
C138 source.n103 a_n1064_n3292# 0.009436f
C139 source.n104 a_n1064_n3292# 0.01756f
C140 source.n105 a_n1064_n3292# 0.01756f
C141 source.n106 a_n1064_n3292# 0.009436f
C142 source.n107 a_n1064_n3292# 0.009991f
C143 source.n108 a_n1064_n3292# 0.022304f
C144 source.n109 a_n1064_n3292# 0.022304f
C145 source.n110 a_n1064_n3292# 0.022304f
C146 source.n111 a_n1064_n3292# 0.009714f
C147 source.n112 a_n1064_n3292# 0.009436f
C148 source.n113 a_n1064_n3292# 0.01756f
C149 source.n114 a_n1064_n3292# 0.01756f
C150 source.n115 a_n1064_n3292# 0.009436f
C151 source.n116 a_n1064_n3292# 0.009991f
C152 source.n117 a_n1064_n3292# 0.022304f
C153 source.n118 a_n1064_n3292# 0.022304f
C154 source.n119 a_n1064_n3292# 0.009991f
C155 source.n120 a_n1064_n3292# 0.009436f
C156 source.n121 a_n1064_n3292# 0.01756f
C157 source.n122 a_n1064_n3292# 0.01756f
C158 source.n123 a_n1064_n3292# 0.009436f
C159 source.n124 a_n1064_n3292# 0.009991f
C160 source.n125 a_n1064_n3292# 0.022304f
C161 source.n126 a_n1064_n3292# 0.04577f
C162 source.n127 a_n1064_n3292# 0.009991f
C163 source.n128 a_n1064_n3292# 0.009436f
C164 source.n129 a_n1064_n3292# 0.037712f
C165 source.n130 a_n1064_n3292# 0.02526f
C166 source.n131 a_n1064_n3292# 0.068253f
C167 source.n132 a_n1064_n3292# 0.023261f
C168 source.n133 a_n1064_n3292# 0.01756f
C169 source.n134 a_n1064_n3292# 0.009436f
C170 source.n135 a_n1064_n3292# 0.022304f
C171 source.n136 a_n1064_n3292# 0.009991f
C172 source.n137 a_n1064_n3292# 0.01756f
C173 source.n138 a_n1064_n3292# 0.009436f
C174 source.n139 a_n1064_n3292# 0.022304f
C175 source.n140 a_n1064_n3292# 0.009991f
C176 source.n141 a_n1064_n3292# 0.01756f
C177 source.n142 a_n1064_n3292# 0.009714f
C178 source.n143 a_n1064_n3292# 0.022304f
C179 source.n144 a_n1064_n3292# 0.009436f
C180 source.n145 a_n1064_n3292# 0.009991f
C181 source.n146 a_n1064_n3292# 0.01756f
C182 source.n147 a_n1064_n3292# 0.009436f
C183 source.n148 a_n1064_n3292# 0.022304f
C184 source.n149 a_n1064_n3292# 0.009991f
C185 source.n150 a_n1064_n3292# 0.01756f
C186 source.n151 a_n1064_n3292# 0.009436f
C187 source.n152 a_n1064_n3292# 0.016728f
C188 source.n153 a_n1064_n3292# 0.015767f
C189 source.t7 a_n1064_n3292# 0.03767f
C190 source.n154 a_n1064_n3292# 0.126609f
C191 source.n155 a_n1064_n3292# 0.885899f
C192 source.n156 a_n1064_n3292# 0.009436f
C193 source.n157 a_n1064_n3292# 0.009991f
C194 source.n158 a_n1064_n3292# 0.022304f
C195 source.n159 a_n1064_n3292# 0.022304f
C196 source.n160 a_n1064_n3292# 0.009991f
C197 source.n161 a_n1064_n3292# 0.009436f
C198 source.n162 a_n1064_n3292# 0.01756f
C199 source.n163 a_n1064_n3292# 0.01756f
C200 source.n164 a_n1064_n3292# 0.009436f
C201 source.n165 a_n1064_n3292# 0.009991f
C202 source.n166 a_n1064_n3292# 0.022304f
C203 source.n167 a_n1064_n3292# 0.022304f
C204 source.n168 a_n1064_n3292# 0.009991f
C205 source.n169 a_n1064_n3292# 0.009436f
C206 source.n170 a_n1064_n3292# 0.01756f
C207 source.n171 a_n1064_n3292# 0.01756f
C208 source.n172 a_n1064_n3292# 0.009436f
C209 source.n173 a_n1064_n3292# 0.009991f
C210 source.n174 a_n1064_n3292# 0.022304f
C211 source.n175 a_n1064_n3292# 0.022304f
C212 source.n176 a_n1064_n3292# 0.022304f
C213 source.n177 a_n1064_n3292# 0.009714f
C214 source.n178 a_n1064_n3292# 0.009436f
C215 source.n179 a_n1064_n3292# 0.01756f
C216 source.n180 a_n1064_n3292# 0.01756f
C217 source.n181 a_n1064_n3292# 0.009436f
C218 source.n182 a_n1064_n3292# 0.009991f
C219 source.n183 a_n1064_n3292# 0.022304f
C220 source.n184 a_n1064_n3292# 0.022304f
C221 source.n185 a_n1064_n3292# 0.009991f
C222 source.n186 a_n1064_n3292# 0.009436f
C223 source.n187 a_n1064_n3292# 0.01756f
C224 source.n188 a_n1064_n3292# 0.01756f
C225 source.n189 a_n1064_n3292# 0.009436f
C226 source.n190 a_n1064_n3292# 0.009991f
C227 source.n191 a_n1064_n3292# 0.022304f
C228 source.n192 a_n1064_n3292# 0.04577f
C229 source.n193 a_n1064_n3292# 0.009991f
C230 source.n194 a_n1064_n3292# 0.009436f
C231 source.n195 a_n1064_n3292# 0.037712f
C232 source.n196 a_n1064_n3292# 0.02526f
C233 source.n197 a_n1064_n3292# 0.068253f
C234 source.n198 a_n1064_n3292# 0.023261f
C235 source.n199 a_n1064_n3292# 0.01756f
C236 source.n200 a_n1064_n3292# 0.009436f
C237 source.n201 a_n1064_n3292# 0.022304f
C238 source.n202 a_n1064_n3292# 0.009991f
C239 source.n203 a_n1064_n3292# 0.01756f
C240 source.n204 a_n1064_n3292# 0.009436f
C241 source.n205 a_n1064_n3292# 0.022304f
C242 source.n206 a_n1064_n3292# 0.009991f
C243 source.n207 a_n1064_n3292# 0.01756f
C244 source.n208 a_n1064_n3292# 0.009714f
C245 source.n209 a_n1064_n3292# 0.022304f
C246 source.n210 a_n1064_n3292# 0.009436f
C247 source.n211 a_n1064_n3292# 0.009991f
C248 source.n212 a_n1064_n3292# 0.01756f
C249 source.n213 a_n1064_n3292# 0.009436f
C250 source.n214 a_n1064_n3292# 0.022304f
C251 source.n215 a_n1064_n3292# 0.009991f
C252 source.n216 a_n1064_n3292# 0.01756f
C253 source.n217 a_n1064_n3292# 0.009436f
C254 source.n218 a_n1064_n3292# 0.016728f
C255 source.n219 a_n1064_n3292# 0.015767f
C256 source.t5 a_n1064_n3292# 0.03767f
C257 source.n220 a_n1064_n3292# 0.126609f
C258 source.n221 a_n1064_n3292# 0.885899f
C259 source.n222 a_n1064_n3292# 0.009436f
C260 source.n223 a_n1064_n3292# 0.009991f
C261 source.n224 a_n1064_n3292# 0.022304f
C262 source.n225 a_n1064_n3292# 0.022304f
C263 source.n226 a_n1064_n3292# 0.009991f
C264 source.n227 a_n1064_n3292# 0.009436f
C265 source.n228 a_n1064_n3292# 0.01756f
C266 source.n229 a_n1064_n3292# 0.01756f
C267 source.n230 a_n1064_n3292# 0.009436f
C268 source.n231 a_n1064_n3292# 0.009991f
C269 source.n232 a_n1064_n3292# 0.022304f
C270 source.n233 a_n1064_n3292# 0.022304f
C271 source.n234 a_n1064_n3292# 0.009991f
C272 source.n235 a_n1064_n3292# 0.009436f
C273 source.n236 a_n1064_n3292# 0.01756f
C274 source.n237 a_n1064_n3292# 0.01756f
C275 source.n238 a_n1064_n3292# 0.009436f
C276 source.n239 a_n1064_n3292# 0.009991f
C277 source.n240 a_n1064_n3292# 0.022304f
C278 source.n241 a_n1064_n3292# 0.022304f
C279 source.n242 a_n1064_n3292# 0.022304f
C280 source.n243 a_n1064_n3292# 0.009714f
C281 source.n244 a_n1064_n3292# 0.009436f
C282 source.n245 a_n1064_n3292# 0.01756f
C283 source.n246 a_n1064_n3292# 0.01756f
C284 source.n247 a_n1064_n3292# 0.009436f
C285 source.n248 a_n1064_n3292# 0.009991f
C286 source.n249 a_n1064_n3292# 0.022304f
C287 source.n250 a_n1064_n3292# 0.022304f
C288 source.n251 a_n1064_n3292# 0.009991f
C289 source.n252 a_n1064_n3292# 0.009436f
C290 source.n253 a_n1064_n3292# 0.01756f
C291 source.n254 a_n1064_n3292# 0.01756f
C292 source.n255 a_n1064_n3292# 0.009436f
C293 source.n256 a_n1064_n3292# 0.009991f
C294 source.n257 a_n1064_n3292# 0.022304f
C295 source.n258 a_n1064_n3292# 0.04577f
C296 source.n259 a_n1064_n3292# 0.009991f
C297 source.n260 a_n1064_n3292# 0.009436f
C298 source.n261 a_n1064_n3292# 0.037712f
C299 source.n262 a_n1064_n3292# 0.02526f
C300 source.n263 a_n1064_n3292# 0.97908f
C301 source.n264 a_n1064_n3292# 0.023261f
C302 source.n265 a_n1064_n3292# 0.01756f
C303 source.n266 a_n1064_n3292# 0.009436f
C304 source.n267 a_n1064_n3292# 0.022304f
C305 source.n268 a_n1064_n3292# 0.009991f
C306 source.n269 a_n1064_n3292# 0.01756f
C307 source.n270 a_n1064_n3292# 0.009436f
C308 source.n271 a_n1064_n3292# 0.022304f
C309 source.n272 a_n1064_n3292# 0.009991f
C310 source.n273 a_n1064_n3292# 0.01756f
C311 source.n274 a_n1064_n3292# 0.009714f
C312 source.n275 a_n1064_n3292# 0.022304f
C313 source.n276 a_n1064_n3292# 0.009991f
C314 source.n277 a_n1064_n3292# 0.01756f
C315 source.n278 a_n1064_n3292# 0.009436f
C316 source.n279 a_n1064_n3292# 0.022304f
C317 source.n280 a_n1064_n3292# 0.009991f
C318 source.n281 a_n1064_n3292# 0.01756f
C319 source.n282 a_n1064_n3292# 0.009436f
C320 source.n283 a_n1064_n3292# 0.016728f
C321 source.n284 a_n1064_n3292# 0.015767f
C322 source.t0 a_n1064_n3292# 0.03767f
C323 source.n285 a_n1064_n3292# 0.126609f
C324 source.n286 a_n1064_n3292# 0.885899f
C325 source.n287 a_n1064_n3292# 0.009436f
C326 source.n288 a_n1064_n3292# 0.009991f
C327 source.n289 a_n1064_n3292# 0.022304f
C328 source.n290 a_n1064_n3292# 0.022304f
C329 source.n291 a_n1064_n3292# 0.009991f
C330 source.n292 a_n1064_n3292# 0.009436f
C331 source.n293 a_n1064_n3292# 0.01756f
C332 source.n294 a_n1064_n3292# 0.01756f
C333 source.n295 a_n1064_n3292# 0.009436f
C334 source.n296 a_n1064_n3292# 0.009991f
C335 source.n297 a_n1064_n3292# 0.022304f
C336 source.n298 a_n1064_n3292# 0.022304f
C337 source.n299 a_n1064_n3292# 0.009991f
C338 source.n300 a_n1064_n3292# 0.009436f
C339 source.n301 a_n1064_n3292# 0.01756f
C340 source.n302 a_n1064_n3292# 0.01756f
C341 source.n303 a_n1064_n3292# 0.009436f
C342 source.n304 a_n1064_n3292# 0.009436f
C343 source.n305 a_n1064_n3292# 0.009991f
C344 source.n306 a_n1064_n3292# 0.022304f
C345 source.n307 a_n1064_n3292# 0.022304f
C346 source.n308 a_n1064_n3292# 0.022304f
C347 source.n309 a_n1064_n3292# 0.009714f
C348 source.n310 a_n1064_n3292# 0.009436f
C349 source.n311 a_n1064_n3292# 0.01756f
C350 source.n312 a_n1064_n3292# 0.01756f
C351 source.n313 a_n1064_n3292# 0.009436f
C352 source.n314 a_n1064_n3292# 0.009991f
C353 source.n315 a_n1064_n3292# 0.022304f
C354 source.n316 a_n1064_n3292# 0.022304f
C355 source.n317 a_n1064_n3292# 0.009991f
C356 source.n318 a_n1064_n3292# 0.009436f
C357 source.n319 a_n1064_n3292# 0.01756f
C358 source.n320 a_n1064_n3292# 0.01756f
C359 source.n321 a_n1064_n3292# 0.009436f
C360 source.n322 a_n1064_n3292# 0.009991f
C361 source.n323 a_n1064_n3292# 0.022304f
C362 source.n324 a_n1064_n3292# 0.04577f
C363 source.n325 a_n1064_n3292# 0.009991f
C364 source.n326 a_n1064_n3292# 0.009436f
C365 source.n327 a_n1064_n3292# 0.037712f
C366 source.n328 a_n1064_n3292# 0.02526f
C367 source.n329 a_n1064_n3292# 0.97908f
C368 source.n330 a_n1064_n3292# 0.023261f
C369 source.n331 a_n1064_n3292# 0.01756f
C370 source.n332 a_n1064_n3292# 0.009436f
C371 source.n333 a_n1064_n3292# 0.022304f
C372 source.n334 a_n1064_n3292# 0.009991f
C373 source.n335 a_n1064_n3292# 0.01756f
C374 source.n336 a_n1064_n3292# 0.009436f
C375 source.n337 a_n1064_n3292# 0.022304f
C376 source.n338 a_n1064_n3292# 0.009991f
C377 source.n339 a_n1064_n3292# 0.01756f
C378 source.n340 a_n1064_n3292# 0.009714f
C379 source.n341 a_n1064_n3292# 0.022304f
C380 source.n342 a_n1064_n3292# 0.009991f
C381 source.n343 a_n1064_n3292# 0.01756f
C382 source.n344 a_n1064_n3292# 0.009436f
C383 source.n345 a_n1064_n3292# 0.022304f
C384 source.n346 a_n1064_n3292# 0.009991f
C385 source.n347 a_n1064_n3292# 0.01756f
C386 source.n348 a_n1064_n3292# 0.009436f
C387 source.n349 a_n1064_n3292# 0.016728f
C388 source.n350 a_n1064_n3292# 0.015767f
C389 source.t1 a_n1064_n3292# 0.03767f
C390 source.n351 a_n1064_n3292# 0.126609f
C391 source.n352 a_n1064_n3292# 0.885899f
C392 source.n353 a_n1064_n3292# 0.009436f
C393 source.n354 a_n1064_n3292# 0.009991f
C394 source.n355 a_n1064_n3292# 0.022304f
C395 source.n356 a_n1064_n3292# 0.022304f
C396 source.n357 a_n1064_n3292# 0.009991f
C397 source.n358 a_n1064_n3292# 0.009436f
C398 source.n359 a_n1064_n3292# 0.01756f
C399 source.n360 a_n1064_n3292# 0.01756f
C400 source.n361 a_n1064_n3292# 0.009436f
C401 source.n362 a_n1064_n3292# 0.009991f
C402 source.n363 a_n1064_n3292# 0.022304f
C403 source.n364 a_n1064_n3292# 0.022304f
C404 source.n365 a_n1064_n3292# 0.009991f
C405 source.n366 a_n1064_n3292# 0.009436f
C406 source.n367 a_n1064_n3292# 0.01756f
C407 source.n368 a_n1064_n3292# 0.01756f
C408 source.n369 a_n1064_n3292# 0.009436f
C409 source.n370 a_n1064_n3292# 0.009436f
C410 source.n371 a_n1064_n3292# 0.009991f
C411 source.n372 a_n1064_n3292# 0.022304f
C412 source.n373 a_n1064_n3292# 0.022304f
C413 source.n374 a_n1064_n3292# 0.022304f
C414 source.n375 a_n1064_n3292# 0.009714f
C415 source.n376 a_n1064_n3292# 0.009436f
C416 source.n377 a_n1064_n3292# 0.01756f
C417 source.n378 a_n1064_n3292# 0.01756f
C418 source.n379 a_n1064_n3292# 0.009436f
C419 source.n380 a_n1064_n3292# 0.009991f
C420 source.n381 a_n1064_n3292# 0.022304f
C421 source.n382 a_n1064_n3292# 0.022304f
C422 source.n383 a_n1064_n3292# 0.009991f
C423 source.n384 a_n1064_n3292# 0.009436f
C424 source.n385 a_n1064_n3292# 0.01756f
C425 source.n386 a_n1064_n3292# 0.01756f
C426 source.n387 a_n1064_n3292# 0.009436f
C427 source.n388 a_n1064_n3292# 0.009991f
C428 source.n389 a_n1064_n3292# 0.022304f
C429 source.n390 a_n1064_n3292# 0.04577f
C430 source.n391 a_n1064_n3292# 0.009991f
C431 source.n392 a_n1064_n3292# 0.009436f
C432 source.n393 a_n1064_n3292# 0.037712f
C433 source.n394 a_n1064_n3292# 0.02526f
C434 source.n395 a_n1064_n3292# 0.068253f
C435 source.n396 a_n1064_n3292# 0.023261f
C436 source.n397 a_n1064_n3292# 0.01756f
C437 source.n398 a_n1064_n3292# 0.009436f
C438 source.n399 a_n1064_n3292# 0.022304f
C439 source.n400 a_n1064_n3292# 0.009991f
C440 source.n401 a_n1064_n3292# 0.01756f
C441 source.n402 a_n1064_n3292# 0.009436f
C442 source.n403 a_n1064_n3292# 0.022304f
C443 source.n404 a_n1064_n3292# 0.009991f
C444 source.n405 a_n1064_n3292# 0.01756f
C445 source.n406 a_n1064_n3292# 0.009714f
C446 source.n407 a_n1064_n3292# 0.022304f
C447 source.n408 a_n1064_n3292# 0.009991f
C448 source.n409 a_n1064_n3292# 0.01756f
C449 source.n410 a_n1064_n3292# 0.009436f
C450 source.n411 a_n1064_n3292# 0.022304f
C451 source.n412 a_n1064_n3292# 0.009991f
C452 source.n413 a_n1064_n3292# 0.01756f
C453 source.n414 a_n1064_n3292# 0.009436f
C454 source.n415 a_n1064_n3292# 0.016728f
C455 source.n416 a_n1064_n3292# 0.015767f
C456 source.t4 a_n1064_n3292# 0.03767f
C457 source.n417 a_n1064_n3292# 0.126609f
C458 source.n418 a_n1064_n3292# 0.885899f
C459 source.n419 a_n1064_n3292# 0.009436f
C460 source.n420 a_n1064_n3292# 0.009991f
C461 source.n421 a_n1064_n3292# 0.022304f
C462 source.n422 a_n1064_n3292# 0.022304f
C463 source.n423 a_n1064_n3292# 0.009991f
C464 source.n424 a_n1064_n3292# 0.009436f
C465 source.n425 a_n1064_n3292# 0.01756f
C466 source.n426 a_n1064_n3292# 0.01756f
C467 source.n427 a_n1064_n3292# 0.009436f
C468 source.n428 a_n1064_n3292# 0.009991f
C469 source.n429 a_n1064_n3292# 0.022304f
C470 source.n430 a_n1064_n3292# 0.022304f
C471 source.n431 a_n1064_n3292# 0.009991f
C472 source.n432 a_n1064_n3292# 0.009436f
C473 source.n433 a_n1064_n3292# 0.01756f
C474 source.n434 a_n1064_n3292# 0.01756f
C475 source.n435 a_n1064_n3292# 0.009436f
C476 source.n436 a_n1064_n3292# 0.009436f
C477 source.n437 a_n1064_n3292# 0.009991f
C478 source.n438 a_n1064_n3292# 0.022304f
C479 source.n439 a_n1064_n3292# 0.022304f
C480 source.n440 a_n1064_n3292# 0.022304f
C481 source.n441 a_n1064_n3292# 0.009714f
C482 source.n442 a_n1064_n3292# 0.009436f
C483 source.n443 a_n1064_n3292# 0.01756f
C484 source.n444 a_n1064_n3292# 0.01756f
C485 source.n445 a_n1064_n3292# 0.009436f
C486 source.n446 a_n1064_n3292# 0.009991f
C487 source.n447 a_n1064_n3292# 0.022304f
C488 source.n448 a_n1064_n3292# 0.022304f
C489 source.n449 a_n1064_n3292# 0.009991f
C490 source.n450 a_n1064_n3292# 0.009436f
C491 source.n451 a_n1064_n3292# 0.01756f
C492 source.n452 a_n1064_n3292# 0.01756f
C493 source.n453 a_n1064_n3292# 0.009436f
C494 source.n454 a_n1064_n3292# 0.009991f
C495 source.n455 a_n1064_n3292# 0.022304f
C496 source.n456 a_n1064_n3292# 0.04577f
C497 source.n457 a_n1064_n3292# 0.009991f
C498 source.n458 a_n1064_n3292# 0.009436f
C499 source.n459 a_n1064_n3292# 0.037712f
C500 source.n460 a_n1064_n3292# 0.02526f
C501 source.n461 a_n1064_n3292# 0.068253f
C502 source.n462 a_n1064_n3292# 0.023261f
C503 source.n463 a_n1064_n3292# 0.01756f
C504 source.n464 a_n1064_n3292# 0.009436f
C505 source.n465 a_n1064_n3292# 0.022304f
C506 source.n466 a_n1064_n3292# 0.009991f
C507 source.n467 a_n1064_n3292# 0.01756f
C508 source.n468 a_n1064_n3292# 0.009436f
C509 source.n469 a_n1064_n3292# 0.022304f
C510 source.n470 a_n1064_n3292# 0.009991f
C511 source.n471 a_n1064_n3292# 0.01756f
C512 source.n472 a_n1064_n3292# 0.009714f
C513 source.n473 a_n1064_n3292# 0.022304f
C514 source.n474 a_n1064_n3292# 0.009991f
C515 source.n475 a_n1064_n3292# 0.01756f
C516 source.n476 a_n1064_n3292# 0.009436f
C517 source.n477 a_n1064_n3292# 0.022304f
C518 source.n478 a_n1064_n3292# 0.009991f
C519 source.n479 a_n1064_n3292# 0.01756f
C520 source.n480 a_n1064_n3292# 0.009436f
C521 source.n481 a_n1064_n3292# 0.016728f
C522 source.n482 a_n1064_n3292# 0.015767f
C523 source.t6 a_n1064_n3292# 0.03767f
C524 source.n483 a_n1064_n3292# 0.126609f
C525 source.n484 a_n1064_n3292# 0.885899f
C526 source.n485 a_n1064_n3292# 0.009436f
C527 source.n486 a_n1064_n3292# 0.009991f
C528 source.n487 a_n1064_n3292# 0.022304f
C529 source.n488 a_n1064_n3292# 0.022304f
C530 source.n489 a_n1064_n3292# 0.009991f
C531 source.n490 a_n1064_n3292# 0.009436f
C532 source.n491 a_n1064_n3292# 0.01756f
C533 source.n492 a_n1064_n3292# 0.01756f
C534 source.n493 a_n1064_n3292# 0.009436f
C535 source.n494 a_n1064_n3292# 0.009991f
C536 source.n495 a_n1064_n3292# 0.022304f
C537 source.n496 a_n1064_n3292# 0.022304f
C538 source.n497 a_n1064_n3292# 0.009991f
C539 source.n498 a_n1064_n3292# 0.009436f
C540 source.n499 a_n1064_n3292# 0.01756f
C541 source.n500 a_n1064_n3292# 0.01756f
C542 source.n501 a_n1064_n3292# 0.009436f
C543 source.n502 a_n1064_n3292# 0.009436f
C544 source.n503 a_n1064_n3292# 0.009991f
C545 source.n504 a_n1064_n3292# 0.022304f
C546 source.n505 a_n1064_n3292# 0.022304f
C547 source.n506 a_n1064_n3292# 0.022304f
C548 source.n507 a_n1064_n3292# 0.009714f
C549 source.n508 a_n1064_n3292# 0.009436f
C550 source.n509 a_n1064_n3292# 0.01756f
C551 source.n510 a_n1064_n3292# 0.01756f
C552 source.n511 a_n1064_n3292# 0.009436f
C553 source.n512 a_n1064_n3292# 0.009991f
C554 source.n513 a_n1064_n3292# 0.022304f
C555 source.n514 a_n1064_n3292# 0.022304f
C556 source.n515 a_n1064_n3292# 0.009991f
C557 source.n516 a_n1064_n3292# 0.009436f
C558 source.n517 a_n1064_n3292# 0.01756f
C559 source.n518 a_n1064_n3292# 0.01756f
C560 source.n519 a_n1064_n3292# 0.009436f
C561 source.n520 a_n1064_n3292# 0.009991f
C562 source.n521 a_n1064_n3292# 0.022304f
C563 source.n522 a_n1064_n3292# 0.04577f
C564 source.n523 a_n1064_n3292# 0.009991f
C565 source.n524 a_n1064_n3292# 0.009436f
C566 source.n525 a_n1064_n3292# 0.037712f
C567 source.n526 a_n1064_n3292# 0.02526f
C568 source.n527 a_n1064_n3292# 0.16543f
C569 source.n528 a_n1064_n3292# 1.10151f
C570 minus.t2 a_n1064_n3292# 0.311011f
C571 minus.t0 a_n1064_n3292# 0.311011f
C572 minus.n0 a_n1064_n3292# 0.445498f
C573 minus.t1 a_n1064_n3292# 0.311011f
C574 minus.t3 a_n1064_n3292# 0.311011f
C575 minus.n1 a_n1064_n3292# 0.264251f
C576 minus.n2 a_n1064_n3292# 2.52242f
.ends

