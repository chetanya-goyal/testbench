* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t19 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X1 a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X2 a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X3 drain_right.t13 minus.t0 source.t6 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X4 drain_right.t12 minus.t1 source.t8 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X5 drain_right.t11 minus.t2 source.t4 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X6 source.t9 minus.t3 drain_right.t10 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X7 source.t24 plus.t1 drain_left.t12 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X8 drain_left.t11 plus.t2 source.t20 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X9 source.t25 plus.t3 drain_left.t10 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X10 drain_right.t9 minus.t4 source.t10 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X11 drain_left.t9 plus.t4 source.t23 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X12 source.t2 minus.t5 drain_right.t8 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X13 source.t0 minus.t6 drain_right.t7 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X14 drain_right.t6 minus.t7 source.t1 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X15 drain_left.t8 plus.t5 source.t14 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X16 a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X17 source.t15 plus.t6 drain_left.t7 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X18 drain_left.t6 plus.t7 source.t22 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X19 source.t3 minus.t8 drain_right.t5 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X20 source.t18 plus.t8 drain_left.t5 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X21 source.t26 plus.t9 drain_left.t4 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X22 drain_right.t4 minus.t9 source.t11 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X23 drain_right.t3 minus.t10 source.t7 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X24 drain_left.t3 plus.t10 source.t16 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X25 a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X26 drain_left.t2 plus.t11 source.t27 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X27 source.t17 plus.t12 drain_left.t1 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X28 source.t12 minus.t11 drain_right.t2 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X29 source.t13 minus.t12 drain_right.t1 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X30 drain_left.t0 plus.t13 source.t21 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X31 drain_right.t0 minus.t13 source.t5 a_n1564_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n3 plus.t7 567.812
R1 plus.n14 plus.t2 567.812
R2 plus.n19 plus.t4 567.812
R3 plus.n30 plus.t5 567.812
R4 plus.n4 plus.t3 518.15
R5 plus.n6 plus.t13 518.15
R6 plus.n1 plus.t12 518.15
R7 plus.n11 plus.t11 518.15
R8 plus.n13 plus.t6 518.15
R9 plus.n20 plus.t9 518.15
R10 plus.n22 plus.t0 518.15
R11 plus.n17 plus.t8 518.15
R12 plus.n27 plus.t10 518.15
R13 plus.n29 plus.t1 518.15
R14 plus.n3 plus.n2 161.489
R15 plus.n19 plus.n18 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n10 plus.n9 161.3
R19 plus.n12 plus.n0 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n21 plus.n18 161.3
R22 plus.n24 plus.n23 161.3
R23 plus.n26 plus.n25 161.3
R24 plus.n28 plus.n16 161.3
R25 plus.n31 plus.n30 161.3
R26 plus.n5 plus.n4 45.2793
R27 plus.n13 plus.n12 45.2793
R28 plus.n29 plus.n28 45.2793
R29 plus.n21 plus.n20 45.2793
R30 plus.n7 plus.n6 40.8975
R31 plus.n11 plus.n10 40.8975
R32 plus.n27 plus.n26 40.8975
R33 plus.n23 plus.n22 40.8975
R34 plus.n7 plus.n1 36.5157
R35 plus.n10 plus.n1 36.5157
R36 plus.n26 plus.n17 36.5157
R37 plus.n23 plus.n17 36.5157
R38 plus.n6 plus.n5 32.1338
R39 plus.n12 plus.n11 32.1338
R40 plus.n28 plus.n27 32.1338
R41 plus.n22 plus.n21 32.1338
R42 plus.n4 plus.n3 27.752
R43 plus.n14 plus.n13 27.752
R44 plus.n30 plus.n29 27.752
R45 plus.n20 plus.n19 27.752
R46 plus plus.n31 25.4782
R47 plus plus.n15 8.69558
R48 plus.n8 plus.n2 0.189894
R49 plus.n9 plus.n8 0.189894
R50 plus.n9 plus.n0 0.189894
R51 plus.n15 plus.n0 0.189894
R52 plus.n31 plus.n16 0.189894
R53 plus.n25 plus.n16 0.189894
R54 plus.n25 plus.n24 0.189894
R55 plus.n24 plus.n18 0.189894
R56 source.n0 source.t20 69.6943
R57 source.n7 source.t11 69.6943
R58 source.n27 source.t4 69.6942
R59 source.n20 source.t23 69.6942
R60 source.n2 source.n1 63.0943
R61 source.n4 source.n3 63.0943
R62 source.n6 source.n5 63.0943
R63 source.n9 source.n8 63.0943
R64 source.n11 source.n10 63.0943
R65 source.n13 source.n12 63.0943
R66 source.n26 source.n25 63.0942
R67 source.n24 source.n23 63.0942
R68 source.n22 source.n21 63.0942
R69 source.n19 source.n18 63.0942
R70 source.n17 source.n16 63.0942
R71 source.n15 source.n14 63.0942
R72 source.n15 source.n13 15.3833
R73 source.n28 source.n0 9.43506
R74 source.n25 source.t1 6.6005
R75 source.n25 source.t13 6.6005
R76 source.n23 source.t5 6.6005
R77 source.n23 source.t9 6.6005
R78 source.n21 source.t10 6.6005
R79 source.n21 source.t3 6.6005
R80 source.n18 source.t19 6.6005
R81 source.n18 source.t26 6.6005
R82 source.n16 source.t16 6.6005
R83 source.n16 source.t18 6.6005
R84 source.n14 source.t14 6.6005
R85 source.n14 source.t24 6.6005
R86 source.n1 source.t27 6.6005
R87 source.n1 source.t15 6.6005
R88 source.n3 source.t21 6.6005
R89 source.n3 source.t17 6.6005
R90 source.n5 source.t22 6.6005
R91 source.n5 source.t25 6.6005
R92 source.n8 source.t6 6.6005
R93 source.n8 source.t0 6.6005
R94 source.n10 source.t7 6.6005
R95 source.n10 source.t12 6.6005
R96 source.n12 source.t8 6.6005
R97 source.n12 source.t2 6.6005
R98 source.n28 source.n27 5.49188
R99 source.n7 source.n6 0.698776
R100 source.n22 source.n20 0.698776
R101 source.n13 source.n11 0.457397
R102 source.n11 source.n9 0.457397
R103 source.n9 source.n7 0.457397
R104 source.n6 source.n4 0.457397
R105 source.n4 source.n2 0.457397
R106 source.n2 source.n0 0.457397
R107 source.n17 source.n15 0.457397
R108 source.n19 source.n17 0.457397
R109 source.n20 source.n19 0.457397
R110 source.n24 source.n22 0.457397
R111 source.n26 source.n24 0.457397
R112 source.n27 source.n26 0.457397
R113 source source.n28 0.188
R114 drain_left.n7 drain_left.t6 86.83
R115 drain_left.n1 drain_left.t8 86.8299
R116 drain_left.n4 drain_left.n2 80.2299
R117 drain_left.n11 drain_left.n10 79.7731
R118 drain_left.n9 drain_left.n8 79.7731
R119 drain_left.n7 drain_left.n6 79.7731
R120 drain_left.n4 drain_left.n3 79.773
R121 drain_left.n1 drain_left.n0 79.773
R122 drain_left drain_left.n5 23.176
R123 drain_left.n2 drain_left.t4 6.6005
R124 drain_left.n2 drain_left.t9 6.6005
R125 drain_left.n3 drain_left.t5 6.6005
R126 drain_left.n3 drain_left.t13 6.6005
R127 drain_left.n0 drain_left.t12 6.6005
R128 drain_left.n0 drain_left.t3 6.6005
R129 drain_left.n10 drain_left.t7 6.6005
R130 drain_left.n10 drain_left.t11 6.6005
R131 drain_left.n8 drain_left.t1 6.6005
R132 drain_left.n8 drain_left.t2 6.6005
R133 drain_left.n6 drain_left.t10 6.6005
R134 drain_left.n6 drain_left.t0 6.6005
R135 drain_left drain_left.n11 6.11011
R136 drain_left.n9 drain_left.n7 0.457397
R137 drain_left.n11 drain_left.n9 0.457397
R138 drain_left.n5 drain_left.n1 0.287826
R139 drain_left.n5 drain_left.n4 0.0593781
R140 minus.n14 minus.t1 567.812
R141 minus.n3 minus.t9 567.812
R142 minus.n30 minus.t2 567.812
R143 minus.n19 minus.t4 567.812
R144 minus.n13 minus.t5 518.15
R145 minus.n11 minus.t10 518.15
R146 minus.n1 minus.t11 518.15
R147 minus.n6 minus.t0 518.15
R148 minus.n4 minus.t6 518.15
R149 minus.n29 minus.t12 518.15
R150 minus.n27 minus.t7 518.15
R151 minus.n17 minus.t3 518.15
R152 minus.n22 minus.t13 518.15
R153 minus.n20 minus.t8 518.15
R154 minus.n3 minus.n2 161.489
R155 minus.n19 minus.n18 161.489
R156 minus.n15 minus.n14 161.3
R157 minus.n12 minus.n0 161.3
R158 minus.n10 minus.n9 161.3
R159 minus.n8 minus.n7 161.3
R160 minus.n5 minus.n2 161.3
R161 minus.n31 minus.n30 161.3
R162 minus.n28 minus.n16 161.3
R163 minus.n26 minus.n25 161.3
R164 minus.n24 minus.n23 161.3
R165 minus.n21 minus.n18 161.3
R166 minus.n13 minus.n12 45.2793
R167 minus.n5 minus.n4 45.2793
R168 minus.n21 minus.n20 45.2793
R169 minus.n29 minus.n28 45.2793
R170 minus.n11 minus.n10 40.8975
R171 minus.n7 minus.n6 40.8975
R172 minus.n23 minus.n22 40.8975
R173 minus.n27 minus.n26 40.8975
R174 minus.n10 minus.n1 36.5157
R175 minus.n7 minus.n1 36.5157
R176 minus.n23 minus.n17 36.5157
R177 minus.n26 minus.n17 36.5157
R178 minus.n12 minus.n11 32.1338
R179 minus.n6 minus.n5 32.1338
R180 minus.n22 minus.n21 32.1338
R181 minus.n28 minus.n27 32.1338
R182 minus.n32 minus.n15 28.188
R183 minus.n14 minus.n13 27.752
R184 minus.n4 minus.n3 27.752
R185 minus.n20 minus.n19 27.752
R186 minus.n30 minus.n29 27.752
R187 minus.n32 minus.n31 6.46073
R188 minus.n15 minus.n0 0.189894
R189 minus.n9 minus.n0 0.189894
R190 minus.n9 minus.n8 0.189894
R191 minus.n8 minus.n2 0.189894
R192 minus.n24 minus.n18 0.189894
R193 minus.n25 minus.n24 0.189894
R194 minus.n25 minus.n16 0.189894
R195 minus.n31 minus.n16 0.189894
R196 minus minus.n32 0.188
R197 drain_right.n1 drain_right.t9 86.8299
R198 drain_right.n11 drain_right.t12 86.3731
R199 drain_right.n8 drain_right.n6 80.23
R200 drain_right.n4 drain_right.n2 80.2299
R201 drain_right.n8 drain_right.n7 79.7731
R202 drain_right.n10 drain_right.n9 79.7731
R203 drain_right.n4 drain_right.n3 79.773
R204 drain_right.n1 drain_right.n0 79.773
R205 drain_right drain_right.n5 22.6228
R206 drain_right.n2 drain_right.t1 6.6005
R207 drain_right.n2 drain_right.t11 6.6005
R208 drain_right.n3 drain_right.t10 6.6005
R209 drain_right.n3 drain_right.t6 6.6005
R210 drain_right.n0 drain_right.t5 6.6005
R211 drain_right.n0 drain_right.t0 6.6005
R212 drain_right.n6 drain_right.t7 6.6005
R213 drain_right.n6 drain_right.t4 6.6005
R214 drain_right.n7 drain_right.t2 6.6005
R215 drain_right.n7 drain_right.t13 6.6005
R216 drain_right.n9 drain_right.t8 6.6005
R217 drain_right.n9 drain_right.t3 6.6005
R218 drain_right drain_right.n11 5.88166
R219 drain_right.n11 drain_right.n10 0.457397
R220 drain_right.n10 drain_right.n8 0.457397
R221 drain_right.n5 drain_right.n1 0.287826
R222 drain_right.n5 drain_right.n4 0.0593781
C0 drain_right drain_left 0.791509f
C1 drain_right minus 1.33777f
C2 drain_left minus 0.176194f
C3 drain_right source 10.268901f
C4 drain_left source 10.272901f
C5 source minus 1.38222f
C6 drain_right plus 0.309995f
C7 drain_left plus 1.48703f
C8 plus minus 3.44498f
C9 plus source 1.3964f
C10 drain_right a_n1564_n1488# 4.27778f
C11 drain_left a_n1564_n1488# 4.5137f
C12 source a_n1564_n1488# 2.841442f
C13 minus a_n1564_n1488# 5.336717f
C14 plus a_n1564_n1488# 6.008798f
C15 drain_right.t9 a_n1564_n1488# 0.645365f
C16 drain_right.t5 a_n1564_n1488# 0.069532f
C17 drain_right.t0 a_n1564_n1488# 0.069532f
C18 drain_right.n0 a_n1564_n1488# 0.501454f
C19 drain_right.n1 a_n1564_n1488# 0.642972f
C20 drain_right.t1 a_n1564_n1488# 0.069532f
C21 drain_right.t11 a_n1564_n1488# 0.069532f
C22 drain_right.n2 a_n1564_n1488# 0.50335f
C23 drain_right.t10 a_n1564_n1488# 0.069532f
C24 drain_right.t6 a_n1564_n1488# 0.069532f
C25 drain_right.n3 a_n1564_n1488# 0.501454f
C26 drain_right.n4 a_n1564_n1488# 0.626128f
C27 drain_right.n5 a_n1564_n1488# 0.733257f
C28 drain_right.t7 a_n1564_n1488# 0.069532f
C29 drain_right.t4 a_n1564_n1488# 0.069532f
C30 drain_right.n6 a_n1564_n1488# 0.503352f
C31 drain_right.t2 a_n1564_n1488# 0.069532f
C32 drain_right.t13 a_n1564_n1488# 0.069532f
C33 drain_right.n7 a_n1564_n1488# 0.501456f
C34 drain_right.n8 a_n1564_n1488# 0.65219f
C35 drain_right.t8 a_n1564_n1488# 0.069532f
C36 drain_right.t3 a_n1564_n1488# 0.069532f
C37 drain_right.n9 a_n1564_n1488# 0.501456f
C38 drain_right.n10 a_n1564_n1488# 0.321136f
C39 drain_right.t12 a_n1564_n1488# 0.643592f
C40 drain_right.n11 a_n1564_n1488# 0.575649f
C41 minus.n0 a_n1564_n1488# 0.029842f
C42 minus.t1 a_n1564_n1488# 0.054817f
C43 minus.t5 a_n1564_n1488# 0.051851f
C44 minus.t10 a_n1564_n1488# 0.051851f
C45 minus.t11 a_n1564_n1488# 0.051851f
C46 minus.n1 a_n1564_n1488# 0.033174f
C47 minus.n2 a_n1564_n1488# 0.066632f
C48 minus.t0 a_n1564_n1488# 0.051851f
C49 minus.t6 a_n1564_n1488# 0.051851f
C50 minus.t9 a_n1564_n1488# 0.054817f
C51 minus.n3 a_n1564_n1488# 0.041439f
C52 minus.n4 a_n1564_n1488# 0.033174f
C53 minus.n5 a_n1564_n1488# 0.010451f
C54 minus.n6 a_n1564_n1488# 0.033174f
C55 minus.n7 a_n1564_n1488# 0.010451f
C56 minus.n8 a_n1564_n1488# 0.029842f
C57 minus.n9 a_n1564_n1488# 0.029842f
C58 minus.n10 a_n1564_n1488# 0.010451f
C59 minus.n11 a_n1564_n1488# 0.033174f
C60 minus.n12 a_n1564_n1488# 0.010451f
C61 minus.n13 a_n1564_n1488# 0.033174f
C62 minus.n14 a_n1564_n1488# 0.041395f
C63 minus.n15 a_n1564_n1488# 0.695598f
C64 minus.n16 a_n1564_n1488# 0.029842f
C65 minus.t12 a_n1564_n1488# 0.051851f
C66 minus.t7 a_n1564_n1488# 0.051851f
C67 minus.t3 a_n1564_n1488# 0.051851f
C68 minus.n17 a_n1564_n1488# 0.033174f
C69 minus.n18 a_n1564_n1488# 0.066632f
C70 minus.t13 a_n1564_n1488# 0.051851f
C71 minus.t8 a_n1564_n1488# 0.051851f
C72 minus.t4 a_n1564_n1488# 0.054817f
C73 minus.n19 a_n1564_n1488# 0.041439f
C74 minus.n20 a_n1564_n1488# 0.033174f
C75 minus.n21 a_n1564_n1488# 0.010451f
C76 minus.n22 a_n1564_n1488# 0.033174f
C77 minus.n23 a_n1564_n1488# 0.010451f
C78 minus.n24 a_n1564_n1488# 0.029842f
C79 minus.n25 a_n1564_n1488# 0.029842f
C80 minus.n26 a_n1564_n1488# 0.010451f
C81 minus.n27 a_n1564_n1488# 0.033174f
C82 minus.n28 a_n1564_n1488# 0.010451f
C83 minus.n29 a_n1564_n1488# 0.033174f
C84 minus.t2 a_n1564_n1488# 0.054817f
C85 minus.n30 a_n1564_n1488# 0.041395f
C86 minus.n31 a_n1564_n1488# 0.192332f
C87 minus.n32 a_n1564_n1488# 0.861362f
C88 drain_left.t8 a_n1564_n1488# 0.638255f
C89 drain_left.t12 a_n1564_n1488# 0.068766f
C90 drain_left.t3 a_n1564_n1488# 0.068766f
C91 drain_left.n0 a_n1564_n1488# 0.49593f
C92 drain_left.n1 a_n1564_n1488# 0.635889f
C93 drain_left.t4 a_n1564_n1488# 0.068766f
C94 drain_left.t9 a_n1564_n1488# 0.068766f
C95 drain_left.n2 a_n1564_n1488# 0.497805f
C96 drain_left.t5 a_n1564_n1488# 0.068766f
C97 drain_left.t13 a_n1564_n1488# 0.068766f
C98 drain_left.n3 a_n1564_n1488# 0.49593f
C99 drain_left.n4 a_n1564_n1488# 0.61923f
C100 drain_left.n5 a_n1564_n1488# 0.782851f
C101 drain_left.t6 a_n1564_n1488# 0.638258f
C102 drain_left.t10 a_n1564_n1488# 0.068766f
C103 drain_left.t0 a_n1564_n1488# 0.068766f
C104 drain_left.n6 a_n1564_n1488# 0.495932f
C105 drain_left.n7 a_n1564_n1488# 0.649393f
C106 drain_left.t1 a_n1564_n1488# 0.068766f
C107 drain_left.t2 a_n1564_n1488# 0.068766f
C108 drain_left.n8 a_n1564_n1488# 0.495932f
C109 drain_left.n9 a_n1564_n1488# 0.317598f
C110 drain_left.t7 a_n1564_n1488# 0.068766f
C111 drain_left.t11 a_n1564_n1488# 0.068766f
C112 drain_left.n10 a_n1564_n1488# 0.495932f
C113 drain_left.n11 a_n1564_n1488# 0.554989f
C114 source.t20 a_n1564_n1488# 0.663449f
C115 source.n0 a_n1564_n1488# 0.888667f
C116 source.t27 a_n1564_n1488# 0.079897f
C117 source.t15 a_n1564_n1488# 0.079897f
C118 source.n1 a_n1564_n1488# 0.506591f
C119 source.n2 a_n1564_n1488# 0.39282f
C120 source.t21 a_n1564_n1488# 0.079897f
C121 source.t17 a_n1564_n1488# 0.079897f
C122 source.n3 a_n1564_n1488# 0.506591f
C123 source.n4 a_n1564_n1488# 0.39282f
C124 source.t22 a_n1564_n1488# 0.079897f
C125 source.t25 a_n1564_n1488# 0.079897f
C126 source.n5 a_n1564_n1488# 0.506591f
C127 source.n6 a_n1564_n1488# 0.419033f
C128 source.t11 a_n1564_n1488# 0.663449f
C129 source.n7 a_n1564_n1488# 0.480076f
C130 source.t6 a_n1564_n1488# 0.079897f
C131 source.t0 a_n1564_n1488# 0.079897f
C132 source.n8 a_n1564_n1488# 0.506591f
C133 source.n9 a_n1564_n1488# 0.39282f
C134 source.t7 a_n1564_n1488# 0.079897f
C135 source.t12 a_n1564_n1488# 0.079897f
C136 source.n10 a_n1564_n1488# 0.506591f
C137 source.n11 a_n1564_n1488# 0.39282f
C138 source.t8 a_n1564_n1488# 0.079897f
C139 source.t2 a_n1564_n1488# 0.079897f
C140 source.n12 a_n1564_n1488# 0.506591f
C141 source.n13 a_n1564_n1488# 1.22631f
C142 source.t14 a_n1564_n1488# 0.079897f
C143 source.t24 a_n1564_n1488# 0.079897f
C144 source.n14 a_n1564_n1488# 0.506588f
C145 source.n15 a_n1564_n1488# 1.22632f
C146 source.t16 a_n1564_n1488# 0.079897f
C147 source.t18 a_n1564_n1488# 0.079897f
C148 source.n16 a_n1564_n1488# 0.506588f
C149 source.n17 a_n1564_n1488# 0.392824f
C150 source.t19 a_n1564_n1488# 0.079897f
C151 source.t26 a_n1564_n1488# 0.079897f
C152 source.n18 a_n1564_n1488# 0.506588f
C153 source.n19 a_n1564_n1488# 0.392824f
C154 source.t23 a_n1564_n1488# 0.663445f
C155 source.n20 a_n1564_n1488# 0.480079f
C156 source.t10 a_n1564_n1488# 0.079897f
C157 source.t3 a_n1564_n1488# 0.079897f
C158 source.n21 a_n1564_n1488# 0.506588f
C159 source.n22 a_n1564_n1488# 0.419036f
C160 source.t5 a_n1564_n1488# 0.079897f
C161 source.t9 a_n1564_n1488# 0.079897f
C162 source.n23 a_n1564_n1488# 0.506588f
C163 source.n24 a_n1564_n1488# 0.392824f
C164 source.t1 a_n1564_n1488# 0.079897f
C165 source.t13 a_n1564_n1488# 0.079897f
C166 source.n25 a_n1564_n1488# 0.506588f
C167 source.n26 a_n1564_n1488# 0.392824f
C168 source.t4 a_n1564_n1488# 0.663445f
C169 source.n27 a_n1564_n1488# 0.638013f
C170 source.n28 a_n1564_n1488# 0.972773f
C171 plus.n0 a_n1564_n1488# 0.030381f
C172 plus.t6 a_n1564_n1488# 0.052788f
C173 plus.t11 a_n1564_n1488# 0.052788f
C174 plus.t12 a_n1564_n1488# 0.052788f
C175 plus.n1 a_n1564_n1488# 0.033773f
C176 plus.n2 a_n1564_n1488# 0.067836f
C177 plus.t13 a_n1564_n1488# 0.052788f
C178 plus.t3 a_n1564_n1488# 0.052788f
C179 plus.t7 a_n1564_n1488# 0.055808f
C180 plus.n3 a_n1564_n1488# 0.042187f
C181 plus.n4 a_n1564_n1488# 0.033773f
C182 plus.n5 a_n1564_n1488# 0.01064f
C183 plus.n6 a_n1564_n1488# 0.033773f
C184 plus.n7 a_n1564_n1488# 0.01064f
C185 plus.n8 a_n1564_n1488# 0.030381f
C186 plus.n9 a_n1564_n1488# 0.030381f
C187 plus.n10 a_n1564_n1488# 0.01064f
C188 plus.n11 a_n1564_n1488# 0.033773f
C189 plus.n12 a_n1564_n1488# 0.01064f
C190 plus.n13 a_n1564_n1488# 0.033773f
C191 plus.t2 a_n1564_n1488# 0.055808f
C192 plus.n14 a_n1564_n1488# 0.042143f
C193 plus.n15 a_n1564_n1488# 0.223981f
C194 plus.n16 a_n1564_n1488# 0.030381f
C195 plus.t5 a_n1564_n1488# 0.055808f
C196 plus.t1 a_n1564_n1488# 0.052788f
C197 plus.t10 a_n1564_n1488# 0.052788f
C198 plus.t8 a_n1564_n1488# 0.052788f
C199 plus.n17 a_n1564_n1488# 0.033773f
C200 plus.n18 a_n1564_n1488# 0.067836f
C201 plus.t0 a_n1564_n1488# 0.052788f
C202 plus.t9 a_n1564_n1488# 0.052788f
C203 plus.t4 a_n1564_n1488# 0.055808f
C204 plus.n19 a_n1564_n1488# 0.042187f
C205 plus.n20 a_n1564_n1488# 0.033773f
C206 plus.n21 a_n1564_n1488# 0.01064f
C207 plus.n22 a_n1564_n1488# 0.033773f
C208 plus.n23 a_n1564_n1488# 0.01064f
C209 plus.n24 a_n1564_n1488# 0.030381f
C210 plus.n25 a_n1564_n1488# 0.030381f
C211 plus.n26 a_n1564_n1488# 0.01064f
C212 plus.n27 a_n1564_n1488# 0.033773f
C213 plus.n28 a_n1564_n1488# 0.01064f
C214 plus.n29 a_n1564_n1488# 0.033773f
C215 plus.n30 a_n1564_n1488# 0.042143f
C216 plus.n31 a_n1564_n1488# 0.667436f
.ends

