* NGSPICE file created from diffpair279.ext - technology: sky130A

.subckt diffpair279 minus drain_right drain_left source plus
X0 source.t33 plus.t0 drain_left.t1 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t46 minus.t0 drain_right.t23 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 source.t6 minus.t1 drain_right.t22 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X3 a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X4 drain_left.t0 plus.t1 source.t32 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X5 source.t2 minus.t2 drain_right.t21 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X6 drain_right.t20 minus.t3 source.t5 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 drain_right.t19 minus.t4 source.t7 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X8 source.t34 minus.t5 drain_right.t18 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X9 source.t38 minus.t6 drain_right.t17 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 drain_left.t2 plus.t2 source.t31 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X11 source.t30 plus.t3 drain_left.t3 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X12 source.t29 plus.t4 drain_left.t15 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X13 source.t28 plus.t5 drain_left.t22 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 source.t27 plus.t6 drain_left.t20 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X15 drain_left.t19 plus.t7 source.t26 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X16 a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X17 drain_right.t16 minus.t7 source.t0 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X18 drain_right.t15 minus.t8 source.t1 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X19 drain_right.t14 minus.t9 source.t39 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X20 source.t41 minus.t10 drain_right.t13 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X21 source.t44 minus.t11 drain_right.t12 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X22 a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X23 drain_right.t11 minus.t12 source.t35 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X24 source.t25 plus.t8 drain_left.t13 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X25 source.t24 plus.t9 drain_left.t14 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X26 drain_right.t10 minus.t13 source.t40 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X27 source.t23 plus.t10 drain_left.t23 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X28 drain_left.t5 plus.t11 source.t22 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X29 drain_left.t8 plus.t12 source.t21 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X30 drain_left.t11 plus.t13 source.t20 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X31 source.t9 minus.t14 drain_right.t9 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X32 source.t19 plus.t14 drain_left.t17 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X33 drain_right.t8 minus.t15 source.t43 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X34 drain_left.t6 plus.t15 source.t18 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X35 source.t47 minus.t16 drain_right.t7 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X36 source.t36 minus.t17 drain_right.t6 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X37 source.t17 plus.t16 drain_left.t9 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X38 drain_right.t5 minus.t18 source.t4 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X39 drain_right.t4 minus.t19 source.t8 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X40 source.t16 plus.t17 drain_left.t4 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X41 drain_left.t16 plus.t18 source.t15 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X42 drain_left.t12 plus.t19 source.t14 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X43 drain_right.t3 minus.t20 source.t37 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X44 drain_right.t2 minus.t21 source.t42 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X45 a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X46 drain_left.t21 plus.t20 source.t13 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X47 drain_left.t18 plus.t21 source.t12 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X48 source.t45 minus.t22 drain_right.t1 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X49 source.t3 minus.t23 drain_right.t0 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X50 source.t11 plus.t22 drain_left.t7 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X51 drain_left.t10 plus.t23 source.t10 a_n2354_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 plus.n9 plus.t4 617.837
R1 plus.n35 plus.t7 617.837
R2 plus.n46 plus.t12 617.837
R3 plus.n72 plus.t17 617.837
R4 plus.n8 plus.t11 586.433
R5 plus.n13 plus.t16 586.433
R6 plus.n15 plus.t23 586.433
R7 plus.n5 plus.t10 586.433
R8 plus.n20 plus.t15 586.433
R9 plus.n3 plus.t22 586.433
R10 plus.n26 plus.t1 586.433
R11 plus.n28 plus.t14 586.433
R12 plus.n1 plus.t19 586.433
R13 plus.n34 plus.t0 586.433
R14 plus.n45 plus.t3 586.433
R15 plus.n50 plus.t13 586.433
R16 plus.n52 plus.t5 586.433
R17 plus.n42 plus.t20 586.433
R18 plus.n57 plus.t6 586.433
R19 plus.n40 plus.t21 586.433
R20 plus.n63 plus.t8 586.433
R21 plus.n65 plus.t18 586.433
R22 plus.n38 plus.t9 586.433
R23 plus.n71 plus.t2 586.433
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 29.6164
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus.n8 plus.n7 12.4157
R88 plus.n34 plus.n33 12.4157
R89 plus.n71 plus.n70 12.4157
R90 plus.n45 plus.n44 12.4157
R91 plus plus.n36 9.84141
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 drain_left.n13 drain_left.n11 67.7339
R125 drain_left.n7 drain_left.n5 67.7338
R126 drain_left.n2 drain_left.n0 67.7338
R127 drain_left.n19 drain_left.n18 67.1908
R128 drain_left.n17 drain_left.n16 67.1908
R129 drain_left.n15 drain_left.n14 67.1908
R130 drain_left.n13 drain_left.n12 67.1908
R131 drain_left.n21 drain_left.n20 67.1907
R132 drain_left.n7 drain_left.n6 67.1907
R133 drain_left.n9 drain_left.n8 67.1907
R134 drain_left.n4 drain_left.n3 67.1907
R135 drain_left.n2 drain_left.n1 67.1907
R136 drain_left drain_left.n10 27.9811
R137 drain_left drain_left.n21 6.19632
R138 drain_left.n5 drain_left.t3 3.3005
R139 drain_left.n5 drain_left.t8 3.3005
R140 drain_left.n6 drain_left.t22 3.3005
R141 drain_left.n6 drain_left.t11 3.3005
R142 drain_left.n8 drain_left.t20 3.3005
R143 drain_left.n8 drain_left.t21 3.3005
R144 drain_left.n3 drain_left.t13 3.3005
R145 drain_left.n3 drain_left.t18 3.3005
R146 drain_left.n1 drain_left.t14 3.3005
R147 drain_left.n1 drain_left.t16 3.3005
R148 drain_left.n0 drain_left.t4 3.3005
R149 drain_left.n0 drain_left.t2 3.3005
R150 drain_left.n20 drain_left.t1 3.3005
R151 drain_left.n20 drain_left.t19 3.3005
R152 drain_left.n18 drain_left.t17 3.3005
R153 drain_left.n18 drain_left.t12 3.3005
R154 drain_left.n16 drain_left.t7 3.3005
R155 drain_left.n16 drain_left.t0 3.3005
R156 drain_left.n14 drain_left.t23 3.3005
R157 drain_left.n14 drain_left.t6 3.3005
R158 drain_left.n12 drain_left.t9 3.3005
R159 drain_left.n12 drain_left.t10 3.3005
R160 drain_left.n11 drain_left.t15 3.3005
R161 drain_left.n11 drain_left.t5 3.3005
R162 drain_left.n9 drain_left.n7 0.543603
R163 drain_left.n4 drain_left.n2 0.543603
R164 drain_left.n15 drain_left.n13 0.543603
R165 drain_left.n17 drain_left.n15 0.543603
R166 drain_left.n19 drain_left.n17 0.543603
R167 drain_left.n21 drain_left.n19 0.543603
R168 drain_left.n10 drain_left.n9 0.216706
R169 drain_left.n10 drain_left.n4 0.216706
R170 source.n290 source.n264 289.615
R171 source.n248 source.n222 289.615
R172 source.n216 source.n190 289.615
R173 source.n174 source.n148 289.615
R174 source.n26 source.n0 289.615
R175 source.n68 source.n42 289.615
R176 source.n100 source.n74 289.615
R177 source.n142 source.n116 289.615
R178 source.n275 source.n274 185
R179 source.n272 source.n271 185
R180 source.n281 source.n280 185
R181 source.n283 source.n282 185
R182 source.n268 source.n267 185
R183 source.n289 source.n288 185
R184 source.n291 source.n290 185
R185 source.n233 source.n232 185
R186 source.n230 source.n229 185
R187 source.n239 source.n238 185
R188 source.n241 source.n240 185
R189 source.n226 source.n225 185
R190 source.n247 source.n246 185
R191 source.n249 source.n248 185
R192 source.n201 source.n200 185
R193 source.n198 source.n197 185
R194 source.n207 source.n206 185
R195 source.n209 source.n208 185
R196 source.n194 source.n193 185
R197 source.n215 source.n214 185
R198 source.n217 source.n216 185
R199 source.n159 source.n158 185
R200 source.n156 source.n155 185
R201 source.n165 source.n164 185
R202 source.n167 source.n166 185
R203 source.n152 source.n151 185
R204 source.n173 source.n172 185
R205 source.n175 source.n174 185
R206 source.n27 source.n26 185
R207 source.n25 source.n24 185
R208 source.n4 source.n3 185
R209 source.n19 source.n18 185
R210 source.n17 source.n16 185
R211 source.n8 source.n7 185
R212 source.n11 source.n10 185
R213 source.n69 source.n68 185
R214 source.n67 source.n66 185
R215 source.n46 source.n45 185
R216 source.n61 source.n60 185
R217 source.n59 source.n58 185
R218 source.n50 source.n49 185
R219 source.n53 source.n52 185
R220 source.n101 source.n100 185
R221 source.n99 source.n98 185
R222 source.n78 source.n77 185
R223 source.n93 source.n92 185
R224 source.n91 source.n90 185
R225 source.n82 source.n81 185
R226 source.n85 source.n84 185
R227 source.n143 source.n142 185
R228 source.n141 source.n140 185
R229 source.n120 source.n119 185
R230 source.n135 source.n134 185
R231 source.n133 source.n132 185
R232 source.n124 source.n123 185
R233 source.n127 source.n126 185
R234 source.t4 source.n273 147.661
R235 source.t36 source.n231 147.661
R236 source.t21 source.n199 147.661
R237 source.t16 source.n157 147.661
R238 source.t26 source.n9 147.661
R239 source.t29 source.n51 147.661
R240 source.t43 source.n83 147.661
R241 source.t34 source.n125 147.661
R242 source.n274 source.n271 104.615
R243 source.n281 source.n271 104.615
R244 source.n282 source.n281 104.615
R245 source.n282 source.n267 104.615
R246 source.n289 source.n267 104.615
R247 source.n290 source.n289 104.615
R248 source.n232 source.n229 104.615
R249 source.n239 source.n229 104.615
R250 source.n240 source.n239 104.615
R251 source.n240 source.n225 104.615
R252 source.n247 source.n225 104.615
R253 source.n248 source.n247 104.615
R254 source.n200 source.n197 104.615
R255 source.n207 source.n197 104.615
R256 source.n208 source.n207 104.615
R257 source.n208 source.n193 104.615
R258 source.n215 source.n193 104.615
R259 source.n216 source.n215 104.615
R260 source.n158 source.n155 104.615
R261 source.n165 source.n155 104.615
R262 source.n166 source.n165 104.615
R263 source.n166 source.n151 104.615
R264 source.n173 source.n151 104.615
R265 source.n174 source.n173 104.615
R266 source.n26 source.n25 104.615
R267 source.n25 source.n3 104.615
R268 source.n18 source.n3 104.615
R269 source.n18 source.n17 104.615
R270 source.n17 source.n7 104.615
R271 source.n10 source.n7 104.615
R272 source.n68 source.n67 104.615
R273 source.n67 source.n45 104.615
R274 source.n60 source.n45 104.615
R275 source.n60 source.n59 104.615
R276 source.n59 source.n49 104.615
R277 source.n52 source.n49 104.615
R278 source.n100 source.n99 104.615
R279 source.n99 source.n77 104.615
R280 source.n92 source.n77 104.615
R281 source.n92 source.n91 104.615
R282 source.n91 source.n81 104.615
R283 source.n84 source.n81 104.615
R284 source.n142 source.n141 104.615
R285 source.n141 source.n119 104.615
R286 source.n134 source.n119 104.615
R287 source.n134 source.n133 104.615
R288 source.n133 source.n123 104.615
R289 source.n126 source.n123 104.615
R290 source.n274 source.t4 52.3082
R291 source.n232 source.t36 52.3082
R292 source.n200 source.t21 52.3082
R293 source.n158 source.t16 52.3082
R294 source.n10 source.t26 52.3082
R295 source.n52 source.t29 52.3082
R296 source.n84 source.t43 52.3082
R297 source.n126 source.t34 52.3082
R298 source.n33 source.n32 50.512
R299 source.n35 source.n34 50.512
R300 source.n37 source.n36 50.512
R301 source.n39 source.n38 50.512
R302 source.n41 source.n40 50.512
R303 source.n107 source.n106 50.512
R304 source.n109 source.n108 50.512
R305 source.n111 source.n110 50.512
R306 source.n113 source.n112 50.512
R307 source.n115 source.n114 50.512
R308 source.n263 source.n262 50.5119
R309 source.n261 source.n260 50.5119
R310 source.n259 source.n258 50.5119
R311 source.n257 source.n256 50.5119
R312 source.n255 source.n254 50.5119
R313 source.n189 source.n188 50.5119
R314 source.n187 source.n186 50.5119
R315 source.n185 source.n184 50.5119
R316 source.n183 source.n182 50.5119
R317 source.n181 source.n180 50.5119
R318 source.n295 source.n294 32.1853
R319 source.n253 source.n252 32.1853
R320 source.n221 source.n220 32.1853
R321 source.n179 source.n178 32.1853
R322 source.n31 source.n30 32.1853
R323 source.n73 source.n72 32.1853
R324 source.n105 source.n104 32.1853
R325 source.n147 source.n146 32.1853
R326 source.n179 source.n147 17.2854
R327 source.n275 source.n273 15.6674
R328 source.n233 source.n231 15.6674
R329 source.n201 source.n199 15.6674
R330 source.n159 source.n157 15.6674
R331 source.n11 source.n9 15.6674
R332 source.n53 source.n51 15.6674
R333 source.n85 source.n83 15.6674
R334 source.n127 source.n125 15.6674
R335 source.n276 source.n272 12.8005
R336 source.n234 source.n230 12.8005
R337 source.n202 source.n198 12.8005
R338 source.n160 source.n156 12.8005
R339 source.n12 source.n8 12.8005
R340 source.n54 source.n50 12.8005
R341 source.n86 source.n82 12.8005
R342 source.n128 source.n124 12.8005
R343 source.n280 source.n279 12.0247
R344 source.n238 source.n237 12.0247
R345 source.n206 source.n205 12.0247
R346 source.n164 source.n163 12.0247
R347 source.n16 source.n15 12.0247
R348 source.n58 source.n57 12.0247
R349 source.n90 source.n89 12.0247
R350 source.n132 source.n131 12.0247
R351 source.n296 source.n31 11.7509
R352 source.n283 source.n270 11.249
R353 source.n241 source.n228 11.249
R354 source.n209 source.n196 11.249
R355 source.n167 source.n154 11.249
R356 source.n19 source.n6 11.249
R357 source.n61 source.n48 11.249
R358 source.n93 source.n80 11.249
R359 source.n135 source.n122 11.249
R360 source.n284 source.n268 10.4732
R361 source.n242 source.n226 10.4732
R362 source.n210 source.n194 10.4732
R363 source.n168 source.n152 10.4732
R364 source.n20 source.n4 10.4732
R365 source.n62 source.n46 10.4732
R366 source.n94 source.n78 10.4732
R367 source.n136 source.n120 10.4732
R368 source.n288 source.n287 9.69747
R369 source.n246 source.n245 9.69747
R370 source.n214 source.n213 9.69747
R371 source.n172 source.n171 9.69747
R372 source.n24 source.n23 9.69747
R373 source.n66 source.n65 9.69747
R374 source.n98 source.n97 9.69747
R375 source.n140 source.n139 9.69747
R376 source.n294 source.n293 9.45567
R377 source.n252 source.n251 9.45567
R378 source.n220 source.n219 9.45567
R379 source.n178 source.n177 9.45567
R380 source.n30 source.n29 9.45567
R381 source.n72 source.n71 9.45567
R382 source.n104 source.n103 9.45567
R383 source.n146 source.n145 9.45567
R384 source.n293 source.n292 9.3005
R385 source.n266 source.n265 9.3005
R386 source.n287 source.n286 9.3005
R387 source.n285 source.n284 9.3005
R388 source.n270 source.n269 9.3005
R389 source.n279 source.n278 9.3005
R390 source.n277 source.n276 9.3005
R391 source.n251 source.n250 9.3005
R392 source.n224 source.n223 9.3005
R393 source.n245 source.n244 9.3005
R394 source.n243 source.n242 9.3005
R395 source.n228 source.n227 9.3005
R396 source.n237 source.n236 9.3005
R397 source.n235 source.n234 9.3005
R398 source.n219 source.n218 9.3005
R399 source.n192 source.n191 9.3005
R400 source.n213 source.n212 9.3005
R401 source.n211 source.n210 9.3005
R402 source.n196 source.n195 9.3005
R403 source.n205 source.n204 9.3005
R404 source.n203 source.n202 9.3005
R405 source.n177 source.n176 9.3005
R406 source.n150 source.n149 9.3005
R407 source.n171 source.n170 9.3005
R408 source.n169 source.n168 9.3005
R409 source.n154 source.n153 9.3005
R410 source.n163 source.n162 9.3005
R411 source.n161 source.n160 9.3005
R412 source.n29 source.n28 9.3005
R413 source.n2 source.n1 9.3005
R414 source.n23 source.n22 9.3005
R415 source.n21 source.n20 9.3005
R416 source.n6 source.n5 9.3005
R417 source.n15 source.n14 9.3005
R418 source.n13 source.n12 9.3005
R419 source.n71 source.n70 9.3005
R420 source.n44 source.n43 9.3005
R421 source.n65 source.n64 9.3005
R422 source.n63 source.n62 9.3005
R423 source.n48 source.n47 9.3005
R424 source.n57 source.n56 9.3005
R425 source.n55 source.n54 9.3005
R426 source.n103 source.n102 9.3005
R427 source.n76 source.n75 9.3005
R428 source.n97 source.n96 9.3005
R429 source.n95 source.n94 9.3005
R430 source.n80 source.n79 9.3005
R431 source.n89 source.n88 9.3005
R432 source.n87 source.n86 9.3005
R433 source.n145 source.n144 9.3005
R434 source.n118 source.n117 9.3005
R435 source.n139 source.n138 9.3005
R436 source.n137 source.n136 9.3005
R437 source.n122 source.n121 9.3005
R438 source.n131 source.n130 9.3005
R439 source.n129 source.n128 9.3005
R440 source.n291 source.n266 8.92171
R441 source.n249 source.n224 8.92171
R442 source.n217 source.n192 8.92171
R443 source.n175 source.n150 8.92171
R444 source.n27 source.n2 8.92171
R445 source.n69 source.n44 8.92171
R446 source.n101 source.n76 8.92171
R447 source.n143 source.n118 8.92171
R448 source.n292 source.n264 8.14595
R449 source.n250 source.n222 8.14595
R450 source.n218 source.n190 8.14595
R451 source.n176 source.n148 8.14595
R452 source.n28 source.n0 8.14595
R453 source.n70 source.n42 8.14595
R454 source.n102 source.n74 8.14595
R455 source.n144 source.n116 8.14595
R456 source.n294 source.n264 5.81868
R457 source.n252 source.n222 5.81868
R458 source.n220 source.n190 5.81868
R459 source.n178 source.n148 5.81868
R460 source.n30 source.n0 5.81868
R461 source.n72 source.n42 5.81868
R462 source.n104 source.n74 5.81868
R463 source.n146 source.n116 5.81868
R464 source.n296 source.n295 5.53498
R465 source.n292 source.n291 5.04292
R466 source.n250 source.n249 5.04292
R467 source.n218 source.n217 5.04292
R468 source.n176 source.n175 5.04292
R469 source.n28 source.n27 5.04292
R470 source.n70 source.n69 5.04292
R471 source.n102 source.n101 5.04292
R472 source.n144 source.n143 5.04292
R473 source.n277 source.n273 4.38594
R474 source.n235 source.n231 4.38594
R475 source.n203 source.n199 4.38594
R476 source.n161 source.n157 4.38594
R477 source.n13 source.n9 4.38594
R478 source.n55 source.n51 4.38594
R479 source.n87 source.n83 4.38594
R480 source.n129 source.n125 4.38594
R481 source.n288 source.n266 4.26717
R482 source.n246 source.n224 4.26717
R483 source.n214 source.n192 4.26717
R484 source.n172 source.n150 4.26717
R485 source.n24 source.n2 4.26717
R486 source.n66 source.n44 4.26717
R487 source.n98 source.n76 4.26717
R488 source.n140 source.n118 4.26717
R489 source.n287 source.n268 3.49141
R490 source.n245 source.n226 3.49141
R491 source.n213 source.n194 3.49141
R492 source.n171 source.n152 3.49141
R493 source.n23 source.n4 3.49141
R494 source.n65 source.n46 3.49141
R495 source.n97 source.n78 3.49141
R496 source.n139 source.n120 3.49141
R497 source.n262 source.t8 3.3005
R498 source.n262 source.t38 3.3005
R499 source.n260 source.t35 3.3005
R500 source.n260 source.t44 3.3005
R501 source.n258 source.t40 3.3005
R502 source.n258 source.t46 3.3005
R503 source.n256 source.t1 3.3005
R504 source.n256 source.t6 3.3005
R505 source.n254 source.t39 3.3005
R506 source.n254 source.t47 3.3005
R507 source.n188 source.t20 3.3005
R508 source.n188 source.t30 3.3005
R509 source.n186 source.t13 3.3005
R510 source.n186 source.t28 3.3005
R511 source.n184 source.t12 3.3005
R512 source.n184 source.t27 3.3005
R513 source.n182 source.t15 3.3005
R514 source.n182 source.t25 3.3005
R515 source.n180 source.t31 3.3005
R516 source.n180 source.t24 3.3005
R517 source.n32 source.t14 3.3005
R518 source.n32 source.t33 3.3005
R519 source.n34 source.t32 3.3005
R520 source.n34 source.t19 3.3005
R521 source.n36 source.t18 3.3005
R522 source.n36 source.t11 3.3005
R523 source.n38 source.t10 3.3005
R524 source.n38 source.t23 3.3005
R525 source.n40 source.t22 3.3005
R526 source.n40 source.t17 3.3005
R527 source.n106 source.t5 3.3005
R528 source.n106 source.t45 3.3005
R529 source.n108 source.t37 3.3005
R530 source.n108 source.t9 3.3005
R531 source.n110 source.t0 3.3005
R532 source.n110 source.t2 3.3005
R533 source.n112 source.t7 3.3005
R534 source.n112 source.t3 3.3005
R535 source.n114 source.t42 3.3005
R536 source.n114 source.t41 3.3005
R537 source.n284 source.n283 2.71565
R538 source.n242 source.n241 2.71565
R539 source.n210 source.n209 2.71565
R540 source.n168 source.n167 2.71565
R541 source.n20 source.n19 2.71565
R542 source.n62 source.n61 2.71565
R543 source.n94 source.n93 2.71565
R544 source.n136 source.n135 2.71565
R545 source.n280 source.n270 1.93989
R546 source.n238 source.n228 1.93989
R547 source.n206 source.n196 1.93989
R548 source.n164 source.n154 1.93989
R549 source.n16 source.n6 1.93989
R550 source.n58 source.n48 1.93989
R551 source.n90 source.n80 1.93989
R552 source.n132 source.n122 1.93989
R553 source.n279 source.n272 1.16414
R554 source.n237 source.n230 1.16414
R555 source.n205 source.n198 1.16414
R556 source.n163 source.n156 1.16414
R557 source.n15 source.n8 1.16414
R558 source.n57 source.n50 1.16414
R559 source.n89 source.n82 1.16414
R560 source.n131 source.n124 1.16414
R561 source.n147 source.n115 0.543603
R562 source.n115 source.n113 0.543603
R563 source.n113 source.n111 0.543603
R564 source.n111 source.n109 0.543603
R565 source.n109 source.n107 0.543603
R566 source.n107 source.n105 0.543603
R567 source.n73 source.n41 0.543603
R568 source.n41 source.n39 0.543603
R569 source.n39 source.n37 0.543603
R570 source.n37 source.n35 0.543603
R571 source.n35 source.n33 0.543603
R572 source.n33 source.n31 0.543603
R573 source.n181 source.n179 0.543603
R574 source.n183 source.n181 0.543603
R575 source.n185 source.n183 0.543603
R576 source.n187 source.n185 0.543603
R577 source.n189 source.n187 0.543603
R578 source.n221 source.n189 0.543603
R579 source.n255 source.n253 0.543603
R580 source.n257 source.n255 0.543603
R581 source.n259 source.n257 0.543603
R582 source.n261 source.n259 0.543603
R583 source.n263 source.n261 0.543603
R584 source.n295 source.n263 0.543603
R585 source.n105 source.n73 0.470328
R586 source.n253 source.n221 0.470328
R587 source.n276 source.n275 0.388379
R588 source.n234 source.n233 0.388379
R589 source.n202 source.n201 0.388379
R590 source.n160 source.n159 0.388379
R591 source.n12 source.n11 0.388379
R592 source.n54 source.n53 0.388379
R593 source.n86 source.n85 0.388379
R594 source.n128 source.n127 0.388379
R595 source source.n296 0.188
R596 source.n278 source.n277 0.155672
R597 source.n278 source.n269 0.155672
R598 source.n285 source.n269 0.155672
R599 source.n286 source.n285 0.155672
R600 source.n286 source.n265 0.155672
R601 source.n293 source.n265 0.155672
R602 source.n236 source.n235 0.155672
R603 source.n236 source.n227 0.155672
R604 source.n243 source.n227 0.155672
R605 source.n244 source.n243 0.155672
R606 source.n244 source.n223 0.155672
R607 source.n251 source.n223 0.155672
R608 source.n204 source.n203 0.155672
R609 source.n204 source.n195 0.155672
R610 source.n211 source.n195 0.155672
R611 source.n212 source.n211 0.155672
R612 source.n212 source.n191 0.155672
R613 source.n219 source.n191 0.155672
R614 source.n162 source.n161 0.155672
R615 source.n162 source.n153 0.155672
R616 source.n169 source.n153 0.155672
R617 source.n170 source.n169 0.155672
R618 source.n170 source.n149 0.155672
R619 source.n177 source.n149 0.155672
R620 source.n29 source.n1 0.155672
R621 source.n22 source.n1 0.155672
R622 source.n22 source.n21 0.155672
R623 source.n21 source.n5 0.155672
R624 source.n14 source.n5 0.155672
R625 source.n14 source.n13 0.155672
R626 source.n71 source.n43 0.155672
R627 source.n64 source.n43 0.155672
R628 source.n64 source.n63 0.155672
R629 source.n63 source.n47 0.155672
R630 source.n56 source.n47 0.155672
R631 source.n56 source.n55 0.155672
R632 source.n103 source.n75 0.155672
R633 source.n96 source.n75 0.155672
R634 source.n96 source.n95 0.155672
R635 source.n95 source.n79 0.155672
R636 source.n88 source.n79 0.155672
R637 source.n88 source.n87 0.155672
R638 source.n145 source.n117 0.155672
R639 source.n138 source.n117 0.155672
R640 source.n138 source.n137 0.155672
R641 source.n137 source.n121 0.155672
R642 source.n130 source.n121 0.155672
R643 source.n130 source.n129 0.155672
R644 minus.n35 minus.t5 617.837
R645 minus.n9 minus.t15 617.837
R646 minus.n72 minus.t18 617.837
R647 minus.n46 minus.t17 617.837
R648 minus.n34 minus.t21 586.433
R649 minus.n1 minus.t10 586.433
R650 minus.n28 minus.t4 586.433
R651 minus.n26 minus.t23 586.433
R652 minus.n3 minus.t7 586.433
R653 minus.n20 minus.t2 586.433
R654 minus.n5 minus.t20 586.433
R655 minus.n15 minus.t14 586.433
R656 minus.n13 minus.t3 586.433
R657 minus.n8 minus.t22 586.433
R658 minus.n71 minus.t6 586.433
R659 minus.n38 minus.t19 586.433
R660 minus.n65 minus.t11 586.433
R661 minus.n63 minus.t12 586.433
R662 minus.n40 minus.t0 586.433
R663 minus.n57 minus.t13 586.433
R664 minus.n42 minus.t1 586.433
R665 minus.n52 minus.t8 586.433
R666 minus.n50 minus.t16 586.433
R667 minus.n45 minus.t9 586.433
R668 minus.n10 minus.n9 161.489
R669 minus.n47 minus.n46 161.489
R670 minus.n36 minus.n35 161.3
R671 minus.n33 minus.n0 161.3
R672 minus.n32 minus.n31 161.3
R673 minus.n30 minus.n29 161.3
R674 minus.n27 minus.n2 161.3
R675 minus.n25 minus.n24 161.3
R676 minus.n23 minus.n22 161.3
R677 minus.n21 minus.n4 161.3
R678 minus.n19 minus.n18 161.3
R679 minus.n17 minus.n16 161.3
R680 minus.n14 minus.n6 161.3
R681 minus.n12 minus.n11 161.3
R682 minus.n10 minus.n7 161.3
R683 minus.n73 minus.n72 161.3
R684 minus.n70 minus.n37 161.3
R685 minus.n69 minus.n68 161.3
R686 minus.n67 minus.n66 161.3
R687 minus.n64 minus.n39 161.3
R688 minus.n62 minus.n61 161.3
R689 minus.n60 minus.n59 161.3
R690 minus.n58 minus.n41 161.3
R691 minus.n56 minus.n55 161.3
R692 minus.n54 minus.n53 161.3
R693 minus.n51 minus.n43 161.3
R694 minus.n49 minus.n48 161.3
R695 minus.n47 minus.n44 161.3
R696 minus.n33 minus.n32 73.0308
R697 minus.n22 minus.n21 73.0308
R698 minus.n12 minus.n7 73.0308
R699 minus.n49 minus.n44 73.0308
R700 minus.n59 minus.n58 73.0308
R701 minus.n70 minus.n69 73.0308
R702 minus.n29 minus.n1 66.4581
R703 minus.n14 minus.n13 66.4581
R704 minus.n51 minus.n50 66.4581
R705 minus.n66 minus.n38 66.4581
R706 minus.n25 minus.n3 63.5369
R707 minus.n20 minus.n19 63.5369
R708 minus.n57 minus.n56 63.5369
R709 minus.n62 minus.n40 63.5369
R710 minus.n35 minus.n34 60.6157
R711 minus.n9 minus.n8 60.6157
R712 minus.n46 minus.n45 60.6157
R713 minus.n72 minus.n71 60.6157
R714 minus.n28 minus.n27 47.4702
R715 minus.n16 minus.n15 47.4702
R716 minus.n53 minus.n52 47.4702
R717 minus.n65 minus.n64 47.4702
R718 minus.n27 minus.n26 44.549
R719 minus.n16 minus.n5 44.549
R720 minus.n53 minus.n42 44.549
R721 minus.n64 minus.n63 44.549
R722 minus.n74 minus.n36 33.4626
R723 minus.n26 minus.n25 28.4823
R724 minus.n19 minus.n5 28.4823
R725 minus.n56 minus.n42 28.4823
R726 minus.n63 minus.n62 28.4823
R727 minus.n29 minus.n28 25.5611
R728 minus.n15 minus.n14 25.5611
R729 minus.n52 minus.n51 25.5611
R730 minus.n66 minus.n65 25.5611
R731 minus.n34 minus.n33 12.4157
R732 minus.n8 minus.n7 12.4157
R733 minus.n45 minus.n44 12.4157
R734 minus.n71 minus.n70 12.4157
R735 minus.n22 minus.n3 9.49444
R736 minus.n21 minus.n20 9.49444
R737 minus.n58 minus.n57 9.49444
R738 minus.n59 minus.n40 9.49444
R739 minus.n32 minus.n1 6.57323
R740 minus.n13 minus.n12 6.57323
R741 minus.n50 minus.n49 6.57323
R742 minus.n69 minus.n38 6.57323
R743 minus.n74 minus.n73 6.4702
R744 minus.n36 minus.n0 0.189894
R745 minus.n31 minus.n0 0.189894
R746 minus.n31 minus.n30 0.189894
R747 minus.n30 minus.n2 0.189894
R748 minus.n24 minus.n2 0.189894
R749 minus.n24 minus.n23 0.189894
R750 minus.n23 minus.n4 0.189894
R751 minus.n18 minus.n4 0.189894
R752 minus.n18 minus.n17 0.189894
R753 minus.n17 minus.n6 0.189894
R754 minus.n11 minus.n6 0.189894
R755 minus.n11 minus.n10 0.189894
R756 minus.n48 minus.n47 0.189894
R757 minus.n48 minus.n43 0.189894
R758 minus.n54 minus.n43 0.189894
R759 minus.n55 minus.n54 0.189894
R760 minus.n55 minus.n41 0.189894
R761 minus.n60 minus.n41 0.189894
R762 minus.n61 minus.n60 0.189894
R763 minus.n61 minus.n39 0.189894
R764 minus.n67 minus.n39 0.189894
R765 minus.n68 minus.n67 0.189894
R766 minus.n68 minus.n37 0.189894
R767 minus.n73 minus.n37 0.189894
R768 minus minus.n74 0.188
R769 drain_right.n7 drain_right.n5 67.7338
R770 drain_right.n2 drain_right.n0 67.7338
R771 drain_right.n13 drain_right.n11 67.7338
R772 drain_right.n13 drain_right.n12 67.1908
R773 drain_right.n15 drain_right.n14 67.1908
R774 drain_right.n17 drain_right.n16 67.1908
R775 drain_right.n19 drain_right.n18 67.1908
R776 drain_right.n21 drain_right.n20 67.1908
R777 drain_right.n7 drain_right.n6 67.1907
R778 drain_right.n9 drain_right.n8 67.1907
R779 drain_right.n4 drain_right.n3 67.1907
R780 drain_right.n2 drain_right.n1 67.1907
R781 drain_right drain_right.n10 27.4279
R782 drain_right drain_right.n21 6.19632
R783 drain_right.n5 drain_right.t17 3.3005
R784 drain_right.n5 drain_right.t5 3.3005
R785 drain_right.n6 drain_right.t12 3.3005
R786 drain_right.n6 drain_right.t4 3.3005
R787 drain_right.n8 drain_right.t23 3.3005
R788 drain_right.n8 drain_right.t11 3.3005
R789 drain_right.n3 drain_right.t22 3.3005
R790 drain_right.n3 drain_right.t10 3.3005
R791 drain_right.n1 drain_right.t7 3.3005
R792 drain_right.n1 drain_right.t15 3.3005
R793 drain_right.n0 drain_right.t6 3.3005
R794 drain_right.n0 drain_right.t14 3.3005
R795 drain_right.n11 drain_right.t1 3.3005
R796 drain_right.n11 drain_right.t8 3.3005
R797 drain_right.n12 drain_right.t9 3.3005
R798 drain_right.n12 drain_right.t20 3.3005
R799 drain_right.n14 drain_right.t21 3.3005
R800 drain_right.n14 drain_right.t3 3.3005
R801 drain_right.n16 drain_right.t0 3.3005
R802 drain_right.n16 drain_right.t16 3.3005
R803 drain_right.n18 drain_right.t13 3.3005
R804 drain_right.n18 drain_right.t19 3.3005
R805 drain_right.n20 drain_right.t18 3.3005
R806 drain_right.n20 drain_right.t2 3.3005
R807 drain_right.n9 drain_right.n7 0.543603
R808 drain_right.n4 drain_right.n2 0.543603
R809 drain_right.n21 drain_right.n19 0.543603
R810 drain_right.n19 drain_right.n17 0.543603
R811 drain_right.n17 drain_right.n15 0.543603
R812 drain_right.n15 drain_right.n13 0.543603
R813 drain_right.n10 drain_right.n9 0.216706
R814 drain_right.n10 drain_right.n4 0.216706
C0 source drain_left 24.123802f
C1 plus minus 4.9829f
C2 drain_right minus 4.55793f
C3 source plus 4.7077f
C4 source drain_right 24.1244f
C5 drain_left plus 4.79013f
C6 drain_right drain_left 1.26597f
C7 source minus 4.69368f
C8 drain_right plus 0.387992f
C9 drain_left minus 0.172624f
C10 drain_right a_n2354_n2088# 6.01797f
C11 drain_left a_n2354_n2088# 6.37083f
C12 source a_n2354_n2088# 5.543537f
C13 minus a_n2354_n2088# 8.787163f
C14 plus a_n2354_n2088# 10.468611f
C15 drain_right.t6 a_n2354_n2088# 0.159782f
C16 drain_right.t14 a_n2354_n2088# 0.159782f
C17 drain_right.n0 a_n2354_n2088# 1.33583f
C18 drain_right.t7 a_n2354_n2088# 0.159782f
C19 drain_right.t15 a_n2354_n2088# 0.159782f
C20 drain_right.n1 a_n2354_n2088# 1.33259f
C21 drain_right.n2 a_n2354_n2088# 0.793257f
C22 drain_right.t22 a_n2354_n2088# 0.159782f
C23 drain_right.t10 a_n2354_n2088# 0.159782f
C24 drain_right.n3 a_n2354_n2088# 1.33259f
C25 drain_right.n4 a_n2354_n2088# 0.359582f
C26 drain_right.t17 a_n2354_n2088# 0.159782f
C27 drain_right.t5 a_n2354_n2088# 0.159782f
C28 drain_right.n5 a_n2354_n2088# 1.33583f
C29 drain_right.t12 a_n2354_n2088# 0.159782f
C30 drain_right.t4 a_n2354_n2088# 0.159782f
C31 drain_right.n6 a_n2354_n2088# 1.33259f
C32 drain_right.n7 a_n2354_n2088# 0.793257f
C33 drain_right.t23 a_n2354_n2088# 0.159782f
C34 drain_right.t11 a_n2354_n2088# 0.159782f
C35 drain_right.n8 a_n2354_n2088# 1.33259f
C36 drain_right.n9 a_n2354_n2088# 0.359582f
C37 drain_right.n10 a_n2354_n2088# 1.31787f
C38 drain_right.t1 a_n2354_n2088# 0.159782f
C39 drain_right.t8 a_n2354_n2088# 0.159782f
C40 drain_right.n11 a_n2354_n2088# 1.33583f
C41 drain_right.t9 a_n2354_n2088# 0.159782f
C42 drain_right.t20 a_n2354_n2088# 0.159782f
C43 drain_right.n12 a_n2354_n2088# 1.33259f
C44 drain_right.n13 a_n2354_n2088# 0.793251f
C45 drain_right.t21 a_n2354_n2088# 0.159782f
C46 drain_right.t3 a_n2354_n2088# 0.159782f
C47 drain_right.n14 a_n2354_n2088# 1.33259f
C48 drain_right.n15 a_n2354_n2088# 0.391459f
C49 drain_right.t0 a_n2354_n2088# 0.159782f
C50 drain_right.t16 a_n2354_n2088# 0.159782f
C51 drain_right.n16 a_n2354_n2088# 1.33259f
C52 drain_right.n17 a_n2354_n2088# 0.391459f
C53 drain_right.t13 a_n2354_n2088# 0.159782f
C54 drain_right.t19 a_n2354_n2088# 0.159782f
C55 drain_right.n18 a_n2354_n2088# 1.33259f
C56 drain_right.n19 a_n2354_n2088# 0.391459f
C57 drain_right.t18 a_n2354_n2088# 0.159782f
C58 drain_right.t2 a_n2354_n2088# 0.159782f
C59 drain_right.n20 a_n2354_n2088# 1.33259f
C60 drain_right.n21 a_n2354_n2088# 0.671961f
C61 minus.n0 a_n2354_n2088# 0.048734f
C62 minus.t5 a_n2354_n2088# 0.255785f
C63 minus.t21 a_n2354_n2088# 0.249932f
C64 minus.t10 a_n2354_n2088# 0.249932f
C65 minus.n1 a_n2354_n2088# 0.114723f
C66 minus.n2 a_n2354_n2088# 0.048734f
C67 minus.t4 a_n2354_n2088# 0.249932f
C68 minus.t23 a_n2354_n2088# 0.249932f
C69 minus.t7 a_n2354_n2088# 0.249932f
C70 minus.n3 a_n2354_n2088# 0.114723f
C71 minus.n4 a_n2354_n2088# 0.048734f
C72 minus.t2 a_n2354_n2088# 0.249932f
C73 minus.t20 a_n2354_n2088# 0.249932f
C74 minus.n5 a_n2354_n2088# 0.114723f
C75 minus.n6 a_n2354_n2088# 0.048734f
C76 minus.t14 a_n2354_n2088# 0.249932f
C77 minus.t3 a_n2354_n2088# 0.249932f
C78 minus.n7 a_n2354_n2088# 0.018721f
C79 minus.t22 a_n2354_n2088# 0.249932f
C80 minus.n8 a_n2354_n2088# 0.114723f
C81 minus.t15 a_n2354_n2088# 0.255785f
C82 minus.n9 a_n2354_n2088# 0.129457f
C83 minus.n10 a_n2354_n2088# 0.104313f
C84 minus.n11 a_n2354_n2088# 0.048734f
C85 minus.n12 a_n2354_n2088# 0.017519f
C86 minus.n13 a_n2354_n2088# 0.114723f
C87 minus.n14 a_n2354_n2088# 0.020073f
C88 minus.n15 a_n2354_n2088# 0.114723f
C89 minus.n16 a_n2354_n2088# 0.020073f
C90 minus.n17 a_n2354_n2088# 0.048734f
C91 minus.n18 a_n2354_n2088# 0.048734f
C92 minus.n19 a_n2354_n2088# 0.020073f
C93 minus.n20 a_n2354_n2088# 0.114723f
C94 minus.n21 a_n2354_n2088# 0.01812f
C95 minus.n22 a_n2354_n2088# 0.01812f
C96 minus.n23 a_n2354_n2088# 0.048734f
C97 minus.n24 a_n2354_n2088# 0.048734f
C98 minus.n25 a_n2354_n2088# 0.020073f
C99 minus.n26 a_n2354_n2088# 0.114723f
C100 minus.n27 a_n2354_n2088# 0.020073f
C101 minus.n28 a_n2354_n2088# 0.114723f
C102 minus.n29 a_n2354_n2088# 0.020073f
C103 minus.n30 a_n2354_n2088# 0.048734f
C104 minus.n31 a_n2354_n2088# 0.048734f
C105 minus.n32 a_n2354_n2088# 0.017519f
C106 minus.n33 a_n2354_n2088# 0.018721f
C107 minus.n34 a_n2354_n2088# 0.114723f
C108 minus.n35 a_n2354_n2088# 0.129392f
C109 minus.n36 a_n2354_n2088# 1.51898f
C110 minus.n37 a_n2354_n2088# 0.048734f
C111 minus.t6 a_n2354_n2088# 0.249932f
C112 minus.t19 a_n2354_n2088# 0.249932f
C113 minus.n38 a_n2354_n2088# 0.114723f
C114 minus.n39 a_n2354_n2088# 0.048734f
C115 minus.t11 a_n2354_n2088# 0.249932f
C116 minus.t12 a_n2354_n2088# 0.249932f
C117 minus.t0 a_n2354_n2088# 0.249932f
C118 minus.n40 a_n2354_n2088# 0.114723f
C119 minus.n41 a_n2354_n2088# 0.048734f
C120 minus.t13 a_n2354_n2088# 0.249932f
C121 minus.t1 a_n2354_n2088# 0.249932f
C122 minus.n42 a_n2354_n2088# 0.114723f
C123 minus.n43 a_n2354_n2088# 0.048734f
C124 minus.t8 a_n2354_n2088# 0.249932f
C125 minus.t16 a_n2354_n2088# 0.249932f
C126 minus.n44 a_n2354_n2088# 0.018721f
C127 minus.t17 a_n2354_n2088# 0.255785f
C128 minus.t9 a_n2354_n2088# 0.249932f
C129 minus.n45 a_n2354_n2088# 0.114723f
C130 minus.n46 a_n2354_n2088# 0.129457f
C131 minus.n47 a_n2354_n2088# 0.104313f
C132 minus.n48 a_n2354_n2088# 0.048734f
C133 minus.n49 a_n2354_n2088# 0.017519f
C134 minus.n50 a_n2354_n2088# 0.114723f
C135 minus.n51 a_n2354_n2088# 0.020073f
C136 minus.n52 a_n2354_n2088# 0.114723f
C137 minus.n53 a_n2354_n2088# 0.020073f
C138 minus.n54 a_n2354_n2088# 0.048734f
C139 minus.n55 a_n2354_n2088# 0.048734f
C140 minus.n56 a_n2354_n2088# 0.020073f
C141 minus.n57 a_n2354_n2088# 0.114723f
C142 minus.n58 a_n2354_n2088# 0.01812f
C143 minus.n59 a_n2354_n2088# 0.01812f
C144 minus.n60 a_n2354_n2088# 0.048734f
C145 minus.n61 a_n2354_n2088# 0.048734f
C146 minus.n62 a_n2354_n2088# 0.020073f
C147 minus.n63 a_n2354_n2088# 0.114723f
C148 minus.n64 a_n2354_n2088# 0.020073f
C149 minus.n65 a_n2354_n2088# 0.114723f
C150 minus.n66 a_n2354_n2088# 0.020073f
C151 minus.n67 a_n2354_n2088# 0.048734f
C152 minus.n68 a_n2354_n2088# 0.048734f
C153 minus.n69 a_n2354_n2088# 0.017519f
C154 minus.n70 a_n2354_n2088# 0.018721f
C155 minus.n71 a_n2354_n2088# 0.114723f
C156 minus.t18 a_n2354_n2088# 0.255785f
C157 minus.n72 a_n2354_n2088# 0.129392f
C158 minus.n73 a_n2354_n2088# 0.315182f
C159 minus.n74 a_n2354_n2088# 1.86083f
C160 source.n0 a_n2354_n2088# 0.044486f
C161 source.n1 a_n2354_n2088# 0.03165f
C162 source.n2 a_n2354_n2088# 0.017007f
C163 source.n3 a_n2354_n2088# 0.040199f
C164 source.n4 a_n2354_n2088# 0.018008f
C165 source.n5 a_n2354_n2088# 0.03165f
C166 source.n6 a_n2354_n2088# 0.017007f
C167 source.n7 a_n2354_n2088# 0.040199f
C168 source.n8 a_n2354_n2088# 0.018008f
C169 source.n9 a_n2354_n2088# 0.135438f
C170 source.t26 a_n2354_n2088# 0.065518f
C171 source.n10 a_n2354_n2088# 0.030149f
C172 source.n11 a_n2354_n2088# 0.023745f
C173 source.n12 a_n2354_n2088# 0.017007f
C174 source.n13 a_n2354_n2088# 0.753071f
C175 source.n14 a_n2354_n2088# 0.03165f
C176 source.n15 a_n2354_n2088# 0.017007f
C177 source.n16 a_n2354_n2088# 0.018008f
C178 source.n17 a_n2354_n2088# 0.040199f
C179 source.n18 a_n2354_n2088# 0.040199f
C180 source.n19 a_n2354_n2088# 0.018008f
C181 source.n20 a_n2354_n2088# 0.017007f
C182 source.n21 a_n2354_n2088# 0.03165f
C183 source.n22 a_n2354_n2088# 0.03165f
C184 source.n23 a_n2354_n2088# 0.017007f
C185 source.n24 a_n2354_n2088# 0.018008f
C186 source.n25 a_n2354_n2088# 0.040199f
C187 source.n26 a_n2354_n2088# 0.087023f
C188 source.n27 a_n2354_n2088# 0.018008f
C189 source.n28 a_n2354_n2088# 0.017007f
C190 source.n29 a_n2354_n2088# 0.073156f
C191 source.n30 a_n2354_n2088# 0.048693f
C192 source.n31 a_n2354_n2088# 0.766616f
C193 source.t14 a_n2354_n2088# 0.150063f
C194 source.t33 a_n2354_n2088# 0.150063f
C195 source.n32 a_n2354_n2088# 1.1687f
C196 source.n33 a_n2354_n2088# 0.407458f
C197 source.t32 a_n2354_n2088# 0.150063f
C198 source.t19 a_n2354_n2088# 0.150063f
C199 source.n34 a_n2354_n2088# 1.1687f
C200 source.n35 a_n2354_n2088# 0.407458f
C201 source.t18 a_n2354_n2088# 0.150063f
C202 source.t11 a_n2354_n2088# 0.150063f
C203 source.n36 a_n2354_n2088# 1.1687f
C204 source.n37 a_n2354_n2088# 0.407458f
C205 source.t10 a_n2354_n2088# 0.150063f
C206 source.t23 a_n2354_n2088# 0.150063f
C207 source.n38 a_n2354_n2088# 1.1687f
C208 source.n39 a_n2354_n2088# 0.407458f
C209 source.t22 a_n2354_n2088# 0.150063f
C210 source.t17 a_n2354_n2088# 0.150063f
C211 source.n40 a_n2354_n2088# 1.1687f
C212 source.n41 a_n2354_n2088# 0.407458f
C213 source.n42 a_n2354_n2088# 0.044486f
C214 source.n43 a_n2354_n2088# 0.03165f
C215 source.n44 a_n2354_n2088# 0.017007f
C216 source.n45 a_n2354_n2088# 0.040199f
C217 source.n46 a_n2354_n2088# 0.018008f
C218 source.n47 a_n2354_n2088# 0.03165f
C219 source.n48 a_n2354_n2088# 0.017007f
C220 source.n49 a_n2354_n2088# 0.040199f
C221 source.n50 a_n2354_n2088# 0.018008f
C222 source.n51 a_n2354_n2088# 0.135438f
C223 source.t29 a_n2354_n2088# 0.065518f
C224 source.n52 a_n2354_n2088# 0.030149f
C225 source.n53 a_n2354_n2088# 0.023745f
C226 source.n54 a_n2354_n2088# 0.017007f
C227 source.n55 a_n2354_n2088# 0.753071f
C228 source.n56 a_n2354_n2088# 0.03165f
C229 source.n57 a_n2354_n2088# 0.017007f
C230 source.n58 a_n2354_n2088# 0.018008f
C231 source.n59 a_n2354_n2088# 0.040199f
C232 source.n60 a_n2354_n2088# 0.040199f
C233 source.n61 a_n2354_n2088# 0.018008f
C234 source.n62 a_n2354_n2088# 0.017007f
C235 source.n63 a_n2354_n2088# 0.03165f
C236 source.n64 a_n2354_n2088# 0.03165f
C237 source.n65 a_n2354_n2088# 0.017007f
C238 source.n66 a_n2354_n2088# 0.018008f
C239 source.n67 a_n2354_n2088# 0.040199f
C240 source.n68 a_n2354_n2088# 0.087023f
C241 source.n69 a_n2354_n2088# 0.018008f
C242 source.n70 a_n2354_n2088# 0.017007f
C243 source.n71 a_n2354_n2088# 0.073156f
C244 source.n72 a_n2354_n2088# 0.048693f
C245 source.n73 a_n2354_n2088# 0.130332f
C246 source.n74 a_n2354_n2088# 0.044486f
C247 source.n75 a_n2354_n2088# 0.03165f
C248 source.n76 a_n2354_n2088# 0.017007f
C249 source.n77 a_n2354_n2088# 0.040199f
C250 source.n78 a_n2354_n2088# 0.018008f
C251 source.n79 a_n2354_n2088# 0.03165f
C252 source.n80 a_n2354_n2088# 0.017007f
C253 source.n81 a_n2354_n2088# 0.040199f
C254 source.n82 a_n2354_n2088# 0.018008f
C255 source.n83 a_n2354_n2088# 0.135438f
C256 source.t43 a_n2354_n2088# 0.065518f
C257 source.n84 a_n2354_n2088# 0.030149f
C258 source.n85 a_n2354_n2088# 0.023745f
C259 source.n86 a_n2354_n2088# 0.017007f
C260 source.n87 a_n2354_n2088# 0.753071f
C261 source.n88 a_n2354_n2088# 0.03165f
C262 source.n89 a_n2354_n2088# 0.017007f
C263 source.n90 a_n2354_n2088# 0.018008f
C264 source.n91 a_n2354_n2088# 0.040199f
C265 source.n92 a_n2354_n2088# 0.040199f
C266 source.n93 a_n2354_n2088# 0.018008f
C267 source.n94 a_n2354_n2088# 0.017007f
C268 source.n95 a_n2354_n2088# 0.03165f
C269 source.n96 a_n2354_n2088# 0.03165f
C270 source.n97 a_n2354_n2088# 0.017007f
C271 source.n98 a_n2354_n2088# 0.018008f
C272 source.n99 a_n2354_n2088# 0.040199f
C273 source.n100 a_n2354_n2088# 0.087023f
C274 source.n101 a_n2354_n2088# 0.018008f
C275 source.n102 a_n2354_n2088# 0.017007f
C276 source.n103 a_n2354_n2088# 0.073156f
C277 source.n104 a_n2354_n2088# 0.048693f
C278 source.n105 a_n2354_n2088# 0.130332f
C279 source.t5 a_n2354_n2088# 0.150063f
C280 source.t45 a_n2354_n2088# 0.150063f
C281 source.n106 a_n2354_n2088# 1.1687f
C282 source.n107 a_n2354_n2088# 0.407458f
C283 source.t37 a_n2354_n2088# 0.150063f
C284 source.t9 a_n2354_n2088# 0.150063f
C285 source.n108 a_n2354_n2088# 1.1687f
C286 source.n109 a_n2354_n2088# 0.407458f
C287 source.t0 a_n2354_n2088# 0.150063f
C288 source.t2 a_n2354_n2088# 0.150063f
C289 source.n110 a_n2354_n2088# 1.1687f
C290 source.n111 a_n2354_n2088# 0.407458f
C291 source.t7 a_n2354_n2088# 0.150063f
C292 source.t3 a_n2354_n2088# 0.150063f
C293 source.n112 a_n2354_n2088# 1.1687f
C294 source.n113 a_n2354_n2088# 0.407458f
C295 source.t42 a_n2354_n2088# 0.150063f
C296 source.t41 a_n2354_n2088# 0.150063f
C297 source.n114 a_n2354_n2088# 1.1687f
C298 source.n115 a_n2354_n2088# 0.407458f
C299 source.n116 a_n2354_n2088# 0.044486f
C300 source.n117 a_n2354_n2088# 0.03165f
C301 source.n118 a_n2354_n2088# 0.017007f
C302 source.n119 a_n2354_n2088# 0.040199f
C303 source.n120 a_n2354_n2088# 0.018008f
C304 source.n121 a_n2354_n2088# 0.03165f
C305 source.n122 a_n2354_n2088# 0.017007f
C306 source.n123 a_n2354_n2088# 0.040199f
C307 source.n124 a_n2354_n2088# 0.018008f
C308 source.n125 a_n2354_n2088# 0.135438f
C309 source.t34 a_n2354_n2088# 0.065518f
C310 source.n126 a_n2354_n2088# 0.030149f
C311 source.n127 a_n2354_n2088# 0.023745f
C312 source.n128 a_n2354_n2088# 0.017007f
C313 source.n129 a_n2354_n2088# 0.753071f
C314 source.n130 a_n2354_n2088# 0.03165f
C315 source.n131 a_n2354_n2088# 0.017007f
C316 source.n132 a_n2354_n2088# 0.018008f
C317 source.n133 a_n2354_n2088# 0.040199f
C318 source.n134 a_n2354_n2088# 0.040199f
C319 source.n135 a_n2354_n2088# 0.018008f
C320 source.n136 a_n2354_n2088# 0.017007f
C321 source.n137 a_n2354_n2088# 0.03165f
C322 source.n138 a_n2354_n2088# 0.03165f
C323 source.n139 a_n2354_n2088# 0.017007f
C324 source.n140 a_n2354_n2088# 0.018008f
C325 source.n141 a_n2354_n2088# 0.040199f
C326 source.n142 a_n2354_n2088# 0.087023f
C327 source.n143 a_n2354_n2088# 0.018008f
C328 source.n144 a_n2354_n2088# 0.017007f
C329 source.n145 a_n2354_n2088# 0.073156f
C330 source.n146 a_n2354_n2088# 0.048693f
C331 source.n147 a_n2354_n2088# 1.17407f
C332 source.n148 a_n2354_n2088# 0.044486f
C333 source.n149 a_n2354_n2088# 0.03165f
C334 source.n150 a_n2354_n2088# 0.017007f
C335 source.n151 a_n2354_n2088# 0.040199f
C336 source.n152 a_n2354_n2088# 0.018008f
C337 source.n153 a_n2354_n2088# 0.03165f
C338 source.n154 a_n2354_n2088# 0.017007f
C339 source.n155 a_n2354_n2088# 0.040199f
C340 source.n156 a_n2354_n2088# 0.018008f
C341 source.n157 a_n2354_n2088# 0.135438f
C342 source.t16 a_n2354_n2088# 0.065518f
C343 source.n158 a_n2354_n2088# 0.030149f
C344 source.n159 a_n2354_n2088# 0.023745f
C345 source.n160 a_n2354_n2088# 0.017007f
C346 source.n161 a_n2354_n2088# 0.753071f
C347 source.n162 a_n2354_n2088# 0.03165f
C348 source.n163 a_n2354_n2088# 0.017007f
C349 source.n164 a_n2354_n2088# 0.018008f
C350 source.n165 a_n2354_n2088# 0.040199f
C351 source.n166 a_n2354_n2088# 0.040199f
C352 source.n167 a_n2354_n2088# 0.018008f
C353 source.n168 a_n2354_n2088# 0.017007f
C354 source.n169 a_n2354_n2088# 0.03165f
C355 source.n170 a_n2354_n2088# 0.03165f
C356 source.n171 a_n2354_n2088# 0.017007f
C357 source.n172 a_n2354_n2088# 0.018008f
C358 source.n173 a_n2354_n2088# 0.040199f
C359 source.n174 a_n2354_n2088# 0.087023f
C360 source.n175 a_n2354_n2088# 0.018008f
C361 source.n176 a_n2354_n2088# 0.017007f
C362 source.n177 a_n2354_n2088# 0.073156f
C363 source.n178 a_n2354_n2088# 0.048693f
C364 source.n179 a_n2354_n2088# 1.17407f
C365 source.t31 a_n2354_n2088# 0.150063f
C366 source.t24 a_n2354_n2088# 0.150063f
C367 source.n180 a_n2354_n2088# 1.16869f
C368 source.n181 a_n2354_n2088# 0.407466f
C369 source.t15 a_n2354_n2088# 0.150063f
C370 source.t25 a_n2354_n2088# 0.150063f
C371 source.n182 a_n2354_n2088# 1.16869f
C372 source.n183 a_n2354_n2088# 0.407466f
C373 source.t12 a_n2354_n2088# 0.150063f
C374 source.t27 a_n2354_n2088# 0.150063f
C375 source.n184 a_n2354_n2088# 1.16869f
C376 source.n185 a_n2354_n2088# 0.407466f
C377 source.t13 a_n2354_n2088# 0.150063f
C378 source.t28 a_n2354_n2088# 0.150063f
C379 source.n186 a_n2354_n2088# 1.16869f
C380 source.n187 a_n2354_n2088# 0.407466f
C381 source.t20 a_n2354_n2088# 0.150063f
C382 source.t30 a_n2354_n2088# 0.150063f
C383 source.n188 a_n2354_n2088# 1.16869f
C384 source.n189 a_n2354_n2088# 0.407466f
C385 source.n190 a_n2354_n2088# 0.044486f
C386 source.n191 a_n2354_n2088# 0.03165f
C387 source.n192 a_n2354_n2088# 0.017007f
C388 source.n193 a_n2354_n2088# 0.040199f
C389 source.n194 a_n2354_n2088# 0.018008f
C390 source.n195 a_n2354_n2088# 0.03165f
C391 source.n196 a_n2354_n2088# 0.017007f
C392 source.n197 a_n2354_n2088# 0.040199f
C393 source.n198 a_n2354_n2088# 0.018008f
C394 source.n199 a_n2354_n2088# 0.135438f
C395 source.t21 a_n2354_n2088# 0.065518f
C396 source.n200 a_n2354_n2088# 0.030149f
C397 source.n201 a_n2354_n2088# 0.023745f
C398 source.n202 a_n2354_n2088# 0.017007f
C399 source.n203 a_n2354_n2088# 0.753071f
C400 source.n204 a_n2354_n2088# 0.03165f
C401 source.n205 a_n2354_n2088# 0.017007f
C402 source.n206 a_n2354_n2088# 0.018008f
C403 source.n207 a_n2354_n2088# 0.040199f
C404 source.n208 a_n2354_n2088# 0.040199f
C405 source.n209 a_n2354_n2088# 0.018008f
C406 source.n210 a_n2354_n2088# 0.017007f
C407 source.n211 a_n2354_n2088# 0.03165f
C408 source.n212 a_n2354_n2088# 0.03165f
C409 source.n213 a_n2354_n2088# 0.017007f
C410 source.n214 a_n2354_n2088# 0.018008f
C411 source.n215 a_n2354_n2088# 0.040199f
C412 source.n216 a_n2354_n2088# 0.087023f
C413 source.n217 a_n2354_n2088# 0.018008f
C414 source.n218 a_n2354_n2088# 0.017007f
C415 source.n219 a_n2354_n2088# 0.073156f
C416 source.n220 a_n2354_n2088# 0.048693f
C417 source.n221 a_n2354_n2088# 0.130332f
C418 source.n222 a_n2354_n2088# 0.044486f
C419 source.n223 a_n2354_n2088# 0.03165f
C420 source.n224 a_n2354_n2088# 0.017007f
C421 source.n225 a_n2354_n2088# 0.040199f
C422 source.n226 a_n2354_n2088# 0.018008f
C423 source.n227 a_n2354_n2088# 0.03165f
C424 source.n228 a_n2354_n2088# 0.017007f
C425 source.n229 a_n2354_n2088# 0.040199f
C426 source.n230 a_n2354_n2088# 0.018008f
C427 source.n231 a_n2354_n2088# 0.135438f
C428 source.t36 a_n2354_n2088# 0.065518f
C429 source.n232 a_n2354_n2088# 0.030149f
C430 source.n233 a_n2354_n2088# 0.023745f
C431 source.n234 a_n2354_n2088# 0.017007f
C432 source.n235 a_n2354_n2088# 0.753071f
C433 source.n236 a_n2354_n2088# 0.03165f
C434 source.n237 a_n2354_n2088# 0.017007f
C435 source.n238 a_n2354_n2088# 0.018008f
C436 source.n239 a_n2354_n2088# 0.040199f
C437 source.n240 a_n2354_n2088# 0.040199f
C438 source.n241 a_n2354_n2088# 0.018008f
C439 source.n242 a_n2354_n2088# 0.017007f
C440 source.n243 a_n2354_n2088# 0.03165f
C441 source.n244 a_n2354_n2088# 0.03165f
C442 source.n245 a_n2354_n2088# 0.017007f
C443 source.n246 a_n2354_n2088# 0.018008f
C444 source.n247 a_n2354_n2088# 0.040199f
C445 source.n248 a_n2354_n2088# 0.087023f
C446 source.n249 a_n2354_n2088# 0.018008f
C447 source.n250 a_n2354_n2088# 0.017007f
C448 source.n251 a_n2354_n2088# 0.073156f
C449 source.n252 a_n2354_n2088# 0.048693f
C450 source.n253 a_n2354_n2088# 0.130332f
C451 source.t39 a_n2354_n2088# 0.150063f
C452 source.t47 a_n2354_n2088# 0.150063f
C453 source.n254 a_n2354_n2088# 1.16869f
C454 source.n255 a_n2354_n2088# 0.407466f
C455 source.t1 a_n2354_n2088# 0.150063f
C456 source.t6 a_n2354_n2088# 0.150063f
C457 source.n256 a_n2354_n2088# 1.16869f
C458 source.n257 a_n2354_n2088# 0.407466f
C459 source.t40 a_n2354_n2088# 0.150063f
C460 source.t46 a_n2354_n2088# 0.150063f
C461 source.n258 a_n2354_n2088# 1.16869f
C462 source.n259 a_n2354_n2088# 0.407466f
C463 source.t35 a_n2354_n2088# 0.150063f
C464 source.t44 a_n2354_n2088# 0.150063f
C465 source.n260 a_n2354_n2088# 1.16869f
C466 source.n261 a_n2354_n2088# 0.407466f
C467 source.t8 a_n2354_n2088# 0.150063f
C468 source.t38 a_n2354_n2088# 0.150063f
C469 source.n262 a_n2354_n2088# 1.16869f
C470 source.n263 a_n2354_n2088# 0.407466f
C471 source.n264 a_n2354_n2088# 0.044486f
C472 source.n265 a_n2354_n2088# 0.03165f
C473 source.n266 a_n2354_n2088# 0.017007f
C474 source.n267 a_n2354_n2088# 0.040199f
C475 source.n268 a_n2354_n2088# 0.018008f
C476 source.n269 a_n2354_n2088# 0.03165f
C477 source.n270 a_n2354_n2088# 0.017007f
C478 source.n271 a_n2354_n2088# 0.040199f
C479 source.n272 a_n2354_n2088# 0.018008f
C480 source.n273 a_n2354_n2088# 0.135438f
C481 source.t4 a_n2354_n2088# 0.065518f
C482 source.n274 a_n2354_n2088# 0.030149f
C483 source.n275 a_n2354_n2088# 0.023745f
C484 source.n276 a_n2354_n2088# 0.017007f
C485 source.n277 a_n2354_n2088# 0.753071f
C486 source.n278 a_n2354_n2088# 0.03165f
C487 source.n279 a_n2354_n2088# 0.017007f
C488 source.n280 a_n2354_n2088# 0.018008f
C489 source.n281 a_n2354_n2088# 0.040199f
C490 source.n282 a_n2354_n2088# 0.040199f
C491 source.n283 a_n2354_n2088# 0.018008f
C492 source.n284 a_n2354_n2088# 0.017007f
C493 source.n285 a_n2354_n2088# 0.03165f
C494 source.n286 a_n2354_n2088# 0.03165f
C495 source.n287 a_n2354_n2088# 0.017007f
C496 source.n288 a_n2354_n2088# 0.018008f
C497 source.n289 a_n2354_n2088# 0.040199f
C498 source.n290 a_n2354_n2088# 0.087023f
C499 source.n291 a_n2354_n2088# 0.018008f
C500 source.n292 a_n2354_n2088# 0.017007f
C501 source.n293 a_n2354_n2088# 0.073156f
C502 source.n294 a_n2354_n2088# 0.048693f
C503 source.n295 a_n2354_n2088# 0.308993f
C504 source.n296 a_n2354_n2088# 1.29504f
C505 drain_left.t4 a_n2354_n2088# 0.16016f
C506 drain_left.t2 a_n2354_n2088# 0.16016f
C507 drain_left.n0 a_n2354_n2088# 1.33899f
C508 drain_left.t14 a_n2354_n2088# 0.16016f
C509 drain_left.t16 a_n2354_n2088# 0.16016f
C510 drain_left.n1 a_n2354_n2088# 1.33574f
C511 drain_left.n2 a_n2354_n2088# 0.795133f
C512 drain_left.t13 a_n2354_n2088# 0.16016f
C513 drain_left.t18 a_n2354_n2088# 0.16016f
C514 drain_left.n3 a_n2354_n2088# 1.33574f
C515 drain_left.n4 a_n2354_n2088# 0.360432f
C516 drain_left.t3 a_n2354_n2088# 0.16016f
C517 drain_left.t8 a_n2354_n2088# 0.16016f
C518 drain_left.n5 a_n2354_n2088# 1.33899f
C519 drain_left.t22 a_n2354_n2088# 0.16016f
C520 drain_left.t11 a_n2354_n2088# 0.16016f
C521 drain_left.n6 a_n2354_n2088# 1.33574f
C522 drain_left.n7 a_n2354_n2088# 0.795133f
C523 drain_left.t20 a_n2354_n2088# 0.16016f
C524 drain_left.t21 a_n2354_n2088# 0.16016f
C525 drain_left.n8 a_n2354_n2088# 1.33574f
C526 drain_left.n9 a_n2354_n2088# 0.360432f
C527 drain_left.n10 a_n2354_n2088# 1.38899f
C528 drain_left.t15 a_n2354_n2088# 0.16016f
C529 drain_left.t5 a_n2354_n2088# 0.16016f
C530 drain_left.n11 a_n2354_n2088# 1.339f
C531 drain_left.t9 a_n2354_n2088# 0.16016f
C532 drain_left.t10 a_n2354_n2088# 0.16016f
C533 drain_left.n12 a_n2354_n2088# 1.33574f
C534 drain_left.n13 a_n2354_n2088# 0.79512f
C535 drain_left.t23 a_n2354_n2088# 0.16016f
C536 drain_left.t6 a_n2354_n2088# 0.16016f
C537 drain_left.n14 a_n2354_n2088# 1.33574f
C538 drain_left.n15 a_n2354_n2088# 0.392385f
C539 drain_left.t7 a_n2354_n2088# 0.16016f
C540 drain_left.t0 a_n2354_n2088# 0.16016f
C541 drain_left.n16 a_n2354_n2088# 1.33574f
C542 drain_left.n17 a_n2354_n2088# 0.392385f
C543 drain_left.t17 a_n2354_n2088# 0.16016f
C544 drain_left.t12 a_n2354_n2088# 0.16016f
C545 drain_left.n18 a_n2354_n2088# 1.33574f
C546 drain_left.n19 a_n2354_n2088# 0.392385f
C547 drain_left.t1 a_n2354_n2088# 0.16016f
C548 drain_left.t19 a_n2354_n2088# 0.16016f
C549 drain_left.n20 a_n2354_n2088# 1.33574f
C550 drain_left.n21 a_n2354_n2088# 0.673556f
C551 plus.n0 a_n2354_n2088# 0.049758f
C552 plus.t0 a_n2354_n2088# 0.255186f
C553 plus.t19 a_n2354_n2088# 0.255186f
C554 plus.n1 a_n2354_n2088# 0.117134f
C555 plus.n2 a_n2354_n2088# 0.049758f
C556 plus.t14 a_n2354_n2088# 0.255186f
C557 plus.t1 a_n2354_n2088# 0.255186f
C558 plus.t22 a_n2354_n2088# 0.255186f
C559 plus.n3 a_n2354_n2088# 0.117134f
C560 plus.n4 a_n2354_n2088# 0.049758f
C561 plus.t15 a_n2354_n2088# 0.255186f
C562 plus.t10 a_n2354_n2088# 0.255186f
C563 plus.n5 a_n2354_n2088# 0.117134f
C564 plus.n6 a_n2354_n2088# 0.049758f
C565 plus.t23 a_n2354_n2088# 0.255186f
C566 plus.t16 a_n2354_n2088# 0.255186f
C567 plus.n7 a_n2354_n2088# 0.019114f
C568 plus.t4 a_n2354_n2088# 0.261163f
C569 plus.t11 a_n2354_n2088# 0.255186f
C570 plus.n8 a_n2354_n2088# 0.117134f
C571 plus.n9 a_n2354_n2088# 0.132179f
C572 plus.n10 a_n2354_n2088# 0.106506f
C573 plus.n11 a_n2354_n2088# 0.049758f
C574 plus.n12 a_n2354_n2088# 0.017887f
C575 plus.n13 a_n2354_n2088# 0.117134f
C576 plus.n14 a_n2354_n2088# 0.020495f
C577 plus.n15 a_n2354_n2088# 0.117134f
C578 plus.n16 a_n2354_n2088# 0.020495f
C579 plus.n17 a_n2354_n2088# 0.049758f
C580 plus.n18 a_n2354_n2088# 0.049758f
C581 plus.n19 a_n2354_n2088# 0.020495f
C582 plus.n20 a_n2354_n2088# 0.117134f
C583 plus.n21 a_n2354_n2088# 0.0185f
C584 plus.n22 a_n2354_n2088# 0.0185f
C585 plus.n23 a_n2354_n2088# 0.049758f
C586 plus.n24 a_n2354_n2088# 0.049758f
C587 plus.n25 a_n2354_n2088# 0.020495f
C588 plus.n26 a_n2354_n2088# 0.117134f
C589 plus.n27 a_n2354_n2088# 0.020495f
C590 plus.n28 a_n2354_n2088# 0.117134f
C591 plus.n29 a_n2354_n2088# 0.020495f
C592 plus.n30 a_n2354_n2088# 0.049758f
C593 plus.n31 a_n2354_n2088# 0.049758f
C594 plus.n32 a_n2354_n2088# 0.017887f
C595 plus.n33 a_n2354_n2088# 0.019114f
C596 plus.n34 a_n2354_n2088# 0.117134f
C597 plus.t7 a_n2354_n2088# 0.261163f
C598 plus.n35 a_n2354_n2088# 0.132112f
C599 plus.n36 a_n2354_n2088# 0.422727f
C600 plus.n37 a_n2354_n2088# 0.049758f
C601 plus.t17 a_n2354_n2088# 0.261163f
C602 plus.t2 a_n2354_n2088# 0.255186f
C603 plus.t9 a_n2354_n2088# 0.255186f
C604 plus.n38 a_n2354_n2088# 0.117134f
C605 plus.n39 a_n2354_n2088# 0.049758f
C606 plus.t18 a_n2354_n2088# 0.255186f
C607 plus.t8 a_n2354_n2088# 0.255186f
C608 plus.t21 a_n2354_n2088# 0.255186f
C609 plus.n40 a_n2354_n2088# 0.117134f
C610 plus.n41 a_n2354_n2088# 0.049758f
C611 plus.t6 a_n2354_n2088# 0.255186f
C612 plus.t20 a_n2354_n2088# 0.255186f
C613 plus.n42 a_n2354_n2088# 0.117134f
C614 plus.n43 a_n2354_n2088# 0.049758f
C615 plus.t5 a_n2354_n2088# 0.255186f
C616 plus.t13 a_n2354_n2088# 0.255186f
C617 plus.n44 a_n2354_n2088# 0.019114f
C618 plus.t3 a_n2354_n2088# 0.255186f
C619 plus.n45 a_n2354_n2088# 0.117134f
C620 plus.t12 a_n2354_n2088# 0.261163f
C621 plus.n46 a_n2354_n2088# 0.132179f
C622 plus.n47 a_n2354_n2088# 0.106506f
C623 plus.n48 a_n2354_n2088# 0.049758f
C624 plus.n49 a_n2354_n2088# 0.017887f
C625 plus.n50 a_n2354_n2088# 0.117134f
C626 plus.n51 a_n2354_n2088# 0.020495f
C627 plus.n52 a_n2354_n2088# 0.117134f
C628 plus.n53 a_n2354_n2088# 0.020495f
C629 plus.n54 a_n2354_n2088# 0.049758f
C630 plus.n55 a_n2354_n2088# 0.049758f
C631 plus.n56 a_n2354_n2088# 0.020495f
C632 plus.n57 a_n2354_n2088# 0.117134f
C633 plus.n58 a_n2354_n2088# 0.0185f
C634 plus.n59 a_n2354_n2088# 0.0185f
C635 plus.n60 a_n2354_n2088# 0.049758f
C636 plus.n61 a_n2354_n2088# 0.049758f
C637 plus.n62 a_n2354_n2088# 0.020495f
C638 plus.n63 a_n2354_n2088# 0.117134f
C639 plus.n64 a_n2354_n2088# 0.020495f
C640 plus.n65 a_n2354_n2088# 0.117134f
C641 plus.n66 a_n2354_n2088# 0.020495f
C642 plus.n67 a_n2354_n2088# 0.049758f
C643 plus.n68 a_n2354_n2088# 0.049758f
C644 plus.n69 a_n2354_n2088# 0.017887f
C645 plus.n70 a_n2354_n2088# 0.019114f
C646 plus.n71 a_n2354_n2088# 0.117134f
C647 plus.n72 a_n2354_n2088# 0.132112f
C648 plus.n73 a_n2354_n2088# 1.40167f
.ends

