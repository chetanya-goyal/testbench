* NGSPICE file created from diffpair407.ext - technology: sky130A

.subckt diffpair407 minus drain_right drain_left source plus
X0 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X1 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X2 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X3 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X4 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X5 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X6 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X7 a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X8 a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X9 a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X10 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X11 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X12 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X14 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X15 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X16 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X18 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X20 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X21 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X22 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X23 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X24 a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X25 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X26 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X27 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X28 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X29 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X30 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X31 source minus drain_right a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X32 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X33 drain_left plus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X34 source plus drain_left a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X35 drain_right minus source a_n1886_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
.ends

