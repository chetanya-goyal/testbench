* NGSPICE file created from diffpair605.ext - technology: sky130A

.subckt diffpair605 minus drain_right drain_left source plus
X0 a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X1 drain_left.t11 plus.t0 source.t19 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X2 source.t18 plus.t1 drain_left.t10 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X3 source.t3 minus.t0 drain_right.t11 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X4 source.t17 plus.t2 drain_left.t9 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X5 drain_left.t8 plus.t3 source.t14 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t15 plus.t4 drain_left.t7 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X7 drain_right.t10 minus.t1 source.t2 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 source.t7 minus.t2 drain_right.t9 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X9 drain_right.t8 minus.t3 source.t1 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X11 drain_right.t7 minus.t4 source.t6 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X12 source.t22 minus.t5 drain_right.t6 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X13 drain_left.t6 plus.t5 source.t20 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X14 drain_left.t5 plus.t6 source.t9 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 source.t21 minus.t6 drain_right.t5 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X16 a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X17 source.t11 plus.t7 drain_left.t4 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X18 drain_right.t4 minus.t7 source.t8 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 drain_right.t3 minus.t8 source.t0 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X20 source.t23 minus.t9 drain_right.t2 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X21 a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X22 drain_left.t3 plus.t8 source.t13 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 drain_right.t1 minus.t10 source.t5 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X24 source.t4 minus.t11 drain_right.t0 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X25 source.t16 plus.t9 drain_left.t2 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X26 source.t10 plus.t10 drain_left.t1 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X27 drain_left.t0 plus.t11 source.t12 a_n1878_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
R0 plus.n5 plus.t4 1069.23
R1 plus.n19 plus.t0 1069.23
R2 plus.n12 plus.t11 1042.57
R3 plus.n10 plus.t9 1042.57
R4 plus.n9 plus.t5 1042.57
R5 plus.n3 plus.t10 1042.57
R6 plus.n4 plus.t8 1042.57
R7 plus.n26 plus.t7 1042.57
R8 plus.n24 plus.t3 1042.57
R9 plus.n23 plus.t2 1042.57
R10 plus.n17 plus.t6 1042.57
R11 plus.n18 plus.t1 1042.57
R12 plus.n6 plus.n3 161.3
R13 plus.n8 plus.n7 161.3
R14 plus.n9 plus.n2 161.3
R15 plus.n10 plus.n1 161.3
R16 plus.n11 plus.n0 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n20 plus.n17 161.3
R19 plus.n22 plus.n21 161.3
R20 plus.n23 plus.n16 161.3
R21 plus.n24 plus.n15 161.3
R22 plus.n25 plus.n14 161.3
R23 plus.n27 plus.n26 161.3
R24 plus.n10 plus.n9 48.2005
R25 plus.n4 plus.n3 48.2005
R26 plus.n24 plus.n23 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n12 plus.n11 47.4702
R29 plus.n26 plus.n25 47.4702
R30 plus.n6 plus.n5 45.1192
R31 plus.n20 plus.n19 45.1192
R32 plus plus.n27 33.1771
R33 plus.n8 plus.n3 24.1005
R34 plus.n9 plus.n8 24.1005
R35 plus.n23 plus.n22 24.1005
R36 plus.n22 plus.n17 24.1005
R37 plus plus.n13 15.205
R38 plus.n5 plus.n4 13.6377
R39 plus.n19 plus.n18 13.6377
R40 plus.n11 plus.n10 0.730803
R41 plus.n25 plus.n24 0.730803
R42 plus.n7 plus.n6 0.189894
R43 plus.n7 plus.n2 0.189894
R44 plus.n2 plus.n1 0.189894
R45 plus.n1 plus.n0 0.189894
R46 plus.n13 plus.n0 0.189894
R47 plus.n27 plus.n14 0.189894
R48 plus.n15 plus.n14 0.189894
R49 plus.n16 plus.n15 0.189894
R50 plus.n21 plus.n16 0.189894
R51 plus.n21 plus.n20 0.189894
R52 source.n0 source.t12 44.1297
R53 source.n5 source.t15 44.1296
R54 source.n6 source.t0 44.1296
R55 source.n11 source.t21 44.1296
R56 source.n23 source.t5 44.1295
R57 source.n18 source.t7 44.1295
R58 source.n17 source.t19 44.1295
R59 source.n12 source.t11 44.1295
R60 source.n2 source.n1 43.1397
R61 source.n4 source.n3 43.1397
R62 source.n8 source.n7 43.1397
R63 source.n10 source.n9 43.1397
R64 source.n22 source.n21 43.1396
R65 source.n20 source.n19 43.1396
R66 source.n16 source.n15 43.1396
R67 source.n14 source.n13 43.1396
R68 source.n12 source.n11 28.0638
R69 source.n24 source.n0 22.4432
R70 source.n24 source.n23 5.62119
R71 source.n21 source.t8 0.9905
R72 source.n21 source.t22 0.9905
R73 source.n19 source.t2 0.9905
R74 source.n19 source.t23 0.9905
R75 source.n15 source.t9 0.9905
R76 source.n15 source.t18 0.9905
R77 source.n13 source.t14 0.9905
R78 source.n13 source.t17 0.9905
R79 source.n1 source.t20 0.9905
R80 source.n1 source.t16 0.9905
R81 source.n3 source.t13 0.9905
R82 source.n3 source.t10 0.9905
R83 source.n7 source.t6 0.9905
R84 source.n7 source.t3 0.9905
R85 source.n9 source.t1 0.9905
R86 source.n9 source.t4 0.9905
R87 source.n11 source.n10 0.716017
R88 source.n10 source.n8 0.716017
R89 source.n8 source.n6 0.716017
R90 source.n5 source.n4 0.716017
R91 source.n4 source.n2 0.716017
R92 source.n2 source.n0 0.716017
R93 source.n14 source.n12 0.716017
R94 source.n16 source.n14 0.716017
R95 source.n17 source.n16 0.716017
R96 source.n20 source.n18 0.716017
R97 source.n22 source.n20 0.716017
R98 source.n23 source.n22 0.716017
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 60.534
R103 drain_left.n3 drain_left.n2 60.4786
R104 drain_left.n3 drain_left.n0 60.4786
R105 drain_left.n8 drain_left.n7 59.8185
R106 drain_left.n6 drain_left.n5 59.8185
R107 drain_left.n3 drain_left.n1 59.8184
R108 drain_left drain_left.n3 37.0053
R109 drain_left drain_left.n8 6.36873
R110 drain_left.n1 drain_left.t9 0.9905
R111 drain_left.n1 drain_left.t5 0.9905
R112 drain_left.n2 drain_left.t10 0.9905
R113 drain_left.n2 drain_left.t11 0.9905
R114 drain_left.n0 drain_left.t4 0.9905
R115 drain_left.n0 drain_left.t8 0.9905
R116 drain_left.n7 drain_left.t2 0.9905
R117 drain_left.n7 drain_left.t0 0.9905
R118 drain_left.n5 drain_left.t1 0.9905
R119 drain_left.n5 drain_left.t6 0.9905
R120 drain_left.n4 drain_left.t7 0.9905
R121 drain_left.n4 drain_left.t3 0.9905
R122 drain_left.n8 drain_left.n6 0.716017
R123 minus.n3 minus.t8 1069.23
R124 minus.n17 minus.t2 1069.23
R125 minus.n4 minus.t0 1042.57
R126 minus.n5 minus.t4 1042.57
R127 minus.n1 minus.t11 1042.57
R128 minus.n10 minus.t3 1042.57
R129 minus.n12 minus.t6 1042.57
R130 minus.n18 minus.t1 1042.57
R131 minus.n19 minus.t9 1042.57
R132 minus.n15 minus.t7 1042.57
R133 minus.n24 minus.t5 1042.57
R134 minus.n26 minus.t10 1042.57
R135 minus.n13 minus.n12 161.3
R136 minus.n11 minus.n0 161.3
R137 minus.n10 minus.n9 161.3
R138 minus.n8 minus.n1 161.3
R139 minus.n7 minus.n6 161.3
R140 minus.n5 minus.n2 161.3
R141 minus.n27 minus.n26 161.3
R142 minus.n25 minus.n14 161.3
R143 minus.n24 minus.n23 161.3
R144 minus.n22 minus.n15 161.3
R145 minus.n21 minus.n20 161.3
R146 minus.n19 minus.n16 161.3
R147 minus.n5 minus.n4 48.2005
R148 minus.n10 minus.n1 48.2005
R149 minus.n19 minus.n18 48.2005
R150 minus.n24 minus.n15 48.2005
R151 minus.n12 minus.n11 47.4702
R152 minus.n26 minus.n25 47.4702
R153 minus.n3 minus.n2 45.1192
R154 minus.n17 minus.n16 45.1192
R155 minus.n28 minus.n13 42.3263
R156 minus.n6 minus.n1 24.1005
R157 minus.n6 minus.n5 24.1005
R158 minus.n20 minus.n19 24.1005
R159 minus.n20 minus.n15 24.1005
R160 minus.n4 minus.n3 13.6377
R161 minus.n18 minus.n17 13.6377
R162 minus.n28 minus.n27 6.5308
R163 minus.n11 minus.n10 0.730803
R164 minus.n25 minus.n24 0.730803
R165 minus.n13 minus.n0 0.189894
R166 minus.n9 minus.n0 0.189894
R167 minus.n9 minus.n8 0.189894
R168 minus.n8 minus.n7 0.189894
R169 minus.n7 minus.n2 0.189894
R170 minus.n21 minus.n16 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n14 0.189894
R174 minus.n27 minus.n14 0.189894
R175 minus minus.n28 0.188
R176 drain_right.n6 drain_right.n4 60.534
R177 drain_right.n3 drain_right.n2 60.4786
R178 drain_right.n3 drain_right.n0 60.4786
R179 drain_right.n6 drain_right.n5 59.8185
R180 drain_right.n8 drain_right.n7 59.8185
R181 drain_right.n3 drain_right.n1 59.8184
R182 drain_right drain_right.n3 36.452
R183 drain_right drain_right.n8 6.36873
R184 drain_right.n1 drain_right.t2 0.9905
R185 drain_right.n1 drain_right.t4 0.9905
R186 drain_right.n2 drain_right.t6 0.9905
R187 drain_right.n2 drain_right.t1 0.9905
R188 drain_right.n0 drain_right.t9 0.9905
R189 drain_right.n0 drain_right.t10 0.9905
R190 drain_right.n4 drain_right.t11 0.9905
R191 drain_right.n4 drain_right.t3 0.9905
R192 drain_right.n5 drain_right.t0 0.9905
R193 drain_right.n5 drain_right.t7 0.9905
R194 drain_right.n7 drain_right.t5 0.9905
R195 drain_right.n7 drain_right.t8 0.9905
R196 drain_right.n8 drain_right.n6 0.716017
C0 source drain_left 28.8063f
C1 drain_left plus 10.6735f
C2 source plus 9.95609f
C3 drain_right minus 10.4909f
C4 drain_right drain_left 0.936346f
C5 drain_right source 28.807299f
C6 minus drain_left 0.171641f
C7 minus source 9.94205f
C8 drain_right plus 0.337327f
C9 minus plus 6.97471f
C10 drain_right a_n1878_n4888# 7.63563f
C11 drain_left a_n1878_n4888# 7.91663f
C12 source a_n1878_n4888# 13.317128f
C13 minus a_n1878_n4888# 7.900587f
C14 plus a_n1878_n4888# 10.20076f
C15 drain_right.t9 a_n1878_n4888# 0.464323f
C16 drain_right.t10 a_n1878_n4888# 0.464323f
C17 drain_right.n0 a_n1878_n4888# 4.24921f
C18 drain_right.t2 a_n1878_n4888# 0.464323f
C19 drain_right.t4 a_n1878_n4888# 0.464323f
C20 drain_right.n1 a_n1878_n4888# 4.24494f
C21 drain_right.t6 a_n1878_n4888# 0.464323f
C22 drain_right.t1 a_n1878_n4888# 0.464323f
C23 drain_right.n2 a_n1878_n4888# 4.24921f
C24 drain_right.n3 a_n1878_n4888# 3.07041f
C25 drain_right.t11 a_n1878_n4888# 0.464323f
C26 drain_right.t3 a_n1878_n4888# 0.464323f
C27 drain_right.n4 a_n1878_n4888# 4.24961f
C28 drain_right.t0 a_n1878_n4888# 0.464323f
C29 drain_right.t7 a_n1878_n4888# 0.464323f
C30 drain_right.n5 a_n1878_n4888# 4.24494f
C31 drain_right.n6 a_n1878_n4888# 0.773945f
C32 drain_right.t5 a_n1878_n4888# 0.464323f
C33 drain_right.t8 a_n1878_n4888# 0.464323f
C34 drain_right.n7 a_n1878_n4888# 4.24494f
C35 drain_right.n8 a_n1878_n4888# 0.635798f
C36 minus.n0 a_n1878_n4888# 0.046365f
C37 minus.t11 a_n1878_n4888# 1.313f
C38 minus.n1 a_n1878_n4888# 0.497949f
C39 minus.t3 a_n1878_n4888# 1.313f
C40 minus.n2 a_n1878_n4888# 0.188827f
C41 minus.t8 a_n1878_n4888# 1.3253f
C42 minus.n3 a_n1878_n4888# 0.482065f
C43 minus.t0 a_n1878_n4888# 1.313f
C44 minus.n4 a_n1878_n4888# 0.503538f
C45 minus.t4 a_n1878_n4888# 1.313f
C46 minus.n5 a_n1878_n4888# 0.497949f
C47 minus.n6 a_n1878_n4888# 0.010521f
C48 minus.n7 a_n1878_n4888# 0.046365f
C49 minus.n8 a_n1878_n4888# 0.046365f
C50 minus.n9 a_n1878_n4888# 0.046365f
C51 minus.n10 a_n1878_n4888# 0.493375f
C52 minus.n11 a_n1878_n4888# 0.010521f
C53 minus.t6 a_n1878_n4888# 1.313f
C54 minus.n12 a_n1878_n4888# 0.493089f
C55 minus.n13 a_n1878_n4888# 2.07777f
C56 minus.n14 a_n1878_n4888# 0.046365f
C57 minus.t7 a_n1878_n4888# 1.313f
C58 minus.n15 a_n1878_n4888# 0.497949f
C59 minus.n16 a_n1878_n4888# 0.188827f
C60 minus.t2 a_n1878_n4888# 1.3253f
C61 minus.n17 a_n1878_n4888# 0.482065f
C62 minus.t1 a_n1878_n4888# 1.313f
C63 minus.n18 a_n1878_n4888# 0.503538f
C64 minus.t9 a_n1878_n4888# 1.313f
C65 minus.n19 a_n1878_n4888# 0.497949f
C66 minus.n20 a_n1878_n4888# 0.010521f
C67 minus.n21 a_n1878_n4888# 0.046365f
C68 minus.n22 a_n1878_n4888# 0.046365f
C69 minus.n23 a_n1878_n4888# 0.046365f
C70 minus.t5 a_n1878_n4888# 1.313f
C71 minus.n24 a_n1878_n4888# 0.493375f
C72 minus.n25 a_n1878_n4888# 0.010521f
C73 minus.t10 a_n1878_n4888# 1.313f
C74 minus.n26 a_n1878_n4888# 0.493089f
C75 minus.n27 a_n1878_n4888# 0.306481f
C76 minus.n28 a_n1878_n4888# 2.4781f
C77 drain_left.t4 a_n1878_n4888# 0.465325f
C78 drain_left.t8 a_n1878_n4888# 0.465325f
C79 drain_left.n0 a_n1878_n4888# 4.25838f
C80 drain_left.t9 a_n1878_n4888# 0.465325f
C81 drain_left.t5 a_n1878_n4888# 0.465325f
C82 drain_left.n1 a_n1878_n4888# 4.2541f
C83 drain_left.t10 a_n1878_n4888# 0.465325f
C84 drain_left.t11 a_n1878_n4888# 0.465325f
C85 drain_left.n2 a_n1878_n4888# 4.25838f
C86 drain_left.n3 a_n1878_n4888# 3.1383f
C87 drain_left.t7 a_n1878_n4888# 0.465325f
C88 drain_left.t3 a_n1878_n4888# 0.465325f
C89 drain_left.n4 a_n1878_n4888# 4.25878f
C90 drain_left.t1 a_n1878_n4888# 0.465325f
C91 drain_left.t6 a_n1878_n4888# 0.465325f
C92 drain_left.n5 a_n1878_n4888# 4.2541f
C93 drain_left.n6 a_n1878_n4888# 0.775616f
C94 drain_left.t2 a_n1878_n4888# 0.465325f
C95 drain_left.t0 a_n1878_n4888# 0.465325f
C96 drain_left.n7 a_n1878_n4888# 4.2541f
C97 drain_left.n8 a_n1878_n4888# 0.63717f
C98 source.t12 a_n1878_n4888# 4.11252f
C99 source.n0 a_n1878_n4888# 1.76913f
C100 source.t20 a_n1878_n4888# 0.359852f
C101 source.t16 a_n1878_n4888# 0.359852f
C102 source.n1 a_n1878_n4888# 3.21723f
C103 source.n2 a_n1878_n4888# 0.338793f
C104 source.t13 a_n1878_n4888# 0.359852f
C105 source.t10 a_n1878_n4888# 0.359852f
C106 source.n3 a_n1878_n4888# 3.21723f
C107 source.n4 a_n1878_n4888# 0.338793f
C108 source.t15 a_n1878_n4888# 4.11253f
C109 source.n5 a_n1878_n4888# 0.406879f
C110 source.t0 a_n1878_n4888# 4.11253f
C111 source.n6 a_n1878_n4888# 0.406879f
C112 source.t6 a_n1878_n4888# 0.359852f
C113 source.t3 a_n1878_n4888# 0.359852f
C114 source.n7 a_n1878_n4888# 3.21723f
C115 source.n8 a_n1878_n4888# 0.338793f
C116 source.t1 a_n1878_n4888# 0.359852f
C117 source.t4 a_n1878_n4888# 0.359852f
C118 source.n9 a_n1878_n4888# 3.21723f
C119 source.n10 a_n1878_n4888# 0.338793f
C120 source.t21 a_n1878_n4888# 4.11253f
C121 source.n11 a_n1878_n4888# 2.17798f
C122 source.t11 a_n1878_n4888# 4.11251f
C123 source.n12 a_n1878_n4888# 2.178f
C124 source.t14 a_n1878_n4888# 0.359852f
C125 source.t17 a_n1878_n4888# 0.359852f
C126 source.n13 a_n1878_n4888# 3.21723f
C127 source.n14 a_n1878_n4888# 0.338787f
C128 source.t9 a_n1878_n4888# 0.359852f
C129 source.t18 a_n1878_n4888# 0.359852f
C130 source.n15 a_n1878_n4888# 3.21723f
C131 source.n16 a_n1878_n4888# 0.338787f
C132 source.t19 a_n1878_n4888# 4.11251f
C133 source.n17 a_n1878_n4888# 0.406902f
C134 source.t7 a_n1878_n4888# 4.11251f
C135 source.n18 a_n1878_n4888# 0.406902f
C136 source.t2 a_n1878_n4888# 0.359852f
C137 source.t23 a_n1878_n4888# 0.359852f
C138 source.n19 a_n1878_n4888# 3.21723f
C139 source.n20 a_n1878_n4888# 0.338787f
C140 source.t8 a_n1878_n4888# 0.359852f
C141 source.t22 a_n1878_n4888# 0.359852f
C142 source.n21 a_n1878_n4888# 3.21723f
C143 source.n22 a_n1878_n4888# 0.338787f
C144 source.t5 a_n1878_n4888# 4.11251f
C145 source.n23 a_n1878_n4888# 0.545484f
C146 source.n24 a_n1878_n4888# 2.05757f
C147 plus.n0 a_n1878_n4888# 0.047033f
C148 plus.t11 a_n1878_n4888# 1.33193f
C149 plus.t9 a_n1878_n4888# 1.33193f
C150 plus.n1 a_n1878_n4888# 0.047033f
C151 plus.t5 a_n1878_n4888# 1.33193f
C152 plus.n2 a_n1878_n4888# 0.047033f
C153 plus.t10 a_n1878_n4888# 1.33193f
C154 plus.n3 a_n1878_n4888# 0.50513f
C155 plus.t8 a_n1878_n4888# 1.33193f
C156 plus.n4 a_n1878_n4888# 0.510799f
C157 plus.t4 a_n1878_n4888# 1.34442f
C158 plus.n5 a_n1878_n4888# 0.489017f
C159 plus.n6 a_n1878_n4888# 0.19155f
C160 plus.n7 a_n1878_n4888# 0.047033f
C161 plus.n8 a_n1878_n4888# 0.010673f
C162 plus.n9 a_n1878_n4888# 0.50513f
C163 plus.n10 a_n1878_n4888# 0.50049f
C164 plus.n11 a_n1878_n4888# 0.010673f
C165 plus.n12 a_n1878_n4888# 0.5002f
C166 plus.n13 a_n1878_n4888# 0.7175f
C167 plus.n14 a_n1878_n4888# 0.047033f
C168 plus.t7 a_n1878_n4888# 1.33193f
C169 plus.n15 a_n1878_n4888# 0.047033f
C170 plus.t3 a_n1878_n4888# 1.33193f
C171 plus.n16 a_n1878_n4888# 0.047033f
C172 plus.t2 a_n1878_n4888# 1.33193f
C173 plus.t6 a_n1878_n4888# 1.33193f
C174 plus.n17 a_n1878_n4888# 0.50513f
C175 plus.t0 a_n1878_n4888# 1.34442f
C176 plus.t1 a_n1878_n4888# 1.33193f
C177 plus.n18 a_n1878_n4888# 0.510799f
C178 plus.n19 a_n1878_n4888# 0.489017f
C179 plus.n20 a_n1878_n4888# 0.19155f
C180 plus.n21 a_n1878_n4888# 0.047033f
C181 plus.n22 a_n1878_n4888# 0.010673f
C182 plus.n23 a_n1878_n4888# 0.50513f
C183 plus.n24 a_n1878_n4888# 0.50049f
C184 plus.n25 a_n1878_n4888# 0.010673f
C185 plus.n26 a_n1878_n4888# 0.5002f
C186 plus.n27 a_n1878_n4888# 1.66854f
.ends

