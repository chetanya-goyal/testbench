* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.2
X1 a_n928_n1092# a_n928_n1092# a_n928_n1092# a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.2
X2 a_n928_n1092# a_n928_n1092# a_n928_n1092# a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X3 a_n928_n1092# a_n928_n1092# a_n928_n1092# a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X4 a_n928_n1092# a_n928_n1092# a_n928_n1092# a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X5 drain_left.t1 plus.t0 source.t0 a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.2
X6 drain_right.t0 minus.t1 source.t3 a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.2
X7 drain_left.t0 plus.t1 source.t1 a_n928_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.2
R0 minus.n0 minus.t0 486.7
R1 minus.n0 minus.t1 468.882
R2 minus minus.n0 0.188
R3 source.n0 source.t0 243.255
R4 source.n1 source.t2 243.255
R5 source.n3 source.t3 243.254
R6 source.n2 source.t1 243.254
R7 source.n2 source.n1 13.8833
R8 source.n4 source.n0 7.93506
R9 source.n4 source.n3 5.49188
R10 source.n1 source.n0 0.698776
R11 source.n3 source.n2 0.698776
R12 source source.n4 0.188
R13 drain_right drain_right.t0 279.058
R14 drain_right drain_right.t1 265.815
R15 plus plus.t1 484.748
R16 plus plus.t0 470.36
R17 drain_left drain_left.t0 279.611
R18 drain_left drain_left.t1 266.043
C0 drain_right plus 0.246532f
C1 source drain_left 1.69177f
C2 source minus 0.359719f
C3 drain_left minus 0.178971f
C4 source plus 0.37364f
C5 drain_right source 1.69098f
C6 drain_left plus 0.405547f
C7 drain_right drain_left 0.417605f
C8 minus plus 2.29562f
C9 drain_right minus 0.322041f
C10 drain_right a_n928_n1092# 1.51996f
C11 drain_left a_n928_n1092# 1.61303f
C12 source a_n928_n1092# 1.62037f
C13 minus a_n928_n1092# 2.71731f
C14 plus a_n928_n1092# 4.70505f
C15 plus.t0 a_n928_n1092# 0.052412f
C16 plus.t1 a_n928_n1092# 0.086621f
C17 minus.t0 a_n928_n1092# 0.086705f
C18 minus.t1 a_n928_n1092# 0.049025f
C19 minus.n0 a_n928_n1092# 2.1331f
.ends

