* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t20 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 drain_left.t19 plus.t0 source.t4 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 source.t28 minus.t1 drain_right.t18 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X3 source.t3 plus.t1 drain_left.t18 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 drain_right.t17 minus.t2 source.t19 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X5 source.t5 plus.t2 drain_left.t17 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X6 drain_right.t16 minus.t3 source.t21 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X7 a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X8 source.t22 minus.t4 drain_right.t15 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X9 source.t2 plus.t3 drain_left.t16 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X10 drain_left.t15 plus.t4 source.t1 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X11 drain_right.t14 minus.t5 source.t13 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X12 source.t23 minus.t6 drain_right.t13 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X14 drain_right.t12 minus.t7 source.t26 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X15 drain_right.t11 minus.t8 source.t27 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 source.t18 minus.t9 drain_right.t10 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X17 drain_left.t14 plus.t5 source.t0 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X18 source.t15 minus.t10 drain_right.t9 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X19 drain_right.t8 minus.t11 source.t10 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X20 source.t16 minus.t12 drain_right.t7 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X21 a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X22 drain_left.t13 plus.t6 source.t31 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X23 source.t39 plus.t7 drain_left.t12 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X24 drain_right.t6 minus.t13 source.t12 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X25 drain_right.t5 minus.t14 source.t11 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X26 source.t14 minus.t15 drain_right.t4 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X27 drain_right.t3 minus.t16 source.t17 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X28 source.t36 plus.t8 drain_left.t11 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X29 drain_left.t10 plus.t9 source.t30 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X30 source.t25 minus.t17 drain_right.t2 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X32 drain_left.t9 plus.t10 source.t9 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X33 drain_left.t8 plus.t11 source.t8 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X34 source.t37 plus.t12 drain_left.t7 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X35 source.t35 plus.t13 drain_left.t6 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X36 source.t24 minus.t18 drain_right.t1 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X37 source.t29 minus.t19 drain_right.t0 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X38 source.t33 plus.t14 drain_left.t5 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X39 drain_left.t4 plus.t15 source.t6 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X40 drain_left.t3 plus.t16 source.t7 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X41 drain_left.t2 plus.t17 source.t32 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X42 source.t38 plus.t18 drain_left.t1 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X43 source.t34 plus.t19 drain_left.t0 a_n2146_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
R0 minus.n27 minus.t18 431.61
R1 minus.n7 minus.t7 431.61
R2 minus.n56 minus.t16 431.61
R3 minus.n35 minus.t12 431.61
R4 minus.n26 minus.t11 369.534
R5 minus.n24 minus.t15 369.534
R6 minus.n3 minus.t14 369.534
R7 minus.n18 minus.t17 369.534
R8 minus.n16 minus.t8 369.534
R9 minus.n4 minus.t10 369.534
R10 minus.n10 minus.t13 369.534
R11 minus.n6 minus.t6 369.534
R12 minus.n55 minus.t19 369.534
R13 minus.n53 minus.t2 369.534
R14 minus.n47 minus.t4 369.534
R15 minus.n46 minus.t5 369.534
R16 minus.n44 minus.t9 369.534
R17 minus.n32 minus.t0 369.534
R18 minus.n38 minus.t1 369.534
R19 minus.n34 minus.t3 369.534
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 69.3793
R47 minus.n15 minus.n4 69.3793
R48 minus.n43 minus.n32 69.3793
R49 minus.n48 minus.n47 69.3793
R50 minus.n25 minus.n24 54.7732
R51 minus.n10 minus.n9 54.7732
R52 minus.n38 minus.n37 54.7732
R53 minus.n54 minus.n53 54.7732
R54 minus.n18 minus.n17 47.4702
R55 minus.n17 minus.n16 47.4702
R56 minus.n45 minus.n44 47.4702
R57 minus.n46 minus.n45 47.4702
R58 minus.n26 minus.n25 40.1672
R59 minus.n9 minus.n6 40.1672
R60 minus.n37 minus.n34 40.1672
R61 minus.n55 minus.n54 40.1672
R62 minus.n27 minus.n26 32.8641
R63 minus.n7 minus.n6 32.8641
R64 minus.n35 minus.n34 32.8641
R65 minus.n56 minus.n55 32.8641
R66 minus.n58 minus.n28 28.9778
R67 minus.n19 minus.n18 25.5611
R68 minus.n16 minus.n15 25.5611
R69 minus.n44 minus.n43 25.5611
R70 minus.n48 minus.n46 25.5611
R71 minus.n24 minus.n23 18.2581
R72 minus.n11 minus.n10 18.2581
R73 minus.n39 minus.n38 18.2581
R74 minus.n53 minus.n52 18.2581
R75 minus.n58 minus.n57 6.56111
R76 minus.n3 minus.n1 3.65202
R77 minus.n12 minus.n4 3.65202
R78 minus.n40 minus.n32 3.65202
R79 minus.n47 minus.n30 3.65202
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 source.n0 source.t8 253.454
R100 source.n9 source.t39 253.454
R101 source.n10 source.t26 253.454
R102 source.n19 source.t24 253.454
R103 source.n39 source.t17 253.453
R104 source.n30 source.t16 253.453
R105 source.n29 source.t1 253.453
R106 source.n20 source.t2 253.453
R107 source.n2 source.n1 223.454
R108 source.n4 source.n3 223.454
R109 source.n6 source.n5 223.454
R110 source.n8 source.n7 223.454
R111 source.n12 source.n11 223.454
R112 source.n14 source.n13 223.454
R113 source.n16 source.n15 223.454
R114 source.n18 source.n17 223.454
R115 source.n38 source.n37 223.453
R116 source.n36 source.n35 223.453
R117 source.n34 source.n33 223.453
R118 source.n32 source.n31 223.453
R119 source.n28 source.n27 223.453
R120 source.n26 source.n25 223.453
R121 source.n24 source.n23 223.453
R122 source.n22 source.n21 223.453
R123 source.n37 source.t19 30.0005
R124 source.n37 source.t29 30.0005
R125 source.n35 source.t13 30.0005
R126 source.n35 source.t22 30.0005
R127 source.n33 source.t20 30.0005
R128 source.n33 source.t18 30.0005
R129 source.n31 source.t21 30.0005
R130 source.n31 source.t28 30.0005
R131 source.n27 source.t32 30.0005
R132 source.n27 source.t5 30.0005
R133 source.n25 source.t0 30.0005
R134 source.n25 source.t36 30.0005
R135 source.n23 source.t4 30.0005
R136 source.n23 source.t3 30.0005
R137 source.n21 source.t9 30.0005
R138 source.n21 source.t38 30.0005
R139 source.n1 source.t31 30.0005
R140 source.n1 source.t33 30.0005
R141 source.n3 source.t6 30.0005
R142 source.n3 source.t37 30.0005
R143 source.n5 source.t30 30.0005
R144 source.n5 source.t34 30.0005
R145 source.n7 source.t7 30.0005
R146 source.n7 source.t35 30.0005
R147 source.n11 source.t12 30.0005
R148 source.n11 source.t23 30.0005
R149 source.n13 source.t27 30.0005
R150 source.n13 source.t15 30.0005
R151 source.n15 source.t11 30.0005
R152 source.n15 source.t25 30.0005
R153 source.n17 source.t10 30.0005
R154 source.n17 source.t14 30.0005
R155 source.n20 source.n19 13.5147
R156 source.n40 source.n0 7.97163
R157 source.n40 source.n39 5.5436
R158 source.n19 source.n18 0.560845
R159 source.n18 source.n16 0.560845
R160 source.n16 source.n14 0.560845
R161 source.n14 source.n12 0.560845
R162 source.n12 source.n10 0.560845
R163 source.n9 source.n8 0.560845
R164 source.n8 source.n6 0.560845
R165 source.n6 source.n4 0.560845
R166 source.n4 source.n2 0.560845
R167 source.n2 source.n0 0.560845
R168 source.n22 source.n20 0.560845
R169 source.n24 source.n22 0.560845
R170 source.n26 source.n24 0.560845
R171 source.n28 source.n26 0.560845
R172 source.n29 source.n28 0.560845
R173 source.n32 source.n30 0.560845
R174 source.n34 source.n32 0.560845
R175 source.n36 source.n34 0.560845
R176 source.n38 source.n36 0.560845
R177 source.n39 source.n38 0.560845
R178 source.n10 source.n9 0.470328
R179 source.n30 source.n29 0.470328
R180 source source.n40 0.188
R181 drain_right.n10 drain_right.n8 240.694
R182 drain_right.n6 drain_right.n4 240.692
R183 drain_right.n2 drain_right.n0 240.692
R184 drain_right.n10 drain_right.n9 240.132
R185 drain_right.n12 drain_right.n11 240.132
R186 drain_right.n14 drain_right.n13 240.132
R187 drain_right.n16 drain_right.n15 240.132
R188 drain_right.n7 drain_right.n3 240.131
R189 drain_right.n6 drain_right.n5 240.131
R190 drain_right.n2 drain_right.n1 240.131
R191 drain_right.n3 drain_right.t10 30.0005
R192 drain_right.n3 drain_right.t14 30.0005
R193 drain_right.n4 drain_right.t0 30.0005
R194 drain_right.n4 drain_right.t3 30.0005
R195 drain_right.n5 drain_right.t15 30.0005
R196 drain_right.n5 drain_right.t17 30.0005
R197 drain_right.n1 drain_right.t18 30.0005
R198 drain_right.n1 drain_right.t19 30.0005
R199 drain_right.n0 drain_right.t7 30.0005
R200 drain_right.n0 drain_right.t16 30.0005
R201 drain_right.n8 drain_right.t13 30.0005
R202 drain_right.n8 drain_right.t12 30.0005
R203 drain_right.n9 drain_right.t9 30.0005
R204 drain_right.n9 drain_right.t6 30.0005
R205 drain_right.n11 drain_right.t2 30.0005
R206 drain_right.n11 drain_right.t11 30.0005
R207 drain_right.n13 drain_right.t4 30.0005
R208 drain_right.n13 drain_right.t5 30.0005
R209 drain_right.n15 drain_right.t1 30.0005
R210 drain_right.n15 drain_right.t8 30.0005
R211 drain_right drain_right.n7 22.9633
R212 drain_right drain_right.n16 6.21356
R213 drain_right.n16 drain_right.n14 0.560845
R214 drain_right.n14 drain_right.n12 0.560845
R215 drain_right.n12 drain_right.n10 0.560845
R216 drain_right.n7 drain_right.n6 0.505499
R217 drain_right.n7 drain_right.n2 0.505499
R218 plus.n6 plus.t7 431.61
R219 plus.n27 plus.t11 431.61
R220 plus.n36 plus.t4 431.61
R221 plus.n56 plus.t3 431.61
R222 plus.n5 plus.t16 369.534
R223 plus.n9 plus.t13 369.534
R224 plus.n3 plus.t9 369.534
R225 plus.n15 plus.t19 369.534
R226 plus.n17 plus.t15 369.534
R227 plus.n18 plus.t12 369.534
R228 plus.n24 plus.t6 369.534
R229 plus.n26 plus.t14 369.534
R230 plus.n35 plus.t2 369.534
R231 plus.n39 plus.t17 369.534
R232 plus.n33 plus.t8 369.534
R233 plus.n45 plus.t5 369.534
R234 plus.n47 plus.t1 369.534
R235 plus.n32 plus.t0 369.534
R236 plus.n53 plus.t18 369.534
R237 plus.n55 plus.t10 369.534
R238 plus.n7 plus.n6 161.489
R239 plus.n37 plus.n36 161.489
R240 plus.n8 plus.n7 161.3
R241 plus.n10 plus.n4 161.3
R242 plus.n12 plus.n11 161.3
R243 plus.n14 plus.n13 161.3
R244 plus.n16 plus.n2 161.3
R245 plus.n20 plus.n19 161.3
R246 plus.n21 plus.n1 161.3
R247 plus.n23 plus.n22 161.3
R248 plus.n25 plus.n0 161.3
R249 plus.n28 plus.n27 161.3
R250 plus.n38 plus.n37 161.3
R251 plus.n40 plus.n34 161.3
R252 plus.n42 plus.n41 161.3
R253 plus.n44 plus.n43 161.3
R254 plus.n46 plus.n31 161.3
R255 plus.n49 plus.n48 161.3
R256 plus.n50 plus.n30 161.3
R257 plus.n52 plus.n51 161.3
R258 plus.n54 plus.n29 161.3
R259 plus.n57 plus.n56 161.3
R260 plus.n11 plus.n10 73.0308
R261 plus.n23 plus.n1 73.0308
R262 plus.n52 plus.n30 73.0308
R263 plus.n41 plus.n40 73.0308
R264 plus.n14 plus.n3 69.3793
R265 plus.n19 plus.n18 69.3793
R266 plus.n48 plus.n32 69.3793
R267 plus.n44 plus.n33 69.3793
R268 plus.n9 plus.n8 54.7732
R269 plus.n25 plus.n24 54.7732
R270 plus.n54 plus.n53 54.7732
R271 plus.n39 plus.n38 54.7732
R272 plus.n16 plus.n15 47.4702
R273 plus.n17 plus.n16 47.4702
R274 plus.n47 plus.n46 47.4702
R275 plus.n46 plus.n45 47.4702
R276 plus.n8 plus.n5 40.1672
R277 plus.n26 plus.n25 40.1672
R278 plus.n55 plus.n54 40.1672
R279 plus.n38 plus.n35 40.1672
R280 plus.n6 plus.n5 32.8641
R281 plus.n27 plus.n26 32.8641
R282 plus.n56 plus.n55 32.8641
R283 plus.n36 plus.n35 32.8641
R284 plus plus.n57 27.0255
R285 plus.n15 plus.n14 25.5611
R286 plus.n19 plus.n17 25.5611
R287 plus.n48 plus.n47 25.5611
R288 plus.n45 plus.n44 25.5611
R289 plus.n10 plus.n9 18.2581
R290 plus.n24 plus.n23 18.2581
R291 plus.n53 plus.n52 18.2581
R292 plus.n40 plus.n39 18.2581
R293 plus plus.n28 8.03838
R294 plus.n11 plus.n3 3.65202
R295 plus.n18 plus.n1 3.65202
R296 plus.n32 plus.n30 3.65202
R297 plus.n41 plus.n33 3.65202
R298 plus.n7 plus.n4 0.189894
R299 plus.n12 plus.n4 0.189894
R300 plus.n13 plus.n12 0.189894
R301 plus.n13 plus.n2 0.189894
R302 plus.n20 plus.n2 0.189894
R303 plus.n21 plus.n20 0.189894
R304 plus.n22 plus.n21 0.189894
R305 plus.n22 plus.n0 0.189894
R306 plus.n28 plus.n0 0.189894
R307 plus.n57 plus.n29 0.189894
R308 plus.n51 plus.n29 0.189894
R309 plus.n51 plus.n50 0.189894
R310 plus.n50 plus.n49 0.189894
R311 plus.n49 plus.n31 0.189894
R312 plus.n43 plus.n31 0.189894
R313 plus.n43 plus.n42 0.189894
R314 plus.n42 plus.n34 0.189894
R315 plus.n37 plus.n34 0.189894
R316 drain_left.n10 drain_left.n8 240.694
R317 drain_left.n6 drain_left.n4 240.692
R318 drain_left.n2 drain_left.n0 240.692
R319 drain_left.n16 drain_left.n15 240.132
R320 drain_left.n14 drain_left.n13 240.132
R321 drain_left.n12 drain_left.n11 240.132
R322 drain_left.n10 drain_left.n9 240.132
R323 drain_left.n7 drain_left.n3 240.131
R324 drain_left.n6 drain_left.n5 240.131
R325 drain_left.n2 drain_left.n1 240.131
R326 drain_left.n3 drain_left.t18 30.0005
R327 drain_left.n3 drain_left.t14 30.0005
R328 drain_left.n4 drain_left.t17 30.0005
R329 drain_left.n4 drain_left.t15 30.0005
R330 drain_left.n5 drain_left.t11 30.0005
R331 drain_left.n5 drain_left.t2 30.0005
R332 drain_left.n1 drain_left.t1 30.0005
R333 drain_left.n1 drain_left.t19 30.0005
R334 drain_left.n0 drain_left.t16 30.0005
R335 drain_left.n0 drain_left.t9 30.0005
R336 drain_left.n15 drain_left.t5 30.0005
R337 drain_left.n15 drain_left.t8 30.0005
R338 drain_left.n13 drain_left.t7 30.0005
R339 drain_left.n13 drain_left.t13 30.0005
R340 drain_left.n11 drain_left.t0 30.0005
R341 drain_left.n11 drain_left.t4 30.0005
R342 drain_left.n9 drain_left.t6 30.0005
R343 drain_left.n9 drain_left.t10 30.0005
R344 drain_left.n8 drain_left.t12 30.0005
R345 drain_left.n8 drain_left.t3 30.0005
R346 drain_left drain_left.n7 23.5165
R347 drain_left drain_left.n16 6.21356
R348 drain_left.n12 drain_left.n10 0.560845
R349 drain_left.n14 drain_left.n12 0.560845
R350 drain_left.n16 drain_left.n14 0.560845
R351 drain_left.n7 drain_left.n6 0.505499
R352 drain_left.n7 drain_left.n2 0.505499
C0 plus minus 3.78614f
C1 drain_left source 6.27021f
C2 plus source 1.15913f
C3 minus source 1.14526f
C4 drain_left drain_right 1.13612f
C5 drain_right plus 0.373605f
C6 drain_right minus 0.87893f
C7 drain_right source 6.2707f
C8 drain_left plus 1.08952f
C9 drain_left minus 0.178941f
C10 drain_right a_n2146_n1088# 4.06904f
C11 drain_left a_n2146_n1088# 4.3547f
C12 source a_n2146_n1088# 2.771954f
C13 minus a_n2146_n1088# 7.034099f
C14 plus a_n2146_n1088# 7.830209f
C15 drain_left.t16 a_n2146_n1088# 0.028926f
C16 drain_left.t9 a_n2146_n1088# 0.028926f
C17 drain_left.n0 a_n2146_n1088# 0.094472f
C18 drain_left.t1 a_n2146_n1088# 0.028926f
C19 drain_left.t19 a_n2146_n1088# 0.028926f
C20 drain_left.n1 a_n2146_n1088# 0.093853f
C21 drain_left.n2 a_n2146_n1088# 0.518291f
C22 drain_left.t18 a_n2146_n1088# 0.028926f
C23 drain_left.t14 a_n2146_n1088# 0.028926f
C24 drain_left.n3 a_n2146_n1088# 0.093853f
C25 drain_left.t17 a_n2146_n1088# 0.028926f
C26 drain_left.t15 a_n2146_n1088# 0.028926f
C27 drain_left.n4 a_n2146_n1088# 0.094472f
C28 drain_left.t11 a_n2146_n1088# 0.028926f
C29 drain_left.t2 a_n2146_n1088# 0.028926f
C30 drain_left.n5 a_n2146_n1088# 0.093853f
C31 drain_left.n6 a_n2146_n1088# 0.518291f
C32 drain_left.n7 a_n2146_n1088# 0.93692f
C33 drain_left.t12 a_n2146_n1088# 0.028926f
C34 drain_left.t3 a_n2146_n1088# 0.028926f
C35 drain_left.n8 a_n2146_n1088# 0.094472f
C36 drain_left.t6 a_n2146_n1088# 0.028926f
C37 drain_left.t10 a_n2146_n1088# 0.028926f
C38 drain_left.n9 a_n2146_n1088# 0.093853f
C39 drain_left.n10 a_n2146_n1088# 0.52149f
C40 drain_left.t0 a_n2146_n1088# 0.028926f
C41 drain_left.t4 a_n2146_n1088# 0.028926f
C42 drain_left.n11 a_n2146_n1088# 0.093853f
C43 drain_left.n12 a_n2146_n1088# 0.256189f
C44 drain_left.t7 a_n2146_n1088# 0.028926f
C45 drain_left.t13 a_n2146_n1088# 0.028926f
C46 drain_left.n13 a_n2146_n1088# 0.093853f
C47 drain_left.n14 a_n2146_n1088# 0.256189f
C48 drain_left.t5 a_n2146_n1088# 0.028926f
C49 drain_left.t8 a_n2146_n1088# 0.028926f
C50 drain_left.n15 a_n2146_n1088# 0.093853f
C51 drain_left.n16 a_n2146_n1088# 0.457944f
C52 plus.n0 a_n2146_n1088# 0.033997f
C53 plus.t14 a_n2146_n1088# 0.01572f
C54 plus.t6 a_n2146_n1088# 0.01572f
C55 plus.n1 a_n2146_n1088# 0.011802f
C56 plus.n2 a_n2146_n1088# 0.033997f
C57 plus.t15 a_n2146_n1088# 0.01572f
C58 plus.t19 a_n2146_n1088# 0.01572f
C59 plus.t9 a_n2146_n1088# 0.01572f
C60 plus.n3 a_n2146_n1088# 0.021437f
C61 plus.n4 a_n2146_n1088# 0.033997f
C62 plus.t13 a_n2146_n1088# 0.01572f
C63 plus.t16 a_n2146_n1088# 0.01572f
C64 plus.n5 a_n2146_n1088# 0.021437f
C65 plus.t7 a_n2146_n1088# 0.01903f
C66 plus.n6 a_n2146_n1088# 0.034174f
C67 plus.n7 a_n2146_n1088# 0.078422f
C68 plus.n8 a_n2146_n1088# 0.014422f
C69 plus.n9 a_n2146_n1088# 0.021437f
C70 plus.n10 a_n2146_n1088# 0.013898f
C71 plus.n11 a_n2146_n1088# 0.011802f
C72 plus.n12 a_n2146_n1088# 0.033997f
C73 plus.n13 a_n2146_n1088# 0.033997f
C74 plus.n14 a_n2146_n1088# 0.014422f
C75 plus.n15 a_n2146_n1088# 0.021437f
C76 plus.n16 a_n2146_n1088# 0.014422f
C77 plus.n17 a_n2146_n1088# 0.021437f
C78 plus.t12 a_n2146_n1088# 0.01572f
C79 plus.n18 a_n2146_n1088# 0.021437f
C80 plus.n19 a_n2146_n1088# 0.014422f
C81 plus.n20 a_n2146_n1088# 0.033997f
C82 plus.n21 a_n2146_n1088# 0.033997f
C83 plus.n22 a_n2146_n1088# 0.033997f
C84 plus.n23 a_n2146_n1088# 0.013898f
C85 plus.n24 a_n2146_n1088# 0.021437f
C86 plus.n25 a_n2146_n1088# 0.014422f
C87 plus.n26 a_n2146_n1088# 0.021437f
C88 plus.t11 a_n2146_n1088# 0.01903f
C89 plus.n27 a_n2146_n1088# 0.034122f
C90 plus.n28 a_n2146_n1088# 0.238227f
C91 plus.n29 a_n2146_n1088# 0.033997f
C92 plus.t3 a_n2146_n1088# 0.01903f
C93 plus.t10 a_n2146_n1088# 0.01572f
C94 plus.t18 a_n2146_n1088# 0.01572f
C95 plus.n30 a_n2146_n1088# 0.011802f
C96 plus.n31 a_n2146_n1088# 0.033997f
C97 plus.t0 a_n2146_n1088# 0.01572f
C98 plus.n32 a_n2146_n1088# 0.021437f
C99 plus.t1 a_n2146_n1088# 0.01572f
C100 plus.t5 a_n2146_n1088# 0.01572f
C101 plus.t8 a_n2146_n1088# 0.01572f
C102 plus.n33 a_n2146_n1088# 0.021437f
C103 plus.n34 a_n2146_n1088# 0.033997f
C104 plus.t17 a_n2146_n1088# 0.01572f
C105 plus.t2 a_n2146_n1088# 0.01572f
C106 plus.n35 a_n2146_n1088# 0.021437f
C107 plus.t4 a_n2146_n1088# 0.01903f
C108 plus.n36 a_n2146_n1088# 0.034174f
C109 plus.n37 a_n2146_n1088# 0.078422f
C110 plus.n38 a_n2146_n1088# 0.014422f
C111 plus.n39 a_n2146_n1088# 0.021437f
C112 plus.n40 a_n2146_n1088# 0.013898f
C113 plus.n41 a_n2146_n1088# 0.011802f
C114 plus.n42 a_n2146_n1088# 0.033997f
C115 plus.n43 a_n2146_n1088# 0.033997f
C116 plus.n44 a_n2146_n1088# 0.014422f
C117 plus.n45 a_n2146_n1088# 0.021437f
C118 plus.n46 a_n2146_n1088# 0.014422f
C119 plus.n47 a_n2146_n1088# 0.021437f
C120 plus.n48 a_n2146_n1088# 0.014422f
C121 plus.n49 a_n2146_n1088# 0.033997f
C122 plus.n50 a_n2146_n1088# 0.033997f
C123 plus.n51 a_n2146_n1088# 0.033997f
C124 plus.n52 a_n2146_n1088# 0.013898f
C125 plus.n53 a_n2146_n1088# 0.021437f
C126 plus.n54 a_n2146_n1088# 0.014422f
C127 plus.n55 a_n2146_n1088# 0.021437f
C128 plus.n56 a_n2146_n1088# 0.034122f
C129 plus.n57 a_n2146_n1088# 0.807685f
C130 drain_right.t7 a_n2146_n1088# 0.029367f
C131 drain_right.t16 a_n2146_n1088# 0.029367f
C132 drain_right.n0 a_n2146_n1088# 0.095911f
C133 drain_right.t18 a_n2146_n1088# 0.029367f
C134 drain_right.t19 a_n2146_n1088# 0.029367f
C135 drain_right.n1 a_n2146_n1088# 0.095282f
C136 drain_right.n2 a_n2146_n1088# 0.526184f
C137 drain_right.t10 a_n2146_n1088# 0.029367f
C138 drain_right.t14 a_n2146_n1088# 0.029367f
C139 drain_right.n3 a_n2146_n1088# 0.095282f
C140 drain_right.t0 a_n2146_n1088# 0.029367f
C141 drain_right.t3 a_n2146_n1088# 0.029367f
C142 drain_right.n4 a_n2146_n1088# 0.095911f
C143 drain_right.t15 a_n2146_n1088# 0.029367f
C144 drain_right.t17 a_n2146_n1088# 0.029367f
C145 drain_right.n5 a_n2146_n1088# 0.095282f
C146 drain_right.n6 a_n2146_n1088# 0.526184f
C147 drain_right.n7 a_n2146_n1088# 0.903883f
C148 drain_right.t13 a_n2146_n1088# 0.029367f
C149 drain_right.t12 a_n2146_n1088# 0.029367f
C150 drain_right.n8 a_n2146_n1088# 0.095911f
C151 drain_right.t9 a_n2146_n1088# 0.029367f
C152 drain_right.t6 a_n2146_n1088# 0.029367f
C153 drain_right.n9 a_n2146_n1088# 0.095282f
C154 drain_right.n10 a_n2146_n1088# 0.529432f
C155 drain_right.t2 a_n2146_n1088# 0.029367f
C156 drain_right.t11 a_n2146_n1088# 0.029367f
C157 drain_right.n11 a_n2146_n1088# 0.095282f
C158 drain_right.n12 a_n2146_n1088# 0.260091f
C159 drain_right.t4 a_n2146_n1088# 0.029367f
C160 drain_right.t5 a_n2146_n1088# 0.029367f
C161 drain_right.n13 a_n2146_n1088# 0.095282f
C162 drain_right.n14 a_n2146_n1088# 0.260091f
C163 drain_right.t1 a_n2146_n1088# 0.029367f
C164 drain_right.t8 a_n2146_n1088# 0.029367f
C165 drain_right.n15 a_n2146_n1088# 0.095282f
C166 drain_right.n16 a_n2146_n1088# 0.464918f
C167 source.t8 a_n2146_n1088# 0.143844f
C168 source.n0 a_n2146_n1088# 0.549644f
C169 source.t31 a_n2146_n1088# 0.034314f
C170 source.t33 a_n2146_n1088# 0.034314f
C171 source.n1 a_n2146_n1088# 0.096783f
C172 source.n2 a_n2146_n1088# 0.279508f
C173 source.t6 a_n2146_n1088# 0.034314f
C174 source.t37 a_n2146_n1088# 0.034314f
C175 source.n3 a_n2146_n1088# 0.096783f
C176 source.n4 a_n2146_n1088# 0.279508f
C177 source.t30 a_n2146_n1088# 0.034314f
C178 source.t34 a_n2146_n1088# 0.034314f
C179 source.n5 a_n2146_n1088# 0.096783f
C180 source.n6 a_n2146_n1088# 0.279508f
C181 source.t7 a_n2146_n1088# 0.034314f
C182 source.t35 a_n2146_n1088# 0.034314f
C183 source.n7 a_n2146_n1088# 0.096783f
C184 source.n8 a_n2146_n1088# 0.279508f
C185 source.t39 a_n2146_n1088# 0.143844f
C186 source.n9 a_n2146_n1088# 0.285854f
C187 source.t26 a_n2146_n1088# 0.143844f
C188 source.n10 a_n2146_n1088# 0.285854f
C189 source.t12 a_n2146_n1088# 0.034314f
C190 source.t23 a_n2146_n1088# 0.034314f
C191 source.n11 a_n2146_n1088# 0.096783f
C192 source.n12 a_n2146_n1088# 0.279508f
C193 source.t27 a_n2146_n1088# 0.034314f
C194 source.t15 a_n2146_n1088# 0.034314f
C195 source.n13 a_n2146_n1088# 0.096783f
C196 source.n14 a_n2146_n1088# 0.279508f
C197 source.t11 a_n2146_n1088# 0.034314f
C198 source.t25 a_n2146_n1088# 0.034314f
C199 source.n15 a_n2146_n1088# 0.096783f
C200 source.n16 a_n2146_n1088# 0.279508f
C201 source.t10 a_n2146_n1088# 0.034314f
C202 source.t14 a_n2146_n1088# 0.034314f
C203 source.n17 a_n2146_n1088# 0.096783f
C204 source.n18 a_n2146_n1088# 0.279508f
C205 source.t24 a_n2146_n1088# 0.143844f
C206 source.n19 a_n2146_n1088# 0.779623f
C207 source.t2 a_n2146_n1088# 0.143844f
C208 source.n20 a_n2146_n1088# 0.779623f
C209 source.t9 a_n2146_n1088# 0.034314f
C210 source.t38 a_n2146_n1088# 0.034314f
C211 source.n21 a_n2146_n1088# 0.096783f
C212 source.n22 a_n2146_n1088# 0.279508f
C213 source.t4 a_n2146_n1088# 0.034314f
C214 source.t3 a_n2146_n1088# 0.034314f
C215 source.n23 a_n2146_n1088# 0.096783f
C216 source.n24 a_n2146_n1088# 0.279508f
C217 source.t0 a_n2146_n1088# 0.034314f
C218 source.t36 a_n2146_n1088# 0.034314f
C219 source.n25 a_n2146_n1088# 0.096783f
C220 source.n26 a_n2146_n1088# 0.279508f
C221 source.t32 a_n2146_n1088# 0.034314f
C222 source.t5 a_n2146_n1088# 0.034314f
C223 source.n27 a_n2146_n1088# 0.096783f
C224 source.n28 a_n2146_n1088# 0.279508f
C225 source.t1 a_n2146_n1088# 0.143844f
C226 source.n29 a_n2146_n1088# 0.285854f
C227 source.t16 a_n2146_n1088# 0.143844f
C228 source.n30 a_n2146_n1088# 0.285854f
C229 source.t21 a_n2146_n1088# 0.034314f
C230 source.t28 a_n2146_n1088# 0.034314f
C231 source.n31 a_n2146_n1088# 0.096783f
C232 source.n32 a_n2146_n1088# 0.279508f
C233 source.t20 a_n2146_n1088# 0.034314f
C234 source.t18 a_n2146_n1088# 0.034314f
C235 source.n33 a_n2146_n1088# 0.096783f
C236 source.n34 a_n2146_n1088# 0.279508f
C237 source.t13 a_n2146_n1088# 0.034314f
C238 source.t22 a_n2146_n1088# 0.034314f
C239 source.n35 a_n2146_n1088# 0.096783f
C240 source.n36 a_n2146_n1088# 0.279508f
C241 source.t19 a_n2146_n1088# 0.034314f
C242 source.t29 a_n2146_n1088# 0.034314f
C243 source.n37 a_n2146_n1088# 0.096783f
C244 source.n38 a_n2146_n1088# 0.279508f
C245 source.t17 a_n2146_n1088# 0.143844f
C246 source.n39 a_n2146_n1088# 0.448907f
C247 source.n40 a_n2146_n1088# 0.58108f
C248 minus.n0 a_n2146_n1088# 0.033393f
C249 minus.t18 a_n2146_n1088# 0.018692f
C250 minus.t11 a_n2146_n1088# 0.015441f
C251 minus.t15 a_n2146_n1088# 0.015441f
C252 minus.n1 a_n2146_n1088# 0.011592f
C253 minus.n2 a_n2146_n1088# 0.033393f
C254 minus.t14 a_n2146_n1088# 0.015441f
C255 minus.n3 a_n2146_n1088# 0.021056f
C256 minus.t17 a_n2146_n1088# 0.015441f
C257 minus.t8 a_n2146_n1088# 0.015441f
C258 minus.t10 a_n2146_n1088# 0.015441f
C259 minus.n4 a_n2146_n1088# 0.021056f
C260 minus.n5 a_n2146_n1088# 0.033393f
C261 minus.t13 a_n2146_n1088# 0.015441f
C262 minus.t6 a_n2146_n1088# 0.015441f
C263 minus.n6 a_n2146_n1088# 0.021056f
C264 minus.t7 a_n2146_n1088# 0.018692f
C265 minus.n7 a_n2146_n1088# 0.033567f
C266 minus.n8 a_n2146_n1088# 0.077029f
C267 minus.n9 a_n2146_n1088# 0.014166f
C268 minus.n10 a_n2146_n1088# 0.021056f
C269 minus.n11 a_n2146_n1088# 0.013651f
C270 minus.n12 a_n2146_n1088# 0.011592f
C271 minus.n13 a_n2146_n1088# 0.033393f
C272 minus.n14 a_n2146_n1088# 0.033393f
C273 minus.n15 a_n2146_n1088# 0.014166f
C274 minus.n16 a_n2146_n1088# 0.021056f
C275 minus.n17 a_n2146_n1088# 0.014166f
C276 minus.n18 a_n2146_n1088# 0.021056f
C277 minus.n19 a_n2146_n1088# 0.014166f
C278 minus.n20 a_n2146_n1088# 0.033393f
C279 minus.n21 a_n2146_n1088# 0.033393f
C280 minus.n22 a_n2146_n1088# 0.033393f
C281 minus.n23 a_n2146_n1088# 0.013651f
C282 minus.n24 a_n2146_n1088# 0.021056f
C283 minus.n25 a_n2146_n1088# 0.014166f
C284 minus.n26 a_n2146_n1088# 0.021056f
C285 minus.n27 a_n2146_n1088# 0.033515f
C286 minus.n28 a_n2146_n1088# 0.820289f
C287 minus.n29 a_n2146_n1088# 0.033393f
C288 minus.t19 a_n2146_n1088# 0.015441f
C289 minus.t2 a_n2146_n1088# 0.015441f
C290 minus.n30 a_n2146_n1088# 0.011592f
C291 minus.n31 a_n2146_n1088# 0.033393f
C292 minus.t5 a_n2146_n1088# 0.015441f
C293 minus.t9 a_n2146_n1088# 0.015441f
C294 minus.t0 a_n2146_n1088# 0.015441f
C295 minus.n32 a_n2146_n1088# 0.021056f
C296 minus.n33 a_n2146_n1088# 0.033393f
C297 minus.t1 a_n2146_n1088# 0.015441f
C298 minus.t3 a_n2146_n1088# 0.015441f
C299 minus.n34 a_n2146_n1088# 0.021056f
C300 minus.t12 a_n2146_n1088# 0.018692f
C301 minus.n35 a_n2146_n1088# 0.033567f
C302 minus.n36 a_n2146_n1088# 0.077029f
C303 minus.n37 a_n2146_n1088# 0.014166f
C304 minus.n38 a_n2146_n1088# 0.021056f
C305 minus.n39 a_n2146_n1088# 0.013651f
C306 minus.n40 a_n2146_n1088# 0.011592f
C307 minus.n41 a_n2146_n1088# 0.033393f
C308 minus.n42 a_n2146_n1088# 0.033393f
C309 minus.n43 a_n2146_n1088# 0.014166f
C310 minus.n44 a_n2146_n1088# 0.021056f
C311 minus.n45 a_n2146_n1088# 0.014166f
C312 minus.n46 a_n2146_n1088# 0.021056f
C313 minus.t4 a_n2146_n1088# 0.015441f
C314 minus.n47 a_n2146_n1088# 0.021056f
C315 minus.n48 a_n2146_n1088# 0.014166f
C316 minus.n49 a_n2146_n1088# 0.033393f
C317 minus.n50 a_n2146_n1088# 0.033393f
C318 minus.n51 a_n2146_n1088# 0.033393f
C319 minus.n52 a_n2146_n1088# 0.013651f
C320 minus.n53 a_n2146_n1088# 0.021056f
C321 minus.n54 a_n2146_n1088# 0.014166f
C322 minus.n55 a_n2146_n1088# 0.021056f
C323 minus.t16 a_n2146_n1088# 0.018692f
C324 minus.n56 a_n2146_n1088# 0.033515f
C325 minus.n57 a_n2146_n1088# 0.223108f
C326 minus.n58 a_n2146_n1088# 1.01081f
.ends

