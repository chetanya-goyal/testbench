* NGSPICE file created from diffpair675.ext - technology: sky130A

.subckt diffpair675 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t1 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X1 drain_right.t0 minus.t1 source.t22 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X2 source.t21 minus.t2 drain_right.t5 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X3 source.t20 minus.t3 drain_right.t4 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X4 a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X5 source.t9 plus.t0 drain_left.t11 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X6 drain_left.t10 plus.t1 source.t0 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X7 a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X8 a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X9 a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X10 source.t8 plus.t2 drain_left.t9 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X11 drain_left.t8 plus.t3 source.t11 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X12 source.t19 minus.t4 drain_right.t7 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X13 source.t18 minus.t5 drain_right.t6 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X14 source.t1 plus.t4 drain_left.t7 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X15 drain_right.t3 minus.t6 source.t17 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X16 drain_left.t6 plus.t5 source.t2 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X17 source.t3 plus.t6 drain_left.t5 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X18 source.t7 plus.t7 drain_left.t4 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X19 source.t10 plus.t8 drain_left.t3 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X20 drain_right.t2 minus.t7 source.t16 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X21 drain_right.t9 minus.t8 source.t15 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X22 drain_right.t8 minus.t9 source.t14 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X23 source.t13 minus.t10 drain_right.t11 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X24 drain_right.t10 minus.t11 source.t12 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X25 drain_left.t2 plus.t9 source.t4 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X26 drain_left.t1 plus.t10 source.t6 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X27 drain_left.t0 plus.t11 source.t5 a_n1598_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
R0 minus.n13 minus.t0 2160.24
R1 minus.n2 minus.t6 2160.24
R2 minus.n28 minus.t11 2160.24
R3 minus.n17 minus.t3 2160.24
R4 minus.n12 minus.t9 2112.77
R5 minus.n10 minus.t5 2112.77
R6 minus.n3 minus.t1 2112.77
R7 minus.n4 minus.t10 2112.77
R8 minus.n27 minus.t4 2112.77
R9 minus.n25 minus.t7 2112.77
R10 minus.n19 minus.t2 2112.77
R11 minus.n18 minus.t8 2112.77
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n30 minus.n14 45.0346
R31 minus.n13 minus.n12 44.549
R32 minus.n4 minus.n2 44.549
R33 minus.n18 minus.n17 44.549
R34 minus.n28 minus.n27 44.549
R35 minus.n12 minus.n11 28.4823
R36 minus.n5 minus.n4 28.4823
R37 minus.n20 minus.n18 28.4823
R38 minus.n27 minus.n26 28.4823
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 59.2584
R54 drain_right.n3 drain_right.n2 59.2032
R55 drain_right.n3 drain_right.n0 59.2032
R56 drain_right.n3 drain_right.n1 58.7154
R57 drain_right.n6 drain_right.n5 58.7154
R58 drain_right.n8 drain_right.n7 58.7154
R59 drain_right drain_right.n3 39.3778
R60 drain_right drain_right.n8 6.19632
R61 drain_right.n1 drain_right.t5 0.7925
R62 drain_right.n1 drain_right.t2 0.7925
R63 drain_right.n2 drain_right.t7 0.7925
R64 drain_right.n2 drain_right.t10 0.7925
R65 drain_right.n0 drain_right.t4 0.7925
R66 drain_right.n0 drain_right.t9 0.7925
R67 drain_right.n4 drain_right.t11 0.7925
R68 drain_right.n4 drain_right.t3 0.7925
R69 drain_right.n5 drain_right.t6 0.7925
R70 drain_right.n5 drain_right.t0 0.7925
R71 drain_right.n7 drain_right.t1 0.7925
R72 drain_right.n7 drain_right.t8 0.7925
R73 drain_right.n8 drain_right.n6 0.543603
R74 source.n1130 source.n996 289.615
R75 source.n986 source.n852 289.615
R76 source.n846 source.n712 289.615
R77 source.n702 source.n568 289.615
R78 source.n134 source.n0 289.615
R79 source.n278 source.n144 289.615
R80 source.n418 source.n284 289.615
R81 source.n562 source.n428 289.615
R82 source.n1040 source.n1039 185
R83 source.n1045 source.n1044 185
R84 source.n1047 source.n1046 185
R85 source.n1036 source.n1035 185
R86 source.n1053 source.n1052 185
R87 source.n1055 source.n1054 185
R88 source.n1032 source.n1031 185
R89 source.n1062 source.n1061 185
R90 source.n1063 source.n1030 185
R91 source.n1065 source.n1064 185
R92 source.n1028 source.n1027 185
R93 source.n1071 source.n1070 185
R94 source.n1073 source.n1072 185
R95 source.n1024 source.n1023 185
R96 source.n1079 source.n1078 185
R97 source.n1081 source.n1080 185
R98 source.n1020 source.n1019 185
R99 source.n1087 source.n1086 185
R100 source.n1089 source.n1088 185
R101 source.n1016 source.n1015 185
R102 source.n1095 source.n1094 185
R103 source.n1097 source.n1096 185
R104 source.n1012 source.n1011 185
R105 source.n1103 source.n1102 185
R106 source.n1106 source.n1105 185
R107 source.n1104 source.n1008 185
R108 source.n1111 source.n1007 185
R109 source.n1113 source.n1112 185
R110 source.n1115 source.n1114 185
R111 source.n1004 source.n1003 185
R112 source.n1121 source.n1120 185
R113 source.n1123 source.n1122 185
R114 source.n1000 source.n999 185
R115 source.n1129 source.n1128 185
R116 source.n1131 source.n1130 185
R117 source.n896 source.n895 185
R118 source.n901 source.n900 185
R119 source.n903 source.n902 185
R120 source.n892 source.n891 185
R121 source.n909 source.n908 185
R122 source.n911 source.n910 185
R123 source.n888 source.n887 185
R124 source.n918 source.n917 185
R125 source.n919 source.n886 185
R126 source.n921 source.n920 185
R127 source.n884 source.n883 185
R128 source.n927 source.n926 185
R129 source.n929 source.n928 185
R130 source.n880 source.n879 185
R131 source.n935 source.n934 185
R132 source.n937 source.n936 185
R133 source.n876 source.n875 185
R134 source.n943 source.n942 185
R135 source.n945 source.n944 185
R136 source.n872 source.n871 185
R137 source.n951 source.n950 185
R138 source.n953 source.n952 185
R139 source.n868 source.n867 185
R140 source.n959 source.n958 185
R141 source.n962 source.n961 185
R142 source.n960 source.n864 185
R143 source.n967 source.n863 185
R144 source.n969 source.n968 185
R145 source.n971 source.n970 185
R146 source.n860 source.n859 185
R147 source.n977 source.n976 185
R148 source.n979 source.n978 185
R149 source.n856 source.n855 185
R150 source.n985 source.n984 185
R151 source.n987 source.n986 185
R152 source.n756 source.n755 185
R153 source.n761 source.n760 185
R154 source.n763 source.n762 185
R155 source.n752 source.n751 185
R156 source.n769 source.n768 185
R157 source.n771 source.n770 185
R158 source.n748 source.n747 185
R159 source.n778 source.n777 185
R160 source.n779 source.n746 185
R161 source.n781 source.n780 185
R162 source.n744 source.n743 185
R163 source.n787 source.n786 185
R164 source.n789 source.n788 185
R165 source.n740 source.n739 185
R166 source.n795 source.n794 185
R167 source.n797 source.n796 185
R168 source.n736 source.n735 185
R169 source.n803 source.n802 185
R170 source.n805 source.n804 185
R171 source.n732 source.n731 185
R172 source.n811 source.n810 185
R173 source.n813 source.n812 185
R174 source.n728 source.n727 185
R175 source.n819 source.n818 185
R176 source.n822 source.n821 185
R177 source.n820 source.n724 185
R178 source.n827 source.n723 185
R179 source.n829 source.n828 185
R180 source.n831 source.n830 185
R181 source.n720 source.n719 185
R182 source.n837 source.n836 185
R183 source.n839 source.n838 185
R184 source.n716 source.n715 185
R185 source.n845 source.n844 185
R186 source.n847 source.n846 185
R187 source.n612 source.n611 185
R188 source.n617 source.n616 185
R189 source.n619 source.n618 185
R190 source.n608 source.n607 185
R191 source.n625 source.n624 185
R192 source.n627 source.n626 185
R193 source.n604 source.n603 185
R194 source.n634 source.n633 185
R195 source.n635 source.n602 185
R196 source.n637 source.n636 185
R197 source.n600 source.n599 185
R198 source.n643 source.n642 185
R199 source.n645 source.n644 185
R200 source.n596 source.n595 185
R201 source.n651 source.n650 185
R202 source.n653 source.n652 185
R203 source.n592 source.n591 185
R204 source.n659 source.n658 185
R205 source.n661 source.n660 185
R206 source.n588 source.n587 185
R207 source.n667 source.n666 185
R208 source.n669 source.n668 185
R209 source.n584 source.n583 185
R210 source.n675 source.n674 185
R211 source.n678 source.n677 185
R212 source.n676 source.n580 185
R213 source.n683 source.n579 185
R214 source.n685 source.n684 185
R215 source.n687 source.n686 185
R216 source.n576 source.n575 185
R217 source.n693 source.n692 185
R218 source.n695 source.n694 185
R219 source.n572 source.n571 185
R220 source.n701 source.n700 185
R221 source.n703 source.n702 185
R222 source.n135 source.n134 185
R223 source.n133 source.n132 185
R224 source.n4 source.n3 185
R225 source.n127 source.n126 185
R226 source.n125 source.n124 185
R227 source.n8 source.n7 185
R228 source.n119 source.n118 185
R229 source.n117 source.n116 185
R230 source.n115 source.n11 185
R231 source.n15 source.n12 185
R232 source.n110 source.n109 185
R233 source.n108 source.n107 185
R234 source.n17 source.n16 185
R235 source.n102 source.n101 185
R236 source.n100 source.n99 185
R237 source.n21 source.n20 185
R238 source.n94 source.n93 185
R239 source.n92 source.n91 185
R240 source.n25 source.n24 185
R241 source.n86 source.n85 185
R242 source.n84 source.n83 185
R243 source.n29 source.n28 185
R244 source.n78 source.n77 185
R245 source.n76 source.n75 185
R246 source.n33 source.n32 185
R247 source.n70 source.n69 185
R248 source.n68 source.n35 185
R249 source.n67 source.n66 185
R250 source.n38 source.n36 185
R251 source.n61 source.n60 185
R252 source.n59 source.n58 185
R253 source.n42 source.n41 185
R254 source.n53 source.n52 185
R255 source.n51 source.n50 185
R256 source.n46 source.n45 185
R257 source.n279 source.n278 185
R258 source.n277 source.n276 185
R259 source.n148 source.n147 185
R260 source.n271 source.n270 185
R261 source.n269 source.n268 185
R262 source.n152 source.n151 185
R263 source.n263 source.n262 185
R264 source.n261 source.n260 185
R265 source.n259 source.n155 185
R266 source.n159 source.n156 185
R267 source.n254 source.n253 185
R268 source.n252 source.n251 185
R269 source.n161 source.n160 185
R270 source.n246 source.n245 185
R271 source.n244 source.n243 185
R272 source.n165 source.n164 185
R273 source.n238 source.n237 185
R274 source.n236 source.n235 185
R275 source.n169 source.n168 185
R276 source.n230 source.n229 185
R277 source.n228 source.n227 185
R278 source.n173 source.n172 185
R279 source.n222 source.n221 185
R280 source.n220 source.n219 185
R281 source.n177 source.n176 185
R282 source.n214 source.n213 185
R283 source.n212 source.n179 185
R284 source.n211 source.n210 185
R285 source.n182 source.n180 185
R286 source.n205 source.n204 185
R287 source.n203 source.n202 185
R288 source.n186 source.n185 185
R289 source.n197 source.n196 185
R290 source.n195 source.n194 185
R291 source.n190 source.n189 185
R292 source.n419 source.n418 185
R293 source.n417 source.n416 185
R294 source.n288 source.n287 185
R295 source.n411 source.n410 185
R296 source.n409 source.n408 185
R297 source.n292 source.n291 185
R298 source.n403 source.n402 185
R299 source.n401 source.n400 185
R300 source.n399 source.n295 185
R301 source.n299 source.n296 185
R302 source.n394 source.n393 185
R303 source.n392 source.n391 185
R304 source.n301 source.n300 185
R305 source.n386 source.n385 185
R306 source.n384 source.n383 185
R307 source.n305 source.n304 185
R308 source.n378 source.n377 185
R309 source.n376 source.n375 185
R310 source.n309 source.n308 185
R311 source.n370 source.n369 185
R312 source.n368 source.n367 185
R313 source.n313 source.n312 185
R314 source.n362 source.n361 185
R315 source.n360 source.n359 185
R316 source.n317 source.n316 185
R317 source.n354 source.n353 185
R318 source.n352 source.n319 185
R319 source.n351 source.n350 185
R320 source.n322 source.n320 185
R321 source.n345 source.n344 185
R322 source.n343 source.n342 185
R323 source.n326 source.n325 185
R324 source.n337 source.n336 185
R325 source.n335 source.n334 185
R326 source.n330 source.n329 185
R327 source.n563 source.n562 185
R328 source.n561 source.n560 185
R329 source.n432 source.n431 185
R330 source.n555 source.n554 185
R331 source.n553 source.n552 185
R332 source.n436 source.n435 185
R333 source.n547 source.n546 185
R334 source.n545 source.n544 185
R335 source.n543 source.n439 185
R336 source.n443 source.n440 185
R337 source.n538 source.n537 185
R338 source.n536 source.n535 185
R339 source.n445 source.n444 185
R340 source.n530 source.n529 185
R341 source.n528 source.n527 185
R342 source.n449 source.n448 185
R343 source.n522 source.n521 185
R344 source.n520 source.n519 185
R345 source.n453 source.n452 185
R346 source.n514 source.n513 185
R347 source.n512 source.n511 185
R348 source.n457 source.n456 185
R349 source.n506 source.n505 185
R350 source.n504 source.n503 185
R351 source.n461 source.n460 185
R352 source.n498 source.n497 185
R353 source.n496 source.n463 185
R354 source.n495 source.n494 185
R355 source.n466 source.n464 185
R356 source.n489 source.n488 185
R357 source.n487 source.n486 185
R358 source.n470 source.n469 185
R359 source.n481 source.n480 185
R360 source.n479 source.n478 185
R361 source.n474 source.n473 185
R362 source.n1041 source.t12 149.524
R363 source.n897 source.t20 149.524
R364 source.n757 source.t6 149.524
R365 source.n613 source.t10 149.524
R366 source.n47 source.t2 149.524
R367 source.n191 source.t9 149.524
R368 source.n331 source.t17 149.524
R369 source.n475 source.t23 149.524
R370 source.n1045 source.n1039 104.615
R371 source.n1046 source.n1045 104.615
R372 source.n1046 source.n1035 104.615
R373 source.n1053 source.n1035 104.615
R374 source.n1054 source.n1053 104.615
R375 source.n1054 source.n1031 104.615
R376 source.n1062 source.n1031 104.615
R377 source.n1063 source.n1062 104.615
R378 source.n1064 source.n1063 104.615
R379 source.n1064 source.n1027 104.615
R380 source.n1071 source.n1027 104.615
R381 source.n1072 source.n1071 104.615
R382 source.n1072 source.n1023 104.615
R383 source.n1079 source.n1023 104.615
R384 source.n1080 source.n1079 104.615
R385 source.n1080 source.n1019 104.615
R386 source.n1087 source.n1019 104.615
R387 source.n1088 source.n1087 104.615
R388 source.n1088 source.n1015 104.615
R389 source.n1095 source.n1015 104.615
R390 source.n1096 source.n1095 104.615
R391 source.n1096 source.n1011 104.615
R392 source.n1103 source.n1011 104.615
R393 source.n1105 source.n1103 104.615
R394 source.n1105 source.n1104 104.615
R395 source.n1104 source.n1007 104.615
R396 source.n1113 source.n1007 104.615
R397 source.n1114 source.n1113 104.615
R398 source.n1114 source.n1003 104.615
R399 source.n1121 source.n1003 104.615
R400 source.n1122 source.n1121 104.615
R401 source.n1122 source.n999 104.615
R402 source.n1129 source.n999 104.615
R403 source.n1130 source.n1129 104.615
R404 source.n901 source.n895 104.615
R405 source.n902 source.n901 104.615
R406 source.n902 source.n891 104.615
R407 source.n909 source.n891 104.615
R408 source.n910 source.n909 104.615
R409 source.n910 source.n887 104.615
R410 source.n918 source.n887 104.615
R411 source.n919 source.n918 104.615
R412 source.n920 source.n919 104.615
R413 source.n920 source.n883 104.615
R414 source.n927 source.n883 104.615
R415 source.n928 source.n927 104.615
R416 source.n928 source.n879 104.615
R417 source.n935 source.n879 104.615
R418 source.n936 source.n935 104.615
R419 source.n936 source.n875 104.615
R420 source.n943 source.n875 104.615
R421 source.n944 source.n943 104.615
R422 source.n944 source.n871 104.615
R423 source.n951 source.n871 104.615
R424 source.n952 source.n951 104.615
R425 source.n952 source.n867 104.615
R426 source.n959 source.n867 104.615
R427 source.n961 source.n959 104.615
R428 source.n961 source.n960 104.615
R429 source.n960 source.n863 104.615
R430 source.n969 source.n863 104.615
R431 source.n970 source.n969 104.615
R432 source.n970 source.n859 104.615
R433 source.n977 source.n859 104.615
R434 source.n978 source.n977 104.615
R435 source.n978 source.n855 104.615
R436 source.n985 source.n855 104.615
R437 source.n986 source.n985 104.615
R438 source.n761 source.n755 104.615
R439 source.n762 source.n761 104.615
R440 source.n762 source.n751 104.615
R441 source.n769 source.n751 104.615
R442 source.n770 source.n769 104.615
R443 source.n770 source.n747 104.615
R444 source.n778 source.n747 104.615
R445 source.n779 source.n778 104.615
R446 source.n780 source.n779 104.615
R447 source.n780 source.n743 104.615
R448 source.n787 source.n743 104.615
R449 source.n788 source.n787 104.615
R450 source.n788 source.n739 104.615
R451 source.n795 source.n739 104.615
R452 source.n796 source.n795 104.615
R453 source.n796 source.n735 104.615
R454 source.n803 source.n735 104.615
R455 source.n804 source.n803 104.615
R456 source.n804 source.n731 104.615
R457 source.n811 source.n731 104.615
R458 source.n812 source.n811 104.615
R459 source.n812 source.n727 104.615
R460 source.n819 source.n727 104.615
R461 source.n821 source.n819 104.615
R462 source.n821 source.n820 104.615
R463 source.n820 source.n723 104.615
R464 source.n829 source.n723 104.615
R465 source.n830 source.n829 104.615
R466 source.n830 source.n719 104.615
R467 source.n837 source.n719 104.615
R468 source.n838 source.n837 104.615
R469 source.n838 source.n715 104.615
R470 source.n845 source.n715 104.615
R471 source.n846 source.n845 104.615
R472 source.n617 source.n611 104.615
R473 source.n618 source.n617 104.615
R474 source.n618 source.n607 104.615
R475 source.n625 source.n607 104.615
R476 source.n626 source.n625 104.615
R477 source.n626 source.n603 104.615
R478 source.n634 source.n603 104.615
R479 source.n635 source.n634 104.615
R480 source.n636 source.n635 104.615
R481 source.n636 source.n599 104.615
R482 source.n643 source.n599 104.615
R483 source.n644 source.n643 104.615
R484 source.n644 source.n595 104.615
R485 source.n651 source.n595 104.615
R486 source.n652 source.n651 104.615
R487 source.n652 source.n591 104.615
R488 source.n659 source.n591 104.615
R489 source.n660 source.n659 104.615
R490 source.n660 source.n587 104.615
R491 source.n667 source.n587 104.615
R492 source.n668 source.n667 104.615
R493 source.n668 source.n583 104.615
R494 source.n675 source.n583 104.615
R495 source.n677 source.n675 104.615
R496 source.n677 source.n676 104.615
R497 source.n676 source.n579 104.615
R498 source.n685 source.n579 104.615
R499 source.n686 source.n685 104.615
R500 source.n686 source.n575 104.615
R501 source.n693 source.n575 104.615
R502 source.n694 source.n693 104.615
R503 source.n694 source.n571 104.615
R504 source.n701 source.n571 104.615
R505 source.n702 source.n701 104.615
R506 source.n134 source.n133 104.615
R507 source.n133 source.n3 104.615
R508 source.n126 source.n3 104.615
R509 source.n126 source.n125 104.615
R510 source.n125 source.n7 104.615
R511 source.n118 source.n7 104.615
R512 source.n118 source.n117 104.615
R513 source.n117 source.n11 104.615
R514 source.n15 source.n11 104.615
R515 source.n109 source.n15 104.615
R516 source.n109 source.n108 104.615
R517 source.n108 source.n16 104.615
R518 source.n101 source.n16 104.615
R519 source.n101 source.n100 104.615
R520 source.n100 source.n20 104.615
R521 source.n93 source.n20 104.615
R522 source.n93 source.n92 104.615
R523 source.n92 source.n24 104.615
R524 source.n85 source.n24 104.615
R525 source.n85 source.n84 104.615
R526 source.n84 source.n28 104.615
R527 source.n77 source.n28 104.615
R528 source.n77 source.n76 104.615
R529 source.n76 source.n32 104.615
R530 source.n69 source.n32 104.615
R531 source.n69 source.n68 104.615
R532 source.n68 source.n67 104.615
R533 source.n67 source.n36 104.615
R534 source.n60 source.n36 104.615
R535 source.n60 source.n59 104.615
R536 source.n59 source.n41 104.615
R537 source.n52 source.n41 104.615
R538 source.n52 source.n51 104.615
R539 source.n51 source.n45 104.615
R540 source.n278 source.n277 104.615
R541 source.n277 source.n147 104.615
R542 source.n270 source.n147 104.615
R543 source.n270 source.n269 104.615
R544 source.n269 source.n151 104.615
R545 source.n262 source.n151 104.615
R546 source.n262 source.n261 104.615
R547 source.n261 source.n155 104.615
R548 source.n159 source.n155 104.615
R549 source.n253 source.n159 104.615
R550 source.n253 source.n252 104.615
R551 source.n252 source.n160 104.615
R552 source.n245 source.n160 104.615
R553 source.n245 source.n244 104.615
R554 source.n244 source.n164 104.615
R555 source.n237 source.n164 104.615
R556 source.n237 source.n236 104.615
R557 source.n236 source.n168 104.615
R558 source.n229 source.n168 104.615
R559 source.n229 source.n228 104.615
R560 source.n228 source.n172 104.615
R561 source.n221 source.n172 104.615
R562 source.n221 source.n220 104.615
R563 source.n220 source.n176 104.615
R564 source.n213 source.n176 104.615
R565 source.n213 source.n212 104.615
R566 source.n212 source.n211 104.615
R567 source.n211 source.n180 104.615
R568 source.n204 source.n180 104.615
R569 source.n204 source.n203 104.615
R570 source.n203 source.n185 104.615
R571 source.n196 source.n185 104.615
R572 source.n196 source.n195 104.615
R573 source.n195 source.n189 104.615
R574 source.n418 source.n417 104.615
R575 source.n417 source.n287 104.615
R576 source.n410 source.n287 104.615
R577 source.n410 source.n409 104.615
R578 source.n409 source.n291 104.615
R579 source.n402 source.n291 104.615
R580 source.n402 source.n401 104.615
R581 source.n401 source.n295 104.615
R582 source.n299 source.n295 104.615
R583 source.n393 source.n299 104.615
R584 source.n393 source.n392 104.615
R585 source.n392 source.n300 104.615
R586 source.n385 source.n300 104.615
R587 source.n385 source.n384 104.615
R588 source.n384 source.n304 104.615
R589 source.n377 source.n304 104.615
R590 source.n377 source.n376 104.615
R591 source.n376 source.n308 104.615
R592 source.n369 source.n308 104.615
R593 source.n369 source.n368 104.615
R594 source.n368 source.n312 104.615
R595 source.n361 source.n312 104.615
R596 source.n361 source.n360 104.615
R597 source.n360 source.n316 104.615
R598 source.n353 source.n316 104.615
R599 source.n353 source.n352 104.615
R600 source.n352 source.n351 104.615
R601 source.n351 source.n320 104.615
R602 source.n344 source.n320 104.615
R603 source.n344 source.n343 104.615
R604 source.n343 source.n325 104.615
R605 source.n336 source.n325 104.615
R606 source.n336 source.n335 104.615
R607 source.n335 source.n329 104.615
R608 source.n562 source.n561 104.615
R609 source.n561 source.n431 104.615
R610 source.n554 source.n431 104.615
R611 source.n554 source.n553 104.615
R612 source.n553 source.n435 104.615
R613 source.n546 source.n435 104.615
R614 source.n546 source.n545 104.615
R615 source.n545 source.n439 104.615
R616 source.n443 source.n439 104.615
R617 source.n537 source.n443 104.615
R618 source.n537 source.n536 104.615
R619 source.n536 source.n444 104.615
R620 source.n529 source.n444 104.615
R621 source.n529 source.n528 104.615
R622 source.n528 source.n448 104.615
R623 source.n521 source.n448 104.615
R624 source.n521 source.n520 104.615
R625 source.n520 source.n452 104.615
R626 source.n513 source.n452 104.615
R627 source.n513 source.n512 104.615
R628 source.n512 source.n456 104.615
R629 source.n505 source.n456 104.615
R630 source.n505 source.n504 104.615
R631 source.n504 source.n460 104.615
R632 source.n497 source.n460 104.615
R633 source.n497 source.n496 104.615
R634 source.n496 source.n495 104.615
R635 source.n495 source.n464 104.615
R636 source.n488 source.n464 104.615
R637 source.n488 source.n487 104.615
R638 source.n487 source.n469 104.615
R639 source.n480 source.n469 104.615
R640 source.n480 source.n479 104.615
R641 source.n479 source.n473 104.615
R642 source.t12 source.n1039 52.3082
R643 source.t20 source.n895 52.3082
R644 source.t6 source.n755 52.3082
R645 source.t10 source.n611 52.3082
R646 source.t2 source.n45 52.3082
R647 source.t9 source.n189 52.3082
R648 source.t17 source.n329 52.3082
R649 source.t23 source.n473 52.3082
R650 source.n995 source.n994 42.0366
R651 source.n993 source.n992 42.0366
R652 source.n711 source.n710 42.0366
R653 source.n709 source.n708 42.0366
R654 source.n141 source.n140 42.0366
R655 source.n143 source.n142 42.0366
R656 source.n425 source.n424 42.0366
R657 source.n427 source.n426 42.0366
R658 source.n707 source.n567 31.6793
R659 source.n1135 source.n1134 30.6338
R660 source.n991 source.n990 30.6338
R661 source.n851 source.n850 30.6338
R662 source.n707 source.n706 30.6338
R663 source.n139 source.n138 30.6338
R664 source.n283 source.n282 30.6338
R665 source.n423 source.n422 30.6338
R666 source.n567 source.n566 30.6338
R667 source.n1136 source.n139 26.1448
R668 source.n1065 source.n1030 13.1884
R669 source.n1112 source.n1111 13.1884
R670 source.n921 source.n886 13.1884
R671 source.n968 source.n967 13.1884
R672 source.n781 source.n746 13.1884
R673 source.n828 source.n827 13.1884
R674 source.n637 source.n602 13.1884
R675 source.n684 source.n683 13.1884
R676 source.n116 source.n115 13.1884
R677 source.n70 source.n35 13.1884
R678 source.n260 source.n259 13.1884
R679 source.n214 source.n179 13.1884
R680 source.n400 source.n399 13.1884
R681 source.n354 source.n319 13.1884
R682 source.n544 source.n543 13.1884
R683 source.n498 source.n463 13.1884
R684 source.n1061 source.n1060 12.8005
R685 source.n1066 source.n1028 12.8005
R686 source.n1110 source.n1008 12.8005
R687 source.n1115 source.n1006 12.8005
R688 source.n917 source.n916 12.8005
R689 source.n922 source.n884 12.8005
R690 source.n966 source.n864 12.8005
R691 source.n971 source.n862 12.8005
R692 source.n777 source.n776 12.8005
R693 source.n782 source.n744 12.8005
R694 source.n826 source.n724 12.8005
R695 source.n831 source.n722 12.8005
R696 source.n633 source.n632 12.8005
R697 source.n638 source.n600 12.8005
R698 source.n682 source.n580 12.8005
R699 source.n687 source.n578 12.8005
R700 source.n119 source.n10 12.8005
R701 source.n114 source.n12 12.8005
R702 source.n71 source.n33 12.8005
R703 source.n66 source.n37 12.8005
R704 source.n263 source.n154 12.8005
R705 source.n258 source.n156 12.8005
R706 source.n215 source.n177 12.8005
R707 source.n210 source.n181 12.8005
R708 source.n403 source.n294 12.8005
R709 source.n398 source.n296 12.8005
R710 source.n355 source.n317 12.8005
R711 source.n350 source.n321 12.8005
R712 source.n547 source.n438 12.8005
R713 source.n542 source.n440 12.8005
R714 source.n499 source.n461 12.8005
R715 source.n494 source.n465 12.8005
R716 source.n1059 source.n1032 12.0247
R717 source.n1070 source.n1069 12.0247
R718 source.n1107 source.n1106 12.0247
R719 source.n1116 source.n1004 12.0247
R720 source.n915 source.n888 12.0247
R721 source.n926 source.n925 12.0247
R722 source.n963 source.n962 12.0247
R723 source.n972 source.n860 12.0247
R724 source.n775 source.n748 12.0247
R725 source.n786 source.n785 12.0247
R726 source.n823 source.n822 12.0247
R727 source.n832 source.n720 12.0247
R728 source.n631 source.n604 12.0247
R729 source.n642 source.n641 12.0247
R730 source.n679 source.n678 12.0247
R731 source.n688 source.n576 12.0247
R732 source.n120 source.n8 12.0247
R733 source.n111 source.n110 12.0247
R734 source.n75 source.n74 12.0247
R735 source.n65 source.n38 12.0247
R736 source.n264 source.n152 12.0247
R737 source.n255 source.n254 12.0247
R738 source.n219 source.n218 12.0247
R739 source.n209 source.n182 12.0247
R740 source.n404 source.n292 12.0247
R741 source.n395 source.n394 12.0247
R742 source.n359 source.n358 12.0247
R743 source.n349 source.n322 12.0247
R744 source.n548 source.n436 12.0247
R745 source.n539 source.n538 12.0247
R746 source.n503 source.n502 12.0247
R747 source.n493 source.n466 12.0247
R748 source.n1056 source.n1055 11.249
R749 source.n1073 source.n1026 11.249
R750 source.n1102 source.n1010 11.249
R751 source.n1120 source.n1119 11.249
R752 source.n912 source.n911 11.249
R753 source.n929 source.n882 11.249
R754 source.n958 source.n866 11.249
R755 source.n976 source.n975 11.249
R756 source.n772 source.n771 11.249
R757 source.n789 source.n742 11.249
R758 source.n818 source.n726 11.249
R759 source.n836 source.n835 11.249
R760 source.n628 source.n627 11.249
R761 source.n645 source.n598 11.249
R762 source.n674 source.n582 11.249
R763 source.n692 source.n691 11.249
R764 source.n124 source.n123 11.249
R765 source.n107 source.n14 11.249
R766 source.n78 source.n31 11.249
R767 source.n62 source.n61 11.249
R768 source.n268 source.n267 11.249
R769 source.n251 source.n158 11.249
R770 source.n222 source.n175 11.249
R771 source.n206 source.n205 11.249
R772 source.n408 source.n407 11.249
R773 source.n391 source.n298 11.249
R774 source.n362 source.n315 11.249
R775 source.n346 source.n345 11.249
R776 source.n552 source.n551 11.249
R777 source.n535 source.n442 11.249
R778 source.n506 source.n459 11.249
R779 source.n490 source.n489 11.249
R780 source.n1052 source.n1034 10.4732
R781 source.n1074 source.n1024 10.4732
R782 source.n1101 source.n1012 10.4732
R783 source.n1123 source.n1002 10.4732
R784 source.n908 source.n890 10.4732
R785 source.n930 source.n880 10.4732
R786 source.n957 source.n868 10.4732
R787 source.n979 source.n858 10.4732
R788 source.n768 source.n750 10.4732
R789 source.n790 source.n740 10.4732
R790 source.n817 source.n728 10.4732
R791 source.n839 source.n718 10.4732
R792 source.n624 source.n606 10.4732
R793 source.n646 source.n596 10.4732
R794 source.n673 source.n584 10.4732
R795 source.n695 source.n574 10.4732
R796 source.n127 source.n6 10.4732
R797 source.n106 source.n17 10.4732
R798 source.n79 source.n29 10.4732
R799 source.n58 source.n40 10.4732
R800 source.n271 source.n150 10.4732
R801 source.n250 source.n161 10.4732
R802 source.n223 source.n173 10.4732
R803 source.n202 source.n184 10.4732
R804 source.n411 source.n290 10.4732
R805 source.n390 source.n301 10.4732
R806 source.n363 source.n313 10.4732
R807 source.n342 source.n324 10.4732
R808 source.n555 source.n434 10.4732
R809 source.n534 source.n445 10.4732
R810 source.n507 source.n457 10.4732
R811 source.n486 source.n468 10.4732
R812 source.n1041 source.n1040 10.2747
R813 source.n897 source.n896 10.2747
R814 source.n757 source.n756 10.2747
R815 source.n613 source.n612 10.2747
R816 source.n47 source.n46 10.2747
R817 source.n191 source.n190 10.2747
R818 source.n331 source.n330 10.2747
R819 source.n475 source.n474 10.2747
R820 source.n1051 source.n1036 9.69747
R821 source.n1078 source.n1077 9.69747
R822 source.n1098 source.n1097 9.69747
R823 source.n1124 source.n1000 9.69747
R824 source.n907 source.n892 9.69747
R825 source.n934 source.n933 9.69747
R826 source.n954 source.n953 9.69747
R827 source.n980 source.n856 9.69747
R828 source.n767 source.n752 9.69747
R829 source.n794 source.n793 9.69747
R830 source.n814 source.n813 9.69747
R831 source.n840 source.n716 9.69747
R832 source.n623 source.n608 9.69747
R833 source.n650 source.n649 9.69747
R834 source.n670 source.n669 9.69747
R835 source.n696 source.n572 9.69747
R836 source.n128 source.n4 9.69747
R837 source.n103 source.n102 9.69747
R838 source.n83 source.n82 9.69747
R839 source.n57 source.n42 9.69747
R840 source.n272 source.n148 9.69747
R841 source.n247 source.n246 9.69747
R842 source.n227 source.n226 9.69747
R843 source.n201 source.n186 9.69747
R844 source.n412 source.n288 9.69747
R845 source.n387 source.n386 9.69747
R846 source.n367 source.n366 9.69747
R847 source.n341 source.n326 9.69747
R848 source.n556 source.n432 9.69747
R849 source.n531 source.n530 9.69747
R850 source.n511 source.n510 9.69747
R851 source.n485 source.n470 9.69747
R852 source.n1134 source.n1133 9.45567
R853 source.n990 source.n989 9.45567
R854 source.n850 source.n849 9.45567
R855 source.n706 source.n705 9.45567
R856 source.n138 source.n137 9.45567
R857 source.n282 source.n281 9.45567
R858 source.n422 source.n421 9.45567
R859 source.n566 source.n565 9.45567
R860 source.n998 source.n997 9.3005
R861 source.n1127 source.n1126 9.3005
R862 source.n1125 source.n1124 9.3005
R863 source.n1002 source.n1001 9.3005
R864 source.n1119 source.n1118 9.3005
R865 source.n1117 source.n1116 9.3005
R866 source.n1006 source.n1005 9.3005
R867 source.n1085 source.n1084 9.3005
R868 source.n1083 source.n1082 9.3005
R869 source.n1022 source.n1021 9.3005
R870 source.n1077 source.n1076 9.3005
R871 source.n1075 source.n1074 9.3005
R872 source.n1026 source.n1025 9.3005
R873 source.n1069 source.n1068 9.3005
R874 source.n1067 source.n1066 9.3005
R875 source.n1043 source.n1042 9.3005
R876 source.n1038 source.n1037 9.3005
R877 source.n1049 source.n1048 9.3005
R878 source.n1051 source.n1050 9.3005
R879 source.n1034 source.n1033 9.3005
R880 source.n1057 source.n1056 9.3005
R881 source.n1059 source.n1058 9.3005
R882 source.n1060 source.n1029 9.3005
R883 source.n1018 source.n1017 9.3005
R884 source.n1091 source.n1090 9.3005
R885 source.n1093 source.n1092 9.3005
R886 source.n1014 source.n1013 9.3005
R887 source.n1099 source.n1098 9.3005
R888 source.n1101 source.n1100 9.3005
R889 source.n1010 source.n1009 9.3005
R890 source.n1108 source.n1107 9.3005
R891 source.n1110 source.n1109 9.3005
R892 source.n1133 source.n1132 9.3005
R893 source.n854 source.n853 9.3005
R894 source.n983 source.n982 9.3005
R895 source.n981 source.n980 9.3005
R896 source.n858 source.n857 9.3005
R897 source.n975 source.n974 9.3005
R898 source.n973 source.n972 9.3005
R899 source.n862 source.n861 9.3005
R900 source.n941 source.n940 9.3005
R901 source.n939 source.n938 9.3005
R902 source.n878 source.n877 9.3005
R903 source.n933 source.n932 9.3005
R904 source.n931 source.n930 9.3005
R905 source.n882 source.n881 9.3005
R906 source.n925 source.n924 9.3005
R907 source.n923 source.n922 9.3005
R908 source.n899 source.n898 9.3005
R909 source.n894 source.n893 9.3005
R910 source.n905 source.n904 9.3005
R911 source.n907 source.n906 9.3005
R912 source.n890 source.n889 9.3005
R913 source.n913 source.n912 9.3005
R914 source.n915 source.n914 9.3005
R915 source.n916 source.n885 9.3005
R916 source.n874 source.n873 9.3005
R917 source.n947 source.n946 9.3005
R918 source.n949 source.n948 9.3005
R919 source.n870 source.n869 9.3005
R920 source.n955 source.n954 9.3005
R921 source.n957 source.n956 9.3005
R922 source.n866 source.n865 9.3005
R923 source.n964 source.n963 9.3005
R924 source.n966 source.n965 9.3005
R925 source.n989 source.n988 9.3005
R926 source.n714 source.n713 9.3005
R927 source.n843 source.n842 9.3005
R928 source.n841 source.n840 9.3005
R929 source.n718 source.n717 9.3005
R930 source.n835 source.n834 9.3005
R931 source.n833 source.n832 9.3005
R932 source.n722 source.n721 9.3005
R933 source.n801 source.n800 9.3005
R934 source.n799 source.n798 9.3005
R935 source.n738 source.n737 9.3005
R936 source.n793 source.n792 9.3005
R937 source.n791 source.n790 9.3005
R938 source.n742 source.n741 9.3005
R939 source.n785 source.n784 9.3005
R940 source.n783 source.n782 9.3005
R941 source.n759 source.n758 9.3005
R942 source.n754 source.n753 9.3005
R943 source.n765 source.n764 9.3005
R944 source.n767 source.n766 9.3005
R945 source.n750 source.n749 9.3005
R946 source.n773 source.n772 9.3005
R947 source.n775 source.n774 9.3005
R948 source.n776 source.n745 9.3005
R949 source.n734 source.n733 9.3005
R950 source.n807 source.n806 9.3005
R951 source.n809 source.n808 9.3005
R952 source.n730 source.n729 9.3005
R953 source.n815 source.n814 9.3005
R954 source.n817 source.n816 9.3005
R955 source.n726 source.n725 9.3005
R956 source.n824 source.n823 9.3005
R957 source.n826 source.n825 9.3005
R958 source.n849 source.n848 9.3005
R959 source.n570 source.n569 9.3005
R960 source.n699 source.n698 9.3005
R961 source.n697 source.n696 9.3005
R962 source.n574 source.n573 9.3005
R963 source.n691 source.n690 9.3005
R964 source.n689 source.n688 9.3005
R965 source.n578 source.n577 9.3005
R966 source.n657 source.n656 9.3005
R967 source.n655 source.n654 9.3005
R968 source.n594 source.n593 9.3005
R969 source.n649 source.n648 9.3005
R970 source.n647 source.n646 9.3005
R971 source.n598 source.n597 9.3005
R972 source.n641 source.n640 9.3005
R973 source.n639 source.n638 9.3005
R974 source.n615 source.n614 9.3005
R975 source.n610 source.n609 9.3005
R976 source.n621 source.n620 9.3005
R977 source.n623 source.n622 9.3005
R978 source.n606 source.n605 9.3005
R979 source.n629 source.n628 9.3005
R980 source.n631 source.n630 9.3005
R981 source.n632 source.n601 9.3005
R982 source.n590 source.n589 9.3005
R983 source.n663 source.n662 9.3005
R984 source.n665 source.n664 9.3005
R985 source.n586 source.n585 9.3005
R986 source.n671 source.n670 9.3005
R987 source.n673 source.n672 9.3005
R988 source.n582 source.n581 9.3005
R989 source.n680 source.n679 9.3005
R990 source.n682 source.n681 9.3005
R991 source.n705 source.n704 9.3005
R992 source.n49 source.n48 9.3005
R993 source.n44 source.n43 9.3005
R994 source.n55 source.n54 9.3005
R995 source.n57 source.n56 9.3005
R996 source.n40 source.n39 9.3005
R997 source.n63 source.n62 9.3005
R998 source.n65 source.n64 9.3005
R999 source.n37 source.n34 9.3005
R1000 source.n96 source.n95 9.3005
R1001 source.n98 source.n97 9.3005
R1002 source.n19 source.n18 9.3005
R1003 source.n104 source.n103 9.3005
R1004 source.n106 source.n105 9.3005
R1005 source.n14 source.n13 9.3005
R1006 source.n112 source.n111 9.3005
R1007 source.n114 source.n113 9.3005
R1008 source.n137 source.n136 9.3005
R1009 source.n2 source.n1 9.3005
R1010 source.n131 source.n130 9.3005
R1011 source.n129 source.n128 9.3005
R1012 source.n6 source.n5 9.3005
R1013 source.n123 source.n122 9.3005
R1014 source.n121 source.n120 9.3005
R1015 source.n10 source.n9 9.3005
R1016 source.n23 source.n22 9.3005
R1017 source.n90 source.n89 9.3005
R1018 source.n88 source.n87 9.3005
R1019 source.n27 source.n26 9.3005
R1020 source.n82 source.n81 9.3005
R1021 source.n80 source.n79 9.3005
R1022 source.n31 source.n30 9.3005
R1023 source.n74 source.n73 9.3005
R1024 source.n72 source.n71 9.3005
R1025 source.n193 source.n192 9.3005
R1026 source.n188 source.n187 9.3005
R1027 source.n199 source.n198 9.3005
R1028 source.n201 source.n200 9.3005
R1029 source.n184 source.n183 9.3005
R1030 source.n207 source.n206 9.3005
R1031 source.n209 source.n208 9.3005
R1032 source.n181 source.n178 9.3005
R1033 source.n240 source.n239 9.3005
R1034 source.n242 source.n241 9.3005
R1035 source.n163 source.n162 9.3005
R1036 source.n248 source.n247 9.3005
R1037 source.n250 source.n249 9.3005
R1038 source.n158 source.n157 9.3005
R1039 source.n256 source.n255 9.3005
R1040 source.n258 source.n257 9.3005
R1041 source.n281 source.n280 9.3005
R1042 source.n146 source.n145 9.3005
R1043 source.n275 source.n274 9.3005
R1044 source.n273 source.n272 9.3005
R1045 source.n150 source.n149 9.3005
R1046 source.n267 source.n266 9.3005
R1047 source.n265 source.n264 9.3005
R1048 source.n154 source.n153 9.3005
R1049 source.n167 source.n166 9.3005
R1050 source.n234 source.n233 9.3005
R1051 source.n232 source.n231 9.3005
R1052 source.n171 source.n170 9.3005
R1053 source.n226 source.n225 9.3005
R1054 source.n224 source.n223 9.3005
R1055 source.n175 source.n174 9.3005
R1056 source.n218 source.n217 9.3005
R1057 source.n216 source.n215 9.3005
R1058 source.n333 source.n332 9.3005
R1059 source.n328 source.n327 9.3005
R1060 source.n339 source.n338 9.3005
R1061 source.n341 source.n340 9.3005
R1062 source.n324 source.n323 9.3005
R1063 source.n347 source.n346 9.3005
R1064 source.n349 source.n348 9.3005
R1065 source.n321 source.n318 9.3005
R1066 source.n380 source.n379 9.3005
R1067 source.n382 source.n381 9.3005
R1068 source.n303 source.n302 9.3005
R1069 source.n388 source.n387 9.3005
R1070 source.n390 source.n389 9.3005
R1071 source.n298 source.n297 9.3005
R1072 source.n396 source.n395 9.3005
R1073 source.n398 source.n397 9.3005
R1074 source.n421 source.n420 9.3005
R1075 source.n286 source.n285 9.3005
R1076 source.n415 source.n414 9.3005
R1077 source.n413 source.n412 9.3005
R1078 source.n290 source.n289 9.3005
R1079 source.n407 source.n406 9.3005
R1080 source.n405 source.n404 9.3005
R1081 source.n294 source.n293 9.3005
R1082 source.n307 source.n306 9.3005
R1083 source.n374 source.n373 9.3005
R1084 source.n372 source.n371 9.3005
R1085 source.n311 source.n310 9.3005
R1086 source.n366 source.n365 9.3005
R1087 source.n364 source.n363 9.3005
R1088 source.n315 source.n314 9.3005
R1089 source.n358 source.n357 9.3005
R1090 source.n356 source.n355 9.3005
R1091 source.n477 source.n476 9.3005
R1092 source.n472 source.n471 9.3005
R1093 source.n483 source.n482 9.3005
R1094 source.n485 source.n484 9.3005
R1095 source.n468 source.n467 9.3005
R1096 source.n491 source.n490 9.3005
R1097 source.n493 source.n492 9.3005
R1098 source.n465 source.n462 9.3005
R1099 source.n524 source.n523 9.3005
R1100 source.n526 source.n525 9.3005
R1101 source.n447 source.n446 9.3005
R1102 source.n532 source.n531 9.3005
R1103 source.n534 source.n533 9.3005
R1104 source.n442 source.n441 9.3005
R1105 source.n540 source.n539 9.3005
R1106 source.n542 source.n541 9.3005
R1107 source.n565 source.n564 9.3005
R1108 source.n430 source.n429 9.3005
R1109 source.n559 source.n558 9.3005
R1110 source.n557 source.n556 9.3005
R1111 source.n434 source.n433 9.3005
R1112 source.n551 source.n550 9.3005
R1113 source.n549 source.n548 9.3005
R1114 source.n438 source.n437 9.3005
R1115 source.n451 source.n450 9.3005
R1116 source.n518 source.n517 9.3005
R1117 source.n516 source.n515 9.3005
R1118 source.n455 source.n454 9.3005
R1119 source.n510 source.n509 9.3005
R1120 source.n508 source.n507 9.3005
R1121 source.n459 source.n458 9.3005
R1122 source.n502 source.n501 9.3005
R1123 source.n500 source.n499 9.3005
R1124 source.n1048 source.n1047 8.92171
R1125 source.n1081 source.n1022 8.92171
R1126 source.n1094 source.n1014 8.92171
R1127 source.n1128 source.n1127 8.92171
R1128 source.n904 source.n903 8.92171
R1129 source.n937 source.n878 8.92171
R1130 source.n950 source.n870 8.92171
R1131 source.n984 source.n983 8.92171
R1132 source.n764 source.n763 8.92171
R1133 source.n797 source.n738 8.92171
R1134 source.n810 source.n730 8.92171
R1135 source.n844 source.n843 8.92171
R1136 source.n620 source.n619 8.92171
R1137 source.n653 source.n594 8.92171
R1138 source.n666 source.n586 8.92171
R1139 source.n700 source.n699 8.92171
R1140 source.n132 source.n131 8.92171
R1141 source.n99 source.n19 8.92171
R1142 source.n86 source.n27 8.92171
R1143 source.n54 source.n53 8.92171
R1144 source.n276 source.n275 8.92171
R1145 source.n243 source.n163 8.92171
R1146 source.n230 source.n171 8.92171
R1147 source.n198 source.n197 8.92171
R1148 source.n416 source.n415 8.92171
R1149 source.n383 source.n303 8.92171
R1150 source.n370 source.n311 8.92171
R1151 source.n338 source.n337 8.92171
R1152 source.n560 source.n559 8.92171
R1153 source.n527 source.n447 8.92171
R1154 source.n514 source.n455 8.92171
R1155 source.n482 source.n481 8.92171
R1156 source.n1044 source.n1038 8.14595
R1157 source.n1082 source.n1020 8.14595
R1158 source.n1093 source.n1016 8.14595
R1159 source.n1131 source.n998 8.14595
R1160 source.n900 source.n894 8.14595
R1161 source.n938 source.n876 8.14595
R1162 source.n949 source.n872 8.14595
R1163 source.n987 source.n854 8.14595
R1164 source.n760 source.n754 8.14595
R1165 source.n798 source.n736 8.14595
R1166 source.n809 source.n732 8.14595
R1167 source.n847 source.n714 8.14595
R1168 source.n616 source.n610 8.14595
R1169 source.n654 source.n592 8.14595
R1170 source.n665 source.n588 8.14595
R1171 source.n703 source.n570 8.14595
R1172 source.n135 source.n2 8.14595
R1173 source.n98 source.n21 8.14595
R1174 source.n87 source.n25 8.14595
R1175 source.n50 source.n44 8.14595
R1176 source.n279 source.n146 8.14595
R1177 source.n242 source.n165 8.14595
R1178 source.n231 source.n169 8.14595
R1179 source.n194 source.n188 8.14595
R1180 source.n419 source.n286 8.14595
R1181 source.n382 source.n305 8.14595
R1182 source.n371 source.n309 8.14595
R1183 source.n334 source.n328 8.14595
R1184 source.n563 source.n430 8.14595
R1185 source.n526 source.n449 8.14595
R1186 source.n515 source.n453 8.14595
R1187 source.n478 source.n472 8.14595
R1188 source.n1043 source.n1040 7.3702
R1189 source.n1086 source.n1085 7.3702
R1190 source.n1090 source.n1089 7.3702
R1191 source.n1132 source.n996 7.3702
R1192 source.n899 source.n896 7.3702
R1193 source.n942 source.n941 7.3702
R1194 source.n946 source.n945 7.3702
R1195 source.n988 source.n852 7.3702
R1196 source.n759 source.n756 7.3702
R1197 source.n802 source.n801 7.3702
R1198 source.n806 source.n805 7.3702
R1199 source.n848 source.n712 7.3702
R1200 source.n615 source.n612 7.3702
R1201 source.n658 source.n657 7.3702
R1202 source.n662 source.n661 7.3702
R1203 source.n704 source.n568 7.3702
R1204 source.n136 source.n0 7.3702
R1205 source.n95 source.n94 7.3702
R1206 source.n91 source.n90 7.3702
R1207 source.n49 source.n46 7.3702
R1208 source.n280 source.n144 7.3702
R1209 source.n239 source.n238 7.3702
R1210 source.n235 source.n234 7.3702
R1211 source.n193 source.n190 7.3702
R1212 source.n420 source.n284 7.3702
R1213 source.n379 source.n378 7.3702
R1214 source.n375 source.n374 7.3702
R1215 source.n333 source.n330 7.3702
R1216 source.n564 source.n428 7.3702
R1217 source.n523 source.n522 7.3702
R1218 source.n519 source.n518 7.3702
R1219 source.n477 source.n474 7.3702
R1220 source.n1086 source.n1018 6.59444
R1221 source.n1089 source.n1018 6.59444
R1222 source.n1134 source.n996 6.59444
R1223 source.n942 source.n874 6.59444
R1224 source.n945 source.n874 6.59444
R1225 source.n990 source.n852 6.59444
R1226 source.n802 source.n734 6.59444
R1227 source.n805 source.n734 6.59444
R1228 source.n850 source.n712 6.59444
R1229 source.n658 source.n590 6.59444
R1230 source.n661 source.n590 6.59444
R1231 source.n706 source.n568 6.59444
R1232 source.n138 source.n0 6.59444
R1233 source.n94 source.n23 6.59444
R1234 source.n91 source.n23 6.59444
R1235 source.n282 source.n144 6.59444
R1236 source.n238 source.n167 6.59444
R1237 source.n235 source.n167 6.59444
R1238 source.n422 source.n284 6.59444
R1239 source.n378 source.n307 6.59444
R1240 source.n375 source.n307 6.59444
R1241 source.n566 source.n428 6.59444
R1242 source.n522 source.n451 6.59444
R1243 source.n519 source.n451 6.59444
R1244 source.n1044 source.n1043 5.81868
R1245 source.n1085 source.n1020 5.81868
R1246 source.n1090 source.n1016 5.81868
R1247 source.n1132 source.n1131 5.81868
R1248 source.n900 source.n899 5.81868
R1249 source.n941 source.n876 5.81868
R1250 source.n946 source.n872 5.81868
R1251 source.n988 source.n987 5.81868
R1252 source.n760 source.n759 5.81868
R1253 source.n801 source.n736 5.81868
R1254 source.n806 source.n732 5.81868
R1255 source.n848 source.n847 5.81868
R1256 source.n616 source.n615 5.81868
R1257 source.n657 source.n592 5.81868
R1258 source.n662 source.n588 5.81868
R1259 source.n704 source.n703 5.81868
R1260 source.n136 source.n135 5.81868
R1261 source.n95 source.n21 5.81868
R1262 source.n90 source.n25 5.81868
R1263 source.n50 source.n49 5.81868
R1264 source.n280 source.n279 5.81868
R1265 source.n239 source.n165 5.81868
R1266 source.n234 source.n169 5.81868
R1267 source.n194 source.n193 5.81868
R1268 source.n420 source.n419 5.81868
R1269 source.n379 source.n305 5.81868
R1270 source.n374 source.n309 5.81868
R1271 source.n334 source.n333 5.81868
R1272 source.n564 source.n563 5.81868
R1273 source.n523 source.n449 5.81868
R1274 source.n518 source.n453 5.81868
R1275 source.n478 source.n477 5.81868
R1276 source.n1136 source.n1135 5.53498
R1277 source.n1047 source.n1038 5.04292
R1278 source.n1082 source.n1081 5.04292
R1279 source.n1094 source.n1093 5.04292
R1280 source.n1128 source.n998 5.04292
R1281 source.n903 source.n894 5.04292
R1282 source.n938 source.n937 5.04292
R1283 source.n950 source.n949 5.04292
R1284 source.n984 source.n854 5.04292
R1285 source.n763 source.n754 5.04292
R1286 source.n798 source.n797 5.04292
R1287 source.n810 source.n809 5.04292
R1288 source.n844 source.n714 5.04292
R1289 source.n619 source.n610 5.04292
R1290 source.n654 source.n653 5.04292
R1291 source.n666 source.n665 5.04292
R1292 source.n700 source.n570 5.04292
R1293 source.n132 source.n2 5.04292
R1294 source.n99 source.n98 5.04292
R1295 source.n87 source.n86 5.04292
R1296 source.n53 source.n44 5.04292
R1297 source.n276 source.n146 5.04292
R1298 source.n243 source.n242 5.04292
R1299 source.n231 source.n230 5.04292
R1300 source.n197 source.n188 5.04292
R1301 source.n416 source.n286 5.04292
R1302 source.n383 source.n382 5.04292
R1303 source.n371 source.n370 5.04292
R1304 source.n337 source.n328 5.04292
R1305 source.n560 source.n430 5.04292
R1306 source.n527 source.n526 5.04292
R1307 source.n515 source.n514 5.04292
R1308 source.n481 source.n472 5.04292
R1309 source.n1048 source.n1036 4.26717
R1310 source.n1078 source.n1022 4.26717
R1311 source.n1097 source.n1014 4.26717
R1312 source.n1127 source.n1000 4.26717
R1313 source.n904 source.n892 4.26717
R1314 source.n934 source.n878 4.26717
R1315 source.n953 source.n870 4.26717
R1316 source.n983 source.n856 4.26717
R1317 source.n764 source.n752 4.26717
R1318 source.n794 source.n738 4.26717
R1319 source.n813 source.n730 4.26717
R1320 source.n843 source.n716 4.26717
R1321 source.n620 source.n608 4.26717
R1322 source.n650 source.n594 4.26717
R1323 source.n669 source.n586 4.26717
R1324 source.n699 source.n572 4.26717
R1325 source.n131 source.n4 4.26717
R1326 source.n102 source.n19 4.26717
R1327 source.n83 source.n27 4.26717
R1328 source.n54 source.n42 4.26717
R1329 source.n275 source.n148 4.26717
R1330 source.n246 source.n163 4.26717
R1331 source.n227 source.n171 4.26717
R1332 source.n198 source.n186 4.26717
R1333 source.n415 source.n288 4.26717
R1334 source.n386 source.n303 4.26717
R1335 source.n367 source.n311 4.26717
R1336 source.n338 source.n326 4.26717
R1337 source.n559 source.n432 4.26717
R1338 source.n530 source.n447 4.26717
R1339 source.n511 source.n455 4.26717
R1340 source.n482 source.n470 4.26717
R1341 source.n1052 source.n1051 3.49141
R1342 source.n1077 source.n1024 3.49141
R1343 source.n1098 source.n1012 3.49141
R1344 source.n1124 source.n1123 3.49141
R1345 source.n908 source.n907 3.49141
R1346 source.n933 source.n880 3.49141
R1347 source.n954 source.n868 3.49141
R1348 source.n980 source.n979 3.49141
R1349 source.n768 source.n767 3.49141
R1350 source.n793 source.n740 3.49141
R1351 source.n814 source.n728 3.49141
R1352 source.n840 source.n839 3.49141
R1353 source.n624 source.n623 3.49141
R1354 source.n649 source.n596 3.49141
R1355 source.n670 source.n584 3.49141
R1356 source.n696 source.n695 3.49141
R1357 source.n128 source.n127 3.49141
R1358 source.n103 source.n17 3.49141
R1359 source.n82 source.n29 3.49141
R1360 source.n58 source.n57 3.49141
R1361 source.n272 source.n271 3.49141
R1362 source.n247 source.n161 3.49141
R1363 source.n226 source.n173 3.49141
R1364 source.n202 source.n201 3.49141
R1365 source.n412 source.n411 3.49141
R1366 source.n387 source.n301 3.49141
R1367 source.n366 source.n313 3.49141
R1368 source.n342 source.n341 3.49141
R1369 source.n556 source.n555 3.49141
R1370 source.n531 source.n445 3.49141
R1371 source.n510 source.n457 3.49141
R1372 source.n486 source.n485 3.49141
R1373 source.n48 source.n47 2.84303
R1374 source.n192 source.n191 2.84303
R1375 source.n332 source.n331 2.84303
R1376 source.n476 source.n475 2.84303
R1377 source.n1042 source.n1041 2.84303
R1378 source.n898 source.n897 2.84303
R1379 source.n758 source.n757 2.84303
R1380 source.n614 source.n613 2.84303
R1381 source.n1055 source.n1034 2.71565
R1382 source.n1074 source.n1073 2.71565
R1383 source.n1102 source.n1101 2.71565
R1384 source.n1120 source.n1002 2.71565
R1385 source.n911 source.n890 2.71565
R1386 source.n930 source.n929 2.71565
R1387 source.n958 source.n957 2.71565
R1388 source.n976 source.n858 2.71565
R1389 source.n771 source.n750 2.71565
R1390 source.n790 source.n789 2.71565
R1391 source.n818 source.n817 2.71565
R1392 source.n836 source.n718 2.71565
R1393 source.n627 source.n606 2.71565
R1394 source.n646 source.n645 2.71565
R1395 source.n674 source.n673 2.71565
R1396 source.n692 source.n574 2.71565
R1397 source.n124 source.n6 2.71565
R1398 source.n107 source.n106 2.71565
R1399 source.n79 source.n78 2.71565
R1400 source.n61 source.n40 2.71565
R1401 source.n268 source.n150 2.71565
R1402 source.n251 source.n250 2.71565
R1403 source.n223 source.n222 2.71565
R1404 source.n205 source.n184 2.71565
R1405 source.n408 source.n290 2.71565
R1406 source.n391 source.n390 2.71565
R1407 source.n363 source.n362 2.71565
R1408 source.n345 source.n324 2.71565
R1409 source.n552 source.n434 2.71565
R1410 source.n535 source.n534 2.71565
R1411 source.n507 source.n506 2.71565
R1412 source.n489 source.n468 2.71565
R1413 source.n1056 source.n1032 1.93989
R1414 source.n1070 source.n1026 1.93989
R1415 source.n1106 source.n1010 1.93989
R1416 source.n1119 source.n1004 1.93989
R1417 source.n912 source.n888 1.93989
R1418 source.n926 source.n882 1.93989
R1419 source.n962 source.n866 1.93989
R1420 source.n975 source.n860 1.93989
R1421 source.n772 source.n748 1.93989
R1422 source.n786 source.n742 1.93989
R1423 source.n822 source.n726 1.93989
R1424 source.n835 source.n720 1.93989
R1425 source.n628 source.n604 1.93989
R1426 source.n642 source.n598 1.93989
R1427 source.n678 source.n582 1.93989
R1428 source.n691 source.n576 1.93989
R1429 source.n123 source.n8 1.93989
R1430 source.n110 source.n14 1.93989
R1431 source.n75 source.n31 1.93989
R1432 source.n62 source.n38 1.93989
R1433 source.n267 source.n152 1.93989
R1434 source.n254 source.n158 1.93989
R1435 source.n219 source.n175 1.93989
R1436 source.n206 source.n182 1.93989
R1437 source.n407 source.n292 1.93989
R1438 source.n394 source.n298 1.93989
R1439 source.n359 source.n315 1.93989
R1440 source.n346 source.n322 1.93989
R1441 source.n551 source.n436 1.93989
R1442 source.n538 source.n442 1.93989
R1443 source.n503 source.n459 1.93989
R1444 source.n490 source.n466 1.93989
R1445 source.n1061 source.n1059 1.16414
R1446 source.n1069 source.n1028 1.16414
R1447 source.n1107 source.n1008 1.16414
R1448 source.n1116 source.n1115 1.16414
R1449 source.n917 source.n915 1.16414
R1450 source.n925 source.n884 1.16414
R1451 source.n963 source.n864 1.16414
R1452 source.n972 source.n971 1.16414
R1453 source.n777 source.n775 1.16414
R1454 source.n785 source.n744 1.16414
R1455 source.n823 source.n724 1.16414
R1456 source.n832 source.n831 1.16414
R1457 source.n633 source.n631 1.16414
R1458 source.n641 source.n600 1.16414
R1459 source.n679 source.n580 1.16414
R1460 source.n688 source.n687 1.16414
R1461 source.n120 source.n119 1.16414
R1462 source.n111 source.n12 1.16414
R1463 source.n74 source.n33 1.16414
R1464 source.n66 source.n65 1.16414
R1465 source.n264 source.n263 1.16414
R1466 source.n255 source.n156 1.16414
R1467 source.n218 source.n177 1.16414
R1468 source.n210 source.n209 1.16414
R1469 source.n404 source.n403 1.16414
R1470 source.n395 source.n296 1.16414
R1471 source.n358 source.n317 1.16414
R1472 source.n350 source.n349 1.16414
R1473 source.n548 source.n547 1.16414
R1474 source.n539 source.n440 1.16414
R1475 source.n502 source.n461 1.16414
R1476 source.n494 source.n493 1.16414
R1477 source.n994 source.t16 0.7925
R1478 source.n994 source.t19 0.7925
R1479 source.n992 source.t15 0.7925
R1480 source.n992 source.t21 0.7925
R1481 source.n710 source.t5 0.7925
R1482 source.n710 source.t1 0.7925
R1483 source.n708 source.t0 0.7925
R1484 source.n708 source.t3 0.7925
R1485 source.n140 source.t4 0.7925
R1486 source.n140 source.t8 0.7925
R1487 source.n142 source.t11 0.7925
R1488 source.n142 source.t7 0.7925
R1489 source.n424 source.t22 0.7925
R1490 source.n424 source.t13 0.7925
R1491 source.n426 source.t14 0.7925
R1492 source.n426 source.t18 0.7925
R1493 source.n567 source.n427 0.543603
R1494 source.n427 source.n425 0.543603
R1495 source.n425 source.n423 0.543603
R1496 source.n283 source.n143 0.543603
R1497 source.n143 source.n141 0.543603
R1498 source.n141 source.n139 0.543603
R1499 source.n709 source.n707 0.543603
R1500 source.n711 source.n709 0.543603
R1501 source.n851 source.n711 0.543603
R1502 source.n993 source.n991 0.543603
R1503 source.n995 source.n993 0.543603
R1504 source.n1135 source.n995 0.543603
R1505 source.n423 source.n283 0.470328
R1506 source.n991 source.n851 0.470328
R1507 source.n1060 source.n1030 0.388379
R1508 source.n1066 source.n1065 0.388379
R1509 source.n1111 source.n1110 0.388379
R1510 source.n1112 source.n1006 0.388379
R1511 source.n916 source.n886 0.388379
R1512 source.n922 source.n921 0.388379
R1513 source.n967 source.n966 0.388379
R1514 source.n968 source.n862 0.388379
R1515 source.n776 source.n746 0.388379
R1516 source.n782 source.n781 0.388379
R1517 source.n827 source.n826 0.388379
R1518 source.n828 source.n722 0.388379
R1519 source.n632 source.n602 0.388379
R1520 source.n638 source.n637 0.388379
R1521 source.n683 source.n682 0.388379
R1522 source.n684 source.n578 0.388379
R1523 source.n116 source.n10 0.388379
R1524 source.n115 source.n114 0.388379
R1525 source.n71 source.n70 0.388379
R1526 source.n37 source.n35 0.388379
R1527 source.n260 source.n154 0.388379
R1528 source.n259 source.n258 0.388379
R1529 source.n215 source.n214 0.388379
R1530 source.n181 source.n179 0.388379
R1531 source.n400 source.n294 0.388379
R1532 source.n399 source.n398 0.388379
R1533 source.n355 source.n354 0.388379
R1534 source.n321 source.n319 0.388379
R1535 source.n544 source.n438 0.388379
R1536 source.n543 source.n542 0.388379
R1537 source.n499 source.n498 0.388379
R1538 source.n465 source.n463 0.388379
R1539 source source.n1136 0.188
R1540 source.n1042 source.n1037 0.155672
R1541 source.n1049 source.n1037 0.155672
R1542 source.n1050 source.n1049 0.155672
R1543 source.n1050 source.n1033 0.155672
R1544 source.n1057 source.n1033 0.155672
R1545 source.n1058 source.n1057 0.155672
R1546 source.n1058 source.n1029 0.155672
R1547 source.n1067 source.n1029 0.155672
R1548 source.n1068 source.n1067 0.155672
R1549 source.n1068 source.n1025 0.155672
R1550 source.n1075 source.n1025 0.155672
R1551 source.n1076 source.n1075 0.155672
R1552 source.n1076 source.n1021 0.155672
R1553 source.n1083 source.n1021 0.155672
R1554 source.n1084 source.n1083 0.155672
R1555 source.n1084 source.n1017 0.155672
R1556 source.n1091 source.n1017 0.155672
R1557 source.n1092 source.n1091 0.155672
R1558 source.n1092 source.n1013 0.155672
R1559 source.n1099 source.n1013 0.155672
R1560 source.n1100 source.n1099 0.155672
R1561 source.n1100 source.n1009 0.155672
R1562 source.n1108 source.n1009 0.155672
R1563 source.n1109 source.n1108 0.155672
R1564 source.n1109 source.n1005 0.155672
R1565 source.n1117 source.n1005 0.155672
R1566 source.n1118 source.n1117 0.155672
R1567 source.n1118 source.n1001 0.155672
R1568 source.n1125 source.n1001 0.155672
R1569 source.n1126 source.n1125 0.155672
R1570 source.n1126 source.n997 0.155672
R1571 source.n1133 source.n997 0.155672
R1572 source.n898 source.n893 0.155672
R1573 source.n905 source.n893 0.155672
R1574 source.n906 source.n905 0.155672
R1575 source.n906 source.n889 0.155672
R1576 source.n913 source.n889 0.155672
R1577 source.n914 source.n913 0.155672
R1578 source.n914 source.n885 0.155672
R1579 source.n923 source.n885 0.155672
R1580 source.n924 source.n923 0.155672
R1581 source.n924 source.n881 0.155672
R1582 source.n931 source.n881 0.155672
R1583 source.n932 source.n931 0.155672
R1584 source.n932 source.n877 0.155672
R1585 source.n939 source.n877 0.155672
R1586 source.n940 source.n939 0.155672
R1587 source.n940 source.n873 0.155672
R1588 source.n947 source.n873 0.155672
R1589 source.n948 source.n947 0.155672
R1590 source.n948 source.n869 0.155672
R1591 source.n955 source.n869 0.155672
R1592 source.n956 source.n955 0.155672
R1593 source.n956 source.n865 0.155672
R1594 source.n964 source.n865 0.155672
R1595 source.n965 source.n964 0.155672
R1596 source.n965 source.n861 0.155672
R1597 source.n973 source.n861 0.155672
R1598 source.n974 source.n973 0.155672
R1599 source.n974 source.n857 0.155672
R1600 source.n981 source.n857 0.155672
R1601 source.n982 source.n981 0.155672
R1602 source.n982 source.n853 0.155672
R1603 source.n989 source.n853 0.155672
R1604 source.n758 source.n753 0.155672
R1605 source.n765 source.n753 0.155672
R1606 source.n766 source.n765 0.155672
R1607 source.n766 source.n749 0.155672
R1608 source.n773 source.n749 0.155672
R1609 source.n774 source.n773 0.155672
R1610 source.n774 source.n745 0.155672
R1611 source.n783 source.n745 0.155672
R1612 source.n784 source.n783 0.155672
R1613 source.n784 source.n741 0.155672
R1614 source.n791 source.n741 0.155672
R1615 source.n792 source.n791 0.155672
R1616 source.n792 source.n737 0.155672
R1617 source.n799 source.n737 0.155672
R1618 source.n800 source.n799 0.155672
R1619 source.n800 source.n733 0.155672
R1620 source.n807 source.n733 0.155672
R1621 source.n808 source.n807 0.155672
R1622 source.n808 source.n729 0.155672
R1623 source.n815 source.n729 0.155672
R1624 source.n816 source.n815 0.155672
R1625 source.n816 source.n725 0.155672
R1626 source.n824 source.n725 0.155672
R1627 source.n825 source.n824 0.155672
R1628 source.n825 source.n721 0.155672
R1629 source.n833 source.n721 0.155672
R1630 source.n834 source.n833 0.155672
R1631 source.n834 source.n717 0.155672
R1632 source.n841 source.n717 0.155672
R1633 source.n842 source.n841 0.155672
R1634 source.n842 source.n713 0.155672
R1635 source.n849 source.n713 0.155672
R1636 source.n614 source.n609 0.155672
R1637 source.n621 source.n609 0.155672
R1638 source.n622 source.n621 0.155672
R1639 source.n622 source.n605 0.155672
R1640 source.n629 source.n605 0.155672
R1641 source.n630 source.n629 0.155672
R1642 source.n630 source.n601 0.155672
R1643 source.n639 source.n601 0.155672
R1644 source.n640 source.n639 0.155672
R1645 source.n640 source.n597 0.155672
R1646 source.n647 source.n597 0.155672
R1647 source.n648 source.n647 0.155672
R1648 source.n648 source.n593 0.155672
R1649 source.n655 source.n593 0.155672
R1650 source.n656 source.n655 0.155672
R1651 source.n656 source.n589 0.155672
R1652 source.n663 source.n589 0.155672
R1653 source.n664 source.n663 0.155672
R1654 source.n664 source.n585 0.155672
R1655 source.n671 source.n585 0.155672
R1656 source.n672 source.n671 0.155672
R1657 source.n672 source.n581 0.155672
R1658 source.n680 source.n581 0.155672
R1659 source.n681 source.n680 0.155672
R1660 source.n681 source.n577 0.155672
R1661 source.n689 source.n577 0.155672
R1662 source.n690 source.n689 0.155672
R1663 source.n690 source.n573 0.155672
R1664 source.n697 source.n573 0.155672
R1665 source.n698 source.n697 0.155672
R1666 source.n698 source.n569 0.155672
R1667 source.n705 source.n569 0.155672
R1668 source.n137 source.n1 0.155672
R1669 source.n130 source.n1 0.155672
R1670 source.n130 source.n129 0.155672
R1671 source.n129 source.n5 0.155672
R1672 source.n122 source.n5 0.155672
R1673 source.n122 source.n121 0.155672
R1674 source.n121 source.n9 0.155672
R1675 source.n113 source.n9 0.155672
R1676 source.n113 source.n112 0.155672
R1677 source.n112 source.n13 0.155672
R1678 source.n105 source.n13 0.155672
R1679 source.n105 source.n104 0.155672
R1680 source.n104 source.n18 0.155672
R1681 source.n97 source.n18 0.155672
R1682 source.n97 source.n96 0.155672
R1683 source.n96 source.n22 0.155672
R1684 source.n89 source.n22 0.155672
R1685 source.n89 source.n88 0.155672
R1686 source.n88 source.n26 0.155672
R1687 source.n81 source.n26 0.155672
R1688 source.n81 source.n80 0.155672
R1689 source.n80 source.n30 0.155672
R1690 source.n73 source.n30 0.155672
R1691 source.n73 source.n72 0.155672
R1692 source.n72 source.n34 0.155672
R1693 source.n64 source.n34 0.155672
R1694 source.n64 source.n63 0.155672
R1695 source.n63 source.n39 0.155672
R1696 source.n56 source.n39 0.155672
R1697 source.n56 source.n55 0.155672
R1698 source.n55 source.n43 0.155672
R1699 source.n48 source.n43 0.155672
R1700 source.n281 source.n145 0.155672
R1701 source.n274 source.n145 0.155672
R1702 source.n274 source.n273 0.155672
R1703 source.n273 source.n149 0.155672
R1704 source.n266 source.n149 0.155672
R1705 source.n266 source.n265 0.155672
R1706 source.n265 source.n153 0.155672
R1707 source.n257 source.n153 0.155672
R1708 source.n257 source.n256 0.155672
R1709 source.n256 source.n157 0.155672
R1710 source.n249 source.n157 0.155672
R1711 source.n249 source.n248 0.155672
R1712 source.n248 source.n162 0.155672
R1713 source.n241 source.n162 0.155672
R1714 source.n241 source.n240 0.155672
R1715 source.n240 source.n166 0.155672
R1716 source.n233 source.n166 0.155672
R1717 source.n233 source.n232 0.155672
R1718 source.n232 source.n170 0.155672
R1719 source.n225 source.n170 0.155672
R1720 source.n225 source.n224 0.155672
R1721 source.n224 source.n174 0.155672
R1722 source.n217 source.n174 0.155672
R1723 source.n217 source.n216 0.155672
R1724 source.n216 source.n178 0.155672
R1725 source.n208 source.n178 0.155672
R1726 source.n208 source.n207 0.155672
R1727 source.n207 source.n183 0.155672
R1728 source.n200 source.n183 0.155672
R1729 source.n200 source.n199 0.155672
R1730 source.n199 source.n187 0.155672
R1731 source.n192 source.n187 0.155672
R1732 source.n421 source.n285 0.155672
R1733 source.n414 source.n285 0.155672
R1734 source.n414 source.n413 0.155672
R1735 source.n413 source.n289 0.155672
R1736 source.n406 source.n289 0.155672
R1737 source.n406 source.n405 0.155672
R1738 source.n405 source.n293 0.155672
R1739 source.n397 source.n293 0.155672
R1740 source.n397 source.n396 0.155672
R1741 source.n396 source.n297 0.155672
R1742 source.n389 source.n297 0.155672
R1743 source.n389 source.n388 0.155672
R1744 source.n388 source.n302 0.155672
R1745 source.n381 source.n302 0.155672
R1746 source.n381 source.n380 0.155672
R1747 source.n380 source.n306 0.155672
R1748 source.n373 source.n306 0.155672
R1749 source.n373 source.n372 0.155672
R1750 source.n372 source.n310 0.155672
R1751 source.n365 source.n310 0.155672
R1752 source.n365 source.n364 0.155672
R1753 source.n364 source.n314 0.155672
R1754 source.n357 source.n314 0.155672
R1755 source.n357 source.n356 0.155672
R1756 source.n356 source.n318 0.155672
R1757 source.n348 source.n318 0.155672
R1758 source.n348 source.n347 0.155672
R1759 source.n347 source.n323 0.155672
R1760 source.n340 source.n323 0.155672
R1761 source.n340 source.n339 0.155672
R1762 source.n339 source.n327 0.155672
R1763 source.n332 source.n327 0.155672
R1764 source.n565 source.n429 0.155672
R1765 source.n558 source.n429 0.155672
R1766 source.n558 source.n557 0.155672
R1767 source.n557 source.n433 0.155672
R1768 source.n550 source.n433 0.155672
R1769 source.n550 source.n549 0.155672
R1770 source.n549 source.n437 0.155672
R1771 source.n541 source.n437 0.155672
R1772 source.n541 source.n540 0.155672
R1773 source.n540 source.n441 0.155672
R1774 source.n533 source.n441 0.155672
R1775 source.n533 source.n532 0.155672
R1776 source.n532 source.n446 0.155672
R1777 source.n525 source.n446 0.155672
R1778 source.n525 source.n524 0.155672
R1779 source.n524 source.n450 0.155672
R1780 source.n517 source.n450 0.155672
R1781 source.n517 source.n516 0.155672
R1782 source.n516 source.n454 0.155672
R1783 source.n509 source.n454 0.155672
R1784 source.n509 source.n508 0.155672
R1785 source.n508 source.n458 0.155672
R1786 source.n501 source.n458 0.155672
R1787 source.n501 source.n500 0.155672
R1788 source.n500 source.n462 0.155672
R1789 source.n492 source.n462 0.155672
R1790 source.n492 source.n491 0.155672
R1791 source.n491 source.n467 0.155672
R1792 source.n484 source.n467 0.155672
R1793 source.n484 source.n483 0.155672
R1794 source.n483 source.n471 0.155672
R1795 source.n476 source.n471 0.155672
R1796 plus.n2 plus.t0 2160.24
R1797 plus.n13 plus.t5 2160.24
R1798 plus.n17 plus.t10 2160.24
R1799 plus.n28 plus.t8 2160.24
R1800 plus.n3 plus.t3 2112.77
R1801 plus.n4 plus.t7 2112.77
R1802 plus.n10 plus.t9 2112.77
R1803 plus.n12 plus.t2 2112.77
R1804 plus.n19 plus.t4 2112.77
R1805 plus.n18 plus.t11 2112.77
R1806 plus.n25 plus.t6 2112.77
R1807 plus.n27 plus.t1 2112.77
R1808 plus.n6 plus.n2 161.489
R1809 plus.n21 plus.n17 161.489
R1810 plus.n6 plus.n5 161.3
R1811 plus.n7 plus.n1 161.3
R1812 plus.n9 plus.n8 161.3
R1813 plus.n11 plus.n0 161.3
R1814 plus.n14 plus.n13 161.3
R1815 plus.n21 plus.n20 161.3
R1816 plus.n22 plus.n16 161.3
R1817 plus.n24 plus.n23 161.3
R1818 plus.n26 plus.n15 161.3
R1819 plus.n29 plus.n28 161.3
R1820 plus.n9 plus.n1 73.0308
R1821 plus.n24 plus.n16 73.0308
R1822 plus.n5 plus.n4 63.5369
R1823 plus.n11 plus.n10 63.5369
R1824 plus.n26 plus.n25 63.5369
R1825 plus.n20 plus.n18 63.5369
R1826 plus.n3 plus.n2 44.549
R1827 plus.n13 plus.n12 44.549
R1828 plus.n28 plus.n27 44.549
R1829 plus.n19 plus.n17 44.549
R1830 plus plus.n29 33.9914
R1831 plus.n5 plus.n3 28.4823
R1832 plus.n12 plus.n11 28.4823
R1833 plus.n27 plus.n26 28.4823
R1834 plus.n20 plus.n19 28.4823
R1835 plus plus.n14 17.08
R1836 plus.n4 plus.n1 9.49444
R1837 plus.n10 plus.n9 9.49444
R1838 plus.n25 plus.n24 9.49444
R1839 plus.n18 plus.n16 9.49444
R1840 plus.n7 plus.n6 0.189894
R1841 plus.n8 plus.n7 0.189894
R1842 plus.n8 plus.n0 0.189894
R1843 plus.n14 plus.n0 0.189894
R1844 plus.n29 plus.n15 0.189894
R1845 plus.n23 plus.n15 0.189894
R1846 plus.n23 plus.n22 0.189894
R1847 plus.n22 plus.n21 0.189894
R1848 drain_left.n6 drain_left.n4 59.2585
R1849 drain_left.n3 drain_left.n2 59.2032
R1850 drain_left.n3 drain_left.n0 59.2032
R1851 drain_left.n3 drain_left.n1 58.7154
R1852 drain_left.n6 drain_left.n5 58.7154
R1853 drain_left.n8 drain_left.n7 58.7153
R1854 drain_left drain_left.n3 39.9311
R1855 drain_left drain_left.n8 6.19632
R1856 drain_left.n1 drain_left.t5 0.7925
R1857 drain_left.n1 drain_left.t0 0.7925
R1858 drain_left.n2 drain_left.t7 0.7925
R1859 drain_left.n2 drain_left.t1 0.7925
R1860 drain_left.n0 drain_left.t3 0.7925
R1861 drain_left.n0 drain_left.t10 0.7925
R1862 drain_left.n7 drain_left.t9 0.7925
R1863 drain_left.n7 drain_left.t6 0.7925
R1864 drain_left.n5 drain_left.t4 0.7925
R1865 drain_left.n5 drain_left.t2 0.7925
R1866 drain_left.n4 drain_left.t11 0.7925
R1867 drain_left.n4 drain_left.t8 0.7925
R1868 drain_left.n8 drain_left.n6 0.543603
C0 plus drain_right 0.30725f
C1 minus plus 7.55094f
C2 plus drain_left 9.34205f
C3 source drain_right 46.5f
C4 minus source 8.26226f
C5 minus drain_right 9.18859f
C6 source drain_left 46.5003f
C7 drain_right drain_left 0.785787f
C8 minus drain_left 0.170859f
C9 plus source 8.276299f
C10 drain_right a_n1598_n5888# 8.90834f
C11 drain_left a_n1598_n5888# 9.1565f
C12 source a_n1598_n5888# 15.700303f
C13 minus a_n1598_n5888# 7.076188f
C14 plus a_n1598_n5888# 9.935321f
C15 drain_left.t3 a_n1598_n5888# 0.674884f
C16 drain_left.t10 a_n1598_n5888# 0.674884f
C17 drain_left.n0 a_n1598_n5888# 6.22322f
C18 drain_left.t5 a_n1598_n5888# 0.674884f
C19 drain_left.t0 a_n1598_n5888# 0.674884f
C20 drain_left.n1 a_n1598_n5888# 6.21978f
C21 drain_left.t7 a_n1598_n5888# 0.674884f
C22 drain_left.t1 a_n1598_n5888# 0.674884f
C23 drain_left.n2 a_n1598_n5888# 6.22322f
C24 drain_left.n3 a_n1598_n5888# 3.88665f
C25 drain_left.t11 a_n1598_n5888# 0.674884f
C26 drain_left.t8 a_n1598_n5888# 0.674884f
C27 drain_left.n4 a_n1598_n5888# 6.22365f
C28 drain_left.t4 a_n1598_n5888# 0.674884f
C29 drain_left.t2 a_n1598_n5888# 0.674884f
C30 drain_left.n5 a_n1598_n5888# 6.21978f
C31 drain_left.n6 a_n1598_n5888# 0.826543f
C32 drain_left.t9 a_n1598_n5888# 0.674884f
C33 drain_left.t6 a_n1598_n5888# 0.674884f
C34 drain_left.n7 a_n1598_n5888# 6.21977f
C35 drain_left.n8 a_n1598_n5888# 0.692687f
C36 plus.n0 a_n1598_n5888# 0.053245f
C37 plus.t2 a_n1598_n5888# 1.12361f
C38 plus.t9 a_n1598_n5888# 1.12361f
C39 plus.n1 a_n1598_n5888# 0.019797f
C40 plus.t0 a_n1598_n5888# 1.13268f
C41 plus.n2 a_n1598_n5888# 0.425896f
C42 plus.t3 a_n1598_n5888# 1.12361f
C43 plus.n3 a_n1598_n5888# 0.408857f
C44 plus.t7 a_n1598_n5888# 1.12361f
C45 plus.n4 a_n1598_n5888# 0.408857f
C46 plus.n5 a_n1598_n5888# 0.021931f
C47 plus.n6 a_n1598_n5888# 0.121183f
C48 plus.n7 a_n1598_n5888# 0.053245f
C49 plus.n8 a_n1598_n5888# 0.053245f
C50 plus.n9 a_n1598_n5888# 0.019797f
C51 plus.n10 a_n1598_n5888# 0.408857f
C52 plus.n11 a_n1598_n5888# 0.021931f
C53 plus.n12 a_n1598_n5888# 0.408857f
C54 plus.t5 a_n1598_n5888# 1.13268f
C55 plus.n13 a_n1598_n5888# 0.425816f
C56 plus.n14 a_n1598_n5888# 0.951878f
C57 plus.n15 a_n1598_n5888# 0.053245f
C58 plus.t8 a_n1598_n5888# 1.13268f
C59 plus.t1 a_n1598_n5888# 1.12361f
C60 plus.t6 a_n1598_n5888# 1.12361f
C61 plus.n16 a_n1598_n5888# 0.019797f
C62 plus.t10 a_n1598_n5888# 1.13268f
C63 plus.n17 a_n1598_n5888# 0.425896f
C64 plus.t11 a_n1598_n5888# 1.12361f
C65 plus.n18 a_n1598_n5888# 0.408857f
C66 plus.t4 a_n1598_n5888# 1.12361f
C67 plus.n19 a_n1598_n5888# 0.408857f
C68 plus.n20 a_n1598_n5888# 0.021931f
C69 plus.n21 a_n1598_n5888# 0.121183f
C70 plus.n22 a_n1598_n5888# 0.053245f
C71 plus.n23 a_n1598_n5888# 0.053245f
C72 plus.n24 a_n1598_n5888# 0.019797f
C73 plus.n25 a_n1598_n5888# 0.408857f
C74 plus.n26 a_n1598_n5888# 0.021931f
C75 plus.n27 a_n1598_n5888# 0.408857f
C76 plus.n28 a_n1598_n5888# 0.425816f
C77 plus.n29 a_n1598_n5888# 1.98897f
C78 source.n0 a_n1598_n5888# 0.035954f
C79 source.n1 a_n1598_n5888# 0.02608f
C80 source.n2 a_n1598_n5888# 0.014014f
C81 source.n3 a_n1598_n5888# 0.033125f
C82 source.n4 a_n1598_n5888# 0.014839f
C83 source.n5 a_n1598_n5888# 0.02608f
C84 source.n6 a_n1598_n5888# 0.014014f
C85 source.n7 a_n1598_n5888# 0.033125f
C86 source.n8 a_n1598_n5888# 0.014839f
C87 source.n9 a_n1598_n5888# 0.02608f
C88 source.n10 a_n1598_n5888# 0.014014f
C89 source.n11 a_n1598_n5888# 0.033125f
C90 source.n12 a_n1598_n5888# 0.014839f
C91 source.n13 a_n1598_n5888# 0.02608f
C92 source.n14 a_n1598_n5888# 0.014014f
C93 source.n15 a_n1598_n5888# 0.033125f
C94 source.n16 a_n1598_n5888# 0.033125f
C95 source.n17 a_n1598_n5888# 0.014839f
C96 source.n18 a_n1598_n5888# 0.02608f
C97 source.n19 a_n1598_n5888# 0.014014f
C98 source.n20 a_n1598_n5888# 0.033125f
C99 source.n21 a_n1598_n5888# 0.014839f
C100 source.n22 a_n1598_n5888# 0.02608f
C101 source.n23 a_n1598_n5888# 0.014014f
C102 source.n24 a_n1598_n5888# 0.033125f
C103 source.n25 a_n1598_n5888# 0.014839f
C104 source.n26 a_n1598_n5888# 0.02608f
C105 source.n27 a_n1598_n5888# 0.014014f
C106 source.n28 a_n1598_n5888# 0.033125f
C107 source.n29 a_n1598_n5888# 0.014839f
C108 source.n30 a_n1598_n5888# 0.02608f
C109 source.n31 a_n1598_n5888# 0.014014f
C110 source.n32 a_n1598_n5888# 0.033125f
C111 source.n33 a_n1598_n5888# 0.014839f
C112 source.n34 a_n1598_n5888# 0.02608f
C113 source.n35 a_n1598_n5888# 0.014427f
C114 source.n36 a_n1598_n5888# 0.033125f
C115 source.n37 a_n1598_n5888# 0.014014f
C116 source.n38 a_n1598_n5888# 0.014839f
C117 source.n39 a_n1598_n5888# 0.02608f
C118 source.n40 a_n1598_n5888# 0.014014f
C119 source.n41 a_n1598_n5888# 0.033125f
C120 source.n42 a_n1598_n5888# 0.014839f
C121 source.n43 a_n1598_n5888# 0.02608f
C122 source.n44 a_n1598_n5888# 0.014014f
C123 source.n45 a_n1598_n5888# 0.024844f
C124 source.n46 a_n1598_n5888# 0.023417f
C125 source.t2 a_n1598_n5888# 0.057772f
C126 source.n47 a_n1598_n5888# 0.318202f
C127 source.n48 a_n1598_n5888# 2.82373f
C128 source.n49 a_n1598_n5888# 0.014014f
C129 source.n50 a_n1598_n5888# 0.014839f
C130 source.n51 a_n1598_n5888# 0.033125f
C131 source.n52 a_n1598_n5888# 0.033125f
C132 source.n53 a_n1598_n5888# 0.014839f
C133 source.n54 a_n1598_n5888# 0.014014f
C134 source.n55 a_n1598_n5888# 0.02608f
C135 source.n56 a_n1598_n5888# 0.02608f
C136 source.n57 a_n1598_n5888# 0.014014f
C137 source.n58 a_n1598_n5888# 0.014839f
C138 source.n59 a_n1598_n5888# 0.033125f
C139 source.n60 a_n1598_n5888# 0.033125f
C140 source.n61 a_n1598_n5888# 0.014839f
C141 source.n62 a_n1598_n5888# 0.014014f
C142 source.n63 a_n1598_n5888# 0.02608f
C143 source.n64 a_n1598_n5888# 0.02608f
C144 source.n65 a_n1598_n5888# 0.014014f
C145 source.n66 a_n1598_n5888# 0.014839f
C146 source.n67 a_n1598_n5888# 0.033125f
C147 source.n68 a_n1598_n5888# 0.033125f
C148 source.n69 a_n1598_n5888# 0.033125f
C149 source.n70 a_n1598_n5888# 0.014427f
C150 source.n71 a_n1598_n5888# 0.014014f
C151 source.n72 a_n1598_n5888# 0.02608f
C152 source.n73 a_n1598_n5888# 0.02608f
C153 source.n74 a_n1598_n5888# 0.014014f
C154 source.n75 a_n1598_n5888# 0.014839f
C155 source.n76 a_n1598_n5888# 0.033125f
C156 source.n77 a_n1598_n5888# 0.033125f
C157 source.n78 a_n1598_n5888# 0.014839f
C158 source.n79 a_n1598_n5888# 0.014014f
C159 source.n80 a_n1598_n5888# 0.02608f
C160 source.n81 a_n1598_n5888# 0.02608f
C161 source.n82 a_n1598_n5888# 0.014014f
C162 source.n83 a_n1598_n5888# 0.014839f
C163 source.n84 a_n1598_n5888# 0.033125f
C164 source.n85 a_n1598_n5888# 0.033125f
C165 source.n86 a_n1598_n5888# 0.014839f
C166 source.n87 a_n1598_n5888# 0.014014f
C167 source.n88 a_n1598_n5888# 0.02608f
C168 source.n89 a_n1598_n5888# 0.02608f
C169 source.n90 a_n1598_n5888# 0.014014f
C170 source.n91 a_n1598_n5888# 0.014839f
C171 source.n92 a_n1598_n5888# 0.033125f
C172 source.n93 a_n1598_n5888# 0.033125f
C173 source.n94 a_n1598_n5888# 0.014839f
C174 source.n95 a_n1598_n5888# 0.014014f
C175 source.n96 a_n1598_n5888# 0.02608f
C176 source.n97 a_n1598_n5888# 0.02608f
C177 source.n98 a_n1598_n5888# 0.014014f
C178 source.n99 a_n1598_n5888# 0.014839f
C179 source.n100 a_n1598_n5888# 0.033125f
C180 source.n101 a_n1598_n5888# 0.033125f
C181 source.n102 a_n1598_n5888# 0.014839f
C182 source.n103 a_n1598_n5888# 0.014014f
C183 source.n104 a_n1598_n5888# 0.02608f
C184 source.n105 a_n1598_n5888# 0.02608f
C185 source.n106 a_n1598_n5888# 0.014014f
C186 source.n107 a_n1598_n5888# 0.014839f
C187 source.n108 a_n1598_n5888# 0.033125f
C188 source.n109 a_n1598_n5888# 0.033125f
C189 source.n110 a_n1598_n5888# 0.014839f
C190 source.n111 a_n1598_n5888# 0.014014f
C191 source.n112 a_n1598_n5888# 0.02608f
C192 source.n113 a_n1598_n5888# 0.02608f
C193 source.n114 a_n1598_n5888# 0.014014f
C194 source.n115 a_n1598_n5888# 0.014427f
C195 source.n116 a_n1598_n5888# 0.014427f
C196 source.n117 a_n1598_n5888# 0.033125f
C197 source.n118 a_n1598_n5888# 0.033125f
C198 source.n119 a_n1598_n5888# 0.014839f
C199 source.n120 a_n1598_n5888# 0.014014f
C200 source.n121 a_n1598_n5888# 0.02608f
C201 source.n122 a_n1598_n5888# 0.02608f
C202 source.n123 a_n1598_n5888# 0.014014f
C203 source.n124 a_n1598_n5888# 0.014839f
C204 source.n125 a_n1598_n5888# 0.033125f
C205 source.n126 a_n1598_n5888# 0.033125f
C206 source.n127 a_n1598_n5888# 0.014839f
C207 source.n128 a_n1598_n5888# 0.014014f
C208 source.n129 a_n1598_n5888# 0.02608f
C209 source.n130 a_n1598_n5888# 0.02608f
C210 source.n131 a_n1598_n5888# 0.014014f
C211 source.n132 a_n1598_n5888# 0.014839f
C212 source.n133 a_n1598_n5888# 0.033125f
C213 source.n134 a_n1598_n5888# 0.070465f
C214 source.n135 a_n1598_n5888# 0.014839f
C215 source.n136 a_n1598_n5888# 0.014014f
C216 source.n137 a_n1598_n5888# 0.057433f
C217 source.n138 a_n1598_n5888# 0.039211f
C218 source.n139 a_n1598_n5888# 2.04971f
C219 source.t4 a_n1598_n5888# 0.515236f
C220 source.t8 a_n1598_n5888# 0.515236f
C221 source.n140 a_n1598_n5888# 4.66296f
C222 source.n141 a_n1598_n5888# 0.361785f
C223 source.t11 a_n1598_n5888# 0.515236f
C224 source.t7 a_n1598_n5888# 0.515236f
C225 source.n142 a_n1598_n5888# 4.66296f
C226 source.n143 a_n1598_n5888# 0.361785f
C227 source.n144 a_n1598_n5888# 0.035954f
C228 source.n145 a_n1598_n5888# 0.02608f
C229 source.n146 a_n1598_n5888# 0.014014f
C230 source.n147 a_n1598_n5888# 0.033125f
C231 source.n148 a_n1598_n5888# 0.014839f
C232 source.n149 a_n1598_n5888# 0.02608f
C233 source.n150 a_n1598_n5888# 0.014014f
C234 source.n151 a_n1598_n5888# 0.033125f
C235 source.n152 a_n1598_n5888# 0.014839f
C236 source.n153 a_n1598_n5888# 0.02608f
C237 source.n154 a_n1598_n5888# 0.014014f
C238 source.n155 a_n1598_n5888# 0.033125f
C239 source.n156 a_n1598_n5888# 0.014839f
C240 source.n157 a_n1598_n5888# 0.02608f
C241 source.n158 a_n1598_n5888# 0.014014f
C242 source.n159 a_n1598_n5888# 0.033125f
C243 source.n160 a_n1598_n5888# 0.033125f
C244 source.n161 a_n1598_n5888# 0.014839f
C245 source.n162 a_n1598_n5888# 0.02608f
C246 source.n163 a_n1598_n5888# 0.014014f
C247 source.n164 a_n1598_n5888# 0.033125f
C248 source.n165 a_n1598_n5888# 0.014839f
C249 source.n166 a_n1598_n5888# 0.02608f
C250 source.n167 a_n1598_n5888# 0.014014f
C251 source.n168 a_n1598_n5888# 0.033125f
C252 source.n169 a_n1598_n5888# 0.014839f
C253 source.n170 a_n1598_n5888# 0.02608f
C254 source.n171 a_n1598_n5888# 0.014014f
C255 source.n172 a_n1598_n5888# 0.033125f
C256 source.n173 a_n1598_n5888# 0.014839f
C257 source.n174 a_n1598_n5888# 0.02608f
C258 source.n175 a_n1598_n5888# 0.014014f
C259 source.n176 a_n1598_n5888# 0.033125f
C260 source.n177 a_n1598_n5888# 0.014839f
C261 source.n178 a_n1598_n5888# 0.02608f
C262 source.n179 a_n1598_n5888# 0.014427f
C263 source.n180 a_n1598_n5888# 0.033125f
C264 source.n181 a_n1598_n5888# 0.014014f
C265 source.n182 a_n1598_n5888# 0.014839f
C266 source.n183 a_n1598_n5888# 0.02608f
C267 source.n184 a_n1598_n5888# 0.014014f
C268 source.n185 a_n1598_n5888# 0.033125f
C269 source.n186 a_n1598_n5888# 0.014839f
C270 source.n187 a_n1598_n5888# 0.02608f
C271 source.n188 a_n1598_n5888# 0.014014f
C272 source.n189 a_n1598_n5888# 0.024844f
C273 source.n190 a_n1598_n5888# 0.023417f
C274 source.t9 a_n1598_n5888# 0.057772f
C275 source.n191 a_n1598_n5888# 0.318202f
C276 source.n192 a_n1598_n5888# 2.82373f
C277 source.n193 a_n1598_n5888# 0.014014f
C278 source.n194 a_n1598_n5888# 0.014839f
C279 source.n195 a_n1598_n5888# 0.033125f
C280 source.n196 a_n1598_n5888# 0.033125f
C281 source.n197 a_n1598_n5888# 0.014839f
C282 source.n198 a_n1598_n5888# 0.014014f
C283 source.n199 a_n1598_n5888# 0.02608f
C284 source.n200 a_n1598_n5888# 0.02608f
C285 source.n201 a_n1598_n5888# 0.014014f
C286 source.n202 a_n1598_n5888# 0.014839f
C287 source.n203 a_n1598_n5888# 0.033125f
C288 source.n204 a_n1598_n5888# 0.033125f
C289 source.n205 a_n1598_n5888# 0.014839f
C290 source.n206 a_n1598_n5888# 0.014014f
C291 source.n207 a_n1598_n5888# 0.02608f
C292 source.n208 a_n1598_n5888# 0.02608f
C293 source.n209 a_n1598_n5888# 0.014014f
C294 source.n210 a_n1598_n5888# 0.014839f
C295 source.n211 a_n1598_n5888# 0.033125f
C296 source.n212 a_n1598_n5888# 0.033125f
C297 source.n213 a_n1598_n5888# 0.033125f
C298 source.n214 a_n1598_n5888# 0.014427f
C299 source.n215 a_n1598_n5888# 0.014014f
C300 source.n216 a_n1598_n5888# 0.02608f
C301 source.n217 a_n1598_n5888# 0.02608f
C302 source.n218 a_n1598_n5888# 0.014014f
C303 source.n219 a_n1598_n5888# 0.014839f
C304 source.n220 a_n1598_n5888# 0.033125f
C305 source.n221 a_n1598_n5888# 0.033125f
C306 source.n222 a_n1598_n5888# 0.014839f
C307 source.n223 a_n1598_n5888# 0.014014f
C308 source.n224 a_n1598_n5888# 0.02608f
C309 source.n225 a_n1598_n5888# 0.02608f
C310 source.n226 a_n1598_n5888# 0.014014f
C311 source.n227 a_n1598_n5888# 0.014839f
C312 source.n228 a_n1598_n5888# 0.033125f
C313 source.n229 a_n1598_n5888# 0.033125f
C314 source.n230 a_n1598_n5888# 0.014839f
C315 source.n231 a_n1598_n5888# 0.014014f
C316 source.n232 a_n1598_n5888# 0.02608f
C317 source.n233 a_n1598_n5888# 0.02608f
C318 source.n234 a_n1598_n5888# 0.014014f
C319 source.n235 a_n1598_n5888# 0.014839f
C320 source.n236 a_n1598_n5888# 0.033125f
C321 source.n237 a_n1598_n5888# 0.033125f
C322 source.n238 a_n1598_n5888# 0.014839f
C323 source.n239 a_n1598_n5888# 0.014014f
C324 source.n240 a_n1598_n5888# 0.02608f
C325 source.n241 a_n1598_n5888# 0.02608f
C326 source.n242 a_n1598_n5888# 0.014014f
C327 source.n243 a_n1598_n5888# 0.014839f
C328 source.n244 a_n1598_n5888# 0.033125f
C329 source.n245 a_n1598_n5888# 0.033125f
C330 source.n246 a_n1598_n5888# 0.014839f
C331 source.n247 a_n1598_n5888# 0.014014f
C332 source.n248 a_n1598_n5888# 0.02608f
C333 source.n249 a_n1598_n5888# 0.02608f
C334 source.n250 a_n1598_n5888# 0.014014f
C335 source.n251 a_n1598_n5888# 0.014839f
C336 source.n252 a_n1598_n5888# 0.033125f
C337 source.n253 a_n1598_n5888# 0.033125f
C338 source.n254 a_n1598_n5888# 0.014839f
C339 source.n255 a_n1598_n5888# 0.014014f
C340 source.n256 a_n1598_n5888# 0.02608f
C341 source.n257 a_n1598_n5888# 0.02608f
C342 source.n258 a_n1598_n5888# 0.014014f
C343 source.n259 a_n1598_n5888# 0.014427f
C344 source.n260 a_n1598_n5888# 0.014427f
C345 source.n261 a_n1598_n5888# 0.033125f
C346 source.n262 a_n1598_n5888# 0.033125f
C347 source.n263 a_n1598_n5888# 0.014839f
C348 source.n264 a_n1598_n5888# 0.014014f
C349 source.n265 a_n1598_n5888# 0.02608f
C350 source.n266 a_n1598_n5888# 0.02608f
C351 source.n267 a_n1598_n5888# 0.014014f
C352 source.n268 a_n1598_n5888# 0.014839f
C353 source.n269 a_n1598_n5888# 0.033125f
C354 source.n270 a_n1598_n5888# 0.033125f
C355 source.n271 a_n1598_n5888# 0.014839f
C356 source.n272 a_n1598_n5888# 0.014014f
C357 source.n273 a_n1598_n5888# 0.02608f
C358 source.n274 a_n1598_n5888# 0.02608f
C359 source.n275 a_n1598_n5888# 0.014014f
C360 source.n276 a_n1598_n5888# 0.014839f
C361 source.n277 a_n1598_n5888# 0.033125f
C362 source.n278 a_n1598_n5888# 0.070465f
C363 source.n279 a_n1598_n5888# 0.014839f
C364 source.n280 a_n1598_n5888# 0.014014f
C365 source.n281 a_n1598_n5888# 0.057433f
C366 source.n282 a_n1598_n5888# 0.039211f
C367 source.n283 a_n1598_n5888# 0.105791f
C368 source.n284 a_n1598_n5888# 0.035954f
C369 source.n285 a_n1598_n5888# 0.02608f
C370 source.n286 a_n1598_n5888# 0.014014f
C371 source.n287 a_n1598_n5888# 0.033125f
C372 source.n288 a_n1598_n5888# 0.014839f
C373 source.n289 a_n1598_n5888# 0.02608f
C374 source.n290 a_n1598_n5888# 0.014014f
C375 source.n291 a_n1598_n5888# 0.033125f
C376 source.n292 a_n1598_n5888# 0.014839f
C377 source.n293 a_n1598_n5888# 0.02608f
C378 source.n294 a_n1598_n5888# 0.014014f
C379 source.n295 a_n1598_n5888# 0.033125f
C380 source.n296 a_n1598_n5888# 0.014839f
C381 source.n297 a_n1598_n5888# 0.02608f
C382 source.n298 a_n1598_n5888# 0.014014f
C383 source.n299 a_n1598_n5888# 0.033125f
C384 source.n300 a_n1598_n5888# 0.033125f
C385 source.n301 a_n1598_n5888# 0.014839f
C386 source.n302 a_n1598_n5888# 0.02608f
C387 source.n303 a_n1598_n5888# 0.014014f
C388 source.n304 a_n1598_n5888# 0.033125f
C389 source.n305 a_n1598_n5888# 0.014839f
C390 source.n306 a_n1598_n5888# 0.02608f
C391 source.n307 a_n1598_n5888# 0.014014f
C392 source.n308 a_n1598_n5888# 0.033125f
C393 source.n309 a_n1598_n5888# 0.014839f
C394 source.n310 a_n1598_n5888# 0.02608f
C395 source.n311 a_n1598_n5888# 0.014014f
C396 source.n312 a_n1598_n5888# 0.033125f
C397 source.n313 a_n1598_n5888# 0.014839f
C398 source.n314 a_n1598_n5888# 0.02608f
C399 source.n315 a_n1598_n5888# 0.014014f
C400 source.n316 a_n1598_n5888# 0.033125f
C401 source.n317 a_n1598_n5888# 0.014839f
C402 source.n318 a_n1598_n5888# 0.02608f
C403 source.n319 a_n1598_n5888# 0.014427f
C404 source.n320 a_n1598_n5888# 0.033125f
C405 source.n321 a_n1598_n5888# 0.014014f
C406 source.n322 a_n1598_n5888# 0.014839f
C407 source.n323 a_n1598_n5888# 0.02608f
C408 source.n324 a_n1598_n5888# 0.014014f
C409 source.n325 a_n1598_n5888# 0.033125f
C410 source.n326 a_n1598_n5888# 0.014839f
C411 source.n327 a_n1598_n5888# 0.02608f
C412 source.n328 a_n1598_n5888# 0.014014f
C413 source.n329 a_n1598_n5888# 0.024844f
C414 source.n330 a_n1598_n5888# 0.023417f
C415 source.t17 a_n1598_n5888# 0.057772f
C416 source.n331 a_n1598_n5888# 0.318202f
C417 source.n332 a_n1598_n5888# 2.82373f
C418 source.n333 a_n1598_n5888# 0.014014f
C419 source.n334 a_n1598_n5888# 0.014839f
C420 source.n335 a_n1598_n5888# 0.033125f
C421 source.n336 a_n1598_n5888# 0.033125f
C422 source.n337 a_n1598_n5888# 0.014839f
C423 source.n338 a_n1598_n5888# 0.014014f
C424 source.n339 a_n1598_n5888# 0.02608f
C425 source.n340 a_n1598_n5888# 0.02608f
C426 source.n341 a_n1598_n5888# 0.014014f
C427 source.n342 a_n1598_n5888# 0.014839f
C428 source.n343 a_n1598_n5888# 0.033125f
C429 source.n344 a_n1598_n5888# 0.033125f
C430 source.n345 a_n1598_n5888# 0.014839f
C431 source.n346 a_n1598_n5888# 0.014014f
C432 source.n347 a_n1598_n5888# 0.02608f
C433 source.n348 a_n1598_n5888# 0.02608f
C434 source.n349 a_n1598_n5888# 0.014014f
C435 source.n350 a_n1598_n5888# 0.014839f
C436 source.n351 a_n1598_n5888# 0.033125f
C437 source.n352 a_n1598_n5888# 0.033125f
C438 source.n353 a_n1598_n5888# 0.033125f
C439 source.n354 a_n1598_n5888# 0.014427f
C440 source.n355 a_n1598_n5888# 0.014014f
C441 source.n356 a_n1598_n5888# 0.02608f
C442 source.n357 a_n1598_n5888# 0.02608f
C443 source.n358 a_n1598_n5888# 0.014014f
C444 source.n359 a_n1598_n5888# 0.014839f
C445 source.n360 a_n1598_n5888# 0.033125f
C446 source.n361 a_n1598_n5888# 0.033125f
C447 source.n362 a_n1598_n5888# 0.014839f
C448 source.n363 a_n1598_n5888# 0.014014f
C449 source.n364 a_n1598_n5888# 0.02608f
C450 source.n365 a_n1598_n5888# 0.02608f
C451 source.n366 a_n1598_n5888# 0.014014f
C452 source.n367 a_n1598_n5888# 0.014839f
C453 source.n368 a_n1598_n5888# 0.033125f
C454 source.n369 a_n1598_n5888# 0.033125f
C455 source.n370 a_n1598_n5888# 0.014839f
C456 source.n371 a_n1598_n5888# 0.014014f
C457 source.n372 a_n1598_n5888# 0.02608f
C458 source.n373 a_n1598_n5888# 0.02608f
C459 source.n374 a_n1598_n5888# 0.014014f
C460 source.n375 a_n1598_n5888# 0.014839f
C461 source.n376 a_n1598_n5888# 0.033125f
C462 source.n377 a_n1598_n5888# 0.033125f
C463 source.n378 a_n1598_n5888# 0.014839f
C464 source.n379 a_n1598_n5888# 0.014014f
C465 source.n380 a_n1598_n5888# 0.02608f
C466 source.n381 a_n1598_n5888# 0.02608f
C467 source.n382 a_n1598_n5888# 0.014014f
C468 source.n383 a_n1598_n5888# 0.014839f
C469 source.n384 a_n1598_n5888# 0.033125f
C470 source.n385 a_n1598_n5888# 0.033125f
C471 source.n386 a_n1598_n5888# 0.014839f
C472 source.n387 a_n1598_n5888# 0.014014f
C473 source.n388 a_n1598_n5888# 0.02608f
C474 source.n389 a_n1598_n5888# 0.02608f
C475 source.n390 a_n1598_n5888# 0.014014f
C476 source.n391 a_n1598_n5888# 0.014839f
C477 source.n392 a_n1598_n5888# 0.033125f
C478 source.n393 a_n1598_n5888# 0.033125f
C479 source.n394 a_n1598_n5888# 0.014839f
C480 source.n395 a_n1598_n5888# 0.014014f
C481 source.n396 a_n1598_n5888# 0.02608f
C482 source.n397 a_n1598_n5888# 0.02608f
C483 source.n398 a_n1598_n5888# 0.014014f
C484 source.n399 a_n1598_n5888# 0.014427f
C485 source.n400 a_n1598_n5888# 0.014427f
C486 source.n401 a_n1598_n5888# 0.033125f
C487 source.n402 a_n1598_n5888# 0.033125f
C488 source.n403 a_n1598_n5888# 0.014839f
C489 source.n404 a_n1598_n5888# 0.014014f
C490 source.n405 a_n1598_n5888# 0.02608f
C491 source.n406 a_n1598_n5888# 0.02608f
C492 source.n407 a_n1598_n5888# 0.014014f
C493 source.n408 a_n1598_n5888# 0.014839f
C494 source.n409 a_n1598_n5888# 0.033125f
C495 source.n410 a_n1598_n5888# 0.033125f
C496 source.n411 a_n1598_n5888# 0.014839f
C497 source.n412 a_n1598_n5888# 0.014014f
C498 source.n413 a_n1598_n5888# 0.02608f
C499 source.n414 a_n1598_n5888# 0.02608f
C500 source.n415 a_n1598_n5888# 0.014014f
C501 source.n416 a_n1598_n5888# 0.014839f
C502 source.n417 a_n1598_n5888# 0.033125f
C503 source.n418 a_n1598_n5888# 0.070465f
C504 source.n419 a_n1598_n5888# 0.014839f
C505 source.n420 a_n1598_n5888# 0.014014f
C506 source.n421 a_n1598_n5888# 0.057433f
C507 source.n422 a_n1598_n5888# 0.039211f
C508 source.n423 a_n1598_n5888# 0.105791f
C509 source.t22 a_n1598_n5888# 0.515236f
C510 source.t13 a_n1598_n5888# 0.515236f
C511 source.n424 a_n1598_n5888# 4.66296f
C512 source.n425 a_n1598_n5888# 0.361785f
C513 source.t14 a_n1598_n5888# 0.515236f
C514 source.t18 a_n1598_n5888# 0.515236f
C515 source.n426 a_n1598_n5888# 4.66296f
C516 source.n427 a_n1598_n5888# 0.361785f
C517 source.n428 a_n1598_n5888# 0.035954f
C518 source.n429 a_n1598_n5888# 0.02608f
C519 source.n430 a_n1598_n5888# 0.014014f
C520 source.n431 a_n1598_n5888# 0.033125f
C521 source.n432 a_n1598_n5888# 0.014839f
C522 source.n433 a_n1598_n5888# 0.02608f
C523 source.n434 a_n1598_n5888# 0.014014f
C524 source.n435 a_n1598_n5888# 0.033125f
C525 source.n436 a_n1598_n5888# 0.014839f
C526 source.n437 a_n1598_n5888# 0.02608f
C527 source.n438 a_n1598_n5888# 0.014014f
C528 source.n439 a_n1598_n5888# 0.033125f
C529 source.n440 a_n1598_n5888# 0.014839f
C530 source.n441 a_n1598_n5888# 0.02608f
C531 source.n442 a_n1598_n5888# 0.014014f
C532 source.n443 a_n1598_n5888# 0.033125f
C533 source.n444 a_n1598_n5888# 0.033125f
C534 source.n445 a_n1598_n5888# 0.014839f
C535 source.n446 a_n1598_n5888# 0.02608f
C536 source.n447 a_n1598_n5888# 0.014014f
C537 source.n448 a_n1598_n5888# 0.033125f
C538 source.n449 a_n1598_n5888# 0.014839f
C539 source.n450 a_n1598_n5888# 0.02608f
C540 source.n451 a_n1598_n5888# 0.014014f
C541 source.n452 a_n1598_n5888# 0.033125f
C542 source.n453 a_n1598_n5888# 0.014839f
C543 source.n454 a_n1598_n5888# 0.02608f
C544 source.n455 a_n1598_n5888# 0.014014f
C545 source.n456 a_n1598_n5888# 0.033125f
C546 source.n457 a_n1598_n5888# 0.014839f
C547 source.n458 a_n1598_n5888# 0.02608f
C548 source.n459 a_n1598_n5888# 0.014014f
C549 source.n460 a_n1598_n5888# 0.033125f
C550 source.n461 a_n1598_n5888# 0.014839f
C551 source.n462 a_n1598_n5888# 0.02608f
C552 source.n463 a_n1598_n5888# 0.014427f
C553 source.n464 a_n1598_n5888# 0.033125f
C554 source.n465 a_n1598_n5888# 0.014014f
C555 source.n466 a_n1598_n5888# 0.014839f
C556 source.n467 a_n1598_n5888# 0.02608f
C557 source.n468 a_n1598_n5888# 0.014014f
C558 source.n469 a_n1598_n5888# 0.033125f
C559 source.n470 a_n1598_n5888# 0.014839f
C560 source.n471 a_n1598_n5888# 0.02608f
C561 source.n472 a_n1598_n5888# 0.014014f
C562 source.n473 a_n1598_n5888# 0.024844f
C563 source.n474 a_n1598_n5888# 0.023417f
C564 source.t23 a_n1598_n5888# 0.057772f
C565 source.n475 a_n1598_n5888# 0.318202f
C566 source.n476 a_n1598_n5888# 2.82373f
C567 source.n477 a_n1598_n5888# 0.014014f
C568 source.n478 a_n1598_n5888# 0.014839f
C569 source.n479 a_n1598_n5888# 0.033125f
C570 source.n480 a_n1598_n5888# 0.033125f
C571 source.n481 a_n1598_n5888# 0.014839f
C572 source.n482 a_n1598_n5888# 0.014014f
C573 source.n483 a_n1598_n5888# 0.02608f
C574 source.n484 a_n1598_n5888# 0.02608f
C575 source.n485 a_n1598_n5888# 0.014014f
C576 source.n486 a_n1598_n5888# 0.014839f
C577 source.n487 a_n1598_n5888# 0.033125f
C578 source.n488 a_n1598_n5888# 0.033125f
C579 source.n489 a_n1598_n5888# 0.014839f
C580 source.n490 a_n1598_n5888# 0.014014f
C581 source.n491 a_n1598_n5888# 0.02608f
C582 source.n492 a_n1598_n5888# 0.02608f
C583 source.n493 a_n1598_n5888# 0.014014f
C584 source.n494 a_n1598_n5888# 0.014839f
C585 source.n495 a_n1598_n5888# 0.033125f
C586 source.n496 a_n1598_n5888# 0.033125f
C587 source.n497 a_n1598_n5888# 0.033125f
C588 source.n498 a_n1598_n5888# 0.014427f
C589 source.n499 a_n1598_n5888# 0.014014f
C590 source.n500 a_n1598_n5888# 0.02608f
C591 source.n501 a_n1598_n5888# 0.02608f
C592 source.n502 a_n1598_n5888# 0.014014f
C593 source.n503 a_n1598_n5888# 0.014839f
C594 source.n504 a_n1598_n5888# 0.033125f
C595 source.n505 a_n1598_n5888# 0.033125f
C596 source.n506 a_n1598_n5888# 0.014839f
C597 source.n507 a_n1598_n5888# 0.014014f
C598 source.n508 a_n1598_n5888# 0.02608f
C599 source.n509 a_n1598_n5888# 0.02608f
C600 source.n510 a_n1598_n5888# 0.014014f
C601 source.n511 a_n1598_n5888# 0.014839f
C602 source.n512 a_n1598_n5888# 0.033125f
C603 source.n513 a_n1598_n5888# 0.033125f
C604 source.n514 a_n1598_n5888# 0.014839f
C605 source.n515 a_n1598_n5888# 0.014014f
C606 source.n516 a_n1598_n5888# 0.02608f
C607 source.n517 a_n1598_n5888# 0.02608f
C608 source.n518 a_n1598_n5888# 0.014014f
C609 source.n519 a_n1598_n5888# 0.014839f
C610 source.n520 a_n1598_n5888# 0.033125f
C611 source.n521 a_n1598_n5888# 0.033125f
C612 source.n522 a_n1598_n5888# 0.014839f
C613 source.n523 a_n1598_n5888# 0.014014f
C614 source.n524 a_n1598_n5888# 0.02608f
C615 source.n525 a_n1598_n5888# 0.02608f
C616 source.n526 a_n1598_n5888# 0.014014f
C617 source.n527 a_n1598_n5888# 0.014839f
C618 source.n528 a_n1598_n5888# 0.033125f
C619 source.n529 a_n1598_n5888# 0.033125f
C620 source.n530 a_n1598_n5888# 0.014839f
C621 source.n531 a_n1598_n5888# 0.014014f
C622 source.n532 a_n1598_n5888# 0.02608f
C623 source.n533 a_n1598_n5888# 0.02608f
C624 source.n534 a_n1598_n5888# 0.014014f
C625 source.n535 a_n1598_n5888# 0.014839f
C626 source.n536 a_n1598_n5888# 0.033125f
C627 source.n537 a_n1598_n5888# 0.033125f
C628 source.n538 a_n1598_n5888# 0.014839f
C629 source.n539 a_n1598_n5888# 0.014014f
C630 source.n540 a_n1598_n5888# 0.02608f
C631 source.n541 a_n1598_n5888# 0.02608f
C632 source.n542 a_n1598_n5888# 0.014014f
C633 source.n543 a_n1598_n5888# 0.014427f
C634 source.n544 a_n1598_n5888# 0.014427f
C635 source.n545 a_n1598_n5888# 0.033125f
C636 source.n546 a_n1598_n5888# 0.033125f
C637 source.n547 a_n1598_n5888# 0.014839f
C638 source.n548 a_n1598_n5888# 0.014014f
C639 source.n549 a_n1598_n5888# 0.02608f
C640 source.n550 a_n1598_n5888# 0.02608f
C641 source.n551 a_n1598_n5888# 0.014014f
C642 source.n552 a_n1598_n5888# 0.014839f
C643 source.n553 a_n1598_n5888# 0.033125f
C644 source.n554 a_n1598_n5888# 0.033125f
C645 source.n555 a_n1598_n5888# 0.014839f
C646 source.n556 a_n1598_n5888# 0.014014f
C647 source.n557 a_n1598_n5888# 0.02608f
C648 source.n558 a_n1598_n5888# 0.02608f
C649 source.n559 a_n1598_n5888# 0.014014f
C650 source.n560 a_n1598_n5888# 0.014839f
C651 source.n561 a_n1598_n5888# 0.033125f
C652 source.n562 a_n1598_n5888# 0.070465f
C653 source.n563 a_n1598_n5888# 0.014839f
C654 source.n564 a_n1598_n5888# 0.014014f
C655 source.n565 a_n1598_n5888# 0.057433f
C656 source.n566 a_n1598_n5888# 0.039211f
C657 source.n567 a_n1598_n5888# 2.53218f
C658 source.n568 a_n1598_n5888# 0.035954f
C659 source.n569 a_n1598_n5888# 0.02608f
C660 source.n570 a_n1598_n5888# 0.014014f
C661 source.n571 a_n1598_n5888# 0.033125f
C662 source.n572 a_n1598_n5888# 0.014839f
C663 source.n573 a_n1598_n5888# 0.02608f
C664 source.n574 a_n1598_n5888# 0.014014f
C665 source.n575 a_n1598_n5888# 0.033125f
C666 source.n576 a_n1598_n5888# 0.014839f
C667 source.n577 a_n1598_n5888# 0.02608f
C668 source.n578 a_n1598_n5888# 0.014014f
C669 source.n579 a_n1598_n5888# 0.033125f
C670 source.n580 a_n1598_n5888# 0.014839f
C671 source.n581 a_n1598_n5888# 0.02608f
C672 source.n582 a_n1598_n5888# 0.014014f
C673 source.n583 a_n1598_n5888# 0.033125f
C674 source.n584 a_n1598_n5888# 0.014839f
C675 source.n585 a_n1598_n5888# 0.02608f
C676 source.n586 a_n1598_n5888# 0.014014f
C677 source.n587 a_n1598_n5888# 0.033125f
C678 source.n588 a_n1598_n5888# 0.014839f
C679 source.n589 a_n1598_n5888# 0.02608f
C680 source.n590 a_n1598_n5888# 0.014014f
C681 source.n591 a_n1598_n5888# 0.033125f
C682 source.n592 a_n1598_n5888# 0.014839f
C683 source.n593 a_n1598_n5888# 0.02608f
C684 source.n594 a_n1598_n5888# 0.014014f
C685 source.n595 a_n1598_n5888# 0.033125f
C686 source.n596 a_n1598_n5888# 0.014839f
C687 source.n597 a_n1598_n5888# 0.02608f
C688 source.n598 a_n1598_n5888# 0.014014f
C689 source.n599 a_n1598_n5888# 0.033125f
C690 source.n600 a_n1598_n5888# 0.014839f
C691 source.n601 a_n1598_n5888# 0.02608f
C692 source.n602 a_n1598_n5888# 0.014427f
C693 source.n603 a_n1598_n5888# 0.033125f
C694 source.n604 a_n1598_n5888# 0.014839f
C695 source.n605 a_n1598_n5888# 0.02608f
C696 source.n606 a_n1598_n5888# 0.014014f
C697 source.n607 a_n1598_n5888# 0.033125f
C698 source.n608 a_n1598_n5888# 0.014839f
C699 source.n609 a_n1598_n5888# 0.02608f
C700 source.n610 a_n1598_n5888# 0.014014f
C701 source.n611 a_n1598_n5888# 0.024844f
C702 source.n612 a_n1598_n5888# 0.023417f
C703 source.t10 a_n1598_n5888# 0.057772f
C704 source.n613 a_n1598_n5888# 0.318202f
C705 source.n614 a_n1598_n5888# 2.82373f
C706 source.n615 a_n1598_n5888# 0.014014f
C707 source.n616 a_n1598_n5888# 0.014839f
C708 source.n617 a_n1598_n5888# 0.033125f
C709 source.n618 a_n1598_n5888# 0.033125f
C710 source.n619 a_n1598_n5888# 0.014839f
C711 source.n620 a_n1598_n5888# 0.014014f
C712 source.n621 a_n1598_n5888# 0.02608f
C713 source.n622 a_n1598_n5888# 0.02608f
C714 source.n623 a_n1598_n5888# 0.014014f
C715 source.n624 a_n1598_n5888# 0.014839f
C716 source.n625 a_n1598_n5888# 0.033125f
C717 source.n626 a_n1598_n5888# 0.033125f
C718 source.n627 a_n1598_n5888# 0.014839f
C719 source.n628 a_n1598_n5888# 0.014014f
C720 source.n629 a_n1598_n5888# 0.02608f
C721 source.n630 a_n1598_n5888# 0.02608f
C722 source.n631 a_n1598_n5888# 0.014014f
C723 source.n632 a_n1598_n5888# 0.014014f
C724 source.n633 a_n1598_n5888# 0.014839f
C725 source.n634 a_n1598_n5888# 0.033125f
C726 source.n635 a_n1598_n5888# 0.033125f
C727 source.n636 a_n1598_n5888# 0.033125f
C728 source.n637 a_n1598_n5888# 0.014427f
C729 source.n638 a_n1598_n5888# 0.014014f
C730 source.n639 a_n1598_n5888# 0.02608f
C731 source.n640 a_n1598_n5888# 0.02608f
C732 source.n641 a_n1598_n5888# 0.014014f
C733 source.n642 a_n1598_n5888# 0.014839f
C734 source.n643 a_n1598_n5888# 0.033125f
C735 source.n644 a_n1598_n5888# 0.033125f
C736 source.n645 a_n1598_n5888# 0.014839f
C737 source.n646 a_n1598_n5888# 0.014014f
C738 source.n647 a_n1598_n5888# 0.02608f
C739 source.n648 a_n1598_n5888# 0.02608f
C740 source.n649 a_n1598_n5888# 0.014014f
C741 source.n650 a_n1598_n5888# 0.014839f
C742 source.n651 a_n1598_n5888# 0.033125f
C743 source.n652 a_n1598_n5888# 0.033125f
C744 source.n653 a_n1598_n5888# 0.014839f
C745 source.n654 a_n1598_n5888# 0.014014f
C746 source.n655 a_n1598_n5888# 0.02608f
C747 source.n656 a_n1598_n5888# 0.02608f
C748 source.n657 a_n1598_n5888# 0.014014f
C749 source.n658 a_n1598_n5888# 0.014839f
C750 source.n659 a_n1598_n5888# 0.033125f
C751 source.n660 a_n1598_n5888# 0.033125f
C752 source.n661 a_n1598_n5888# 0.014839f
C753 source.n662 a_n1598_n5888# 0.014014f
C754 source.n663 a_n1598_n5888# 0.02608f
C755 source.n664 a_n1598_n5888# 0.02608f
C756 source.n665 a_n1598_n5888# 0.014014f
C757 source.n666 a_n1598_n5888# 0.014839f
C758 source.n667 a_n1598_n5888# 0.033125f
C759 source.n668 a_n1598_n5888# 0.033125f
C760 source.n669 a_n1598_n5888# 0.014839f
C761 source.n670 a_n1598_n5888# 0.014014f
C762 source.n671 a_n1598_n5888# 0.02608f
C763 source.n672 a_n1598_n5888# 0.02608f
C764 source.n673 a_n1598_n5888# 0.014014f
C765 source.n674 a_n1598_n5888# 0.014839f
C766 source.n675 a_n1598_n5888# 0.033125f
C767 source.n676 a_n1598_n5888# 0.033125f
C768 source.n677 a_n1598_n5888# 0.033125f
C769 source.n678 a_n1598_n5888# 0.014839f
C770 source.n679 a_n1598_n5888# 0.014014f
C771 source.n680 a_n1598_n5888# 0.02608f
C772 source.n681 a_n1598_n5888# 0.02608f
C773 source.n682 a_n1598_n5888# 0.014014f
C774 source.n683 a_n1598_n5888# 0.014427f
C775 source.n684 a_n1598_n5888# 0.014427f
C776 source.n685 a_n1598_n5888# 0.033125f
C777 source.n686 a_n1598_n5888# 0.033125f
C778 source.n687 a_n1598_n5888# 0.014839f
C779 source.n688 a_n1598_n5888# 0.014014f
C780 source.n689 a_n1598_n5888# 0.02608f
C781 source.n690 a_n1598_n5888# 0.02608f
C782 source.n691 a_n1598_n5888# 0.014014f
C783 source.n692 a_n1598_n5888# 0.014839f
C784 source.n693 a_n1598_n5888# 0.033125f
C785 source.n694 a_n1598_n5888# 0.033125f
C786 source.n695 a_n1598_n5888# 0.014839f
C787 source.n696 a_n1598_n5888# 0.014014f
C788 source.n697 a_n1598_n5888# 0.02608f
C789 source.n698 a_n1598_n5888# 0.02608f
C790 source.n699 a_n1598_n5888# 0.014014f
C791 source.n700 a_n1598_n5888# 0.014839f
C792 source.n701 a_n1598_n5888# 0.033125f
C793 source.n702 a_n1598_n5888# 0.070465f
C794 source.n703 a_n1598_n5888# 0.014839f
C795 source.n704 a_n1598_n5888# 0.014014f
C796 source.n705 a_n1598_n5888# 0.057433f
C797 source.n706 a_n1598_n5888# 0.039211f
C798 source.n707 a_n1598_n5888# 2.53218f
C799 source.t0 a_n1598_n5888# 0.515236f
C800 source.t3 a_n1598_n5888# 0.515236f
C801 source.n708 a_n1598_n5888# 4.66296f
C802 source.n709 a_n1598_n5888# 0.361787f
C803 source.t5 a_n1598_n5888# 0.515236f
C804 source.t1 a_n1598_n5888# 0.515236f
C805 source.n710 a_n1598_n5888# 4.66296f
C806 source.n711 a_n1598_n5888# 0.361787f
C807 source.n712 a_n1598_n5888# 0.035954f
C808 source.n713 a_n1598_n5888# 0.02608f
C809 source.n714 a_n1598_n5888# 0.014014f
C810 source.n715 a_n1598_n5888# 0.033125f
C811 source.n716 a_n1598_n5888# 0.014839f
C812 source.n717 a_n1598_n5888# 0.02608f
C813 source.n718 a_n1598_n5888# 0.014014f
C814 source.n719 a_n1598_n5888# 0.033125f
C815 source.n720 a_n1598_n5888# 0.014839f
C816 source.n721 a_n1598_n5888# 0.02608f
C817 source.n722 a_n1598_n5888# 0.014014f
C818 source.n723 a_n1598_n5888# 0.033125f
C819 source.n724 a_n1598_n5888# 0.014839f
C820 source.n725 a_n1598_n5888# 0.02608f
C821 source.n726 a_n1598_n5888# 0.014014f
C822 source.n727 a_n1598_n5888# 0.033125f
C823 source.n728 a_n1598_n5888# 0.014839f
C824 source.n729 a_n1598_n5888# 0.02608f
C825 source.n730 a_n1598_n5888# 0.014014f
C826 source.n731 a_n1598_n5888# 0.033125f
C827 source.n732 a_n1598_n5888# 0.014839f
C828 source.n733 a_n1598_n5888# 0.02608f
C829 source.n734 a_n1598_n5888# 0.014014f
C830 source.n735 a_n1598_n5888# 0.033125f
C831 source.n736 a_n1598_n5888# 0.014839f
C832 source.n737 a_n1598_n5888# 0.02608f
C833 source.n738 a_n1598_n5888# 0.014014f
C834 source.n739 a_n1598_n5888# 0.033125f
C835 source.n740 a_n1598_n5888# 0.014839f
C836 source.n741 a_n1598_n5888# 0.02608f
C837 source.n742 a_n1598_n5888# 0.014014f
C838 source.n743 a_n1598_n5888# 0.033125f
C839 source.n744 a_n1598_n5888# 0.014839f
C840 source.n745 a_n1598_n5888# 0.02608f
C841 source.n746 a_n1598_n5888# 0.014427f
C842 source.n747 a_n1598_n5888# 0.033125f
C843 source.n748 a_n1598_n5888# 0.014839f
C844 source.n749 a_n1598_n5888# 0.02608f
C845 source.n750 a_n1598_n5888# 0.014014f
C846 source.n751 a_n1598_n5888# 0.033125f
C847 source.n752 a_n1598_n5888# 0.014839f
C848 source.n753 a_n1598_n5888# 0.02608f
C849 source.n754 a_n1598_n5888# 0.014014f
C850 source.n755 a_n1598_n5888# 0.024844f
C851 source.n756 a_n1598_n5888# 0.023417f
C852 source.t6 a_n1598_n5888# 0.057772f
C853 source.n757 a_n1598_n5888# 0.318202f
C854 source.n758 a_n1598_n5888# 2.82373f
C855 source.n759 a_n1598_n5888# 0.014014f
C856 source.n760 a_n1598_n5888# 0.014839f
C857 source.n761 a_n1598_n5888# 0.033125f
C858 source.n762 a_n1598_n5888# 0.033125f
C859 source.n763 a_n1598_n5888# 0.014839f
C860 source.n764 a_n1598_n5888# 0.014014f
C861 source.n765 a_n1598_n5888# 0.02608f
C862 source.n766 a_n1598_n5888# 0.02608f
C863 source.n767 a_n1598_n5888# 0.014014f
C864 source.n768 a_n1598_n5888# 0.014839f
C865 source.n769 a_n1598_n5888# 0.033125f
C866 source.n770 a_n1598_n5888# 0.033125f
C867 source.n771 a_n1598_n5888# 0.014839f
C868 source.n772 a_n1598_n5888# 0.014014f
C869 source.n773 a_n1598_n5888# 0.02608f
C870 source.n774 a_n1598_n5888# 0.02608f
C871 source.n775 a_n1598_n5888# 0.014014f
C872 source.n776 a_n1598_n5888# 0.014014f
C873 source.n777 a_n1598_n5888# 0.014839f
C874 source.n778 a_n1598_n5888# 0.033125f
C875 source.n779 a_n1598_n5888# 0.033125f
C876 source.n780 a_n1598_n5888# 0.033125f
C877 source.n781 a_n1598_n5888# 0.014427f
C878 source.n782 a_n1598_n5888# 0.014014f
C879 source.n783 a_n1598_n5888# 0.02608f
C880 source.n784 a_n1598_n5888# 0.02608f
C881 source.n785 a_n1598_n5888# 0.014014f
C882 source.n786 a_n1598_n5888# 0.014839f
C883 source.n787 a_n1598_n5888# 0.033125f
C884 source.n788 a_n1598_n5888# 0.033125f
C885 source.n789 a_n1598_n5888# 0.014839f
C886 source.n790 a_n1598_n5888# 0.014014f
C887 source.n791 a_n1598_n5888# 0.02608f
C888 source.n792 a_n1598_n5888# 0.02608f
C889 source.n793 a_n1598_n5888# 0.014014f
C890 source.n794 a_n1598_n5888# 0.014839f
C891 source.n795 a_n1598_n5888# 0.033125f
C892 source.n796 a_n1598_n5888# 0.033125f
C893 source.n797 a_n1598_n5888# 0.014839f
C894 source.n798 a_n1598_n5888# 0.014014f
C895 source.n799 a_n1598_n5888# 0.02608f
C896 source.n800 a_n1598_n5888# 0.02608f
C897 source.n801 a_n1598_n5888# 0.014014f
C898 source.n802 a_n1598_n5888# 0.014839f
C899 source.n803 a_n1598_n5888# 0.033125f
C900 source.n804 a_n1598_n5888# 0.033125f
C901 source.n805 a_n1598_n5888# 0.014839f
C902 source.n806 a_n1598_n5888# 0.014014f
C903 source.n807 a_n1598_n5888# 0.02608f
C904 source.n808 a_n1598_n5888# 0.02608f
C905 source.n809 a_n1598_n5888# 0.014014f
C906 source.n810 a_n1598_n5888# 0.014839f
C907 source.n811 a_n1598_n5888# 0.033125f
C908 source.n812 a_n1598_n5888# 0.033125f
C909 source.n813 a_n1598_n5888# 0.014839f
C910 source.n814 a_n1598_n5888# 0.014014f
C911 source.n815 a_n1598_n5888# 0.02608f
C912 source.n816 a_n1598_n5888# 0.02608f
C913 source.n817 a_n1598_n5888# 0.014014f
C914 source.n818 a_n1598_n5888# 0.014839f
C915 source.n819 a_n1598_n5888# 0.033125f
C916 source.n820 a_n1598_n5888# 0.033125f
C917 source.n821 a_n1598_n5888# 0.033125f
C918 source.n822 a_n1598_n5888# 0.014839f
C919 source.n823 a_n1598_n5888# 0.014014f
C920 source.n824 a_n1598_n5888# 0.02608f
C921 source.n825 a_n1598_n5888# 0.02608f
C922 source.n826 a_n1598_n5888# 0.014014f
C923 source.n827 a_n1598_n5888# 0.014427f
C924 source.n828 a_n1598_n5888# 0.014427f
C925 source.n829 a_n1598_n5888# 0.033125f
C926 source.n830 a_n1598_n5888# 0.033125f
C927 source.n831 a_n1598_n5888# 0.014839f
C928 source.n832 a_n1598_n5888# 0.014014f
C929 source.n833 a_n1598_n5888# 0.02608f
C930 source.n834 a_n1598_n5888# 0.02608f
C931 source.n835 a_n1598_n5888# 0.014014f
C932 source.n836 a_n1598_n5888# 0.014839f
C933 source.n837 a_n1598_n5888# 0.033125f
C934 source.n838 a_n1598_n5888# 0.033125f
C935 source.n839 a_n1598_n5888# 0.014839f
C936 source.n840 a_n1598_n5888# 0.014014f
C937 source.n841 a_n1598_n5888# 0.02608f
C938 source.n842 a_n1598_n5888# 0.02608f
C939 source.n843 a_n1598_n5888# 0.014014f
C940 source.n844 a_n1598_n5888# 0.014839f
C941 source.n845 a_n1598_n5888# 0.033125f
C942 source.n846 a_n1598_n5888# 0.070465f
C943 source.n847 a_n1598_n5888# 0.014839f
C944 source.n848 a_n1598_n5888# 0.014014f
C945 source.n849 a_n1598_n5888# 0.057433f
C946 source.n850 a_n1598_n5888# 0.039211f
C947 source.n851 a_n1598_n5888# 0.105791f
C948 source.n852 a_n1598_n5888# 0.035954f
C949 source.n853 a_n1598_n5888# 0.02608f
C950 source.n854 a_n1598_n5888# 0.014014f
C951 source.n855 a_n1598_n5888# 0.033125f
C952 source.n856 a_n1598_n5888# 0.014839f
C953 source.n857 a_n1598_n5888# 0.02608f
C954 source.n858 a_n1598_n5888# 0.014014f
C955 source.n859 a_n1598_n5888# 0.033125f
C956 source.n860 a_n1598_n5888# 0.014839f
C957 source.n861 a_n1598_n5888# 0.02608f
C958 source.n862 a_n1598_n5888# 0.014014f
C959 source.n863 a_n1598_n5888# 0.033125f
C960 source.n864 a_n1598_n5888# 0.014839f
C961 source.n865 a_n1598_n5888# 0.02608f
C962 source.n866 a_n1598_n5888# 0.014014f
C963 source.n867 a_n1598_n5888# 0.033125f
C964 source.n868 a_n1598_n5888# 0.014839f
C965 source.n869 a_n1598_n5888# 0.02608f
C966 source.n870 a_n1598_n5888# 0.014014f
C967 source.n871 a_n1598_n5888# 0.033125f
C968 source.n872 a_n1598_n5888# 0.014839f
C969 source.n873 a_n1598_n5888# 0.02608f
C970 source.n874 a_n1598_n5888# 0.014014f
C971 source.n875 a_n1598_n5888# 0.033125f
C972 source.n876 a_n1598_n5888# 0.014839f
C973 source.n877 a_n1598_n5888# 0.02608f
C974 source.n878 a_n1598_n5888# 0.014014f
C975 source.n879 a_n1598_n5888# 0.033125f
C976 source.n880 a_n1598_n5888# 0.014839f
C977 source.n881 a_n1598_n5888# 0.02608f
C978 source.n882 a_n1598_n5888# 0.014014f
C979 source.n883 a_n1598_n5888# 0.033125f
C980 source.n884 a_n1598_n5888# 0.014839f
C981 source.n885 a_n1598_n5888# 0.02608f
C982 source.n886 a_n1598_n5888# 0.014427f
C983 source.n887 a_n1598_n5888# 0.033125f
C984 source.n888 a_n1598_n5888# 0.014839f
C985 source.n889 a_n1598_n5888# 0.02608f
C986 source.n890 a_n1598_n5888# 0.014014f
C987 source.n891 a_n1598_n5888# 0.033125f
C988 source.n892 a_n1598_n5888# 0.014839f
C989 source.n893 a_n1598_n5888# 0.02608f
C990 source.n894 a_n1598_n5888# 0.014014f
C991 source.n895 a_n1598_n5888# 0.024844f
C992 source.n896 a_n1598_n5888# 0.023417f
C993 source.t20 a_n1598_n5888# 0.057772f
C994 source.n897 a_n1598_n5888# 0.318202f
C995 source.n898 a_n1598_n5888# 2.82373f
C996 source.n899 a_n1598_n5888# 0.014014f
C997 source.n900 a_n1598_n5888# 0.014839f
C998 source.n901 a_n1598_n5888# 0.033125f
C999 source.n902 a_n1598_n5888# 0.033125f
C1000 source.n903 a_n1598_n5888# 0.014839f
C1001 source.n904 a_n1598_n5888# 0.014014f
C1002 source.n905 a_n1598_n5888# 0.02608f
C1003 source.n906 a_n1598_n5888# 0.02608f
C1004 source.n907 a_n1598_n5888# 0.014014f
C1005 source.n908 a_n1598_n5888# 0.014839f
C1006 source.n909 a_n1598_n5888# 0.033125f
C1007 source.n910 a_n1598_n5888# 0.033125f
C1008 source.n911 a_n1598_n5888# 0.014839f
C1009 source.n912 a_n1598_n5888# 0.014014f
C1010 source.n913 a_n1598_n5888# 0.02608f
C1011 source.n914 a_n1598_n5888# 0.02608f
C1012 source.n915 a_n1598_n5888# 0.014014f
C1013 source.n916 a_n1598_n5888# 0.014014f
C1014 source.n917 a_n1598_n5888# 0.014839f
C1015 source.n918 a_n1598_n5888# 0.033125f
C1016 source.n919 a_n1598_n5888# 0.033125f
C1017 source.n920 a_n1598_n5888# 0.033125f
C1018 source.n921 a_n1598_n5888# 0.014427f
C1019 source.n922 a_n1598_n5888# 0.014014f
C1020 source.n923 a_n1598_n5888# 0.02608f
C1021 source.n924 a_n1598_n5888# 0.02608f
C1022 source.n925 a_n1598_n5888# 0.014014f
C1023 source.n926 a_n1598_n5888# 0.014839f
C1024 source.n927 a_n1598_n5888# 0.033125f
C1025 source.n928 a_n1598_n5888# 0.033125f
C1026 source.n929 a_n1598_n5888# 0.014839f
C1027 source.n930 a_n1598_n5888# 0.014014f
C1028 source.n931 a_n1598_n5888# 0.02608f
C1029 source.n932 a_n1598_n5888# 0.02608f
C1030 source.n933 a_n1598_n5888# 0.014014f
C1031 source.n934 a_n1598_n5888# 0.014839f
C1032 source.n935 a_n1598_n5888# 0.033125f
C1033 source.n936 a_n1598_n5888# 0.033125f
C1034 source.n937 a_n1598_n5888# 0.014839f
C1035 source.n938 a_n1598_n5888# 0.014014f
C1036 source.n939 a_n1598_n5888# 0.02608f
C1037 source.n940 a_n1598_n5888# 0.02608f
C1038 source.n941 a_n1598_n5888# 0.014014f
C1039 source.n942 a_n1598_n5888# 0.014839f
C1040 source.n943 a_n1598_n5888# 0.033125f
C1041 source.n944 a_n1598_n5888# 0.033125f
C1042 source.n945 a_n1598_n5888# 0.014839f
C1043 source.n946 a_n1598_n5888# 0.014014f
C1044 source.n947 a_n1598_n5888# 0.02608f
C1045 source.n948 a_n1598_n5888# 0.02608f
C1046 source.n949 a_n1598_n5888# 0.014014f
C1047 source.n950 a_n1598_n5888# 0.014839f
C1048 source.n951 a_n1598_n5888# 0.033125f
C1049 source.n952 a_n1598_n5888# 0.033125f
C1050 source.n953 a_n1598_n5888# 0.014839f
C1051 source.n954 a_n1598_n5888# 0.014014f
C1052 source.n955 a_n1598_n5888# 0.02608f
C1053 source.n956 a_n1598_n5888# 0.02608f
C1054 source.n957 a_n1598_n5888# 0.014014f
C1055 source.n958 a_n1598_n5888# 0.014839f
C1056 source.n959 a_n1598_n5888# 0.033125f
C1057 source.n960 a_n1598_n5888# 0.033125f
C1058 source.n961 a_n1598_n5888# 0.033125f
C1059 source.n962 a_n1598_n5888# 0.014839f
C1060 source.n963 a_n1598_n5888# 0.014014f
C1061 source.n964 a_n1598_n5888# 0.02608f
C1062 source.n965 a_n1598_n5888# 0.02608f
C1063 source.n966 a_n1598_n5888# 0.014014f
C1064 source.n967 a_n1598_n5888# 0.014427f
C1065 source.n968 a_n1598_n5888# 0.014427f
C1066 source.n969 a_n1598_n5888# 0.033125f
C1067 source.n970 a_n1598_n5888# 0.033125f
C1068 source.n971 a_n1598_n5888# 0.014839f
C1069 source.n972 a_n1598_n5888# 0.014014f
C1070 source.n973 a_n1598_n5888# 0.02608f
C1071 source.n974 a_n1598_n5888# 0.02608f
C1072 source.n975 a_n1598_n5888# 0.014014f
C1073 source.n976 a_n1598_n5888# 0.014839f
C1074 source.n977 a_n1598_n5888# 0.033125f
C1075 source.n978 a_n1598_n5888# 0.033125f
C1076 source.n979 a_n1598_n5888# 0.014839f
C1077 source.n980 a_n1598_n5888# 0.014014f
C1078 source.n981 a_n1598_n5888# 0.02608f
C1079 source.n982 a_n1598_n5888# 0.02608f
C1080 source.n983 a_n1598_n5888# 0.014014f
C1081 source.n984 a_n1598_n5888# 0.014839f
C1082 source.n985 a_n1598_n5888# 0.033125f
C1083 source.n986 a_n1598_n5888# 0.070465f
C1084 source.n987 a_n1598_n5888# 0.014839f
C1085 source.n988 a_n1598_n5888# 0.014014f
C1086 source.n989 a_n1598_n5888# 0.057433f
C1087 source.n990 a_n1598_n5888# 0.039211f
C1088 source.n991 a_n1598_n5888# 0.105791f
C1089 source.t15 a_n1598_n5888# 0.515236f
C1090 source.t21 a_n1598_n5888# 0.515236f
C1091 source.n992 a_n1598_n5888# 4.66296f
C1092 source.n993 a_n1598_n5888# 0.361787f
C1093 source.t16 a_n1598_n5888# 0.515236f
C1094 source.t19 a_n1598_n5888# 0.515236f
C1095 source.n994 a_n1598_n5888# 4.66296f
C1096 source.n995 a_n1598_n5888# 0.361787f
C1097 source.n996 a_n1598_n5888# 0.035954f
C1098 source.n997 a_n1598_n5888# 0.02608f
C1099 source.n998 a_n1598_n5888# 0.014014f
C1100 source.n999 a_n1598_n5888# 0.033125f
C1101 source.n1000 a_n1598_n5888# 0.014839f
C1102 source.n1001 a_n1598_n5888# 0.02608f
C1103 source.n1002 a_n1598_n5888# 0.014014f
C1104 source.n1003 a_n1598_n5888# 0.033125f
C1105 source.n1004 a_n1598_n5888# 0.014839f
C1106 source.n1005 a_n1598_n5888# 0.02608f
C1107 source.n1006 a_n1598_n5888# 0.014014f
C1108 source.n1007 a_n1598_n5888# 0.033125f
C1109 source.n1008 a_n1598_n5888# 0.014839f
C1110 source.n1009 a_n1598_n5888# 0.02608f
C1111 source.n1010 a_n1598_n5888# 0.014014f
C1112 source.n1011 a_n1598_n5888# 0.033125f
C1113 source.n1012 a_n1598_n5888# 0.014839f
C1114 source.n1013 a_n1598_n5888# 0.02608f
C1115 source.n1014 a_n1598_n5888# 0.014014f
C1116 source.n1015 a_n1598_n5888# 0.033125f
C1117 source.n1016 a_n1598_n5888# 0.014839f
C1118 source.n1017 a_n1598_n5888# 0.02608f
C1119 source.n1018 a_n1598_n5888# 0.014014f
C1120 source.n1019 a_n1598_n5888# 0.033125f
C1121 source.n1020 a_n1598_n5888# 0.014839f
C1122 source.n1021 a_n1598_n5888# 0.02608f
C1123 source.n1022 a_n1598_n5888# 0.014014f
C1124 source.n1023 a_n1598_n5888# 0.033125f
C1125 source.n1024 a_n1598_n5888# 0.014839f
C1126 source.n1025 a_n1598_n5888# 0.02608f
C1127 source.n1026 a_n1598_n5888# 0.014014f
C1128 source.n1027 a_n1598_n5888# 0.033125f
C1129 source.n1028 a_n1598_n5888# 0.014839f
C1130 source.n1029 a_n1598_n5888# 0.02608f
C1131 source.n1030 a_n1598_n5888# 0.014427f
C1132 source.n1031 a_n1598_n5888# 0.033125f
C1133 source.n1032 a_n1598_n5888# 0.014839f
C1134 source.n1033 a_n1598_n5888# 0.02608f
C1135 source.n1034 a_n1598_n5888# 0.014014f
C1136 source.n1035 a_n1598_n5888# 0.033125f
C1137 source.n1036 a_n1598_n5888# 0.014839f
C1138 source.n1037 a_n1598_n5888# 0.02608f
C1139 source.n1038 a_n1598_n5888# 0.014014f
C1140 source.n1039 a_n1598_n5888# 0.024844f
C1141 source.n1040 a_n1598_n5888# 0.023417f
C1142 source.t12 a_n1598_n5888# 0.057772f
C1143 source.n1041 a_n1598_n5888# 0.318202f
C1144 source.n1042 a_n1598_n5888# 2.82373f
C1145 source.n1043 a_n1598_n5888# 0.014014f
C1146 source.n1044 a_n1598_n5888# 0.014839f
C1147 source.n1045 a_n1598_n5888# 0.033125f
C1148 source.n1046 a_n1598_n5888# 0.033125f
C1149 source.n1047 a_n1598_n5888# 0.014839f
C1150 source.n1048 a_n1598_n5888# 0.014014f
C1151 source.n1049 a_n1598_n5888# 0.02608f
C1152 source.n1050 a_n1598_n5888# 0.02608f
C1153 source.n1051 a_n1598_n5888# 0.014014f
C1154 source.n1052 a_n1598_n5888# 0.014839f
C1155 source.n1053 a_n1598_n5888# 0.033125f
C1156 source.n1054 a_n1598_n5888# 0.033125f
C1157 source.n1055 a_n1598_n5888# 0.014839f
C1158 source.n1056 a_n1598_n5888# 0.014014f
C1159 source.n1057 a_n1598_n5888# 0.02608f
C1160 source.n1058 a_n1598_n5888# 0.02608f
C1161 source.n1059 a_n1598_n5888# 0.014014f
C1162 source.n1060 a_n1598_n5888# 0.014014f
C1163 source.n1061 a_n1598_n5888# 0.014839f
C1164 source.n1062 a_n1598_n5888# 0.033125f
C1165 source.n1063 a_n1598_n5888# 0.033125f
C1166 source.n1064 a_n1598_n5888# 0.033125f
C1167 source.n1065 a_n1598_n5888# 0.014427f
C1168 source.n1066 a_n1598_n5888# 0.014014f
C1169 source.n1067 a_n1598_n5888# 0.02608f
C1170 source.n1068 a_n1598_n5888# 0.02608f
C1171 source.n1069 a_n1598_n5888# 0.014014f
C1172 source.n1070 a_n1598_n5888# 0.014839f
C1173 source.n1071 a_n1598_n5888# 0.033125f
C1174 source.n1072 a_n1598_n5888# 0.033125f
C1175 source.n1073 a_n1598_n5888# 0.014839f
C1176 source.n1074 a_n1598_n5888# 0.014014f
C1177 source.n1075 a_n1598_n5888# 0.02608f
C1178 source.n1076 a_n1598_n5888# 0.02608f
C1179 source.n1077 a_n1598_n5888# 0.014014f
C1180 source.n1078 a_n1598_n5888# 0.014839f
C1181 source.n1079 a_n1598_n5888# 0.033125f
C1182 source.n1080 a_n1598_n5888# 0.033125f
C1183 source.n1081 a_n1598_n5888# 0.014839f
C1184 source.n1082 a_n1598_n5888# 0.014014f
C1185 source.n1083 a_n1598_n5888# 0.02608f
C1186 source.n1084 a_n1598_n5888# 0.02608f
C1187 source.n1085 a_n1598_n5888# 0.014014f
C1188 source.n1086 a_n1598_n5888# 0.014839f
C1189 source.n1087 a_n1598_n5888# 0.033125f
C1190 source.n1088 a_n1598_n5888# 0.033125f
C1191 source.n1089 a_n1598_n5888# 0.014839f
C1192 source.n1090 a_n1598_n5888# 0.014014f
C1193 source.n1091 a_n1598_n5888# 0.02608f
C1194 source.n1092 a_n1598_n5888# 0.02608f
C1195 source.n1093 a_n1598_n5888# 0.014014f
C1196 source.n1094 a_n1598_n5888# 0.014839f
C1197 source.n1095 a_n1598_n5888# 0.033125f
C1198 source.n1096 a_n1598_n5888# 0.033125f
C1199 source.n1097 a_n1598_n5888# 0.014839f
C1200 source.n1098 a_n1598_n5888# 0.014014f
C1201 source.n1099 a_n1598_n5888# 0.02608f
C1202 source.n1100 a_n1598_n5888# 0.02608f
C1203 source.n1101 a_n1598_n5888# 0.014014f
C1204 source.n1102 a_n1598_n5888# 0.014839f
C1205 source.n1103 a_n1598_n5888# 0.033125f
C1206 source.n1104 a_n1598_n5888# 0.033125f
C1207 source.n1105 a_n1598_n5888# 0.033125f
C1208 source.n1106 a_n1598_n5888# 0.014839f
C1209 source.n1107 a_n1598_n5888# 0.014014f
C1210 source.n1108 a_n1598_n5888# 0.02608f
C1211 source.n1109 a_n1598_n5888# 0.02608f
C1212 source.n1110 a_n1598_n5888# 0.014014f
C1213 source.n1111 a_n1598_n5888# 0.014427f
C1214 source.n1112 a_n1598_n5888# 0.014427f
C1215 source.n1113 a_n1598_n5888# 0.033125f
C1216 source.n1114 a_n1598_n5888# 0.033125f
C1217 source.n1115 a_n1598_n5888# 0.014839f
C1218 source.n1116 a_n1598_n5888# 0.014014f
C1219 source.n1117 a_n1598_n5888# 0.02608f
C1220 source.n1118 a_n1598_n5888# 0.02608f
C1221 source.n1119 a_n1598_n5888# 0.014014f
C1222 source.n1120 a_n1598_n5888# 0.014839f
C1223 source.n1121 a_n1598_n5888# 0.033125f
C1224 source.n1122 a_n1598_n5888# 0.033125f
C1225 source.n1123 a_n1598_n5888# 0.014839f
C1226 source.n1124 a_n1598_n5888# 0.014014f
C1227 source.n1125 a_n1598_n5888# 0.02608f
C1228 source.n1126 a_n1598_n5888# 0.02608f
C1229 source.n1127 a_n1598_n5888# 0.014014f
C1230 source.n1128 a_n1598_n5888# 0.014839f
C1231 source.n1129 a_n1598_n5888# 0.033125f
C1232 source.n1130 a_n1598_n5888# 0.070465f
C1233 source.n1131 a_n1598_n5888# 0.014839f
C1234 source.n1132 a_n1598_n5888# 0.014014f
C1235 source.n1133 a_n1598_n5888# 0.057433f
C1236 source.n1134 a_n1598_n5888# 0.039211f
C1237 source.n1135 a_n1598_n5888# 0.253014f
C1238 source.n1136 a_n1598_n5888# 2.7802f
C1239 drain_right.t4 a_n1598_n5888# 0.675292f
C1240 drain_right.t9 a_n1598_n5888# 0.675292f
C1241 drain_right.n0 a_n1598_n5888# 6.22698f
C1242 drain_right.t5 a_n1598_n5888# 0.675292f
C1243 drain_right.t2 a_n1598_n5888# 0.675292f
C1244 drain_right.n1 a_n1598_n5888# 6.22354f
C1245 drain_right.t7 a_n1598_n5888# 0.675292f
C1246 drain_right.t10 a_n1598_n5888# 0.675292f
C1247 drain_right.n2 a_n1598_n5888# 6.22698f
C1248 drain_right.n3 a_n1598_n5888# 3.8179f
C1249 drain_right.t11 a_n1598_n5888# 0.675292f
C1250 drain_right.t3 a_n1598_n5888# 0.675292f
C1251 drain_right.n4 a_n1598_n5888# 6.2274f
C1252 drain_right.t6 a_n1598_n5888# 0.675292f
C1253 drain_right.t0 a_n1598_n5888# 0.675292f
C1254 drain_right.n5 a_n1598_n5888# 6.22354f
C1255 drain_right.n6 a_n1598_n5888# 0.827058f
C1256 drain_right.t1 a_n1598_n5888# 0.675292f
C1257 drain_right.t8 a_n1598_n5888# 0.675292f
C1258 drain_right.n7 a_n1598_n5888# 6.22354f
C1259 drain_right.n8 a_n1598_n5888# 0.693091f
C1260 minus.n0 a_n1598_n5888# 0.052808f
C1261 minus.t0 a_n1598_n5888# 1.12339f
C1262 minus.t9 a_n1598_n5888# 1.11439f
C1263 minus.t5 a_n1598_n5888# 1.11439f
C1264 minus.n1 a_n1598_n5888# 0.019635f
C1265 minus.t6 a_n1598_n5888# 1.12339f
C1266 minus.n2 a_n1598_n5888# 0.422401f
C1267 minus.t1 a_n1598_n5888# 1.11439f
C1268 minus.n3 a_n1598_n5888# 0.405502f
C1269 minus.t10 a_n1598_n5888# 1.11439f
C1270 minus.n4 a_n1598_n5888# 0.405502f
C1271 minus.n5 a_n1598_n5888# 0.021751f
C1272 minus.n6 a_n1598_n5888# 0.120189f
C1273 minus.n7 a_n1598_n5888# 0.052808f
C1274 minus.n8 a_n1598_n5888# 0.052808f
C1275 minus.n9 a_n1598_n5888# 0.019635f
C1276 minus.n10 a_n1598_n5888# 0.405502f
C1277 minus.n11 a_n1598_n5888# 0.021751f
C1278 minus.n12 a_n1598_n5888# 0.405502f
C1279 minus.n13 a_n1598_n5888# 0.422322f
C1280 minus.n14 a_n1598_n5888# 2.58871f
C1281 minus.n15 a_n1598_n5888# 0.052808f
C1282 minus.t4 a_n1598_n5888# 1.11439f
C1283 minus.t7 a_n1598_n5888# 1.11439f
C1284 minus.n16 a_n1598_n5888# 0.019635f
C1285 minus.t3 a_n1598_n5888# 1.12339f
C1286 minus.n17 a_n1598_n5888# 0.422401f
C1287 minus.t8 a_n1598_n5888# 1.11439f
C1288 minus.n18 a_n1598_n5888# 0.405502f
C1289 minus.t2 a_n1598_n5888# 1.11439f
C1290 minus.n19 a_n1598_n5888# 0.405502f
C1291 minus.n20 a_n1598_n5888# 0.021751f
C1292 minus.n21 a_n1598_n5888# 0.120189f
C1293 minus.n22 a_n1598_n5888# 0.052808f
C1294 minus.n23 a_n1598_n5888# 0.052808f
C1295 minus.n24 a_n1598_n5888# 0.019635f
C1296 minus.n25 a_n1598_n5888# 0.405502f
C1297 minus.n26 a_n1598_n5888# 0.021751f
C1298 minus.n27 a_n1598_n5888# 0.405502f
C1299 minus.t11 a_n1598_n5888# 1.12339f
C1300 minus.n28 a_n1598_n5888# 0.422322f
C1301 minus.n29 a_n1598_n5888# 0.346722f
C1302 minus.n30 a_n1598_n5888# 3.06499f
.ends

