* NGSPICE file created from diffpair233.ext - technology: sky130A

.subckt diffpair233 minus drain_right drain_left source plus
X0 source.t15 minus.t0 drain_right.t2 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X1 source.t14 minus.t1 drain_right.t7 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X2 a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X3 drain_left.t7 plus.t0 source.t7 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X4 drain_left.t6 plus.t1 source.t2 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X5 a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X6 a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X7 a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X8 drain_right.t5 minus.t2 source.t13 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X9 drain_right.t4 minus.t3 source.t12 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X10 source.t11 minus.t4 drain_right.t3 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X11 drain_right.t1 minus.t5 source.t10 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X12 drain_right.t0 minus.t6 source.t9 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X13 source.t4 plus.t2 drain_left.t5 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X14 source.t8 minus.t7 drain_right.t6 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X15 source.t3 plus.t3 drain_left.t4 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X16 drain_left.t3 plus.t4 source.t1 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X17 source.t6 plus.t5 drain_left.t2 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X18 drain_left.t1 plus.t6 source.t5 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 source.t0 plus.t7 drain_left.t0 a_n1846_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
R0 minus.n7 minus.n6 161.3
R1 minus.n5 minus.n0 161.3
R2 minus.n15 minus.n14 161.3
R3 minus.n13 minus.n8 161.3
R4 minus.n2 minus.t6 160.082
R5 minus.n10 minus.t0 160.082
R6 minus.n1 minus.t4 139.48
R7 minus.n4 minus.t2 139.48
R8 minus.n6 minus.t7 139.48
R9 minus.n9 minus.t3 139.48
R10 minus.n12 minus.t1 139.48
R11 minus.n14 minus.t5 139.48
R12 minus.n4 minus.n3 80.6037
R13 minus.n12 minus.n11 80.6037
R14 minus.n4 minus.n1 48.2005
R15 minus.n12 minus.n9 48.2005
R16 minus.n5 minus.n4 41.6278
R17 minus.n13 minus.n12 41.6278
R18 minus.n3 minus.n2 31.6158
R19 minus.n11 minus.n10 31.6158
R20 minus.n16 minus.n7 29.4475
R21 minus.n2 minus.n1 17.6494
R22 minus.n10 minus.n9 17.6494
R23 minus.n16 minus.n15 6.65202
R24 minus.n6 minus.n5 6.57323
R25 minus.n14 minus.n13 6.57323
R26 minus.n3 minus.n0 0.285035
R27 minus.n11 minus.n8 0.285035
R28 minus.n7 minus.n0 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 drain_right.n5 drain_right.n3 80.7472
R32 drain_right.n2 drain_right.n1 80.2047
R33 drain_right.n2 drain_right.n0 80.2047
R34 drain_right.n5 drain_right.n4 79.7731
R35 drain_right drain_right.n2 23.4051
R36 drain_right drain_right.n5 6.62735
R37 drain_right.n1 drain_right.t7 6.6005
R38 drain_right.n1 drain_right.t1 6.6005
R39 drain_right.n0 drain_right.t2 6.6005
R40 drain_right.n0 drain_right.t4 6.6005
R41 drain_right.n3 drain_right.t3 6.6005
R42 drain_right.n3 drain_right.t0 6.6005
R43 drain_right.n4 drain_right.t6 6.6005
R44 drain_right.n4 drain_right.t5 6.6005
R45 source.n0 source.t1 69.6943
R46 source.n3 source.t0 69.6943
R47 source.n4 source.t9 69.6943
R48 source.n7 source.t8 69.6943
R49 source.n15 source.t10 69.6942
R50 source.n12 source.t15 69.6942
R51 source.n11 source.t7 69.6942
R52 source.n8 source.t3 69.6942
R53 source.n2 source.n1 63.0943
R54 source.n6 source.n5 63.0943
R55 source.n14 source.n13 63.0942
R56 source.n10 source.n9 63.0942
R57 source.n8 source.n7 15.4437
R58 source.n16 source.n0 9.69368
R59 source.n13 source.t12 6.6005
R60 source.n13 source.t14 6.6005
R61 source.n9 source.t2 6.6005
R62 source.n9 source.t4 6.6005
R63 source.n1 source.t5 6.6005
R64 source.n1 source.t6 6.6005
R65 source.n5 source.t13 6.6005
R66 source.n5 source.t11 6.6005
R67 source.n16 source.n15 5.7505
R68 source.n7 source.n6 0.974638
R69 source.n6 source.n4 0.974638
R70 source.n3 source.n2 0.974638
R71 source.n2 source.n0 0.974638
R72 source.n10 source.n8 0.974638
R73 source.n11 source.n10 0.974638
R74 source.n14 source.n12 0.974638
R75 source.n15 source.n14 0.974638
R76 source.n4 source.n3 0.470328
R77 source.n12 source.n11 0.470328
R78 source source.n16 0.188
R79 plus.n5 plus.n0 161.3
R80 plus.n7 plus.n6 161.3
R81 plus.n13 plus.n8 161.3
R82 plus.n15 plus.n14 161.3
R83 plus.n2 plus.t7 160.082
R84 plus.n10 plus.t0 160.082
R85 plus.n6 plus.t4 139.48
R86 plus.n4 plus.t5 139.48
R87 plus.n3 plus.t6 139.48
R88 plus.n14 plus.t3 139.48
R89 plus.n12 plus.t1 139.48
R90 plus.n11 plus.t2 139.48
R91 plus.n4 plus.n1 80.6037
R92 plus.n12 plus.n9 80.6037
R93 plus.n4 plus.n3 48.2005
R94 plus.n12 plus.n11 48.2005
R95 plus.n5 plus.n4 41.6278
R96 plus.n13 plus.n12 41.6278
R97 plus.n2 plus.n1 31.6158
R98 plus.n10 plus.n9 31.6158
R99 plus plus.n15 26.7377
R100 plus.n3 plus.n2 17.6494
R101 plus.n11 plus.n10 17.6494
R102 plus plus.n7 8.88686
R103 plus.n6 plus.n5 6.57323
R104 plus.n14 plus.n13 6.57323
R105 plus.n1 plus.n0 0.285035
R106 plus.n9 plus.n8 0.285035
R107 plus.n7 plus.n0 0.189894
R108 plus.n15 plus.n8 0.189894
R109 drain_left.n5 drain_left.n3 80.7472
R110 drain_left.n2 drain_left.n1 80.2047
R111 drain_left.n2 drain_left.n0 80.2047
R112 drain_left.n5 drain_left.n4 79.7731
R113 drain_left drain_left.n2 23.9584
R114 drain_left drain_left.n5 6.62735
R115 drain_left.n1 drain_left.t5 6.6005
R116 drain_left.n1 drain_left.t7 6.6005
R117 drain_left.n0 drain_left.t4 6.6005
R118 drain_left.n0 drain_left.t6 6.6005
R119 drain_left.n4 drain_left.t2 6.6005
R120 drain_left.n4 drain_left.t3 6.6005
R121 drain_left.n3 drain_left.t0 6.6005
R122 drain_left.n3 drain_left.t1 6.6005
C0 drain_left plus 1.95129f
C1 source drain_left 4.35266f
C2 minus drain_right 1.77208f
C3 minus plus 3.78307f
C4 source minus 2.02272f
C5 drain_right plus 0.339415f
C6 source drain_right 4.35505f
C7 source plus 2.03671f
C8 minus drain_left 0.176511f
C9 drain_right drain_left 0.873724f
C10 drain_right a_n1846_n1488# 3.52815f
C11 drain_left a_n1846_n1488# 3.75437f
C12 source a_n1846_n1488# 3.728586f
C13 minus a_n1846_n1488# 6.425112f
C14 plus a_n1846_n1488# 7.28147f
C15 drain_left.t4 a_n1846_n1488# 0.042842f
C16 drain_left.t6 a_n1846_n1488# 0.042842f
C17 drain_left.n0 a_n1846_n1488# 0.310233f
C18 drain_left.t5 a_n1846_n1488# 0.042842f
C19 drain_left.t7 a_n1846_n1488# 0.042842f
C20 drain_left.n1 a_n1846_n1488# 0.310233f
C21 drain_left.n2 a_n1846_n1488# 1.03489f
C22 drain_left.t0 a_n1846_n1488# 0.042842f
C23 drain_left.t1 a_n1846_n1488# 0.042842f
C24 drain_left.n3 a_n1846_n1488# 0.312173f
C25 drain_left.t2 a_n1846_n1488# 0.042842f
C26 drain_left.t3 a_n1846_n1488# 0.042842f
C27 drain_left.n4 a_n1846_n1488# 0.308971f
C28 drain_left.n5 a_n1846_n1488# 0.682332f
C29 plus.n0 a_n1846_n1488# 0.046005f
C30 plus.t4 a_n1846_n1488# 0.248123f
C31 plus.t5 a_n1846_n1488# 0.248123f
C32 plus.n1 a_n1846_n1488# 0.197324f
C33 plus.t6 a_n1846_n1488# 0.248123f
C34 plus.t7 a_n1846_n1488# 0.266719f
C35 plus.n2 a_n1846_n1488# 0.12878f
C36 plus.n3 a_n1846_n1488# 0.151552f
C37 plus.n4 a_n1846_n1488# 0.150991f
C38 plus.n5 a_n1846_n1488# 0.007824f
C39 plus.n6 a_n1846_n1488# 0.138065f
C40 plus.n7 a_n1846_n1488# 0.270458f
C41 plus.n8 a_n1846_n1488# 0.046005f
C42 plus.t3 a_n1846_n1488# 0.248123f
C43 plus.n9 a_n1846_n1488# 0.197324f
C44 plus.t1 a_n1846_n1488# 0.248123f
C45 plus.t0 a_n1846_n1488# 0.266719f
C46 plus.n10 a_n1846_n1488# 0.12878f
C47 plus.t2 a_n1846_n1488# 0.248123f
C48 plus.n11 a_n1846_n1488# 0.151552f
C49 plus.n12 a_n1846_n1488# 0.150991f
C50 plus.n13 a_n1846_n1488# 0.007824f
C51 plus.n14 a_n1846_n1488# 0.138065f
C52 plus.n15 a_n1846_n1488# 0.822438f
C53 source.t1 a_n1846_n1488# 0.484696f
C54 source.n0 a_n1846_n1488# 0.721317f
C55 source.t5 a_n1846_n1488# 0.05837f
C56 source.t6 a_n1846_n1488# 0.05837f
C57 source.n1 a_n1846_n1488# 0.370101f
C58 source.n2 a_n1846_n1488# 0.369055f
C59 source.t0 a_n1846_n1488# 0.484696f
C60 source.n3 a_n1846_n1488# 0.373641f
C61 source.t9 a_n1846_n1488# 0.484696f
C62 source.n4 a_n1846_n1488# 0.373641f
C63 source.t13 a_n1846_n1488# 0.05837f
C64 source.t11 a_n1846_n1488# 0.05837f
C65 source.n5 a_n1846_n1488# 0.370101f
C66 source.n6 a_n1846_n1488# 0.369055f
C67 source.t8 a_n1846_n1488# 0.484696f
C68 source.n7 a_n1846_n1488# 0.986329f
C69 source.t3 a_n1846_n1488# 0.484694f
C70 source.n8 a_n1846_n1488# 0.986331f
C71 source.t2 a_n1846_n1488# 0.05837f
C72 source.t4 a_n1846_n1488# 0.05837f
C73 source.n9 a_n1846_n1488# 0.370098f
C74 source.n10 a_n1846_n1488# 0.369058f
C75 source.t7 a_n1846_n1488# 0.484694f
C76 source.n11 a_n1846_n1488# 0.373644f
C77 source.t15 a_n1846_n1488# 0.484694f
C78 source.n12 a_n1846_n1488# 0.373644f
C79 source.t12 a_n1846_n1488# 0.05837f
C80 source.t14 a_n1846_n1488# 0.05837f
C81 source.n13 a_n1846_n1488# 0.370098f
C82 source.n14 a_n1846_n1488# 0.369058f
C83 source.t10 a_n1846_n1488# 0.484694f
C84 source.n15 a_n1846_n1488# 0.539582f
C85 source.n16 a_n1846_n1488# 0.729274f
C86 drain_right.t2 a_n1846_n1488# 0.043541f
C87 drain_right.t4 a_n1846_n1488# 0.043541f
C88 drain_right.n0 a_n1846_n1488# 0.315299f
C89 drain_right.t7 a_n1846_n1488# 0.043541f
C90 drain_right.t1 a_n1846_n1488# 0.043541f
C91 drain_right.n1 a_n1846_n1488# 0.315299f
C92 drain_right.n2 a_n1846_n1488# 1.01539f
C93 drain_right.t3 a_n1846_n1488# 0.043541f
C94 drain_right.t0 a_n1846_n1488# 0.043541f
C95 drain_right.n3 a_n1846_n1488# 0.31727f
C96 drain_right.t6 a_n1846_n1488# 0.043541f
C97 drain_right.t5 a_n1846_n1488# 0.043541f
C98 drain_right.n4 a_n1846_n1488# 0.314016f
C99 drain_right.n5 a_n1846_n1488# 0.693474f
C100 minus.n0 a_n1846_n1488# 0.045459f
C101 minus.t4 a_n1846_n1488# 0.245175f
C102 minus.n1 a_n1846_n1488# 0.149752f
C103 minus.t2 a_n1846_n1488# 0.245175f
C104 minus.t6 a_n1846_n1488# 0.263551f
C105 minus.n2 a_n1846_n1488# 0.12725f
C106 minus.n3 a_n1846_n1488# 0.194981f
C107 minus.n4 a_n1846_n1488# 0.149197f
C108 minus.n5 a_n1846_n1488# 0.007731f
C109 minus.t7 a_n1846_n1488# 0.245175f
C110 minus.n6 a_n1846_n1488# 0.136425f
C111 minus.n7 a_n1846_n1488# 0.863331f
C112 minus.n8 a_n1846_n1488# 0.045459f
C113 minus.t3 a_n1846_n1488# 0.245175f
C114 minus.n9 a_n1846_n1488# 0.149752f
C115 minus.t0 a_n1846_n1488# 0.263551f
C116 minus.n10 a_n1846_n1488# 0.12725f
C117 minus.n11 a_n1846_n1488# 0.194981f
C118 minus.t1 a_n1846_n1488# 0.245175f
C119 minus.n12 a_n1846_n1488# 0.149197f
C120 minus.n13 a_n1846_n1488# 0.007731f
C121 minus.t5 a_n1846_n1488# 0.245175f
C122 minus.n14 a_n1846_n1488# 0.136425f
C123 minus.n15 a_n1846_n1488# 0.234839f
C124 minus.n16 a_n1846_n1488# 1.05972f
.ends

