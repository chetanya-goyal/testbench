* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t33 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X1 source.t5 minus.t0 drain_right.t19 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X2 drain_right.t18 minus.t1 source.t9 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t31 plus.t1 drain_left.t18 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 drain_right.t17 minus.t2 source.t10 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 drain_right.t16 minus.t3 source.t14 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X6 source.t26 plus.t2 drain_left.t17 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X7 source.t34 plus.t3 drain_left.t16 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X8 drain_right.t15 minus.t4 source.t1 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X9 source.t32 plus.t4 drain_left.t15 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X10 drain_left.t14 plus.t5 source.t22 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X11 drain_left.t13 plus.t6 source.t24 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 source.t2 minus.t5 drain_right.t14 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X13 source.t39 minus.t6 drain_right.t13 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X14 drain_left.t12 plus.t7 source.t18 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X15 source.t4 minus.t7 drain_right.t12 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X16 drain_left.t11 plus.t8 source.t29 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X17 source.t21 plus.t9 drain_left.t10 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X18 source.t0 minus.t8 drain_right.t11 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X19 drain_right.t10 minus.t9 source.t3 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X20 source.t23 plus.t10 drain_left.t9 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X21 source.t13 minus.t10 drain_right.t9 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X22 drain_right.t8 minus.t11 source.t11 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X23 drain_left.t8 plus.t11 source.t30 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X24 drain_right.t7 minus.t12 source.t15 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X25 drain_right.t6 minus.t13 source.t38 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X26 a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X27 source.t35 plus.t12 drain_left.t7 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X28 a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X29 source.t12 minus.t14 drain_right.t5 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X30 source.t36 plus.t13 drain_left.t6 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X31 drain_left.t5 plus.t14 source.t20 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X32 drain_right.t4 minus.t15 source.t6 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X33 source.t27 plus.t15 drain_left.t4 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X34 source.t7 minus.t16 drain_right.t3 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X35 source.t17 minus.t17 drain_right.t2 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X36 a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X37 source.t16 minus.t18 drain_right.t1 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X38 drain_left.t3 plus.t16 source.t19 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X39 drain_left.t2 plus.t17 source.t28 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X40 source.t37 plus.t18 drain_left.t1 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X41 a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X42 drain_right.t0 minus.t19 source.t8 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X43 drain_left.t0 plus.t19 source.t25 a_n1882_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 plus.n5 plus.t9 453.884
R1 plus.n23 plus.t7 453.884
R2 plus.n30 plus.t16 453.884
R3 plus.n48 plus.t3 453.884
R4 plus.n6 plus.t5 397.651
R5 plus.n8 plus.t18 397.651
R6 plus.n3 plus.t14 397.651
R7 plus.n13 plus.t13 397.651
R8 plus.n15 plus.t8 397.651
R9 plus.n1 plus.t4 397.651
R10 plus.n20 plus.t17 397.651
R11 plus.n22 plus.t12 397.651
R12 plus.n31 plus.t2 397.651
R13 plus.n33 plus.t11 397.651
R14 plus.n28 plus.t1 397.651
R15 plus.n38 plus.t6 397.651
R16 plus.n40 plus.t15 397.651
R17 plus.n26 plus.t0 397.651
R18 plus.n45 plus.t10 397.651
R19 plus.n47 plus.t19 397.651
R20 plus.n5 plus.n4 161.489
R21 plus.n30 plus.n29 161.489
R22 plus.n7 plus.n4 161.3
R23 plus.n10 plus.n9 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n2 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n0 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n32 plus.n29 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n36 161.3
R33 plus.n39 plus.n27 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n25 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n7 plus.n6 51.852
R39 plus.n22 plus.n21 51.852
R40 plus.n47 plus.n46 51.852
R41 plus.n32 plus.n31 51.852
R42 plus.n9 plus.n8 47.4702
R43 plus.n20 plus.n19 47.4702
R44 plus.n45 plus.n44 47.4702
R45 plus.n34 plus.n33 47.4702
R46 plus.n12 plus.n3 43.0884
R47 plus.n16 plus.n1 43.0884
R48 plus.n41 plus.n26 43.0884
R49 plus.n37 plus.n28 43.0884
R50 plus.n14 plus.n13 38.7066
R51 plus.n15 plus.n14 38.7066
R52 plus.n40 plus.n39 38.7066
R53 plus.n39 plus.n38 38.7066
R54 plus.n13 plus.n12 34.3247
R55 plus.n16 plus.n15 34.3247
R56 plus.n41 plus.n40 34.3247
R57 plus.n38 plus.n37 34.3247
R58 plus.n9 plus.n3 29.9429
R59 plus.n19 plus.n1 29.9429
R60 plus.n44 plus.n26 29.9429
R61 plus.n34 plus.n28 29.9429
R62 plus plus.n49 26.321
R63 plus.n8 plus.n7 25.5611
R64 plus.n21 plus.n20 25.5611
R65 plus.n46 plus.n45 25.5611
R66 plus.n33 plus.n32 25.5611
R67 plus.n6 plus.n5 21.1793
R68 plus.n23 plus.n22 21.1793
R69 plus.n48 plus.n47 21.1793
R70 plus.n31 plus.n30 21.1793
R71 plus plus.n24 8.33383
R72 plus.n10 plus.n4 0.189894
R73 plus.n11 plus.n10 0.189894
R74 plus.n11 plus.n2 0.189894
R75 plus.n17 plus.n2 0.189894
R76 plus.n18 plus.n17 0.189894
R77 plus.n18 plus.n0 0.189894
R78 plus.n24 plus.n0 0.189894
R79 plus.n49 plus.n25 0.189894
R80 plus.n43 plus.n25 0.189894
R81 plus.n43 plus.n42 0.189894
R82 plus.n42 plus.n27 0.189894
R83 plus.n36 plus.n27 0.189894
R84 plus.n36 plus.n35 0.189894
R85 plus.n35 plus.n29 0.189894
R86 source.n90 source.n88 289.615
R87 source.n74 source.n72 289.615
R88 source.n66 source.n64 289.615
R89 source.n50 source.n48 289.615
R90 source.n2 source.n0 289.615
R91 source.n18 source.n16 289.615
R92 source.n26 source.n24 289.615
R93 source.n42 source.n40 289.615
R94 source.n91 source.n90 185
R95 source.n75 source.n74 185
R96 source.n67 source.n66 185
R97 source.n51 source.n50 185
R98 source.n3 source.n2 185
R99 source.n19 source.n18 185
R100 source.n27 source.n26 185
R101 source.n43 source.n42 185
R102 source.t8 source.n89 167.117
R103 source.t16 source.n73 167.117
R104 source.t19 source.n65 167.117
R105 source.t34 source.n49 167.117
R106 source.t18 source.n1 167.117
R107 source.t21 source.n17 167.117
R108 source.t15 source.n25 167.117
R109 source.t4 source.n41 167.117
R110 source.n9 source.n8 84.1169
R111 source.n11 source.n10 84.1169
R112 source.n13 source.n12 84.1169
R113 source.n15 source.n14 84.1169
R114 source.n33 source.n32 84.1169
R115 source.n35 source.n34 84.1169
R116 source.n37 source.n36 84.1169
R117 source.n39 source.n38 84.1169
R118 source.n87 source.n86 84.1168
R119 source.n85 source.n84 84.1168
R120 source.n83 source.n82 84.1168
R121 source.n81 source.n80 84.1168
R122 source.n63 source.n62 84.1168
R123 source.n61 source.n60 84.1168
R124 source.n59 source.n58 84.1168
R125 source.n57 source.n56 84.1168
R126 source.n90 source.t8 52.3082
R127 source.n74 source.t16 52.3082
R128 source.n66 source.t19 52.3082
R129 source.n50 source.t34 52.3082
R130 source.n2 source.t18 52.3082
R131 source.n18 source.t21 52.3082
R132 source.n26 source.t15 52.3082
R133 source.n42 source.t4 52.3082
R134 source.n95 source.n94 31.4096
R135 source.n79 source.n78 31.4096
R136 source.n71 source.n70 31.4096
R137 source.n55 source.n54 31.4096
R138 source.n7 source.n6 31.4096
R139 source.n23 source.n22 31.4096
R140 source.n31 source.n30 31.4096
R141 source.n47 source.n46 31.4096
R142 source.n55 source.n47 14.1689
R143 source.n86 source.t1 9.9005
R144 source.n86 source.t0 9.9005
R145 source.n84 source.t3 9.9005
R146 source.n84 source.t12 9.9005
R147 source.n82 source.t6 9.9005
R148 source.n82 source.t5 9.9005
R149 source.n80 source.t9 9.9005
R150 source.n80 source.t13 9.9005
R151 source.n62 source.t30 9.9005
R152 source.n62 source.t26 9.9005
R153 source.n60 source.t24 9.9005
R154 source.n60 source.t31 9.9005
R155 source.n58 source.t33 9.9005
R156 source.n58 source.t27 9.9005
R157 source.n56 source.t25 9.9005
R158 source.n56 source.t23 9.9005
R159 source.n8 source.t28 9.9005
R160 source.n8 source.t35 9.9005
R161 source.n10 source.t29 9.9005
R162 source.n10 source.t32 9.9005
R163 source.n12 source.t20 9.9005
R164 source.n12 source.t36 9.9005
R165 source.n14 source.t22 9.9005
R166 source.n14 source.t37 9.9005
R167 source.n32 source.t10 9.9005
R168 source.n32 source.t39 9.9005
R169 source.n34 source.t38 9.9005
R170 source.n34 source.t7 9.9005
R171 source.n36 source.t14 9.9005
R172 source.n36 source.t2 9.9005
R173 source.n38 source.t11 9.9005
R174 source.n38 source.t17 9.9005
R175 source.n91 source.n89 9.71174
R176 source.n75 source.n73 9.71174
R177 source.n67 source.n65 9.71174
R178 source.n51 source.n49 9.71174
R179 source.n3 source.n1 9.71174
R180 source.n19 source.n17 9.71174
R181 source.n27 source.n25 9.71174
R182 source.n43 source.n41 9.71174
R183 source.n94 source.n93 9.45567
R184 source.n78 source.n77 9.45567
R185 source.n70 source.n69 9.45567
R186 source.n54 source.n53 9.45567
R187 source.n6 source.n5 9.45567
R188 source.n22 source.n21 9.45567
R189 source.n30 source.n29 9.45567
R190 source.n46 source.n45 9.45567
R191 source.n93 source.n92 9.3005
R192 source.n77 source.n76 9.3005
R193 source.n69 source.n68 9.3005
R194 source.n53 source.n52 9.3005
R195 source.n5 source.n4 9.3005
R196 source.n21 source.n20 9.3005
R197 source.n29 source.n28 9.3005
R198 source.n45 source.n44 9.3005
R199 source.n96 source.n7 8.67749
R200 source.n94 source.n88 8.14595
R201 source.n78 source.n72 8.14595
R202 source.n70 source.n64 8.14595
R203 source.n54 source.n48 8.14595
R204 source.n6 source.n0 8.14595
R205 source.n22 source.n16 8.14595
R206 source.n30 source.n24 8.14595
R207 source.n46 source.n40 8.14595
R208 source.n92 source.n91 7.3702
R209 source.n76 source.n75 7.3702
R210 source.n68 source.n67 7.3702
R211 source.n52 source.n51 7.3702
R212 source.n4 source.n3 7.3702
R213 source.n20 source.n19 7.3702
R214 source.n28 source.n27 7.3702
R215 source.n44 source.n43 7.3702
R216 source.n92 source.n88 5.81868
R217 source.n76 source.n72 5.81868
R218 source.n68 source.n64 5.81868
R219 source.n52 source.n48 5.81868
R220 source.n4 source.n0 5.81868
R221 source.n20 source.n16 5.81868
R222 source.n28 source.n24 5.81868
R223 source.n44 source.n40 5.81868
R224 source.n96 source.n95 5.49188
R225 source.n93 source.n89 3.44771
R226 source.n77 source.n73 3.44771
R227 source.n69 source.n65 3.44771
R228 source.n53 source.n49 3.44771
R229 source.n5 source.n1 3.44771
R230 source.n21 source.n17 3.44771
R231 source.n29 source.n25 3.44771
R232 source.n45 source.n41 3.44771
R233 source.n31 source.n23 0.470328
R234 source.n79 source.n71 0.470328
R235 source.n47 source.n39 0.457397
R236 source.n39 source.n37 0.457397
R237 source.n37 source.n35 0.457397
R238 source.n35 source.n33 0.457397
R239 source.n33 source.n31 0.457397
R240 source.n23 source.n15 0.457397
R241 source.n15 source.n13 0.457397
R242 source.n13 source.n11 0.457397
R243 source.n11 source.n9 0.457397
R244 source.n9 source.n7 0.457397
R245 source.n57 source.n55 0.457397
R246 source.n59 source.n57 0.457397
R247 source.n61 source.n59 0.457397
R248 source.n63 source.n61 0.457397
R249 source.n71 source.n63 0.457397
R250 source.n81 source.n79 0.457397
R251 source.n83 source.n81 0.457397
R252 source.n85 source.n83 0.457397
R253 source.n87 source.n85 0.457397
R254 source.n95 source.n87 0.457397
R255 source source.n96 0.188
R256 drain_left.n10 drain_left.n8 101.252
R257 drain_left.n6 drain_left.n4 101.252
R258 drain_left.n2 drain_left.n0 101.252
R259 drain_left.n16 drain_left.n15 100.796
R260 drain_left.n14 drain_left.n13 100.796
R261 drain_left.n12 drain_left.n11 100.796
R262 drain_left.n10 drain_left.n9 100.796
R263 drain_left.n7 drain_left.n3 100.796
R264 drain_left.n6 drain_left.n5 100.796
R265 drain_left.n2 drain_left.n1 100.796
R266 drain_left drain_left.n7 23.4465
R267 drain_left.n3 drain_left.t4 9.9005
R268 drain_left.n3 drain_left.t13 9.9005
R269 drain_left.n4 drain_left.t17 9.9005
R270 drain_left.n4 drain_left.t3 9.9005
R271 drain_left.n5 drain_left.t18 9.9005
R272 drain_left.n5 drain_left.t8 9.9005
R273 drain_left.n1 drain_left.t9 9.9005
R274 drain_left.n1 drain_left.t19 9.9005
R275 drain_left.n0 drain_left.t16 9.9005
R276 drain_left.n0 drain_left.t0 9.9005
R277 drain_left.n15 drain_left.t7 9.9005
R278 drain_left.n15 drain_left.t12 9.9005
R279 drain_left.n13 drain_left.t15 9.9005
R280 drain_left.n13 drain_left.t2 9.9005
R281 drain_left.n11 drain_left.t6 9.9005
R282 drain_left.n11 drain_left.t11 9.9005
R283 drain_left.n9 drain_left.t1 9.9005
R284 drain_left.n9 drain_left.t5 9.9005
R285 drain_left.n8 drain_left.t10 9.9005
R286 drain_left.n8 drain_left.t14 9.9005
R287 drain_left drain_left.n16 6.11011
R288 drain_left.n12 drain_left.n10 0.457397
R289 drain_left.n14 drain_left.n12 0.457397
R290 drain_left.n16 drain_left.n14 0.457397
R291 drain_left.n7 drain_left.n6 0.402051
R292 drain_left.n7 drain_left.n2 0.402051
R293 minus.n23 minus.t7 453.884
R294 minus.n5 minus.t12 453.884
R295 minus.n48 minus.t19 453.884
R296 minus.n30 minus.t18 453.884
R297 minus.n22 minus.t11 397.651
R298 minus.n20 minus.t17 397.651
R299 minus.n1 minus.t3 397.651
R300 minus.n15 minus.t5 397.651
R301 minus.n13 minus.t13 397.651
R302 minus.n3 minus.t16 397.651
R303 minus.n8 minus.t2 397.651
R304 minus.n6 minus.t6 397.651
R305 minus.n47 minus.t8 397.651
R306 minus.n45 minus.t4 397.651
R307 minus.n26 minus.t14 397.651
R308 minus.n40 minus.t9 397.651
R309 minus.n38 minus.t0 397.651
R310 minus.n28 minus.t15 397.651
R311 minus.n33 minus.t10 397.651
R312 minus.n31 minus.t1 397.651
R313 minus.n5 minus.n4 161.489
R314 minus.n30 minus.n29 161.489
R315 minus.n24 minus.n23 161.3
R316 minus.n21 minus.n0 161.3
R317 minus.n19 minus.n18 161.3
R318 minus.n17 minus.n16 161.3
R319 minus.n14 minus.n2 161.3
R320 minus.n12 minus.n11 161.3
R321 minus.n10 minus.n9 161.3
R322 minus.n7 minus.n4 161.3
R323 minus.n49 minus.n48 161.3
R324 minus.n46 minus.n25 161.3
R325 minus.n44 minus.n43 161.3
R326 minus.n42 minus.n41 161.3
R327 minus.n39 minus.n27 161.3
R328 minus.n37 minus.n36 161.3
R329 minus.n35 minus.n34 161.3
R330 minus.n32 minus.n29 161.3
R331 minus.n22 minus.n21 51.852
R332 minus.n7 minus.n6 51.852
R333 minus.n32 minus.n31 51.852
R334 minus.n47 minus.n46 51.852
R335 minus.n20 minus.n19 47.4702
R336 minus.n9 minus.n8 47.4702
R337 minus.n34 minus.n33 47.4702
R338 minus.n45 minus.n44 47.4702
R339 minus.n16 minus.n1 43.0884
R340 minus.n12 minus.n3 43.0884
R341 minus.n37 minus.n28 43.0884
R342 minus.n41 minus.n26 43.0884
R343 minus.n15 minus.n14 38.7066
R344 minus.n14 minus.n13 38.7066
R345 minus.n39 minus.n38 38.7066
R346 minus.n40 minus.n39 38.7066
R347 minus.n16 minus.n15 34.3247
R348 minus.n13 minus.n12 34.3247
R349 minus.n38 minus.n37 34.3247
R350 minus.n41 minus.n40 34.3247
R351 minus.n19 minus.n1 29.9429
R352 minus.n9 minus.n3 29.9429
R353 minus.n34 minus.n28 29.9429
R354 minus.n44 minus.n26 29.9429
R355 minus.n50 minus.n24 28.652
R356 minus.n21 minus.n20 25.5611
R357 minus.n8 minus.n7 25.5611
R358 minus.n33 minus.n32 25.5611
R359 minus.n46 minus.n45 25.5611
R360 minus.n23 minus.n22 21.1793
R361 minus.n6 minus.n5 21.1793
R362 minus.n31 minus.n30 21.1793
R363 minus.n48 minus.n47 21.1793
R364 minus.n50 minus.n49 6.47777
R365 minus.n24 minus.n0 0.189894
R366 minus.n18 minus.n0 0.189894
R367 minus.n18 minus.n17 0.189894
R368 minus.n17 minus.n2 0.189894
R369 minus.n11 minus.n2 0.189894
R370 minus.n11 minus.n10 0.189894
R371 minus.n10 minus.n4 0.189894
R372 minus.n35 minus.n29 0.189894
R373 minus.n36 minus.n35 0.189894
R374 minus.n36 minus.n27 0.189894
R375 minus.n42 minus.n27 0.189894
R376 minus.n43 minus.n42 0.189894
R377 minus.n43 minus.n25 0.189894
R378 minus.n49 minus.n25 0.189894
R379 minus minus.n50 0.188
R380 drain_right.n10 drain_right.n8 101.252
R381 drain_right.n6 drain_right.n4 101.252
R382 drain_right.n2 drain_right.n0 101.252
R383 drain_right.n10 drain_right.n9 100.796
R384 drain_right.n12 drain_right.n11 100.796
R385 drain_right.n14 drain_right.n13 100.796
R386 drain_right.n16 drain_right.n15 100.796
R387 drain_right.n7 drain_right.n3 100.796
R388 drain_right.n6 drain_right.n5 100.796
R389 drain_right.n2 drain_right.n1 100.796
R390 drain_right drain_right.n7 22.8933
R391 drain_right.n3 drain_right.t19 9.9005
R392 drain_right.n3 drain_right.t10 9.9005
R393 drain_right.n4 drain_right.t11 9.9005
R394 drain_right.n4 drain_right.t0 9.9005
R395 drain_right.n5 drain_right.t5 9.9005
R396 drain_right.n5 drain_right.t15 9.9005
R397 drain_right.n1 drain_right.t9 9.9005
R398 drain_right.n1 drain_right.t4 9.9005
R399 drain_right.n0 drain_right.t1 9.9005
R400 drain_right.n0 drain_right.t18 9.9005
R401 drain_right.n8 drain_right.t13 9.9005
R402 drain_right.n8 drain_right.t7 9.9005
R403 drain_right.n9 drain_right.t3 9.9005
R404 drain_right.n9 drain_right.t17 9.9005
R405 drain_right.n11 drain_right.t14 9.9005
R406 drain_right.n11 drain_right.t6 9.9005
R407 drain_right.n13 drain_right.t2 9.9005
R408 drain_right.n13 drain_right.t16 9.9005
R409 drain_right.n15 drain_right.t12 9.9005
R410 drain_right.n15 drain_right.t8 9.9005
R411 drain_right drain_right.n16 6.11011
R412 drain_right.n16 drain_right.n14 0.457397
R413 drain_right.n14 drain_right.n12 0.457397
R414 drain_right.n12 drain_right.n10 0.457397
R415 drain_right.n7 drain_right.n6 0.402051
R416 drain_right.n7 drain_right.n2 0.402051
C0 drain_right plus 0.343902f
C1 source drain_left 10.1826f
C2 plus drain_left 1.54919f
C3 plus source 1.54652f
C4 drain_right minus 1.36613f
C5 minus drain_left 0.177242f
C6 drain_right drain_left 0.982283f
C7 minus source 1.53256f
C8 drain_right source 10.1826f
C9 minus plus 3.65786f
C10 drain_right a_n1882_n1288# 4.28179f
C11 drain_left a_n1882_n1288# 4.54898f
C12 source a_n1882_n1288# 3.145518f
C13 minus a_n1882_n1288# 6.506308f
C14 plus a_n1882_n1288# 7.171153f
C15 drain_right.t1 a_n1882_n1288# 0.049517f
C16 drain_right.t18 a_n1882_n1288# 0.049517f
C17 drain_right.n0 a_n1882_n1288# 0.312636f
C18 drain_right.t9 a_n1882_n1288# 0.049517f
C19 drain_right.t4 a_n1882_n1288# 0.049517f
C20 drain_right.n1 a_n1882_n1288# 0.311081f
C21 drain_right.n2 a_n1882_n1288# 0.671393f
C22 drain_right.t19 a_n1882_n1288# 0.049517f
C23 drain_right.t10 a_n1882_n1288# 0.049517f
C24 drain_right.n3 a_n1882_n1288# 0.311081f
C25 drain_right.t11 a_n1882_n1288# 0.049517f
C26 drain_right.t0 a_n1882_n1288# 0.049517f
C27 drain_right.n4 a_n1882_n1288# 0.312636f
C28 drain_right.t5 a_n1882_n1288# 0.049517f
C29 drain_right.t15 a_n1882_n1288# 0.049517f
C30 drain_right.n5 a_n1882_n1288# 0.311081f
C31 drain_right.n6 a_n1882_n1288# 0.671393f
C32 drain_right.n7 a_n1882_n1288# 1.12604f
C33 drain_right.t13 a_n1882_n1288# 0.049517f
C34 drain_right.t7 a_n1882_n1288# 0.049517f
C35 drain_right.n8 a_n1882_n1288# 0.312637f
C36 drain_right.t3 a_n1882_n1288# 0.049517f
C37 drain_right.t17 a_n1882_n1288# 0.049517f
C38 drain_right.n9 a_n1882_n1288# 0.311082f
C39 drain_right.n10 a_n1882_n1288# 0.675169f
C40 drain_right.t14 a_n1882_n1288# 0.049517f
C41 drain_right.t6 a_n1882_n1288# 0.049517f
C42 drain_right.n11 a_n1882_n1288# 0.311082f
C43 drain_right.n12 a_n1882_n1288# 0.332053f
C44 drain_right.t2 a_n1882_n1288# 0.049517f
C45 drain_right.t16 a_n1882_n1288# 0.049517f
C46 drain_right.n13 a_n1882_n1288# 0.311082f
C47 drain_right.n14 a_n1882_n1288# 0.332053f
C48 drain_right.t12 a_n1882_n1288# 0.049517f
C49 drain_right.t8 a_n1882_n1288# 0.049517f
C50 drain_right.n15 a_n1882_n1288# 0.311082f
C51 drain_right.n16 a_n1882_n1288# 0.588464f
C52 minus.n0 a_n1882_n1288# 0.029372f
C53 minus.t7 a_n1882_n1288# 0.038128f
C54 minus.t11 a_n1882_n1288# 0.034571f
C55 minus.t17 a_n1882_n1288# 0.034571f
C56 minus.t3 a_n1882_n1288# 0.034571f
C57 minus.n1 a_n1882_n1288# 0.027163f
C58 minus.n2 a_n1882_n1288# 0.029372f
C59 minus.t5 a_n1882_n1288# 0.034571f
C60 minus.t13 a_n1882_n1288# 0.034571f
C61 minus.t16 a_n1882_n1288# 0.034571f
C62 minus.n3 a_n1882_n1288# 0.027163f
C63 minus.n4 a_n1882_n1288# 0.06721f
C64 minus.t2 a_n1882_n1288# 0.034571f
C65 minus.t6 a_n1882_n1288# 0.034571f
C66 minus.t12 a_n1882_n1288# 0.038128f
C67 minus.n5 a_n1882_n1288# 0.035478f
C68 minus.n6 a_n1882_n1288# 0.027163f
C69 minus.n7 a_n1882_n1288# 0.010287f
C70 minus.n8 a_n1882_n1288# 0.027163f
C71 minus.n9 a_n1882_n1288# 0.010287f
C72 minus.n10 a_n1882_n1288# 0.029372f
C73 minus.n11 a_n1882_n1288# 0.029372f
C74 minus.n12 a_n1882_n1288# 0.010287f
C75 minus.n13 a_n1882_n1288# 0.027163f
C76 minus.n14 a_n1882_n1288# 0.010287f
C77 minus.n15 a_n1882_n1288# 0.027163f
C78 minus.n16 a_n1882_n1288# 0.010287f
C79 minus.n17 a_n1882_n1288# 0.029372f
C80 minus.n18 a_n1882_n1288# 0.029372f
C81 minus.n19 a_n1882_n1288# 0.010287f
C82 minus.n20 a_n1882_n1288# 0.027163f
C83 minus.n21 a_n1882_n1288# 0.010287f
C84 minus.n22 a_n1882_n1288# 0.027163f
C85 minus.n23 a_n1882_n1288# 0.035433f
C86 minus.n24 a_n1882_n1288# 0.705095f
C87 minus.n25 a_n1882_n1288# 0.029372f
C88 minus.t8 a_n1882_n1288# 0.034571f
C89 minus.t4 a_n1882_n1288# 0.034571f
C90 minus.t14 a_n1882_n1288# 0.034571f
C91 minus.n26 a_n1882_n1288# 0.027163f
C92 minus.n27 a_n1882_n1288# 0.029372f
C93 minus.t9 a_n1882_n1288# 0.034571f
C94 minus.t0 a_n1882_n1288# 0.034571f
C95 minus.t15 a_n1882_n1288# 0.034571f
C96 minus.n28 a_n1882_n1288# 0.027163f
C97 minus.n29 a_n1882_n1288# 0.06721f
C98 minus.t10 a_n1882_n1288# 0.034571f
C99 minus.t1 a_n1882_n1288# 0.034571f
C100 minus.t18 a_n1882_n1288# 0.038128f
C101 minus.n30 a_n1882_n1288# 0.035478f
C102 minus.n31 a_n1882_n1288# 0.027163f
C103 minus.n32 a_n1882_n1288# 0.010287f
C104 minus.n33 a_n1882_n1288# 0.027163f
C105 minus.n34 a_n1882_n1288# 0.010287f
C106 minus.n35 a_n1882_n1288# 0.029372f
C107 minus.n36 a_n1882_n1288# 0.029372f
C108 minus.n37 a_n1882_n1288# 0.010287f
C109 minus.n38 a_n1882_n1288# 0.027163f
C110 minus.n39 a_n1882_n1288# 0.010287f
C111 minus.n40 a_n1882_n1288# 0.027163f
C112 minus.n41 a_n1882_n1288# 0.010287f
C113 minus.n42 a_n1882_n1288# 0.029372f
C114 minus.n43 a_n1882_n1288# 0.029372f
C115 minus.n44 a_n1882_n1288# 0.010287f
C116 minus.n45 a_n1882_n1288# 0.027163f
C117 minus.n46 a_n1882_n1288# 0.010287f
C118 minus.n47 a_n1882_n1288# 0.027163f
C119 minus.t19 a_n1882_n1288# 0.038128f
C120 minus.n48 a_n1882_n1288# 0.035433f
C121 minus.n49 a_n1882_n1288# 0.190485f
C122 minus.n50 a_n1882_n1288# 0.872146f
C123 drain_left.t16 a_n1882_n1288# 0.048929f
C124 drain_left.t0 a_n1882_n1288# 0.048929f
C125 drain_left.n0 a_n1882_n1288# 0.308924f
C126 drain_left.t9 a_n1882_n1288# 0.048929f
C127 drain_left.t19 a_n1882_n1288# 0.048929f
C128 drain_left.n1 a_n1882_n1288# 0.307387f
C129 drain_left.n2 a_n1882_n1288# 0.663422f
C130 drain_left.t4 a_n1882_n1288# 0.048929f
C131 drain_left.t13 a_n1882_n1288# 0.048929f
C132 drain_left.n3 a_n1882_n1288# 0.307387f
C133 drain_left.t17 a_n1882_n1288# 0.048929f
C134 drain_left.t3 a_n1882_n1288# 0.048929f
C135 drain_left.n4 a_n1882_n1288# 0.308924f
C136 drain_left.t18 a_n1882_n1288# 0.048929f
C137 drain_left.t8 a_n1882_n1288# 0.048929f
C138 drain_left.n5 a_n1882_n1288# 0.307387f
C139 drain_left.n6 a_n1882_n1288# 0.663422f
C140 drain_left.n7 a_n1882_n1288# 1.17329f
C141 drain_left.t10 a_n1882_n1288# 0.048929f
C142 drain_left.t14 a_n1882_n1288# 0.048929f
C143 drain_left.n8 a_n1882_n1288# 0.308925f
C144 drain_left.t1 a_n1882_n1288# 0.048929f
C145 drain_left.t5 a_n1882_n1288# 0.048929f
C146 drain_left.n9 a_n1882_n1288# 0.307388f
C147 drain_left.n10 a_n1882_n1288# 0.667153f
C148 drain_left.t6 a_n1882_n1288# 0.048929f
C149 drain_left.t11 a_n1882_n1288# 0.048929f
C150 drain_left.n11 a_n1882_n1288# 0.307388f
C151 drain_left.n12 a_n1882_n1288# 0.32811f
C152 drain_left.t15 a_n1882_n1288# 0.048929f
C153 drain_left.t2 a_n1882_n1288# 0.048929f
C154 drain_left.n13 a_n1882_n1288# 0.307388f
C155 drain_left.n14 a_n1882_n1288# 0.32811f
C156 drain_left.t7 a_n1882_n1288# 0.048929f
C157 drain_left.t12 a_n1882_n1288# 0.048929f
C158 drain_left.n15 a_n1882_n1288# 0.307388f
C159 drain_left.n16 a_n1882_n1288# 0.581477f
C160 source.n0 a_n1882_n1288# 0.047409f
C161 source.n1 a_n1882_n1288# 0.104898f
C162 source.t18 a_n1882_n1288# 0.078721f
C163 source.n2 a_n1882_n1288# 0.082098f
C164 source.n3 a_n1882_n1288# 0.026465f
C165 source.n4 a_n1882_n1288# 0.017454f
C166 source.n5 a_n1882_n1288# 0.231222f
C167 source.n6 a_n1882_n1288# 0.051971f
C168 source.n7 a_n1882_n1288# 0.474375f
C169 source.t28 a_n1882_n1288# 0.051336f
C170 source.t35 a_n1882_n1288# 0.051336f
C171 source.n8 a_n1882_n1288# 0.274441f
C172 source.n9 a_n1882_n1288# 0.348171f
C173 source.t29 a_n1882_n1288# 0.051336f
C174 source.t32 a_n1882_n1288# 0.051336f
C175 source.n10 a_n1882_n1288# 0.274441f
C176 source.n11 a_n1882_n1288# 0.348171f
C177 source.t20 a_n1882_n1288# 0.051336f
C178 source.t36 a_n1882_n1288# 0.051336f
C179 source.n12 a_n1882_n1288# 0.274441f
C180 source.n13 a_n1882_n1288# 0.348171f
C181 source.t22 a_n1882_n1288# 0.051336f
C182 source.t37 a_n1882_n1288# 0.051336f
C183 source.n14 a_n1882_n1288# 0.274441f
C184 source.n15 a_n1882_n1288# 0.348171f
C185 source.n16 a_n1882_n1288# 0.047409f
C186 source.n17 a_n1882_n1288# 0.104898f
C187 source.t21 a_n1882_n1288# 0.078721f
C188 source.n18 a_n1882_n1288# 0.082098f
C189 source.n19 a_n1882_n1288# 0.026465f
C190 source.n20 a_n1882_n1288# 0.017454f
C191 source.n21 a_n1882_n1288# 0.231222f
C192 source.n22 a_n1882_n1288# 0.051971f
C193 source.n23 a_n1882_n1288# 0.123734f
C194 source.n24 a_n1882_n1288# 0.047409f
C195 source.n25 a_n1882_n1288# 0.104898f
C196 source.t15 a_n1882_n1288# 0.078721f
C197 source.n26 a_n1882_n1288# 0.082098f
C198 source.n27 a_n1882_n1288# 0.026465f
C199 source.n28 a_n1882_n1288# 0.017454f
C200 source.n29 a_n1882_n1288# 0.231222f
C201 source.n30 a_n1882_n1288# 0.051971f
C202 source.n31 a_n1882_n1288# 0.123734f
C203 source.t10 a_n1882_n1288# 0.051336f
C204 source.t39 a_n1882_n1288# 0.051336f
C205 source.n32 a_n1882_n1288# 0.274441f
C206 source.n33 a_n1882_n1288# 0.348171f
C207 source.t38 a_n1882_n1288# 0.051336f
C208 source.t7 a_n1882_n1288# 0.051336f
C209 source.n34 a_n1882_n1288# 0.274441f
C210 source.n35 a_n1882_n1288# 0.348171f
C211 source.t14 a_n1882_n1288# 0.051336f
C212 source.t2 a_n1882_n1288# 0.051336f
C213 source.n36 a_n1882_n1288# 0.274441f
C214 source.n37 a_n1882_n1288# 0.348171f
C215 source.t11 a_n1882_n1288# 0.051336f
C216 source.t17 a_n1882_n1288# 0.051336f
C217 source.n38 a_n1882_n1288# 0.274441f
C218 source.n39 a_n1882_n1288# 0.348171f
C219 source.n40 a_n1882_n1288# 0.047409f
C220 source.n41 a_n1882_n1288# 0.104898f
C221 source.t4 a_n1882_n1288# 0.078721f
C222 source.n42 a_n1882_n1288# 0.082098f
C223 source.n43 a_n1882_n1288# 0.026465f
C224 source.n44 a_n1882_n1288# 0.017454f
C225 source.n45 a_n1882_n1288# 0.231222f
C226 source.n46 a_n1882_n1288# 0.051971f
C227 source.n47 a_n1882_n1288# 0.775204f
C228 source.n48 a_n1882_n1288# 0.047409f
C229 source.n49 a_n1882_n1288# 0.104898f
C230 source.t34 a_n1882_n1288# 0.078721f
C231 source.n50 a_n1882_n1288# 0.082098f
C232 source.n51 a_n1882_n1288# 0.026465f
C233 source.n52 a_n1882_n1288# 0.017454f
C234 source.n53 a_n1882_n1288# 0.231222f
C235 source.n54 a_n1882_n1288# 0.051971f
C236 source.n55 a_n1882_n1288# 0.775204f
C237 source.t25 a_n1882_n1288# 0.051336f
C238 source.t23 a_n1882_n1288# 0.051336f
C239 source.n56 a_n1882_n1288# 0.27444f
C240 source.n57 a_n1882_n1288# 0.348173f
C241 source.t33 a_n1882_n1288# 0.051336f
C242 source.t27 a_n1882_n1288# 0.051336f
C243 source.n58 a_n1882_n1288# 0.27444f
C244 source.n59 a_n1882_n1288# 0.348173f
C245 source.t24 a_n1882_n1288# 0.051336f
C246 source.t31 a_n1882_n1288# 0.051336f
C247 source.n60 a_n1882_n1288# 0.27444f
C248 source.n61 a_n1882_n1288# 0.348173f
C249 source.t30 a_n1882_n1288# 0.051336f
C250 source.t26 a_n1882_n1288# 0.051336f
C251 source.n62 a_n1882_n1288# 0.27444f
C252 source.n63 a_n1882_n1288# 0.348173f
C253 source.n64 a_n1882_n1288# 0.047409f
C254 source.n65 a_n1882_n1288# 0.104898f
C255 source.t19 a_n1882_n1288# 0.078721f
C256 source.n66 a_n1882_n1288# 0.082098f
C257 source.n67 a_n1882_n1288# 0.026465f
C258 source.n68 a_n1882_n1288# 0.017454f
C259 source.n69 a_n1882_n1288# 0.231222f
C260 source.n70 a_n1882_n1288# 0.051971f
C261 source.n71 a_n1882_n1288# 0.123734f
C262 source.n72 a_n1882_n1288# 0.047409f
C263 source.n73 a_n1882_n1288# 0.104898f
C264 source.t16 a_n1882_n1288# 0.078721f
C265 source.n74 a_n1882_n1288# 0.082098f
C266 source.n75 a_n1882_n1288# 0.026465f
C267 source.n76 a_n1882_n1288# 0.017454f
C268 source.n77 a_n1882_n1288# 0.231222f
C269 source.n78 a_n1882_n1288# 0.051971f
C270 source.n79 a_n1882_n1288# 0.123734f
C271 source.t9 a_n1882_n1288# 0.051336f
C272 source.t13 a_n1882_n1288# 0.051336f
C273 source.n80 a_n1882_n1288# 0.27444f
C274 source.n81 a_n1882_n1288# 0.348173f
C275 source.t6 a_n1882_n1288# 0.051336f
C276 source.t5 a_n1882_n1288# 0.051336f
C277 source.n82 a_n1882_n1288# 0.27444f
C278 source.n83 a_n1882_n1288# 0.348173f
C279 source.t3 a_n1882_n1288# 0.051336f
C280 source.t12 a_n1882_n1288# 0.051336f
C281 source.n84 a_n1882_n1288# 0.27444f
C282 source.n85 a_n1882_n1288# 0.348173f
C283 source.t1 a_n1882_n1288# 0.051336f
C284 source.t0 a_n1882_n1288# 0.051336f
C285 source.n86 a_n1882_n1288# 0.27444f
C286 source.n87 a_n1882_n1288# 0.348173f
C287 source.n88 a_n1882_n1288# 0.047409f
C288 source.n89 a_n1882_n1288# 0.104898f
C289 source.t8 a_n1882_n1288# 0.078721f
C290 source.n90 a_n1882_n1288# 0.082098f
C291 source.n91 a_n1882_n1288# 0.026465f
C292 source.n92 a_n1882_n1288# 0.017454f
C293 source.n93 a_n1882_n1288# 0.231222f
C294 source.n94 a_n1882_n1288# 0.051971f
C295 source.n95 a_n1882_n1288# 0.29986f
C296 source.n96 a_n1882_n1288# 0.799277f
C297 plus.n0 a_n1882_n1288# 0.029851f
C298 plus.t12 a_n1882_n1288# 0.035136f
C299 plus.t17 a_n1882_n1288# 0.035136f
C300 plus.t4 a_n1882_n1288# 0.035136f
C301 plus.n1 a_n1882_n1288# 0.027607f
C302 plus.n2 a_n1882_n1288# 0.029851f
C303 plus.t8 a_n1882_n1288# 0.035136f
C304 plus.t13 a_n1882_n1288# 0.035136f
C305 plus.t14 a_n1882_n1288# 0.035136f
C306 plus.n3 a_n1882_n1288# 0.027607f
C307 plus.n4 a_n1882_n1288# 0.068307f
C308 plus.t18 a_n1882_n1288# 0.035136f
C309 plus.t5 a_n1882_n1288# 0.035136f
C310 plus.t9 a_n1882_n1288# 0.03875f
C311 plus.n5 a_n1882_n1288# 0.036057f
C312 plus.n6 a_n1882_n1288# 0.027607f
C313 plus.n7 a_n1882_n1288# 0.010455f
C314 plus.n8 a_n1882_n1288# 0.027607f
C315 plus.n9 a_n1882_n1288# 0.010455f
C316 plus.n10 a_n1882_n1288# 0.029851f
C317 plus.n11 a_n1882_n1288# 0.029851f
C318 plus.n12 a_n1882_n1288# 0.010455f
C319 plus.n13 a_n1882_n1288# 0.027607f
C320 plus.n14 a_n1882_n1288# 0.010455f
C321 plus.n15 a_n1882_n1288# 0.027607f
C322 plus.n16 a_n1882_n1288# 0.010455f
C323 plus.n17 a_n1882_n1288# 0.029851f
C324 plus.n18 a_n1882_n1288# 0.029851f
C325 plus.n19 a_n1882_n1288# 0.010455f
C326 plus.n20 a_n1882_n1288# 0.027607f
C327 plus.n21 a_n1882_n1288# 0.010455f
C328 plus.n22 a_n1882_n1288# 0.027607f
C329 plus.t7 a_n1882_n1288# 0.03875f
C330 plus.n23 a_n1882_n1288# 0.036011f
C331 plus.n24 a_n1882_n1288# 0.211752f
C332 plus.n25 a_n1882_n1288# 0.029851f
C333 plus.t3 a_n1882_n1288# 0.03875f
C334 plus.t19 a_n1882_n1288# 0.035136f
C335 plus.t10 a_n1882_n1288# 0.035136f
C336 plus.t0 a_n1882_n1288# 0.035136f
C337 plus.n26 a_n1882_n1288# 0.027607f
C338 plus.n27 a_n1882_n1288# 0.029851f
C339 plus.t15 a_n1882_n1288# 0.035136f
C340 plus.t6 a_n1882_n1288# 0.035136f
C341 plus.t1 a_n1882_n1288# 0.035136f
C342 plus.n28 a_n1882_n1288# 0.027607f
C343 plus.n29 a_n1882_n1288# 0.068307f
C344 plus.t11 a_n1882_n1288# 0.035136f
C345 plus.t2 a_n1882_n1288# 0.035136f
C346 plus.t16 a_n1882_n1288# 0.03875f
C347 plus.n30 a_n1882_n1288# 0.036057f
C348 plus.n31 a_n1882_n1288# 0.027607f
C349 plus.n32 a_n1882_n1288# 0.010455f
C350 plus.n33 a_n1882_n1288# 0.027607f
C351 plus.n34 a_n1882_n1288# 0.010455f
C352 plus.n35 a_n1882_n1288# 0.029851f
C353 plus.n36 a_n1882_n1288# 0.029851f
C354 plus.n37 a_n1882_n1288# 0.010455f
C355 plus.n38 a_n1882_n1288# 0.027607f
C356 plus.n39 a_n1882_n1288# 0.010455f
C357 plus.n40 a_n1882_n1288# 0.027607f
C358 plus.n41 a_n1882_n1288# 0.010455f
C359 plus.n42 a_n1882_n1288# 0.029851f
C360 plus.n43 a_n1882_n1288# 0.029851f
C361 plus.n44 a_n1882_n1288# 0.010455f
C362 plus.n45 a_n1882_n1288# 0.027607f
C363 plus.n46 a_n1882_n1288# 0.010455f
C364 plus.n47 a_n1882_n1288# 0.027607f
C365 plus.n48 a_n1882_n1288# 0.036011f
C366 plus.n49 a_n1882_n1288# 0.683897f
.ends

