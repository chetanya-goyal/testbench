* NGSPICE file created from diffpair700.ext - technology: sky130A

.subckt diffpair700 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.7
X1 a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.7
X2 a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X3 drain_left.t1 plus.t0 source.t1 a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.7
X4 drain_left.t0 plus.t1 source.t0 a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.7
X5 drain_right.t0 minus.t1 source.t3 a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.7
X6 a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X7 a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# a_n1128_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
R0 minus.n0 minus.t0 1121.51
R1 minus.n0 minus.t1 1084.75
R2 minus minus.n0 0.188
R3 source.n554 source.n420 289.615
R4 source.n414 source.n280 289.615
R5 source.n134 source.n0 289.615
R6 source.n274 source.n140 289.615
R7 source.n464 source.n463 185
R8 source.n469 source.n468 185
R9 source.n471 source.n470 185
R10 source.n460 source.n459 185
R11 source.n477 source.n476 185
R12 source.n479 source.n478 185
R13 source.n456 source.n455 185
R14 source.n486 source.n485 185
R15 source.n487 source.n454 185
R16 source.n489 source.n488 185
R17 source.n452 source.n451 185
R18 source.n495 source.n494 185
R19 source.n497 source.n496 185
R20 source.n448 source.n447 185
R21 source.n503 source.n502 185
R22 source.n505 source.n504 185
R23 source.n444 source.n443 185
R24 source.n511 source.n510 185
R25 source.n513 source.n512 185
R26 source.n440 source.n439 185
R27 source.n519 source.n518 185
R28 source.n521 source.n520 185
R29 source.n436 source.n435 185
R30 source.n527 source.n526 185
R31 source.n530 source.n529 185
R32 source.n528 source.n432 185
R33 source.n535 source.n431 185
R34 source.n537 source.n536 185
R35 source.n539 source.n538 185
R36 source.n428 source.n427 185
R37 source.n545 source.n544 185
R38 source.n547 source.n546 185
R39 source.n424 source.n423 185
R40 source.n553 source.n552 185
R41 source.n555 source.n554 185
R42 source.n324 source.n323 185
R43 source.n329 source.n328 185
R44 source.n331 source.n330 185
R45 source.n320 source.n319 185
R46 source.n337 source.n336 185
R47 source.n339 source.n338 185
R48 source.n316 source.n315 185
R49 source.n346 source.n345 185
R50 source.n347 source.n314 185
R51 source.n349 source.n348 185
R52 source.n312 source.n311 185
R53 source.n355 source.n354 185
R54 source.n357 source.n356 185
R55 source.n308 source.n307 185
R56 source.n363 source.n362 185
R57 source.n365 source.n364 185
R58 source.n304 source.n303 185
R59 source.n371 source.n370 185
R60 source.n373 source.n372 185
R61 source.n300 source.n299 185
R62 source.n379 source.n378 185
R63 source.n381 source.n380 185
R64 source.n296 source.n295 185
R65 source.n387 source.n386 185
R66 source.n390 source.n389 185
R67 source.n388 source.n292 185
R68 source.n395 source.n291 185
R69 source.n397 source.n396 185
R70 source.n399 source.n398 185
R71 source.n288 source.n287 185
R72 source.n405 source.n404 185
R73 source.n407 source.n406 185
R74 source.n284 source.n283 185
R75 source.n413 source.n412 185
R76 source.n415 source.n414 185
R77 source.n135 source.n134 185
R78 source.n133 source.n132 185
R79 source.n4 source.n3 185
R80 source.n127 source.n126 185
R81 source.n125 source.n124 185
R82 source.n8 source.n7 185
R83 source.n119 source.n118 185
R84 source.n117 source.n116 185
R85 source.n115 source.n11 185
R86 source.n15 source.n12 185
R87 source.n110 source.n109 185
R88 source.n108 source.n107 185
R89 source.n17 source.n16 185
R90 source.n102 source.n101 185
R91 source.n100 source.n99 185
R92 source.n21 source.n20 185
R93 source.n94 source.n93 185
R94 source.n92 source.n91 185
R95 source.n25 source.n24 185
R96 source.n86 source.n85 185
R97 source.n84 source.n83 185
R98 source.n29 source.n28 185
R99 source.n78 source.n77 185
R100 source.n76 source.n75 185
R101 source.n33 source.n32 185
R102 source.n70 source.n69 185
R103 source.n68 source.n35 185
R104 source.n67 source.n66 185
R105 source.n38 source.n36 185
R106 source.n61 source.n60 185
R107 source.n59 source.n58 185
R108 source.n42 source.n41 185
R109 source.n53 source.n52 185
R110 source.n51 source.n50 185
R111 source.n46 source.n45 185
R112 source.n275 source.n274 185
R113 source.n273 source.n272 185
R114 source.n144 source.n143 185
R115 source.n267 source.n266 185
R116 source.n265 source.n264 185
R117 source.n148 source.n147 185
R118 source.n259 source.n258 185
R119 source.n257 source.n256 185
R120 source.n255 source.n151 185
R121 source.n155 source.n152 185
R122 source.n250 source.n249 185
R123 source.n248 source.n247 185
R124 source.n157 source.n156 185
R125 source.n242 source.n241 185
R126 source.n240 source.n239 185
R127 source.n161 source.n160 185
R128 source.n234 source.n233 185
R129 source.n232 source.n231 185
R130 source.n165 source.n164 185
R131 source.n226 source.n225 185
R132 source.n224 source.n223 185
R133 source.n169 source.n168 185
R134 source.n218 source.n217 185
R135 source.n216 source.n215 185
R136 source.n173 source.n172 185
R137 source.n210 source.n209 185
R138 source.n208 source.n175 185
R139 source.n207 source.n206 185
R140 source.n178 source.n176 185
R141 source.n201 source.n200 185
R142 source.n199 source.n198 185
R143 source.n182 source.n181 185
R144 source.n193 source.n192 185
R145 source.n191 source.n190 185
R146 source.n186 source.n185 185
R147 source.n465 source.t3 149.524
R148 source.n325 source.t1 149.524
R149 source.n47 source.t0 149.524
R150 source.n187 source.t2 149.524
R151 source.n469 source.n463 104.615
R152 source.n470 source.n469 104.615
R153 source.n470 source.n459 104.615
R154 source.n477 source.n459 104.615
R155 source.n478 source.n477 104.615
R156 source.n478 source.n455 104.615
R157 source.n486 source.n455 104.615
R158 source.n487 source.n486 104.615
R159 source.n488 source.n487 104.615
R160 source.n488 source.n451 104.615
R161 source.n495 source.n451 104.615
R162 source.n496 source.n495 104.615
R163 source.n496 source.n447 104.615
R164 source.n503 source.n447 104.615
R165 source.n504 source.n503 104.615
R166 source.n504 source.n443 104.615
R167 source.n511 source.n443 104.615
R168 source.n512 source.n511 104.615
R169 source.n512 source.n439 104.615
R170 source.n519 source.n439 104.615
R171 source.n520 source.n519 104.615
R172 source.n520 source.n435 104.615
R173 source.n527 source.n435 104.615
R174 source.n529 source.n527 104.615
R175 source.n529 source.n528 104.615
R176 source.n528 source.n431 104.615
R177 source.n537 source.n431 104.615
R178 source.n538 source.n537 104.615
R179 source.n538 source.n427 104.615
R180 source.n545 source.n427 104.615
R181 source.n546 source.n545 104.615
R182 source.n546 source.n423 104.615
R183 source.n553 source.n423 104.615
R184 source.n554 source.n553 104.615
R185 source.n329 source.n323 104.615
R186 source.n330 source.n329 104.615
R187 source.n330 source.n319 104.615
R188 source.n337 source.n319 104.615
R189 source.n338 source.n337 104.615
R190 source.n338 source.n315 104.615
R191 source.n346 source.n315 104.615
R192 source.n347 source.n346 104.615
R193 source.n348 source.n347 104.615
R194 source.n348 source.n311 104.615
R195 source.n355 source.n311 104.615
R196 source.n356 source.n355 104.615
R197 source.n356 source.n307 104.615
R198 source.n363 source.n307 104.615
R199 source.n364 source.n363 104.615
R200 source.n364 source.n303 104.615
R201 source.n371 source.n303 104.615
R202 source.n372 source.n371 104.615
R203 source.n372 source.n299 104.615
R204 source.n379 source.n299 104.615
R205 source.n380 source.n379 104.615
R206 source.n380 source.n295 104.615
R207 source.n387 source.n295 104.615
R208 source.n389 source.n387 104.615
R209 source.n389 source.n388 104.615
R210 source.n388 source.n291 104.615
R211 source.n397 source.n291 104.615
R212 source.n398 source.n397 104.615
R213 source.n398 source.n287 104.615
R214 source.n405 source.n287 104.615
R215 source.n406 source.n405 104.615
R216 source.n406 source.n283 104.615
R217 source.n413 source.n283 104.615
R218 source.n414 source.n413 104.615
R219 source.n134 source.n133 104.615
R220 source.n133 source.n3 104.615
R221 source.n126 source.n3 104.615
R222 source.n126 source.n125 104.615
R223 source.n125 source.n7 104.615
R224 source.n118 source.n7 104.615
R225 source.n118 source.n117 104.615
R226 source.n117 source.n11 104.615
R227 source.n15 source.n11 104.615
R228 source.n109 source.n15 104.615
R229 source.n109 source.n108 104.615
R230 source.n108 source.n16 104.615
R231 source.n101 source.n16 104.615
R232 source.n101 source.n100 104.615
R233 source.n100 source.n20 104.615
R234 source.n93 source.n20 104.615
R235 source.n93 source.n92 104.615
R236 source.n92 source.n24 104.615
R237 source.n85 source.n24 104.615
R238 source.n85 source.n84 104.615
R239 source.n84 source.n28 104.615
R240 source.n77 source.n28 104.615
R241 source.n77 source.n76 104.615
R242 source.n76 source.n32 104.615
R243 source.n69 source.n32 104.615
R244 source.n69 source.n68 104.615
R245 source.n68 source.n67 104.615
R246 source.n67 source.n36 104.615
R247 source.n60 source.n36 104.615
R248 source.n60 source.n59 104.615
R249 source.n59 source.n41 104.615
R250 source.n52 source.n41 104.615
R251 source.n52 source.n51 104.615
R252 source.n51 source.n45 104.615
R253 source.n274 source.n273 104.615
R254 source.n273 source.n143 104.615
R255 source.n266 source.n143 104.615
R256 source.n266 source.n265 104.615
R257 source.n265 source.n147 104.615
R258 source.n258 source.n147 104.615
R259 source.n258 source.n257 104.615
R260 source.n257 source.n151 104.615
R261 source.n155 source.n151 104.615
R262 source.n249 source.n155 104.615
R263 source.n249 source.n248 104.615
R264 source.n248 source.n156 104.615
R265 source.n241 source.n156 104.615
R266 source.n241 source.n240 104.615
R267 source.n240 source.n160 104.615
R268 source.n233 source.n160 104.615
R269 source.n233 source.n232 104.615
R270 source.n232 source.n164 104.615
R271 source.n225 source.n164 104.615
R272 source.n225 source.n224 104.615
R273 source.n224 source.n168 104.615
R274 source.n217 source.n168 104.615
R275 source.n217 source.n216 104.615
R276 source.n216 source.n172 104.615
R277 source.n209 source.n172 104.615
R278 source.n209 source.n208 104.615
R279 source.n208 source.n207 104.615
R280 source.n207 source.n176 104.615
R281 source.n200 source.n176 104.615
R282 source.n200 source.n199 104.615
R283 source.n199 source.n181 104.615
R284 source.n192 source.n181 104.615
R285 source.n192 source.n191 104.615
R286 source.n191 source.n185 104.615
R287 source.t3 source.n463 52.3082
R288 source.t1 source.n323 52.3082
R289 source.t0 source.n45 52.3082
R290 source.t2 source.n185 52.3082
R291 source.n419 source.n279 32.9272
R292 source.n559 source.n558 30.6338
R293 source.n419 source.n418 30.6338
R294 source.n139 source.n138 30.6338
R295 source.n279 source.n278 30.6338
R296 source.n560 source.n139 26.3324
R297 source.n489 source.n454 13.1884
R298 source.n536 source.n535 13.1884
R299 source.n349 source.n314 13.1884
R300 source.n396 source.n395 13.1884
R301 source.n116 source.n115 13.1884
R302 source.n70 source.n35 13.1884
R303 source.n256 source.n255 13.1884
R304 source.n210 source.n175 13.1884
R305 source.n485 source.n484 12.8005
R306 source.n490 source.n452 12.8005
R307 source.n534 source.n432 12.8005
R308 source.n539 source.n430 12.8005
R309 source.n345 source.n344 12.8005
R310 source.n350 source.n312 12.8005
R311 source.n394 source.n292 12.8005
R312 source.n399 source.n290 12.8005
R313 source.n119 source.n10 12.8005
R314 source.n114 source.n12 12.8005
R315 source.n71 source.n33 12.8005
R316 source.n66 source.n37 12.8005
R317 source.n259 source.n150 12.8005
R318 source.n254 source.n152 12.8005
R319 source.n211 source.n173 12.8005
R320 source.n206 source.n177 12.8005
R321 source.n483 source.n456 12.0247
R322 source.n494 source.n493 12.0247
R323 source.n531 source.n530 12.0247
R324 source.n540 source.n428 12.0247
R325 source.n343 source.n316 12.0247
R326 source.n354 source.n353 12.0247
R327 source.n391 source.n390 12.0247
R328 source.n400 source.n288 12.0247
R329 source.n120 source.n8 12.0247
R330 source.n111 source.n110 12.0247
R331 source.n75 source.n74 12.0247
R332 source.n65 source.n38 12.0247
R333 source.n260 source.n148 12.0247
R334 source.n251 source.n250 12.0247
R335 source.n215 source.n214 12.0247
R336 source.n205 source.n178 12.0247
R337 source.n480 source.n479 11.249
R338 source.n497 source.n450 11.249
R339 source.n526 source.n434 11.249
R340 source.n544 source.n543 11.249
R341 source.n340 source.n339 11.249
R342 source.n357 source.n310 11.249
R343 source.n386 source.n294 11.249
R344 source.n404 source.n403 11.249
R345 source.n124 source.n123 11.249
R346 source.n107 source.n14 11.249
R347 source.n78 source.n31 11.249
R348 source.n62 source.n61 11.249
R349 source.n264 source.n263 11.249
R350 source.n247 source.n154 11.249
R351 source.n218 source.n171 11.249
R352 source.n202 source.n201 11.249
R353 source.n476 source.n458 10.4732
R354 source.n498 source.n448 10.4732
R355 source.n525 source.n436 10.4732
R356 source.n547 source.n426 10.4732
R357 source.n336 source.n318 10.4732
R358 source.n358 source.n308 10.4732
R359 source.n385 source.n296 10.4732
R360 source.n407 source.n286 10.4732
R361 source.n127 source.n6 10.4732
R362 source.n106 source.n17 10.4732
R363 source.n79 source.n29 10.4732
R364 source.n58 source.n40 10.4732
R365 source.n267 source.n146 10.4732
R366 source.n246 source.n157 10.4732
R367 source.n219 source.n169 10.4732
R368 source.n198 source.n180 10.4732
R369 source.n465 source.n464 10.2747
R370 source.n325 source.n324 10.2747
R371 source.n47 source.n46 10.2747
R372 source.n187 source.n186 10.2747
R373 source.n475 source.n460 9.69747
R374 source.n502 source.n501 9.69747
R375 source.n522 source.n521 9.69747
R376 source.n548 source.n424 9.69747
R377 source.n335 source.n320 9.69747
R378 source.n362 source.n361 9.69747
R379 source.n382 source.n381 9.69747
R380 source.n408 source.n284 9.69747
R381 source.n128 source.n4 9.69747
R382 source.n103 source.n102 9.69747
R383 source.n83 source.n82 9.69747
R384 source.n57 source.n42 9.69747
R385 source.n268 source.n144 9.69747
R386 source.n243 source.n242 9.69747
R387 source.n223 source.n222 9.69747
R388 source.n197 source.n182 9.69747
R389 source.n558 source.n557 9.45567
R390 source.n418 source.n417 9.45567
R391 source.n138 source.n137 9.45567
R392 source.n278 source.n277 9.45567
R393 source.n422 source.n421 9.3005
R394 source.n551 source.n550 9.3005
R395 source.n549 source.n548 9.3005
R396 source.n426 source.n425 9.3005
R397 source.n543 source.n542 9.3005
R398 source.n541 source.n540 9.3005
R399 source.n430 source.n429 9.3005
R400 source.n509 source.n508 9.3005
R401 source.n507 source.n506 9.3005
R402 source.n446 source.n445 9.3005
R403 source.n501 source.n500 9.3005
R404 source.n499 source.n498 9.3005
R405 source.n450 source.n449 9.3005
R406 source.n493 source.n492 9.3005
R407 source.n491 source.n490 9.3005
R408 source.n467 source.n466 9.3005
R409 source.n462 source.n461 9.3005
R410 source.n473 source.n472 9.3005
R411 source.n475 source.n474 9.3005
R412 source.n458 source.n457 9.3005
R413 source.n481 source.n480 9.3005
R414 source.n483 source.n482 9.3005
R415 source.n484 source.n453 9.3005
R416 source.n442 source.n441 9.3005
R417 source.n515 source.n514 9.3005
R418 source.n517 source.n516 9.3005
R419 source.n438 source.n437 9.3005
R420 source.n523 source.n522 9.3005
R421 source.n525 source.n524 9.3005
R422 source.n434 source.n433 9.3005
R423 source.n532 source.n531 9.3005
R424 source.n534 source.n533 9.3005
R425 source.n557 source.n556 9.3005
R426 source.n282 source.n281 9.3005
R427 source.n411 source.n410 9.3005
R428 source.n409 source.n408 9.3005
R429 source.n286 source.n285 9.3005
R430 source.n403 source.n402 9.3005
R431 source.n401 source.n400 9.3005
R432 source.n290 source.n289 9.3005
R433 source.n369 source.n368 9.3005
R434 source.n367 source.n366 9.3005
R435 source.n306 source.n305 9.3005
R436 source.n361 source.n360 9.3005
R437 source.n359 source.n358 9.3005
R438 source.n310 source.n309 9.3005
R439 source.n353 source.n352 9.3005
R440 source.n351 source.n350 9.3005
R441 source.n327 source.n326 9.3005
R442 source.n322 source.n321 9.3005
R443 source.n333 source.n332 9.3005
R444 source.n335 source.n334 9.3005
R445 source.n318 source.n317 9.3005
R446 source.n341 source.n340 9.3005
R447 source.n343 source.n342 9.3005
R448 source.n344 source.n313 9.3005
R449 source.n302 source.n301 9.3005
R450 source.n375 source.n374 9.3005
R451 source.n377 source.n376 9.3005
R452 source.n298 source.n297 9.3005
R453 source.n383 source.n382 9.3005
R454 source.n385 source.n384 9.3005
R455 source.n294 source.n293 9.3005
R456 source.n392 source.n391 9.3005
R457 source.n394 source.n393 9.3005
R458 source.n417 source.n416 9.3005
R459 source.n49 source.n48 9.3005
R460 source.n44 source.n43 9.3005
R461 source.n55 source.n54 9.3005
R462 source.n57 source.n56 9.3005
R463 source.n40 source.n39 9.3005
R464 source.n63 source.n62 9.3005
R465 source.n65 source.n64 9.3005
R466 source.n37 source.n34 9.3005
R467 source.n96 source.n95 9.3005
R468 source.n98 source.n97 9.3005
R469 source.n19 source.n18 9.3005
R470 source.n104 source.n103 9.3005
R471 source.n106 source.n105 9.3005
R472 source.n14 source.n13 9.3005
R473 source.n112 source.n111 9.3005
R474 source.n114 source.n113 9.3005
R475 source.n137 source.n136 9.3005
R476 source.n2 source.n1 9.3005
R477 source.n131 source.n130 9.3005
R478 source.n129 source.n128 9.3005
R479 source.n6 source.n5 9.3005
R480 source.n123 source.n122 9.3005
R481 source.n121 source.n120 9.3005
R482 source.n10 source.n9 9.3005
R483 source.n23 source.n22 9.3005
R484 source.n90 source.n89 9.3005
R485 source.n88 source.n87 9.3005
R486 source.n27 source.n26 9.3005
R487 source.n82 source.n81 9.3005
R488 source.n80 source.n79 9.3005
R489 source.n31 source.n30 9.3005
R490 source.n74 source.n73 9.3005
R491 source.n72 source.n71 9.3005
R492 source.n189 source.n188 9.3005
R493 source.n184 source.n183 9.3005
R494 source.n195 source.n194 9.3005
R495 source.n197 source.n196 9.3005
R496 source.n180 source.n179 9.3005
R497 source.n203 source.n202 9.3005
R498 source.n205 source.n204 9.3005
R499 source.n177 source.n174 9.3005
R500 source.n236 source.n235 9.3005
R501 source.n238 source.n237 9.3005
R502 source.n159 source.n158 9.3005
R503 source.n244 source.n243 9.3005
R504 source.n246 source.n245 9.3005
R505 source.n154 source.n153 9.3005
R506 source.n252 source.n251 9.3005
R507 source.n254 source.n253 9.3005
R508 source.n277 source.n276 9.3005
R509 source.n142 source.n141 9.3005
R510 source.n271 source.n270 9.3005
R511 source.n269 source.n268 9.3005
R512 source.n146 source.n145 9.3005
R513 source.n263 source.n262 9.3005
R514 source.n261 source.n260 9.3005
R515 source.n150 source.n149 9.3005
R516 source.n163 source.n162 9.3005
R517 source.n230 source.n229 9.3005
R518 source.n228 source.n227 9.3005
R519 source.n167 source.n166 9.3005
R520 source.n222 source.n221 9.3005
R521 source.n220 source.n219 9.3005
R522 source.n171 source.n170 9.3005
R523 source.n214 source.n213 9.3005
R524 source.n212 source.n211 9.3005
R525 source.n472 source.n471 8.92171
R526 source.n505 source.n446 8.92171
R527 source.n518 source.n438 8.92171
R528 source.n552 source.n551 8.92171
R529 source.n332 source.n331 8.92171
R530 source.n365 source.n306 8.92171
R531 source.n378 source.n298 8.92171
R532 source.n412 source.n411 8.92171
R533 source.n132 source.n131 8.92171
R534 source.n99 source.n19 8.92171
R535 source.n86 source.n27 8.92171
R536 source.n54 source.n53 8.92171
R537 source.n272 source.n271 8.92171
R538 source.n239 source.n159 8.92171
R539 source.n226 source.n167 8.92171
R540 source.n194 source.n193 8.92171
R541 source.n468 source.n462 8.14595
R542 source.n506 source.n444 8.14595
R543 source.n517 source.n440 8.14595
R544 source.n555 source.n422 8.14595
R545 source.n328 source.n322 8.14595
R546 source.n366 source.n304 8.14595
R547 source.n377 source.n300 8.14595
R548 source.n415 source.n282 8.14595
R549 source.n135 source.n2 8.14595
R550 source.n98 source.n21 8.14595
R551 source.n87 source.n25 8.14595
R552 source.n50 source.n44 8.14595
R553 source.n275 source.n142 8.14595
R554 source.n238 source.n161 8.14595
R555 source.n227 source.n165 8.14595
R556 source.n190 source.n184 8.14595
R557 source.n467 source.n464 7.3702
R558 source.n510 source.n509 7.3702
R559 source.n514 source.n513 7.3702
R560 source.n556 source.n420 7.3702
R561 source.n327 source.n324 7.3702
R562 source.n370 source.n369 7.3702
R563 source.n374 source.n373 7.3702
R564 source.n416 source.n280 7.3702
R565 source.n136 source.n0 7.3702
R566 source.n95 source.n94 7.3702
R567 source.n91 source.n90 7.3702
R568 source.n49 source.n46 7.3702
R569 source.n276 source.n140 7.3702
R570 source.n235 source.n234 7.3702
R571 source.n231 source.n230 7.3702
R572 source.n189 source.n186 7.3702
R573 source.n510 source.n442 6.59444
R574 source.n513 source.n442 6.59444
R575 source.n558 source.n420 6.59444
R576 source.n370 source.n302 6.59444
R577 source.n373 source.n302 6.59444
R578 source.n418 source.n280 6.59444
R579 source.n138 source.n0 6.59444
R580 source.n94 source.n23 6.59444
R581 source.n91 source.n23 6.59444
R582 source.n278 source.n140 6.59444
R583 source.n234 source.n163 6.59444
R584 source.n231 source.n163 6.59444
R585 source.n468 source.n467 5.81868
R586 source.n509 source.n444 5.81868
R587 source.n514 source.n440 5.81868
R588 source.n556 source.n555 5.81868
R589 source.n328 source.n327 5.81868
R590 source.n369 source.n304 5.81868
R591 source.n374 source.n300 5.81868
R592 source.n416 source.n415 5.81868
R593 source.n136 source.n135 5.81868
R594 source.n95 source.n21 5.81868
R595 source.n90 source.n25 5.81868
R596 source.n50 source.n49 5.81868
R597 source.n276 source.n275 5.81868
R598 source.n235 source.n161 5.81868
R599 source.n230 source.n165 5.81868
R600 source.n190 source.n189 5.81868
R601 source.n560 source.n559 5.7074
R602 source.n471 source.n462 5.04292
R603 source.n506 source.n505 5.04292
R604 source.n518 source.n517 5.04292
R605 source.n552 source.n422 5.04292
R606 source.n331 source.n322 5.04292
R607 source.n366 source.n365 5.04292
R608 source.n378 source.n377 5.04292
R609 source.n412 source.n282 5.04292
R610 source.n132 source.n2 5.04292
R611 source.n99 source.n98 5.04292
R612 source.n87 source.n86 5.04292
R613 source.n53 source.n44 5.04292
R614 source.n272 source.n142 5.04292
R615 source.n239 source.n238 5.04292
R616 source.n227 source.n226 5.04292
R617 source.n193 source.n184 5.04292
R618 source.n472 source.n460 4.26717
R619 source.n502 source.n446 4.26717
R620 source.n521 source.n438 4.26717
R621 source.n551 source.n424 4.26717
R622 source.n332 source.n320 4.26717
R623 source.n362 source.n306 4.26717
R624 source.n381 source.n298 4.26717
R625 source.n411 source.n284 4.26717
R626 source.n131 source.n4 4.26717
R627 source.n102 source.n19 4.26717
R628 source.n83 source.n27 4.26717
R629 source.n54 source.n42 4.26717
R630 source.n271 source.n144 4.26717
R631 source.n242 source.n159 4.26717
R632 source.n223 source.n167 4.26717
R633 source.n194 source.n182 4.26717
R634 source.n476 source.n475 3.49141
R635 source.n501 source.n448 3.49141
R636 source.n522 source.n436 3.49141
R637 source.n548 source.n547 3.49141
R638 source.n336 source.n335 3.49141
R639 source.n361 source.n308 3.49141
R640 source.n382 source.n296 3.49141
R641 source.n408 source.n407 3.49141
R642 source.n128 source.n127 3.49141
R643 source.n103 source.n17 3.49141
R644 source.n82 source.n29 3.49141
R645 source.n58 source.n57 3.49141
R646 source.n268 source.n267 3.49141
R647 source.n243 source.n157 3.49141
R648 source.n222 source.n169 3.49141
R649 source.n198 source.n197 3.49141
R650 source.n48 source.n47 2.84303
R651 source.n188 source.n187 2.84303
R652 source.n466 source.n465 2.84303
R653 source.n326 source.n325 2.84303
R654 source.n479 source.n458 2.71565
R655 source.n498 source.n497 2.71565
R656 source.n526 source.n525 2.71565
R657 source.n544 source.n426 2.71565
R658 source.n339 source.n318 2.71565
R659 source.n358 source.n357 2.71565
R660 source.n386 source.n385 2.71565
R661 source.n404 source.n286 2.71565
R662 source.n124 source.n6 2.71565
R663 source.n107 source.n106 2.71565
R664 source.n79 source.n78 2.71565
R665 source.n61 source.n40 2.71565
R666 source.n264 source.n146 2.71565
R667 source.n247 source.n246 2.71565
R668 source.n219 source.n218 2.71565
R669 source.n201 source.n180 2.71565
R670 source.n480 source.n456 1.93989
R671 source.n494 source.n450 1.93989
R672 source.n530 source.n434 1.93989
R673 source.n543 source.n428 1.93989
R674 source.n340 source.n316 1.93989
R675 source.n354 source.n310 1.93989
R676 source.n390 source.n294 1.93989
R677 source.n403 source.n288 1.93989
R678 source.n123 source.n8 1.93989
R679 source.n110 source.n14 1.93989
R680 source.n75 source.n31 1.93989
R681 source.n62 source.n38 1.93989
R682 source.n263 source.n148 1.93989
R683 source.n250 source.n154 1.93989
R684 source.n215 source.n171 1.93989
R685 source.n202 source.n178 1.93989
R686 source.n485 source.n483 1.16414
R687 source.n493 source.n452 1.16414
R688 source.n531 source.n432 1.16414
R689 source.n540 source.n539 1.16414
R690 source.n345 source.n343 1.16414
R691 source.n353 source.n312 1.16414
R692 source.n391 source.n292 1.16414
R693 source.n400 source.n399 1.16414
R694 source.n120 source.n119 1.16414
R695 source.n111 source.n12 1.16414
R696 source.n74 source.n33 1.16414
R697 source.n66 source.n65 1.16414
R698 source.n260 source.n259 1.16414
R699 source.n251 source.n152 1.16414
R700 source.n214 source.n173 1.16414
R701 source.n206 source.n205 1.16414
R702 source.n279 source.n139 0.914293
R703 source.n559 source.n419 0.914293
R704 source.n484 source.n454 0.388379
R705 source.n490 source.n489 0.388379
R706 source.n535 source.n534 0.388379
R707 source.n536 source.n430 0.388379
R708 source.n344 source.n314 0.388379
R709 source.n350 source.n349 0.388379
R710 source.n395 source.n394 0.388379
R711 source.n396 source.n290 0.388379
R712 source.n116 source.n10 0.388379
R713 source.n115 source.n114 0.388379
R714 source.n71 source.n70 0.388379
R715 source.n37 source.n35 0.388379
R716 source.n256 source.n150 0.388379
R717 source.n255 source.n254 0.388379
R718 source.n211 source.n210 0.388379
R719 source.n177 source.n175 0.388379
R720 source source.n560 0.188
R721 source.n466 source.n461 0.155672
R722 source.n473 source.n461 0.155672
R723 source.n474 source.n473 0.155672
R724 source.n474 source.n457 0.155672
R725 source.n481 source.n457 0.155672
R726 source.n482 source.n481 0.155672
R727 source.n482 source.n453 0.155672
R728 source.n491 source.n453 0.155672
R729 source.n492 source.n491 0.155672
R730 source.n492 source.n449 0.155672
R731 source.n499 source.n449 0.155672
R732 source.n500 source.n499 0.155672
R733 source.n500 source.n445 0.155672
R734 source.n507 source.n445 0.155672
R735 source.n508 source.n507 0.155672
R736 source.n508 source.n441 0.155672
R737 source.n515 source.n441 0.155672
R738 source.n516 source.n515 0.155672
R739 source.n516 source.n437 0.155672
R740 source.n523 source.n437 0.155672
R741 source.n524 source.n523 0.155672
R742 source.n524 source.n433 0.155672
R743 source.n532 source.n433 0.155672
R744 source.n533 source.n532 0.155672
R745 source.n533 source.n429 0.155672
R746 source.n541 source.n429 0.155672
R747 source.n542 source.n541 0.155672
R748 source.n542 source.n425 0.155672
R749 source.n549 source.n425 0.155672
R750 source.n550 source.n549 0.155672
R751 source.n550 source.n421 0.155672
R752 source.n557 source.n421 0.155672
R753 source.n326 source.n321 0.155672
R754 source.n333 source.n321 0.155672
R755 source.n334 source.n333 0.155672
R756 source.n334 source.n317 0.155672
R757 source.n341 source.n317 0.155672
R758 source.n342 source.n341 0.155672
R759 source.n342 source.n313 0.155672
R760 source.n351 source.n313 0.155672
R761 source.n352 source.n351 0.155672
R762 source.n352 source.n309 0.155672
R763 source.n359 source.n309 0.155672
R764 source.n360 source.n359 0.155672
R765 source.n360 source.n305 0.155672
R766 source.n367 source.n305 0.155672
R767 source.n368 source.n367 0.155672
R768 source.n368 source.n301 0.155672
R769 source.n375 source.n301 0.155672
R770 source.n376 source.n375 0.155672
R771 source.n376 source.n297 0.155672
R772 source.n383 source.n297 0.155672
R773 source.n384 source.n383 0.155672
R774 source.n384 source.n293 0.155672
R775 source.n392 source.n293 0.155672
R776 source.n393 source.n392 0.155672
R777 source.n393 source.n289 0.155672
R778 source.n401 source.n289 0.155672
R779 source.n402 source.n401 0.155672
R780 source.n402 source.n285 0.155672
R781 source.n409 source.n285 0.155672
R782 source.n410 source.n409 0.155672
R783 source.n410 source.n281 0.155672
R784 source.n417 source.n281 0.155672
R785 source.n137 source.n1 0.155672
R786 source.n130 source.n1 0.155672
R787 source.n130 source.n129 0.155672
R788 source.n129 source.n5 0.155672
R789 source.n122 source.n5 0.155672
R790 source.n122 source.n121 0.155672
R791 source.n121 source.n9 0.155672
R792 source.n113 source.n9 0.155672
R793 source.n113 source.n112 0.155672
R794 source.n112 source.n13 0.155672
R795 source.n105 source.n13 0.155672
R796 source.n105 source.n104 0.155672
R797 source.n104 source.n18 0.155672
R798 source.n97 source.n18 0.155672
R799 source.n97 source.n96 0.155672
R800 source.n96 source.n22 0.155672
R801 source.n89 source.n22 0.155672
R802 source.n89 source.n88 0.155672
R803 source.n88 source.n26 0.155672
R804 source.n81 source.n26 0.155672
R805 source.n81 source.n80 0.155672
R806 source.n80 source.n30 0.155672
R807 source.n73 source.n30 0.155672
R808 source.n73 source.n72 0.155672
R809 source.n72 source.n34 0.155672
R810 source.n64 source.n34 0.155672
R811 source.n64 source.n63 0.155672
R812 source.n63 source.n39 0.155672
R813 source.n56 source.n39 0.155672
R814 source.n56 source.n55 0.155672
R815 source.n55 source.n43 0.155672
R816 source.n48 source.n43 0.155672
R817 source.n277 source.n141 0.155672
R818 source.n270 source.n141 0.155672
R819 source.n270 source.n269 0.155672
R820 source.n269 source.n145 0.155672
R821 source.n262 source.n145 0.155672
R822 source.n262 source.n261 0.155672
R823 source.n261 source.n149 0.155672
R824 source.n253 source.n149 0.155672
R825 source.n253 source.n252 0.155672
R826 source.n252 source.n153 0.155672
R827 source.n245 source.n153 0.155672
R828 source.n245 source.n244 0.155672
R829 source.n244 source.n158 0.155672
R830 source.n237 source.n158 0.155672
R831 source.n237 source.n236 0.155672
R832 source.n236 source.n162 0.155672
R833 source.n229 source.n162 0.155672
R834 source.n229 source.n228 0.155672
R835 source.n228 source.n166 0.155672
R836 source.n221 source.n166 0.155672
R837 source.n221 source.n220 0.155672
R838 source.n220 source.n170 0.155672
R839 source.n213 source.n170 0.155672
R840 source.n213 source.n212 0.155672
R841 source.n212 source.n174 0.155672
R842 source.n204 source.n174 0.155672
R843 source.n204 source.n203 0.155672
R844 source.n203 source.n179 0.155672
R845 source.n196 source.n179 0.155672
R846 source.n196 source.n195 0.155672
R847 source.n195 source.n183 0.155672
R848 source.n188 source.n183 0.155672
R849 drain_right.n134 drain_right.n0 289.615
R850 drain_right.n273 drain_right.n139 289.615
R851 drain_right.n44 drain_right.n43 185
R852 drain_right.n49 drain_right.n48 185
R853 drain_right.n51 drain_right.n50 185
R854 drain_right.n40 drain_right.n39 185
R855 drain_right.n57 drain_right.n56 185
R856 drain_right.n59 drain_right.n58 185
R857 drain_right.n36 drain_right.n35 185
R858 drain_right.n66 drain_right.n65 185
R859 drain_right.n67 drain_right.n34 185
R860 drain_right.n69 drain_right.n68 185
R861 drain_right.n32 drain_right.n31 185
R862 drain_right.n75 drain_right.n74 185
R863 drain_right.n77 drain_right.n76 185
R864 drain_right.n28 drain_right.n27 185
R865 drain_right.n83 drain_right.n82 185
R866 drain_right.n85 drain_right.n84 185
R867 drain_right.n24 drain_right.n23 185
R868 drain_right.n91 drain_right.n90 185
R869 drain_right.n93 drain_right.n92 185
R870 drain_right.n20 drain_right.n19 185
R871 drain_right.n99 drain_right.n98 185
R872 drain_right.n101 drain_right.n100 185
R873 drain_right.n16 drain_right.n15 185
R874 drain_right.n107 drain_right.n106 185
R875 drain_right.n110 drain_right.n109 185
R876 drain_right.n108 drain_right.n12 185
R877 drain_right.n115 drain_right.n11 185
R878 drain_right.n117 drain_right.n116 185
R879 drain_right.n119 drain_right.n118 185
R880 drain_right.n8 drain_right.n7 185
R881 drain_right.n125 drain_right.n124 185
R882 drain_right.n127 drain_right.n126 185
R883 drain_right.n4 drain_right.n3 185
R884 drain_right.n133 drain_right.n132 185
R885 drain_right.n135 drain_right.n134 185
R886 drain_right.n274 drain_right.n273 185
R887 drain_right.n272 drain_right.n271 185
R888 drain_right.n143 drain_right.n142 185
R889 drain_right.n266 drain_right.n265 185
R890 drain_right.n264 drain_right.n263 185
R891 drain_right.n147 drain_right.n146 185
R892 drain_right.n258 drain_right.n257 185
R893 drain_right.n256 drain_right.n255 185
R894 drain_right.n254 drain_right.n150 185
R895 drain_right.n154 drain_right.n151 185
R896 drain_right.n249 drain_right.n248 185
R897 drain_right.n247 drain_right.n246 185
R898 drain_right.n156 drain_right.n155 185
R899 drain_right.n241 drain_right.n240 185
R900 drain_right.n239 drain_right.n238 185
R901 drain_right.n160 drain_right.n159 185
R902 drain_right.n233 drain_right.n232 185
R903 drain_right.n231 drain_right.n230 185
R904 drain_right.n164 drain_right.n163 185
R905 drain_right.n225 drain_right.n224 185
R906 drain_right.n223 drain_right.n222 185
R907 drain_right.n168 drain_right.n167 185
R908 drain_right.n217 drain_right.n216 185
R909 drain_right.n215 drain_right.n214 185
R910 drain_right.n172 drain_right.n171 185
R911 drain_right.n209 drain_right.n208 185
R912 drain_right.n207 drain_right.n174 185
R913 drain_right.n206 drain_right.n205 185
R914 drain_right.n177 drain_right.n175 185
R915 drain_right.n200 drain_right.n199 185
R916 drain_right.n198 drain_right.n197 185
R917 drain_right.n181 drain_right.n180 185
R918 drain_right.n192 drain_right.n191 185
R919 drain_right.n190 drain_right.n189 185
R920 drain_right.n185 drain_right.n184 185
R921 drain_right.n45 drain_right.t0 149.524
R922 drain_right.n186 drain_right.t1 149.524
R923 drain_right.n49 drain_right.n43 104.615
R924 drain_right.n50 drain_right.n49 104.615
R925 drain_right.n50 drain_right.n39 104.615
R926 drain_right.n57 drain_right.n39 104.615
R927 drain_right.n58 drain_right.n57 104.615
R928 drain_right.n58 drain_right.n35 104.615
R929 drain_right.n66 drain_right.n35 104.615
R930 drain_right.n67 drain_right.n66 104.615
R931 drain_right.n68 drain_right.n67 104.615
R932 drain_right.n68 drain_right.n31 104.615
R933 drain_right.n75 drain_right.n31 104.615
R934 drain_right.n76 drain_right.n75 104.615
R935 drain_right.n76 drain_right.n27 104.615
R936 drain_right.n83 drain_right.n27 104.615
R937 drain_right.n84 drain_right.n83 104.615
R938 drain_right.n84 drain_right.n23 104.615
R939 drain_right.n91 drain_right.n23 104.615
R940 drain_right.n92 drain_right.n91 104.615
R941 drain_right.n92 drain_right.n19 104.615
R942 drain_right.n99 drain_right.n19 104.615
R943 drain_right.n100 drain_right.n99 104.615
R944 drain_right.n100 drain_right.n15 104.615
R945 drain_right.n107 drain_right.n15 104.615
R946 drain_right.n109 drain_right.n107 104.615
R947 drain_right.n109 drain_right.n108 104.615
R948 drain_right.n108 drain_right.n11 104.615
R949 drain_right.n117 drain_right.n11 104.615
R950 drain_right.n118 drain_right.n117 104.615
R951 drain_right.n118 drain_right.n7 104.615
R952 drain_right.n125 drain_right.n7 104.615
R953 drain_right.n126 drain_right.n125 104.615
R954 drain_right.n126 drain_right.n3 104.615
R955 drain_right.n133 drain_right.n3 104.615
R956 drain_right.n134 drain_right.n133 104.615
R957 drain_right.n273 drain_right.n272 104.615
R958 drain_right.n272 drain_right.n142 104.615
R959 drain_right.n265 drain_right.n142 104.615
R960 drain_right.n265 drain_right.n264 104.615
R961 drain_right.n264 drain_right.n146 104.615
R962 drain_right.n257 drain_right.n146 104.615
R963 drain_right.n257 drain_right.n256 104.615
R964 drain_right.n256 drain_right.n150 104.615
R965 drain_right.n154 drain_right.n150 104.615
R966 drain_right.n248 drain_right.n154 104.615
R967 drain_right.n248 drain_right.n247 104.615
R968 drain_right.n247 drain_right.n155 104.615
R969 drain_right.n240 drain_right.n155 104.615
R970 drain_right.n240 drain_right.n239 104.615
R971 drain_right.n239 drain_right.n159 104.615
R972 drain_right.n232 drain_right.n159 104.615
R973 drain_right.n232 drain_right.n231 104.615
R974 drain_right.n231 drain_right.n163 104.615
R975 drain_right.n224 drain_right.n163 104.615
R976 drain_right.n224 drain_right.n223 104.615
R977 drain_right.n223 drain_right.n167 104.615
R978 drain_right.n216 drain_right.n167 104.615
R979 drain_right.n216 drain_right.n215 104.615
R980 drain_right.n215 drain_right.n171 104.615
R981 drain_right.n208 drain_right.n171 104.615
R982 drain_right.n208 drain_right.n207 104.615
R983 drain_right.n207 drain_right.n206 104.615
R984 drain_right.n206 drain_right.n175 104.615
R985 drain_right.n199 drain_right.n175 104.615
R986 drain_right.n199 drain_right.n198 104.615
R987 drain_right.n198 drain_right.n180 104.615
R988 drain_right.n191 drain_right.n180 104.615
R989 drain_right.n191 drain_right.n190 104.615
R990 drain_right.n190 drain_right.n184 104.615
R991 drain_right drain_right.n138 85.2662
R992 drain_right drain_right.n277 53.4093
R993 drain_right.t0 drain_right.n43 52.3082
R994 drain_right.t1 drain_right.n184 52.3082
R995 drain_right.n69 drain_right.n34 13.1884
R996 drain_right.n116 drain_right.n115 13.1884
R997 drain_right.n255 drain_right.n254 13.1884
R998 drain_right.n209 drain_right.n174 13.1884
R999 drain_right.n65 drain_right.n64 12.8005
R1000 drain_right.n70 drain_right.n32 12.8005
R1001 drain_right.n114 drain_right.n12 12.8005
R1002 drain_right.n119 drain_right.n10 12.8005
R1003 drain_right.n258 drain_right.n149 12.8005
R1004 drain_right.n253 drain_right.n151 12.8005
R1005 drain_right.n210 drain_right.n172 12.8005
R1006 drain_right.n205 drain_right.n176 12.8005
R1007 drain_right.n63 drain_right.n36 12.0247
R1008 drain_right.n74 drain_right.n73 12.0247
R1009 drain_right.n111 drain_right.n110 12.0247
R1010 drain_right.n120 drain_right.n8 12.0247
R1011 drain_right.n259 drain_right.n147 12.0247
R1012 drain_right.n250 drain_right.n249 12.0247
R1013 drain_right.n214 drain_right.n213 12.0247
R1014 drain_right.n204 drain_right.n177 12.0247
R1015 drain_right.n60 drain_right.n59 11.249
R1016 drain_right.n77 drain_right.n30 11.249
R1017 drain_right.n106 drain_right.n14 11.249
R1018 drain_right.n124 drain_right.n123 11.249
R1019 drain_right.n263 drain_right.n262 11.249
R1020 drain_right.n246 drain_right.n153 11.249
R1021 drain_right.n217 drain_right.n170 11.249
R1022 drain_right.n201 drain_right.n200 11.249
R1023 drain_right.n56 drain_right.n38 10.4732
R1024 drain_right.n78 drain_right.n28 10.4732
R1025 drain_right.n105 drain_right.n16 10.4732
R1026 drain_right.n127 drain_right.n6 10.4732
R1027 drain_right.n266 drain_right.n145 10.4732
R1028 drain_right.n245 drain_right.n156 10.4732
R1029 drain_right.n218 drain_right.n168 10.4732
R1030 drain_right.n197 drain_right.n179 10.4732
R1031 drain_right.n45 drain_right.n44 10.2747
R1032 drain_right.n186 drain_right.n185 10.2747
R1033 drain_right.n55 drain_right.n40 9.69747
R1034 drain_right.n82 drain_right.n81 9.69747
R1035 drain_right.n102 drain_right.n101 9.69747
R1036 drain_right.n128 drain_right.n4 9.69747
R1037 drain_right.n267 drain_right.n143 9.69747
R1038 drain_right.n242 drain_right.n241 9.69747
R1039 drain_right.n222 drain_right.n221 9.69747
R1040 drain_right.n196 drain_right.n181 9.69747
R1041 drain_right.n138 drain_right.n137 9.45567
R1042 drain_right.n277 drain_right.n276 9.45567
R1043 drain_right.n2 drain_right.n1 9.3005
R1044 drain_right.n131 drain_right.n130 9.3005
R1045 drain_right.n129 drain_right.n128 9.3005
R1046 drain_right.n6 drain_right.n5 9.3005
R1047 drain_right.n123 drain_right.n122 9.3005
R1048 drain_right.n121 drain_right.n120 9.3005
R1049 drain_right.n10 drain_right.n9 9.3005
R1050 drain_right.n89 drain_right.n88 9.3005
R1051 drain_right.n87 drain_right.n86 9.3005
R1052 drain_right.n26 drain_right.n25 9.3005
R1053 drain_right.n81 drain_right.n80 9.3005
R1054 drain_right.n79 drain_right.n78 9.3005
R1055 drain_right.n30 drain_right.n29 9.3005
R1056 drain_right.n73 drain_right.n72 9.3005
R1057 drain_right.n71 drain_right.n70 9.3005
R1058 drain_right.n47 drain_right.n46 9.3005
R1059 drain_right.n42 drain_right.n41 9.3005
R1060 drain_right.n53 drain_right.n52 9.3005
R1061 drain_right.n55 drain_right.n54 9.3005
R1062 drain_right.n38 drain_right.n37 9.3005
R1063 drain_right.n61 drain_right.n60 9.3005
R1064 drain_right.n63 drain_right.n62 9.3005
R1065 drain_right.n64 drain_right.n33 9.3005
R1066 drain_right.n22 drain_right.n21 9.3005
R1067 drain_right.n95 drain_right.n94 9.3005
R1068 drain_right.n97 drain_right.n96 9.3005
R1069 drain_right.n18 drain_right.n17 9.3005
R1070 drain_right.n103 drain_right.n102 9.3005
R1071 drain_right.n105 drain_right.n104 9.3005
R1072 drain_right.n14 drain_right.n13 9.3005
R1073 drain_right.n112 drain_right.n111 9.3005
R1074 drain_right.n114 drain_right.n113 9.3005
R1075 drain_right.n137 drain_right.n136 9.3005
R1076 drain_right.n188 drain_right.n187 9.3005
R1077 drain_right.n183 drain_right.n182 9.3005
R1078 drain_right.n194 drain_right.n193 9.3005
R1079 drain_right.n196 drain_right.n195 9.3005
R1080 drain_right.n179 drain_right.n178 9.3005
R1081 drain_right.n202 drain_right.n201 9.3005
R1082 drain_right.n204 drain_right.n203 9.3005
R1083 drain_right.n176 drain_right.n173 9.3005
R1084 drain_right.n235 drain_right.n234 9.3005
R1085 drain_right.n237 drain_right.n236 9.3005
R1086 drain_right.n158 drain_right.n157 9.3005
R1087 drain_right.n243 drain_right.n242 9.3005
R1088 drain_right.n245 drain_right.n244 9.3005
R1089 drain_right.n153 drain_right.n152 9.3005
R1090 drain_right.n251 drain_right.n250 9.3005
R1091 drain_right.n253 drain_right.n252 9.3005
R1092 drain_right.n276 drain_right.n275 9.3005
R1093 drain_right.n141 drain_right.n140 9.3005
R1094 drain_right.n270 drain_right.n269 9.3005
R1095 drain_right.n268 drain_right.n267 9.3005
R1096 drain_right.n145 drain_right.n144 9.3005
R1097 drain_right.n262 drain_right.n261 9.3005
R1098 drain_right.n260 drain_right.n259 9.3005
R1099 drain_right.n149 drain_right.n148 9.3005
R1100 drain_right.n162 drain_right.n161 9.3005
R1101 drain_right.n229 drain_right.n228 9.3005
R1102 drain_right.n227 drain_right.n226 9.3005
R1103 drain_right.n166 drain_right.n165 9.3005
R1104 drain_right.n221 drain_right.n220 9.3005
R1105 drain_right.n219 drain_right.n218 9.3005
R1106 drain_right.n170 drain_right.n169 9.3005
R1107 drain_right.n213 drain_right.n212 9.3005
R1108 drain_right.n211 drain_right.n210 9.3005
R1109 drain_right.n52 drain_right.n51 8.92171
R1110 drain_right.n85 drain_right.n26 8.92171
R1111 drain_right.n98 drain_right.n18 8.92171
R1112 drain_right.n132 drain_right.n131 8.92171
R1113 drain_right.n271 drain_right.n270 8.92171
R1114 drain_right.n238 drain_right.n158 8.92171
R1115 drain_right.n225 drain_right.n166 8.92171
R1116 drain_right.n193 drain_right.n192 8.92171
R1117 drain_right.n48 drain_right.n42 8.14595
R1118 drain_right.n86 drain_right.n24 8.14595
R1119 drain_right.n97 drain_right.n20 8.14595
R1120 drain_right.n135 drain_right.n2 8.14595
R1121 drain_right.n274 drain_right.n141 8.14595
R1122 drain_right.n237 drain_right.n160 8.14595
R1123 drain_right.n226 drain_right.n164 8.14595
R1124 drain_right.n189 drain_right.n183 8.14595
R1125 drain_right.n47 drain_right.n44 7.3702
R1126 drain_right.n90 drain_right.n89 7.3702
R1127 drain_right.n94 drain_right.n93 7.3702
R1128 drain_right.n136 drain_right.n0 7.3702
R1129 drain_right.n275 drain_right.n139 7.3702
R1130 drain_right.n234 drain_right.n233 7.3702
R1131 drain_right.n230 drain_right.n229 7.3702
R1132 drain_right.n188 drain_right.n185 7.3702
R1133 drain_right.n90 drain_right.n22 6.59444
R1134 drain_right.n93 drain_right.n22 6.59444
R1135 drain_right.n138 drain_right.n0 6.59444
R1136 drain_right.n277 drain_right.n139 6.59444
R1137 drain_right.n233 drain_right.n162 6.59444
R1138 drain_right.n230 drain_right.n162 6.59444
R1139 drain_right.n48 drain_right.n47 5.81868
R1140 drain_right.n89 drain_right.n24 5.81868
R1141 drain_right.n94 drain_right.n20 5.81868
R1142 drain_right.n136 drain_right.n135 5.81868
R1143 drain_right.n275 drain_right.n274 5.81868
R1144 drain_right.n234 drain_right.n160 5.81868
R1145 drain_right.n229 drain_right.n164 5.81868
R1146 drain_right.n189 drain_right.n188 5.81868
R1147 drain_right.n51 drain_right.n42 5.04292
R1148 drain_right.n86 drain_right.n85 5.04292
R1149 drain_right.n98 drain_right.n97 5.04292
R1150 drain_right.n132 drain_right.n2 5.04292
R1151 drain_right.n271 drain_right.n141 5.04292
R1152 drain_right.n238 drain_right.n237 5.04292
R1153 drain_right.n226 drain_right.n225 5.04292
R1154 drain_right.n192 drain_right.n183 5.04292
R1155 drain_right.n52 drain_right.n40 4.26717
R1156 drain_right.n82 drain_right.n26 4.26717
R1157 drain_right.n101 drain_right.n18 4.26717
R1158 drain_right.n131 drain_right.n4 4.26717
R1159 drain_right.n270 drain_right.n143 4.26717
R1160 drain_right.n241 drain_right.n158 4.26717
R1161 drain_right.n222 drain_right.n166 4.26717
R1162 drain_right.n193 drain_right.n181 4.26717
R1163 drain_right.n56 drain_right.n55 3.49141
R1164 drain_right.n81 drain_right.n28 3.49141
R1165 drain_right.n102 drain_right.n16 3.49141
R1166 drain_right.n128 drain_right.n127 3.49141
R1167 drain_right.n267 drain_right.n266 3.49141
R1168 drain_right.n242 drain_right.n156 3.49141
R1169 drain_right.n221 drain_right.n168 3.49141
R1170 drain_right.n197 drain_right.n196 3.49141
R1171 drain_right.n187 drain_right.n186 2.84303
R1172 drain_right.n46 drain_right.n45 2.84303
R1173 drain_right.n59 drain_right.n38 2.71565
R1174 drain_right.n78 drain_right.n77 2.71565
R1175 drain_right.n106 drain_right.n105 2.71565
R1176 drain_right.n124 drain_right.n6 2.71565
R1177 drain_right.n263 drain_right.n145 2.71565
R1178 drain_right.n246 drain_right.n245 2.71565
R1179 drain_right.n218 drain_right.n217 2.71565
R1180 drain_right.n200 drain_right.n179 2.71565
R1181 drain_right.n60 drain_right.n36 1.93989
R1182 drain_right.n74 drain_right.n30 1.93989
R1183 drain_right.n110 drain_right.n14 1.93989
R1184 drain_right.n123 drain_right.n8 1.93989
R1185 drain_right.n262 drain_right.n147 1.93989
R1186 drain_right.n249 drain_right.n153 1.93989
R1187 drain_right.n214 drain_right.n170 1.93989
R1188 drain_right.n201 drain_right.n177 1.93989
R1189 drain_right.n65 drain_right.n63 1.16414
R1190 drain_right.n73 drain_right.n32 1.16414
R1191 drain_right.n111 drain_right.n12 1.16414
R1192 drain_right.n120 drain_right.n119 1.16414
R1193 drain_right.n259 drain_right.n258 1.16414
R1194 drain_right.n250 drain_right.n151 1.16414
R1195 drain_right.n213 drain_right.n172 1.16414
R1196 drain_right.n205 drain_right.n204 1.16414
R1197 drain_right.n64 drain_right.n34 0.388379
R1198 drain_right.n70 drain_right.n69 0.388379
R1199 drain_right.n115 drain_right.n114 0.388379
R1200 drain_right.n116 drain_right.n10 0.388379
R1201 drain_right.n255 drain_right.n149 0.388379
R1202 drain_right.n254 drain_right.n253 0.388379
R1203 drain_right.n210 drain_right.n209 0.388379
R1204 drain_right.n176 drain_right.n174 0.388379
R1205 drain_right.n46 drain_right.n41 0.155672
R1206 drain_right.n53 drain_right.n41 0.155672
R1207 drain_right.n54 drain_right.n53 0.155672
R1208 drain_right.n54 drain_right.n37 0.155672
R1209 drain_right.n61 drain_right.n37 0.155672
R1210 drain_right.n62 drain_right.n61 0.155672
R1211 drain_right.n62 drain_right.n33 0.155672
R1212 drain_right.n71 drain_right.n33 0.155672
R1213 drain_right.n72 drain_right.n71 0.155672
R1214 drain_right.n72 drain_right.n29 0.155672
R1215 drain_right.n79 drain_right.n29 0.155672
R1216 drain_right.n80 drain_right.n79 0.155672
R1217 drain_right.n80 drain_right.n25 0.155672
R1218 drain_right.n87 drain_right.n25 0.155672
R1219 drain_right.n88 drain_right.n87 0.155672
R1220 drain_right.n88 drain_right.n21 0.155672
R1221 drain_right.n95 drain_right.n21 0.155672
R1222 drain_right.n96 drain_right.n95 0.155672
R1223 drain_right.n96 drain_right.n17 0.155672
R1224 drain_right.n103 drain_right.n17 0.155672
R1225 drain_right.n104 drain_right.n103 0.155672
R1226 drain_right.n104 drain_right.n13 0.155672
R1227 drain_right.n112 drain_right.n13 0.155672
R1228 drain_right.n113 drain_right.n112 0.155672
R1229 drain_right.n113 drain_right.n9 0.155672
R1230 drain_right.n121 drain_right.n9 0.155672
R1231 drain_right.n122 drain_right.n121 0.155672
R1232 drain_right.n122 drain_right.n5 0.155672
R1233 drain_right.n129 drain_right.n5 0.155672
R1234 drain_right.n130 drain_right.n129 0.155672
R1235 drain_right.n130 drain_right.n1 0.155672
R1236 drain_right.n137 drain_right.n1 0.155672
R1237 drain_right.n276 drain_right.n140 0.155672
R1238 drain_right.n269 drain_right.n140 0.155672
R1239 drain_right.n269 drain_right.n268 0.155672
R1240 drain_right.n268 drain_right.n144 0.155672
R1241 drain_right.n261 drain_right.n144 0.155672
R1242 drain_right.n261 drain_right.n260 0.155672
R1243 drain_right.n260 drain_right.n148 0.155672
R1244 drain_right.n252 drain_right.n148 0.155672
R1245 drain_right.n252 drain_right.n251 0.155672
R1246 drain_right.n251 drain_right.n152 0.155672
R1247 drain_right.n244 drain_right.n152 0.155672
R1248 drain_right.n244 drain_right.n243 0.155672
R1249 drain_right.n243 drain_right.n157 0.155672
R1250 drain_right.n236 drain_right.n157 0.155672
R1251 drain_right.n236 drain_right.n235 0.155672
R1252 drain_right.n235 drain_right.n161 0.155672
R1253 drain_right.n228 drain_right.n161 0.155672
R1254 drain_right.n228 drain_right.n227 0.155672
R1255 drain_right.n227 drain_right.n165 0.155672
R1256 drain_right.n220 drain_right.n165 0.155672
R1257 drain_right.n220 drain_right.n219 0.155672
R1258 drain_right.n219 drain_right.n169 0.155672
R1259 drain_right.n212 drain_right.n169 0.155672
R1260 drain_right.n212 drain_right.n211 0.155672
R1261 drain_right.n211 drain_right.n173 0.155672
R1262 drain_right.n203 drain_right.n173 0.155672
R1263 drain_right.n203 drain_right.n202 0.155672
R1264 drain_right.n202 drain_right.n178 0.155672
R1265 drain_right.n195 drain_right.n178 0.155672
R1266 drain_right.n195 drain_right.n194 0.155672
R1267 drain_right.n194 drain_right.n182 0.155672
R1268 drain_right.n187 drain_right.n182 0.155672
R1269 plus plus.t0 1110.46
R1270 plus plus.t1 1095.32
R1271 drain_left.n134 drain_left.n0 289.615
R1272 drain_left.n273 drain_left.n139 289.615
R1273 drain_left.n44 drain_left.n43 185
R1274 drain_left.n49 drain_left.n48 185
R1275 drain_left.n51 drain_left.n50 185
R1276 drain_left.n40 drain_left.n39 185
R1277 drain_left.n57 drain_left.n56 185
R1278 drain_left.n59 drain_left.n58 185
R1279 drain_left.n36 drain_left.n35 185
R1280 drain_left.n66 drain_left.n65 185
R1281 drain_left.n67 drain_left.n34 185
R1282 drain_left.n69 drain_left.n68 185
R1283 drain_left.n32 drain_left.n31 185
R1284 drain_left.n75 drain_left.n74 185
R1285 drain_left.n77 drain_left.n76 185
R1286 drain_left.n28 drain_left.n27 185
R1287 drain_left.n83 drain_left.n82 185
R1288 drain_left.n85 drain_left.n84 185
R1289 drain_left.n24 drain_left.n23 185
R1290 drain_left.n91 drain_left.n90 185
R1291 drain_left.n93 drain_left.n92 185
R1292 drain_left.n20 drain_left.n19 185
R1293 drain_left.n99 drain_left.n98 185
R1294 drain_left.n101 drain_left.n100 185
R1295 drain_left.n16 drain_left.n15 185
R1296 drain_left.n107 drain_left.n106 185
R1297 drain_left.n110 drain_left.n109 185
R1298 drain_left.n108 drain_left.n12 185
R1299 drain_left.n115 drain_left.n11 185
R1300 drain_left.n117 drain_left.n116 185
R1301 drain_left.n119 drain_left.n118 185
R1302 drain_left.n8 drain_left.n7 185
R1303 drain_left.n125 drain_left.n124 185
R1304 drain_left.n127 drain_left.n126 185
R1305 drain_left.n4 drain_left.n3 185
R1306 drain_left.n133 drain_left.n132 185
R1307 drain_left.n135 drain_left.n134 185
R1308 drain_left.n274 drain_left.n273 185
R1309 drain_left.n272 drain_left.n271 185
R1310 drain_left.n143 drain_left.n142 185
R1311 drain_left.n266 drain_left.n265 185
R1312 drain_left.n264 drain_left.n263 185
R1313 drain_left.n147 drain_left.n146 185
R1314 drain_left.n258 drain_left.n257 185
R1315 drain_left.n256 drain_left.n255 185
R1316 drain_left.n254 drain_left.n150 185
R1317 drain_left.n154 drain_left.n151 185
R1318 drain_left.n249 drain_left.n248 185
R1319 drain_left.n247 drain_left.n246 185
R1320 drain_left.n156 drain_left.n155 185
R1321 drain_left.n241 drain_left.n240 185
R1322 drain_left.n239 drain_left.n238 185
R1323 drain_left.n160 drain_left.n159 185
R1324 drain_left.n233 drain_left.n232 185
R1325 drain_left.n231 drain_left.n230 185
R1326 drain_left.n164 drain_left.n163 185
R1327 drain_left.n225 drain_left.n224 185
R1328 drain_left.n223 drain_left.n222 185
R1329 drain_left.n168 drain_left.n167 185
R1330 drain_left.n217 drain_left.n216 185
R1331 drain_left.n215 drain_left.n214 185
R1332 drain_left.n172 drain_left.n171 185
R1333 drain_left.n209 drain_left.n208 185
R1334 drain_left.n207 drain_left.n174 185
R1335 drain_left.n206 drain_left.n205 185
R1336 drain_left.n177 drain_left.n175 185
R1337 drain_left.n200 drain_left.n199 185
R1338 drain_left.n198 drain_left.n197 185
R1339 drain_left.n181 drain_left.n180 185
R1340 drain_left.n192 drain_left.n191 185
R1341 drain_left.n190 drain_left.n189 185
R1342 drain_left.n185 drain_left.n184 185
R1343 drain_left.n45 drain_left.t1 149.524
R1344 drain_left.n186 drain_left.t0 149.524
R1345 drain_left.n49 drain_left.n43 104.615
R1346 drain_left.n50 drain_left.n49 104.615
R1347 drain_left.n50 drain_left.n39 104.615
R1348 drain_left.n57 drain_left.n39 104.615
R1349 drain_left.n58 drain_left.n57 104.615
R1350 drain_left.n58 drain_left.n35 104.615
R1351 drain_left.n66 drain_left.n35 104.615
R1352 drain_left.n67 drain_left.n66 104.615
R1353 drain_left.n68 drain_left.n67 104.615
R1354 drain_left.n68 drain_left.n31 104.615
R1355 drain_left.n75 drain_left.n31 104.615
R1356 drain_left.n76 drain_left.n75 104.615
R1357 drain_left.n76 drain_left.n27 104.615
R1358 drain_left.n83 drain_left.n27 104.615
R1359 drain_left.n84 drain_left.n83 104.615
R1360 drain_left.n84 drain_left.n23 104.615
R1361 drain_left.n91 drain_left.n23 104.615
R1362 drain_left.n92 drain_left.n91 104.615
R1363 drain_left.n92 drain_left.n19 104.615
R1364 drain_left.n99 drain_left.n19 104.615
R1365 drain_left.n100 drain_left.n99 104.615
R1366 drain_left.n100 drain_left.n15 104.615
R1367 drain_left.n107 drain_left.n15 104.615
R1368 drain_left.n109 drain_left.n107 104.615
R1369 drain_left.n109 drain_left.n108 104.615
R1370 drain_left.n108 drain_left.n11 104.615
R1371 drain_left.n117 drain_left.n11 104.615
R1372 drain_left.n118 drain_left.n117 104.615
R1373 drain_left.n118 drain_left.n7 104.615
R1374 drain_left.n125 drain_left.n7 104.615
R1375 drain_left.n126 drain_left.n125 104.615
R1376 drain_left.n126 drain_left.n3 104.615
R1377 drain_left.n133 drain_left.n3 104.615
R1378 drain_left.n134 drain_left.n133 104.615
R1379 drain_left.n273 drain_left.n272 104.615
R1380 drain_left.n272 drain_left.n142 104.615
R1381 drain_left.n265 drain_left.n142 104.615
R1382 drain_left.n265 drain_left.n264 104.615
R1383 drain_left.n264 drain_left.n146 104.615
R1384 drain_left.n257 drain_left.n146 104.615
R1385 drain_left.n257 drain_left.n256 104.615
R1386 drain_left.n256 drain_left.n150 104.615
R1387 drain_left.n154 drain_left.n150 104.615
R1388 drain_left.n248 drain_left.n154 104.615
R1389 drain_left.n248 drain_left.n247 104.615
R1390 drain_left.n247 drain_left.n155 104.615
R1391 drain_left.n240 drain_left.n155 104.615
R1392 drain_left.n240 drain_left.n239 104.615
R1393 drain_left.n239 drain_left.n159 104.615
R1394 drain_left.n232 drain_left.n159 104.615
R1395 drain_left.n232 drain_left.n231 104.615
R1396 drain_left.n231 drain_left.n163 104.615
R1397 drain_left.n224 drain_left.n163 104.615
R1398 drain_left.n224 drain_left.n223 104.615
R1399 drain_left.n223 drain_left.n167 104.615
R1400 drain_left.n216 drain_left.n167 104.615
R1401 drain_left.n216 drain_left.n215 104.615
R1402 drain_left.n215 drain_left.n171 104.615
R1403 drain_left.n208 drain_left.n171 104.615
R1404 drain_left.n208 drain_left.n207 104.615
R1405 drain_left.n207 drain_left.n206 104.615
R1406 drain_left.n206 drain_left.n175 104.615
R1407 drain_left.n199 drain_left.n175 104.615
R1408 drain_left.n199 drain_left.n198 104.615
R1409 drain_left.n198 drain_left.n180 104.615
R1410 drain_left.n191 drain_left.n180 104.615
R1411 drain_left.n191 drain_left.n190 104.615
R1412 drain_left.n190 drain_left.n184 104.615
R1413 drain_left drain_left.n138 85.8194
R1414 drain_left drain_left.n277 53.8533
R1415 drain_left.t1 drain_left.n43 52.3082
R1416 drain_left.t0 drain_left.n184 52.3082
R1417 drain_left.n69 drain_left.n34 13.1884
R1418 drain_left.n116 drain_left.n115 13.1884
R1419 drain_left.n255 drain_left.n254 13.1884
R1420 drain_left.n209 drain_left.n174 13.1884
R1421 drain_left.n65 drain_left.n64 12.8005
R1422 drain_left.n70 drain_left.n32 12.8005
R1423 drain_left.n114 drain_left.n12 12.8005
R1424 drain_left.n119 drain_left.n10 12.8005
R1425 drain_left.n258 drain_left.n149 12.8005
R1426 drain_left.n253 drain_left.n151 12.8005
R1427 drain_left.n210 drain_left.n172 12.8005
R1428 drain_left.n205 drain_left.n176 12.8005
R1429 drain_left.n63 drain_left.n36 12.0247
R1430 drain_left.n74 drain_left.n73 12.0247
R1431 drain_left.n111 drain_left.n110 12.0247
R1432 drain_left.n120 drain_left.n8 12.0247
R1433 drain_left.n259 drain_left.n147 12.0247
R1434 drain_left.n250 drain_left.n249 12.0247
R1435 drain_left.n214 drain_left.n213 12.0247
R1436 drain_left.n204 drain_left.n177 12.0247
R1437 drain_left.n60 drain_left.n59 11.249
R1438 drain_left.n77 drain_left.n30 11.249
R1439 drain_left.n106 drain_left.n14 11.249
R1440 drain_left.n124 drain_left.n123 11.249
R1441 drain_left.n263 drain_left.n262 11.249
R1442 drain_left.n246 drain_left.n153 11.249
R1443 drain_left.n217 drain_left.n170 11.249
R1444 drain_left.n201 drain_left.n200 11.249
R1445 drain_left.n56 drain_left.n38 10.4732
R1446 drain_left.n78 drain_left.n28 10.4732
R1447 drain_left.n105 drain_left.n16 10.4732
R1448 drain_left.n127 drain_left.n6 10.4732
R1449 drain_left.n266 drain_left.n145 10.4732
R1450 drain_left.n245 drain_left.n156 10.4732
R1451 drain_left.n218 drain_left.n168 10.4732
R1452 drain_left.n197 drain_left.n179 10.4732
R1453 drain_left.n45 drain_left.n44 10.2747
R1454 drain_left.n186 drain_left.n185 10.2747
R1455 drain_left.n55 drain_left.n40 9.69747
R1456 drain_left.n82 drain_left.n81 9.69747
R1457 drain_left.n102 drain_left.n101 9.69747
R1458 drain_left.n128 drain_left.n4 9.69747
R1459 drain_left.n267 drain_left.n143 9.69747
R1460 drain_left.n242 drain_left.n241 9.69747
R1461 drain_left.n222 drain_left.n221 9.69747
R1462 drain_left.n196 drain_left.n181 9.69747
R1463 drain_left.n138 drain_left.n137 9.45567
R1464 drain_left.n277 drain_left.n276 9.45567
R1465 drain_left.n2 drain_left.n1 9.3005
R1466 drain_left.n131 drain_left.n130 9.3005
R1467 drain_left.n129 drain_left.n128 9.3005
R1468 drain_left.n6 drain_left.n5 9.3005
R1469 drain_left.n123 drain_left.n122 9.3005
R1470 drain_left.n121 drain_left.n120 9.3005
R1471 drain_left.n10 drain_left.n9 9.3005
R1472 drain_left.n89 drain_left.n88 9.3005
R1473 drain_left.n87 drain_left.n86 9.3005
R1474 drain_left.n26 drain_left.n25 9.3005
R1475 drain_left.n81 drain_left.n80 9.3005
R1476 drain_left.n79 drain_left.n78 9.3005
R1477 drain_left.n30 drain_left.n29 9.3005
R1478 drain_left.n73 drain_left.n72 9.3005
R1479 drain_left.n71 drain_left.n70 9.3005
R1480 drain_left.n47 drain_left.n46 9.3005
R1481 drain_left.n42 drain_left.n41 9.3005
R1482 drain_left.n53 drain_left.n52 9.3005
R1483 drain_left.n55 drain_left.n54 9.3005
R1484 drain_left.n38 drain_left.n37 9.3005
R1485 drain_left.n61 drain_left.n60 9.3005
R1486 drain_left.n63 drain_left.n62 9.3005
R1487 drain_left.n64 drain_left.n33 9.3005
R1488 drain_left.n22 drain_left.n21 9.3005
R1489 drain_left.n95 drain_left.n94 9.3005
R1490 drain_left.n97 drain_left.n96 9.3005
R1491 drain_left.n18 drain_left.n17 9.3005
R1492 drain_left.n103 drain_left.n102 9.3005
R1493 drain_left.n105 drain_left.n104 9.3005
R1494 drain_left.n14 drain_left.n13 9.3005
R1495 drain_left.n112 drain_left.n111 9.3005
R1496 drain_left.n114 drain_left.n113 9.3005
R1497 drain_left.n137 drain_left.n136 9.3005
R1498 drain_left.n188 drain_left.n187 9.3005
R1499 drain_left.n183 drain_left.n182 9.3005
R1500 drain_left.n194 drain_left.n193 9.3005
R1501 drain_left.n196 drain_left.n195 9.3005
R1502 drain_left.n179 drain_left.n178 9.3005
R1503 drain_left.n202 drain_left.n201 9.3005
R1504 drain_left.n204 drain_left.n203 9.3005
R1505 drain_left.n176 drain_left.n173 9.3005
R1506 drain_left.n235 drain_left.n234 9.3005
R1507 drain_left.n237 drain_left.n236 9.3005
R1508 drain_left.n158 drain_left.n157 9.3005
R1509 drain_left.n243 drain_left.n242 9.3005
R1510 drain_left.n245 drain_left.n244 9.3005
R1511 drain_left.n153 drain_left.n152 9.3005
R1512 drain_left.n251 drain_left.n250 9.3005
R1513 drain_left.n253 drain_left.n252 9.3005
R1514 drain_left.n276 drain_left.n275 9.3005
R1515 drain_left.n141 drain_left.n140 9.3005
R1516 drain_left.n270 drain_left.n269 9.3005
R1517 drain_left.n268 drain_left.n267 9.3005
R1518 drain_left.n145 drain_left.n144 9.3005
R1519 drain_left.n262 drain_left.n261 9.3005
R1520 drain_left.n260 drain_left.n259 9.3005
R1521 drain_left.n149 drain_left.n148 9.3005
R1522 drain_left.n162 drain_left.n161 9.3005
R1523 drain_left.n229 drain_left.n228 9.3005
R1524 drain_left.n227 drain_left.n226 9.3005
R1525 drain_left.n166 drain_left.n165 9.3005
R1526 drain_left.n221 drain_left.n220 9.3005
R1527 drain_left.n219 drain_left.n218 9.3005
R1528 drain_left.n170 drain_left.n169 9.3005
R1529 drain_left.n213 drain_left.n212 9.3005
R1530 drain_left.n211 drain_left.n210 9.3005
R1531 drain_left.n52 drain_left.n51 8.92171
R1532 drain_left.n85 drain_left.n26 8.92171
R1533 drain_left.n98 drain_left.n18 8.92171
R1534 drain_left.n132 drain_left.n131 8.92171
R1535 drain_left.n271 drain_left.n270 8.92171
R1536 drain_left.n238 drain_left.n158 8.92171
R1537 drain_left.n225 drain_left.n166 8.92171
R1538 drain_left.n193 drain_left.n192 8.92171
R1539 drain_left.n48 drain_left.n42 8.14595
R1540 drain_left.n86 drain_left.n24 8.14595
R1541 drain_left.n97 drain_left.n20 8.14595
R1542 drain_left.n135 drain_left.n2 8.14595
R1543 drain_left.n274 drain_left.n141 8.14595
R1544 drain_left.n237 drain_left.n160 8.14595
R1545 drain_left.n226 drain_left.n164 8.14595
R1546 drain_left.n189 drain_left.n183 8.14595
R1547 drain_left.n47 drain_left.n44 7.3702
R1548 drain_left.n90 drain_left.n89 7.3702
R1549 drain_left.n94 drain_left.n93 7.3702
R1550 drain_left.n136 drain_left.n0 7.3702
R1551 drain_left.n275 drain_left.n139 7.3702
R1552 drain_left.n234 drain_left.n233 7.3702
R1553 drain_left.n230 drain_left.n229 7.3702
R1554 drain_left.n188 drain_left.n185 7.3702
R1555 drain_left.n90 drain_left.n22 6.59444
R1556 drain_left.n93 drain_left.n22 6.59444
R1557 drain_left.n138 drain_left.n0 6.59444
R1558 drain_left.n277 drain_left.n139 6.59444
R1559 drain_left.n233 drain_left.n162 6.59444
R1560 drain_left.n230 drain_left.n162 6.59444
R1561 drain_left.n48 drain_left.n47 5.81868
R1562 drain_left.n89 drain_left.n24 5.81868
R1563 drain_left.n94 drain_left.n20 5.81868
R1564 drain_left.n136 drain_left.n135 5.81868
R1565 drain_left.n275 drain_left.n274 5.81868
R1566 drain_left.n234 drain_left.n160 5.81868
R1567 drain_left.n229 drain_left.n164 5.81868
R1568 drain_left.n189 drain_left.n188 5.81868
R1569 drain_left.n51 drain_left.n42 5.04292
R1570 drain_left.n86 drain_left.n85 5.04292
R1571 drain_left.n98 drain_left.n97 5.04292
R1572 drain_left.n132 drain_left.n2 5.04292
R1573 drain_left.n271 drain_left.n141 5.04292
R1574 drain_left.n238 drain_left.n237 5.04292
R1575 drain_left.n226 drain_left.n225 5.04292
R1576 drain_left.n192 drain_left.n183 5.04292
R1577 drain_left.n52 drain_left.n40 4.26717
R1578 drain_left.n82 drain_left.n26 4.26717
R1579 drain_left.n101 drain_left.n18 4.26717
R1580 drain_left.n131 drain_left.n4 4.26717
R1581 drain_left.n270 drain_left.n143 4.26717
R1582 drain_left.n241 drain_left.n158 4.26717
R1583 drain_left.n222 drain_left.n166 4.26717
R1584 drain_left.n193 drain_left.n181 4.26717
R1585 drain_left.n56 drain_left.n55 3.49141
R1586 drain_left.n81 drain_left.n28 3.49141
R1587 drain_left.n102 drain_left.n16 3.49141
R1588 drain_left.n128 drain_left.n127 3.49141
R1589 drain_left.n267 drain_left.n266 3.49141
R1590 drain_left.n242 drain_left.n156 3.49141
R1591 drain_left.n221 drain_left.n168 3.49141
R1592 drain_left.n197 drain_left.n196 3.49141
R1593 drain_left.n187 drain_left.n186 2.84303
R1594 drain_left.n46 drain_left.n45 2.84303
R1595 drain_left.n59 drain_left.n38 2.71565
R1596 drain_left.n78 drain_left.n77 2.71565
R1597 drain_left.n106 drain_left.n105 2.71565
R1598 drain_left.n124 drain_left.n6 2.71565
R1599 drain_left.n263 drain_left.n145 2.71565
R1600 drain_left.n246 drain_left.n245 2.71565
R1601 drain_left.n218 drain_left.n217 2.71565
R1602 drain_left.n200 drain_left.n179 2.71565
R1603 drain_left.n60 drain_left.n36 1.93989
R1604 drain_left.n74 drain_left.n30 1.93989
R1605 drain_left.n110 drain_left.n14 1.93989
R1606 drain_left.n123 drain_left.n8 1.93989
R1607 drain_left.n262 drain_left.n147 1.93989
R1608 drain_left.n249 drain_left.n153 1.93989
R1609 drain_left.n214 drain_left.n170 1.93989
R1610 drain_left.n201 drain_left.n177 1.93989
R1611 drain_left.n65 drain_left.n63 1.16414
R1612 drain_left.n73 drain_left.n32 1.16414
R1613 drain_left.n111 drain_left.n12 1.16414
R1614 drain_left.n120 drain_left.n119 1.16414
R1615 drain_left.n259 drain_left.n258 1.16414
R1616 drain_left.n250 drain_left.n151 1.16414
R1617 drain_left.n213 drain_left.n172 1.16414
R1618 drain_left.n205 drain_left.n204 1.16414
R1619 drain_left.n64 drain_left.n34 0.388379
R1620 drain_left.n70 drain_left.n69 0.388379
R1621 drain_left.n115 drain_left.n114 0.388379
R1622 drain_left.n116 drain_left.n10 0.388379
R1623 drain_left.n255 drain_left.n149 0.388379
R1624 drain_left.n254 drain_left.n253 0.388379
R1625 drain_left.n210 drain_left.n209 0.388379
R1626 drain_left.n176 drain_left.n174 0.388379
R1627 drain_left.n46 drain_left.n41 0.155672
R1628 drain_left.n53 drain_left.n41 0.155672
R1629 drain_left.n54 drain_left.n53 0.155672
R1630 drain_left.n54 drain_left.n37 0.155672
R1631 drain_left.n61 drain_left.n37 0.155672
R1632 drain_left.n62 drain_left.n61 0.155672
R1633 drain_left.n62 drain_left.n33 0.155672
R1634 drain_left.n71 drain_left.n33 0.155672
R1635 drain_left.n72 drain_left.n71 0.155672
R1636 drain_left.n72 drain_left.n29 0.155672
R1637 drain_left.n79 drain_left.n29 0.155672
R1638 drain_left.n80 drain_left.n79 0.155672
R1639 drain_left.n80 drain_left.n25 0.155672
R1640 drain_left.n87 drain_left.n25 0.155672
R1641 drain_left.n88 drain_left.n87 0.155672
R1642 drain_left.n88 drain_left.n21 0.155672
R1643 drain_left.n95 drain_left.n21 0.155672
R1644 drain_left.n96 drain_left.n95 0.155672
R1645 drain_left.n96 drain_left.n17 0.155672
R1646 drain_left.n103 drain_left.n17 0.155672
R1647 drain_left.n104 drain_left.n103 0.155672
R1648 drain_left.n104 drain_left.n13 0.155672
R1649 drain_left.n112 drain_left.n13 0.155672
R1650 drain_left.n113 drain_left.n112 0.155672
R1651 drain_left.n113 drain_left.n9 0.155672
R1652 drain_left.n121 drain_left.n9 0.155672
R1653 drain_left.n122 drain_left.n121 0.155672
R1654 drain_left.n122 drain_left.n5 0.155672
R1655 drain_left.n129 drain_left.n5 0.155672
R1656 drain_left.n130 drain_left.n129 0.155672
R1657 drain_left.n130 drain_left.n1 0.155672
R1658 drain_left.n137 drain_left.n1 0.155672
R1659 drain_left.n276 drain_left.n140 0.155672
R1660 drain_left.n269 drain_left.n140 0.155672
R1661 drain_left.n269 drain_left.n268 0.155672
R1662 drain_left.n268 drain_left.n144 0.155672
R1663 drain_left.n261 drain_left.n144 0.155672
R1664 drain_left.n261 drain_left.n260 0.155672
R1665 drain_left.n260 drain_left.n148 0.155672
R1666 drain_left.n252 drain_left.n148 0.155672
R1667 drain_left.n252 drain_left.n251 0.155672
R1668 drain_left.n251 drain_left.n152 0.155672
R1669 drain_left.n244 drain_left.n152 0.155672
R1670 drain_left.n244 drain_left.n243 0.155672
R1671 drain_left.n243 drain_left.n157 0.155672
R1672 drain_left.n236 drain_left.n157 0.155672
R1673 drain_left.n236 drain_left.n235 0.155672
R1674 drain_left.n235 drain_left.n161 0.155672
R1675 drain_left.n228 drain_left.n161 0.155672
R1676 drain_left.n228 drain_left.n227 0.155672
R1677 drain_left.n227 drain_left.n165 0.155672
R1678 drain_left.n220 drain_left.n165 0.155672
R1679 drain_left.n220 drain_left.n219 0.155672
R1680 drain_left.n219 drain_left.n169 0.155672
R1681 drain_left.n212 drain_left.n169 0.155672
R1682 drain_left.n212 drain_left.n211 0.155672
R1683 drain_left.n211 drain_left.n173 0.155672
R1684 drain_left.n203 drain_left.n173 0.155672
R1685 drain_left.n203 drain_left.n202 0.155672
R1686 drain_left.n202 drain_left.n178 0.155672
R1687 drain_left.n195 drain_left.n178 0.155672
R1688 drain_left.n195 drain_left.n194 0.155672
R1689 drain_left.n194 drain_left.n182 0.155672
R1690 drain_left.n187 drain_left.n182 0.155672
C0 drain_right minus 3.91523f
C1 source drain_left 10.7091f
C2 plus drain_left 4.01485f
C3 drain_right drain_left 0.465826f
C4 minus drain_left 0.171858f
C5 source plus 2.82323f
C6 drain_right source 10.693f
C7 drain_right plus 0.262954f
C8 source minus 2.80815f
C9 minus plus 6.94959f
C10 drain_right a_n1128_n5892# 10.012061f
C11 drain_left a_n1128_n5892# 10.177171f
C12 source a_n1128_n5892# 11.453456f
C13 minus a_n1128_n5892# 5.025655f
C14 plus a_n1128_n5892# 12.54853f
C15 drain_left.n0 a_n1128_n5892# 0.028337f
C16 drain_left.n1 a_n1128_n5892# 0.020555f
C17 drain_left.n2 a_n1128_n5892# 0.011045f
C18 drain_left.n3 a_n1128_n5892# 0.026107f
C19 drain_left.n4 a_n1128_n5892# 0.011695f
C20 drain_left.n5 a_n1128_n5892# 0.020555f
C21 drain_left.n6 a_n1128_n5892# 0.011045f
C22 drain_left.n7 a_n1128_n5892# 0.026107f
C23 drain_left.n8 a_n1128_n5892# 0.011695f
C24 drain_left.n9 a_n1128_n5892# 0.020555f
C25 drain_left.n10 a_n1128_n5892# 0.011045f
C26 drain_left.n11 a_n1128_n5892# 0.026107f
C27 drain_left.n12 a_n1128_n5892# 0.011695f
C28 drain_left.n13 a_n1128_n5892# 0.020555f
C29 drain_left.n14 a_n1128_n5892# 0.011045f
C30 drain_left.n15 a_n1128_n5892# 0.026107f
C31 drain_left.n16 a_n1128_n5892# 0.011695f
C32 drain_left.n17 a_n1128_n5892# 0.020555f
C33 drain_left.n18 a_n1128_n5892# 0.011045f
C34 drain_left.n19 a_n1128_n5892# 0.026107f
C35 drain_left.n20 a_n1128_n5892# 0.011695f
C36 drain_left.n21 a_n1128_n5892# 0.020555f
C37 drain_left.n22 a_n1128_n5892# 0.011045f
C38 drain_left.n23 a_n1128_n5892# 0.026107f
C39 drain_left.n24 a_n1128_n5892# 0.011695f
C40 drain_left.n25 a_n1128_n5892# 0.020555f
C41 drain_left.n26 a_n1128_n5892# 0.011045f
C42 drain_left.n27 a_n1128_n5892# 0.026107f
C43 drain_left.n28 a_n1128_n5892# 0.011695f
C44 drain_left.n29 a_n1128_n5892# 0.020555f
C45 drain_left.n30 a_n1128_n5892# 0.011045f
C46 drain_left.n31 a_n1128_n5892# 0.026107f
C47 drain_left.n32 a_n1128_n5892# 0.011695f
C48 drain_left.n33 a_n1128_n5892# 0.020555f
C49 drain_left.n34 a_n1128_n5892# 0.01137f
C50 drain_left.n35 a_n1128_n5892# 0.026107f
C51 drain_left.n36 a_n1128_n5892# 0.011695f
C52 drain_left.n37 a_n1128_n5892# 0.020555f
C53 drain_left.n38 a_n1128_n5892# 0.011045f
C54 drain_left.n39 a_n1128_n5892# 0.026107f
C55 drain_left.n40 a_n1128_n5892# 0.011695f
C56 drain_left.n41 a_n1128_n5892# 0.020555f
C57 drain_left.n42 a_n1128_n5892# 0.011045f
C58 drain_left.n43 a_n1128_n5892# 0.01958f
C59 drain_left.n44 a_n1128_n5892# 0.018456f
C60 drain_left.t1 a_n1128_n5892# 0.045532f
C61 drain_left.n45 a_n1128_n5892# 0.250786f
C62 drain_left.n46 a_n1128_n5892# 2.22548f
C63 drain_left.n47 a_n1128_n5892# 0.011045f
C64 drain_left.n48 a_n1128_n5892# 0.011695f
C65 drain_left.n49 a_n1128_n5892# 0.026107f
C66 drain_left.n50 a_n1128_n5892# 0.026107f
C67 drain_left.n51 a_n1128_n5892# 0.011695f
C68 drain_left.n52 a_n1128_n5892# 0.011045f
C69 drain_left.n53 a_n1128_n5892# 0.020555f
C70 drain_left.n54 a_n1128_n5892# 0.020555f
C71 drain_left.n55 a_n1128_n5892# 0.011045f
C72 drain_left.n56 a_n1128_n5892# 0.011695f
C73 drain_left.n57 a_n1128_n5892# 0.026107f
C74 drain_left.n58 a_n1128_n5892# 0.026107f
C75 drain_left.n59 a_n1128_n5892# 0.011695f
C76 drain_left.n60 a_n1128_n5892# 0.011045f
C77 drain_left.n61 a_n1128_n5892# 0.020555f
C78 drain_left.n62 a_n1128_n5892# 0.020555f
C79 drain_left.n63 a_n1128_n5892# 0.011045f
C80 drain_left.n64 a_n1128_n5892# 0.011045f
C81 drain_left.n65 a_n1128_n5892# 0.011695f
C82 drain_left.n66 a_n1128_n5892# 0.026107f
C83 drain_left.n67 a_n1128_n5892# 0.026107f
C84 drain_left.n68 a_n1128_n5892# 0.026107f
C85 drain_left.n69 a_n1128_n5892# 0.01137f
C86 drain_left.n70 a_n1128_n5892# 0.011045f
C87 drain_left.n71 a_n1128_n5892# 0.020555f
C88 drain_left.n72 a_n1128_n5892# 0.020555f
C89 drain_left.n73 a_n1128_n5892# 0.011045f
C90 drain_left.n74 a_n1128_n5892# 0.011695f
C91 drain_left.n75 a_n1128_n5892# 0.026107f
C92 drain_left.n76 a_n1128_n5892# 0.026107f
C93 drain_left.n77 a_n1128_n5892# 0.011695f
C94 drain_left.n78 a_n1128_n5892# 0.011045f
C95 drain_left.n79 a_n1128_n5892# 0.020555f
C96 drain_left.n80 a_n1128_n5892# 0.020555f
C97 drain_left.n81 a_n1128_n5892# 0.011045f
C98 drain_left.n82 a_n1128_n5892# 0.011695f
C99 drain_left.n83 a_n1128_n5892# 0.026107f
C100 drain_left.n84 a_n1128_n5892# 0.026107f
C101 drain_left.n85 a_n1128_n5892# 0.011695f
C102 drain_left.n86 a_n1128_n5892# 0.011045f
C103 drain_left.n87 a_n1128_n5892# 0.020555f
C104 drain_left.n88 a_n1128_n5892# 0.020555f
C105 drain_left.n89 a_n1128_n5892# 0.011045f
C106 drain_left.n90 a_n1128_n5892# 0.011695f
C107 drain_left.n91 a_n1128_n5892# 0.026107f
C108 drain_left.n92 a_n1128_n5892# 0.026107f
C109 drain_left.n93 a_n1128_n5892# 0.011695f
C110 drain_left.n94 a_n1128_n5892# 0.011045f
C111 drain_left.n95 a_n1128_n5892# 0.020555f
C112 drain_left.n96 a_n1128_n5892# 0.020555f
C113 drain_left.n97 a_n1128_n5892# 0.011045f
C114 drain_left.n98 a_n1128_n5892# 0.011695f
C115 drain_left.n99 a_n1128_n5892# 0.026107f
C116 drain_left.n100 a_n1128_n5892# 0.026107f
C117 drain_left.n101 a_n1128_n5892# 0.011695f
C118 drain_left.n102 a_n1128_n5892# 0.011045f
C119 drain_left.n103 a_n1128_n5892# 0.020555f
C120 drain_left.n104 a_n1128_n5892# 0.020555f
C121 drain_left.n105 a_n1128_n5892# 0.011045f
C122 drain_left.n106 a_n1128_n5892# 0.011695f
C123 drain_left.n107 a_n1128_n5892# 0.026107f
C124 drain_left.n108 a_n1128_n5892# 0.026107f
C125 drain_left.n109 a_n1128_n5892# 0.026107f
C126 drain_left.n110 a_n1128_n5892# 0.011695f
C127 drain_left.n111 a_n1128_n5892# 0.011045f
C128 drain_left.n112 a_n1128_n5892# 0.020555f
C129 drain_left.n113 a_n1128_n5892# 0.020555f
C130 drain_left.n114 a_n1128_n5892# 0.011045f
C131 drain_left.n115 a_n1128_n5892# 0.01137f
C132 drain_left.n116 a_n1128_n5892# 0.01137f
C133 drain_left.n117 a_n1128_n5892# 0.026107f
C134 drain_left.n118 a_n1128_n5892# 0.026107f
C135 drain_left.n119 a_n1128_n5892# 0.011695f
C136 drain_left.n120 a_n1128_n5892# 0.011045f
C137 drain_left.n121 a_n1128_n5892# 0.020555f
C138 drain_left.n122 a_n1128_n5892# 0.020555f
C139 drain_left.n123 a_n1128_n5892# 0.011045f
C140 drain_left.n124 a_n1128_n5892# 0.011695f
C141 drain_left.n125 a_n1128_n5892# 0.026107f
C142 drain_left.n126 a_n1128_n5892# 0.026107f
C143 drain_left.n127 a_n1128_n5892# 0.011695f
C144 drain_left.n128 a_n1128_n5892# 0.011045f
C145 drain_left.n129 a_n1128_n5892# 0.020555f
C146 drain_left.n130 a_n1128_n5892# 0.020555f
C147 drain_left.n131 a_n1128_n5892# 0.011045f
C148 drain_left.n132 a_n1128_n5892# 0.011695f
C149 drain_left.n133 a_n1128_n5892# 0.026107f
C150 drain_left.n134 a_n1128_n5892# 0.055536f
C151 drain_left.n135 a_n1128_n5892# 0.011695f
C152 drain_left.n136 a_n1128_n5892# 0.011045f
C153 drain_left.n137 a_n1128_n5892# 0.045265f
C154 drain_left.n138 a_n1128_n5892# 0.733035f
C155 drain_left.n139 a_n1128_n5892# 0.028337f
C156 drain_left.n140 a_n1128_n5892# 0.020555f
C157 drain_left.n141 a_n1128_n5892# 0.011045f
C158 drain_left.n142 a_n1128_n5892# 0.026107f
C159 drain_left.n143 a_n1128_n5892# 0.011695f
C160 drain_left.n144 a_n1128_n5892# 0.020555f
C161 drain_left.n145 a_n1128_n5892# 0.011045f
C162 drain_left.n146 a_n1128_n5892# 0.026107f
C163 drain_left.n147 a_n1128_n5892# 0.011695f
C164 drain_left.n148 a_n1128_n5892# 0.020555f
C165 drain_left.n149 a_n1128_n5892# 0.011045f
C166 drain_left.n150 a_n1128_n5892# 0.026107f
C167 drain_left.n151 a_n1128_n5892# 0.011695f
C168 drain_left.n152 a_n1128_n5892# 0.020555f
C169 drain_left.n153 a_n1128_n5892# 0.011045f
C170 drain_left.n154 a_n1128_n5892# 0.026107f
C171 drain_left.n155 a_n1128_n5892# 0.026107f
C172 drain_left.n156 a_n1128_n5892# 0.011695f
C173 drain_left.n157 a_n1128_n5892# 0.020555f
C174 drain_left.n158 a_n1128_n5892# 0.011045f
C175 drain_left.n159 a_n1128_n5892# 0.026107f
C176 drain_left.n160 a_n1128_n5892# 0.011695f
C177 drain_left.n161 a_n1128_n5892# 0.020555f
C178 drain_left.n162 a_n1128_n5892# 0.011045f
C179 drain_left.n163 a_n1128_n5892# 0.026107f
C180 drain_left.n164 a_n1128_n5892# 0.011695f
C181 drain_left.n165 a_n1128_n5892# 0.020555f
C182 drain_left.n166 a_n1128_n5892# 0.011045f
C183 drain_left.n167 a_n1128_n5892# 0.026107f
C184 drain_left.n168 a_n1128_n5892# 0.011695f
C185 drain_left.n169 a_n1128_n5892# 0.020555f
C186 drain_left.n170 a_n1128_n5892# 0.011045f
C187 drain_left.n171 a_n1128_n5892# 0.026107f
C188 drain_left.n172 a_n1128_n5892# 0.011695f
C189 drain_left.n173 a_n1128_n5892# 0.020555f
C190 drain_left.n174 a_n1128_n5892# 0.01137f
C191 drain_left.n175 a_n1128_n5892# 0.026107f
C192 drain_left.n176 a_n1128_n5892# 0.011045f
C193 drain_left.n177 a_n1128_n5892# 0.011695f
C194 drain_left.n178 a_n1128_n5892# 0.020555f
C195 drain_left.n179 a_n1128_n5892# 0.011045f
C196 drain_left.n180 a_n1128_n5892# 0.026107f
C197 drain_left.n181 a_n1128_n5892# 0.011695f
C198 drain_left.n182 a_n1128_n5892# 0.020555f
C199 drain_left.n183 a_n1128_n5892# 0.011045f
C200 drain_left.n184 a_n1128_n5892# 0.01958f
C201 drain_left.n185 a_n1128_n5892# 0.018456f
C202 drain_left.t0 a_n1128_n5892# 0.045532f
C203 drain_left.n186 a_n1128_n5892# 0.250786f
C204 drain_left.n187 a_n1128_n5892# 2.22548f
C205 drain_left.n188 a_n1128_n5892# 0.011045f
C206 drain_left.n189 a_n1128_n5892# 0.011695f
C207 drain_left.n190 a_n1128_n5892# 0.026107f
C208 drain_left.n191 a_n1128_n5892# 0.026107f
C209 drain_left.n192 a_n1128_n5892# 0.011695f
C210 drain_left.n193 a_n1128_n5892# 0.011045f
C211 drain_left.n194 a_n1128_n5892# 0.020555f
C212 drain_left.n195 a_n1128_n5892# 0.020555f
C213 drain_left.n196 a_n1128_n5892# 0.011045f
C214 drain_left.n197 a_n1128_n5892# 0.011695f
C215 drain_left.n198 a_n1128_n5892# 0.026107f
C216 drain_left.n199 a_n1128_n5892# 0.026107f
C217 drain_left.n200 a_n1128_n5892# 0.011695f
C218 drain_left.n201 a_n1128_n5892# 0.011045f
C219 drain_left.n202 a_n1128_n5892# 0.020555f
C220 drain_left.n203 a_n1128_n5892# 0.020555f
C221 drain_left.n204 a_n1128_n5892# 0.011045f
C222 drain_left.n205 a_n1128_n5892# 0.011695f
C223 drain_left.n206 a_n1128_n5892# 0.026107f
C224 drain_left.n207 a_n1128_n5892# 0.026107f
C225 drain_left.n208 a_n1128_n5892# 0.026107f
C226 drain_left.n209 a_n1128_n5892# 0.01137f
C227 drain_left.n210 a_n1128_n5892# 0.011045f
C228 drain_left.n211 a_n1128_n5892# 0.020555f
C229 drain_left.n212 a_n1128_n5892# 0.020555f
C230 drain_left.n213 a_n1128_n5892# 0.011045f
C231 drain_left.n214 a_n1128_n5892# 0.011695f
C232 drain_left.n215 a_n1128_n5892# 0.026107f
C233 drain_left.n216 a_n1128_n5892# 0.026107f
C234 drain_left.n217 a_n1128_n5892# 0.011695f
C235 drain_left.n218 a_n1128_n5892# 0.011045f
C236 drain_left.n219 a_n1128_n5892# 0.020555f
C237 drain_left.n220 a_n1128_n5892# 0.020555f
C238 drain_left.n221 a_n1128_n5892# 0.011045f
C239 drain_left.n222 a_n1128_n5892# 0.011695f
C240 drain_left.n223 a_n1128_n5892# 0.026107f
C241 drain_left.n224 a_n1128_n5892# 0.026107f
C242 drain_left.n225 a_n1128_n5892# 0.011695f
C243 drain_left.n226 a_n1128_n5892# 0.011045f
C244 drain_left.n227 a_n1128_n5892# 0.020555f
C245 drain_left.n228 a_n1128_n5892# 0.020555f
C246 drain_left.n229 a_n1128_n5892# 0.011045f
C247 drain_left.n230 a_n1128_n5892# 0.011695f
C248 drain_left.n231 a_n1128_n5892# 0.026107f
C249 drain_left.n232 a_n1128_n5892# 0.026107f
C250 drain_left.n233 a_n1128_n5892# 0.011695f
C251 drain_left.n234 a_n1128_n5892# 0.011045f
C252 drain_left.n235 a_n1128_n5892# 0.020555f
C253 drain_left.n236 a_n1128_n5892# 0.020555f
C254 drain_left.n237 a_n1128_n5892# 0.011045f
C255 drain_left.n238 a_n1128_n5892# 0.011695f
C256 drain_left.n239 a_n1128_n5892# 0.026107f
C257 drain_left.n240 a_n1128_n5892# 0.026107f
C258 drain_left.n241 a_n1128_n5892# 0.011695f
C259 drain_left.n242 a_n1128_n5892# 0.011045f
C260 drain_left.n243 a_n1128_n5892# 0.020555f
C261 drain_left.n244 a_n1128_n5892# 0.020555f
C262 drain_left.n245 a_n1128_n5892# 0.011045f
C263 drain_left.n246 a_n1128_n5892# 0.011695f
C264 drain_left.n247 a_n1128_n5892# 0.026107f
C265 drain_left.n248 a_n1128_n5892# 0.026107f
C266 drain_left.n249 a_n1128_n5892# 0.011695f
C267 drain_left.n250 a_n1128_n5892# 0.011045f
C268 drain_left.n251 a_n1128_n5892# 0.020555f
C269 drain_left.n252 a_n1128_n5892# 0.020555f
C270 drain_left.n253 a_n1128_n5892# 0.011045f
C271 drain_left.n254 a_n1128_n5892# 0.01137f
C272 drain_left.n255 a_n1128_n5892# 0.01137f
C273 drain_left.n256 a_n1128_n5892# 0.026107f
C274 drain_left.n257 a_n1128_n5892# 0.026107f
C275 drain_left.n258 a_n1128_n5892# 0.011695f
C276 drain_left.n259 a_n1128_n5892# 0.011045f
C277 drain_left.n260 a_n1128_n5892# 0.020555f
C278 drain_left.n261 a_n1128_n5892# 0.020555f
C279 drain_left.n262 a_n1128_n5892# 0.011045f
C280 drain_left.n263 a_n1128_n5892# 0.011695f
C281 drain_left.n264 a_n1128_n5892# 0.026107f
C282 drain_left.n265 a_n1128_n5892# 0.026107f
C283 drain_left.n266 a_n1128_n5892# 0.011695f
C284 drain_left.n267 a_n1128_n5892# 0.011045f
C285 drain_left.n268 a_n1128_n5892# 0.020555f
C286 drain_left.n269 a_n1128_n5892# 0.020555f
C287 drain_left.n270 a_n1128_n5892# 0.011045f
C288 drain_left.n271 a_n1128_n5892# 0.011695f
C289 drain_left.n272 a_n1128_n5892# 0.026107f
C290 drain_left.n273 a_n1128_n5892# 0.055536f
C291 drain_left.n274 a_n1128_n5892# 0.011695f
C292 drain_left.n275 a_n1128_n5892# 0.011045f
C293 drain_left.n276 a_n1128_n5892# 0.045265f
C294 drain_left.n277 a_n1128_n5892# 0.07899f
C295 plus.t1 a_n1128_n5892# 2.97969f
C296 plus.t0 a_n1128_n5892# 3.03328f
C297 drain_right.n0 a_n1128_n5892# 0.028299f
C298 drain_right.n1 a_n1128_n5892# 0.020527f
C299 drain_right.n2 a_n1128_n5892# 0.011031f
C300 drain_right.n3 a_n1128_n5892# 0.026072f
C301 drain_right.n4 a_n1128_n5892# 0.011679f
C302 drain_right.n5 a_n1128_n5892# 0.020527f
C303 drain_right.n6 a_n1128_n5892# 0.011031f
C304 drain_right.n7 a_n1128_n5892# 0.026072f
C305 drain_right.n8 a_n1128_n5892# 0.011679f
C306 drain_right.n9 a_n1128_n5892# 0.020527f
C307 drain_right.n10 a_n1128_n5892# 0.011031f
C308 drain_right.n11 a_n1128_n5892# 0.026072f
C309 drain_right.n12 a_n1128_n5892# 0.011679f
C310 drain_right.n13 a_n1128_n5892# 0.020527f
C311 drain_right.n14 a_n1128_n5892# 0.011031f
C312 drain_right.n15 a_n1128_n5892# 0.026072f
C313 drain_right.n16 a_n1128_n5892# 0.011679f
C314 drain_right.n17 a_n1128_n5892# 0.020527f
C315 drain_right.n18 a_n1128_n5892# 0.011031f
C316 drain_right.n19 a_n1128_n5892# 0.026072f
C317 drain_right.n20 a_n1128_n5892# 0.011679f
C318 drain_right.n21 a_n1128_n5892# 0.020527f
C319 drain_right.n22 a_n1128_n5892# 0.011031f
C320 drain_right.n23 a_n1128_n5892# 0.026072f
C321 drain_right.n24 a_n1128_n5892# 0.011679f
C322 drain_right.n25 a_n1128_n5892# 0.020527f
C323 drain_right.n26 a_n1128_n5892# 0.011031f
C324 drain_right.n27 a_n1128_n5892# 0.026072f
C325 drain_right.n28 a_n1128_n5892# 0.011679f
C326 drain_right.n29 a_n1128_n5892# 0.020527f
C327 drain_right.n30 a_n1128_n5892# 0.011031f
C328 drain_right.n31 a_n1128_n5892# 0.026072f
C329 drain_right.n32 a_n1128_n5892# 0.011679f
C330 drain_right.n33 a_n1128_n5892# 0.020527f
C331 drain_right.n34 a_n1128_n5892# 0.011355f
C332 drain_right.n35 a_n1128_n5892# 0.026072f
C333 drain_right.n36 a_n1128_n5892# 0.011679f
C334 drain_right.n37 a_n1128_n5892# 0.020527f
C335 drain_right.n38 a_n1128_n5892# 0.011031f
C336 drain_right.n39 a_n1128_n5892# 0.026072f
C337 drain_right.n40 a_n1128_n5892# 0.011679f
C338 drain_right.n41 a_n1128_n5892# 0.020527f
C339 drain_right.n42 a_n1128_n5892# 0.011031f
C340 drain_right.n43 a_n1128_n5892# 0.019554f
C341 drain_right.n44 a_n1128_n5892# 0.018431f
C342 drain_right.t0 a_n1128_n5892# 0.045471f
C343 drain_right.n45 a_n1128_n5892# 0.25045f
C344 drain_right.n46 a_n1128_n5892# 2.2225f
C345 drain_right.n47 a_n1128_n5892# 0.011031f
C346 drain_right.n48 a_n1128_n5892# 0.011679f
C347 drain_right.n49 a_n1128_n5892# 0.026072f
C348 drain_right.n50 a_n1128_n5892# 0.026072f
C349 drain_right.n51 a_n1128_n5892# 0.011679f
C350 drain_right.n52 a_n1128_n5892# 0.011031f
C351 drain_right.n53 a_n1128_n5892# 0.020527f
C352 drain_right.n54 a_n1128_n5892# 0.020527f
C353 drain_right.n55 a_n1128_n5892# 0.011031f
C354 drain_right.n56 a_n1128_n5892# 0.011679f
C355 drain_right.n57 a_n1128_n5892# 0.026072f
C356 drain_right.n58 a_n1128_n5892# 0.026072f
C357 drain_right.n59 a_n1128_n5892# 0.011679f
C358 drain_right.n60 a_n1128_n5892# 0.011031f
C359 drain_right.n61 a_n1128_n5892# 0.020527f
C360 drain_right.n62 a_n1128_n5892# 0.020527f
C361 drain_right.n63 a_n1128_n5892# 0.011031f
C362 drain_right.n64 a_n1128_n5892# 0.011031f
C363 drain_right.n65 a_n1128_n5892# 0.011679f
C364 drain_right.n66 a_n1128_n5892# 0.026072f
C365 drain_right.n67 a_n1128_n5892# 0.026072f
C366 drain_right.n68 a_n1128_n5892# 0.026072f
C367 drain_right.n69 a_n1128_n5892# 0.011355f
C368 drain_right.n70 a_n1128_n5892# 0.011031f
C369 drain_right.n71 a_n1128_n5892# 0.020527f
C370 drain_right.n72 a_n1128_n5892# 0.020527f
C371 drain_right.n73 a_n1128_n5892# 0.011031f
C372 drain_right.n74 a_n1128_n5892# 0.011679f
C373 drain_right.n75 a_n1128_n5892# 0.026072f
C374 drain_right.n76 a_n1128_n5892# 0.026072f
C375 drain_right.n77 a_n1128_n5892# 0.011679f
C376 drain_right.n78 a_n1128_n5892# 0.011031f
C377 drain_right.n79 a_n1128_n5892# 0.020527f
C378 drain_right.n80 a_n1128_n5892# 0.020527f
C379 drain_right.n81 a_n1128_n5892# 0.011031f
C380 drain_right.n82 a_n1128_n5892# 0.011679f
C381 drain_right.n83 a_n1128_n5892# 0.026072f
C382 drain_right.n84 a_n1128_n5892# 0.026072f
C383 drain_right.n85 a_n1128_n5892# 0.011679f
C384 drain_right.n86 a_n1128_n5892# 0.011031f
C385 drain_right.n87 a_n1128_n5892# 0.020527f
C386 drain_right.n88 a_n1128_n5892# 0.020527f
C387 drain_right.n89 a_n1128_n5892# 0.011031f
C388 drain_right.n90 a_n1128_n5892# 0.011679f
C389 drain_right.n91 a_n1128_n5892# 0.026072f
C390 drain_right.n92 a_n1128_n5892# 0.026072f
C391 drain_right.n93 a_n1128_n5892# 0.011679f
C392 drain_right.n94 a_n1128_n5892# 0.011031f
C393 drain_right.n95 a_n1128_n5892# 0.020527f
C394 drain_right.n96 a_n1128_n5892# 0.020527f
C395 drain_right.n97 a_n1128_n5892# 0.011031f
C396 drain_right.n98 a_n1128_n5892# 0.011679f
C397 drain_right.n99 a_n1128_n5892# 0.026072f
C398 drain_right.n100 a_n1128_n5892# 0.026072f
C399 drain_right.n101 a_n1128_n5892# 0.011679f
C400 drain_right.n102 a_n1128_n5892# 0.011031f
C401 drain_right.n103 a_n1128_n5892# 0.020527f
C402 drain_right.n104 a_n1128_n5892# 0.020527f
C403 drain_right.n105 a_n1128_n5892# 0.011031f
C404 drain_right.n106 a_n1128_n5892# 0.011679f
C405 drain_right.n107 a_n1128_n5892# 0.026072f
C406 drain_right.n108 a_n1128_n5892# 0.026072f
C407 drain_right.n109 a_n1128_n5892# 0.026072f
C408 drain_right.n110 a_n1128_n5892# 0.011679f
C409 drain_right.n111 a_n1128_n5892# 0.011031f
C410 drain_right.n112 a_n1128_n5892# 0.020527f
C411 drain_right.n113 a_n1128_n5892# 0.020527f
C412 drain_right.n114 a_n1128_n5892# 0.011031f
C413 drain_right.n115 a_n1128_n5892# 0.011355f
C414 drain_right.n116 a_n1128_n5892# 0.011355f
C415 drain_right.n117 a_n1128_n5892# 0.026072f
C416 drain_right.n118 a_n1128_n5892# 0.026072f
C417 drain_right.n119 a_n1128_n5892# 0.011679f
C418 drain_right.n120 a_n1128_n5892# 0.011031f
C419 drain_right.n121 a_n1128_n5892# 0.020527f
C420 drain_right.n122 a_n1128_n5892# 0.020527f
C421 drain_right.n123 a_n1128_n5892# 0.011031f
C422 drain_right.n124 a_n1128_n5892# 0.011679f
C423 drain_right.n125 a_n1128_n5892# 0.026072f
C424 drain_right.n126 a_n1128_n5892# 0.026072f
C425 drain_right.n127 a_n1128_n5892# 0.011679f
C426 drain_right.n128 a_n1128_n5892# 0.011031f
C427 drain_right.n129 a_n1128_n5892# 0.020527f
C428 drain_right.n130 a_n1128_n5892# 0.020527f
C429 drain_right.n131 a_n1128_n5892# 0.011031f
C430 drain_right.n132 a_n1128_n5892# 0.011679f
C431 drain_right.n133 a_n1128_n5892# 0.026072f
C432 drain_right.n134 a_n1128_n5892# 0.055462f
C433 drain_right.n135 a_n1128_n5892# 0.011679f
C434 drain_right.n136 a_n1128_n5892# 0.011031f
C435 drain_right.n137 a_n1128_n5892# 0.045204f
C436 drain_right.n138 a_n1128_n5892# 0.707483f
C437 drain_right.n139 a_n1128_n5892# 0.028299f
C438 drain_right.n140 a_n1128_n5892# 0.020527f
C439 drain_right.n141 a_n1128_n5892# 0.011031f
C440 drain_right.n142 a_n1128_n5892# 0.026072f
C441 drain_right.n143 a_n1128_n5892# 0.011679f
C442 drain_right.n144 a_n1128_n5892# 0.020527f
C443 drain_right.n145 a_n1128_n5892# 0.011031f
C444 drain_right.n146 a_n1128_n5892# 0.026072f
C445 drain_right.n147 a_n1128_n5892# 0.011679f
C446 drain_right.n148 a_n1128_n5892# 0.020527f
C447 drain_right.n149 a_n1128_n5892# 0.011031f
C448 drain_right.n150 a_n1128_n5892# 0.026072f
C449 drain_right.n151 a_n1128_n5892# 0.011679f
C450 drain_right.n152 a_n1128_n5892# 0.020527f
C451 drain_right.n153 a_n1128_n5892# 0.011031f
C452 drain_right.n154 a_n1128_n5892# 0.026072f
C453 drain_right.n155 a_n1128_n5892# 0.026072f
C454 drain_right.n156 a_n1128_n5892# 0.011679f
C455 drain_right.n157 a_n1128_n5892# 0.020527f
C456 drain_right.n158 a_n1128_n5892# 0.011031f
C457 drain_right.n159 a_n1128_n5892# 0.026072f
C458 drain_right.n160 a_n1128_n5892# 0.011679f
C459 drain_right.n161 a_n1128_n5892# 0.020527f
C460 drain_right.n162 a_n1128_n5892# 0.011031f
C461 drain_right.n163 a_n1128_n5892# 0.026072f
C462 drain_right.n164 a_n1128_n5892# 0.011679f
C463 drain_right.n165 a_n1128_n5892# 0.020527f
C464 drain_right.n166 a_n1128_n5892# 0.011031f
C465 drain_right.n167 a_n1128_n5892# 0.026072f
C466 drain_right.n168 a_n1128_n5892# 0.011679f
C467 drain_right.n169 a_n1128_n5892# 0.020527f
C468 drain_right.n170 a_n1128_n5892# 0.011031f
C469 drain_right.n171 a_n1128_n5892# 0.026072f
C470 drain_right.n172 a_n1128_n5892# 0.011679f
C471 drain_right.n173 a_n1128_n5892# 0.020527f
C472 drain_right.n174 a_n1128_n5892# 0.011355f
C473 drain_right.n175 a_n1128_n5892# 0.026072f
C474 drain_right.n176 a_n1128_n5892# 0.011031f
C475 drain_right.n177 a_n1128_n5892# 0.011679f
C476 drain_right.n178 a_n1128_n5892# 0.020527f
C477 drain_right.n179 a_n1128_n5892# 0.011031f
C478 drain_right.n180 a_n1128_n5892# 0.026072f
C479 drain_right.n181 a_n1128_n5892# 0.011679f
C480 drain_right.n182 a_n1128_n5892# 0.020527f
C481 drain_right.n183 a_n1128_n5892# 0.011031f
C482 drain_right.n184 a_n1128_n5892# 0.019554f
C483 drain_right.n185 a_n1128_n5892# 0.018431f
C484 drain_right.t1 a_n1128_n5892# 0.045471f
C485 drain_right.n186 a_n1128_n5892# 0.25045f
C486 drain_right.n187 a_n1128_n5892# 2.2225f
C487 drain_right.n188 a_n1128_n5892# 0.011031f
C488 drain_right.n189 a_n1128_n5892# 0.011679f
C489 drain_right.n190 a_n1128_n5892# 0.026072f
C490 drain_right.n191 a_n1128_n5892# 0.026072f
C491 drain_right.n192 a_n1128_n5892# 0.011679f
C492 drain_right.n193 a_n1128_n5892# 0.011031f
C493 drain_right.n194 a_n1128_n5892# 0.020527f
C494 drain_right.n195 a_n1128_n5892# 0.020527f
C495 drain_right.n196 a_n1128_n5892# 0.011031f
C496 drain_right.n197 a_n1128_n5892# 0.011679f
C497 drain_right.n198 a_n1128_n5892# 0.026072f
C498 drain_right.n199 a_n1128_n5892# 0.026072f
C499 drain_right.n200 a_n1128_n5892# 0.011679f
C500 drain_right.n201 a_n1128_n5892# 0.011031f
C501 drain_right.n202 a_n1128_n5892# 0.020527f
C502 drain_right.n203 a_n1128_n5892# 0.020527f
C503 drain_right.n204 a_n1128_n5892# 0.011031f
C504 drain_right.n205 a_n1128_n5892# 0.011679f
C505 drain_right.n206 a_n1128_n5892# 0.026072f
C506 drain_right.n207 a_n1128_n5892# 0.026072f
C507 drain_right.n208 a_n1128_n5892# 0.026072f
C508 drain_right.n209 a_n1128_n5892# 0.011355f
C509 drain_right.n210 a_n1128_n5892# 0.011031f
C510 drain_right.n211 a_n1128_n5892# 0.020527f
C511 drain_right.n212 a_n1128_n5892# 0.020527f
C512 drain_right.n213 a_n1128_n5892# 0.011031f
C513 drain_right.n214 a_n1128_n5892# 0.011679f
C514 drain_right.n215 a_n1128_n5892# 0.026072f
C515 drain_right.n216 a_n1128_n5892# 0.026072f
C516 drain_right.n217 a_n1128_n5892# 0.011679f
C517 drain_right.n218 a_n1128_n5892# 0.011031f
C518 drain_right.n219 a_n1128_n5892# 0.020527f
C519 drain_right.n220 a_n1128_n5892# 0.020527f
C520 drain_right.n221 a_n1128_n5892# 0.011031f
C521 drain_right.n222 a_n1128_n5892# 0.011679f
C522 drain_right.n223 a_n1128_n5892# 0.026072f
C523 drain_right.n224 a_n1128_n5892# 0.026072f
C524 drain_right.n225 a_n1128_n5892# 0.011679f
C525 drain_right.n226 a_n1128_n5892# 0.011031f
C526 drain_right.n227 a_n1128_n5892# 0.020527f
C527 drain_right.n228 a_n1128_n5892# 0.020527f
C528 drain_right.n229 a_n1128_n5892# 0.011031f
C529 drain_right.n230 a_n1128_n5892# 0.011679f
C530 drain_right.n231 a_n1128_n5892# 0.026072f
C531 drain_right.n232 a_n1128_n5892# 0.026072f
C532 drain_right.n233 a_n1128_n5892# 0.011679f
C533 drain_right.n234 a_n1128_n5892# 0.011031f
C534 drain_right.n235 a_n1128_n5892# 0.020527f
C535 drain_right.n236 a_n1128_n5892# 0.020527f
C536 drain_right.n237 a_n1128_n5892# 0.011031f
C537 drain_right.n238 a_n1128_n5892# 0.011679f
C538 drain_right.n239 a_n1128_n5892# 0.026072f
C539 drain_right.n240 a_n1128_n5892# 0.026072f
C540 drain_right.n241 a_n1128_n5892# 0.011679f
C541 drain_right.n242 a_n1128_n5892# 0.011031f
C542 drain_right.n243 a_n1128_n5892# 0.020527f
C543 drain_right.n244 a_n1128_n5892# 0.020527f
C544 drain_right.n245 a_n1128_n5892# 0.011031f
C545 drain_right.n246 a_n1128_n5892# 0.011679f
C546 drain_right.n247 a_n1128_n5892# 0.026072f
C547 drain_right.n248 a_n1128_n5892# 0.026072f
C548 drain_right.n249 a_n1128_n5892# 0.011679f
C549 drain_right.n250 a_n1128_n5892# 0.011031f
C550 drain_right.n251 a_n1128_n5892# 0.020527f
C551 drain_right.n252 a_n1128_n5892# 0.020527f
C552 drain_right.n253 a_n1128_n5892# 0.011031f
C553 drain_right.n254 a_n1128_n5892# 0.011355f
C554 drain_right.n255 a_n1128_n5892# 0.011355f
C555 drain_right.n256 a_n1128_n5892# 0.026072f
C556 drain_right.n257 a_n1128_n5892# 0.026072f
C557 drain_right.n258 a_n1128_n5892# 0.011679f
C558 drain_right.n259 a_n1128_n5892# 0.011031f
C559 drain_right.n260 a_n1128_n5892# 0.020527f
C560 drain_right.n261 a_n1128_n5892# 0.020527f
C561 drain_right.n262 a_n1128_n5892# 0.011031f
C562 drain_right.n263 a_n1128_n5892# 0.011679f
C563 drain_right.n264 a_n1128_n5892# 0.026072f
C564 drain_right.n265 a_n1128_n5892# 0.026072f
C565 drain_right.n266 a_n1128_n5892# 0.011679f
C566 drain_right.n267 a_n1128_n5892# 0.011031f
C567 drain_right.n268 a_n1128_n5892# 0.020527f
C568 drain_right.n269 a_n1128_n5892# 0.020527f
C569 drain_right.n270 a_n1128_n5892# 0.011031f
C570 drain_right.n271 a_n1128_n5892# 0.011679f
C571 drain_right.n272 a_n1128_n5892# 0.026072f
C572 drain_right.n273 a_n1128_n5892# 0.055462f
C573 drain_right.n274 a_n1128_n5892# 0.011679f
C574 drain_right.n275 a_n1128_n5892# 0.011031f
C575 drain_right.n276 a_n1128_n5892# 0.045204f
C576 drain_right.n277 a_n1128_n5892# 0.078603f
C577 source.n0 a_n1128_n5892# 0.027071f
C578 source.n1 a_n1128_n5892# 0.019637f
C579 source.n2 a_n1128_n5892# 0.010552f
C580 source.n3 a_n1128_n5892# 0.024941f
C581 source.n4 a_n1128_n5892# 0.011173f
C582 source.n5 a_n1128_n5892# 0.019637f
C583 source.n6 a_n1128_n5892# 0.010552f
C584 source.n7 a_n1128_n5892# 0.024941f
C585 source.n8 a_n1128_n5892# 0.011173f
C586 source.n9 a_n1128_n5892# 0.019637f
C587 source.n10 a_n1128_n5892# 0.010552f
C588 source.n11 a_n1128_n5892# 0.024941f
C589 source.n12 a_n1128_n5892# 0.011173f
C590 source.n13 a_n1128_n5892# 0.019637f
C591 source.n14 a_n1128_n5892# 0.010552f
C592 source.n15 a_n1128_n5892# 0.024941f
C593 source.n16 a_n1128_n5892# 0.024941f
C594 source.n17 a_n1128_n5892# 0.011173f
C595 source.n18 a_n1128_n5892# 0.019637f
C596 source.n19 a_n1128_n5892# 0.010552f
C597 source.n20 a_n1128_n5892# 0.024941f
C598 source.n21 a_n1128_n5892# 0.011173f
C599 source.n22 a_n1128_n5892# 0.019637f
C600 source.n23 a_n1128_n5892# 0.010552f
C601 source.n24 a_n1128_n5892# 0.024941f
C602 source.n25 a_n1128_n5892# 0.011173f
C603 source.n26 a_n1128_n5892# 0.019637f
C604 source.n27 a_n1128_n5892# 0.010552f
C605 source.n28 a_n1128_n5892# 0.024941f
C606 source.n29 a_n1128_n5892# 0.011173f
C607 source.n30 a_n1128_n5892# 0.019637f
C608 source.n31 a_n1128_n5892# 0.010552f
C609 source.n32 a_n1128_n5892# 0.024941f
C610 source.n33 a_n1128_n5892# 0.011173f
C611 source.n34 a_n1128_n5892# 0.019637f
C612 source.n35 a_n1128_n5892# 0.010862f
C613 source.n36 a_n1128_n5892# 0.024941f
C614 source.n37 a_n1128_n5892# 0.010552f
C615 source.n38 a_n1128_n5892# 0.011173f
C616 source.n39 a_n1128_n5892# 0.019637f
C617 source.n40 a_n1128_n5892# 0.010552f
C618 source.n41 a_n1128_n5892# 0.024941f
C619 source.n42 a_n1128_n5892# 0.011173f
C620 source.n43 a_n1128_n5892# 0.019637f
C621 source.n44 a_n1128_n5892# 0.010552f
C622 source.n45 a_n1128_n5892# 0.018706f
C623 source.n46 a_n1128_n5892# 0.017631f
C624 source.t0 a_n1128_n5892# 0.043499f
C625 source.n47 a_n1128_n5892# 0.239586f
C626 source.n48 a_n1128_n5892# 2.12609f
C627 source.n49 a_n1128_n5892# 0.010552f
C628 source.n50 a_n1128_n5892# 0.011173f
C629 source.n51 a_n1128_n5892# 0.024941f
C630 source.n52 a_n1128_n5892# 0.024941f
C631 source.n53 a_n1128_n5892# 0.011173f
C632 source.n54 a_n1128_n5892# 0.010552f
C633 source.n55 a_n1128_n5892# 0.019637f
C634 source.n56 a_n1128_n5892# 0.019637f
C635 source.n57 a_n1128_n5892# 0.010552f
C636 source.n58 a_n1128_n5892# 0.011173f
C637 source.n59 a_n1128_n5892# 0.024941f
C638 source.n60 a_n1128_n5892# 0.024941f
C639 source.n61 a_n1128_n5892# 0.011173f
C640 source.n62 a_n1128_n5892# 0.010552f
C641 source.n63 a_n1128_n5892# 0.019637f
C642 source.n64 a_n1128_n5892# 0.019637f
C643 source.n65 a_n1128_n5892# 0.010552f
C644 source.n66 a_n1128_n5892# 0.011173f
C645 source.n67 a_n1128_n5892# 0.024941f
C646 source.n68 a_n1128_n5892# 0.024941f
C647 source.n69 a_n1128_n5892# 0.024941f
C648 source.n70 a_n1128_n5892# 0.010862f
C649 source.n71 a_n1128_n5892# 0.010552f
C650 source.n72 a_n1128_n5892# 0.019637f
C651 source.n73 a_n1128_n5892# 0.019637f
C652 source.n74 a_n1128_n5892# 0.010552f
C653 source.n75 a_n1128_n5892# 0.011173f
C654 source.n76 a_n1128_n5892# 0.024941f
C655 source.n77 a_n1128_n5892# 0.024941f
C656 source.n78 a_n1128_n5892# 0.011173f
C657 source.n79 a_n1128_n5892# 0.010552f
C658 source.n80 a_n1128_n5892# 0.019637f
C659 source.n81 a_n1128_n5892# 0.019637f
C660 source.n82 a_n1128_n5892# 0.010552f
C661 source.n83 a_n1128_n5892# 0.011173f
C662 source.n84 a_n1128_n5892# 0.024941f
C663 source.n85 a_n1128_n5892# 0.024941f
C664 source.n86 a_n1128_n5892# 0.011173f
C665 source.n87 a_n1128_n5892# 0.010552f
C666 source.n88 a_n1128_n5892# 0.019637f
C667 source.n89 a_n1128_n5892# 0.019637f
C668 source.n90 a_n1128_n5892# 0.010552f
C669 source.n91 a_n1128_n5892# 0.011173f
C670 source.n92 a_n1128_n5892# 0.024941f
C671 source.n93 a_n1128_n5892# 0.024941f
C672 source.n94 a_n1128_n5892# 0.011173f
C673 source.n95 a_n1128_n5892# 0.010552f
C674 source.n96 a_n1128_n5892# 0.019637f
C675 source.n97 a_n1128_n5892# 0.019637f
C676 source.n98 a_n1128_n5892# 0.010552f
C677 source.n99 a_n1128_n5892# 0.011173f
C678 source.n100 a_n1128_n5892# 0.024941f
C679 source.n101 a_n1128_n5892# 0.024941f
C680 source.n102 a_n1128_n5892# 0.011173f
C681 source.n103 a_n1128_n5892# 0.010552f
C682 source.n104 a_n1128_n5892# 0.019637f
C683 source.n105 a_n1128_n5892# 0.019637f
C684 source.n106 a_n1128_n5892# 0.010552f
C685 source.n107 a_n1128_n5892# 0.011173f
C686 source.n108 a_n1128_n5892# 0.024941f
C687 source.n109 a_n1128_n5892# 0.024941f
C688 source.n110 a_n1128_n5892# 0.011173f
C689 source.n111 a_n1128_n5892# 0.010552f
C690 source.n112 a_n1128_n5892# 0.019637f
C691 source.n113 a_n1128_n5892# 0.019637f
C692 source.n114 a_n1128_n5892# 0.010552f
C693 source.n115 a_n1128_n5892# 0.010862f
C694 source.n116 a_n1128_n5892# 0.010862f
C695 source.n117 a_n1128_n5892# 0.024941f
C696 source.n118 a_n1128_n5892# 0.024941f
C697 source.n119 a_n1128_n5892# 0.011173f
C698 source.n120 a_n1128_n5892# 0.010552f
C699 source.n121 a_n1128_n5892# 0.019637f
C700 source.n122 a_n1128_n5892# 0.019637f
C701 source.n123 a_n1128_n5892# 0.010552f
C702 source.n124 a_n1128_n5892# 0.011173f
C703 source.n125 a_n1128_n5892# 0.024941f
C704 source.n126 a_n1128_n5892# 0.024941f
C705 source.n127 a_n1128_n5892# 0.011173f
C706 source.n128 a_n1128_n5892# 0.010552f
C707 source.n129 a_n1128_n5892# 0.019637f
C708 source.n130 a_n1128_n5892# 0.019637f
C709 source.n131 a_n1128_n5892# 0.010552f
C710 source.n132 a_n1128_n5892# 0.011173f
C711 source.n133 a_n1128_n5892# 0.024941f
C712 source.n134 a_n1128_n5892# 0.053056f
C713 source.n135 a_n1128_n5892# 0.011173f
C714 source.n136 a_n1128_n5892# 0.010552f
C715 source.n137 a_n1128_n5892# 0.043244f
C716 source.n138 a_n1128_n5892# 0.029523f
C717 source.n139 a_n1128_n5892# 1.57991f
C718 source.n140 a_n1128_n5892# 0.027071f
C719 source.n141 a_n1128_n5892# 0.019637f
C720 source.n142 a_n1128_n5892# 0.010552f
C721 source.n143 a_n1128_n5892# 0.024941f
C722 source.n144 a_n1128_n5892# 0.011173f
C723 source.n145 a_n1128_n5892# 0.019637f
C724 source.n146 a_n1128_n5892# 0.010552f
C725 source.n147 a_n1128_n5892# 0.024941f
C726 source.n148 a_n1128_n5892# 0.011173f
C727 source.n149 a_n1128_n5892# 0.019637f
C728 source.n150 a_n1128_n5892# 0.010552f
C729 source.n151 a_n1128_n5892# 0.024941f
C730 source.n152 a_n1128_n5892# 0.011173f
C731 source.n153 a_n1128_n5892# 0.019637f
C732 source.n154 a_n1128_n5892# 0.010552f
C733 source.n155 a_n1128_n5892# 0.024941f
C734 source.n156 a_n1128_n5892# 0.024941f
C735 source.n157 a_n1128_n5892# 0.011173f
C736 source.n158 a_n1128_n5892# 0.019637f
C737 source.n159 a_n1128_n5892# 0.010552f
C738 source.n160 a_n1128_n5892# 0.024941f
C739 source.n161 a_n1128_n5892# 0.011173f
C740 source.n162 a_n1128_n5892# 0.019637f
C741 source.n163 a_n1128_n5892# 0.010552f
C742 source.n164 a_n1128_n5892# 0.024941f
C743 source.n165 a_n1128_n5892# 0.011173f
C744 source.n166 a_n1128_n5892# 0.019637f
C745 source.n167 a_n1128_n5892# 0.010552f
C746 source.n168 a_n1128_n5892# 0.024941f
C747 source.n169 a_n1128_n5892# 0.011173f
C748 source.n170 a_n1128_n5892# 0.019637f
C749 source.n171 a_n1128_n5892# 0.010552f
C750 source.n172 a_n1128_n5892# 0.024941f
C751 source.n173 a_n1128_n5892# 0.011173f
C752 source.n174 a_n1128_n5892# 0.019637f
C753 source.n175 a_n1128_n5892# 0.010862f
C754 source.n176 a_n1128_n5892# 0.024941f
C755 source.n177 a_n1128_n5892# 0.010552f
C756 source.n178 a_n1128_n5892# 0.011173f
C757 source.n179 a_n1128_n5892# 0.019637f
C758 source.n180 a_n1128_n5892# 0.010552f
C759 source.n181 a_n1128_n5892# 0.024941f
C760 source.n182 a_n1128_n5892# 0.011173f
C761 source.n183 a_n1128_n5892# 0.019637f
C762 source.n184 a_n1128_n5892# 0.010552f
C763 source.n185 a_n1128_n5892# 0.018706f
C764 source.n186 a_n1128_n5892# 0.017631f
C765 source.t2 a_n1128_n5892# 0.043499f
C766 source.n187 a_n1128_n5892# 0.239586f
C767 source.n188 a_n1128_n5892# 2.12609f
C768 source.n189 a_n1128_n5892# 0.010552f
C769 source.n190 a_n1128_n5892# 0.011173f
C770 source.n191 a_n1128_n5892# 0.024941f
C771 source.n192 a_n1128_n5892# 0.024941f
C772 source.n193 a_n1128_n5892# 0.011173f
C773 source.n194 a_n1128_n5892# 0.010552f
C774 source.n195 a_n1128_n5892# 0.019637f
C775 source.n196 a_n1128_n5892# 0.019637f
C776 source.n197 a_n1128_n5892# 0.010552f
C777 source.n198 a_n1128_n5892# 0.011173f
C778 source.n199 a_n1128_n5892# 0.024941f
C779 source.n200 a_n1128_n5892# 0.024941f
C780 source.n201 a_n1128_n5892# 0.011173f
C781 source.n202 a_n1128_n5892# 0.010552f
C782 source.n203 a_n1128_n5892# 0.019637f
C783 source.n204 a_n1128_n5892# 0.019637f
C784 source.n205 a_n1128_n5892# 0.010552f
C785 source.n206 a_n1128_n5892# 0.011173f
C786 source.n207 a_n1128_n5892# 0.024941f
C787 source.n208 a_n1128_n5892# 0.024941f
C788 source.n209 a_n1128_n5892# 0.024941f
C789 source.n210 a_n1128_n5892# 0.010862f
C790 source.n211 a_n1128_n5892# 0.010552f
C791 source.n212 a_n1128_n5892# 0.019637f
C792 source.n213 a_n1128_n5892# 0.019637f
C793 source.n214 a_n1128_n5892# 0.010552f
C794 source.n215 a_n1128_n5892# 0.011173f
C795 source.n216 a_n1128_n5892# 0.024941f
C796 source.n217 a_n1128_n5892# 0.024941f
C797 source.n218 a_n1128_n5892# 0.011173f
C798 source.n219 a_n1128_n5892# 0.010552f
C799 source.n220 a_n1128_n5892# 0.019637f
C800 source.n221 a_n1128_n5892# 0.019637f
C801 source.n222 a_n1128_n5892# 0.010552f
C802 source.n223 a_n1128_n5892# 0.011173f
C803 source.n224 a_n1128_n5892# 0.024941f
C804 source.n225 a_n1128_n5892# 0.024941f
C805 source.n226 a_n1128_n5892# 0.011173f
C806 source.n227 a_n1128_n5892# 0.010552f
C807 source.n228 a_n1128_n5892# 0.019637f
C808 source.n229 a_n1128_n5892# 0.019637f
C809 source.n230 a_n1128_n5892# 0.010552f
C810 source.n231 a_n1128_n5892# 0.011173f
C811 source.n232 a_n1128_n5892# 0.024941f
C812 source.n233 a_n1128_n5892# 0.024941f
C813 source.n234 a_n1128_n5892# 0.011173f
C814 source.n235 a_n1128_n5892# 0.010552f
C815 source.n236 a_n1128_n5892# 0.019637f
C816 source.n237 a_n1128_n5892# 0.019637f
C817 source.n238 a_n1128_n5892# 0.010552f
C818 source.n239 a_n1128_n5892# 0.011173f
C819 source.n240 a_n1128_n5892# 0.024941f
C820 source.n241 a_n1128_n5892# 0.024941f
C821 source.n242 a_n1128_n5892# 0.011173f
C822 source.n243 a_n1128_n5892# 0.010552f
C823 source.n244 a_n1128_n5892# 0.019637f
C824 source.n245 a_n1128_n5892# 0.019637f
C825 source.n246 a_n1128_n5892# 0.010552f
C826 source.n247 a_n1128_n5892# 0.011173f
C827 source.n248 a_n1128_n5892# 0.024941f
C828 source.n249 a_n1128_n5892# 0.024941f
C829 source.n250 a_n1128_n5892# 0.011173f
C830 source.n251 a_n1128_n5892# 0.010552f
C831 source.n252 a_n1128_n5892# 0.019637f
C832 source.n253 a_n1128_n5892# 0.019637f
C833 source.n254 a_n1128_n5892# 0.010552f
C834 source.n255 a_n1128_n5892# 0.010862f
C835 source.n256 a_n1128_n5892# 0.010862f
C836 source.n257 a_n1128_n5892# 0.024941f
C837 source.n258 a_n1128_n5892# 0.024941f
C838 source.n259 a_n1128_n5892# 0.011173f
C839 source.n260 a_n1128_n5892# 0.010552f
C840 source.n261 a_n1128_n5892# 0.019637f
C841 source.n262 a_n1128_n5892# 0.019637f
C842 source.n263 a_n1128_n5892# 0.010552f
C843 source.n264 a_n1128_n5892# 0.011173f
C844 source.n265 a_n1128_n5892# 0.024941f
C845 source.n266 a_n1128_n5892# 0.024941f
C846 source.n267 a_n1128_n5892# 0.011173f
C847 source.n268 a_n1128_n5892# 0.010552f
C848 source.n269 a_n1128_n5892# 0.019637f
C849 source.n270 a_n1128_n5892# 0.019637f
C850 source.n271 a_n1128_n5892# 0.010552f
C851 source.n272 a_n1128_n5892# 0.011173f
C852 source.n273 a_n1128_n5892# 0.024941f
C853 source.n274 a_n1128_n5892# 0.053056f
C854 source.n275 a_n1128_n5892# 0.011173f
C855 source.n276 a_n1128_n5892# 0.010552f
C856 source.n277 a_n1128_n5892# 0.043244f
C857 source.n278 a_n1128_n5892# 0.029523f
C858 source.n279 a_n1128_n5892# 2.00928f
C859 source.n280 a_n1128_n5892# 0.027071f
C860 source.n281 a_n1128_n5892# 0.019637f
C861 source.n282 a_n1128_n5892# 0.010552f
C862 source.n283 a_n1128_n5892# 0.024941f
C863 source.n284 a_n1128_n5892# 0.011173f
C864 source.n285 a_n1128_n5892# 0.019637f
C865 source.n286 a_n1128_n5892# 0.010552f
C866 source.n287 a_n1128_n5892# 0.024941f
C867 source.n288 a_n1128_n5892# 0.011173f
C868 source.n289 a_n1128_n5892# 0.019637f
C869 source.n290 a_n1128_n5892# 0.010552f
C870 source.n291 a_n1128_n5892# 0.024941f
C871 source.n292 a_n1128_n5892# 0.011173f
C872 source.n293 a_n1128_n5892# 0.019637f
C873 source.n294 a_n1128_n5892# 0.010552f
C874 source.n295 a_n1128_n5892# 0.024941f
C875 source.n296 a_n1128_n5892# 0.011173f
C876 source.n297 a_n1128_n5892# 0.019637f
C877 source.n298 a_n1128_n5892# 0.010552f
C878 source.n299 a_n1128_n5892# 0.024941f
C879 source.n300 a_n1128_n5892# 0.011173f
C880 source.n301 a_n1128_n5892# 0.019637f
C881 source.n302 a_n1128_n5892# 0.010552f
C882 source.n303 a_n1128_n5892# 0.024941f
C883 source.n304 a_n1128_n5892# 0.011173f
C884 source.n305 a_n1128_n5892# 0.019637f
C885 source.n306 a_n1128_n5892# 0.010552f
C886 source.n307 a_n1128_n5892# 0.024941f
C887 source.n308 a_n1128_n5892# 0.011173f
C888 source.n309 a_n1128_n5892# 0.019637f
C889 source.n310 a_n1128_n5892# 0.010552f
C890 source.n311 a_n1128_n5892# 0.024941f
C891 source.n312 a_n1128_n5892# 0.011173f
C892 source.n313 a_n1128_n5892# 0.019637f
C893 source.n314 a_n1128_n5892# 0.010862f
C894 source.n315 a_n1128_n5892# 0.024941f
C895 source.n316 a_n1128_n5892# 0.011173f
C896 source.n317 a_n1128_n5892# 0.019637f
C897 source.n318 a_n1128_n5892# 0.010552f
C898 source.n319 a_n1128_n5892# 0.024941f
C899 source.n320 a_n1128_n5892# 0.011173f
C900 source.n321 a_n1128_n5892# 0.019637f
C901 source.n322 a_n1128_n5892# 0.010552f
C902 source.n323 a_n1128_n5892# 0.018706f
C903 source.n324 a_n1128_n5892# 0.017631f
C904 source.t1 a_n1128_n5892# 0.043499f
C905 source.n325 a_n1128_n5892# 0.239586f
C906 source.n326 a_n1128_n5892# 2.12609f
C907 source.n327 a_n1128_n5892# 0.010552f
C908 source.n328 a_n1128_n5892# 0.011173f
C909 source.n329 a_n1128_n5892# 0.024941f
C910 source.n330 a_n1128_n5892# 0.024941f
C911 source.n331 a_n1128_n5892# 0.011173f
C912 source.n332 a_n1128_n5892# 0.010552f
C913 source.n333 a_n1128_n5892# 0.019637f
C914 source.n334 a_n1128_n5892# 0.019637f
C915 source.n335 a_n1128_n5892# 0.010552f
C916 source.n336 a_n1128_n5892# 0.011173f
C917 source.n337 a_n1128_n5892# 0.024941f
C918 source.n338 a_n1128_n5892# 0.024941f
C919 source.n339 a_n1128_n5892# 0.011173f
C920 source.n340 a_n1128_n5892# 0.010552f
C921 source.n341 a_n1128_n5892# 0.019637f
C922 source.n342 a_n1128_n5892# 0.019637f
C923 source.n343 a_n1128_n5892# 0.010552f
C924 source.n344 a_n1128_n5892# 0.010552f
C925 source.n345 a_n1128_n5892# 0.011173f
C926 source.n346 a_n1128_n5892# 0.024941f
C927 source.n347 a_n1128_n5892# 0.024941f
C928 source.n348 a_n1128_n5892# 0.024941f
C929 source.n349 a_n1128_n5892# 0.010862f
C930 source.n350 a_n1128_n5892# 0.010552f
C931 source.n351 a_n1128_n5892# 0.019637f
C932 source.n352 a_n1128_n5892# 0.019637f
C933 source.n353 a_n1128_n5892# 0.010552f
C934 source.n354 a_n1128_n5892# 0.011173f
C935 source.n355 a_n1128_n5892# 0.024941f
C936 source.n356 a_n1128_n5892# 0.024941f
C937 source.n357 a_n1128_n5892# 0.011173f
C938 source.n358 a_n1128_n5892# 0.010552f
C939 source.n359 a_n1128_n5892# 0.019637f
C940 source.n360 a_n1128_n5892# 0.019637f
C941 source.n361 a_n1128_n5892# 0.010552f
C942 source.n362 a_n1128_n5892# 0.011173f
C943 source.n363 a_n1128_n5892# 0.024941f
C944 source.n364 a_n1128_n5892# 0.024941f
C945 source.n365 a_n1128_n5892# 0.011173f
C946 source.n366 a_n1128_n5892# 0.010552f
C947 source.n367 a_n1128_n5892# 0.019637f
C948 source.n368 a_n1128_n5892# 0.019637f
C949 source.n369 a_n1128_n5892# 0.010552f
C950 source.n370 a_n1128_n5892# 0.011173f
C951 source.n371 a_n1128_n5892# 0.024941f
C952 source.n372 a_n1128_n5892# 0.024941f
C953 source.n373 a_n1128_n5892# 0.011173f
C954 source.n374 a_n1128_n5892# 0.010552f
C955 source.n375 a_n1128_n5892# 0.019637f
C956 source.n376 a_n1128_n5892# 0.019637f
C957 source.n377 a_n1128_n5892# 0.010552f
C958 source.n378 a_n1128_n5892# 0.011173f
C959 source.n379 a_n1128_n5892# 0.024941f
C960 source.n380 a_n1128_n5892# 0.024941f
C961 source.n381 a_n1128_n5892# 0.011173f
C962 source.n382 a_n1128_n5892# 0.010552f
C963 source.n383 a_n1128_n5892# 0.019637f
C964 source.n384 a_n1128_n5892# 0.019637f
C965 source.n385 a_n1128_n5892# 0.010552f
C966 source.n386 a_n1128_n5892# 0.011173f
C967 source.n387 a_n1128_n5892# 0.024941f
C968 source.n388 a_n1128_n5892# 0.024941f
C969 source.n389 a_n1128_n5892# 0.024941f
C970 source.n390 a_n1128_n5892# 0.011173f
C971 source.n391 a_n1128_n5892# 0.010552f
C972 source.n392 a_n1128_n5892# 0.019637f
C973 source.n393 a_n1128_n5892# 0.019637f
C974 source.n394 a_n1128_n5892# 0.010552f
C975 source.n395 a_n1128_n5892# 0.010862f
C976 source.n396 a_n1128_n5892# 0.010862f
C977 source.n397 a_n1128_n5892# 0.024941f
C978 source.n398 a_n1128_n5892# 0.024941f
C979 source.n399 a_n1128_n5892# 0.011173f
C980 source.n400 a_n1128_n5892# 0.010552f
C981 source.n401 a_n1128_n5892# 0.019637f
C982 source.n402 a_n1128_n5892# 0.019637f
C983 source.n403 a_n1128_n5892# 0.010552f
C984 source.n404 a_n1128_n5892# 0.011173f
C985 source.n405 a_n1128_n5892# 0.024941f
C986 source.n406 a_n1128_n5892# 0.024941f
C987 source.n407 a_n1128_n5892# 0.011173f
C988 source.n408 a_n1128_n5892# 0.010552f
C989 source.n409 a_n1128_n5892# 0.019637f
C990 source.n410 a_n1128_n5892# 0.019637f
C991 source.n411 a_n1128_n5892# 0.010552f
C992 source.n412 a_n1128_n5892# 0.011173f
C993 source.n413 a_n1128_n5892# 0.024941f
C994 source.n414 a_n1128_n5892# 0.053056f
C995 source.n415 a_n1128_n5892# 0.011173f
C996 source.n416 a_n1128_n5892# 0.010552f
C997 source.n417 a_n1128_n5892# 0.043244f
C998 source.n418 a_n1128_n5892# 0.029523f
C999 source.n419 a_n1128_n5892# 2.00928f
C1000 source.n420 a_n1128_n5892# 0.027071f
C1001 source.n421 a_n1128_n5892# 0.019637f
C1002 source.n422 a_n1128_n5892# 0.010552f
C1003 source.n423 a_n1128_n5892# 0.024941f
C1004 source.n424 a_n1128_n5892# 0.011173f
C1005 source.n425 a_n1128_n5892# 0.019637f
C1006 source.n426 a_n1128_n5892# 0.010552f
C1007 source.n427 a_n1128_n5892# 0.024941f
C1008 source.n428 a_n1128_n5892# 0.011173f
C1009 source.n429 a_n1128_n5892# 0.019637f
C1010 source.n430 a_n1128_n5892# 0.010552f
C1011 source.n431 a_n1128_n5892# 0.024941f
C1012 source.n432 a_n1128_n5892# 0.011173f
C1013 source.n433 a_n1128_n5892# 0.019637f
C1014 source.n434 a_n1128_n5892# 0.010552f
C1015 source.n435 a_n1128_n5892# 0.024941f
C1016 source.n436 a_n1128_n5892# 0.011173f
C1017 source.n437 a_n1128_n5892# 0.019637f
C1018 source.n438 a_n1128_n5892# 0.010552f
C1019 source.n439 a_n1128_n5892# 0.024941f
C1020 source.n440 a_n1128_n5892# 0.011173f
C1021 source.n441 a_n1128_n5892# 0.019637f
C1022 source.n442 a_n1128_n5892# 0.010552f
C1023 source.n443 a_n1128_n5892# 0.024941f
C1024 source.n444 a_n1128_n5892# 0.011173f
C1025 source.n445 a_n1128_n5892# 0.019637f
C1026 source.n446 a_n1128_n5892# 0.010552f
C1027 source.n447 a_n1128_n5892# 0.024941f
C1028 source.n448 a_n1128_n5892# 0.011173f
C1029 source.n449 a_n1128_n5892# 0.019637f
C1030 source.n450 a_n1128_n5892# 0.010552f
C1031 source.n451 a_n1128_n5892# 0.024941f
C1032 source.n452 a_n1128_n5892# 0.011173f
C1033 source.n453 a_n1128_n5892# 0.019637f
C1034 source.n454 a_n1128_n5892# 0.010862f
C1035 source.n455 a_n1128_n5892# 0.024941f
C1036 source.n456 a_n1128_n5892# 0.011173f
C1037 source.n457 a_n1128_n5892# 0.019637f
C1038 source.n458 a_n1128_n5892# 0.010552f
C1039 source.n459 a_n1128_n5892# 0.024941f
C1040 source.n460 a_n1128_n5892# 0.011173f
C1041 source.n461 a_n1128_n5892# 0.019637f
C1042 source.n462 a_n1128_n5892# 0.010552f
C1043 source.n463 a_n1128_n5892# 0.018706f
C1044 source.n464 a_n1128_n5892# 0.017631f
C1045 source.t3 a_n1128_n5892# 0.043499f
C1046 source.n465 a_n1128_n5892# 0.239586f
C1047 source.n466 a_n1128_n5892# 2.12609f
C1048 source.n467 a_n1128_n5892# 0.010552f
C1049 source.n468 a_n1128_n5892# 0.011173f
C1050 source.n469 a_n1128_n5892# 0.024941f
C1051 source.n470 a_n1128_n5892# 0.024941f
C1052 source.n471 a_n1128_n5892# 0.011173f
C1053 source.n472 a_n1128_n5892# 0.010552f
C1054 source.n473 a_n1128_n5892# 0.019637f
C1055 source.n474 a_n1128_n5892# 0.019637f
C1056 source.n475 a_n1128_n5892# 0.010552f
C1057 source.n476 a_n1128_n5892# 0.011173f
C1058 source.n477 a_n1128_n5892# 0.024941f
C1059 source.n478 a_n1128_n5892# 0.024941f
C1060 source.n479 a_n1128_n5892# 0.011173f
C1061 source.n480 a_n1128_n5892# 0.010552f
C1062 source.n481 a_n1128_n5892# 0.019637f
C1063 source.n482 a_n1128_n5892# 0.019637f
C1064 source.n483 a_n1128_n5892# 0.010552f
C1065 source.n484 a_n1128_n5892# 0.010552f
C1066 source.n485 a_n1128_n5892# 0.011173f
C1067 source.n486 a_n1128_n5892# 0.024941f
C1068 source.n487 a_n1128_n5892# 0.024941f
C1069 source.n488 a_n1128_n5892# 0.024941f
C1070 source.n489 a_n1128_n5892# 0.010862f
C1071 source.n490 a_n1128_n5892# 0.010552f
C1072 source.n491 a_n1128_n5892# 0.019637f
C1073 source.n492 a_n1128_n5892# 0.019637f
C1074 source.n493 a_n1128_n5892# 0.010552f
C1075 source.n494 a_n1128_n5892# 0.011173f
C1076 source.n495 a_n1128_n5892# 0.024941f
C1077 source.n496 a_n1128_n5892# 0.024941f
C1078 source.n497 a_n1128_n5892# 0.011173f
C1079 source.n498 a_n1128_n5892# 0.010552f
C1080 source.n499 a_n1128_n5892# 0.019637f
C1081 source.n500 a_n1128_n5892# 0.019637f
C1082 source.n501 a_n1128_n5892# 0.010552f
C1083 source.n502 a_n1128_n5892# 0.011173f
C1084 source.n503 a_n1128_n5892# 0.024941f
C1085 source.n504 a_n1128_n5892# 0.024941f
C1086 source.n505 a_n1128_n5892# 0.011173f
C1087 source.n506 a_n1128_n5892# 0.010552f
C1088 source.n507 a_n1128_n5892# 0.019637f
C1089 source.n508 a_n1128_n5892# 0.019637f
C1090 source.n509 a_n1128_n5892# 0.010552f
C1091 source.n510 a_n1128_n5892# 0.011173f
C1092 source.n511 a_n1128_n5892# 0.024941f
C1093 source.n512 a_n1128_n5892# 0.024941f
C1094 source.n513 a_n1128_n5892# 0.011173f
C1095 source.n514 a_n1128_n5892# 0.010552f
C1096 source.n515 a_n1128_n5892# 0.019637f
C1097 source.n516 a_n1128_n5892# 0.019637f
C1098 source.n517 a_n1128_n5892# 0.010552f
C1099 source.n518 a_n1128_n5892# 0.011173f
C1100 source.n519 a_n1128_n5892# 0.024941f
C1101 source.n520 a_n1128_n5892# 0.024941f
C1102 source.n521 a_n1128_n5892# 0.011173f
C1103 source.n522 a_n1128_n5892# 0.010552f
C1104 source.n523 a_n1128_n5892# 0.019637f
C1105 source.n524 a_n1128_n5892# 0.019637f
C1106 source.n525 a_n1128_n5892# 0.010552f
C1107 source.n526 a_n1128_n5892# 0.011173f
C1108 source.n527 a_n1128_n5892# 0.024941f
C1109 source.n528 a_n1128_n5892# 0.024941f
C1110 source.n529 a_n1128_n5892# 0.024941f
C1111 source.n530 a_n1128_n5892# 0.011173f
C1112 source.n531 a_n1128_n5892# 0.010552f
C1113 source.n532 a_n1128_n5892# 0.019637f
C1114 source.n533 a_n1128_n5892# 0.019637f
C1115 source.n534 a_n1128_n5892# 0.010552f
C1116 source.n535 a_n1128_n5892# 0.010862f
C1117 source.n536 a_n1128_n5892# 0.010862f
C1118 source.n537 a_n1128_n5892# 0.024941f
C1119 source.n538 a_n1128_n5892# 0.024941f
C1120 source.n539 a_n1128_n5892# 0.011173f
C1121 source.n540 a_n1128_n5892# 0.010552f
C1122 source.n541 a_n1128_n5892# 0.019637f
C1123 source.n542 a_n1128_n5892# 0.019637f
C1124 source.n543 a_n1128_n5892# 0.010552f
C1125 source.n544 a_n1128_n5892# 0.011173f
C1126 source.n545 a_n1128_n5892# 0.024941f
C1127 source.n546 a_n1128_n5892# 0.024941f
C1128 source.n547 a_n1128_n5892# 0.011173f
C1129 source.n548 a_n1128_n5892# 0.010552f
C1130 source.n549 a_n1128_n5892# 0.019637f
C1131 source.n550 a_n1128_n5892# 0.019637f
C1132 source.n551 a_n1128_n5892# 0.010552f
C1133 source.n552 a_n1128_n5892# 0.011173f
C1134 source.n553 a_n1128_n5892# 0.024941f
C1135 source.n554 a_n1128_n5892# 0.053056f
C1136 source.n555 a_n1128_n5892# 0.011173f
C1137 source.n556 a_n1128_n5892# 0.010552f
C1138 source.n557 a_n1128_n5892# 0.043244f
C1139 source.n558 a_n1128_n5892# 0.029523f
C1140 source.n559 a_n1128_n5892# 0.231201f
C1141 source.n560 a_n1128_n5892# 2.10905f
C1142 minus.t0 a_n1128_n5892# 3.0374f
C1143 minus.t1 a_n1128_n5892# 2.91174f
C1144 minus.n0 a_n1128_n5892# 7.61428f
.ends

