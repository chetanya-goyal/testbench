* NGSPICE file created from diffpair639.ext - technology: sky130A

.subckt diffpair639 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t38 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 drain_right.t23 minus.t0 source.t12 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X2 source.t16 minus.t1 drain_right.t22 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X3 source.t14 minus.t2 drain_right.t21 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X4 source.t37 plus.t1 drain_left.t22 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X5 source.t36 plus.t2 drain_left.t21 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X6 drain_right.t20 minus.t3 source.t6 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X7 drain_right.t19 minus.t4 source.t11 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X8 a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X9 source.t23 plus.t3 drain_left.t20 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 drain_right.t18 minus.t5 source.t8 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X11 source.t47 minus.t6 drain_right.t17 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 drain_left.t19 plus.t4 source.t35 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X13 a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X14 drain_right.t16 minus.t7 source.t15 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X15 source.t30 plus.t5 drain_left.t18 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X16 source.t29 plus.t6 drain_left.t17 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_right.t15 minus.t8 source.t45 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X18 source.t3 minus.t9 drain_right.t14 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X19 drain_left.t16 plus.t7 source.t28 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 drain_left.t15 plus.t8 source.t39 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X21 source.t4 minus.t10 drain_right.t13 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X22 source.t46 minus.t11 drain_right.t12 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X23 source.t27 plus.t9 drain_left.t14 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X24 drain_right.t11 minus.t12 source.t44 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X25 drain_right.t10 minus.t13 source.t0 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X26 drain_left.t13 plus.t10 source.t22 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X27 drain_right.t9 minus.t14 source.t7 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X28 drain_right.t8 minus.t15 source.t5 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X29 drain_left.t12 plus.t11 source.t26 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X30 source.t25 plus.t12 drain_left.t11 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X31 source.t10 minus.t16 drain_right.t7 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X32 drain_left.t10 plus.t13 source.t40 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X33 source.t19 minus.t17 drain_right.t6 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X34 drain_right.t5 minus.t18 source.t13 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X35 drain_right.t4 minus.t19 source.t17 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X36 source.t42 plus.t14 drain_left.t9 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X37 a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X38 drain_left.t8 plus.t15 source.t41 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X39 drain_left.t7 plus.t16 source.t43 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X40 source.t1 minus.t20 drain_right.t3 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X41 source.t24 plus.t17 drain_left.t6 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X42 drain_left.t5 plus.t18 source.t34 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X43 drain_left.t4 plus.t19 source.t33 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X44 source.t32 plus.t20 drain_left.t3 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X45 drain_left.t2 plus.t21 source.t31 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X46 source.t18 minus.t21 drain_right.t2 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X47 a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X48 source.t9 minus.t22 drain_right.t1 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X49 source.t21 plus.t22 drain_left.t1 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X50 source.t2 minus.t23 drain_right.t0 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X51 source.t20 plus.t23 drain_left.t0 a_n3654_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n10 plus.t22 673.04
R1 plus.n46 plus.t0 673.04
R2 plus.n34 plus.t4 651.605
R3 plus.n32 plus.t6 651.605
R4 plus.n31 plus.t8 651.605
R5 plus.n3 plus.t12 651.605
R6 plus.n25 plus.t13 651.605
R7 plus.n5 plus.t14 651.605
R8 plus.n20 plus.t15 651.605
R9 plus.n18 plus.t20 651.605
R10 plus.n8 plus.t16 651.605
R11 plus.n12 plus.t17 651.605
R12 plus.n11 plus.t21 651.605
R13 plus.n70 plus.t2 651.605
R14 plus.n68 plus.t10 651.605
R15 plus.n67 plus.t23 651.605
R16 plus.n39 plus.t7 651.605
R17 plus.n61 plus.t3 651.605
R18 plus.n41 plus.t11 651.605
R19 plus.n56 plus.t1 651.605
R20 plus.n54 plus.t18 651.605
R21 plus.n44 plus.t5 651.605
R22 plus.n48 plus.t19 651.605
R23 plus.n47 plus.t9 651.605
R24 plus.n14 plus.n13 161.3
R25 plus.n15 plus.n8 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n18 plus.n7 161.3
R28 plus.n19 plus.n6 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n25 plus.n4 161.3
R31 plus.n27 plus.n26 161.3
R32 plus.n28 plus.n3 161.3
R33 plus.n30 plus.n29 161.3
R34 plus.n33 plus.n0 161.3
R35 plus.n35 plus.n34 161.3
R36 plus.n50 plus.n49 161.3
R37 plus.n51 plus.n44 161.3
R38 plus.n53 plus.n52 161.3
R39 plus.n54 plus.n43 161.3
R40 plus.n55 plus.n42 161.3
R41 plus.n60 plus.n59 161.3
R42 plus.n61 plus.n40 161.3
R43 plus.n63 plus.n62 161.3
R44 plus.n64 plus.n39 161.3
R45 plus.n66 plus.n65 161.3
R46 plus.n69 plus.n36 161.3
R47 plus.n71 plus.n70 161.3
R48 plus.n12 plus.n9 80.6037
R49 plus.n21 plus.n20 80.6037
R50 plus.n22 plus.n5 80.6037
R51 plus.n31 plus.n2 80.6037
R52 plus.n32 plus.n1 80.6037
R53 plus.n48 plus.n45 80.6037
R54 plus.n57 plus.n56 80.6037
R55 plus.n58 plus.n41 80.6037
R56 plus.n67 plus.n38 80.6037
R57 plus.n68 plus.n37 80.6037
R58 plus.n32 plus.n31 48.2005
R59 plus.n20 plus.n5 48.2005
R60 plus.n12 plus.n11 48.2005
R61 plus.n68 plus.n67 48.2005
R62 plus.n56 plus.n41 48.2005
R63 plus.n48 plus.n47 48.2005
R64 plus.n31 plus.n30 44.549
R65 plus.n13 plus.n12 44.549
R66 plus.n67 plus.n66 44.549
R67 plus.n49 plus.n48 44.549
R68 plus.n24 plus.n5 41.6278
R69 plus.n20 plus.n19 41.6278
R70 plus.n60 plus.n41 41.6278
R71 plus.n56 plus.n55 41.6278
R72 plus plus.n71 40.0331
R73 plus.n33 plus.n32 38.7066
R74 plus.n69 plus.n68 38.7066
R75 plus.n10 plus.n9 31.6825
R76 plus.n46 plus.n45 31.6825
R77 plus.n26 plus.n3 25.5611
R78 plus.n17 plus.n8 25.5611
R79 plus.n62 plus.n39 25.5611
R80 plus.n53 plus.n44 25.5611
R81 plus.n26 plus.n25 22.6399
R82 plus.n18 plus.n17 22.6399
R83 plus.n62 plus.n61 22.6399
R84 plus.n54 plus.n53 22.6399
R85 plus.n11 plus.n10 17.2341
R86 plus.n47 plus.n46 17.2341
R87 plus plus.n35 15.3338
R88 plus.n34 plus.n33 9.49444
R89 plus.n70 plus.n69 9.49444
R90 plus.n25 plus.n24 6.57323
R91 plus.n19 plus.n18 6.57323
R92 plus.n61 plus.n60 6.57323
R93 plus.n55 plus.n54 6.57323
R94 plus.n30 plus.n3 3.65202
R95 plus.n13 plus.n8 3.65202
R96 plus.n66 plus.n39 3.65202
R97 plus.n49 plus.n44 3.65202
R98 plus.n22 plus.n21 0.380177
R99 plus.n2 plus.n1 0.380177
R100 plus.n38 plus.n37 0.380177
R101 plus.n58 plus.n57 0.380177
R102 plus.n14 plus.n9 0.285035
R103 plus.n21 plus.n6 0.285035
R104 plus.n23 plus.n22 0.285035
R105 plus.n29 plus.n2 0.285035
R106 plus.n1 plus.n0 0.285035
R107 plus.n37 plus.n36 0.285035
R108 plus.n65 plus.n38 0.285035
R109 plus.n59 plus.n58 0.285035
R110 plus.n57 plus.n42 0.285035
R111 plus.n50 plus.n45 0.285035
R112 plus.n15 plus.n14 0.189894
R113 plus.n16 plus.n15 0.189894
R114 plus.n16 plus.n7 0.189894
R115 plus.n7 plus.n6 0.189894
R116 plus.n23 plus.n4 0.189894
R117 plus.n27 plus.n4 0.189894
R118 plus.n28 plus.n27 0.189894
R119 plus.n29 plus.n28 0.189894
R120 plus.n35 plus.n0 0.189894
R121 plus.n71 plus.n36 0.189894
R122 plus.n65 plus.n64 0.189894
R123 plus.n64 plus.n63 0.189894
R124 plus.n63 plus.n40 0.189894
R125 plus.n59 plus.n40 0.189894
R126 plus.n43 plus.n42 0.189894
R127 plus.n52 plus.n43 0.189894
R128 plus.n52 plus.n51 0.189894
R129 plus.n51 plus.n50 0.189894
R130 source.n0 source.t35 44.1297
R131 source.n11 source.t21 44.1296
R132 source.n12 source.t7 44.1296
R133 source.n23 source.t46 44.1296
R134 source.n47 source.t12 44.1295
R135 source.n36 source.t14 44.1295
R136 source.n35 source.t38 44.1295
R137 source.n24 source.t36 44.1295
R138 source.n2 source.n1 43.1397
R139 source.n4 source.n3 43.1397
R140 source.n6 source.n5 43.1397
R141 source.n8 source.n7 43.1397
R142 source.n10 source.n9 43.1397
R143 source.n14 source.n13 43.1397
R144 source.n16 source.n15 43.1397
R145 source.n18 source.n17 43.1397
R146 source.n20 source.n19 43.1397
R147 source.n22 source.n21 43.1397
R148 source.n46 source.n45 43.1396
R149 source.n44 source.n43 43.1396
R150 source.n42 source.n41 43.1396
R151 source.n40 source.n39 43.1396
R152 source.n38 source.n37 43.1396
R153 source.n34 source.n33 43.1396
R154 source.n32 source.n31 43.1396
R155 source.n30 source.n29 43.1396
R156 source.n28 source.n27 43.1396
R157 source.n26 source.n25 43.1396
R158 source.n24 source.n23 28.3225
R159 source.n48 source.n0 22.5725
R160 source.n48 source.n47 5.7505
R161 source.n45 source.t11 0.9905
R162 source.n45 source.t3 0.9905
R163 source.n43 source.t6 0.9905
R164 source.n43 source.t2 0.9905
R165 source.n41 source.t8 0.9905
R166 source.n41 source.t18 0.9905
R167 source.n39 source.t15 0.9905
R168 source.n39 source.t16 0.9905
R169 source.n37 source.t5 0.9905
R170 source.n37 source.t9 0.9905
R171 source.n33 source.t33 0.9905
R172 source.n33 source.t27 0.9905
R173 source.n31 source.t34 0.9905
R174 source.n31 source.t30 0.9905
R175 source.n29 source.t26 0.9905
R176 source.n29 source.t37 0.9905
R177 source.n27 source.t28 0.9905
R178 source.n27 source.t23 0.9905
R179 source.n25 source.t22 0.9905
R180 source.n25 source.t20 0.9905
R181 source.n1 source.t39 0.9905
R182 source.n1 source.t29 0.9905
R183 source.n3 source.t40 0.9905
R184 source.n3 source.t25 0.9905
R185 source.n5 source.t41 0.9905
R186 source.n5 source.t42 0.9905
R187 source.n7 source.t43 0.9905
R188 source.n7 source.t32 0.9905
R189 source.n9 source.t31 0.9905
R190 source.n9 source.t24 0.9905
R191 source.n13 source.t45 0.9905
R192 source.n13 source.t4 0.9905
R193 source.n15 source.t17 0.9905
R194 source.n15 source.t19 0.9905
R195 source.n17 source.t44 0.9905
R196 source.n17 source.t10 0.9905
R197 source.n19 source.t13 0.9905
R198 source.n19 source.t1 0.9905
R199 source.n21 source.t0 0.9905
R200 source.n21 source.t47 0.9905
R201 source.n23 source.n22 0.974638
R202 source.n22 source.n20 0.974638
R203 source.n20 source.n18 0.974638
R204 source.n18 source.n16 0.974638
R205 source.n16 source.n14 0.974638
R206 source.n14 source.n12 0.974638
R207 source.n11 source.n10 0.974638
R208 source.n10 source.n8 0.974638
R209 source.n8 source.n6 0.974638
R210 source.n6 source.n4 0.974638
R211 source.n4 source.n2 0.974638
R212 source.n2 source.n0 0.974638
R213 source.n26 source.n24 0.974638
R214 source.n28 source.n26 0.974638
R215 source.n30 source.n28 0.974638
R216 source.n32 source.n30 0.974638
R217 source.n34 source.n32 0.974638
R218 source.n35 source.n34 0.974638
R219 source.n38 source.n36 0.974638
R220 source.n40 source.n38 0.974638
R221 source.n42 source.n40 0.974638
R222 source.n44 source.n42 0.974638
R223 source.n46 source.n44 0.974638
R224 source.n47 source.n46 0.974638
R225 source.n12 source.n11 0.470328
R226 source.n36 source.n35 0.470328
R227 source source.n48 0.188
R228 drain_left.n13 drain_left.n11 60.7926
R229 drain_left.n7 drain_left.n5 60.7925
R230 drain_left.n2 drain_left.n0 60.7925
R231 drain_left.n21 drain_left.n20 59.8185
R232 drain_left.n19 drain_left.n18 59.8185
R233 drain_left.n17 drain_left.n16 59.8185
R234 drain_left.n15 drain_left.n14 59.8185
R235 drain_left.n13 drain_left.n12 59.8185
R236 drain_left.n7 drain_left.n6 59.8184
R237 drain_left.n9 drain_left.n8 59.8184
R238 drain_left.n4 drain_left.n3 59.8184
R239 drain_left.n2 drain_left.n1 59.8184
R240 drain_left drain_left.n10 42.682
R241 drain_left drain_left.n21 6.62735
R242 drain_left.n5 drain_left.t14 0.9905
R243 drain_left.n5 drain_left.t23 0.9905
R244 drain_left.n6 drain_left.t18 0.9905
R245 drain_left.n6 drain_left.t4 0.9905
R246 drain_left.n8 drain_left.t22 0.9905
R247 drain_left.n8 drain_left.t5 0.9905
R248 drain_left.n3 drain_left.t20 0.9905
R249 drain_left.n3 drain_left.t12 0.9905
R250 drain_left.n1 drain_left.t0 0.9905
R251 drain_left.n1 drain_left.t16 0.9905
R252 drain_left.n0 drain_left.t21 0.9905
R253 drain_left.n0 drain_left.t13 0.9905
R254 drain_left.n20 drain_left.t17 0.9905
R255 drain_left.n20 drain_left.t19 0.9905
R256 drain_left.n18 drain_left.t11 0.9905
R257 drain_left.n18 drain_left.t15 0.9905
R258 drain_left.n16 drain_left.t9 0.9905
R259 drain_left.n16 drain_left.t10 0.9905
R260 drain_left.n14 drain_left.t3 0.9905
R261 drain_left.n14 drain_left.t8 0.9905
R262 drain_left.n12 drain_left.t6 0.9905
R263 drain_left.n12 drain_left.t7 0.9905
R264 drain_left.n11 drain_left.t1 0.9905
R265 drain_left.n11 drain_left.t2 0.9905
R266 drain_left.n9 drain_left.n7 0.974638
R267 drain_left.n4 drain_left.n2 0.974638
R268 drain_left.n15 drain_left.n13 0.974638
R269 drain_left.n17 drain_left.n15 0.974638
R270 drain_left.n19 drain_left.n17 0.974638
R271 drain_left.n21 drain_left.n19 0.974638
R272 drain_left.n10 drain_left.n9 0.432223
R273 drain_left.n10 drain_left.n4 0.432223
R274 minus.n8 minus.t14 673.04
R275 minus.n44 minus.t2 673.04
R276 minus.n9 minus.t10 651.605
R277 minus.n10 minus.t8 651.605
R278 minus.n14 minus.t17 651.605
R279 minus.n16 minus.t19 651.605
R280 minus.n20 minus.t16 651.605
R281 minus.n21 minus.t12 651.605
R282 minus.n3 minus.t20 651.605
R283 minus.n27 minus.t18 651.605
R284 minus.n1 minus.t6 651.605
R285 minus.n32 minus.t13 651.605
R286 minus.n34 minus.t11 651.605
R287 minus.n45 minus.t15 651.605
R288 minus.n46 minus.t22 651.605
R289 minus.n50 minus.t7 651.605
R290 minus.n52 minus.t1 651.605
R291 minus.n56 minus.t5 651.605
R292 minus.n57 minus.t21 651.605
R293 minus.n39 minus.t3 651.605
R294 minus.n63 minus.t23 651.605
R295 minus.n37 minus.t4 651.605
R296 minus.n68 minus.t9 651.605
R297 minus.n70 minus.t0 651.605
R298 minus.n35 minus.n34 161.3
R299 minus.n33 minus.n0 161.3
R300 minus.n29 minus.n28 161.3
R301 minus.n27 minus.n2 161.3
R302 minus.n26 minus.n25 161.3
R303 minus.n24 minus.n3 161.3
R304 minus.n23 minus.n22 161.3
R305 minus.n18 minus.n5 161.3
R306 minus.n17 minus.n16 161.3
R307 minus.n15 minus.n6 161.3
R308 minus.n14 minus.n13 161.3
R309 minus.n12 minus.n7 161.3
R310 minus.n71 minus.n70 161.3
R311 minus.n69 minus.n36 161.3
R312 minus.n65 minus.n64 161.3
R313 minus.n63 minus.n38 161.3
R314 minus.n62 minus.n61 161.3
R315 minus.n60 minus.n39 161.3
R316 minus.n59 minus.n58 161.3
R317 minus.n54 minus.n41 161.3
R318 minus.n53 minus.n52 161.3
R319 minus.n51 minus.n42 161.3
R320 minus.n50 minus.n49 161.3
R321 minus.n48 minus.n43 161.3
R322 minus.n32 minus.n31 80.6037
R323 minus.n30 minus.n1 80.6037
R324 minus.n21 minus.n4 80.6037
R325 minus.n20 minus.n19 80.6037
R326 minus.n11 minus.n10 80.6037
R327 minus.n68 minus.n67 80.6037
R328 minus.n66 minus.n37 80.6037
R329 minus.n57 minus.n40 80.6037
R330 minus.n56 minus.n55 80.6037
R331 minus.n47 minus.n46 80.6037
R332 minus.n72 minus.n35 49.1823
R333 minus.n10 minus.n9 48.2005
R334 minus.n21 minus.n20 48.2005
R335 minus.n32 minus.n1 48.2005
R336 minus.n46 minus.n45 48.2005
R337 minus.n57 minus.n56 48.2005
R338 minus.n68 minus.n37 48.2005
R339 minus.n10 minus.n7 44.549
R340 minus.n28 minus.n1 44.549
R341 minus.n46 minus.n43 44.549
R342 minus.n64 minus.n37 44.549
R343 minus.n20 minus.n5 41.6278
R344 minus.n22 minus.n21 41.6278
R345 minus.n56 minus.n41 41.6278
R346 minus.n58 minus.n57 41.6278
R347 minus.n33 minus.n32 38.7066
R348 minus.n69 minus.n68 38.7066
R349 minus.n11 minus.n8 31.6825
R350 minus.n47 minus.n44 31.6825
R351 minus.n15 minus.n14 25.5611
R352 minus.n27 minus.n26 25.5611
R353 minus.n51 minus.n50 25.5611
R354 minus.n63 minus.n62 25.5611
R355 minus.n16 minus.n15 22.6399
R356 minus.n26 minus.n3 22.6399
R357 minus.n52 minus.n51 22.6399
R358 minus.n62 minus.n39 22.6399
R359 minus.n9 minus.n8 17.2341
R360 minus.n45 minus.n44 17.2341
R361 minus.n34 minus.n33 9.49444
R362 minus.n70 minus.n69 9.49444
R363 minus.n72 minus.n71 6.65959
R364 minus.n16 minus.n5 6.57323
R365 minus.n22 minus.n3 6.57323
R366 minus.n52 minus.n41 6.57323
R367 minus.n58 minus.n39 6.57323
R368 minus.n14 minus.n7 3.65202
R369 minus.n28 minus.n27 3.65202
R370 minus.n50 minus.n43 3.65202
R371 minus.n64 minus.n63 3.65202
R372 minus.n31 minus.n30 0.380177
R373 minus.n19 minus.n4 0.380177
R374 minus.n55 minus.n40 0.380177
R375 minus.n67 minus.n66 0.380177
R376 minus.n31 minus.n0 0.285035
R377 minus.n30 minus.n29 0.285035
R378 minus.n23 minus.n4 0.285035
R379 minus.n19 minus.n18 0.285035
R380 minus.n12 minus.n11 0.285035
R381 minus.n48 minus.n47 0.285035
R382 minus.n55 minus.n54 0.285035
R383 minus.n59 minus.n40 0.285035
R384 minus.n66 minus.n65 0.285035
R385 minus.n67 minus.n36 0.285035
R386 minus.n35 minus.n0 0.189894
R387 minus.n29 minus.n2 0.189894
R388 minus.n25 minus.n2 0.189894
R389 minus.n25 minus.n24 0.189894
R390 minus.n24 minus.n23 0.189894
R391 minus.n18 minus.n17 0.189894
R392 minus.n17 minus.n6 0.189894
R393 minus.n13 minus.n6 0.189894
R394 minus.n13 minus.n12 0.189894
R395 minus.n49 minus.n48 0.189894
R396 minus.n49 minus.n42 0.189894
R397 minus.n53 minus.n42 0.189894
R398 minus.n54 minus.n53 0.189894
R399 minus.n60 minus.n59 0.189894
R400 minus.n61 minus.n60 0.189894
R401 minus.n61 minus.n38 0.189894
R402 minus.n65 minus.n38 0.189894
R403 minus.n71 minus.n36 0.189894
R404 minus minus.n72 0.188
R405 drain_right.n13 drain_right.n11 60.7926
R406 drain_right.n7 drain_right.n5 60.7925
R407 drain_right.n2 drain_right.n0 60.7925
R408 drain_right.n13 drain_right.n12 59.8185
R409 drain_right.n15 drain_right.n14 59.8185
R410 drain_right.n17 drain_right.n16 59.8185
R411 drain_right.n19 drain_right.n18 59.8185
R412 drain_right.n21 drain_right.n20 59.8185
R413 drain_right.n7 drain_right.n6 59.8184
R414 drain_right.n9 drain_right.n8 59.8184
R415 drain_right.n4 drain_right.n3 59.8184
R416 drain_right.n2 drain_right.n1 59.8184
R417 drain_right drain_right.n10 42.1288
R418 drain_right drain_right.n21 6.62735
R419 drain_right.n5 drain_right.t14 0.9905
R420 drain_right.n5 drain_right.t23 0.9905
R421 drain_right.n6 drain_right.t0 0.9905
R422 drain_right.n6 drain_right.t19 0.9905
R423 drain_right.n8 drain_right.t2 0.9905
R424 drain_right.n8 drain_right.t20 0.9905
R425 drain_right.n3 drain_right.t22 0.9905
R426 drain_right.n3 drain_right.t18 0.9905
R427 drain_right.n1 drain_right.t1 0.9905
R428 drain_right.n1 drain_right.t16 0.9905
R429 drain_right.n0 drain_right.t21 0.9905
R430 drain_right.n0 drain_right.t8 0.9905
R431 drain_right.n11 drain_right.t13 0.9905
R432 drain_right.n11 drain_right.t9 0.9905
R433 drain_right.n12 drain_right.t6 0.9905
R434 drain_right.n12 drain_right.t15 0.9905
R435 drain_right.n14 drain_right.t7 0.9905
R436 drain_right.n14 drain_right.t4 0.9905
R437 drain_right.n16 drain_right.t3 0.9905
R438 drain_right.n16 drain_right.t11 0.9905
R439 drain_right.n18 drain_right.t17 0.9905
R440 drain_right.n18 drain_right.t5 0.9905
R441 drain_right.n20 drain_right.t12 0.9905
R442 drain_right.n20 drain_right.t10 0.9905
R443 drain_right.n9 drain_right.n7 0.974638
R444 drain_right.n4 drain_right.n2 0.974638
R445 drain_right.n21 drain_right.n19 0.974638
R446 drain_right.n19 drain_right.n17 0.974638
R447 drain_right.n17 drain_right.n15 0.974638
R448 drain_right.n15 drain_right.n13 0.974638
R449 drain_right.n10 drain_right.n9 0.432223
R450 drain_right.n10 drain_right.n4 0.432223
C0 plus drain_right 0.526806f
C1 source drain_right 40.760002f
C2 minus drain_right 26.2523f
C3 plus drain_left 26.6198f
C4 source drain_left 40.756897f
C5 source plus 26.3601f
C6 minus drain_left 0.175388f
C7 minus plus 9.190269f
C8 source minus 26.3461f
C9 drain_left drain_right 2.02887f
C10 drain_right a_n3654_n4888# 9.65481f
C11 drain_left a_n3654_n4888# 10.15036f
C12 source a_n3654_n4888# 14.218859f
C13 minus a_n3654_n4888# 15.413514f
C14 plus a_n3654_n4888# 17.61322f
C15 drain_right.t21 a_n3654_n4888# 0.43166f
C16 drain_right.t8 a_n3654_n4888# 0.43166f
C17 drain_right.n0 a_n3654_n4888# 3.95295f
C18 drain_right.t1 a_n3654_n4888# 0.43166f
C19 drain_right.t16 a_n3654_n4888# 0.43166f
C20 drain_right.n1 a_n3654_n4888# 3.94633f
C21 drain_right.n2 a_n3654_n4888# 0.808258f
C22 drain_right.t22 a_n3654_n4888# 0.43166f
C23 drain_right.t18 a_n3654_n4888# 0.43166f
C24 drain_right.n3 a_n3654_n4888# 3.94633f
C25 drain_right.n4 a_n3654_n4888# 0.355668f
C26 drain_right.t14 a_n3654_n4888# 0.43166f
C27 drain_right.t23 a_n3654_n4888# 0.43166f
C28 drain_right.n5 a_n3654_n4888# 3.95295f
C29 drain_right.t0 a_n3654_n4888# 0.43166f
C30 drain_right.t19 a_n3654_n4888# 0.43166f
C31 drain_right.n6 a_n3654_n4888# 3.94633f
C32 drain_right.n7 a_n3654_n4888# 0.808258f
C33 drain_right.t2 a_n3654_n4888# 0.43166f
C34 drain_right.t20 a_n3654_n4888# 0.43166f
C35 drain_right.n8 a_n3654_n4888# 3.94633f
C36 drain_right.n9 a_n3654_n4888# 0.355668f
C37 drain_right.n10 a_n3654_n4888# 2.36315f
C38 drain_right.t13 a_n3654_n4888# 0.43166f
C39 drain_right.t9 a_n3654_n4888# 0.43166f
C40 drain_right.n11 a_n3654_n4888# 3.95294f
C41 drain_right.t6 a_n3654_n4888# 0.43166f
C42 drain_right.t15 a_n3654_n4888# 0.43166f
C43 drain_right.n12 a_n3654_n4888# 3.94632f
C44 drain_right.n13 a_n3654_n4888# 0.808269f
C45 drain_right.t7 a_n3654_n4888# 0.43166f
C46 drain_right.t4 a_n3654_n4888# 0.43166f
C47 drain_right.n14 a_n3654_n4888# 3.94632f
C48 drain_right.n15 a_n3654_n4888# 0.401943f
C49 drain_right.t3 a_n3654_n4888# 0.43166f
C50 drain_right.t11 a_n3654_n4888# 0.43166f
C51 drain_right.n16 a_n3654_n4888# 3.94632f
C52 drain_right.n17 a_n3654_n4888# 0.401943f
C53 drain_right.t17 a_n3654_n4888# 0.43166f
C54 drain_right.t5 a_n3654_n4888# 0.43166f
C55 drain_right.n18 a_n3654_n4888# 3.94632f
C56 drain_right.n19 a_n3654_n4888# 0.401943f
C57 drain_right.t12 a_n3654_n4888# 0.43166f
C58 drain_right.t10 a_n3654_n4888# 0.43166f
C59 drain_right.n20 a_n3654_n4888# 3.94632f
C60 drain_right.n21 a_n3654_n4888# 0.64685f
C61 minus.n0 a_n3654_n4888# 0.049204f
C62 minus.t6 a_n3654_n4888# 1.67079f
C63 minus.n1 a_n3654_n4888# 0.630416f
C64 minus.t13 a_n3654_n4888# 1.67079f
C65 minus.n2 a_n3654_n4888# 0.036874f
C66 minus.t20 a_n3654_n4888# 1.67079f
C67 minus.n3 a_n3654_n4888# 0.619662f
C68 minus.n4 a_n3654_n4888# 0.061419f
C69 minus.n5 a_n3654_n4888# 0.008368f
C70 minus.t16 a_n3654_n4888# 1.67079f
C71 minus.n6 a_n3654_n4888# 0.036874f
C72 minus.n7 a_n3654_n4888# 0.008368f
C73 minus.t17 a_n3654_n4888# 1.67079f
C74 minus.t14 a_n3654_n4888# 1.69063f
C75 minus.n8 a_n3654_n4888# 0.60644f
C76 minus.t10 a_n3654_n4888# 1.67079f
C77 minus.n9 a_n3654_n4888# 0.630397f
C78 minus.t8 a_n3654_n4888# 1.67079f
C79 minus.n10 a_n3654_n4888# 0.630416f
C80 minus.n11 a_n3654_n4888# 0.21194f
C81 minus.n12 a_n3654_n4888# 0.049204f
C82 minus.n13 a_n3654_n4888# 0.036874f
C83 minus.n14 a_n3654_n4888# 0.619662f
C84 minus.n15 a_n3654_n4888# 0.008368f
C85 minus.t19 a_n3654_n4888# 1.67079f
C86 minus.n16 a_n3654_n4888# 0.619662f
C87 minus.n17 a_n3654_n4888# 0.036874f
C88 minus.n18 a_n3654_n4888# 0.049204f
C89 minus.n19 a_n3654_n4888# 0.061419f
C90 minus.n20 a_n3654_n4888# 0.629962f
C91 minus.t12 a_n3654_n4888# 1.67079f
C92 minus.n21 a_n3654_n4888# 0.629962f
C93 minus.n22 a_n3654_n4888# 0.008368f
C94 minus.n23 a_n3654_n4888# 0.049204f
C95 minus.n24 a_n3654_n4888# 0.036874f
C96 minus.n25 a_n3654_n4888# 0.036874f
C97 minus.n26 a_n3654_n4888# 0.008368f
C98 minus.t18 a_n3654_n4888# 1.67079f
C99 minus.n27 a_n3654_n4888# 0.619662f
C100 minus.n28 a_n3654_n4888# 0.008368f
C101 minus.n29 a_n3654_n4888# 0.049204f
C102 minus.n30 a_n3654_n4888# 0.061419f
C103 minus.n31 a_n3654_n4888# 0.061419f
C104 minus.n32 a_n3654_n4888# 0.629507f
C105 minus.n33 a_n3654_n4888# 0.008368f
C106 minus.t11 a_n3654_n4888# 1.67079f
C107 minus.n34 a_n3654_n4888# 0.616592f
C108 minus.n35 a_n3654_n4888# 2.0505f
C109 minus.n36 a_n3654_n4888# 0.049204f
C110 minus.t4 a_n3654_n4888# 1.67079f
C111 minus.n37 a_n3654_n4888# 0.630416f
C112 minus.n38 a_n3654_n4888# 0.036874f
C113 minus.t3 a_n3654_n4888# 1.67079f
C114 minus.n39 a_n3654_n4888# 0.619662f
C115 minus.n40 a_n3654_n4888# 0.061419f
C116 minus.n41 a_n3654_n4888# 0.008368f
C117 minus.n42 a_n3654_n4888# 0.036874f
C118 minus.n43 a_n3654_n4888# 0.008368f
C119 minus.t2 a_n3654_n4888# 1.69063f
C120 minus.n44 a_n3654_n4888# 0.60644f
C121 minus.t15 a_n3654_n4888# 1.67079f
C122 minus.n45 a_n3654_n4888# 0.630397f
C123 minus.t22 a_n3654_n4888# 1.67079f
C124 minus.n46 a_n3654_n4888# 0.630416f
C125 minus.n47 a_n3654_n4888# 0.21194f
C126 minus.n48 a_n3654_n4888# 0.049204f
C127 minus.n49 a_n3654_n4888# 0.036874f
C128 minus.t7 a_n3654_n4888# 1.67079f
C129 minus.n50 a_n3654_n4888# 0.619662f
C130 minus.n51 a_n3654_n4888# 0.008368f
C131 minus.t1 a_n3654_n4888# 1.67079f
C132 minus.n52 a_n3654_n4888# 0.619662f
C133 minus.n53 a_n3654_n4888# 0.036874f
C134 minus.n54 a_n3654_n4888# 0.049204f
C135 minus.n55 a_n3654_n4888# 0.061419f
C136 minus.t5 a_n3654_n4888# 1.67079f
C137 minus.n56 a_n3654_n4888# 0.629962f
C138 minus.t21 a_n3654_n4888# 1.67079f
C139 minus.n57 a_n3654_n4888# 0.629962f
C140 minus.n58 a_n3654_n4888# 0.008368f
C141 minus.n59 a_n3654_n4888# 0.049204f
C142 minus.n60 a_n3654_n4888# 0.036874f
C143 minus.n61 a_n3654_n4888# 0.036874f
C144 minus.n62 a_n3654_n4888# 0.008368f
C145 minus.t23 a_n3654_n4888# 1.67079f
C146 minus.n63 a_n3654_n4888# 0.619662f
C147 minus.n64 a_n3654_n4888# 0.008368f
C148 minus.n65 a_n3654_n4888# 0.049204f
C149 minus.n66 a_n3654_n4888# 0.061419f
C150 minus.n67 a_n3654_n4888# 0.061419f
C151 minus.t9 a_n3654_n4888# 1.67079f
C152 minus.n68 a_n3654_n4888# 0.629507f
C153 minus.n69 a_n3654_n4888# 0.008368f
C154 minus.t0 a_n3654_n4888# 1.67079f
C155 minus.n70 a_n3654_n4888# 0.616592f
C156 minus.n71 a_n3654_n4888# 0.254837f
C157 minus.n72 a_n3654_n4888# 2.40021f
C158 drain_left.t21 a_n3654_n4888# 0.432865f
C159 drain_left.t13 a_n3654_n4888# 0.432865f
C160 drain_left.n0 a_n3654_n4888# 3.96398f
C161 drain_left.t0 a_n3654_n4888# 0.432865f
C162 drain_left.t16 a_n3654_n4888# 0.432865f
C163 drain_left.n1 a_n3654_n4888# 3.95734f
C164 drain_left.n2 a_n3654_n4888# 0.810514f
C165 drain_left.t20 a_n3654_n4888# 0.432865f
C166 drain_left.t12 a_n3654_n4888# 0.432865f
C167 drain_left.n3 a_n3654_n4888# 3.95734f
C168 drain_left.n4 a_n3654_n4888# 0.35666f
C169 drain_left.t14 a_n3654_n4888# 0.432865f
C170 drain_left.t23 a_n3654_n4888# 0.432865f
C171 drain_left.n5 a_n3654_n4888# 3.96398f
C172 drain_left.t18 a_n3654_n4888# 0.432865f
C173 drain_left.t4 a_n3654_n4888# 0.432865f
C174 drain_left.n6 a_n3654_n4888# 3.95734f
C175 drain_left.n7 a_n3654_n4888# 0.810514f
C176 drain_left.t22 a_n3654_n4888# 0.432865f
C177 drain_left.t5 a_n3654_n4888# 0.432865f
C178 drain_left.n8 a_n3654_n4888# 3.95734f
C179 drain_left.n9 a_n3654_n4888# 0.35666f
C180 drain_left.n10 a_n3654_n4888# 2.42542f
C181 drain_left.t1 a_n3654_n4888# 0.432865f
C182 drain_left.t2 a_n3654_n4888# 0.432865f
C183 drain_left.n11 a_n3654_n4888# 3.96397f
C184 drain_left.t6 a_n3654_n4888# 0.432865f
C185 drain_left.t7 a_n3654_n4888# 0.432865f
C186 drain_left.n12 a_n3654_n4888# 3.95734f
C187 drain_left.n13 a_n3654_n4888# 0.810525f
C188 drain_left.t3 a_n3654_n4888# 0.432865f
C189 drain_left.t8 a_n3654_n4888# 0.432865f
C190 drain_left.n14 a_n3654_n4888# 3.95734f
C191 drain_left.n15 a_n3654_n4888# 0.403064f
C192 drain_left.t9 a_n3654_n4888# 0.432865f
C193 drain_left.t10 a_n3654_n4888# 0.432865f
C194 drain_left.n16 a_n3654_n4888# 3.95734f
C195 drain_left.n17 a_n3654_n4888# 0.403064f
C196 drain_left.t11 a_n3654_n4888# 0.432865f
C197 drain_left.t15 a_n3654_n4888# 0.432865f
C198 drain_left.n18 a_n3654_n4888# 3.95734f
C199 drain_left.n19 a_n3654_n4888# 0.403064f
C200 drain_left.t17 a_n3654_n4888# 0.432865f
C201 drain_left.t19 a_n3654_n4888# 0.432865f
C202 drain_left.n20 a_n3654_n4888# 3.95734f
C203 drain_left.n21 a_n3654_n4888# 0.648655f
C204 source.t35 a_n3654_n4888# 4.25525f
C205 source.n0 a_n3654_n4888# 1.86146f
C206 source.t39 a_n3654_n4888# 0.372341f
C207 source.t29 a_n3654_n4888# 0.372341f
C208 source.n1 a_n3654_n4888# 3.32888f
C209 source.n2 a_n3654_n4888# 0.389817f
C210 source.t40 a_n3654_n4888# 0.372341f
C211 source.t25 a_n3654_n4888# 0.372341f
C212 source.n3 a_n3654_n4888# 3.32888f
C213 source.n4 a_n3654_n4888# 0.389817f
C214 source.t41 a_n3654_n4888# 0.372341f
C215 source.t42 a_n3654_n4888# 0.372341f
C216 source.n5 a_n3654_n4888# 3.32888f
C217 source.n6 a_n3654_n4888# 0.389817f
C218 source.t43 a_n3654_n4888# 0.372341f
C219 source.t32 a_n3654_n4888# 0.372341f
C220 source.n7 a_n3654_n4888# 3.32888f
C221 source.n8 a_n3654_n4888# 0.389817f
C222 source.t31 a_n3654_n4888# 0.372341f
C223 source.t24 a_n3654_n4888# 0.372341f
C224 source.n9 a_n3654_n4888# 3.32888f
C225 source.n10 a_n3654_n4888# 0.389817f
C226 source.t21 a_n3654_n4888# 4.25526f
C227 source.n11 a_n3654_n4888# 0.440633f
C228 source.t7 a_n3654_n4888# 4.25526f
C229 source.n12 a_n3654_n4888# 0.440633f
C230 source.t45 a_n3654_n4888# 0.372341f
C231 source.t4 a_n3654_n4888# 0.372341f
C232 source.n13 a_n3654_n4888# 3.32888f
C233 source.n14 a_n3654_n4888# 0.389817f
C234 source.t17 a_n3654_n4888# 0.372341f
C235 source.t19 a_n3654_n4888# 0.372341f
C236 source.n15 a_n3654_n4888# 3.32888f
C237 source.n16 a_n3654_n4888# 0.389817f
C238 source.t44 a_n3654_n4888# 0.372341f
C239 source.t10 a_n3654_n4888# 0.372341f
C240 source.n17 a_n3654_n4888# 3.32888f
C241 source.n18 a_n3654_n4888# 0.389817f
C242 source.t13 a_n3654_n4888# 0.372341f
C243 source.t1 a_n3654_n4888# 0.372341f
C244 source.n19 a_n3654_n4888# 3.32888f
C245 source.n20 a_n3654_n4888# 0.389817f
C246 source.t0 a_n3654_n4888# 0.372341f
C247 source.t47 a_n3654_n4888# 0.372341f
C248 source.n21 a_n3654_n4888# 3.32888f
C249 source.n22 a_n3654_n4888# 0.389817f
C250 source.t46 a_n3654_n4888# 4.25526f
C251 source.n23 a_n3654_n4888# 2.29284f
C252 source.t36 a_n3654_n4888# 4.25524f
C253 source.n24 a_n3654_n4888# 2.29286f
C254 source.t22 a_n3654_n4888# 0.372341f
C255 source.t20 a_n3654_n4888# 0.372341f
C256 source.n25 a_n3654_n4888# 3.32889f
C257 source.n26 a_n3654_n4888# 0.38981f
C258 source.t28 a_n3654_n4888# 0.372341f
C259 source.t23 a_n3654_n4888# 0.372341f
C260 source.n27 a_n3654_n4888# 3.32889f
C261 source.n28 a_n3654_n4888# 0.38981f
C262 source.t26 a_n3654_n4888# 0.372341f
C263 source.t37 a_n3654_n4888# 0.372341f
C264 source.n29 a_n3654_n4888# 3.32889f
C265 source.n30 a_n3654_n4888# 0.38981f
C266 source.t34 a_n3654_n4888# 0.372341f
C267 source.t30 a_n3654_n4888# 0.372341f
C268 source.n31 a_n3654_n4888# 3.32889f
C269 source.n32 a_n3654_n4888# 0.38981f
C270 source.t33 a_n3654_n4888# 0.372341f
C271 source.t27 a_n3654_n4888# 0.372341f
C272 source.n33 a_n3654_n4888# 3.32889f
C273 source.n34 a_n3654_n4888# 0.38981f
C274 source.t38 a_n3654_n4888# 4.25524f
C275 source.n35 a_n3654_n4888# 0.440656f
C276 source.t14 a_n3654_n4888# 4.25524f
C277 source.n36 a_n3654_n4888# 0.440656f
C278 source.t5 a_n3654_n4888# 0.372341f
C279 source.t9 a_n3654_n4888# 0.372341f
C280 source.n37 a_n3654_n4888# 3.32889f
C281 source.n38 a_n3654_n4888# 0.38981f
C282 source.t15 a_n3654_n4888# 0.372341f
C283 source.t16 a_n3654_n4888# 0.372341f
C284 source.n39 a_n3654_n4888# 3.32889f
C285 source.n40 a_n3654_n4888# 0.38981f
C286 source.t8 a_n3654_n4888# 0.372341f
C287 source.t18 a_n3654_n4888# 0.372341f
C288 source.n41 a_n3654_n4888# 3.32889f
C289 source.n42 a_n3654_n4888# 0.38981f
C290 source.t6 a_n3654_n4888# 0.372341f
C291 source.t2 a_n3654_n4888# 0.372341f
C292 source.n43 a_n3654_n4888# 3.32889f
C293 source.n44 a_n3654_n4888# 0.38981f
C294 source.t11 a_n3654_n4888# 0.372341f
C295 source.t3 a_n3654_n4888# 0.372341f
C296 source.n45 a_n3654_n4888# 3.32889f
C297 source.n46 a_n3654_n4888# 0.38981f
C298 source.t12 a_n3654_n4888# 4.25524f
C299 source.n47 a_n3654_n4888# 0.599433f
C300 source.n48 a_n3654_n4888# 2.14157f
C301 plus.n0 a_n3654_n4888# 0.049583f
C302 plus.t4 a_n3654_n4888# 1.68364f
C303 plus.t6 a_n3654_n4888# 1.68364f
C304 plus.n1 a_n3654_n4888# 0.061891f
C305 plus.t8 a_n3654_n4888# 1.68364f
C306 plus.n2 a_n3654_n4888# 0.061891f
C307 plus.t12 a_n3654_n4888# 1.68364f
C308 plus.n3 a_n3654_n4888# 0.624426f
C309 plus.n4 a_n3654_n4888# 0.037158f
C310 plus.t13 a_n3654_n4888# 1.68364f
C311 plus.t14 a_n3654_n4888# 1.68364f
C312 plus.n5 a_n3654_n4888# 0.634805f
C313 plus.n6 a_n3654_n4888# 0.049583f
C314 plus.t15 a_n3654_n4888# 1.68364f
C315 plus.t20 a_n3654_n4888# 1.68364f
C316 plus.n7 a_n3654_n4888# 0.037158f
C317 plus.t16 a_n3654_n4888# 1.68364f
C318 plus.n8 a_n3654_n4888# 0.624426f
C319 plus.n9 a_n3654_n4888# 0.21357f
C320 plus.t17 a_n3654_n4888# 1.68364f
C321 plus.t21 a_n3654_n4888# 1.68364f
C322 plus.t22 a_n3654_n4888# 1.70363f
C323 plus.n10 a_n3654_n4888# 0.611102f
C324 plus.n11 a_n3654_n4888# 0.635244f
C325 plus.n12 a_n3654_n4888# 0.635263f
C326 plus.n13 a_n3654_n4888# 0.008432f
C327 plus.n14 a_n3654_n4888# 0.049583f
C328 plus.n15 a_n3654_n4888# 0.037158f
C329 plus.n16 a_n3654_n4888# 0.037158f
C330 plus.n17 a_n3654_n4888# 0.008432f
C331 plus.n18 a_n3654_n4888# 0.624426f
C332 plus.n19 a_n3654_n4888# 0.008432f
C333 plus.n20 a_n3654_n4888# 0.634805f
C334 plus.n21 a_n3654_n4888# 0.061891f
C335 plus.n22 a_n3654_n4888# 0.061891f
C336 plus.n23 a_n3654_n4888# 0.049583f
C337 plus.n24 a_n3654_n4888# 0.008432f
C338 plus.n25 a_n3654_n4888# 0.624426f
C339 plus.n26 a_n3654_n4888# 0.008432f
C340 plus.n27 a_n3654_n4888# 0.037158f
C341 plus.n28 a_n3654_n4888# 0.037158f
C342 plus.n29 a_n3654_n4888# 0.049583f
C343 plus.n30 a_n3654_n4888# 0.008432f
C344 plus.n31 a_n3654_n4888# 0.635263f
C345 plus.n32 a_n3654_n4888# 0.634347f
C346 plus.n33 a_n3654_n4888# 0.008432f
C347 plus.n34 a_n3654_n4888# 0.621333f
C348 plus.n35 a_n3654_n4888# 0.577817f
C349 plus.n36 a_n3654_n4888# 0.049583f
C350 plus.t2 a_n3654_n4888# 1.68364f
C351 plus.n37 a_n3654_n4888# 0.061891f
C352 plus.t10 a_n3654_n4888# 1.68364f
C353 plus.n38 a_n3654_n4888# 0.061891f
C354 plus.t23 a_n3654_n4888# 1.68364f
C355 plus.t7 a_n3654_n4888# 1.68364f
C356 plus.n39 a_n3654_n4888# 0.624426f
C357 plus.n40 a_n3654_n4888# 0.037158f
C358 plus.t3 a_n3654_n4888# 1.68364f
C359 plus.t11 a_n3654_n4888# 1.68364f
C360 plus.n41 a_n3654_n4888# 0.634805f
C361 plus.n42 a_n3654_n4888# 0.049583f
C362 plus.t1 a_n3654_n4888# 1.68364f
C363 plus.n43 a_n3654_n4888# 0.037158f
C364 plus.t18 a_n3654_n4888# 1.68364f
C365 plus.t5 a_n3654_n4888# 1.68364f
C366 plus.n44 a_n3654_n4888# 0.624426f
C367 plus.n45 a_n3654_n4888# 0.21357f
C368 plus.t19 a_n3654_n4888# 1.68364f
C369 plus.t0 a_n3654_n4888# 1.70363f
C370 plus.n46 a_n3654_n4888# 0.611102f
C371 plus.t9 a_n3654_n4888# 1.68364f
C372 plus.n47 a_n3654_n4888# 0.635244f
C373 plus.n48 a_n3654_n4888# 0.635263f
C374 plus.n49 a_n3654_n4888# 0.008432f
C375 plus.n50 a_n3654_n4888# 0.049583f
C376 plus.n51 a_n3654_n4888# 0.037158f
C377 plus.n52 a_n3654_n4888# 0.037158f
C378 plus.n53 a_n3654_n4888# 0.008432f
C379 plus.n54 a_n3654_n4888# 0.624426f
C380 plus.n55 a_n3654_n4888# 0.008432f
C381 plus.n56 a_n3654_n4888# 0.634805f
C382 plus.n57 a_n3654_n4888# 0.061891f
C383 plus.n58 a_n3654_n4888# 0.061891f
C384 plus.n59 a_n3654_n4888# 0.049583f
C385 plus.n60 a_n3654_n4888# 0.008432f
C386 plus.n61 a_n3654_n4888# 0.624426f
C387 plus.n62 a_n3654_n4888# 0.008432f
C388 plus.n63 a_n3654_n4888# 0.037158f
C389 plus.n64 a_n3654_n4888# 0.037158f
C390 plus.n65 a_n3654_n4888# 0.049583f
C391 plus.n66 a_n3654_n4888# 0.008432f
C392 plus.n67 a_n3654_n4888# 0.635263f
C393 plus.n68 a_n3654_n4888# 0.634347f
C394 plus.n69 a_n3654_n4888# 0.008432f
C395 plus.n70 a_n3654_n4888# 0.621333f
C396 plus.n71 a_n3654_n4888# 1.68084f
.ends

