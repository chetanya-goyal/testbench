* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t22 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X1 drain_right.t13 minus.t0 source.t13 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X2 source.t9 minus.t1 drain_right.t12 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t17 plus.t1 drain_left.t12 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 drain_right.t11 minus.t2 source.t4 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 drain_right.t10 minus.t3 source.t7 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X6 source.t16 plus.t2 drain_left.t11 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X7 drain_left.t10 plus.t3 source.t23 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X8 source.t27 plus.t4 drain_left.t9 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X9 drain_left.t8 plus.t5 source.t25 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X10 source.t10 minus.t4 drain_right.t9 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X11 source.t0 minus.t5 drain_right.t8 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X13 source.t21 plus.t6 drain_left.t7 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X14 drain_left.t6 plus.t7 source.t19 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X15 source.t11 minus.t6 drain_right.t7 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X16 drain_right.t6 minus.t7 source.t1 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X17 drain_left.t5 plus.t8 source.t15 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X18 drain_right.t5 minus.t8 source.t6 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X19 drain_right.t4 minus.t9 source.t2 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X20 a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X21 a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X22 a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X23 drain_right.t3 minus.t10 source.t3 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X24 drain_left.t4 plus.t9 source.t26 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X25 source.t20 plus.t10 drain_left.t3 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X26 source.t12 minus.t11 drain_right.t2 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X27 source.t18 plus.t11 drain_left.t2 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X28 source.t5 minus.t12 drain_right.t1 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X29 drain_right.t0 minus.t13 source.t8 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X30 drain_left.t1 plus.t12 source.t14 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X31 drain_left.t0 plus.t13 source.t24 a_n1564_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 plus.n3 plus.t7 447.312
R1 plus.n14 plus.t3 447.312
R2 plus.n19 plus.t12 447.312
R3 plus.n30 plus.t0 447.312
R4 plus.n4 plus.t4 397.651
R5 plus.n6 plus.t13 397.651
R6 plus.n1 plus.t10 397.651
R7 plus.n11 plus.t9 397.651
R8 plus.n13 plus.t6 397.651
R9 plus.n20 plus.t2 397.651
R10 plus.n22 plus.t8 397.651
R11 plus.n17 plus.t1 397.651
R12 plus.n27 plus.t5 397.651
R13 plus.n29 plus.t11 397.651
R14 plus.n3 plus.n2 161.489
R15 plus.n19 plus.n18 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n10 plus.n9 161.3
R19 plus.n12 plus.n0 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n21 plus.n18 161.3
R22 plus.n24 plus.n23 161.3
R23 plus.n26 plus.n25 161.3
R24 plus.n28 plus.n16 161.3
R25 plus.n31 plus.n30 161.3
R26 plus.n5 plus.n4 45.2793
R27 plus.n13 plus.n12 45.2793
R28 plus.n29 plus.n28 45.2793
R29 plus.n21 plus.n20 45.2793
R30 plus.n7 plus.n6 40.8975
R31 plus.n11 plus.n10 40.8975
R32 plus.n27 plus.n26 40.8975
R33 plus.n23 plus.n22 40.8975
R34 plus.n7 plus.n1 36.5157
R35 plus.n10 plus.n1 36.5157
R36 plus.n26 plus.n17 36.5157
R37 plus.n23 plus.n17 36.5157
R38 plus.n6 plus.n5 32.1338
R39 plus.n12 plus.n11 32.1338
R40 plus.n28 plus.n27 32.1338
R41 plus.n22 plus.n21 32.1338
R42 plus.n4 plus.n3 27.752
R43 plus.n14 plus.n13 27.752
R44 plus.n30 plus.n29 27.752
R45 plus.n20 plus.n19 27.752
R46 plus plus.n31 25.0994
R47 plus plus.n15 8.31679
R48 plus.n8 plus.n2 0.189894
R49 plus.n9 plus.n8 0.189894
R50 plus.n9 plus.n0 0.189894
R51 plus.n15 plus.n0 0.189894
R52 plus.n31 plus.n16 0.189894
R53 plus.n25 plus.n16 0.189894
R54 plus.n25 plus.n24 0.189894
R55 plus.n24 plus.n18 0.189894
R56 source.n50 source.n48 289.615
R57 source.n36 source.n34 289.615
R58 source.n2 source.n0 289.615
R59 source.n16 source.n14 289.615
R60 source.n51 source.n50 185
R61 source.n37 source.n36 185
R62 source.n3 source.n2 185
R63 source.n17 source.n16 185
R64 source.t3 source.n49 167.117
R65 source.t14 source.n35 167.117
R66 source.t23 source.n1 167.117
R67 source.t6 source.n15 167.117
R68 source.n9 source.n8 84.1169
R69 source.n11 source.n10 84.1169
R70 source.n13 source.n12 84.1169
R71 source.n23 source.n22 84.1169
R72 source.n25 source.n24 84.1169
R73 source.n27 source.n26 84.1169
R74 source.n47 source.n46 84.1168
R75 source.n45 source.n44 84.1168
R76 source.n43 source.n42 84.1168
R77 source.n33 source.n32 84.1168
R78 source.n31 source.n30 84.1168
R79 source.n29 source.n28 84.1168
R80 source.n50 source.t3 52.3082
R81 source.n36 source.t14 52.3082
R82 source.n2 source.t23 52.3082
R83 source.n16 source.t6 52.3082
R84 source.n55 source.n54 31.4096
R85 source.n41 source.n40 31.4096
R86 source.n7 source.n6 31.4096
R87 source.n21 source.n20 31.4096
R88 source.n29 source.n27 14.6258
R89 source.n46 source.t13 9.9005
R90 source.n46 source.t11 9.9005
R91 source.n44 source.t1 9.9005
R92 source.n44 source.t12 9.9005
R93 source.n42 source.t8 9.9005
R94 source.n42 source.t9 9.9005
R95 source.n32 source.t15 9.9005
R96 source.n32 source.t16 9.9005
R97 source.n30 source.t25 9.9005
R98 source.n30 source.t17 9.9005
R99 source.n28 source.t22 9.9005
R100 source.n28 source.t18 9.9005
R101 source.n8 source.t26 9.9005
R102 source.n8 source.t21 9.9005
R103 source.n10 source.t24 9.9005
R104 source.n10 source.t20 9.9005
R105 source.n12 source.t19 9.9005
R106 source.n12 source.t27 9.9005
R107 source.n22 source.t4 9.9005
R108 source.n22 source.t0 9.9005
R109 source.n24 source.t2 9.9005
R110 source.n24 source.t5 9.9005
R111 source.n26 source.t7 9.9005
R112 source.n26 source.t10 9.9005
R113 source.n51 source.n49 9.71174
R114 source.n37 source.n35 9.71174
R115 source.n3 source.n1 9.71174
R116 source.n17 source.n15 9.71174
R117 source.n54 source.n53 9.45567
R118 source.n40 source.n39 9.45567
R119 source.n6 source.n5 9.45567
R120 source.n20 source.n19 9.45567
R121 source.n53 source.n52 9.3005
R122 source.n39 source.n38 9.3005
R123 source.n5 source.n4 9.3005
R124 source.n19 source.n18 9.3005
R125 source.n56 source.n7 8.67749
R126 source.n54 source.n48 8.14595
R127 source.n40 source.n34 8.14595
R128 source.n6 source.n0 8.14595
R129 source.n20 source.n14 8.14595
R130 source.n52 source.n51 7.3702
R131 source.n38 source.n37 7.3702
R132 source.n4 source.n3 7.3702
R133 source.n18 source.n17 7.3702
R134 source.n52 source.n48 5.81868
R135 source.n38 source.n34 5.81868
R136 source.n4 source.n0 5.81868
R137 source.n18 source.n14 5.81868
R138 source.n56 source.n55 5.49188
R139 source.n53 source.n49 3.44771
R140 source.n39 source.n35 3.44771
R141 source.n5 source.n1 3.44771
R142 source.n19 source.n15 3.44771
R143 source.n21 source.n13 0.698776
R144 source.n43 source.n41 0.698776
R145 source.n27 source.n25 0.457397
R146 source.n25 source.n23 0.457397
R147 source.n23 source.n21 0.457397
R148 source.n13 source.n11 0.457397
R149 source.n11 source.n9 0.457397
R150 source.n9 source.n7 0.457397
R151 source.n31 source.n29 0.457397
R152 source.n33 source.n31 0.457397
R153 source.n41 source.n33 0.457397
R154 source.n45 source.n43 0.457397
R155 source.n47 source.n45 0.457397
R156 source.n55 source.n47 0.457397
R157 source source.n56 0.188
R158 drain_left.n2 drain_left.n0 289.615
R159 drain_left.n15 drain_left.n13 289.615
R160 drain_left.n3 drain_left.n2 185
R161 drain_left.n16 drain_left.n15 185
R162 drain_left.t13 drain_left.n1 167.117
R163 drain_left.t6 drain_left.n14 167.117
R164 drain_left.n11 drain_left.n9 101.252
R165 drain_left.n25 drain_left.n24 100.796
R166 drain_left.n23 drain_left.n22 100.796
R167 drain_left.n21 drain_left.n20 100.796
R168 drain_left.n11 drain_left.n10 100.796
R169 drain_left.n8 drain_left.n7 100.796
R170 drain_left.n2 drain_left.t13 52.3082
R171 drain_left.n15 drain_left.t6 52.3082
R172 drain_left.n8 drain_left.n6 48.5453
R173 drain_left.n21 drain_left.n19 48.5453
R174 drain_left drain_left.n12 22.4185
R175 drain_left.n9 drain_left.t11 9.9005
R176 drain_left.n9 drain_left.t1 9.9005
R177 drain_left.n10 drain_left.t12 9.9005
R178 drain_left.n10 drain_left.t5 9.9005
R179 drain_left.n7 drain_left.t2 9.9005
R180 drain_left.n7 drain_left.t8 9.9005
R181 drain_left.n24 drain_left.t7 9.9005
R182 drain_left.n24 drain_left.t10 9.9005
R183 drain_left.n22 drain_left.t3 9.9005
R184 drain_left.n22 drain_left.t4 9.9005
R185 drain_left.n20 drain_left.t9 9.9005
R186 drain_left.n20 drain_left.t0 9.9005
R187 drain_left.n3 drain_left.n1 9.71174
R188 drain_left.n16 drain_left.n14 9.71174
R189 drain_left.n6 drain_left.n5 9.45567
R190 drain_left.n19 drain_left.n18 9.45567
R191 drain_left.n5 drain_left.n4 9.3005
R192 drain_left.n18 drain_left.n17 9.3005
R193 drain_left.n6 drain_left.n0 8.14595
R194 drain_left.n19 drain_left.n13 8.14595
R195 drain_left.n4 drain_left.n3 7.3702
R196 drain_left.n17 drain_left.n16 7.3702
R197 drain_left drain_left.n25 6.11011
R198 drain_left.n4 drain_left.n0 5.81868
R199 drain_left.n17 drain_left.n13 5.81868
R200 drain_left.n5 drain_left.n1 3.44771
R201 drain_left.n18 drain_left.n14 3.44771
R202 drain_left.n23 drain_left.n21 0.457397
R203 drain_left.n25 drain_left.n23 0.457397
R204 drain_left.n12 drain_left.n8 0.287826
R205 drain_left.n12 drain_left.n11 0.0593781
R206 minus.n14 minus.t3 447.312
R207 minus.n3 minus.t8 447.312
R208 minus.n30 minus.t10 447.312
R209 minus.n19 minus.t13 447.312
R210 minus.n13 minus.t4 397.651
R211 minus.n11 minus.t9 397.651
R212 minus.n1 minus.t12 397.651
R213 minus.n6 minus.t2 397.651
R214 minus.n4 minus.t5 397.651
R215 minus.n29 minus.t6 397.651
R216 minus.n27 minus.t0 397.651
R217 minus.n17 minus.t11 397.651
R218 minus.n22 minus.t7 397.651
R219 minus.n20 minus.t1 397.651
R220 minus.n3 minus.n2 161.489
R221 minus.n19 minus.n18 161.489
R222 minus.n15 minus.n14 161.3
R223 minus.n12 minus.n0 161.3
R224 minus.n10 minus.n9 161.3
R225 minus.n8 minus.n7 161.3
R226 minus.n5 minus.n2 161.3
R227 minus.n31 minus.n30 161.3
R228 minus.n28 minus.n16 161.3
R229 minus.n26 minus.n25 161.3
R230 minus.n24 minus.n23 161.3
R231 minus.n21 minus.n18 161.3
R232 minus.n13 minus.n12 45.2793
R233 minus.n5 minus.n4 45.2793
R234 minus.n21 minus.n20 45.2793
R235 minus.n29 minus.n28 45.2793
R236 minus.n11 minus.n10 40.8975
R237 minus.n7 minus.n6 40.8975
R238 minus.n23 minus.n22 40.8975
R239 minus.n27 minus.n26 40.8975
R240 minus.n10 minus.n1 36.5157
R241 minus.n7 minus.n1 36.5157
R242 minus.n23 minus.n17 36.5157
R243 minus.n26 minus.n17 36.5157
R244 minus.n12 minus.n11 32.1338
R245 minus.n6 minus.n5 32.1338
R246 minus.n22 minus.n21 32.1338
R247 minus.n28 minus.n27 32.1338
R248 minus.n14 minus.n13 27.752
R249 minus.n4 minus.n3 27.752
R250 minus.n20 minus.n19 27.752
R251 minus.n30 minus.n29 27.752
R252 minus.n32 minus.n15 27.4304
R253 minus.n32 minus.n31 6.46073
R254 minus.n15 minus.n0 0.189894
R255 minus.n9 minus.n0 0.189894
R256 minus.n9 minus.n8 0.189894
R257 minus.n8 minus.n2 0.189894
R258 minus.n24 minus.n18 0.189894
R259 minus.n25 minus.n24 0.189894
R260 minus.n25 minus.n16 0.189894
R261 minus.n31 minus.n16 0.189894
R262 minus minus.n32 0.188
R263 drain_right.n2 drain_right.n0 289.615
R264 drain_right.n20 drain_right.n18 289.615
R265 drain_right.n3 drain_right.n2 185
R266 drain_right.n21 drain_right.n20 185
R267 drain_right.t0 drain_right.n1 167.117
R268 drain_right.t10 drain_right.n19 167.117
R269 drain_right.n15 drain_right.n13 101.252
R270 drain_right.n11 drain_right.n9 101.252
R271 drain_right.n15 drain_right.n14 100.796
R272 drain_right.n17 drain_right.n16 100.796
R273 drain_right.n11 drain_right.n10 100.796
R274 drain_right.n8 drain_right.n7 100.796
R275 drain_right.n2 drain_right.t0 52.3082
R276 drain_right.n20 drain_right.t10 52.3082
R277 drain_right.n8 drain_right.n6 48.5453
R278 drain_right.n25 drain_right.n24 48.0884
R279 drain_right drain_right.n12 21.8652
R280 drain_right.n9 drain_right.t7 9.9005
R281 drain_right.n9 drain_right.t3 9.9005
R282 drain_right.n10 drain_right.t2 9.9005
R283 drain_right.n10 drain_right.t13 9.9005
R284 drain_right.n7 drain_right.t12 9.9005
R285 drain_right.n7 drain_right.t6 9.9005
R286 drain_right.n13 drain_right.t8 9.9005
R287 drain_right.n13 drain_right.t5 9.9005
R288 drain_right.n14 drain_right.t1 9.9005
R289 drain_right.n14 drain_right.t11 9.9005
R290 drain_right.n16 drain_right.t9 9.9005
R291 drain_right.n16 drain_right.t4 9.9005
R292 drain_right.n3 drain_right.n1 9.71174
R293 drain_right.n21 drain_right.n19 9.71174
R294 drain_right.n6 drain_right.n5 9.45567
R295 drain_right.n24 drain_right.n23 9.45567
R296 drain_right.n5 drain_right.n4 9.3005
R297 drain_right.n23 drain_right.n22 9.3005
R298 drain_right.n6 drain_right.n0 8.14595
R299 drain_right.n24 drain_right.n18 8.14595
R300 drain_right.n4 drain_right.n3 7.3702
R301 drain_right.n22 drain_right.n21 7.3702
R302 drain_right drain_right.n25 5.88166
R303 drain_right.n4 drain_right.n0 5.81868
R304 drain_right.n22 drain_right.n18 5.81868
R305 drain_right.n5 drain_right.n1 3.44771
R306 drain_right.n23 drain_right.n19 3.44771
R307 drain_right.n25 drain_right.n17 0.457397
R308 drain_right.n17 drain_right.n15 0.457397
R309 drain_right.n12 drain_right.n8 0.287826
R310 drain_right.n12 drain_right.n11 0.0593781
C0 drain_left plus 1.19378f
C1 source minus 1.15225f
C2 plus minus 3.26097f
C3 source drain_right 7.69488f
C4 drain_right plus 0.311104f
C5 drain_left minus 0.177298f
C6 drain_left drain_right 0.79113f
C7 source plus 1.16633f
C8 drain_right minus 1.04427f
C9 source drain_left 7.69807f
C10 drain_right a_n1564_n1288# 3.91448f
C11 drain_left a_n1564_n1288# 4.14639f
C12 source a_n1564_n1288# 2.479108f
C13 minus a_n1564_n1288# 5.254964f
C14 plus a_n1564_n1288# 5.950367f
C15 drain_right.n0 a_n1564_n1288# 0.041484f
C16 drain_right.n1 a_n1564_n1288# 0.091789f
C17 drain_right.t0 a_n1564_n1288# 0.068883f
C18 drain_right.n2 a_n1564_n1288# 0.071838f
C19 drain_right.n3 a_n1564_n1288# 0.023158f
C20 drain_right.n4 a_n1564_n1288# 0.015273f
C21 drain_right.n5 a_n1564_n1288# 0.202326f
C22 drain_right.n6 a_n1564_n1288# 0.066015f
C23 drain_right.t12 a_n1564_n1288# 0.044921f
C24 drain_right.t6 a_n1564_n1288# 0.044921f
C25 drain_right.n7 a_n1564_n1288# 0.282205f
C26 drain_right.n8 a_n1564_n1288# 0.382779f
C27 drain_right.t7 a_n1564_n1288# 0.044921f
C28 drain_right.t3 a_n1564_n1288# 0.044921f
C29 drain_right.n9 a_n1564_n1288# 0.283616f
C30 drain_right.t2 a_n1564_n1288# 0.044921f
C31 drain_right.t13 a_n1564_n1288# 0.044921f
C32 drain_right.n10 a_n1564_n1288# 0.282205f
C33 drain_right.n11 a_n1564_n1288# 0.58724f
C34 drain_right.n12 a_n1564_n1288# 0.663077f
C35 drain_right.t8 a_n1564_n1288# 0.044921f
C36 drain_right.t5 a_n1564_n1288# 0.044921f
C37 drain_right.n13 a_n1564_n1288# 0.283617f
C38 drain_right.t1 a_n1564_n1288# 0.044921f
C39 drain_right.t11 a_n1564_n1288# 0.044921f
C40 drain_right.n14 a_n1564_n1288# 0.282206f
C41 drain_right.n15 a_n1564_n1288# 0.612498f
C42 drain_right.t9 a_n1564_n1288# 0.044921f
C43 drain_right.t4 a_n1564_n1288# 0.044921f
C44 drain_right.n16 a_n1564_n1288# 0.282206f
C45 drain_right.n17 a_n1564_n1288# 0.30123f
C46 drain_right.n18 a_n1564_n1288# 0.041484f
C47 drain_right.n19 a_n1564_n1288# 0.091789f
C48 drain_right.t10 a_n1564_n1288# 0.068883f
C49 drain_right.n20 a_n1564_n1288# 0.071838f
C50 drain_right.n21 a_n1564_n1288# 0.023158f
C51 drain_right.n22 a_n1564_n1288# 0.015273f
C52 drain_right.n23 a_n1564_n1288# 0.202326f
C53 drain_right.n24 a_n1564_n1288# 0.065114f
C54 drain_right.n25 a_n1564_n1288# 0.326696f
C55 minus.n0 a_n1564_n1288# 0.032672f
C56 minus.t3 a_n1564_n1288# 0.0419f
C57 minus.t4 a_n1564_n1288# 0.038456f
C58 minus.t9 a_n1564_n1288# 0.038456f
C59 minus.t12 a_n1564_n1288# 0.038456f
C60 minus.n1 a_n1564_n1288# 0.030215f
C61 minus.n2 a_n1564_n1288# 0.07295f
C62 minus.t2 a_n1564_n1288# 0.038456f
C63 minus.t5 a_n1564_n1288# 0.038456f
C64 minus.t8 a_n1564_n1288# 0.0419f
C65 minus.n3 a_n1564_n1288# 0.039067f
C66 minus.n4 a_n1564_n1288# 0.030215f
C67 minus.n5 a_n1564_n1288# 0.011443f
C68 minus.n6 a_n1564_n1288# 0.030215f
C69 minus.n7 a_n1564_n1288# 0.011443f
C70 minus.n8 a_n1564_n1288# 0.032672f
C71 minus.n9 a_n1564_n1288# 0.032672f
C72 minus.n10 a_n1564_n1288# 0.011443f
C73 minus.n11 a_n1564_n1288# 0.030215f
C74 minus.n12 a_n1564_n1288# 0.011443f
C75 minus.n13 a_n1564_n1288# 0.030215f
C76 minus.n14 a_n1564_n1288# 0.039019f
C77 minus.n15 a_n1564_n1288# 0.72547f
C78 minus.n16 a_n1564_n1288# 0.032672f
C79 minus.t6 a_n1564_n1288# 0.038456f
C80 minus.t0 a_n1564_n1288# 0.038456f
C81 minus.t11 a_n1564_n1288# 0.038456f
C82 minus.n17 a_n1564_n1288# 0.030215f
C83 minus.n18 a_n1564_n1288# 0.07295f
C84 minus.t7 a_n1564_n1288# 0.038456f
C85 minus.t1 a_n1564_n1288# 0.038456f
C86 minus.t13 a_n1564_n1288# 0.0419f
C87 minus.n19 a_n1564_n1288# 0.039067f
C88 minus.n20 a_n1564_n1288# 0.030215f
C89 minus.n21 a_n1564_n1288# 0.011443f
C90 minus.n22 a_n1564_n1288# 0.030215f
C91 minus.n23 a_n1564_n1288# 0.011443f
C92 minus.n24 a_n1564_n1288# 0.032672f
C93 minus.n25 a_n1564_n1288# 0.032672f
C94 minus.n26 a_n1564_n1288# 0.011443f
C95 minus.n27 a_n1564_n1288# 0.030215f
C96 minus.n28 a_n1564_n1288# 0.011443f
C97 minus.n29 a_n1564_n1288# 0.030215f
C98 minus.t10 a_n1564_n1288# 0.0419f
C99 minus.n30 a_n1564_n1288# 0.039019f
C100 minus.n31 a_n1564_n1288# 0.21057f
C101 minus.n32 a_n1564_n1288# 0.898554f
C102 drain_left.n0 a_n1564_n1288# 0.040894f
C103 drain_left.n1 a_n1564_n1288# 0.090483f
C104 drain_left.t13 a_n1564_n1288# 0.067903f
C105 drain_left.n2 a_n1564_n1288# 0.070815f
C106 drain_left.n3 a_n1564_n1288# 0.022828f
C107 drain_left.n4 a_n1564_n1288# 0.015056f
C108 drain_left.n5 a_n1564_n1288# 0.199446f
C109 drain_left.n6 a_n1564_n1288# 0.065075f
C110 drain_left.t2 a_n1564_n1288# 0.044281f
C111 drain_left.t8 a_n1564_n1288# 0.044281f
C112 drain_left.n7 a_n1564_n1288# 0.278188f
C113 drain_left.n8 a_n1564_n1288# 0.377331f
C114 drain_left.t11 a_n1564_n1288# 0.044281f
C115 drain_left.t1 a_n1564_n1288# 0.044281f
C116 drain_left.n9 a_n1564_n1288# 0.279579f
C117 drain_left.t12 a_n1564_n1288# 0.044281f
C118 drain_left.t5 a_n1564_n1288# 0.044281f
C119 drain_left.n10 a_n1564_n1288# 0.278188f
C120 drain_left.n11 a_n1564_n1288# 0.578881f
C121 drain_left.n12 a_n1564_n1288# 0.708679f
C122 drain_left.n13 a_n1564_n1288# 0.040894f
C123 drain_left.n14 a_n1564_n1288# 0.090483f
C124 drain_left.t6 a_n1564_n1288# 0.067903f
C125 drain_left.n15 a_n1564_n1288# 0.070815f
C126 drain_left.n16 a_n1564_n1288# 0.022828f
C127 drain_left.n17 a_n1564_n1288# 0.015056f
C128 drain_left.n18 a_n1564_n1288# 0.199446f
C129 drain_left.n19 a_n1564_n1288# 0.065075f
C130 drain_left.t9 a_n1564_n1288# 0.044281f
C131 drain_left.t0 a_n1564_n1288# 0.044281f
C132 drain_left.n20 a_n1564_n1288# 0.278189f
C133 drain_left.n21 a_n1564_n1288# 0.390378f
C134 drain_left.t3 a_n1564_n1288# 0.044281f
C135 drain_left.t4 a_n1564_n1288# 0.044281f
C136 drain_left.n22 a_n1564_n1288# 0.278189f
C137 drain_left.n23 a_n1564_n1288# 0.296943f
C138 drain_left.t7 a_n1564_n1288# 0.044281f
C139 drain_left.t10 a_n1564_n1288# 0.044281f
C140 drain_left.n24 a_n1564_n1288# 0.278189f
C141 drain_left.n25 a_n1564_n1288# 0.526243f
C142 source.n0 a_n1564_n1288# 0.049871f
C143 source.n1 a_n1564_n1288# 0.110347f
C144 source.t23 a_n1564_n1288# 0.082809f
C145 source.n2 a_n1564_n1288# 0.086361f
C146 source.n3 a_n1564_n1288# 0.02784f
C147 source.n4 a_n1564_n1288# 0.018361f
C148 source.n5 a_n1564_n1288# 0.243231f
C149 source.n6 a_n1564_n1288# 0.054671f
C150 source.n7 a_n1564_n1288# 0.499012f
C151 source.t26 a_n1564_n1288# 0.054002f
C152 source.t21 a_n1564_n1288# 0.054002f
C153 source.n8 a_n1564_n1288# 0.288695f
C154 source.n9 a_n1564_n1288# 0.366254f
C155 source.t24 a_n1564_n1288# 0.054002f
C156 source.t20 a_n1564_n1288# 0.054002f
C157 source.n10 a_n1564_n1288# 0.288695f
C158 source.n11 a_n1564_n1288# 0.366254f
C159 source.t19 a_n1564_n1288# 0.054002f
C160 source.t27 a_n1564_n1288# 0.054002f
C161 source.n12 a_n1564_n1288# 0.288695f
C162 source.n13 a_n1564_n1288# 0.39283f
C163 source.n14 a_n1564_n1288# 0.049871f
C164 source.n15 a_n1564_n1288# 0.110346f
C165 source.t6 a_n1564_n1288# 0.082809f
C166 source.n16 a_n1564_n1288# 0.086361f
C167 source.n17 a_n1564_n1288# 0.02784f
C168 source.n18 a_n1564_n1288# 0.018361f
C169 source.n19 a_n1564_n1288# 0.243231f
C170 source.n20 a_n1564_n1288# 0.054671f
C171 source.n21 a_n1564_n1288# 0.155313f
C172 source.t4 a_n1564_n1288# 0.054002f
C173 source.t0 a_n1564_n1288# 0.054002f
C174 source.n22 a_n1564_n1288# 0.288695f
C175 source.n23 a_n1564_n1288# 0.366254f
C176 source.t2 a_n1564_n1288# 0.054002f
C177 source.t5 a_n1564_n1288# 0.054002f
C178 source.n24 a_n1564_n1288# 0.288695f
C179 source.n25 a_n1564_n1288# 0.366254f
C180 source.t7 a_n1564_n1288# 0.054002f
C181 source.t10 a_n1564_n1288# 0.054002f
C182 source.n26 a_n1564_n1288# 0.288695f
C183 source.n27 a_n1564_n1288# 1.10329f
C184 source.t22 a_n1564_n1288# 0.054002f
C185 source.t18 a_n1564_n1288# 0.054002f
C186 source.n28 a_n1564_n1288# 0.288693f
C187 source.n29 a_n1564_n1288# 1.10329f
C188 source.t25 a_n1564_n1288# 0.054002f
C189 source.t17 a_n1564_n1288# 0.054002f
C190 source.n30 a_n1564_n1288# 0.288693f
C191 source.n31 a_n1564_n1288# 0.366256f
C192 source.t15 a_n1564_n1288# 0.054002f
C193 source.t16 a_n1564_n1288# 0.054002f
C194 source.n32 a_n1564_n1288# 0.288693f
C195 source.n33 a_n1564_n1288# 0.366256f
C196 source.n34 a_n1564_n1288# 0.049871f
C197 source.n35 a_n1564_n1288# 0.110346f
C198 source.t14 a_n1564_n1288# 0.082809f
C199 source.n36 a_n1564_n1288# 0.086361f
C200 source.n37 a_n1564_n1288# 0.02784f
C201 source.n38 a_n1564_n1288# 0.018361f
C202 source.n39 a_n1564_n1288# 0.243231f
C203 source.n40 a_n1564_n1288# 0.054671f
C204 source.n41 a_n1564_n1288# 0.155313f
C205 source.t8 a_n1564_n1288# 0.054002f
C206 source.t9 a_n1564_n1288# 0.054002f
C207 source.n42 a_n1564_n1288# 0.288693f
C208 source.n43 a_n1564_n1288# 0.392832f
C209 source.t1 a_n1564_n1288# 0.054002f
C210 source.t12 a_n1564_n1288# 0.054002f
C211 source.n44 a_n1564_n1288# 0.288693f
C212 source.n45 a_n1564_n1288# 0.366256f
C213 source.t13 a_n1564_n1288# 0.054002f
C214 source.t11 a_n1564_n1288# 0.054002f
C215 source.n46 a_n1564_n1288# 0.288693f
C216 source.n47 a_n1564_n1288# 0.366256f
C217 source.n48 a_n1564_n1288# 0.049871f
C218 source.n49 a_n1564_n1288# 0.110346f
C219 source.t3 a_n1564_n1288# 0.082809f
C220 source.n50 a_n1564_n1288# 0.086361f
C221 source.n51 a_n1564_n1288# 0.02784f
C222 source.n52 a_n1564_n1288# 0.018361f
C223 source.n53 a_n1564_n1288# 0.243231f
C224 source.n54 a_n1564_n1288# 0.054671f
C225 source.n55 a_n1564_n1288# 0.315434f
C226 source.n56 a_n1564_n1288# 0.840789f
C227 plus.n0 a_n1564_n1288# 0.033339f
C228 plus.t6 a_n1564_n1288# 0.039241f
C229 plus.t9 a_n1564_n1288# 0.039241f
C230 plus.t10 a_n1564_n1288# 0.039241f
C231 plus.n1 a_n1564_n1288# 0.030832f
C232 plus.n2 a_n1564_n1288# 0.074441f
C233 plus.t13 a_n1564_n1288# 0.039241f
C234 plus.t4 a_n1564_n1288# 0.039241f
C235 plus.t7 a_n1564_n1288# 0.042756f
C236 plus.n3 a_n1564_n1288# 0.039865f
C237 plus.n4 a_n1564_n1288# 0.030832f
C238 plus.n5 a_n1564_n1288# 0.011676f
C239 plus.n6 a_n1564_n1288# 0.030832f
C240 plus.n7 a_n1564_n1288# 0.011676f
C241 plus.n8 a_n1564_n1288# 0.033339f
C242 plus.n9 a_n1564_n1288# 0.033339f
C243 plus.n10 a_n1564_n1288# 0.011676f
C244 plus.n11 a_n1564_n1288# 0.030832f
C245 plus.n12 a_n1564_n1288# 0.011676f
C246 plus.n13 a_n1564_n1288# 0.030832f
C247 plus.t3 a_n1564_n1288# 0.042756f
C248 plus.n14 a_n1564_n1288# 0.039817f
C249 plus.n15 a_n1564_n1288# 0.235082f
C250 plus.n16 a_n1564_n1288# 0.033339f
C251 plus.t0 a_n1564_n1288# 0.042756f
C252 plus.t11 a_n1564_n1288# 0.039241f
C253 plus.t5 a_n1564_n1288# 0.039241f
C254 plus.t1 a_n1564_n1288# 0.039241f
C255 plus.n17 a_n1564_n1288# 0.030832f
C256 plus.n18 a_n1564_n1288# 0.074441f
C257 plus.t8 a_n1564_n1288# 0.039241f
C258 plus.t2 a_n1564_n1288# 0.039241f
C259 plus.t12 a_n1564_n1288# 0.042756f
C260 plus.n19 a_n1564_n1288# 0.039865f
C261 plus.n20 a_n1564_n1288# 0.030832f
C262 plus.n21 a_n1564_n1288# 0.011676f
C263 plus.n22 a_n1564_n1288# 0.030832f
C264 plus.n23 a_n1564_n1288# 0.011676f
C265 plus.n24 a_n1564_n1288# 0.033339f
C266 plus.n25 a_n1564_n1288# 0.033339f
C267 plus.n26 a_n1564_n1288# 0.011676f
C268 plus.n27 a_n1564_n1288# 0.030832f
C269 plus.n28 a_n1564_n1288# 0.011676f
C270 plus.n29 a_n1564_n1288# 0.030832f
C271 plus.n30 a_n1564_n1288# 0.039817f
C272 plus.n31 a_n1564_n1288# 0.708727f
.ends

