* NGSPICE file created from diffpair333.ext - technology: sky130A

.subckt diffpair333 minus drain_right drain_left source plus
X0 source.t13 minus.t0 drain_right.t3 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 source.t12 minus.t1 drain_right.t5 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 drain_right.t0 minus.t2 source.t11 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X3 drain_right.t2 minus.t3 source.t10 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X4 drain_right.t4 minus.t4 source.t9 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X6 drain_left.t7 plus.t0 source.t14 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X7 a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X8 a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X9 source.t8 minus.t5 drain_right.t7 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X10 source.t3 plus.t1 drain_left.t6 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X11 source.t0 plus.t2 drain_left.t5 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X12 a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X13 drain_right.t6 minus.t6 source.t7 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X14 drain_left.t4 plus.t3 source.t15 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X15 drain_left.t3 plus.t4 source.t1 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X16 drain_left.t2 plus.t5 source.t2 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X17 source.t5 plus.t6 drain_left.t1 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X18 source.t6 minus.t7 drain_right.t1 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X19 source.t4 plus.t7 drain_left.t0 a_n1246_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n5 minus.t7 1284.24
R1 minus.n1 minus.t6 1284.24
R2 minus.n12 minus.t3 1284.24
R3 minus.n8 minus.t1 1284.24
R4 minus.n4 minus.t2 1241.15
R5 minus.n2 minus.t5 1241.15
R6 minus.n11 minus.t0 1241.15
R7 minus.n9 minus.t4 1241.15
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 38.7066
R15 minus.n3 minus.n2 38.7066
R16 minus.n10 minus.n9 38.7066
R17 minus.n11 minus.n10 38.7066
R18 minus.n5 minus.n4 34.3247
R19 minus.n2 minus.n1 34.3247
R20 minus.n9 minus.n8 34.3247
R21 minus.n12 minus.n11 34.3247
R22 minus.n14 minus.n6 31.5119
R23 minus.n14 minus.n13 6.44368
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 drain_right.n5 drain_right.n3 65.9943
R28 drain_right.n2 drain_right.n1 65.7104
R29 drain_right.n2 drain_right.n0 65.7104
R30 drain_right.n5 drain_right.n4 65.5376
R31 drain_right drain_right.n2 26.1403
R32 drain_right drain_right.n5 6.11011
R33 drain_right.n1 drain_right.t3 2.2005
R34 drain_right.n1 drain_right.t2 2.2005
R35 drain_right.n0 drain_right.t5 2.2005
R36 drain_right.n0 drain_right.t4 2.2005
R37 drain_right.n3 drain_right.t7 2.2005
R38 drain_right.n3 drain_right.t6 2.2005
R39 drain_right.n4 drain_right.t1 2.2005
R40 drain_right.n4 drain_right.t0 2.2005
R41 source.n3 source.t3 51.0588
R42 source.n4 source.t7 51.0588
R43 source.n7 source.t6 51.0588
R44 source.n15 source.t10 51.0586
R45 source.n12 source.t12 51.0586
R46 source.n11 source.t15 51.0586
R47 source.n8 source.t0 51.0586
R48 source.n0 source.t2 51.0586
R49 source.n2 source.n1 48.8588
R50 source.n6 source.n5 48.8588
R51 source.n14 source.n13 48.8586
R52 source.n10 source.n9 48.8586
R53 source.n8 source.n7 19.4719
R54 source.n16 source.n0 13.9805
R55 source.n16 source.n15 5.49188
R56 source.n13 source.t9 2.2005
R57 source.n13 source.t13 2.2005
R58 source.n9 source.t1 2.2005
R59 source.n9 source.t5 2.2005
R60 source.n1 source.t14 2.2005
R61 source.n1 source.t4 2.2005
R62 source.n5 source.t11 2.2005
R63 source.n5 source.t8 2.2005
R64 source.n4 source.n3 0.470328
R65 source.n12 source.n11 0.470328
R66 source.n7 source.n6 0.457397
R67 source.n6 source.n4 0.457397
R68 source.n3 source.n2 0.457397
R69 source.n2 source.n0 0.457397
R70 source.n10 source.n8 0.457397
R71 source.n11 source.n10 0.457397
R72 source.n14 source.n12 0.457397
R73 source.n15 source.n14 0.457397
R74 source source.n16 0.188
R75 plus.n1 plus.t1 1284.24
R76 plus.n5 plus.t5 1284.24
R77 plus.n8 plus.t3 1284.24
R78 plus.n12 plus.t2 1284.24
R79 plus.n2 plus.t0 1241.15
R80 plus.n4 plus.t7 1241.15
R81 plus.n9 plus.t6 1241.15
R82 plus.n11 plus.t4 1241.15
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 38.7066
R90 plus.n4 plus.n3 38.7066
R91 plus.n11 plus.n10 38.7066
R92 plus.n10 plus.n9 38.7066
R93 plus.n2 plus.n1 34.3247
R94 plus.n5 plus.n4 34.3247
R95 plus.n12 plus.n11 34.3247
R96 plus.n9 plus.n8 34.3247
R97 plus plus.n13 26.5293
R98 plus plus.n6 10.9513
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 65.9945
R102 drain_left.n2 drain_left.n1 65.7104
R103 drain_left.n2 drain_left.n0 65.7104
R104 drain_left.n5 drain_left.n4 65.5374
R105 drain_left drain_left.n2 26.6935
R106 drain_left drain_left.n5 6.11011
R107 drain_left.n1 drain_left.t1 2.2005
R108 drain_left.n1 drain_left.t4 2.2005
R109 drain_left.n0 drain_left.t5 2.2005
R110 drain_left.n0 drain_left.t3 2.2005
R111 drain_left.n4 drain_left.t0 2.2005
R112 drain_left.n4 drain_left.t2 2.2005
R113 drain_left.n3 drain_left.t6 2.2005
R114 drain_left.n3 drain_left.t7 2.2005
C0 drain_right source 15.182799f
C1 drain_right plus 0.269775f
C2 drain_right minus 2.05464f
C3 source drain_left 15.1842f
C4 drain_left plus 2.17144f
C5 drain_left minus 0.17017f
C6 source plus 1.7027f
C7 source minus 1.68866f
C8 minus plus 4.15279f
C9 drain_right drain_left 0.58123f
C10 drain_right a_n1246_n2688# 5.28044f
C11 drain_left a_n1246_n2688# 5.47136f
C12 source a_n1246_n2688# 6.764269f
C13 minus a_n1246_n2688# 4.582671f
C14 plus a_n1246_n2688# 6.04456f
C15 drain_left.t5 a_n1246_n2688# 0.261554f
C16 drain_left.t3 a_n1246_n2688# 0.261554f
C17 drain_left.n0 a_n1246_n2688# 2.28875f
C18 drain_left.t1 a_n1246_n2688# 0.261554f
C19 drain_left.t4 a_n1246_n2688# 0.261554f
C20 drain_left.n1 a_n1246_n2688# 2.28875f
C21 drain_left.n2 a_n1246_n2688# 2.09132f
C22 drain_left.t6 a_n1246_n2688# 0.261554f
C23 drain_left.t7 a_n1246_n2688# 0.261554f
C24 drain_left.n3 a_n1246_n2688# 2.29062f
C25 drain_left.t0 a_n1246_n2688# 0.261554f
C26 drain_left.t2 a_n1246_n2688# 0.261554f
C27 drain_left.n4 a_n1246_n2688# 2.28772f
C28 drain_left.n5 a_n1246_n2688# 1.11863f
C29 plus.n0 a_n1246_n2688# 0.104676f
C30 plus.t7 a_n1246_n2688# 0.245198f
C31 plus.t0 a_n1246_n2688# 0.245198f
C32 plus.t1 a_n1246_n2688# 0.248794f
C33 plus.n1 a_n1246_n2688# 0.120489f
C34 plus.n2 a_n1246_n2688# 0.10733f
C35 plus.n3 a_n1246_n2688# 0.016837f
C36 plus.n4 a_n1246_n2688# 0.10733f
C37 plus.t5 a_n1246_n2688# 0.248794f
C38 plus.n5 a_n1246_n2688# 0.120423f
C39 plus.n6 a_n1246_n2688# 0.465646f
C40 plus.n7 a_n1246_n2688# 0.104676f
C41 plus.t2 a_n1246_n2688# 0.248794f
C42 plus.t4 a_n1246_n2688# 0.245198f
C43 plus.t6 a_n1246_n2688# 0.245198f
C44 plus.t3 a_n1246_n2688# 0.248794f
C45 plus.n8 a_n1246_n2688# 0.120489f
C46 plus.n9 a_n1246_n2688# 0.10733f
C47 plus.n10 a_n1246_n2688# 0.016837f
C48 plus.n11 a_n1246_n2688# 0.10733f
C49 plus.n12 a_n1246_n2688# 0.120423f
C50 plus.n13 a_n1246_n2688# 1.18027f
C51 source.t2 a_n1246_n2688# 1.85159f
C52 source.n0 a_n1246_n2688# 1.05336f
C53 source.t14 a_n1246_n2688# 0.173639f
C54 source.t4 a_n1246_n2688# 0.173639f
C55 source.n1 a_n1246_n2688# 1.45359f
C56 source.n2 a_n1246_n2688# 0.299436f
C57 source.t3 a_n1246_n2688# 1.85159f
C58 source.n3 a_n1246_n2688# 0.376008f
C59 source.t7 a_n1246_n2688# 1.85159f
C60 source.n4 a_n1246_n2688# 0.376008f
C61 source.t11 a_n1246_n2688# 0.173639f
C62 source.t8 a_n1246_n2688# 0.173639f
C63 source.n5 a_n1246_n2688# 1.45359f
C64 source.n6 a_n1246_n2688# 0.299436f
C65 source.t6 a_n1246_n2688# 1.85159f
C66 source.n7 a_n1246_n2688# 1.40589f
C67 source.t0 a_n1246_n2688# 1.85159f
C68 source.n8 a_n1246_n2688# 1.40589f
C69 source.t1 a_n1246_n2688# 0.173639f
C70 source.t5 a_n1246_n2688# 0.173639f
C71 source.n9 a_n1246_n2688# 1.45358f
C72 source.n10 a_n1246_n2688# 0.29944f
C73 source.t15 a_n1246_n2688# 1.85159f
C74 source.n11 a_n1246_n2688# 0.376013f
C75 source.t12 a_n1246_n2688# 1.85159f
C76 source.n12 a_n1246_n2688# 0.376013f
C77 source.t9 a_n1246_n2688# 0.173639f
C78 source.t13 a_n1246_n2688# 0.173639f
C79 source.n13 a_n1246_n2688# 1.45358f
C80 source.n14 a_n1246_n2688# 0.29944f
C81 source.t10 a_n1246_n2688# 1.85159f
C82 source.n15 a_n1246_n2688# 0.508397f
C83 source.n16 a_n1246_n2688# 1.2674f
C84 drain_right.t5 a_n1246_n2688# 0.262219f
C85 drain_right.t4 a_n1246_n2688# 0.262219f
C86 drain_right.n0 a_n1246_n2688# 2.29456f
C87 drain_right.t3 a_n1246_n2688# 0.262219f
C88 drain_right.t2 a_n1246_n2688# 0.262219f
C89 drain_right.n1 a_n1246_n2688# 2.29456f
C90 drain_right.n2 a_n1246_n2688# 2.01989f
C91 drain_right.t7 a_n1246_n2688# 0.262219f
C92 drain_right.t6 a_n1246_n2688# 0.262219f
C93 drain_right.n3 a_n1246_n2688# 2.29643f
C94 drain_right.t1 a_n1246_n2688# 0.262219f
C95 drain_right.t0 a_n1246_n2688# 0.262219f
C96 drain_right.n4 a_n1246_n2688# 2.29354f
C97 drain_right.n5 a_n1246_n2688# 1.12147f
C98 minus.n0 a_n1246_n2688# 0.101499f
C99 minus.t7 a_n1246_n2688# 0.241243f
C100 minus.t2 a_n1246_n2688# 0.237756f
C101 minus.t5 a_n1246_n2688# 0.237756f
C102 minus.t6 a_n1246_n2688# 0.241243f
C103 minus.n1 a_n1246_n2688# 0.116832f
C104 minus.n2 a_n1246_n2688# 0.104072f
C105 minus.n3 a_n1246_n2688# 0.016326f
C106 minus.n4 a_n1246_n2688# 0.104072f
C107 minus.n5 a_n1246_n2688# 0.116768f
C108 minus.n6 a_n1246_n2688# 1.31515f
C109 minus.n7 a_n1246_n2688# 0.101499f
C110 minus.t0 a_n1246_n2688# 0.237756f
C111 minus.t4 a_n1246_n2688# 0.237756f
C112 minus.t1 a_n1246_n2688# 0.241243f
C113 minus.n8 a_n1246_n2688# 0.116832f
C114 minus.n9 a_n1246_n2688# 0.104072f
C115 minus.n10 a_n1246_n2688# 0.016326f
C116 minus.n11 a_n1246_n2688# 0.104072f
C117 minus.t3 a_n1246_n2688# 0.241243f
C118 minus.n12 a_n1246_n2688# 0.116768f
C119 minus.n13 a_n1246_n2688# 0.29855f
C120 minus.n14 a_n1246_n2688# 1.62055f
.ends

