* NGSPICE file created from diffpair159.ext - technology: sky130A

.subckt diffpair159 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t17 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X1 source.t6 plus.t0 drain_left.t23 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X2 drain_right.t7 minus.t1 source.t46 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 drain_right.t10 minus.t2 source.t45 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X4 source.t3 plus.t1 drain_left.t22 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X5 drain_right.t21 minus.t3 source.t44 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X6 drain_right.t3 minus.t4 source.t43 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X7 source.t10 plus.t2 drain_left.t21 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X8 source.t4 plus.t3 drain_left.t20 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X9 source.t13 plus.t4 drain_left.t19 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X10 source.t42 minus.t5 drain_right.t14 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X11 drain_right.t5 minus.t6 source.t41 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X12 drain_right.t16 minus.t7 source.t40 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X13 drain_left.t18 plus.t5 source.t1 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X14 source.t16 plus.t6 drain_left.t17 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X15 source.t23 plus.t7 drain_left.t16 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X16 drain_right.t6 minus.t8 source.t39 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X17 drain_left.t15 plus.t8 source.t14 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X18 source.t38 minus.t9 drain_right.t22 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X19 source.t37 minus.t10 drain_right.t20 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X20 a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X21 drain_right.t19 minus.t11 source.t36 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X22 drain_right.t18 minus.t12 source.t35 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X23 drain_right.t8 minus.t13 source.t34 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X24 source.t33 minus.t14 drain_right.t11 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X25 a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X26 source.t18 plus.t9 drain_left.t14 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X27 source.t32 minus.t15 drain_right.t23 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X28 source.t31 minus.t16 drain_right.t4 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X29 drain_left.t13 plus.t10 source.t22 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X30 drain_left.t12 plus.t11 source.t19 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X31 source.t30 minus.t17 drain_right.t15 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X32 drain_right.t9 minus.t18 source.t29 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X33 drain_left.t11 plus.t12 source.t17 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X34 drain_right.t0 minus.t19 source.t28 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X35 drain_left.t10 plus.t13 source.t7 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X36 source.t20 plus.t14 drain_left.t9 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X37 a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X38 source.t27 minus.t20 drain_right.t2 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X39 drain_left.t8 plus.t15 source.t21 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X40 drain_left.t7 plus.t16 source.t0 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X41 source.t26 minus.t21 drain_right.t13 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X42 source.t25 minus.t22 drain_right.t12 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X43 source.t15 plus.t17 drain_left.t6 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X44 source.t24 minus.t23 drain_right.t1 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X45 drain_left.t5 plus.t18 source.t2 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X46 source.t9 plus.t19 drain_left.t4 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X47 drain_left.t3 plus.t20 source.t12 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X48 a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X49 drain_left.t2 plus.t21 source.t5 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X50 source.t8 plus.t22 drain_left.t1 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X51 drain_left.t0 plus.t23 source.t11 a_n3654_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n35 minus.n34 161.3
R1 minus.n33 minus.n0 161.3
R2 minus.n29 minus.n28 161.3
R3 minus.n27 minus.n2 161.3
R4 minus.n26 minus.n25 161.3
R5 minus.n24 minus.n3 161.3
R6 minus.n23 minus.n22 161.3
R7 minus.n18 minus.n5 161.3
R8 minus.n17 minus.n16 161.3
R9 minus.n15 minus.n6 161.3
R10 minus.n14 minus.n13 161.3
R11 minus.n12 minus.n7 161.3
R12 minus.n71 minus.n70 161.3
R13 minus.n69 minus.n36 161.3
R14 minus.n65 minus.n64 161.3
R15 minus.n63 minus.n38 161.3
R16 minus.n62 minus.n61 161.3
R17 minus.n60 minus.n39 161.3
R18 minus.n59 minus.n58 161.3
R19 minus.n54 minus.n41 161.3
R20 minus.n53 minus.n52 161.3
R21 minus.n51 minus.n42 161.3
R22 minus.n50 minus.n49 161.3
R23 minus.n48 minus.n43 161.3
R24 minus.n8 minus.t13 130.791
R25 minus.n44 minus.t22 130.791
R26 minus.n9 minus.t9 109.355
R27 minus.n10 minus.t8 109.355
R28 minus.n14 minus.t17 109.355
R29 minus.n16 minus.t19 109.355
R30 minus.n20 minus.t15 109.355
R31 minus.n21 minus.t11 109.355
R32 minus.n3 minus.t21 109.355
R33 minus.n27 minus.t18 109.355
R34 minus.n1 minus.t5 109.355
R35 minus.n32 minus.t12 109.355
R36 minus.n34 minus.t10 109.355
R37 minus.n45 minus.t1 109.355
R38 minus.n46 minus.t23 109.355
R39 minus.n50 minus.t2 109.355
R40 minus.n52 minus.t14 109.355
R41 minus.n56 minus.t3 109.355
R42 minus.n57 minus.t16 109.355
R43 minus.n39 minus.t4 109.355
R44 minus.n63 minus.t20 109.355
R45 minus.n37 minus.t7 109.355
R46 minus.n68 minus.t0 109.355
R47 minus.n70 minus.t6 109.355
R48 minus.n32 minus.n31 80.6037
R49 minus.n30 minus.n1 80.6037
R50 minus.n21 minus.n4 80.6037
R51 minus.n20 minus.n19 80.6037
R52 minus.n11 minus.n10 80.6037
R53 minus.n68 minus.n67 80.6037
R54 minus.n66 minus.n37 80.6037
R55 minus.n57 minus.n40 80.6037
R56 minus.n56 minus.n55 80.6037
R57 minus.n47 minus.n46 80.6037
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n20 minus.n5 41.6278
R69 minus.n22 minus.n21 41.6278
R70 minus.n56 minus.n41 41.6278
R71 minus.n58 minus.n57 41.6278
R72 minus.n33 minus.n32 38.7066
R73 minus.n69 minus.n68 38.7066
R74 minus.n72 minus.n35 35.546
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 drain_right.n13 drain_right.n11 101.769
R132 drain_right.n7 drain_right.n5 101.769
R133 drain_right.n2 drain_right.n0 101.769
R134 drain_right.n13 drain_right.n12 100.796
R135 drain_right.n15 drain_right.n14 100.796
R136 drain_right.n17 drain_right.n16 100.796
R137 drain_right.n19 drain_right.n18 100.796
R138 drain_right.n21 drain_right.n20 100.796
R139 drain_right.n7 drain_right.n6 100.796
R140 drain_right.n9 drain_right.n8 100.796
R141 drain_right.n4 drain_right.n3 100.796
R142 drain_right.n2 drain_right.n1 100.796
R143 drain_right drain_right.n10 28.4924
R144 drain_right.n5 drain_right.t17 9.9005
R145 drain_right.n5 drain_right.t5 9.9005
R146 drain_right.n6 drain_right.t2 9.9005
R147 drain_right.n6 drain_right.t16 9.9005
R148 drain_right.n8 drain_right.t4 9.9005
R149 drain_right.n8 drain_right.t3 9.9005
R150 drain_right.n3 drain_right.t11 9.9005
R151 drain_right.n3 drain_right.t21 9.9005
R152 drain_right.n1 drain_right.t1 9.9005
R153 drain_right.n1 drain_right.t10 9.9005
R154 drain_right.n0 drain_right.t12 9.9005
R155 drain_right.n0 drain_right.t7 9.9005
R156 drain_right.n11 drain_right.t22 9.9005
R157 drain_right.n11 drain_right.t8 9.9005
R158 drain_right.n12 drain_right.t15 9.9005
R159 drain_right.n12 drain_right.t6 9.9005
R160 drain_right.n14 drain_right.t23 9.9005
R161 drain_right.n14 drain_right.t0 9.9005
R162 drain_right.n16 drain_right.t13 9.9005
R163 drain_right.n16 drain_right.t19 9.9005
R164 drain_right.n18 drain_right.t14 9.9005
R165 drain_right.n18 drain_right.t9 9.9005
R166 drain_right.n20 drain_right.t20 9.9005
R167 drain_right.n20 drain_right.t18 9.9005
R168 drain_right drain_right.n21 6.62735
R169 drain_right.n9 drain_right.n7 0.974638
R170 drain_right.n4 drain_right.n2 0.974638
R171 drain_right.n21 drain_right.n19 0.974638
R172 drain_right.n19 drain_right.n17 0.974638
R173 drain_right.n17 drain_right.n15 0.974638
R174 drain_right.n15 drain_right.n13 0.974638
R175 drain_right.n10 drain_right.n9 0.432223
R176 drain_right.n10 drain_right.n4 0.432223
R177 source.n98 source.n96 289.615
R178 source.n80 source.n78 289.615
R179 source.n72 source.n70 289.615
R180 source.n54 source.n52 289.615
R181 source.n2 source.n0 289.615
R182 source.n20 source.n18 289.615
R183 source.n28 source.n26 289.615
R184 source.n46 source.n44 289.615
R185 source.n99 source.n98 185
R186 source.n81 source.n80 185
R187 source.n73 source.n72 185
R188 source.n55 source.n54 185
R189 source.n3 source.n2 185
R190 source.n21 source.n20 185
R191 source.n29 source.n28 185
R192 source.n47 source.n46 185
R193 source.t41 source.n97 167.117
R194 source.t25 source.n79 167.117
R195 source.t5 source.n71 167.117
R196 source.t3 source.n53 167.117
R197 source.t1 source.n1 167.117
R198 source.t8 source.n19 167.117
R199 source.t34 source.n27 167.117
R200 source.t37 source.n45 167.117
R201 source.n9 source.n8 84.1169
R202 source.n11 source.n10 84.1169
R203 source.n13 source.n12 84.1169
R204 source.n15 source.n14 84.1169
R205 source.n17 source.n16 84.1169
R206 source.n35 source.n34 84.1169
R207 source.n37 source.n36 84.1169
R208 source.n39 source.n38 84.1169
R209 source.n41 source.n40 84.1169
R210 source.n43 source.n42 84.1169
R211 source.n95 source.n94 84.1168
R212 source.n93 source.n92 84.1168
R213 source.n91 source.n90 84.1168
R214 source.n89 source.n88 84.1168
R215 source.n87 source.n86 84.1168
R216 source.n69 source.n68 84.1168
R217 source.n67 source.n66 84.1168
R218 source.n65 source.n64 84.1168
R219 source.n63 source.n62 84.1168
R220 source.n61 source.n60 84.1168
R221 source.n98 source.t41 52.3082
R222 source.n80 source.t25 52.3082
R223 source.n72 source.t5 52.3082
R224 source.n54 source.t3 52.3082
R225 source.n2 source.t1 52.3082
R226 source.n20 source.t8 52.3082
R227 source.n28 source.t34 52.3082
R228 source.n46 source.t37 52.3082
R229 source.n103 source.n102 31.4096
R230 source.n85 source.n84 31.4096
R231 source.n77 source.n76 31.4096
R232 source.n59 source.n58 31.4096
R233 source.n7 source.n6 31.4096
R234 source.n25 source.n24 31.4096
R235 source.n33 source.n32 31.4096
R236 source.n51 source.n50 31.4096
R237 source.n59 source.n51 14.6861
R238 source.n94 source.t40 9.9005
R239 source.n94 source.t47 9.9005
R240 source.n92 source.t43 9.9005
R241 source.n92 source.t27 9.9005
R242 source.n90 source.t44 9.9005
R243 source.n90 source.t31 9.9005
R244 source.n88 source.t45 9.9005
R245 source.n88 source.t33 9.9005
R246 source.n86 source.t46 9.9005
R247 source.n86 source.t24 9.9005
R248 source.n68 source.t11 9.9005
R249 source.n68 source.t10 9.9005
R250 source.n66 source.t22 9.9005
R251 source.n66 source.t4 9.9005
R252 source.n64 source.t17 9.9005
R253 source.n64 source.t13 9.9005
R254 source.n62 source.t7 9.9005
R255 source.n62 source.t6 9.9005
R256 source.n60 source.t2 9.9005
R257 source.n60 source.t16 9.9005
R258 source.n8 source.t14 9.9005
R259 source.n8 source.t23 9.9005
R260 source.n10 source.t19 9.9005
R261 source.n10 source.t18 9.9005
R262 source.n12 source.t21 9.9005
R263 source.n12 source.t20 9.9005
R264 source.n14 source.t0 9.9005
R265 source.n14 source.t9 9.9005
R266 source.n16 source.t12 9.9005
R267 source.n16 source.t15 9.9005
R268 source.n34 source.t39 9.9005
R269 source.n34 source.t38 9.9005
R270 source.n36 source.t28 9.9005
R271 source.n36 source.t30 9.9005
R272 source.n38 source.t36 9.9005
R273 source.n38 source.t32 9.9005
R274 source.n40 source.t29 9.9005
R275 source.n40 source.t26 9.9005
R276 source.n42 source.t35 9.9005
R277 source.n42 source.t42 9.9005
R278 source.n99 source.n97 9.71174
R279 source.n81 source.n79 9.71174
R280 source.n73 source.n71 9.71174
R281 source.n55 source.n53 9.71174
R282 source.n3 source.n1 9.71174
R283 source.n21 source.n19 9.71174
R284 source.n29 source.n27 9.71174
R285 source.n47 source.n45 9.71174
R286 source.n102 source.n101 9.45567
R287 source.n84 source.n83 9.45567
R288 source.n76 source.n75 9.45567
R289 source.n58 source.n57 9.45567
R290 source.n6 source.n5 9.45567
R291 source.n24 source.n23 9.45567
R292 source.n32 source.n31 9.45567
R293 source.n50 source.n49 9.45567
R294 source.n101 source.n100 9.3005
R295 source.n83 source.n82 9.3005
R296 source.n75 source.n74 9.3005
R297 source.n57 source.n56 9.3005
R298 source.n5 source.n4 9.3005
R299 source.n23 source.n22 9.3005
R300 source.n31 source.n30 9.3005
R301 source.n49 source.n48 9.3005
R302 source.n104 source.n7 8.93611
R303 source.n102 source.n96 8.14595
R304 source.n84 source.n78 8.14595
R305 source.n76 source.n70 8.14595
R306 source.n58 source.n52 8.14595
R307 source.n6 source.n0 8.14595
R308 source.n24 source.n18 8.14595
R309 source.n32 source.n26 8.14595
R310 source.n50 source.n44 8.14595
R311 source.n100 source.n99 7.3702
R312 source.n82 source.n81 7.3702
R313 source.n74 source.n73 7.3702
R314 source.n56 source.n55 7.3702
R315 source.n4 source.n3 7.3702
R316 source.n22 source.n21 7.3702
R317 source.n30 source.n29 7.3702
R318 source.n48 source.n47 7.3702
R319 source.n100 source.n96 5.81868
R320 source.n82 source.n78 5.81868
R321 source.n74 source.n70 5.81868
R322 source.n56 source.n52 5.81868
R323 source.n4 source.n0 5.81868
R324 source.n22 source.n18 5.81868
R325 source.n30 source.n26 5.81868
R326 source.n48 source.n44 5.81868
R327 source.n104 source.n103 5.7505
R328 source.n101 source.n97 3.44771
R329 source.n83 source.n79 3.44771
R330 source.n75 source.n71 3.44771
R331 source.n57 source.n53 3.44771
R332 source.n5 source.n1 3.44771
R333 source.n23 source.n19 3.44771
R334 source.n31 source.n27 3.44771
R335 source.n49 source.n45 3.44771
R336 source.n51 source.n43 0.974638
R337 source.n43 source.n41 0.974638
R338 source.n41 source.n39 0.974638
R339 source.n39 source.n37 0.974638
R340 source.n37 source.n35 0.974638
R341 source.n35 source.n33 0.974638
R342 source.n25 source.n17 0.974638
R343 source.n17 source.n15 0.974638
R344 source.n15 source.n13 0.974638
R345 source.n13 source.n11 0.974638
R346 source.n11 source.n9 0.974638
R347 source.n9 source.n7 0.974638
R348 source.n61 source.n59 0.974638
R349 source.n63 source.n61 0.974638
R350 source.n65 source.n63 0.974638
R351 source.n67 source.n65 0.974638
R352 source.n69 source.n67 0.974638
R353 source.n77 source.n69 0.974638
R354 source.n87 source.n85 0.974638
R355 source.n89 source.n87 0.974638
R356 source.n91 source.n89 0.974638
R357 source.n93 source.n91 0.974638
R358 source.n95 source.n93 0.974638
R359 source.n103 source.n95 0.974638
R360 source.n33 source.n25 0.470328
R361 source.n85 source.n77 0.470328
R362 source source.n104 0.188
R363 plus.n14 plus.n13 161.3
R364 plus.n15 plus.n8 161.3
R365 plus.n17 plus.n16 161.3
R366 plus.n18 plus.n7 161.3
R367 plus.n19 plus.n6 161.3
R368 plus.n24 plus.n23 161.3
R369 plus.n25 plus.n4 161.3
R370 plus.n27 plus.n26 161.3
R371 plus.n28 plus.n3 161.3
R372 plus.n30 plus.n29 161.3
R373 plus.n33 plus.n0 161.3
R374 plus.n35 plus.n34 161.3
R375 plus.n50 plus.n49 161.3
R376 plus.n51 plus.n44 161.3
R377 plus.n53 plus.n52 161.3
R378 plus.n54 plus.n43 161.3
R379 plus.n55 plus.n42 161.3
R380 plus.n60 plus.n59 161.3
R381 plus.n61 plus.n40 161.3
R382 plus.n63 plus.n62 161.3
R383 plus.n64 plus.n39 161.3
R384 plus.n66 plus.n65 161.3
R385 plus.n69 plus.n36 161.3
R386 plus.n71 plus.n70 161.3
R387 plus.n10 plus.t22 130.791
R388 plus.n46 plus.t21 130.791
R389 plus.n34 plus.t5 109.355
R390 plus.n32 plus.t7 109.355
R391 plus.n31 plus.t8 109.355
R392 plus.n3 plus.t9 109.355
R393 plus.n25 plus.t11 109.355
R394 plus.n5 plus.t14 109.355
R395 plus.n20 plus.t15 109.355
R396 plus.n18 plus.t19 109.355
R397 plus.n8 plus.t16 109.355
R398 plus.n12 plus.t17 109.355
R399 plus.n11 plus.t20 109.355
R400 plus.n70 plus.t1 109.355
R401 plus.n68 plus.t18 109.355
R402 plus.n67 plus.t6 109.355
R403 plus.n39 plus.t13 109.355
R404 plus.n61 plus.t0 109.355
R405 plus.n41 plus.t12 109.355
R406 plus.n56 plus.t4 109.355
R407 plus.n54 plus.t10 109.355
R408 plus.n44 plus.t3 109.355
R409 plus.n48 plus.t23 109.355
R410 plus.n47 plus.t2 109.355
R411 plus.n12 plus.n9 80.6037
R412 plus.n21 plus.n20 80.6037
R413 plus.n22 plus.n5 80.6037
R414 plus.n31 plus.n2 80.6037
R415 plus.n32 plus.n1 80.6037
R416 plus.n48 plus.n45 80.6037
R417 plus.n57 plus.n56 80.6037
R418 plus.n58 plus.n41 80.6037
R419 plus.n67 plus.n38 80.6037
R420 plus.n68 plus.n37 80.6037
R421 plus.n32 plus.n31 48.2005
R422 plus.n20 plus.n5 48.2005
R423 plus.n12 plus.n11 48.2005
R424 plus.n68 plus.n67 48.2005
R425 plus.n56 plus.n41 48.2005
R426 plus.n48 plus.n47 48.2005
R427 plus.n31 plus.n30 44.549
R428 plus.n13 plus.n12 44.549
R429 plus.n67 plus.n66 44.549
R430 plus.n49 plus.n48 44.549
R431 plus.n24 plus.n5 41.6278
R432 plus.n20 plus.n19 41.6278
R433 plus.n60 plus.n41 41.6278
R434 plus.n56 plus.n55 41.6278
R435 plus.n33 plus.n32 38.7066
R436 plus.n69 plus.n68 38.7066
R437 plus plus.n71 33.2149
R438 plus.n10 plus.n9 31.6825
R439 plus.n46 plus.n45 31.6825
R440 plus.n26 plus.n3 25.5611
R441 plus.n17 plus.n8 25.5611
R442 plus.n62 plus.n39 25.5611
R443 plus.n53 plus.n44 25.5611
R444 plus.n26 plus.n25 22.6399
R445 plus.n18 plus.n17 22.6399
R446 plus.n62 plus.n61 22.6399
R447 plus.n54 plus.n53 22.6399
R448 plus.n11 plus.n10 17.2341
R449 plus.n47 plus.n46 17.2341
R450 plus.n34 plus.n33 9.49444
R451 plus.n70 plus.n69 9.49444
R452 plus plus.n35 8.51565
R453 plus.n25 plus.n24 6.57323
R454 plus.n19 plus.n18 6.57323
R455 plus.n61 plus.n60 6.57323
R456 plus.n55 plus.n54 6.57323
R457 plus.n30 plus.n3 3.65202
R458 plus.n13 plus.n8 3.65202
R459 plus.n66 plus.n39 3.65202
R460 plus.n49 plus.n44 3.65202
R461 plus.n22 plus.n21 0.380177
R462 plus.n2 plus.n1 0.380177
R463 plus.n38 plus.n37 0.380177
R464 plus.n58 plus.n57 0.380177
R465 plus.n14 plus.n9 0.285035
R466 plus.n21 plus.n6 0.285035
R467 plus.n23 plus.n22 0.285035
R468 plus.n29 plus.n2 0.285035
R469 plus.n1 plus.n0 0.285035
R470 plus.n37 plus.n36 0.285035
R471 plus.n65 plus.n38 0.285035
R472 plus.n59 plus.n58 0.285035
R473 plus.n57 plus.n42 0.285035
R474 plus.n50 plus.n45 0.285035
R475 plus.n15 plus.n14 0.189894
R476 plus.n16 plus.n15 0.189894
R477 plus.n16 plus.n7 0.189894
R478 plus.n7 plus.n6 0.189894
R479 plus.n23 plus.n4 0.189894
R480 plus.n27 plus.n4 0.189894
R481 plus.n28 plus.n27 0.189894
R482 plus.n29 plus.n28 0.189894
R483 plus.n35 plus.n0 0.189894
R484 plus.n71 plus.n36 0.189894
R485 plus.n65 plus.n64 0.189894
R486 plus.n64 plus.n63 0.189894
R487 plus.n63 plus.n40 0.189894
R488 plus.n59 plus.n40 0.189894
R489 plus.n43 plus.n42 0.189894
R490 plus.n52 plus.n43 0.189894
R491 plus.n52 plus.n51 0.189894
R492 plus.n51 plus.n50 0.189894
R493 drain_left.n13 drain_left.n11 101.769
R494 drain_left.n7 drain_left.n5 101.769
R495 drain_left.n2 drain_left.n0 101.769
R496 drain_left.n21 drain_left.n20 100.796
R497 drain_left.n19 drain_left.n18 100.796
R498 drain_left.n17 drain_left.n16 100.796
R499 drain_left.n15 drain_left.n14 100.796
R500 drain_left.n13 drain_left.n12 100.796
R501 drain_left.n7 drain_left.n6 100.796
R502 drain_left.n9 drain_left.n8 100.796
R503 drain_left.n4 drain_left.n3 100.796
R504 drain_left.n2 drain_left.n1 100.796
R505 drain_left drain_left.n10 29.0456
R506 drain_left.n5 drain_left.t21 9.9005
R507 drain_left.n5 drain_left.t2 9.9005
R508 drain_left.n6 drain_left.t20 9.9005
R509 drain_left.n6 drain_left.t0 9.9005
R510 drain_left.n8 drain_left.t19 9.9005
R511 drain_left.n8 drain_left.t13 9.9005
R512 drain_left.n3 drain_left.t23 9.9005
R513 drain_left.n3 drain_left.t11 9.9005
R514 drain_left.n1 drain_left.t17 9.9005
R515 drain_left.n1 drain_left.t10 9.9005
R516 drain_left.n0 drain_left.t22 9.9005
R517 drain_left.n0 drain_left.t5 9.9005
R518 drain_left.n20 drain_left.t16 9.9005
R519 drain_left.n20 drain_left.t18 9.9005
R520 drain_left.n18 drain_left.t14 9.9005
R521 drain_left.n18 drain_left.t15 9.9005
R522 drain_left.n16 drain_left.t9 9.9005
R523 drain_left.n16 drain_left.t12 9.9005
R524 drain_left.n14 drain_left.t4 9.9005
R525 drain_left.n14 drain_left.t8 9.9005
R526 drain_left.n12 drain_left.t6 9.9005
R527 drain_left.n12 drain_left.t7 9.9005
R528 drain_left.n11 drain_left.t1 9.9005
R529 drain_left.n11 drain_left.t3 9.9005
R530 drain_left drain_left.n21 6.62735
R531 drain_left.n9 drain_left.n7 0.974638
R532 drain_left.n4 drain_left.n2 0.974638
R533 drain_left.n15 drain_left.n13 0.974638
R534 drain_left.n17 drain_left.n15 0.974638
R535 drain_left.n19 drain_left.n17 0.974638
R536 drain_left.n21 drain_left.n19 0.974638
R537 drain_left.n10 drain_left.n9 0.432223
R538 drain_left.n10 drain_left.n4 0.432223
C0 drain_left minus 0.181449f
C1 drain_right minus 3.34573f
C2 source minus 4.36704f
C3 plus minus 5.86513f
C4 drain_left drain_right 2.02887f
C5 drain_left source 8.592389f
C6 source drain_right 8.59548f
C7 plus drain_left 3.71298f
C8 plus drain_right 0.533985f
C9 plus source 4.381f
C10 drain_right a_n3654_n1288# 6.56749f
C11 drain_left a_n3654_n1288# 7.10875f
C12 source a_n3654_n1288# 3.750305f
C13 minus a_n3654_n1288# 14.011654f
C14 plus a_n3654_n1288# 15.472549f
C15 drain_left.t22 a_n3654_n1288# 0.049716f
C16 drain_left.t5 a_n3654_n1288# 0.049716f
C17 drain_left.n0 a_n3654_n1288# 0.316645f
C18 drain_left.t17 a_n3654_n1288# 0.049716f
C19 drain_left.t10 a_n3654_n1288# 0.049716f
C20 drain_left.n1 a_n3654_n1288# 0.312329f
C21 drain_left.n2 a_n3654_n1288# 0.884835f
C22 drain_left.t23 a_n3654_n1288# 0.049716f
C23 drain_left.t11 a_n3654_n1288# 0.049716f
C24 drain_left.n3 a_n3654_n1288# 0.312329f
C25 drain_left.n4 a_n3654_n1288# 0.384951f
C26 drain_left.t21 a_n3654_n1288# 0.049716f
C27 drain_left.t2 a_n3654_n1288# 0.049716f
C28 drain_left.n5 a_n3654_n1288# 0.316645f
C29 drain_left.t20 a_n3654_n1288# 0.049716f
C30 drain_left.t0 a_n3654_n1288# 0.049716f
C31 drain_left.n6 a_n3654_n1288# 0.312329f
C32 drain_left.n7 a_n3654_n1288# 0.884835f
C33 drain_left.t19 a_n3654_n1288# 0.049716f
C34 drain_left.t13 a_n3654_n1288# 0.049716f
C35 drain_left.n8 a_n3654_n1288# 0.312329f
C36 drain_left.n9 a_n3654_n1288# 0.384951f
C37 drain_left.n10 a_n3654_n1288# 1.49978f
C38 drain_left.t1 a_n3654_n1288# 0.049716f
C39 drain_left.t3 a_n3654_n1288# 0.049716f
C40 drain_left.n11 a_n3654_n1288# 0.316646f
C41 drain_left.t6 a_n3654_n1288# 0.049716f
C42 drain_left.t7 a_n3654_n1288# 0.049716f
C43 drain_left.n12 a_n3654_n1288# 0.31233f
C44 drain_left.n13 a_n3654_n1288# 0.884833f
C45 drain_left.t4 a_n3654_n1288# 0.049716f
C46 drain_left.t8 a_n3654_n1288# 0.049716f
C47 drain_left.n14 a_n3654_n1288# 0.31233f
C48 drain_left.n15 a_n3654_n1288# 0.438239f
C49 drain_left.t9 a_n3654_n1288# 0.049716f
C50 drain_left.t12 a_n3654_n1288# 0.049716f
C51 drain_left.n16 a_n3654_n1288# 0.31233f
C52 drain_left.n17 a_n3654_n1288# 0.438239f
C53 drain_left.t14 a_n3654_n1288# 0.049716f
C54 drain_left.t15 a_n3654_n1288# 0.049716f
C55 drain_left.n18 a_n3654_n1288# 0.31233f
C56 drain_left.n19 a_n3654_n1288# 0.438239f
C57 drain_left.t16 a_n3654_n1288# 0.049716f
C58 drain_left.t18 a_n3654_n1288# 0.049716f
C59 drain_left.n20 a_n3654_n1288# 0.31233f
C60 drain_left.n21 a_n3654_n1288# 0.720307f
C61 plus.n0 a_n3654_n1288# 0.055243f
C62 plus.t5 a_n3654_n1288# 0.205125f
C63 plus.t7 a_n3654_n1288# 0.205125f
C64 plus.n1 a_n3654_n1288# 0.068956f
C65 plus.t8 a_n3654_n1288# 0.205125f
C66 plus.n2 a_n3654_n1288# 0.068956f
C67 plus.t9 a_n3654_n1288# 0.205125f
C68 plus.n3 a_n3654_n1288# 0.138804f
C69 plus.n4 a_n3654_n1288# 0.0414f
C70 plus.t11 a_n3654_n1288# 0.205125f
C71 plus.t14 a_n3654_n1288# 0.205125f
C72 plus.n5 a_n3654_n1288# 0.150368f
C73 plus.n6 a_n3654_n1288# 0.055243f
C74 plus.t15 a_n3654_n1288# 0.205125f
C75 plus.t19 a_n3654_n1288# 0.205125f
C76 plus.n7 a_n3654_n1288# 0.0414f
C77 plus.t16 a_n3654_n1288# 0.205125f
C78 plus.n8 a_n3654_n1288# 0.138804f
C79 plus.n9 a_n3654_n1288# 0.237949f
C80 plus.t17 a_n3654_n1288# 0.205125f
C81 plus.t20 a_n3654_n1288# 0.205125f
C82 plus.t22 a_n3654_n1288# 0.228446f
C83 plus.n10 a_n3654_n1288# 0.122907f
C84 plus.n11 a_n3654_n1288# 0.150857f
C85 plus.n12 a_n3654_n1288# 0.150879f
C86 plus.n13 a_n3654_n1288# 0.009394f
C87 plus.n14 a_n3654_n1288# 0.055243f
C88 plus.n15 a_n3654_n1288# 0.0414f
C89 plus.n16 a_n3654_n1288# 0.0414f
C90 plus.n17 a_n3654_n1288# 0.009394f
C91 plus.n18 a_n3654_n1288# 0.138804f
C92 plus.n19 a_n3654_n1288# 0.009394f
C93 plus.n20 a_n3654_n1288# 0.150368f
C94 plus.n21 a_n3654_n1288# 0.068956f
C95 plus.n22 a_n3654_n1288# 0.068956f
C96 plus.n23 a_n3654_n1288# 0.055243f
C97 plus.n24 a_n3654_n1288# 0.009394f
C98 plus.n25 a_n3654_n1288# 0.138804f
C99 plus.n26 a_n3654_n1288# 0.009394f
C100 plus.n27 a_n3654_n1288# 0.0414f
C101 plus.n28 a_n3654_n1288# 0.0414f
C102 plus.n29 a_n3654_n1288# 0.055243f
C103 plus.n30 a_n3654_n1288# 0.009394f
C104 plus.n31 a_n3654_n1288# 0.150879f
C105 plus.n32 a_n3654_n1288# 0.149858f
C106 plus.n33 a_n3654_n1288# 0.009394f
C107 plus.n34 a_n3654_n1288# 0.135358f
C108 plus.n35 a_n3654_n1288# 0.312258f
C109 plus.n36 a_n3654_n1288# 0.055243f
C110 plus.t1 a_n3654_n1288# 0.205125f
C111 plus.n37 a_n3654_n1288# 0.068956f
C112 plus.t18 a_n3654_n1288# 0.205125f
C113 plus.n38 a_n3654_n1288# 0.068956f
C114 plus.t6 a_n3654_n1288# 0.205125f
C115 plus.t13 a_n3654_n1288# 0.205125f
C116 plus.n39 a_n3654_n1288# 0.138804f
C117 plus.n40 a_n3654_n1288# 0.0414f
C118 plus.t0 a_n3654_n1288# 0.205125f
C119 plus.t12 a_n3654_n1288# 0.205125f
C120 plus.n41 a_n3654_n1288# 0.150368f
C121 plus.n42 a_n3654_n1288# 0.055243f
C122 plus.t4 a_n3654_n1288# 0.205125f
C123 plus.n43 a_n3654_n1288# 0.0414f
C124 plus.t10 a_n3654_n1288# 0.205125f
C125 plus.t3 a_n3654_n1288# 0.205125f
C126 plus.n44 a_n3654_n1288# 0.138804f
C127 plus.n45 a_n3654_n1288# 0.237949f
C128 plus.t23 a_n3654_n1288# 0.205125f
C129 plus.t21 a_n3654_n1288# 0.228446f
C130 plus.n46 a_n3654_n1288# 0.122907f
C131 plus.t2 a_n3654_n1288# 0.205125f
C132 plus.n47 a_n3654_n1288# 0.150857f
C133 plus.n48 a_n3654_n1288# 0.150879f
C134 plus.n49 a_n3654_n1288# 0.009394f
C135 plus.n50 a_n3654_n1288# 0.055243f
C136 plus.n51 a_n3654_n1288# 0.0414f
C137 plus.n52 a_n3654_n1288# 0.0414f
C138 plus.n53 a_n3654_n1288# 0.009394f
C139 plus.n54 a_n3654_n1288# 0.138804f
C140 plus.n55 a_n3654_n1288# 0.009394f
C141 plus.n56 a_n3654_n1288# 0.150368f
C142 plus.n57 a_n3654_n1288# 0.068956f
C143 plus.n58 a_n3654_n1288# 0.068956f
C144 plus.n59 a_n3654_n1288# 0.055243f
C145 plus.n60 a_n3654_n1288# 0.009394f
C146 plus.n61 a_n3654_n1288# 0.138804f
C147 plus.n62 a_n3654_n1288# 0.009394f
C148 plus.n63 a_n3654_n1288# 0.0414f
C149 plus.n64 a_n3654_n1288# 0.0414f
C150 plus.n65 a_n3654_n1288# 0.055243f
C151 plus.n66 a_n3654_n1288# 0.009394f
C152 plus.n67 a_n3654_n1288# 0.150879f
C153 plus.n68 a_n3654_n1288# 0.149858f
C154 plus.n69 a_n3654_n1288# 0.009394f
C155 plus.n70 a_n3654_n1288# 0.135358f
C156 plus.n71 a_n3654_n1288# 1.35668f
C157 source.n0 a_n3654_n1288# 0.047198f
C158 source.n1 a_n3654_n1288# 0.104432f
C159 source.t1 a_n3654_n1288# 0.078371f
C160 source.n2 a_n3654_n1288# 0.081732f
C161 source.n3 a_n3654_n1288# 0.026347f
C162 source.n4 a_n3654_n1288# 0.017377f
C163 source.n5 a_n3654_n1288# 0.230193f
C164 source.n6 a_n3654_n1288# 0.05174f
C165 source.n7 a_n3654_n1288# 0.567754f
C166 source.t14 a_n3654_n1288# 0.051108f
C167 source.t23 a_n3654_n1288# 0.051108f
C168 source.n8 a_n3654_n1288# 0.27322f
C169 source.n9 a_n3654_n1288# 0.454412f
C170 source.t19 a_n3654_n1288# 0.051108f
C171 source.t18 a_n3654_n1288# 0.051108f
C172 source.n10 a_n3654_n1288# 0.27322f
C173 source.n11 a_n3654_n1288# 0.454412f
C174 source.t21 a_n3654_n1288# 0.051108f
C175 source.t20 a_n3654_n1288# 0.051108f
C176 source.n12 a_n3654_n1288# 0.27322f
C177 source.n13 a_n3654_n1288# 0.454412f
C178 source.t0 a_n3654_n1288# 0.051108f
C179 source.t9 a_n3654_n1288# 0.051108f
C180 source.n14 a_n3654_n1288# 0.27322f
C181 source.n15 a_n3654_n1288# 0.454412f
C182 source.t12 a_n3654_n1288# 0.051108f
C183 source.t15 a_n3654_n1288# 0.051108f
C184 source.n16 a_n3654_n1288# 0.27322f
C185 source.n17 a_n3654_n1288# 0.454412f
C186 source.n18 a_n3654_n1288# 0.047198f
C187 source.n19 a_n3654_n1288# 0.104432f
C188 source.t8 a_n3654_n1288# 0.078371f
C189 source.n20 a_n3654_n1288# 0.081732f
C190 source.n21 a_n3654_n1288# 0.026347f
C191 source.n22 a_n3654_n1288# 0.017377f
C192 source.n23 a_n3654_n1288# 0.230193f
C193 source.n24 a_n3654_n1288# 0.05174f
C194 source.n25 a_n3654_n1288# 0.177079f
C195 source.n26 a_n3654_n1288# 0.047198f
C196 source.n27 a_n3654_n1288# 0.104432f
C197 source.t34 a_n3654_n1288# 0.078371f
C198 source.n28 a_n3654_n1288# 0.081732f
C199 source.n29 a_n3654_n1288# 0.026347f
C200 source.n30 a_n3654_n1288# 0.017377f
C201 source.n31 a_n3654_n1288# 0.230193f
C202 source.n32 a_n3654_n1288# 0.05174f
C203 source.n33 a_n3654_n1288# 0.177079f
C204 source.t39 a_n3654_n1288# 0.051108f
C205 source.t38 a_n3654_n1288# 0.051108f
C206 source.n34 a_n3654_n1288# 0.27322f
C207 source.n35 a_n3654_n1288# 0.454412f
C208 source.t28 a_n3654_n1288# 0.051108f
C209 source.t30 a_n3654_n1288# 0.051108f
C210 source.n36 a_n3654_n1288# 0.27322f
C211 source.n37 a_n3654_n1288# 0.454412f
C212 source.t36 a_n3654_n1288# 0.051108f
C213 source.t32 a_n3654_n1288# 0.051108f
C214 source.n38 a_n3654_n1288# 0.27322f
C215 source.n39 a_n3654_n1288# 0.454412f
C216 source.t29 a_n3654_n1288# 0.051108f
C217 source.t26 a_n3654_n1288# 0.051108f
C218 source.n40 a_n3654_n1288# 0.27322f
C219 source.n41 a_n3654_n1288# 0.454412f
C220 source.t35 a_n3654_n1288# 0.051108f
C221 source.t42 a_n3654_n1288# 0.051108f
C222 source.n42 a_n3654_n1288# 0.27322f
C223 source.n43 a_n3654_n1288# 0.454412f
C224 source.n44 a_n3654_n1288# 0.047198f
C225 source.n45 a_n3654_n1288# 0.104432f
C226 source.t37 a_n3654_n1288# 0.078371f
C227 source.n46 a_n3654_n1288# 0.081732f
C228 source.n47 a_n3654_n1288# 0.026347f
C229 source.n48 a_n3654_n1288# 0.017377f
C230 source.n49 a_n3654_n1288# 0.230193f
C231 source.n50 a_n3654_n1288# 0.05174f
C232 source.n51 a_n3654_n1288# 0.879545f
C233 source.n52 a_n3654_n1288# 0.047198f
C234 source.n53 a_n3654_n1288# 0.104432f
C235 source.t3 a_n3654_n1288# 0.078371f
C236 source.n54 a_n3654_n1288# 0.081732f
C237 source.n55 a_n3654_n1288# 0.026347f
C238 source.n56 a_n3654_n1288# 0.017377f
C239 source.n57 a_n3654_n1288# 0.230193f
C240 source.n58 a_n3654_n1288# 0.05174f
C241 source.n59 a_n3654_n1288# 0.879545f
C242 source.t2 a_n3654_n1288# 0.051108f
C243 source.t16 a_n3654_n1288# 0.051108f
C244 source.n60 a_n3654_n1288# 0.273218f
C245 source.n61 a_n3654_n1288# 0.454414f
C246 source.t7 a_n3654_n1288# 0.051108f
C247 source.t6 a_n3654_n1288# 0.051108f
C248 source.n62 a_n3654_n1288# 0.273218f
C249 source.n63 a_n3654_n1288# 0.454414f
C250 source.t17 a_n3654_n1288# 0.051108f
C251 source.t13 a_n3654_n1288# 0.051108f
C252 source.n64 a_n3654_n1288# 0.273218f
C253 source.n65 a_n3654_n1288# 0.454414f
C254 source.t22 a_n3654_n1288# 0.051108f
C255 source.t4 a_n3654_n1288# 0.051108f
C256 source.n66 a_n3654_n1288# 0.273218f
C257 source.n67 a_n3654_n1288# 0.454414f
C258 source.t11 a_n3654_n1288# 0.051108f
C259 source.t10 a_n3654_n1288# 0.051108f
C260 source.n68 a_n3654_n1288# 0.273218f
C261 source.n69 a_n3654_n1288# 0.454414f
C262 source.n70 a_n3654_n1288# 0.047198f
C263 source.n71 a_n3654_n1288# 0.104432f
C264 source.t5 a_n3654_n1288# 0.078371f
C265 source.n72 a_n3654_n1288# 0.081732f
C266 source.n73 a_n3654_n1288# 0.026347f
C267 source.n74 a_n3654_n1288# 0.017377f
C268 source.n75 a_n3654_n1288# 0.230193f
C269 source.n76 a_n3654_n1288# 0.05174f
C270 source.n77 a_n3654_n1288# 0.177079f
C271 source.n78 a_n3654_n1288# 0.047198f
C272 source.n79 a_n3654_n1288# 0.104432f
C273 source.t25 a_n3654_n1288# 0.078371f
C274 source.n80 a_n3654_n1288# 0.081732f
C275 source.n81 a_n3654_n1288# 0.026347f
C276 source.n82 a_n3654_n1288# 0.017377f
C277 source.n83 a_n3654_n1288# 0.230193f
C278 source.n84 a_n3654_n1288# 0.05174f
C279 source.n85 a_n3654_n1288# 0.177079f
C280 source.t46 a_n3654_n1288# 0.051108f
C281 source.t24 a_n3654_n1288# 0.051108f
C282 source.n86 a_n3654_n1288# 0.273218f
C283 source.n87 a_n3654_n1288# 0.454414f
C284 source.t45 a_n3654_n1288# 0.051108f
C285 source.t33 a_n3654_n1288# 0.051108f
C286 source.n88 a_n3654_n1288# 0.273218f
C287 source.n89 a_n3654_n1288# 0.454414f
C288 source.t44 a_n3654_n1288# 0.051108f
C289 source.t31 a_n3654_n1288# 0.051108f
C290 source.n90 a_n3654_n1288# 0.273218f
C291 source.n91 a_n3654_n1288# 0.454414f
C292 source.t43 a_n3654_n1288# 0.051108f
C293 source.t27 a_n3654_n1288# 0.051108f
C294 source.n92 a_n3654_n1288# 0.273218f
C295 source.n93 a_n3654_n1288# 0.454414f
C296 source.t40 a_n3654_n1288# 0.051108f
C297 source.t47 a_n3654_n1288# 0.051108f
C298 source.n94 a_n3654_n1288# 0.273218f
C299 source.n95 a_n3654_n1288# 0.454414f
C300 source.n96 a_n3654_n1288# 0.047198f
C301 source.n97 a_n3654_n1288# 0.104432f
C302 source.t41 a_n3654_n1288# 0.078371f
C303 source.n98 a_n3654_n1288# 0.081732f
C304 source.n99 a_n3654_n1288# 0.026347f
C305 source.n100 a_n3654_n1288# 0.017377f
C306 source.n101 a_n3654_n1288# 0.230193f
C307 source.n102 a_n3654_n1288# 0.05174f
C308 source.n103 a_n3654_n1288# 0.395016f
C309 source.n104 a_n3654_n1288# 0.81932f
C310 drain_right.t12 a_n3654_n1288# 0.048744f
C311 drain_right.t7 a_n3654_n1288# 0.048744f
C312 drain_right.n0 a_n3654_n1288# 0.310459f
C313 drain_right.t1 a_n3654_n1288# 0.048744f
C314 drain_right.t10 a_n3654_n1288# 0.048744f
C315 drain_right.n1 a_n3654_n1288# 0.306227f
C316 drain_right.n2 a_n3654_n1288# 0.86755f
C317 drain_right.t11 a_n3654_n1288# 0.048744f
C318 drain_right.t21 a_n3654_n1288# 0.048744f
C319 drain_right.n3 a_n3654_n1288# 0.306227f
C320 drain_right.n4 a_n3654_n1288# 0.377431f
C321 drain_right.t17 a_n3654_n1288# 0.048744f
C322 drain_right.t5 a_n3654_n1288# 0.048744f
C323 drain_right.n5 a_n3654_n1288# 0.310459f
C324 drain_right.t2 a_n3654_n1288# 0.048744f
C325 drain_right.t16 a_n3654_n1288# 0.048744f
C326 drain_right.n6 a_n3654_n1288# 0.306227f
C327 drain_right.n7 a_n3654_n1288# 0.86755f
C328 drain_right.t4 a_n3654_n1288# 0.048744f
C329 drain_right.t3 a_n3654_n1288# 0.048744f
C330 drain_right.n8 a_n3654_n1288# 0.306227f
C331 drain_right.n9 a_n3654_n1288# 0.377431f
C332 drain_right.n10 a_n3654_n1288# 1.41106f
C333 drain_right.t22 a_n3654_n1288# 0.048744f
C334 drain_right.t8 a_n3654_n1288# 0.048744f
C335 drain_right.n11 a_n3654_n1288# 0.31046f
C336 drain_right.t15 a_n3654_n1288# 0.048744f
C337 drain_right.t6 a_n3654_n1288# 0.048744f
C338 drain_right.n12 a_n3654_n1288# 0.306229f
C339 drain_right.n13 a_n3654_n1288# 0.867547f
C340 drain_right.t23 a_n3654_n1288# 0.048744f
C341 drain_right.t0 a_n3654_n1288# 0.048744f
C342 drain_right.n14 a_n3654_n1288# 0.306229f
C343 drain_right.n15 a_n3654_n1288# 0.429678f
C344 drain_right.t13 a_n3654_n1288# 0.048744f
C345 drain_right.t19 a_n3654_n1288# 0.048744f
C346 drain_right.n16 a_n3654_n1288# 0.306229f
C347 drain_right.n17 a_n3654_n1288# 0.429678f
C348 drain_right.t14 a_n3654_n1288# 0.048744f
C349 drain_right.t9 a_n3654_n1288# 0.048744f
C350 drain_right.n18 a_n3654_n1288# 0.306229f
C351 drain_right.n19 a_n3654_n1288# 0.429678f
C352 drain_right.t20 a_n3654_n1288# 0.048744f
C353 drain_right.t18 a_n3654_n1288# 0.048744f
C354 drain_right.n20 a_n3654_n1288# 0.306229f
C355 drain_right.n21 a_n3654_n1288# 0.706236f
C356 minus.n0 a_n3654_n1288# 0.053345f
C357 minus.t5 a_n3654_n1288# 0.19808f
C358 minus.n1 a_n3654_n1288# 0.145697f
C359 minus.t12 a_n3654_n1288# 0.19808f
C360 minus.n2 a_n3654_n1288# 0.039978f
C361 minus.t21 a_n3654_n1288# 0.19808f
C362 minus.n3 a_n3654_n1288# 0.134037f
C363 minus.n4 a_n3654_n1288# 0.066588f
C364 minus.n5 a_n3654_n1288# 0.009072f
C365 minus.t15 a_n3654_n1288# 0.19808f
C366 minus.n6 a_n3654_n1288# 0.039978f
C367 minus.n7 a_n3654_n1288# 0.009072f
C368 minus.t17 a_n3654_n1288# 0.19808f
C369 minus.t13 a_n3654_n1288# 0.2206f
C370 minus.n8 a_n3654_n1288# 0.118686f
C371 minus.t9 a_n3654_n1288# 0.19808f
C372 minus.n9 a_n3654_n1288# 0.145676f
C373 minus.t8 a_n3654_n1288# 0.19808f
C374 minus.n10 a_n3654_n1288# 0.145697f
C375 minus.n11 a_n3654_n1288# 0.229777f
C376 minus.n12 a_n3654_n1288# 0.053345f
C377 minus.n13 a_n3654_n1288# 0.039978f
C378 minus.n14 a_n3654_n1288# 0.134037f
C379 minus.n15 a_n3654_n1288# 0.009072f
C380 minus.t19 a_n3654_n1288# 0.19808f
C381 minus.n16 a_n3654_n1288# 0.134037f
C382 minus.n17 a_n3654_n1288# 0.039978f
C383 minus.n18 a_n3654_n1288# 0.053345f
C384 minus.n19 a_n3654_n1288# 0.066588f
C385 minus.n20 a_n3654_n1288# 0.145204f
C386 minus.t11 a_n3654_n1288# 0.19808f
C387 minus.n21 a_n3654_n1288# 0.145204f
C388 minus.n22 a_n3654_n1288# 0.009072f
C389 minus.n23 a_n3654_n1288# 0.053345f
C390 minus.n24 a_n3654_n1288# 0.039978f
C391 minus.n25 a_n3654_n1288# 0.039978f
C392 minus.n26 a_n3654_n1288# 0.009072f
C393 minus.t18 a_n3654_n1288# 0.19808f
C394 minus.n27 a_n3654_n1288# 0.134037f
C395 minus.n28 a_n3654_n1288# 0.009072f
C396 minus.n29 a_n3654_n1288# 0.053345f
C397 minus.n30 a_n3654_n1288# 0.066588f
C398 minus.n31 a_n3654_n1288# 0.066588f
C399 minus.n32 a_n3654_n1288# 0.144711f
C400 minus.n33 a_n3654_n1288# 0.009072f
C401 minus.t10 a_n3654_n1288# 0.19808f
C402 minus.n34 a_n3654_n1288# 0.130709f
C403 minus.n35 a_n3654_n1288# 1.37837f
C404 minus.n36 a_n3654_n1288# 0.053345f
C405 minus.t7 a_n3654_n1288# 0.19808f
C406 minus.n37 a_n3654_n1288# 0.145697f
C407 minus.n38 a_n3654_n1288# 0.039978f
C408 minus.t4 a_n3654_n1288# 0.19808f
C409 minus.n39 a_n3654_n1288# 0.134037f
C410 minus.n40 a_n3654_n1288# 0.066588f
C411 minus.n41 a_n3654_n1288# 0.009072f
C412 minus.n42 a_n3654_n1288# 0.039978f
C413 minus.n43 a_n3654_n1288# 0.009072f
C414 minus.t22 a_n3654_n1288# 0.2206f
C415 minus.n44 a_n3654_n1288# 0.118686f
C416 minus.t1 a_n3654_n1288# 0.19808f
C417 minus.n45 a_n3654_n1288# 0.145676f
C418 minus.t23 a_n3654_n1288# 0.19808f
C419 minus.n46 a_n3654_n1288# 0.145697f
C420 minus.n47 a_n3654_n1288# 0.229777f
C421 minus.n48 a_n3654_n1288# 0.053345f
C422 minus.n49 a_n3654_n1288# 0.039978f
C423 minus.t2 a_n3654_n1288# 0.19808f
C424 minus.n50 a_n3654_n1288# 0.134037f
C425 minus.n51 a_n3654_n1288# 0.009072f
C426 minus.t14 a_n3654_n1288# 0.19808f
C427 minus.n52 a_n3654_n1288# 0.134037f
C428 minus.n53 a_n3654_n1288# 0.039978f
C429 minus.n54 a_n3654_n1288# 0.053345f
C430 minus.n55 a_n3654_n1288# 0.066588f
C431 minus.t3 a_n3654_n1288# 0.19808f
C432 minus.n56 a_n3654_n1288# 0.145204f
C433 minus.t16 a_n3654_n1288# 0.19808f
C434 minus.n57 a_n3654_n1288# 0.145204f
C435 minus.n58 a_n3654_n1288# 0.009072f
C436 minus.n59 a_n3654_n1288# 0.053345f
C437 minus.n60 a_n3654_n1288# 0.039978f
C438 minus.n61 a_n3654_n1288# 0.039978f
C439 minus.n62 a_n3654_n1288# 0.009072f
C440 minus.t20 a_n3654_n1288# 0.19808f
C441 minus.n63 a_n3654_n1288# 0.134037f
C442 minus.n64 a_n3654_n1288# 0.009072f
C443 minus.n65 a_n3654_n1288# 0.053345f
C444 minus.n66 a_n3654_n1288# 0.066588f
C445 minus.n67 a_n3654_n1288# 0.066588f
C446 minus.t0 a_n3654_n1288# 0.19808f
C447 minus.n68 a_n3654_n1288# 0.144711f
C448 minus.n69 a_n3654_n1288# 0.009072f
C449 minus.t6 a_n3654_n1288# 0.19808f
C450 minus.n70 a_n3654_n1288# 0.130709f
C451 minus.n71 a_n3654_n1288# 0.276283f
C452 minus.n72 a_n3654_n1288# 1.67223f
.ends

