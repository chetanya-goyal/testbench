* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t16 minus.t0 drain_right.t6 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X2 source.t18 plus.t0 drain_left.t9 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 source.t15 minus.t1 drain_right.t8 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X4 drain_left.t8 plus.t1 source.t19 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X5 source.t1 plus.t2 drain_left.t7 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X6 a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X7 drain_right.t1 minus.t2 source.t14 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X8 drain_right.t7 minus.t3 source.t13 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X9 drain_right.t9 minus.t4 source.t12 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X10 source.t0 plus.t3 drain_left.t6 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 drain_left.t5 plus.t4 source.t4 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X12 a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X13 a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X14 drain_right.t3 minus.t5 source.t11 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X15 source.t2 plus.t5 drain_left.t4 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X16 drain_right.t4 minus.t6 source.t10 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X17 source.t9 minus.t7 drain_right.t2 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X18 drain_left.t3 plus.t6 source.t6 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X19 drain_right.t5 minus.t8 source.t8 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X20 drain_left.t2 plus.t7 source.t3 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X21 source.t7 minus.t9 drain_right.t0 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X22 drain_left.t1 plus.t8 source.t17 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X23 drain_left.t0 plus.t9 source.t5 a_n1712_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
R0 minus.n2 minus.t5 195.948
R1 minus.n14 minus.t8 195.948
R2 minus.n3 minus.t1 174.966
R3 minus.n1 minus.t3 174.966
R4 minus.n9 minus.t7 174.966
R5 minus.n10 minus.t2 174.966
R6 minus.n15 minus.t0 174.966
R7 minus.n13 minus.t6 174.966
R8 minus.n21 minus.t9 174.966
R9 minus.n22 minus.t4 174.966
R10 minus.n11 minus.n10 161.3
R11 minus.n9 minus.n0 161.3
R12 minus.n8 minus.n7 161.3
R13 minus.n6 minus.n1 161.3
R14 minus.n5 minus.n4 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n18 minus.n13 161.3
R19 minus.n17 minus.n16 161.3
R20 minus.n5 minus.n2 70.4033
R21 minus.n17 minus.n14 70.4033
R22 minus.n10 minus.n9 48.2005
R23 minus.n22 minus.n21 48.2005
R24 minus.n4 minus.n1 36.5157
R25 minus.n8 minus.n1 36.5157
R26 minus.n16 minus.n13 36.5157
R27 minus.n20 minus.n13 36.5157
R28 minus.n24 minus.n11 28.0933
R29 minus.n3 minus.n2 20.9576
R30 minus.n15 minus.n14 20.9576
R31 minus.n4 minus.n3 11.6853
R32 minus.n9 minus.n8 11.6853
R33 minus.n16 minus.n15 11.6853
R34 minus.n21 minus.n20 11.6853
R35 minus.n24 minus.n23 6.563
R36 minus.n11 minus.n0 0.189894
R37 minus.n7 minus.n0 0.189894
R38 minus.n7 minus.n6 0.189894
R39 minus.n6 minus.n5 0.189894
R40 minus.n18 minus.n17 0.189894
R41 minus.n19 minus.n18 0.189894
R42 minus.n19 minus.n12 0.189894
R43 minus.n23 minus.n12 0.189894
R44 minus minus.n24 0.188
R45 drain_right.n2 drain_right.n0 289.615
R46 drain_right.n16 drain_right.n14 289.615
R47 drain_right.n3 drain_right.n2 185
R48 drain_right.n17 drain_right.n16 185
R49 drain_right.t5 drain_right.n1 167.117
R50 drain_right.t1 drain_right.n15 167.117
R51 drain_right.n13 drain_right.n11 101.511
R52 drain_right.n10 drain_right.n9 101.276
R53 drain_right.n13 drain_right.n12 100.796
R54 drain_right.n8 drain_right.n7 100.796
R55 drain_right.n2 drain_right.t5 52.3082
R56 drain_right.n16 drain_right.t1 52.3082
R57 drain_right.n8 drain_right.n6 48.8039
R58 drain_right.n21 drain_right.n20 48.0884
R59 drain_right drain_right.n10 22.279
R60 drain_right.n9 drain_right.t0 9.9005
R61 drain_right.n9 drain_right.t9 9.9005
R62 drain_right.n7 drain_right.t6 9.9005
R63 drain_right.n7 drain_right.t4 9.9005
R64 drain_right.n11 drain_right.t8 9.9005
R65 drain_right.n11 drain_right.t3 9.9005
R66 drain_right.n12 drain_right.t2 9.9005
R67 drain_right.n12 drain_right.t7 9.9005
R68 drain_right.n3 drain_right.n1 9.71174
R69 drain_right.n17 drain_right.n15 9.71174
R70 drain_right.n6 drain_right.n5 9.45567
R71 drain_right.n20 drain_right.n19 9.45567
R72 drain_right.n5 drain_right.n4 9.3005
R73 drain_right.n19 drain_right.n18 9.3005
R74 drain_right.n6 drain_right.n0 8.14595
R75 drain_right.n20 drain_right.n14 8.14595
R76 drain_right.n4 drain_right.n3 7.3702
R77 drain_right.n18 drain_right.n17 7.3702
R78 drain_right drain_right.n21 6.01097
R79 drain_right.n4 drain_right.n0 5.81868
R80 drain_right.n18 drain_right.n14 5.81868
R81 drain_right.n5 drain_right.n1 3.44771
R82 drain_right.n19 drain_right.n15 3.44771
R83 drain_right.n21 drain_right.n13 0.716017
R84 drain_right.n10 drain_right.n8 0.124033
R85 source.n42 source.n40 289.615
R86 source.n30 source.n28 289.615
R87 source.n2 source.n0 289.615
R88 source.n14 source.n12 289.615
R89 source.n43 source.n42 185
R90 source.n31 source.n30 185
R91 source.n3 source.n2 185
R92 source.n15 source.n14 185
R93 source.t12 source.n41 167.117
R94 source.t5 source.n29 167.117
R95 source.t3 source.n1 167.117
R96 source.t11 source.n13 167.117
R97 source.n9 source.n8 84.1169
R98 source.n11 source.n10 84.1169
R99 source.n21 source.n20 84.1169
R100 source.n23 source.n22 84.1169
R101 source.n39 source.n38 84.1168
R102 source.n37 source.n36 84.1168
R103 source.n27 source.n26 84.1168
R104 source.n25 source.n24 84.1168
R105 source.n42 source.t12 52.3082
R106 source.n30 source.t5 52.3082
R107 source.n2 source.t3 52.3082
R108 source.n14 source.t11 52.3082
R109 source.n47 source.n46 31.4096
R110 source.n35 source.n34 31.4096
R111 source.n7 source.n6 31.4096
R112 source.n19 source.n18 31.4096
R113 source.n25 source.n23 15.143
R114 source.n38 source.t10 9.9005
R115 source.n38 source.t7 9.9005
R116 source.n36 source.t8 9.9005
R117 source.n36 source.t16 9.9005
R118 source.n26 source.t6 9.9005
R119 source.n26 source.t18 9.9005
R120 source.n24 source.t4 9.9005
R121 source.n24 source.t1 9.9005
R122 source.n8 source.t17 9.9005
R123 source.n8 source.t0 9.9005
R124 source.n10 source.t19 9.9005
R125 source.n10 source.t2 9.9005
R126 source.n20 source.t13 9.9005
R127 source.n20 source.t15 9.9005
R128 source.n22 source.t14 9.9005
R129 source.n22 source.t9 9.9005
R130 source.n43 source.n41 9.71174
R131 source.n31 source.n29 9.71174
R132 source.n3 source.n1 9.71174
R133 source.n15 source.n13 9.71174
R134 source.n46 source.n45 9.45567
R135 source.n34 source.n33 9.45567
R136 source.n6 source.n5 9.45567
R137 source.n18 source.n17 9.45567
R138 source.n45 source.n44 9.3005
R139 source.n33 source.n32 9.3005
R140 source.n5 source.n4 9.3005
R141 source.n17 source.n16 9.3005
R142 source.n48 source.n7 8.8068
R143 source.n46 source.n40 8.14595
R144 source.n34 source.n28 8.14595
R145 source.n6 source.n0 8.14595
R146 source.n18 source.n12 8.14595
R147 source.n44 source.n43 7.3702
R148 source.n32 source.n31 7.3702
R149 source.n4 source.n3 7.3702
R150 source.n16 source.n15 7.3702
R151 source.n44 source.n40 5.81868
R152 source.n32 source.n28 5.81868
R153 source.n4 source.n0 5.81868
R154 source.n16 source.n12 5.81868
R155 source.n48 source.n47 5.62119
R156 source.n45 source.n41 3.44771
R157 source.n33 source.n29 3.44771
R158 source.n5 source.n1 3.44771
R159 source.n17 source.n13 3.44771
R160 source.n19 source.n11 0.828086
R161 source.n37 source.n35 0.828086
R162 source.n23 source.n21 0.716017
R163 source.n21 source.n19 0.716017
R164 source.n11 source.n9 0.716017
R165 source.n9 source.n7 0.716017
R166 source.n27 source.n25 0.716017
R167 source.n35 source.n27 0.716017
R168 source.n39 source.n37 0.716017
R169 source.n47 source.n39 0.716017
R170 source source.n48 0.188
R171 plus.n2 plus.t1 195.948
R172 plus.n14 plus.t9 195.948
R173 plus.n10 plus.t7 174.966
R174 plus.n9 plus.t3 174.966
R175 plus.n1 plus.t8 174.966
R176 plus.n3 plus.t5 174.966
R177 plus.n22 plus.t4 174.966
R178 plus.n21 plus.t2 174.966
R179 plus.n13 plus.t6 174.966
R180 plus.n15 plus.t0 174.966
R181 plus.n5 plus.n4 161.3
R182 plus.n6 plus.n1 161.3
R183 plus.n8 plus.n7 161.3
R184 plus.n9 plus.n0 161.3
R185 plus.n11 plus.n10 161.3
R186 plus.n17 plus.n16 161.3
R187 plus.n18 plus.n13 161.3
R188 plus.n20 plus.n19 161.3
R189 plus.n21 plus.n12 161.3
R190 plus.n23 plus.n22 161.3
R191 plus.n5 plus.n2 70.4033
R192 plus.n17 plus.n14 70.4033
R193 plus.n10 plus.n9 48.2005
R194 plus.n22 plus.n21 48.2005
R195 plus.n8 plus.n1 36.5157
R196 plus.n4 plus.n1 36.5157
R197 plus.n20 plus.n13 36.5157
R198 plus.n16 plus.n13 36.5157
R199 plus plus.n23 25.7623
R200 plus.n3 plus.n2 20.9576
R201 plus.n15 plus.n14 20.9576
R202 plus.n9 plus.n8 11.6853
R203 plus.n4 plus.n3 11.6853
R204 plus.n21 plus.n20 11.6853
R205 plus.n16 plus.n15 11.6853
R206 plus plus.n11 8.41906
R207 plus.n6 plus.n5 0.189894
R208 plus.n7 plus.n6 0.189894
R209 plus.n7 plus.n0 0.189894
R210 plus.n11 plus.n0 0.189894
R211 plus.n23 plus.n12 0.189894
R212 plus.n19 plus.n12 0.189894
R213 plus.n19 plus.n18 0.189894
R214 plus.n18 plus.n17 0.189894
R215 drain_left.n2 drain_left.n0 289.615
R216 drain_left.n13 drain_left.n11 289.615
R217 drain_left.n3 drain_left.n2 185
R218 drain_left.n14 drain_left.n13 185
R219 drain_left.t5 drain_left.n1 167.117
R220 drain_left.t8 drain_left.n12 167.117
R221 drain_left.n10 drain_left.n9 101.276
R222 drain_left.n21 drain_left.n20 100.796
R223 drain_left.n19 drain_left.n18 100.796
R224 drain_left.n8 drain_left.n7 100.796
R225 drain_left.n2 drain_left.t5 52.3082
R226 drain_left.n13 drain_left.t8 52.3082
R227 drain_left.n8 drain_left.n6 48.8039
R228 drain_left.n19 drain_left.n17 48.8039
R229 drain_left drain_left.n10 22.8323
R230 drain_left.n9 drain_left.t9 9.9005
R231 drain_left.n9 drain_left.t0 9.9005
R232 drain_left.n7 drain_left.t7 9.9005
R233 drain_left.n7 drain_left.t3 9.9005
R234 drain_left.n20 drain_left.t6 9.9005
R235 drain_left.n20 drain_left.t2 9.9005
R236 drain_left.n18 drain_left.t4 9.9005
R237 drain_left.n18 drain_left.t1 9.9005
R238 drain_left.n3 drain_left.n1 9.71174
R239 drain_left.n14 drain_left.n12 9.71174
R240 drain_left.n6 drain_left.n5 9.45567
R241 drain_left.n17 drain_left.n16 9.45567
R242 drain_left.n5 drain_left.n4 9.3005
R243 drain_left.n16 drain_left.n15 9.3005
R244 drain_left.n6 drain_left.n0 8.14595
R245 drain_left.n17 drain_left.n11 8.14595
R246 drain_left.n4 drain_left.n3 7.3702
R247 drain_left.n15 drain_left.n14 7.3702
R248 drain_left drain_left.n21 6.36873
R249 drain_left.n4 drain_left.n0 5.81868
R250 drain_left.n15 drain_left.n11 5.81868
R251 drain_left.n5 drain_left.n1 3.44771
R252 drain_left.n16 drain_left.n12 3.44771
R253 drain_left.n21 drain_left.n19 0.716017
R254 drain_left.n10 drain_left.n8 0.124033
C0 drain_right source 4.73486f
C1 drain_right drain_left 0.843613f
C2 drain_left source 4.73642f
C3 drain_right minus 1.27063f
C4 minus source 1.51072f
C5 minus drain_left 0.17817f
C6 drain_right plus 0.327566f
C7 plus source 1.52478f
C8 plus drain_left 1.43545f
C9 minus plus 3.4383f
C10 drain_right a_n1712_n1288# 3.60592f
C11 drain_left a_n1712_n1288# 3.8381f
C12 source a_n1712_n1288# 2.533259f
C13 minus a_n1712_n1288# 5.852321f
C14 plus a_n1712_n1288# 6.422613f
C15 drain_left.n0 a_n1712_n1288# 0.028669f
C16 drain_left.n1 a_n1712_n1288# 0.063434f
C17 drain_left.t5 a_n1712_n1288# 0.047604f
C18 drain_left.n2 a_n1712_n1288# 0.049646f
C19 drain_left.n3 a_n1712_n1288# 0.016004f
C20 drain_left.n4 a_n1712_n1288# 0.010555f
C21 drain_left.n5 a_n1712_n1288# 0.139823f
C22 drain_left.n6 a_n1712_n1288# 0.046209f
C23 drain_left.t7 a_n1712_n1288# 0.031044f
C24 drain_left.t3 a_n1712_n1288# 0.031044f
C25 drain_left.n7 a_n1712_n1288# 0.195026f
C26 drain_left.n8 a_n1712_n1288# 0.288415f
C27 drain_left.t9 a_n1712_n1288# 0.031044f
C28 drain_left.t0 a_n1712_n1288# 0.031044f
C29 drain_left.n9 a_n1712_n1288# 0.196142f
C30 drain_left.n10 a_n1712_n1288# 0.776332f
C31 drain_left.n11 a_n1712_n1288# 0.028669f
C32 drain_left.n12 a_n1712_n1288# 0.063434f
C33 drain_left.t8 a_n1712_n1288# 0.047604f
C34 drain_left.n13 a_n1712_n1288# 0.049646f
C35 drain_left.n14 a_n1712_n1288# 0.016004f
C36 drain_left.n15 a_n1712_n1288# 0.010555f
C37 drain_left.n16 a_n1712_n1288# 0.139823f
C38 drain_left.n17 a_n1712_n1288# 0.046209f
C39 drain_left.t4 a_n1712_n1288# 0.031044f
C40 drain_left.t1 a_n1712_n1288# 0.031044f
C41 drain_left.n18 a_n1712_n1288# 0.195027f
C42 drain_left.n19 a_n1712_n1288# 0.322196f
C43 drain_left.t6 a_n1712_n1288# 0.031044f
C44 drain_left.t2 a_n1712_n1288# 0.031044f
C45 drain_left.n20 a_n1712_n1288# 0.195027f
C46 drain_left.n21 a_n1712_n1288# 0.409664f
C47 plus.n0 a_n1712_n1288# 0.027362f
C48 plus.t7 a_n1712_n1288# 0.084732f
C49 plus.t3 a_n1712_n1288# 0.084732f
C50 plus.t8 a_n1712_n1288# 0.084732f
C51 plus.n1 a_n1712_n1288# 0.063903f
C52 plus.t1 a_n1712_n1288# 0.091271f
C53 plus.n2 a_n1712_n1288# 0.054696f
C54 plus.t5 a_n1712_n1288# 0.084732f
C55 plus.n3 a_n1712_n1288# 0.062385f
C56 plus.n4 a_n1712_n1288# 0.006209f
C57 plus.n5 a_n1712_n1288# 0.087283f
C58 plus.n6 a_n1712_n1288# 0.027362f
C59 plus.n7 a_n1712_n1288# 0.027362f
C60 plus.n8 a_n1712_n1288# 0.006209f
C61 plus.n9 a_n1712_n1288# 0.062385f
C62 plus.n10 a_n1712_n1288# 0.061035f
C63 plus.n11 a_n1712_n1288# 0.199875f
C64 plus.n12 a_n1712_n1288# 0.027362f
C65 plus.t4 a_n1712_n1288# 0.084732f
C66 plus.t2 a_n1712_n1288# 0.084732f
C67 plus.t6 a_n1712_n1288# 0.084732f
C68 plus.n13 a_n1712_n1288# 0.063903f
C69 plus.t9 a_n1712_n1288# 0.091271f
C70 plus.n14 a_n1712_n1288# 0.054696f
C71 plus.t0 a_n1712_n1288# 0.084732f
C72 plus.n15 a_n1712_n1288# 0.062385f
C73 plus.n16 a_n1712_n1288# 0.006209f
C74 plus.n17 a_n1712_n1288# 0.087283f
C75 plus.n18 a_n1712_n1288# 0.027362f
C76 plus.n19 a_n1712_n1288# 0.027362f
C77 plus.n20 a_n1712_n1288# 0.006209f
C78 plus.n21 a_n1712_n1288# 0.062385f
C79 plus.n22 a_n1712_n1288# 0.061035f
C80 plus.n23 a_n1712_n1288# 0.608842f
C81 source.n0 a_n1712_n1288# 0.035974f
C82 source.n1 a_n1712_n1288# 0.079596f
C83 source.t3 a_n1712_n1288# 0.059733f
C84 source.n2 a_n1712_n1288# 0.062295f
C85 source.n3 a_n1712_n1288# 0.020081f
C86 source.n4 a_n1712_n1288# 0.013244f
C87 source.n5 a_n1712_n1288# 0.175449f
C88 source.n6 a_n1712_n1288# 0.039435f
C89 source.n7 a_n1712_n1288# 0.396423f
C90 source.t17 a_n1712_n1288# 0.038953f
C91 source.t0 a_n1712_n1288# 0.038953f
C92 source.n8 a_n1712_n1288# 0.208243f
C93 source.n9 a_n1712_n1288# 0.305266f
C94 source.t19 a_n1712_n1288# 0.038953f
C95 source.t2 a_n1712_n1288# 0.038953f
C96 source.n10 a_n1712_n1288# 0.208243f
C97 source.n11 a_n1712_n1288# 0.314167f
C98 source.n12 a_n1712_n1288# 0.035974f
C99 source.n13 a_n1712_n1288# 0.079596f
C100 source.t11 a_n1712_n1288# 0.059733f
C101 source.n14 a_n1712_n1288# 0.062295f
C102 source.n15 a_n1712_n1288# 0.020081f
C103 source.n16 a_n1712_n1288# 0.013244f
C104 source.n17 a_n1712_n1288# 0.175449f
C105 source.n18 a_n1712_n1288# 0.039435f
C106 source.n19 a_n1712_n1288# 0.14284f
C107 source.t13 a_n1712_n1288# 0.038953f
C108 source.t15 a_n1712_n1288# 0.038953f
C109 source.n20 a_n1712_n1288# 0.208243f
C110 source.n21 a_n1712_n1288# 0.305266f
C111 source.t14 a_n1712_n1288# 0.038953f
C112 source.t9 a_n1712_n1288# 0.038953f
C113 source.n22 a_n1712_n1288# 0.208243f
C114 source.n23 a_n1712_n1288# 0.857446f
C115 source.t4 a_n1712_n1288# 0.038953f
C116 source.t1 a_n1712_n1288# 0.038953f
C117 source.n24 a_n1712_n1288# 0.208242f
C118 source.n25 a_n1712_n1288# 0.857447f
C119 source.t6 a_n1712_n1288# 0.038953f
C120 source.t18 a_n1712_n1288# 0.038953f
C121 source.n26 a_n1712_n1288# 0.208242f
C122 source.n27 a_n1712_n1288# 0.305268f
C123 source.n28 a_n1712_n1288# 0.035974f
C124 source.n29 a_n1712_n1288# 0.079596f
C125 source.t5 a_n1712_n1288# 0.059733f
C126 source.n30 a_n1712_n1288# 0.062295f
C127 source.n31 a_n1712_n1288# 0.020081f
C128 source.n32 a_n1712_n1288# 0.013244f
C129 source.n33 a_n1712_n1288# 0.175449f
C130 source.n34 a_n1712_n1288# 0.039435f
C131 source.n35 a_n1712_n1288# 0.14284f
C132 source.t8 a_n1712_n1288# 0.038953f
C133 source.t16 a_n1712_n1288# 0.038953f
C134 source.n36 a_n1712_n1288# 0.208242f
C135 source.n37 a_n1712_n1288# 0.314168f
C136 source.t10 a_n1712_n1288# 0.038953f
C137 source.t7 a_n1712_n1288# 0.038953f
C138 source.n38 a_n1712_n1288# 0.208242f
C139 source.n39 a_n1712_n1288# 0.305268f
C140 source.n40 a_n1712_n1288# 0.035974f
C141 source.n41 a_n1712_n1288# 0.079596f
C142 source.t12 a_n1712_n1288# 0.059733f
C143 source.n42 a_n1712_n1288# 0.062295f
C144 source.n43 a_n1712_n1288# 0.020081f
C145 source.n44 a_n1712_n1288# 0.013244f
C146 source.n45 a_n1712_n1288# 0.175449f
C147 source.n46 a_n1712_n1288# 0.039435f
C148 source.n47 a_n1712_n1288# 0.264439f
C149 source.n48 a_n1712_n1288# 0.615257f
C150 drain_right.n0 a_n1712_n1288# 0.029145f
C151 drain_right.n1 a_n1712_n1288# 0.064488f
C152 drain_right.t5 a_n1712_n1288# 0.048395f
C153 drain_right.n2 a_n1712_n1288# 0.050471f
C154 drain_right.n3 a_n1712_n1288# 0.01627f
C155 drain_right.n4 a_n1712_n1288# 0.01073f
C156 drain_right.n5 a_n1712_n1288# 0.142147f
C157 drain_right.n6 a_n1712_n1288# 0.046976f
C158 drain_right.t6 a_n1712_n1288# 0.03156f
C159 drain_right.t4 a_n1712_n1288# 0.03156f
C160 drain_right.n7 a_n1712_n1288# 0.198267f
C161 drain_right.n8 a_n1712_n1288# 0.293209f
C162 drain_right.t0 a_n1712_n1288# 0.03156f
C163 drain_right.t9 a_n1712_n1288# 0.03156f
C164 drain_right.n9 a_n1712_n1288# 0.199402f
C165 drain_right.n10 a_n1712_n1288# 0.750059f
C166 drain_right.t8 a_n1712_n1288# 0.03156f
C167 drain_right.t3 a_n1712_n1288# 0.03156f
C168 drain_right.n11 a_n1712_n1288# 0.200051f
C169 drain_right.t2 a_n1712_n1288# 0.03156f
C170 drain_right.t7 a_n1712_n1288# 0.03156f
C171 drain_right.n12 a_n1712_n1288# 0.198268f
C172 drain_right.n13 a_n1712_n1288# 0.49609f
C173 drain_right.n14 a_n1712_n1288# 0.029145f
C174 drain_right.n15 a_n1712_n1288# 0.064488f
C175 drain_right.t1 a_n1712_n1288# 0.048395f
C176 drain_right.n16 a_n1712_n1288# 0.050471f
C177 drain_right.n17 a_n1712_n1288# 0.01627f
C178 drain_right.n18 a_n1712_n1288# 0.01073f
C179 drain_right.n19 a_n1712_n1288# 0.142147f
C180 drain_right.n20 a_n1712_n1288# 0.045747f
C181 drain_right.n21 a_n1712_n1288# 0.258962f
C182 minus.n0 a_n1712_n1288# 0.026924f
C183 minus.t3 a_n1712_n1288# 0.083375f
C184 minus.n1 a_n1712_n1288# 0.06288f
C185 minus.t5 a_n1712_n1288# 0.08981f
C186 minus.n2 a_n1712_n1288# 0.05382f
C187 minus.t1 a_n1712_n1288# 0.083375f
C188 minus.n3 a_n1712_n1288# 0.061386f
C189 minus.n4 a_n1712_n1288# 0.00611f
C190 minus.n5 a_n1712_n1288# 0.085886f
C191 minus.n6 a_n1712_n1288# 0.026924f
C192 minus.n7 a_n1712_n1288# 0.026924f
C193 minus.n8 a_n1712_n1288# 0.00611f
C194 minus.t7 a_n1712_n1288# 0.083375f
C195 minus.n9 a_n1712_n1288# 0.061386f
C196 minus.t2 a_n1712_n1288# 0.083375f
C197 minus.n10 a_n1712_n1288# 0.060058f
C198 minus.n11 a_n1712_n1288# 0.626582f
C199 minus.n12 a_n1712_n1288# 0.026924f
C200 minus.t6 a_n1712_n1288# 0.083375f
C201 minus.n13 a_n1712_n1288# 0.06288f
C202 minus.t8 a_n1712_n1288# 0.08981f
C203 minus.n14 a_n1712_n1288# 0.05382f
C204 minus.t0 a_n1712_n1288# 0.083375f
C205 minus.n15 a_n1712_n1288# 0.061386f
C206 minus.n16 a_n1712_n1288# 0.00611f
C207 minus.n17 a_n1712_n1288# 0.085886f
C208 minus.n18 a_n1712_n1288# 0.026924f
C209 minus.n19 a_n1712_n1288# 0.026924f
C210 minus.n20 a_n1712_n1288# 0.00611f
C211 minus.t9 a_n1712_n1288# 0.083375f
C212 minus.n21 a_n1712_n1288# 0.061386f
C213 minus.t4 a_n1712_n1288# 0.083375f
C214 minus.n22 a_n1712_n1288# 0.060058f
C215 minus.n23 a_n1712_n1288# 0.180004f
C216 minus.n24 a_n1712_n1288# 0.772303f
.ends

