* NGSPICE file created from diffpair199.ext - technology: sky130A

.subckt diffpair199 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t22 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 source.t9 plus.t0 drain_left.t23 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X2 drain_right.t2 minus.t1 source.t46 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X3 drain_left.t22 plus.t1 source.t4 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X4 drain_left.t21 plus.t2 source.t10 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X5 source.t45 minus.t2 drain_right.t0 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X6 drain_right.t1 minus.t3 source.t44 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X7 drain_left.t20 plus.t3 source.t14 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X8 drain_right.t23 minus.t4 source.t43 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X9 drain_right.t3 minus.t5 source.t42 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X10 source.t41 minus.t6 drain_right.t4 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X11 source.t40 minus.t7 drain_right.t5 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X12 source.t6 plus.t4 drain_left.t19 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X13 source.t19 plus.t5 drain_left.t18 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X14 a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X15 drain_left.t17 plus.t6 source.t23 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X16 drain_left.t16 plus.t7 source.t13 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X17 a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X18 drain_right.t6 minus.t8 source.t39 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X19 drain_left.t15 plus.t8 source.t0 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X20 source.t38 minus.t9 drain_right.t7 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X21 drain_right.t8 minus.t10 source.t37 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X22 source.t36 minus.t11 drain_right.t9 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X23 source.t20 plus.t9 drain_left.t14 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X24 a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X25 source.t12 plus.t10 drain_left.t13 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X26 drain_left.t12 plus.t11 source.t16 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X27 drain_right.t10 minus.t12 source.t35 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X28 source.t34 minus.t13 drain_right.t11 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X29 drain_left.t11 plus.t12 source.t21 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X30 source.t1 plus.t13 drain_left.t10 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X31 drain_right.t12 minus.t14 source.t33 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X32 drain_right.t13 minus.t15 source.t32 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X33 drain_left.t9 plus.t14 source.t8 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X34 source.t11 plus.t15 drain_left.t8 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X35 source.t31 minus.t16 drain_right.t14 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X36 source.t15 plus.t16 drain_left.t7 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X37 source.t30 minus.t17 drain_right.t15 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X38 drain_left.t6 plus.t17 source.t5 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X39 drain_left.t5 plus.t18 source.t3 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X40 drain_right.t16 minus.t18 source.t29 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X41 drain_right.t19 minus.t19 source.t28 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X42 a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X43 source.t27 minus.t20 drain_right.t20 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X44 source.t26 minus.t21 drain_right.t17 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X45 drain_right.t21 minus.t22 source.t25 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X46 source.t24 minus.t23 drain_right.t18 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X47 source.t18 plus.t19 drain_left.t4 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X48 source.t17 plus.t20 drain_left.t3 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X49 source.t22 plus.t21 drain_left.t2 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X50 source.t2 plus.t22 drain_left.t1 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X51 drain_left.t0 plus.t23 source.t7 a_n2354_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n35 minus.t6 376.837
R1 minus.n9 minus.t14 376.837
R2 minus.n72 minus.t10 376.837
R3 minus.n46 minus.t11 376.837
R4 minus.n34 minus.t19 345.433
R5 minus.n1 minus.t9 345.433
R6 minus.n28 minus.t5 345.433
R7 minus.n26 minus.t21 345.433
R8 minus.n3 minus.t8 345.433
R9 minus.n20 minus.t2 345.433
R10 minus.n5 minus.t18 345.433
R11 minus.n15 minus.t13 345.433
R12 minus.n13 minus.t4 345.433
R13 minus.n8 minus.t20 345.433
R14 minus.n71 minus.t17 345.433
R15 minus.n38 minus.t22 345.433
R16 minus.n65 minus.t0 345.433
R17 minus.n63 minus.t15 345.433
R18 minus.n40 minus.t16 345.433
R19 minus.n57 minus.t3 345.433
R20 minus.n42 minus.t7 345.433
R21 minus.n52 minus.t12 345.433
R22 minus.n50 minus.t23 345.433
R23 minus.n45 minus.t1 345.433
R24 minus.n10 minus.n9 161.489
R25 minus.n47 minus.n46 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n32 minus.n31 161.3
R29 minus.n30 minus.n29 161.3
R30 minus.n27 minus.n2 161.3
R31 minus.n25 minus.n24 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n19 minus.n18 161.3
R35 minus.n17 minus.n16 161.3
R36 minus.n14 minus.n6 161.3
R37 minus.n12 minus.n11 161.3
R38 minus.n10 minus.n7 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n69 minus.n68 161.3
R42 minus.n67 minus.n66 161.3
R43 minus.n64 minus.n39 161.3
R44 minus.n62 minus.n61 161.3
R45 minus.n60 minus.n59 161.3
R46 minus.n58 minus.n41 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n54 minus.n53 161.3
R49 minus.n51 minus.n43 161.3
R50 minus.n49 minus.n48 161.3
R51 minus.n47 minus.n44 161.3
R52 minus.n33 minus.n32 73.0308
R53 minus.n22 minus.n21 73.0308
R54 minus.n12 minus.n7 73.0308
R55 minus.n49 minus.n44 73.0308
R56 minus.n59 minus.n58 73.0308
R57 minus.n70 minus.n69 73.0308
R58 minus.n29 minus.n1 66.4581
R59 minus.n14 minus.n13 66.4581
R60 minus.n51 minus.n50 66.4581
R61 minus.n66 minus.n38 66.4581
R62 minus.n25 minus.n3 63.5369
R63 minus.n20 minus.n19 63.5369
R64 minus.n57 minus.n56 63.5369
R65 minus.n62 minus.n40 63.5369
R66 minus.n35 minus.n34 60.6157
R67 minus.n9 minus.n8 60.6157
R68 minus.n46 minus.n45 60.6157
R69 minus.n72 minus.n71 60.6157
R70 minus.n28 minus.n27 47.4702
R71 minus.n16 minus.n15 47.4702
R72 minus.n53 minus.n52 47.4702
R73 minus.n65 minus.n64 47.4702
R74 minus.n27 minus.n26 44.549
R75 minus.n16 minus.n5 44.549
R76 minus.n53 minus.n42 44.549
R77 minus.n64 minus.n63 44.549
R78 minus.n74 minus.n36 31.1899
R79 minus.n26 minus.n25 28.4823
R80 minus.n19 minus.n5 28.4823
R81 minus.n56 minus.n42 28.4823
R82 minus.n63 minus.n62 28.4823
R83 minus.n29 minus.n28 25.5611
R84 minus.n15 minus.n14 25.5611
R85 minus.n52 minus.n51 25.5611
R86 minus.n66 minus.n65 25.5611
R87 minus.n34 minus.n33 12.4157
R88 minus.n8 minus.n7 12.4157
R89 minus.n45 minus.n44 12.4157
R90 minus.n71 minus.n70 12.4157
R91 minus.n22 minus.n3 9.49444
R92 minus.n21 minus.n20 9.49444
R93 minus.n58 minus.n57 9.49444
R94 minus.n59 minus.n40 9.49444
R95 minus.n32 minus.n1 6.57323
R96 minus.n13 minus.n12 6.57323
R97 minus.n50 minus.n49 6.57323
R98 minus.n69 minus.n38 6.57323
R99 minus.n74 minus.n73 6.4702
R100 minus.n36 minus.n0 0.189894
R101 minus.n31 minus.n0 0.189894
R102 minus.n31 minus.n30 0.189894
R103 minus.n30 minus.n2 0.189894
R104 minus.n24 minus.n2 0.189894
R105 minus.n24 minus.n23 0.189894
R106 minus.n23 minus.n4 0.189894
R107 minus.n18 minus.n4 0.189894
R108 minus.n18 minus.n17 0.189894
R109 minus.n17 minus.n6 0.189894
R110 minus.n11 minus.n6 0.189894
R111 minus.n11 minus.n10 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n48 minus.n43 0.189894
R114 minus.n54 minus.n43 0.189894
R115 minus.n55 minus.n54 0.189894
R116 minus.n55 minus.n41 0.189894
R117 minus.n60 minus.n41 0.189894
R118 minus.n61 minus.n60 0.189894
R119 minus.n61 minus.n39 0.189894
R120 minus.n67 minus.n39 0.189894
R121 minus.n68 minus.n67 0.189894
R122 minus.n68 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 drain_right.n13 drain_right.n11 80.3162
R126 drain_right.n7 drain_right.n5 80.3161
R127 drain_right.n2 drain_right.n0 80.3161
R128 drain_right.n13 drain_right.n12 79.7731
R129 drain_right.n15 drain_right.n14 79.7731
R130 drain_right.n17 drain_right.n16 79.7731
R131 drain_right.n19 drain_right.n18 79.7731
R132 drain_right.n21 drain_right.n20 79.7731
R133 drain_right.n7 drain_right.n6 79.773
R134 drain_right.n9 drain_right.n8 79.773
R135 drain_right.n4 drain_right.n3 79.773
R136 drain_right.n2 drain_right.n1 79.773
R137 drain_right drain_right.n10 25.1551
R138 drain_right.n5 drain_right.t15 6.6005
R139 drain_right.n5 drain_right.t8 6.6005
R140 drain_right.n6 drain_right.t22 6.6005
R141 drain_right.n6 drain_right.t21 6.6005
R142 drain_right.n8 drain_right.t14 6.6005
R143 drain_right.n8 drain_right.t13 6.6005
R144 drain_right.n3 drain_right.t5 6.6005
R145 drain_right.n3 drain_right.t1 6.6005
R146 drain_right.n1 drain_right.t18 6.6005
R147 drain_right.n1 drain_right.t10 6.6005
R148 drain_right.n0 drain_right.t9 6.6005
R149 drain_right.n0 drain_right.t2 6.6005
R150 drain_right.n11 drain_right.t20 6.6005
R151 drain_right.n11 drain_right.t12 6.6005
R152 drain_right.n12 drain_right.t11 6.6005
R153 drain_right.n12 drain_right.t23 6.6005
R154 drain_right.n14 drain_right.t0 6.6005
R155 drain_right.n14 drain_right.t16 6.6005
R156 drain_right.n16 drain_right.t17 6.6005
R157 drain_right.n16 drain_right.t6 6.6005
R158 drain_right.n18 drain_right.t7 6.6005
R159 drain_right.n18 drain_right.t3 6.6005
R160 drain_right.n20 drain_right.t4 6.6005
R161 drain_right.n20 drain_right.t19 6.6005
R162 drain_right drain_right.n21 6.19632
R163 drain_right.n9 drain_right.n7 0.543603
R164 drain_right.n4 drain_right.n2 0.543603
R165 drain_right.n21 drain_right.n19 0.543603
R166 drain_right.n19 drain_right.n17 0.543603
R167 drain_right.n17 drain_right.n15 0.543603
R168 drain_right.n15 drain_right.n13 0.543603
R169 drain_right.n10 drain_right.n9 0.216706
R170 drain_right.n10 drain_right.n4 0.216706
R171 source.n0 source.t23 69.6943
R172 source.n11 source.t19 69.6943
R173 source.n12 source.t33 69.6943
R174 source.n23 source.t41 69.6943
R175 source.n47 source.t37 69.6942
R176 source.n36 source.t36 69.6942
R177 source.n35 source.t13 69.6942
R178 source.n24 source.t2 69.6942
R179 source.n2 source.n1 63.0943
R180 source.n4 source.n3 63.0943
R181 source.n6 source.n5 63.0943
R182 source.n8 source.n7 63.0943
R183 source.n10 source.n9 63.0943
R184 source.n14 source.n13 63.0943
R185 source.n16 source.n15 63.0943
R186 source.n18 source.n17 63.0943
R187 source.n20 source.n19 63.0943
R188 source.n22 source.n21 63.0943
R189 source.n46 source.n45 63.0942
R190 source.n44 source.n43 63.0942
R191 source.n42 source.n41 63.0942
R192 source.n40 source.n39 63.0942
R193 source.n38 source.n37 63.0942
R194 source.n34 source.n33 63.0942
R195 source.n32 source.n31 63.0942
R196 source.n30 source.n29 63.0942
R197 source.n28 source.n27 63.0942
R198 source.n26 source.n25 63.0942
R199 source.n24 source.n23 15.0126
R200 source.n48 source.n0 9.47816
R201 source.n45 source.t25 6.6005
R202 source.n45 source.t30 6.6005
R203 source.n43 source.t32 6.6005
R204 source.n43 source.t47 6.6005
R205 source.n41 source.t44 6.6005
R206 source.n41 source.t31 6.6005
R207 source.n39 source.t35 6.6005
R208 source.n39 source.t40 6.6005
R209 source.n37 source.t46 6.6005
R210 source.n37 source.t24 6.6005
R211 source.n33 source.t5 6.6005
R212 source.n33 source.t18 6.6005
R213 source.n31 source.t14 6.6005
R214 source.n31 source.t12 6.6005
R215 source.n29 source.t21 6.6005
R216 source.n29 source.t22 6.6005
R217 source.n27 source.t4 6.6005
R218 source.n27 source.t6 6.6005
R219 source.n25 source.t0 6.6005
R220 source.n25 source.t11 6.6005
R221 source.n1 source.t3 6.6005
R222 source.n1 source.t9 6.6005
R223 source.n3 source.t10 6.6005
R224 source.n3 source.t1 6.6005
R225 source.n5 source.t8 6.6005
R226 source.n5 source.t17 6.6005
R227 source.n7 source.t7 6.6005
R228 source.n7 source.t20 6.6005
R229 source.n9 source.t16 6.6005
R230 source.n9 source.t15 6.6005
R231 source.n13 source.t43 6.6005
R232 source.n13 source.t27 6.6005
R233 source.n15 source.t29 6.6005
R234 source.n15 source.t34 6.6005
R235 source.n17 source.t39 6.6005
R236 source.n17 source.t45 6.6005
R237 source.n19 source.t42 6.6005
R238 source.n19 source.t26 6.6005
R239 source.n21 source.t28 6.6005
R240 source.n21 source.t38 6.6005
R241 source.n48 source.n47 5.53498
R242 source.n23 source.n22 0.543603
R243 source.n22 source.n20 0.543603
R244 source.n20 source.n18 0.543603
R245 source.n18 source.n16 0.543603
R246 source.n16 source.n14 0.543603
R247 source.n14 source.n12 0.543603
R248 source.n11 source.n10 0.543603
R249 source.n10 source.n8 0.543603
R250 source.n8 source.n6 0.543603
R251 source.n6 source.n4 0.543603
R252 source.n4 source.n2 0.543603
R253 source.n2 source.n0 0.543603
R254 source.n26 source.n24 0.543603
R255 source.n28 source.n26 0.543603
R256 source.n30 source.n28 0.543603
R257 source.n32 source.n30 0.543603
R258 source.n34 source.n32 0.543603
R259 source.n35 source.n34 0.543603
R260 source.n38 source.n36 0.543603
R261 source.n40 source.n38 0.543603
R262 source.n42 source.n40 0.543603
R263 source.n44 source.n42 0.543603
R264 source.n46 source.n44 0.543603
R265 source.n47 source.n46 0.543603
R266 source.n12 source.n11 0.470328
R267 source.n36 source.n35 0.470328
R268 source source.n48 0.188
R269 plus.n9 plus.t5 376.837
R270 plus.n35 plus.t6 376.837
R271 plus.n46 plus.t7 376.837
R272 plus.n72 plus.t22 376.837
R273 plus.n8 plus.t11 345.433
R274 plus.n13 plus.t16 345.433
R275 plus.n15 plus.t23 345.433
R276 plus.n5 plus.t9 345.433
R277 plus.n20 plus.t14 345.433
R278 plus.n3 plus.t20 345.433
R279 plus.n26 plus.t2 345.433
R280 plus.n28 plus.t13 345.433
R281 plus.n1 plus.t18 345.433
R282 plus.n34 plus.t0 345.433
R283 plus.n45 plus.t19 345.433
R284 plus.n50 plus.t17 345.433
R285 plus.n52 plus.t10 345.433
R286 plus.n42 plus.t3 345.433
R287 plus.n57 plus.t21 345.433
R288 plus.n40 plus.t12 345.433
R289 plus.n63 plus.t4 345.433
R290 plus.n65 plus.t1 345.433
R291 plus.n38 plus.t15 345.433
R292 plus.n71 plus.t8 345.433
R293 plus.n10 plus.n9 161.489
R294 plus.n47 plus.n46 161.489
R295 plus.n10 plus.n7 161.3
R296 plus.n12 plus.n11 161.3
R297 plus.n14 plus.n6 161.3
R298 plus.n17 plus.n16 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n21 plus.n4 161.3
R301 plus.n23 plus.n22 161.3
R302 plus.n25 plus.n24 161.3
R303 plus.n27 plus.n2 161.3
R304 plus.n30 plus.n29 161.3
R305 plus.n32 plus.n31 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n47 plus.n44 161.3
R309 plus.n49 plus.n48 161.3
R310 plus.n51 plus.n43 161.3
R311 plus.n54 plus.n53 161.3
R312 plus.n56 plus.n55 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n61 161.3
R316 plus.n64 plus.n39 161.3
R317 plus.n67 plus.n66 161.3
R318 plus.n69 plus.n68 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n12 plus.n7 73.0308
R322 plus.n22 plus.n21 73.0308
R323 plus.n33 plus.n32 73.0308
R324 plus.n70 plus.n69 73.0308
R325 plus.n59 plus.n58 73.0308
R326 plus.n49 plus.n44 73.0308
R327 plus.n14 plus.n13 66.4581
R328 plus.n29 plus.n1 66.4581
R329 plus.n66 plus.n38 66.4581
R330 plus.n51 plus.n50 66.4581
R331 plus.n20 plus.n19 63.5369
R332 plus.n25 plus.n3 63.5369
R333 plus.n62 plus.n40 63.5369
R334 plus.n57 plus.n56 63.5369
R335 plus.n9 plus.n8 60.6157
R336 plus.n35 plus.n34 60.6157
R337 plus.n72 plus.n71 60.6157
R338 plus.n46 plus.n45 60.6157
R339 plus.n16 plus.n15 47.4702
R340 plus.n28 plus.n27 47.4702
R341 plus.n65 plus.n64 47.4702
R342 plus.n53 plus.n52 47.4702
R343 plus.n16 plus.n5 44.549
R344 plus.n27 plus.n26 44.549
R345 plus.n64 plus.n63 44.549
R346 plus.n53 plus.n42 44.549
R347 plus.n19 plus.n5 28.4823
R348 plus.n26 plus.n25 28.4823
R349 plus.n63 plus.n62 28.4823
R350 plus.n56 plus.n42 28.4823
R351 plus plus.n73 28.4801
R352 plus.n15 plus.n14 25.5611
R353 plus.n29 plus.n28 25.5611
R354 plus.n66 plus.n65 25.5611
R355 plus.n52 plus.n51 25.5611
R356 plus.n8 plus.n7 12.4157
R357 plus.n34 plus.n33 12.4157
R358 plus.n71 plus.n70 12.4157
R359 plus.n45 plus.n44 12.4157
R360 plus.n21 plus.n20 9.49444
R361 plus.n22 plus.n3 9.49444
R362 plus.n59 plus.n40 9.49444
R363 plus.n58 plus.n57 9.49444
R364 plus plus.n36 8.70505
R365 plus.n13 plus.n12 6.57323
R366 plus.n32 plus.n1 6.57323
R367 plus.n69 plus.n38 6.57323
R368 plus.n50 plus.n49 6.57323
R369 plus.n11 plus.n10 0.189894
R370 plus.n11 plus.n6 0.189894
R371 plus.n17 plus.n6 0.189894
R372 plus.n18 plus.n17 0.189894
R373 plus.n18 plus.n4 0.189894
R374 plus.n23 plus.n4 0.189894
R375 plus.n24 plus.n23 0.189894
R376 plus.n24 plus.n2 0.189894
R377 plus.n30 plus.n2 0.189894
R378 plus.n31 plus.n30 0.189894
R379 plus.n31 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n68 plus.n37 0.189894
R383 plus.n68 plus.n67 0.189894
R384 plus.n67 plus.n39 0.189894
R385 plus.n61 plus.n39 0.189894
R386 plus.n61 plus.n60 0.189894
R387 plus.n60 plus.n41 0.189894
R388 plus.n55 plus.n41 0.189894
R389 plus.n55 plus.n54 0.189894
R390 plus.n54 plus.n43 0.189894
R391 plus.n48 plus.n43 0.189894
R392 plus.n48 plus.n47 0.189894
R393 drain_left.n13 drain_left.n11 80.3162
R394 drain_left.n7 drain_left.n5 80.3161
R395 drain_left.n2 drain_left.n0 80.3161
R396 drain_left.n21 drain_left.n20 79.7731
R397 drain_left.n19 drain_left.n18 79.7731
R398 drain_left.n17 drain_left.n16 79.7731
R399 drain_left.n15 drain_left.n14 79.7731
R400 drain_left.n13 drain_left.n12 79.7731
R401 drain_left.n7 drain_left.n6 79.773
R402 drain_left.n9 drain_left.n8 79.773
R403 drain_left.n4 drain_left.n3 79.773
R404 drain_left.n2 drain_left.n1 79.773
R405 drain_left drain_left.n10 25.7084
R406 drain_left.n5 drain_left.t4 6.6005
R407 drain_left.n5 drain_left.t16 6.6005
R408 drain_left.n6 drain_left.t13 6.6005
R409 drain_left.n6 drain_left.t6 6.6005
R410 drain_left.n8 drain_left.t2 6.6005
R411 drain_left.n8 drain_left.t20 6.6005
R412 drain_left.n3 drain_left.t19 6.6005
R413 drain_left.n3 drain_left.t11 6.6005
R414 drain_left.n1 drain_left.t8 6.6005
R415 drain_left.n1 drain_left.t22 6.6005
R416 drain_left.n0 drain_left.t1 6.6005
R417 drain_left.n0 drain_left.t15 6.6005
R418 drain_left.n20 drain_left.t23 6.6005
R419 drain_left.n20 drain_left.t17 6.6005
R420 drain_left.n18 drain_left.t10 6.6005
R421 drain_left.n18 drain_left.t5 6.6005
R422 drain_left.n16 drain_left.t3 6.6005
R423 drain_left.n16 drain_left.t21 6.6005
R424 drain_left.n14 drain_left.t14 6.6005
R425 drain_left.n14 drain_left.t9 6.6005
R426 drain_left.n12 drain_left.t7 6.6005
R427 drain_left.n12 drain_left.t0 6.6005
R428 drain_left.n11 drain_left.t18 6.6005
R429 drain_left.n11 drain_left.t12 6.6005
R430 drain_left drain_left.n21 6.19632
R431 drain_left.n9 drain_left.n7 0.543603
R432 drain_left.n4 drain_left.n2 0.543603
R433 drain_left.n15 drain_left.n13 0.543603
R434 drain_left.n17 drain_left.n15 0.543603
R435 drain_left.n19 drain_left.n17 0.543603
R436 drain_left.n21 drain_left.n19 0.543603
R437 drain_left.n10 drain_left.n9 0.216706
R438 drain_left.n10 drain_left.n4 0.216706
C0 minus source 2.90545f
C1 drain_left plus 2.84846f
C2 plus drain_right 0.393643f
C3 drain_left drain_right 1.26597f
C4 plus minus 4.43426f
C5 drain_left minus 0.177748f
C6 drain_right minus 2.6163f
C7 plus source 2.91945f
C8 drain_left source 13.968699f
C9 drain_right source 13.969299f
C10 drain_right a_n2354_n1488# 5.28769f
C11 drain_left a_n2354_n1488# 5.64379f
C12 source a_n2354_n1488# 3.9098f
C13 minus a_n2354_n1488# 8.553863f
C14 plus a_n2354_n1488# 10.01044f
C15 drain_left.t1 a_n2354_n1488# 0.078246f
C16 drain_left.t15 a_n2354_n1488# 0.078246f
C17 drain_left.n0 a_n2354_n1488# 0.566961f
C18 drain_left.t8 a_n2354_n1488# 0.078246f
C19 drain_left.t22 a_n2354_n1488# 0.078246f
C20 drain_left.n1 a_n2354_n1488# 0.564303f
C21 drain_left.n2 a_n2354_n1488# 0.770086f
C22 drain_left.t19 a_n2354_n1488# 0.078246f
C23 drain_left.t11 a_n2354_n1488# 0.078246f
C24 drain_left.n3 a_n2354_n1488# 0.564303f
C25 drain_left.n4 a_n2354_n1488# 0.348498f
C26 drain_left.t4 a_n2354_n1488# 0.078246f
C27 drain_left.t16 a_n2354_n1488# 0.078246f
C28 drain_left.n5 a_n2354_n1488# 0.566961f
C29 drain_left.t13 a_n2354_n1488# 0.078246f
C30 drain_left.t6 a_n2354_n1488# 0.078246f
C31 drain_left.n6 a_n2354_n1488# 0.564303f
C32 drain_left.n7 a_n2354_n1488# 0.770086f
C33 drain_left.t2 a_n2354_n1488# 0.078246f
C34 drain_left.t20 a_n2354_n1488# 0.078246f
C35 drain_left.n8 a_n2354_n1488# 0.564303f
C36 drain_left.n9 a_n2354_n1488# 0.348498f
C37 drain_left.n10 a_n2354_n1488# 1.16597f
C38 drain_left.t18 a_n2354_n1488# 0.078246f
C39 drain_left.t12 a_n2354_n1488# 0.078246f
C40 drain_left.n11 a_n2354_n1488# 0.566963f
C41 drain_left.t7 a_n2354_n1488# 0.078246f
C42 drain_left.t0 a_n2354_n1488# 0.078246f
C43 drain_left.n12 a_n2354_n1488# 0.564306f
C44 drain_left.n13 a_n2354_n1488# 0.77008f
C45 drain_left.t14 a_n2354_n1488# 0.078246f
C46 drain_left.t9 a_n2354_n1488# 0.078246f
C47 drain_left.n14 a_n2354_n1488# 0.564306f
C48 drain_left.n15 a_n2354_n1488# 0.379722f
C49 drain_left.t3 a_n2354_n1488# 0.078246f
C50 drain_left.t21 a_n2354_n1488# 0.078246f
C51 drain_left.n16 a_n2354_n1488# 0.564306f
C52 drain_left.n17 a_n2354_n1488# 0.379722f
C53 drain_left.t10 a_n2354_n1488# 0.078246f
C54 drain_left.t5 a_n2354_n1488# 0.078246f
C55 drain_left.n18 a_n2354_n1488# 0.564306f
C56 drain_left.n19 a_n2354_n1488# 0.379722f
C57 drain_left.t23 a_n2354_n1488# 0.078246f
C58 drain_left.t17 a_n2354_n1488# 0.078246f
C59 drain_left.n20 a_n2354_n1488# 0.564306f
C60 drain_left.n21 a_n2354_n1488# 0.654448f
C61 plus.n0 a_n2354_n1488# 0.04968f
C62 plus.t0 a_n2354_n1488# 0.129482f
C63 plus.t18 a_n2354_n1488# 0.129482f
C64 plus.n1 a_n2354_n1488# 0.075183f
C65 plus.n2 a_n2354_n1488# 0.04968f
C66 plus.t13 a_n2354_n1488# 0.129482f
C67 plus.t2 a_n2354_n1488# 0.129482f
C68 plus.t20 a_n2354_n1488# 0.129482f
C69 plus.n3 a_n2354_n1488# 0.075183f
C70 plus.n4 a_n2354_n1488# 0.04968f
C71 plus.t14 a_n2354_n1488# 0.129482f
C72 plus.t9 a_n2354_n1488# 0.129482f
C73 plus.n5 a_n2354_n1488# 0.075183f
C74 plus.n6 a_n2354_n1488# 0.04968f
C75 plus.t23 a_n2354_n1488# 0.129482f
C76 plus.t16 a_n2354_n1488# 0.129482f
C77 plus.n7 a_n2354_n1488# 0.019084f
C78 plus.t5 a_n2354_n1488# 0.135785f
C79 plus.t11 a_n2354_n1488# 0.129482f
C80 plus.n8 a_n2354_n1488# 0.075183f
C81 plus.n9 a_n2354_n1488# 0.089868f
C82 plus.n10 a_n2354_n1488# 0.106339f
C83 plus.n11 a_n2354_n1488# 0.04968f
C84 plus.n12 a_n2354_n1488# 0.017859f
C85 plus.n13 a_n2354_n1488# 0.075183f
C86 plus.n14 a_n2354_n1488# 0.020462f
C87 plus.n15 a_n2354_n1488# 0.075183f
C88 plus.n16 a_n2354_n1488# 0.020462f
C89 plus.n17 a_n2354_n1488# 0.04968f
C90 plus.n18 a_n2354_n1488# 0.04968f
C91 plus.n19 a_n2354_n1488# 0.020462f
C92 plus.n20 a_n2354_n1488# 0.075183f
C93 plus.n21 a_n2354_n1488# 0.018472f
C94 plus.n22 a_n2354_n1488# 0.018472f
C95 plus.n23 a_n2354_n1488# 0.04968f
C96 plus.n24 a_n2354_n1488# 0.04968f
C97 plus.n25 a_n2354_n1488# 0.020462f
C98 plus.n26 a_n2354_n1488# 0.075183f
C99 plus.n27 a_n2354_n1488# 0.020462f
C100 plus.n28 a_n2354_n1488# 0.075183f
C101 plus.n29 a_n2354_n1488# 0.020462f
C102 plus.n30 a_n2354_n1488# 0.04968f
C103 plus.n31 a_n2354_n1488# 0.04968f
C104 plus.n32 a_n2354_n1488# 0.017859f
C105 plus.n33 a_n2354_n1488# 0.019084f
C106 plus.n34 a_n2354_n1488# 0.075183f
C107 plus.t6 a_n2354_n1488# 0.135785f
C108 plus.n35 a_n2354_n1488# 0.089801f
C109 plus.n36 a_n2354_n1488# 0.367432f
C110 plus.n37 a_n2354_n1488# 0.04968f
C111 plus.t22 a_n2354_n1488# 0.135785f
C112 plus.t8 a_n2354_n1488# 0.129482f
C113 plus.t15 a_n2354_n1488# 0.129482f
C114 plus.n38 a_n2354_n1488# 0.075183f
C115 plus.n39 a_n2354_n1488# 0.04968f
C116 plus.t1 a_n2354_n1488# 0.129482f
C117 plus.t4 a_n2354_n1488# 0.129482f
C118 plus.t12 a_n2354_n1488# 0.129482f
C119 plus.n40 a_n2354_n1488# 0.075183f
C120 plus.n41 a_n2354_n1488# 0.04968f
C121 plus.t21 a_n2354_n1488# 0.129482f
C122 plus.t3 a_n2354_n1488# 0.129482f
C123 plus.n42 a_n2354_n1488# 0.075183f
C124 plus.n43 a_n2354_n1488# 0.04968f
C125 plus.t10 a_n2354_n1488# 0.129482f
C126 plus.t17 a_n2354_n1488# 0.129482f
C127 plus.n44 a_n2354_n1488# 0.019084f
C128 plus.t19 a_n2354_n1488# 0.129482f
C129 plus.n45 a_n2354_n1488# 0.075183f
C130 plus.t7 a_n2354_n1488# 0.135785f
C131 plus.n46 a_n2354_n1488# 0.089868f
C132 plus.n47 a_n2354_n1488# 0.106339f
C133 plus.n48 a_n2354_n1488# 0.04968f
C134 plus.n49 a_n2354_n1488# 0.017859f
C135 plus.n50 a_n2354_n1488# 0.075183f
C136 plus.n51 a_n2354_n1488# 0.020462f
C137 plus.n52 a_n2354_n1488# 0.075183f
C138 plus.n53 a_n2354_n1488# 0.020462f
C139 plus.n54 a_n2354_n1488# 0.04968f
C140 plus.n55 a_n2354_n1488# 0.04968f
C141 plus.n56 a_n2354_n1488# 0.020462f
C142 plus.n57 a_n2354_n1488# 0.075183f
C143 plus.n58 a_n2354_n1488# 0.018472f
C144 plus.n59 a_n2354_n1488# 0.018472f
C145 plus.n60 a_n2354_n1488# 0.04968f
C146 plus.n61 a_n2354_n1488# 0.04968f
C147 plus.n62 a_n2354_n1488# 0.020462f
C148 plus.n63 a_n2354_n1488# 0.075183f
C149 plus.n64 a_n2354_n1488# 0.020462f
C150 plus.n65 a_n2354_n1488# 0.075183f
C151 plus.n66 a_n2354_n1488# 0.020462f
C152 plus.n67 a_n2354_n1488# 0.04968f
C153 plus.n68 a_n2354_n1488# 0.04968f
C154 plus.n69 a_n2354_n1488# 0.017859f
C155 plus.n70 a_n2354_n1488# 0.019084f
C156 plus.n71 a_n2354_n1488# 0.075183f
C157 plus.n72 a_n2354_n1488# 0.089801f
C158 plus.n73 a_n2354_n1488# 1.29417f
C159 source.t23 a_n2354_n1488# 0.662836f
C160 source.n0 a_n2354_n1488# 0.904331f
C161 source.t3 a_n2354_n1488# 0.079823f
C162 source.t9 a_n2354_n1488# 0.079823f
C163 source.n1 a_n2354_n1488# 0.506124f
C164 source.n2 a_n2354_n1488# 0.411164f
C165 source.t10 a_n2354_n1488# 0.079823f
C166 source.t1 a_n2354_n1488# 0.079823f
C167 source.n3 a_n2354_n1488# 0.506124f
C168 source.n4 a_n2354_n1488# 0.411164f
C169 source.t8 a_n2354_n1488# 0.079823f
C170 source.t17 a_n2354_n1488# 0.079823f
C171 source.n5 a_n2354_n1488# 0.506124f
C172 source.n6 a_n2354_n1488# 0.411164f
C173 source.t7 a_n2354_n1488# 0.079823f
C174 source.t20 a_n2354_n1488# 0.079823f
C175 source.n7 a_n2354_n1488# 0.506124f
C176 source.n8 a_n2354_n1488# 0.411164f
C177 source.t16 a_n2354_n1488# 0.079823f
C178 source.t15 a_n2354_n1488# 0.079823f
C179 source.n9 a_n2354_n1488# 0.506124f
C180 source.n10 a_n2354_n1488# 0.411164f
C181 source.t19 a_n2354_n1488# 0.662836f
C182 source.n11 a_n2354_n1488# 0.4642f
C183 source.t33 a_n2354_n1488# 0.662836f
C184 source.n12 a_n2354_n1488# 0.4642f
C185 source.t43 a_n2354_n1488# 0.079823f
C186 source.t27 a_n2354_n1488# 0.079823f
C187 source.n13 a_n2354_n1488# 0.506124f
C188 source.n14 a_n2354_n1488# 0.411164f
C189 source.t29 a_n2354_n1488# 0.079823f
C190 source.t34 a_n2354_n1488# 0.079823f
C191 source.n15 a_n2354_n1488# 0.506124f
C192 source.n16 a_n2354_n1488# 0.411164f
C193 source.t39 a_n2354_n1488# 0.079823f
C194 source.t45 a_n2354_n1488# 0.079823f
C195 source.n17 a_n2354_n1488# 0.506124f
C196 source.n18 a_n2354_n1488# 0.411164f
C197 source.t42 a_n2354_n1488# 0.079823f
C198 source.t26 a_n2354_n1488# 0.079823f
C199 source.n19 a_n2354_n1488# 0.506124f
C200 source.n20 a_n2354_n1488# 0.411164f
C201 source.t28 a_n2354_n1488# 0.079823f
C202 source.t38 a_n2354_n1488# 0.079823f
C203 source.n21 a_n2354_n1488# 0.506124f
C204 source.n22 a_n2354_n1488# 0.411164f
C205 source.t41 a_n2354_n1488# 0.662836f
C206 source.n23 a_n2354_n1488# 1.2553f
C207 source.t2 a_n2354_n1488# 0.662833f
C208 source.n24 a_n2354_n1488# 1.25531f
C209 source.t0 a_n2354_n1488# 0.079823f
C210 source.t11 a_n2354_n1488# 0.079823f
C211 source.n25 a_n2354_n1488# 0.50612f
C212 source.n26 a_n2354_n1488# 0.411167f
C213 source.t4 a_n2354_n1488# 0.079823f
C214 source.t6 a_n2354_n1488# 0.079823f
C215 source.n27 a_n2354_n1488# 0.50612f
C216 source.n28 a_n2354_n1488# 0.411167f
C217 source.t21 a_n2354_n1488# 0.079823f
C218 source.t22 a_n2354_n1488# 0.079823f
C219 source.n29 a_n2354_n1488# 0.50612f
C220 source.n30 a_n2354_n1488# 0.411167f
C221 source.t14 a_n2354_n1488# 0.079823f
C222 source.t12 a_n2354_n1488# 0.079823f
C223 source.n31 a_n2354_n1488# 0.50612f
C224 source.n32 a_n2354_n1488# 0.411167f
C225 source.t5 a_n2354_n1488# 0.079823f
C226 source.t18 a_n2354_n1488# 0.079823f
C227 source.n33 a_n2354_n1488# 0.50612f
C228 source.n34 a_n2354_n1488# 0.411167f
C229 source.t13 a_n2354_n1488# 0.662833f
C230 source.n35 a_n2354_n1488# 0.464204f
C231 source.t36 a_n2354_n1488# 0.662833f
C232 source.n36 a_n2354_n1488# 0.464204f
C233 source.t46 a_n2354_n1488# 0.079823f
C234 source.t24 a_n2354_n1488# 0.079823f
C235 source.n37 a_n2354_n1488# 0.50612f
C236 source.n38 a_n2354_n1488# 0.411167f
C237 source.t35 a_n2354_n1488# 0.079823f
C238 source.t40 a_n2354_n1488# 0.079823f
C239 source.n39 a_n2354_n1488# 0.50612f
C240 source.n40 a_n2354_n1488# 0.411167f
C241 source.t44 a_n2354_n1488# 0.079823f
C242 source.t31 a_n2354_n1488# 0.079823f
C243 source.n41 a_n2354_n1488# 0.50612f
C244 source.n42 a_n2354_n1488# 0.411167f
C245 source.t32 a_n2354_n1488# 0.079823f
C246 source.t47 a_n2354_n1488# 0.079823f
C247 source.n43 a_n2354_n1488# 0.50612f
C248 source.n44 a_n2354_n1488# 0.411167f
C249 source.t25 a_n2354_n1488# 0.079823f
C250 source.t30 a_n2354_n1488# 0.079823f
C251 source.n45 a_n2354_n1488# 0.50612f
C252 source.n46 a_n2354_n1488# 0.411167f
C253 source.t37 a_n2354_n1488# 0.662833f
C254 source.n47 a_n2354_n1488# 0.654275f
C255 source.n48 a_n2354_n1488# 0.975953f
C256 drain_right.t9 a_n2354_n1488# 0.077913f
C257 drain_right.t2 a_n2354_n1488# 0.077913f
C258 drain_right.n0 a_n2354_n1488# 0.56455f
C259 drain_right.t18 a_n2354_n1488# 0.077913f
C260 drain_right.t10 a_n2354_n1488# 0.077913f
C261 drain_right.n1 a_n2354_n1488# 0.561904f
C262 drain_right.n2 a_n2354_n1488# 0.766811f
C263 drain_right.t5 a_n2354_n1488# 0.077913f
C264 drain_right.t1 a_n2354_n1488# 0.077913f
C265 drain_right.n3 a_n2354_n1488# 0.561904f
C266 drain_right.n4 a_n2354_n1488# 0.347016f
C267 drain_right.t15 a_n2354_n1488# 0.077913f
C268 drain_right.t8 a_n2354_n1488# 0.077913f
C269 drain_right.n5 a_n2354_n1488# 0.56455f
C270 drain_right.t22 a_n2354_n1488# 0.077913f
C271 drain_right.t21 a_n2354_n1488# 0.077913f
C272 drain_right.n6 a_n2354_n1488# 0.561904f
C273 drain_right.n7 a_n2354_n1488# 0.766811f
C274 drain_right.t14 a_n2354_n1488# 0.077913f
C275 drain_right.t13 a_n2354_n1488# 0.077913f
C276 drain_right.n8 a_n2354_n1488# 0.561904f
C277 drain_right.n9 a_n2354_n1488# 0.347016f
C278 drain_right.n10 a_n2354_n1488# 1.0963f
C279 drain_right.t20 a_n2354_n1488# 0.077913f
C280 drain_right.t12 a_n2354_n1488# 0.077913f
C281 drain_right.n11 a_n2354_n1488# 0.564553f
C282 drain_right.t11 a_n2354_n1488# 0.077913f
C283 drain_right.t23 a_n2354_n1488# 0.077913f
C284 drain_right.n12 a_n2354_n1488# 0.561906f
C285 drain_right.n13 a_n2354_n1488# 0.766806f
C286 drain_right.t0 a_n2354_n1488# 0.077913f
C287 drain_right.t16 a_n2354_n1488# 0.077913f
C288 drain_right.n14 a_n2354_n1488# 0.561906f
C289 drain_right.n15 a_n2354_n1488# 0.378107f
C290 drain_right.t17 a_n2354_n1488# 0.077913f
C291 drain_right.t6 a_n2354_n1488# 0.077913f
C292 drain_right.n16 a_n2354_n1488# 0.561906f
C293 drain_right.n17 a_n2354_n1488# 0.378107f
C294 drain_right.t7 a_n2354_n1488# 0.077913f
C295 drain_right.t3 a_n2354_n1488# 0.077913f
C296 drain_right.n18 a_n2354_n1488# 0.561906f
C297 drain_right.n19 a_n2354_n1488# 0.378107f
C298 drain_right.t4 a_n2354_n1488# 0.077913f
C299 drain_right.t19 a_n2354_n1488# 0.077913f
C300 drain_right.n20 a_n2354_n1488# 0.561906f
C301 drain_right.n21 a_n2354_n1488# 0.651665f
C302 minus.n0 a_n2354_n1488# 0.048217f
C303 minus.t6 a_n2354_n1488# 0.131786f
C304 minus.t19 a_n2354_n1488# 0.125668f
C305 minus.t9 a_n2354_n1488# 0.125668f
C306 minus.n1 a_n2354_n1488# 0.072968f
C307 minus.n2 a_n2354_n1488# 0.048217f
C308 minus.t5 a_n2354_n1488# 0.125668f
C309 minus.t21 a_n2354_n1488# 0.125668f
C310 minus.t8 a_n2354_n1488# 0.125668f
C311 minus.n3 a_n2354_n1488# 0.072968f
C312 minus.n4 a_n2354_n1488# 0.048217f
C313 minus.t2 a_n2354_n1488# 0.125668f
C314 minus.t18 a_n2354_n1488# 0.125668f
C315 minus.n5 a_n2354_n1488# 0.072968f
C316 minus.n6 a_n2354_n1488# 0.048217f
C317 minus.t13 a_n2354_n1488# 0.125668f
C318 minus.t4 a_n2354_n1488# 0.125668f
C319 minus.n7 a_n2354_n1488# 0.018522f
C320 minus.t20 a_n2354_n1488# 0.125668f
C321 minus.n8 a_n2354_n1488# 0.072968f
C322 minus.t14 a_n2354_n1488# 0.131786f
C323 minus.n9 a_n2354_n1488# 0.087221f
C324 minus.n10 a_n2354_n1488# 0.103207f
C325 minus.n11 a_n2354_n1488# 0.048217f
C326 minus.n12 a_n2354_n1488# 0.017333f
C327 minus.n13 a_n2354_n1488# 0.072968f
C328 minus.n14 a_n2354_n1488# 0.01986f
C329 minus.n15 a_n2354_n1488# 0.072968f
C330 minus.n16 a_n2354_n1488# 0.01986f
C331 minus.n17 a_n2354_n1488# 0.048217f
C332 minus.n18 a_n2354_n1488# 0.048217f
C333 minus.n19 a_n2354_n1488# 0.01986f
C334 minus.n20 a_n2354_n1488# 0.072968f
C335 minus.n21 a_n2354_n1488# 0.017927f
C336 minus.n22 a_n2354_n1488# 0.017927f
C337 minus.n23 a_n2354_n1488# 0.048217f
C338 minus.n24 a_n2354_n1488# 0.048217f
C339 minus.n25 a_n2354_n1488# 0.01986f
C340 minus.n26 a_n2354_n1488# 0.072968f
C341 minus.n27 a_n2354_n1488# 0.01986f
C342 minus.n28 a_n2354_n1488# 0.072968f
C343 minus.n29 a_n2354_n1488# 0.01986f
C344 minus.n30 a_n2354_n1488# 0.048217f
C345 minus.n31 a_n2354_n1488# 0.048217f
C346 minus.n32 a_n2354_n1488# 0.017333f
C347 minus.n33 a_n2354_n1488# 0.018522f
C348 minus.n34 a_n2354_n1488# 0.072968f
C349 minus.n35 a_n2354_n1488# 0.087156f
C350 minus.n36 a_n2354_n1488# 1.33831f
C351 minus.n37 a_n2354_n1488# 0.048217f
C352 minus.t17 a_n2354_n1488# 0.125668f
C353 minus.t22 a_n2354_n1488# 0.125668f
C354 minus.n38 a_n2354_n1488# 0.072968f
C355 minus.n39 a_n2354_n1488# 0.048217f
C356 minus.t0 a_n2354_n1488# 0.125668f
C357 minus.t15 a_n2354_n1488# 0.125668f
C358 minus.t16 a_n2354_n1488# 0.125668f
C359 minus.n40 a_n2354_n1488# 0.072968f
C360 minus.n41 a_n2354_n1488# 0.048217f
C361 minus.t3 a_n2354_n1488# 0.125668f
C362 minus.t7 a_n2354_n1488# 0.125668f
C363 minus.n42 a_n2354_n1488# 0.072968f
C364 minus.n43 a_n2354_n1488# 0.048217f
C365 minus.t12 a_n2354_n1488# 0.125668f
C366 minus.t23 a_n2354_n1488# 0.125668f
C367 minus.n44 a_n2354_n1488# 0.018522f
C368 minus.t11 a_n2354_n1488# 0.131786f
C369 minus.t1 a_n2354_n1488# 0.125668f
C370 minus.n45 a_n2354_n1488# 0.072968f
C371 minus.n46 a_n2354_n1488# 0.087221f
C372 minus.n47 a_n2354_n1488# 0.103207f
C373 minus.n48 a_n2354_n1488# 0.048217f
C374 minus.n49 a_n2354_n1488# 0.017333f
C375 minus.n50 a_n2354_n1488# 0.072968f
C376 minus.n51 a_n2354_n1488# 0.01986f
C377 minus.n52 a_n2354_n1488# 0.072968f
C378 minus.n53 a_n2354_n1488# 0.01986f
C379 minus.n54 a_n2354_n1488# 0.048217f
C380 minus.n55 a_n2354_n1488# 0.048217f
C381 minus.n56 a_n2354_n1488# 0.01986f
C382 minus.n57 a_n2354_n1488# 0.072968f
C383 minus.n58 a_n2354_n1488# 0.017927f
C384 minus.n59 a_n2354_n1488# 0.017927f
C385 minus.n60 a_n2354_n1488# 0.048217f
C386 minus.n61 a_n2354_n1488# 0.048217f
C387 minus.n62 a_n2354_n1488# 0.01986f
C388 minus.n63 a_n2354_n1488# 0.072968f
C389 minus.n64 a_n2354_n1488# 0.01986f
C390 minus.n65 a_n2354_n1488# 0.072968f
C391 minus.n66 a_n2354_n1488# 0.01986f
C392 minus.n67 a_n2354_n1488# 0.048217f
C393 minus.n68 a_n2354_n1488# 0.048217f
C394 minus.n69 a_n2354_n1488# 0.017333f
C395 minus.n70 a_n2354_n1488# 0.018522f
C396 minus.n71 a_n2354_n1488# 0.072968f
C397 minus.t10 a_n2354_n1488# 0.131786f
C398 minus.n72 a_n2354_n1488# 0.087156f
C399 minus.n73 a_n2354_n1488# 0.31184f
C400 minus.n74 a_n2354_n1488# 1.64893f
.ends

