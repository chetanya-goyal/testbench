* NGSPICE file created from diffpair429.ext - technology: sky130A

.subckt diffpair429 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t31 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 drain_left.t22 plus.t1 source.t39 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 drain_left.t21 plus.t2 source.t24 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X3 drain_left.t20 plus.t3 source.t47 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X4 source.t11 minus.t0 drain_right.t23 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X5 drain_left.t19 plus.t4 source.t36 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 source.t15 minus.t1 drain_right.t22 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X7 drain_right.t21 minus.t2 source.t0 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X8 drain_right.t20 minus.t3 source.t1 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X9 drain_right.t19 minus.t4 source.t7 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 drain_left.t18 plus.t5 source.t46 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X11 source.t45 plus.t6 drain_left.t17 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X12 source.t2 minus.t5 drain_right.t18 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X13 source.t33 plus.t7 drain_left.t16 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X14 source.t21 minus.t6 drain_right.t17 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X15 source.t12 minus.t7 drain_right.t16 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X16 drain_left.t15 plus.t8 source.t32 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X17 a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X18 source.t17 minus.t8 drain_right.t15 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X19 source.t40 plus.t9 drain_left.t14 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X20 source.t27 plus.t10 drain_left.t13 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X21 source.t29 plus.t11 drain_left.t12 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X22 source.t42 plus.t12 drain_left.t11 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X23 a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X24 source.t9 minus.t9 drain_right.t14 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X25 drain_left.t10 plus.t13 source.t41 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X26 source.t43 plus.t14 drain_left.t9 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X27 drain_right.t13 minus.t10 source.t20 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X28 source.t25 plus.t15 drain_left.t8 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X29 source.t37 plus.t16 drain_left.t7 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X30 drain_right.t12 minus.t11 source.t23 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X31 drain_right.t11 minus.t12 source.t16 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X32 source.t18 minus.t13 drain_right.t10 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X33 a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X34 drain_right.t9 minus.t14 source.t8 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X35 drain_left.t6 plus.t17 source.t38 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X36 drain_right.t8 minus.t15 source.t14 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X37 source.t30 plus.t18 drain_left.t5 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X38 drain_left.t4 plus.t19 source.t28 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X39 source.t19 minus.t16 drain_right.t7 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X40 source.t22 minus.t17 drain_right.t6 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X41 source.t4 minus.t18 drain_right.t5 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X42 source.t26 plus.t20 drain_left.t3 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X43 drain_right.t4 minus.t19 source.t10 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X44 drain_right.t3 minus.t20 source.t13 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X45 drain_left.t2 plus.t21 source.t44 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X46 drain_right.t2 minus.t21 source.t5 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X47 drain_right.t1 minus.t22 source.t3 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X48 drain_left.t1 plus.t22 source.t35 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X49 source.t6 minus.t23 drain_right.t0 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X50 source.t34 plus.t23 drain_left.t0 a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X51 a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# a_n2224_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
R0 plus.n6 plus.t6 1309.87
R1 plus.n33 plus.t2 1309.87
R2 plus.n42 plus.t21 1309.87
R3 plus.n68 plus.t9 1309.87
R4 plus.n7 plus.t1 1282.12
R5 plus.n8 plus.t12 1282.12
R6 plus.n14 plus.t0 1282.12
R7 plus.n16 plus.t11 1282.12
R8 plus.n3 plus.t22 1282.12
R9 plus.n21 plus.t10 1282.12
R10 plus.n23 plus.t4 1282.12
R11 plus.n24 plus.t16 1282.12
R12 plus.n30 plus.t3 1282.12
R13 plus.n32 plus.t14 1282.12
R14 plus.n44 plus.t18 1282.12
R15 plus.n43 plus.t8 1282.12
R16 plus.n50 plus.t23 1282.12
R17 plus.n52 plus.t5 1282.12
R18 plus.n39 plus.t20 1282.12
R19 plus.n57 plus.t17 1282.12
R20 plus.n59 plus.t7 1282.12
R21 plus.n38 plus.t19 1282.12
R22 plus.n65 plus.t15 1282.12
R23 plus.n67 plus.t13 1282.12
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus plus.n69 31.3589
R75 plus.n17 plus.n3 30.6732
R76 plus.n22 plus.n21 30.6732
R77 plus.n58 plus.n57 30.6732
R78 plus.n53 plus.n39 30.6732
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 12.0763
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n562 source.n502 289.615
R119 source.n486 source.n426 289.615
R120 source.n420 source.n360 289.615
R121 source.n344 source.n284 289.615
R122 source.n60 source.n0 289.615
R123 source.n136 source.n76 289.615
R124 source.n202 source.n142 289.615
R125 source.n278 source.n218 289.615
R126 source.n522 source.n521 185
R127 source.n527 source.n526 185
R128 source.n529 source.n528 185
R129 source.n518 source.n517 185
R130 source.n535 source.n534 185
R131 source.n537 source.n536 185
R132 source.n514 source.n513 185
R133 source.n544 source.n543 185
R134 source.n545 source.n512 185
R135 source.n547 source.n546 185
R136 source.n510 source.n509 185
R137 source.n553 source.n552 185
R138 source.n555 source.n554 185
R139 source.n506 source.n505 185
R140 source.n561 source.n560 185
R141 source.n563 source.n562 185
R142 source.n446 source.n445 185
R143 source.n451 source.n450 185
R144 source.n453 source.n452 185
R145 source.n442 source.n441 185
R146 source.n459 source.n458 185
R147 source.n461 source.n460 185
R148 source.n438 source.n437 185
R149 source.n468 source.n467 185
R150 source.n469 source.n436 185
R151 source.n471 source.n470 185
R152 source.n434 source.n433 185
R153 source.n477 source.n476 185
R154 source.n479 source.n478 185
R155 source.n430 source.n429 185
R156 source.n485 source.n484 185
R157 source.n487 source.n486 185
R158 source.n380 source.n379 185
R159 source.n385 source.n384 185
R160 source.n387 source.n386 185
R161 source.n376 source.n375 185
R162 source.n393 source.n392 185
R163 source.n395 source.n394 185
R164 source.n372 source.n371 185
R165 source.n402 source.n401 185
R166 source.n403 source.n370 185
R167 source.n405 source.n404 185
R168 source.n368 source.n367 185
R169 source.n411 source.n410 185
R170 source.n413 source.n412 185
R171 source.n364 source.n363 185
R172 source.n419 source.n418 185
R173 source.n421 source.n420 185
R174 source.n304 source.n303 185
R175 source.n309 source.n308 185
R176 source.n311 source.n310 185
R177 source.n300 source.n299 185
R178 source.n317 source.n316 185
R179 source.n319 source.n318 185
R180 source.n296 source.n295 185
R181 source.n326 source.n325 185
R182 source.n327 source.n294 185
R183 source.n329 source.n328 185
R184 source.n292 source.n291 185
R185 source.n335 source.n334 185
R186 source.n337 source.n336 185
R187 source.n288 source.n287 185
R188 source.n343 source.n342 185
R189 source.n345 source.n344 185
R190 source.n61 source.n60 185
R191 source.n59 source.n58 185
R192 source.n4 source.n3 185
R193 source.n53 source.n52 185
R194 source.n51 source.n50 185
R195 source.n8 source.n7 185
R196 source.n45 source.n44 185
R197 source.n43 source.n10 185
R198 source.n42 source.n41 185
R199 source.n13 source.n11 185
R200 source.n36 source.n35 185
R201 source.n34 source.n33 185
R202 source.n17 source.n16 185
R203 source.n28 source.n27 185
R204 source.n26 source.n25 185
R205 source.n21 source.n20 185
R206 source.n137 source.n136 185
R207 source.n135 source.n134 185
R208 source.n80 source.n79 185
R209 source.n129 source.n128 185
R210 source.n127 source.n126 185
R211 source.n84 source.n83 185
R212 source.n121 source.n120 185
R213 source.n119 source.n86 185
R214 source.n118 source.n117 185
R215 source.n89 source.n87 185
R216 source.n112 source.n111 185
R217 source.n110 source.n109 185
R218 source.n93 source.n92 185
R219 source.n104 source.n103 185
R220 source.n102 source.n101 185
R221 source.n97 source.n96 185
R222 source.n203 source.n202 185
R223 source.n201 source.n200 185
R224 source.n146 source.n145 185
R225 source.n195 source.n194 185
R226 source.n193 source.n192 185
R227 source.n150 source.n149 185
R228 source.n187 source.n186 185
R229 source.n185 source.n152 185
R230 source.n184 source.n183 185
R231 source.n155 source.n153 185
R232 source.n178 source.n177 185
R233 source.n176 source.n175 185
R234 source.n159 source.n158 185
R235 source.n170 source.n169 185
R236 source.n168 source.n167 185
R237 source.n163 source.n162 185
R238 source.n279 source.n278 185
R239 source.n277 source.n276 185
R240 source.n222 source.n221 185
R241 source.n271 source.n270 185
R242 source.n269 source.n268 185
R243 source.n226 source.n225 185
R244 source.n263 source.n262 185
R245 source.n261 source.n228 185
R246 source.n260 source.n259 185
R247 source.n231 source.n229 185
R248 source.n254 source.n253 185
R249 source.n252 source.n251 185
R250 source.n235 source.n234 185
R251 source.n246 source.n245 185
R252 source.n244 source.n243 185
R253 source.n239 source.n238 185
R254 source.n523 source.t8 149.524
R255 source.n447 source.t6 149.524
R256 source.n381 source.t44 149.524
R257 source.n305 source.t40 149.524
R258 source.n22 source.t24 149.524
R259 source.n98 source.t45 149.524
R260 source.n164 source.t23 149.524
R261 source.n240 source.t18 149.524
R262 source.n527 source.n521 104.615
R263 source.n528 source.n527 104.615
R264 source.n528 source.n517 104.615
R265 source.n535 source.n517 104.615
R266 source.n536 source.n535 104.615
R267 source.n536 source.n513 104.615
R268 source.n544 source.n513 104.615
R269 source.n545 source.n544 104.615
R270 source.n546 source.n545 104.615
R271 source.n546 source.n509 104.615
R272 source.n553 source.n509 104.615
R273 source.n554 source.n553 104.615
R274 source.n554 source.n505 104.615
R275 source.n561 source.n505 104.615
R276 source.n562 source.n561 104.615
R277 source.n451 source.n445 104.615
R278 source.n452 source.n451 104.615
R279 source.n452 source.n441 104.615
R280 source.n459 source.n441 104.615
R281 source.n460 source.n459 104.615
R282 source.n460 source.n437 104.615
R283 source.n468 source.n437 104.615
R284 source.n469 source.n468 104.615
R285 source.n470 source.n469 104.615
R286 source.n470 source.n433 104.615
R287 source.n477 source.n433 104.615
R288 source.n478 source.n477 104.615
R289 source.n478 source.n429 104.615
R290 source.n485 source.n429 104.615
R291 source.n486 source.n485 104.615
R292 source.n385 source.n379 104.615
R293 source.n386 source.n385 104.615
R294 source.n386 source.n375 104.615
R295 source.n393 source.n375 104.615
R296 source.n394 source.n393 104.615
R297 source.n394 source.n371 104.615
R298 source.n402 source.n371 104.615
R299 source.n403 source.n402 104.615
R300 source.n404 source.n403 104.615
R301 source.n404 source.n367 104.615
R302 source.n411 source.n367 104.615
R303 source.n412 source.n411 104.615
R304 source.n412 source.n363 104.615
R305 source.n419 source.n363 104.615
R306 source.n420 source.n419 104.615
R307 source.n309 source.n303 104.615
R308 source.n310 source.n309 104.615
R309 source.n310 source.n299 104.615
R310 source.n317 source.n299 104.615
R311 source.n318 source.n317 104.615
R312 source.n318 source.n295 104.615
R313 source.n326 source.n295 104.615
R314 source.n327 source.n326 104.615
R315 source.n328 source.n327 104.615
R316 source.n328 source.n291 104.615
R317 source.n335 source.n291 104.615
R318 source.n336 source.n335 104.615
R319 source.n336 source.n287 104.615
R320 source.n343 source.n287 104.615
R321 source.n344 source.n343 104.615
R322 source.n60 source.n59 104.615
R323 source.n59 source.n3 104.615
R324 source.n52 source.n3 104.615
R325 source.n52 source.n51 104.615
R326 source.n51 source.n7 104.615
R327 source.n44 source.n7 104.615
R328 source.n44 source.n43 104.615
R329 source.n43 source.n42 104.615
R330 source.n42 source.n11 104.615
R331 source.n35 source.n11 104.615
R332 source.n35 source.n34 104.615
R333 source.n34 source.n16 104.615
R334 source.n27 source.n16 104.615
R335 source.n27 source.n26 104.615
R336 source.n26 source.n20 104.615
R337 source.n136 source.n135 104.615
R338 source.n135 source.n79 104.615
R339 source.n128 source.n79 104.615
R340 source.n128 source.n127 104.615
R341 source.n127 source.n83 104.615
R342 source.n120 source.n83 104.615
R343 source.n120 source.n119 104.615
R344 source.n119 source.n118 104.615
R345 source.n118 source.n87 104.615
R346 source.n111 source.n87 104.615
R347 source.n111 source.n110 104.615
R348 source.n110 source.n92 104.615
R349 source.n103 source.n92 104.615
R350 source.n103 source.n102 104.615
R351 source.n102 source.n96 104.615
R352 source.n202 source.n201 104.615
R353 source.n201 source.n145 104.615
R354 source.n194 source.n145 104.615
R355 source.n194 source.n193 104.615
R356 source.n193 source.n149 104.615
R357 source.n186 source.n149 104.615
R358 source.n186 source.n185 104.615
R359 source.n185 source.n184 104.615
R360 source.n184 source.n153 104.615
R361 source.n177 source.n153 104.615
R362 source.n177 source.n176 104.615
R363 source.n176 source.n158 104.615
R364 source.n169 source.n158 104.615
R365 source.n169 source.n168 104.615
R366 source.n168 source.n162 104.615
R367 source.n278 source.n277 104.615
R368 source.n277 source.n221 104.615
R369 source.n270 source.n221 104.615
R370 source.n270 source.n269 104.615
R371 source.n269 source.n225 104.615
R372 source.n262 source.n225 104.615
R373 source.n262 source.n261 104.615
R374 source.n261 source.n260 104.615
R375 source.n260 source.n229 104.615
R376 source.n253 source.n229 104.615
R377 source.n253 source.n252 104.615
R378 source.n252 source.n234 104.615
R379 source.n245 source.n234 104.615
R380 source.n245 source.n244 104.615
R381 source.n244 source.n238 104.615
R382 source.t8 source.n521 52.3082
R383 source.t6 source.n445 52.3082
R384 source.t44 source.n379 52.3082
R385 source.t40 source.n303 52.3082
R386 source.t24 source.n20 52.3082
R387 source.t45 source.n96 52.3082
R388 source.t23 source.n162 52.3082
R389 source.t18 source.n238 52.3082
R390 source.n67 source.n66 42.8739
R391 source.n69 source.n68 42.8739
R392 source.n71 source.n70 42.8739
R393 source.n73 source.n72 42.8739
R394 source.n75 source.n74 42.8739
R395 source.n209 source.n208 42.8739
R396 source.n211 source.n210 42.8739
R397 source.n213 source.n212 42.8739
R398 source.n215 source.n214 42.8739
R399 source.n217 source.n216 42.8739
R400 source.n501 source.n500 42.8737
R401 source.n499 source.n498 42.8737
R402 source.n497 source.n496 42.8737
R403 source.n495 source.n494 42.8737
R404 source.n493 source.n492 42.8737
R405 source.n359 source.n358 42.8737
R406 source.n357 source.n356 42.8737
R407 source.n355 source.n354 42.8737
R408 source.n353 source.n352 42.8737
R409 source.n351 source.n350 42.8737
R410 source.n567 source.n566 29.8581
R411 source.n491 source.n490 29.8581
R412 source.n425 source.n424 29.8581
R413 source.n349 source.n348 29.8581
R414 source.n65 source.n64 29.8581
R415 source.n141 source.n140 29.8581
R416 source.n207 source.n206 29.8581
R417 source.n283 source.n282 29.8581
R418 source.n349 source.n283 21.7877
R419 source.n568 source.n65 16.2748
R420 source.n547 source.n512 13.1884
R421 source.n471 source.n436 13.1884
R422 source.n405 source.n370 13.1884
R423 source.n329 source.n294 13.1884
R424 source.n45 source.n10 13.1884
R425 source.n121 source.n86 13.1884
R426 source.n187 source.n152 13.1884
R427 source.n263 source.n228 13.1884
R428 source.n543 source.n542 12.8005
R429 source.n548 source.n510 12.8005
R430 source.n467 source.n466 12.8005
R431 source.n472 source.n434 12.8005
R432 source.n401 source.n400 12.8005
R433 source.n406 source.n368 12.8005
R434 source.n325 source.n324 12.8005
R435 source.n330 source.n292 12.8005
R436 source.n46 source.n8 12.8005
R437 source.n41 source.n12 12.8005
R438 source.n122 source.n84 12.8005
R439 source.n117 source.n88 12.8005
R440 source.n188 source.n150 12.8005
R441 source.n183 source.n154 12.8005
R442 source.n264 source.n226 12.8005
R443 source.n259 source.n230 12.8005
R444 source.n541 source.n514 12.0247
R445 source.n552 source.n551 12.0247
R446 source.n465 source.n438 12.0247
R447 source.n476 source.n475 12.0247
R448 source.n399 source.n372 12.0247
R449 source.n410 source.n409 12.0247
R450 source.n323 source.n296 12.0247
R451 source.n334 source.n333 12.0247
R452 source.n50 source.n49 12.0247
R453 source.n40 source.n13 12.0247
R454 source.n126 source.n125 12.0247
R455 source.n116 source.n89 12.0247
R456 source.n192 source.n191 12.0247
R457 source.n182 source.n155 12.0247
R458 source.n268 source.n267 12.0247
R459 source.n258 source.n231 12.0247
R460 source.n538 source.n537 11.249
R461 source.n555 source.n508 11.249
R462 source.n462 source.n461 11.249
R463 source.n479 source.n432 11.249
R464 source.n396 source.n395 11.249
R465 source.n413 source.n366 11.249
R466 source.n320 source.n319 11.249
R467 source.n337 source.n290 11.249
R468 source.n53 source.n6 11.249
R469 source.n37 source.n36 11.249
R470 source.n129 source.n82 11.249
R471 source.n113 source.n112 11.249
R472 source.n195 source.n148 11.249
R473 source.n179 source.n178 11.249
R474 source.n271 source.n224 11.249
R475 source.n255 source.n254 11.249
R476 source.n534 source.n516 10.4732
R477 source.n556 source.n506 10.4732
R478 source.n458 source.n440 10.4732
R479 source.n480 source.n430 10.4732
R480 source.n392 source.n374 10.4732
R481 source.n414 source.n364 10.4732
R482 source.n316 source.n298 10.4732
R483 source.n338 source.n288 10.4732
R484 source.n54 source.n4 10.4732
R485 source.n33 source.n15 10.4732
R486 source.n130 source.n80 10.4732
R487 source.n109 source.n91 10.4732
R488 source.n196 source.n146 10.4732
R489 source.n175 source.n157 10.4732
R490 source.n272 source.n222 10.4732
R491 source.n251 source.n233 10.4732
R492 source.n523 source.n522 10.2747
R493 source.n447 source.n446 10.2747
R494 source.n381 source.n380 10.2747
R495 source.n305 source.n304 10.2747
R496 source.n22 source.n21 10.2747
R497 source.n98 source.n97 10.2747
R498 source.n164 source.n163 10.2747
R499 source.n240 source.n239 10.2747
R500 source.n533 source.n518 9.69747
R501 source.n560 source.n559 9.69747
R502 source.n457 source.n442 9.69747
R503 source.n484 source.n483 9.69747
R504 source.n391 source.n376 9.69747
R505 source.n418 source.n417 9.69747
R506 source.n315 source.n300 9.69747
R507 source.n342 source.n341 9.69747
R508 source.n58 source.n57 9.69747
R509 source.n32 source.n17 9.69747
R510 source.n134 source.n133 9.69747
R511 source.n108 source.n93 9.69747
R512 source.n200 source.n199 9.69747
R513 source.n174 source.n159 9.69747
R514 source.n276 source.n275 9.69747
R515 source.n250 source.n235 9.69747
R516 source.n566 source.n565 9.45567
R517 source.n490 source.n489 9.45567
R518 source.n424 source.n423 9.45567
R519 source.n348 source.n347 9.45567
R520 source.n64 source.n63 9.45567
R521 source.n140 source.n139 9.45567
R522 source.n206 source.n205 9.45567
R523 source.n282 source.n281 9.45567
R524 source.n565 source.n564 9.3005
R525 source.n504 source.n503 9.3005
R526 source.n559 source.n558 9.3005
R527 source.n557 source.n556 9.3005
R528 source.n508 source.n507 9.3005
R529 source.n551 source.n550 9.3005
R530 source.n549 source.n548 9.3005
R531 source.n525 source.n524 9.3005
R532 source.n520 source.n519 9.3005
R533 source.n531 source.n530 9.3005
R534 source.n533 source.n532 9.3005
R535 source.n516 source.n515 9.3005
R536 source.n539 source.n538 9.3005
R537 source.n541 source.n540 9.3005
R538 source.n542 source.n511 9.3005
R539 source.n489 source.n488 9.3005
R540 source.n428 source.n427 9.3005
R541 source.n483 source.n482 9.3005
R542 source.n481 source.n480 9.3005
R543 source.n432 source.n431 9.3005
R544 source.n475 source.n474 9.3005
R545 source.n473 source.n472 9.3005
R546 source.n449 source.n448 9.3005
R547 source.n444 source.n443 9.3005
R548 source.n455 source.n454 9.3005
R549 source.n457 source.n456 9.3005
R550 source.n440 source.n439 9.3005
R551 source.n463 source.n462 9.3005
R552 source.n465 source.n464 9.3005
R553 source.n466 source.n435 9.3005
R554 source.n423 source.n422 9.3005
R555 source.n362 source.n361 9.3005
R556 source.n417 source.n416 9.3005
R557 source.n415 source.n414 9.3005
R558 source.n366 source.n365 9.3005
R559 source.n409 source.n408 9.3005
R560 source.n407 source.n406 9.3005
R561 source.n383 source.n382 9.3005
R562 source.n378 source.n377 9.3005
R563 source.n389 source.n388 9.3005
R564 source.n391 source.n390 9.3005
R565 source.n374 source.n373 9.3005
R566 source.n397 source.n396 9.3005
R567 source.n399 source.n398 9.3005
R568 source.n400 source.n369 9.3005
R569 source.n347 source.n346 9.3005
R570 source.n286 source.n285 9.3005
R571 source.n341 source.n340 9.3005
R572 source.n339 source.n338 9.3005
R573 source.n290 source.n289 9.3005
R574 source.n333 source.n332 9.3005
R575 source.n331 source.n330 9.3005
R576 source.n307 source.n306 9.3005
R577 source.n302 source.n301 9.3005
R578 source.n313 source.n312 9.3005
R579 source.n315 source.n314 9.3005
R580 source.n298 source.n297 9.3005
R581 source.n321 source.n320 9.3005
R582 source.n323 source.n322 9.3005
R583 source.n324 source.n293 9.3005
R584 source.n24 source.n23 9.3005
R585 source.n19 source.n18 9.3005
R586 source.n30 source.n29 9.3005
R587 source.n32 source.n31 9.3005
R588 source.n15 source.n14 9.3005
R589 source.n38 source.n37 9.3005
R590 source.n40 source.n39 9.3005
R591 source.n12 source.n9 9.3005
R592 source.n63 source.n62 9.3005
R593 source.n2 source.n1 9.3005
R594 source.n57 source.n56 9.3005
R595 source.n55 source.n54 9.3005
R596 source.n6 source.n5 9.3005
R597 source.n49 source.n48 9.3005
R598 source.n47 source.n46 9.3005
R599 source.n100 source.n99 9.3005
R600 source.n95 source.n94 9.3005
R601 source.n106 source.n105 9.3005
R602 source.n108 source.n107 9.3005
R603 source.n91 source.n90 9.3005
R604 source.n114 source.n113 9.3005
R605 source.n116 source.n115 9.3005
R606 source.n88 source.n85 9.3005
R607 source.n139 source.n138 9.3005
R608 source.n78 source.n77 9.3005
R609 source.n133 source.n132 9.3005
R610 source.n131 source.n130 9.3005
R611 source.n82 source.n81 9.3005
R612 source.n125 source.n124 9.3005
R613 source.n123 source.n122 9.3005
R614 source.n166 source.n165 9.3005
R615 source.n161 source.n160 9.3005
R616 source.n172 source.n171 9.3005
R617 source.n174 source.n173 9.3005
R618 source.n157 source.n156 9.3005
R619 source.n180 source.n179 9.3005
R620 source.n182 source.n181 9.3005
R621 source.n154 source.n151 9.3005
R622 source.n205 source.n204 9.3005
R623 source.n144 source.n143 9.3005
R624 source.n199 source.n198 9.3005
R625 source.n197 source.n196 9.3005
R626 source.n148 source.n147 9.3005
R627 source.n191 source.n190 9.3005
R628 source.n189 source.n188 9.3005
R629 source.n242 source.n241 9.3005
R630 source.n237 source.n236 9.3005
R631 source.n248 source.n247 9.3005
R632 source.n250 source.n249 9.3005
R633 source.n233 source.n232 9.3005
R634 source.n256 source.n255 9.3005
R635 source.n258 source.n257 9.3005
R636 source.n230 source.n227 9.3005
R637 source.n281 source.n280 9.3005
R638 source.n220 source.n219 9.3005
R639 source.n275 source.n274 9.3005
R640 source.n273 source.n272 9.3005
R641 source.n224 source.n223 9.3005
R642 source.n267 source.n266 9.3005
R643 source.n265 source.n264 9.3005
R644 source.n530 source.n529 8.92171
R645 source.n563 source.n504 8.92171
R646 source.n454 source.n453 8.92171
R647 source.n487 source.n428 8.92171
R648 source.n388 source.n387 8.92171
R649 source.n421 source.n362 8.92171
R650 source.n312 source.n311 8.92171
R651 source.n345 source.n286 8.92171
R652 source.n61 source.n2 8.92171
R653 source.n29 source.n28 8.92171
R654 source.n137 source.n78 8.92171
R655 source.n105 source.n104 8.92171
R656 source.n203 source.n144 8.92171
R657 source.n171 source.n170 8.92171
R658 source.n279 source.n220 8.92171
R659 source.n247 source.n246 8.92171
R660 source.n526 source.n520 8.14595
R661 source.n564 source.n502 8.14595
R662 source.n450 source.n444 8.14595
R663 source.n488 source.n426 8.14595
R664 source.n384 source.n378 8.14595
R665 source.n422 source.n360 8.14595
R666 source.n308 source.n302 8.14595
R667 source.n346 source.n284 8.14595
R668 source.n62 source.n0 8.14595
R669 source.n25 source.n19 8.14595
R670 source.n138 source.n76 8.14595
R671 source.n101 source.n95 8.14595
R672 source.n204 source.n142 8.14595
R673 source.n167 source.n161 8.14595
R674 source.n280 source.n218 8.14595
R675 source.n243 source.n237 8.14595
R676 source.n525 source.n522 7.3702
R677 source.n449 source.n446 7.3702
R678 source.n383 source.n380 7.3702
R679 source.n307 source.n304 7.3702
R680 source.n24 source.n21 7.3702
R681 source.n100 source.n97 7.3702
R682 source.n166 source.n163 7.3702
R683 source.n242 source.n239 7.3702
R684 source.n526 source.n525 5.81868
R685 source.n566 source.n502 5.81868
R686 source.n450 source.n449 5.81868
R687 source.n490 source.n426 5.81868
R688 source.n384 source.n383 5.81868
R689 source.n424 source.n360 5.81868
R690 source.n308 source.n307 5.81868
R691 source.n348 source.n284 5.81868
R692 source.n64 source.n0 5.81868
R693 source.n25 source.n24 5.81868
R694 source.n140 source.n76 5.81868
R695 source.n101 source.n100 5.81868
R696 source.n206 source.n142 5.81868
R697 source.n167 source.n166 5.81868
R698 source.n282 source.n218 5.81868
R699 source.n243 source.n242 5.81868
R700 source.n568 source.n567 5.51343
R701 source.n529 source.n520 5.04292
R702 source.n564 source.n563 5.04292
R703 source.n453 source.n444 5.04292
R704 source.n488 source.n487 5.04292
R705 source.n387 source.n378 5.04292
R706 source.n422 source.n421 5.04292
R707 source.n311 source.n302 5.04292
R708 source.n346 source.n345 5.04292
R709 source.n62 source.n61 5.04292
R710 source.n28 source.n19 5.04292
R711 source.n138 source.n137 5.04292
R712 source.n104 source.n95 5.04292
R713 source.n204 source.n203 5.04292
R714 source.n170 source.n161 5.04292
R715 source.n280 source.n279 5.04292
R716 source.n246 source.n237 5.04292
R717 source.n530 source.n518 4.26717
R718 source.n560 source.n504 4.26717
R719 source.n454 source.n442 4.26717
R720 source.n484 source.n428 4.26717
R721 source.n388 source.n376 4.26717
R722 source.n418 source.n362 4.26717
R723 source.n312 source.n300 4.26717
R724 source.n342 source.n286 4.26717
R725 source.n58 source.n2 4.26717
R726 source.n29 source.n17 4.26717
R727 source.n134 source.n78 4.26717
R728 source.n105 source.n93 4.26717
R729 source.n200 source.n144 4.26717
R730 source.n171 source.n159 4.26717
R731 source.n276 source.n220 4.26717
R732 source.n247 source.n235 4.26717
R733 source.n534 source.n533 3.49141
R734 source.n559 source.n506 3.49141
R735 source.n458 source.n457 3.49141
R736 source.n483 source.n430 3.49141
R737 source.n392 source.n391 3.49141
R738 source.n417 source.n364 3.49141
R739 source.n316 source.n315 3.49141
R740 source.n341 source.n288 3.49141
R741 source.n57 source.n4 3.49141
R742 source.n33 source.n32 3.49141
R743 source.n133 source.n80 3.49141
R744 source.n109 source.n108 3.49141
R745 source.n199 source.n146 3.49141
R746 source.n175 source.n174 3.49141
R747 source.n275 source.n222 3.49141
R748 source.n251 source.n250 3.49141
R749 source.n524 source.n523 2.84303
R750 source.n448 source.n447 2.84303
R751 source.n382 source.n381 2.84303
R752 source.n306 source.n305 2.84303
R753 source.n23 source.n22 2.84303
R754 source.n99 source.n98 2.84303
R755 source.n165 source.n164 2.84303
R756 source.n241 source.n240 2.84303
R757 source.n537 source.n516 2.71565
R758 source.n556 source.n555 2.71565
R759 source.n461 source.n440 2.71565
R760 source.n480 source.n479 2.71565
R761 source.n395 source.n374 2.71565
R762 source.n414 source.n413 2.71565
R763 source.n319 source.n298 2.71565
R764 source.n338 source.n337 2.71565
R765 source.n54 source.n53 2.71565
R766 source.n36 source.n15 2.71565
R767 source.n130 source.n129 2.71565
R768 source.n112 source.n91 2.71565
R769 source.n196 source.n195 2.71565
R770 source.n178 source.n157 2.71565
R771 source.n272 source.n271 2.71565
R772 source.n254 source.n233 2.71565
R773 source.n538 source.n514 1.93989
R774 source.n552 source.n508 1.93989
R775 source.n462 source.n438 1.93989
R776 source.n476 source.n432 1.93989
R777 source.n396 source.n372 1.93989
R778 source.n410 source.n366 1.93989
R779 source.n320 source.n296 1.93989
R780 source.n334 source.n290 1.93989
R781 source.n50 source.n6 1.93989
R782 source.n37 source.n13 1.93989
R783 source.n126 source.n82 1.93989
R784 source.n113 source.n89 1.93989
R785 source.n192 source.n148 1.93989
R786 source.n179 source.n155 1.93989
R787 source.n268 source.n224 1.93989
R788 source.n255 source.n231 1.93989
R789 source.n500 source.t7 1.6505
R790 source.n500 source.t4 1.6505
R791 source.n498 source.t14 1.6505
R792 source.n498 source.t9 1.6505
R793 source.n496 source.t3 1.6505
R794 source.n496 source.t19 1.6505
R795 source.n494 source.t16 1.6505
R796 source.n494 source.t2 1.6505
R797 source.n492 source.t1 1.6505
R798 source.n492 source.t22 1.6505
R799 source.n358 source.t32 1.6505
R800 source.n358 source.t30 1.6505
R801 source.n356 source.t46 1.6505
R802 source.n356 source.t34 1.6505
R803 source.n354 source.t38 1.6505
R804 source.n354 source.t26 1.6505
R805 source.n352 source.t28 1.6505
R806 source.n352 source.t33 1.6505
R807 source.n350 source.t41 1.6505
R808 source.n350 source.t25 1.6505
R809 source.n66 source.t47 1.6505
R810 source.n66 source.t43 1.6505
R811 source.n68 source.t36 1.6505
R812 source.n68 source.t37 1.6505
R813 source.n70 source.t35 1.6505
R814 source.n70 source.t27 1.6505
R815 source.n72 source.t31 1.6505
R816 source.n72 source.t29 1.6505
R817 source.n74 source.t39 1.6505
R818 source.n74 source.t42 1.6505
R819 source.n208 source.t20 1.6505
R820 source.n208 source.t15 1.6505
R821 source.n210 source.t10 1.6505
R822 source.n210 source.t11 1.6505
R823 source.n212 source.t13 1.6505
R824 source.n212 source.t12 1.6505
R825 source.n214 source.t5 1.6505
R826 source.n214 source.t21 1.6505
R827 source.n216 source.t0 1.6505
R828 source.n216 source.t17 1.6505
R829 source.n543 source.n541 1.16414
R830 source.n551 source.n510 1.16414
R831 source.n467 source.n465 1.16414
R832 source.n475 source.n434 1.16414
R833 source.n401 source.n399 1.16414
R834 source.n409 source.n368 1.16414
R835 source.n325 source.n323 1.16414
R836 source.n333 source.n292 1.16414
R837 source.n49 source.n8 1.16414
R838 source.n41 source.n40 1.16414
R839 source.n125 source.n84 1.16414
R840 source.n117 source.n116 1.16414
R841 source.n191 source.n150 1.16414
R842 source.n183 source.n182 1.16414
R843 source.n267 source.n226 1.16414
R844 source.n259 source.n258 1.16414
R845 source.n283 source.n217 0.5005
R846 source.n217 source.n215 0.5005
R847 source.n215 source.n213 0.5005
R848 source.n213 source.n211 0.5005
R849 source.n211 source.n209 0.5005
R850 source.n209 source.n207 0.5005
R851 source.n141 source.n75 0.5005
R852 source.n75 source.n73 0.5005
R853 source.n73 source.n71 0.5005
R854 source.n71 source.n69 0.5005
R855 source.n69 source.n67 0.5005
R856 source.n67 source.n65 0.5005
R857 source.n351 source.n349 0.5005
R858 source.n353 source.n351 0.5005
R859 source.n355 source.n353 0.5005
R860 source.n357 source.n355 0.5005
R861 source.n359 source.n357 0.5005
R862 source.n425 source.n359 0.5005
R863 source.n493 source.n491 0.5005
R864 source.n495 source.n493 0.5005
R865 source.n497 source.n495 0.5005
R866 source.n499 source.n497 0.5005
R867 source.n501 source.n499 0.5005
R868 source.n567 source.n501 0.5005
R869 source.n207 source.n141 0.470328
R870 source.n491 source.n425 0.470328
R871 source.n542 source.n512 0.388379
R872 source.n548 source.n547 0.388379
R873 source.n466 source.n436 0.388379
R874 source.n472 source.n471 0.388379
R875 source.n400 source.n370 0.388379
R876 source.n406 source.n405 0.388379
R877 source.n324 source.n294 0.388379
R878 source.n330 source.n329 0.388379
R879 source.n46 source.n45 0.388379
R880 source.n12 source.n10 0.388379
R881 source.n122 source.n121 0.388379
R882 source.n88 source.n86 0.388379
R883 source.n188 source.n187 0.388379
R884 source.n154 source.n152 0.388379
R885 source.n264 source.n263 0.388379
R886 source.n230 source.n228 0.388379
R887 source source.n568 0.188
R888 source.n524 source.n519 0.155672
R889 source.n531 source.n519 0.155672
R890 source.n532 source.n531 0.155672
R891 source.n532 source.n515 0.155672
R892 source.n539 source.n515 0.155672
R893 source.n540 source.n539 0.155672
R894 source.n540 source.n511 0.155672
R895 source.n549 source.n511 0.155672
R896 source.n550 source.n549 0.155672
R897 source.n550 source.n507 0.155672
R898 source.n557 source.n507 0.155672
R899 source.n558 source.n557 0.155672
R900 source.n558 source.n503 0.155672
R901 source.n565 source.n503 0.155672
R902 source.n448 source.n443 0.155672
R903 source.n455 source.n443 0.155672
R904 source.n456 source.n455 0.155672
R905 source.n456 source.n439 0.155672
R906 source.n463 source.n439 0.155672
R907 source.n464 source.n463 0.155672
R908 source.n464 source.n435 0.155672
R909 source.n473 source.n435 0.155672
R910 source.n474 source.n473 0.155672
R911 source.n474 source.n431 0.155672
R912 source.n481 source.n431 0.155672
R913 source.n482 source.n481 0.155672
R914 source.n482 source.n427 0.155672
R915 source.n489 source.n427 0.155672
R916 source.n382 source.n377 0.155672
R917 source.n389 source.n377 0.155672
R918 source.n390 source.n389 0.155672
R919 source.n390 source.n373 0.155672
R920 source.n397 source.n373 0.155672
R921 source.n398 source.n397 0.155672
R922 source.n398 source.n369 0.155672
R923 source.n407 source.n369 0.155672
R924 source.n408 source.n407 0.155672
R925 source.n408 source.n365 0.155672
R926 source.n415 source.n365 0.155672
R927 source.n416 source.n415 0.155672
R928 source.n416 source.n361 0.155672
R929 source.n423 source.n361 0.155672
R930 source.n306 source.n301 0.155672
R931 source.n313 source.n301 0.155672
R932 source.n314 source.n313 0.155672
R933 source.n314 source.n297 0.155672
R934 source.n321 source.n297 0.155672
R935 source.n322 source.n321 0.155672
R936 source.n322 source.n293 0.155672
R937 source.n331 source.n293 0.155672
R938 source.n332 source.n331 0.155672
R939 source.n332 source.n289 0.155672
R940 source.n339 source.n289 0.155672
R941 source.n340 source.n339 0.155672
R942 source.n340 source.n285 0.155672
R943 source.n347 source.n285 0.155672
R944 source.n63 source.n1 0.155672
R945 source.n56 source.n1 0.155672
R946 source.n56 source.n55 0.155672
R947 source.n55 source.n5 0.155672
R948 source.n48 source.n5 0.155672
R949 source.n48 source.n47 0.155672
R950 source.n47 source.n9 0.155672
R951 source.n39 source.n9 0.155672
R952 source.n39 source.n38 0.155672
R953 source.n38 source.n14 0.155672
R954 source.n31 source.n14 0.155672
R955 source.n31 source.n30 0.155672
R956 source.n30 source.n18 0.155672
R957 source.n23 source.n18 0.155672
R958 source.n139 source.n77 0.155672
R959 source.n132 source.n77 0.155672
R960 source.n132 source.n131 0.155672
R961 source.n131 source.n81 0.155672
R962 source.n124 source.n81 0.155672
R963 source.n124 source.n123 0.155672
R964 source.n123 source.n85 0.155672
R965 source.n115 source.n85 0.155672
R966 source.n115 source.n114 0.155672
R967 source.n114 source.n90 0.155672
R968 source.n107 source.n90 0.155672
R969 source.n107 source.n106 0.155672
R970 source.n106 source.n94 0.155672
R971 source.n99 source.n94 0.155672
R972 source.n205 source.n143 0.155672
R973 source.n198 source.n143 0.155672
R974 source.n198 source.n197 0.155672
R975 source.n197 source.n147 0.155672
R976 source.n190 source.n147 0.155672
R977 source.n190 source.n189 0.155672
R978 source.n189 source.n151 0.155672
R979 source.n181 source.n151 0.155672
R980 source.n181 source.n180 0.155672
R981 source.n180 source.n156 0.155672
R982 source.n173 source.n156 0.155672
R983 source.n173 source.n172 0.155672
R984 source.n172 source.n160 0.155672
R985 source.n165 source.n160 0.155672
R986 source.n281 source.n219 0.155672
R987 source.n274 source.n219 0.155672
R988 source.n274 source.n273 0.155672
R989 source.n273 source.n223 0.155672
R990 source.n266 source.n223 0.155672
R991 source.n266 source.n265 0.155672
R992 source.n265 source.n227 0.155672
R993 source.n257 source.n227 0.155672
R994 source.n257 source.n256 0.155672
R995 source.n256 source.n232 0.155672
R996 source.n249 source.n232 0.155672
R997 source.n249 source.n248 0.155672
R998 source.n248 source.n236 0.155672
R999 source.n241 source.n236 0.155672
R1000 drain_left.n13 drain_left.n11 60.0527
R1001 drain_left.n7 drain_left.n5 60.0525
R1002 drain_left.n2 drain_left.n0 60.0525
R1003 drain_left.n19 drain_left.n18 59.5527
R1004 drain_left.n17 drain_left.n16 59.5527
R1005 drain_left.n15 drain_left.n14 59.5527
R1006 drain_left.n13 drain_left.n12 59.5527
R1007 drain_left.n7 drain_left.n6 59.5525
R1008 drain_left.n9 drain_left.n8 59.5525
R1009 drain_left.n4 drain_left.n3 59.5525
R1010 drain_left.n2 drain_left.n1 59.5525
R1011 drain_left.n21 drain_left.n20 59.5525
R1012 drain_left drain_left.n10 32.1171
R1013 drain_left drain_left.n21 6.15322
R1014 drain_left.n5 drain_left.t5 1.6505
R1015 drain_left.n5 drain_left.t2 1.6505
R1016 drain_left.n6 drain_left.t0 1.6505
R1017 drain_left.n6 drain_left.t15 1.6505
R1018 drain_left.n8 drain_left.t3 1.6505
R1019 drain_left.n8 drain_left.t18 1.6505
R1020 drain_left.n3 drain_left.t16 1.6505
R1021 drain_left.n3 drain_left.t6 1.6505
R1022 drain_left.n1 drain_left.t8 1.6505
R1023 drain_left.n1 drain_left.t4 1.6505
R1024 drain_left.n0 drain_left.t14 1.6505
R1025 drain_left.n0 drain_left.t10 1.6505
R1026 drain_left.n20 drain_left.t9 1.6505
R1027 drain_left.n20 drain_left.t21 1.6505
R1028 drain_left.n18 drain_left.t7 1.6505
R1029 drain_left.n18 drain_left.t20 1.6505
R1030 drain_left.n16 drain_left.t13 1.6505
R1031 drain_left.n16 drain_left.t19 1.6505
R1032 drain_left.n14 drain_left.t12 1.6505
R1033 drain_left.n14 drain_left.t1 1.6505
R1034 drain_left.n12 drain_left.t11 1.6505
R1035 drain_left.n12 drain_left.t23 1.6505
R1036 drain_left.n11 drain_left.t17 1.6505
R1037 drain_left.n11 drain_left.t22 1.6505
R1038 drain_left.n9 drain_left.n7 0.5005
R1039 drain_left.n4 drain_left.n2 0.5005
R1040 drain_left.n15 drain_left.n13 0.5005
R1041 drain_left.n17 drain_left.n15 0.5005
R1042 drain_left.n19 drain_left.n17 0.5005
R1043 drain_left.n21 drain_left.n19 0.5005
R1044 drain_left.n10 drain_left.n9 0.195154
R1045 drain_left.n10 drain_left.n4 0.195154
R1046 minus.n33 minus.t13 1309.87
R1047 minus.n7 minus.t11 1309.87
R1048 minus.n68 minus.t14 1309.87
R1049 minus.n41 minus.t23 1309.87
R1050 minus.n32 minus.t2 1282.12
R1051 minus.n30 minus.t8 1282.12
R1052 minus.n3 minus.t21 1282.12
R1053 minus.n24 minus.t6 1282.12
R1054 minus.n22 minus.t20 1282.12
R1055 minus.n4 minus.t7 1282.12
R1056 minus.n17 minus.t19 1282.12
R1057 minus.n15 minus.t0 1282.12
R1058 minus.n8 minus.t10 1282.12
R1059 minus.n9 minus.t1 1282.12
R1060 minus.n67 minus.t18 1282.12
R1061 minus.n65 minus.t4 1282.12
R1062 minus.n59 minus.t9 1282.12
R1063 minus.n58 minus.t15 1282.12
R1064 minus.n56 minus.t16 1282.12
R1065 minus.n38 minus.t22 1282.12
R1066 minus.n51 minus.t5 1282.12
R1067 minus.n49 minus.t12 1282.12
R1068 minus.n43 minus.t17 1282.12
R1069 minus.n42 minus.t3 1282.12
R1070 minus.n11 minus.n7 161.489
R1071 minus.n45 minus.n41 161.489
R1072 minus.n34 minus.n33 161.3
R1073 minus.n31 minus.n0 161.3
R1074 minus.n29 minus.n28 161.3
R1075 minus.n27 minus.n1 161.3
R1076 minus.n26 minus.n25 161.3
R1077 minus.n23 minus.n2 161.3
R1078 minus.n21 minus.n20 161.3
R1079 minus.n19 minus.n18 161.3
R1080 minus.n16 minus.n5 161.3
R1081 minus.n14 minus.n13 161.3
R1082 minus.n12 minus.n6 161.3
R1083 minus.n11 minus.n10 161.3
R1084 minus.n69 minus.n68 161.3
R1085 minus.n66 minus.n35 161.3
R1086 minus.n64 minus.n63 161.3
R1087 minus.n62 minus.n36 161.3
R1088 minus.n61 minus.n60 161.3
R1089 minus.n57 minus.n37 161.3
R1090 minus.n55 minus.n54 161.3
R1091 minus.n53 minus.n52 161.3
R1092 minus.n50 minus.n39 161.3
R1093 minus.n48 minus.n47 161.3
R1094 minus.n46 minus.n40 161.3
R1095 minus.n45 minus.n44 161.3
R1096 minus.n29 minus.n1 73.0308
R1097 minus.n14 minus.n6 73.0308
R1098 minus.n48 minus.n40 73.0308
R1099 minus.n64 minus.n36 73.0308
R1100 minus.n31 minus.n30 68.649
R1101 minus.n10 minus.n8 68.649
R1102 minus.n44 minus.n43 68.649
R1103 minus.n66 minus.n65 68.649
R1104 minus.n25 minus.n3 65.7278
R1105 minus.n16 minus.n15 65.7278
R1106 minus.n50 minus.n49 65.7278
R1107 minus.n60 minus.n59 65.7278
R1108 minus.n33 minus.n32 56.9641
R1109 minus.n9 minus.n7 56.9641
R1110 minus.n42 minus.n41 56.9641
R1111 minus.n68 minus.n67 56.9641
R1112 minus.n24 minus.n23 54.0429
R1113 minus.n18 minus.n17 54.0429
R1114 minus.n52 minus.n51 54.0429
R1115 minus.n58 minus.n57 54.0429
R1116 minus.n22 minus.n21 42.3581
R1117 minus.n21 minus.n4 42.3581
R1118 minus.n55 minus.n38 42.3581
R1119 minus.n56 minus.n55 42.3581
R1120 minus.n70 minus.n34 37.4778
R1121 minus.n23 minus.n22 30.6732
R1122 minus.n18 minus.n4 30.6732
R1123 minus.n52 minus.n38 30.6732
R1124 minus.n57 minus.n56 30.6732
R1125 minus.n25 minus.n24 18.9884
R1126 minus.n17 minus.n16 18.9884
R1127 minus.n51 minus.n50 18.9884
R1128 minus.n60 minus.n58 18.9884
R1129 minus.n32 minus.n31 16.0672
R1130 minus.n10 minus.n9 16.0672
R1131 minus.n44 minus.n42 16.0672
R1132 minus.n67 minus.n66 16.0672
R1133 minus.n3 minus.n1 7.30353
R1134 minus.n15 minus.n14 7.30353
R1135 minus.n49 minus.n48 7.30353
R1136 minus.n59 minus.n36 7.30353
R1137 minus.n70 minus.n69 6.43232
R1138 minus.n30 minus.n29 4.38232
R1139 minus.n8 minus.n6 4.38232
R1140 minus.n43 minus.n40 4.38232
R1141 minus.n65 minus.n64 4.38232
R1142 minus.n34 minus.n0 0.189894
R1143 minus.n28 minus.n0 0.189894
R1144 minus.n28 minus.n27 0.189894
R1145 minus.n27 minus.n26 0.189894
R1146 minus.n26 minus.n2 0.189894
R1147 minus.n20 minus.n2 0.189894
R1148 minus.n20 minus.n19 0.189894
R1149 minus.n19 minus.n5 0.189894
R1150 minus.n13 minus.n5 0.189894
R1151 minus.n13 minus.n12 0.189894
R1152 minus.n12 minus.n11 0.189894
R1153 minus.n46 minus.n45 0.189894
R1154 minus.n47 minus.n46 0.189894
R1155 minus.n47 minus.n39 0.189894
R1156 minus.n53 minus.n39 0.189894
R1157 minus.n54 minus.n53 0.189894
R1158 minus.n54 minus.n37 0.189894
R1159 minus.n61 minus.n37 0.189894
R1160 minus.n62 minus.n61 0.189894
R1161 minus.n63 minus.n62 0.189894
R1162 minus.n63 minus.n35 0.189894
R1163 minus.n69 minus.n35 0.189894
R1164 minus minus.n70 0.188
R1165 drain_right.n7 drain_right.n5 60.0525
R1166 drain_right.n2 drain_right.n0 60.0525
R1167 drain_right.n13 drain_right.n11 60.0525
R1168 drain_right.n13 drain_right.n12 59.5527
R1169 drain_right.n15 drain_right.n14 59.5527
R1170 drain_right.n17 drain_right.n16 59.5527
R1171 drain_right.n19 drain_right.n18 59.5527
R1172 drain_right.n21 drain_right.n20 59.5527
R1173 drain_right.n7 drain_right.n6 59.5525
R1174 drain_right.n9 drain_right.n8 59.5525
R1175 drain_right.n4 drain_right.n3 59.5525
R1176 drain_right.n2 drain_right.n1 59.5525
R1177 drain_right drain_right.n10 31.5638
R1178 drain_right drain_right.n21 6.15322
R1179 drain_right.n5 drain_right.t5 1.6505
R1180 drain_right.n5 drain_right.t9 1.6505
R1181 drain_right.n6 drain_right.t14 1.6505
R1182 drain_right.n6 drain_right.t19 1.6505
R1183 drain_right.n8 drain_right.t7 1.6505
R1184 drain_right.n8 drain_right.t8 1.6505
R1185 drain_right.n3 drain_right.t18 1.6505
R1186 drain_right.n3 drain_right.t1 1.6505
R1187 drain_right.n1 drain_right.t6 1.6505
R1188 drain_right.n1 drain_right.t11 1.6505
R1189 drain_right.n0 drain_right.t0 1.6505
R1190 drain_right.n0 drain_right.t20 1.6505
R1191 drain_right.n11 drain_right.t22 1.6505
R1192 drain_right.n11 drain_right.t12 1.6505
R1193 drain_right.n12 drain_right.t23 1.6505
R1194 drain_right.n12 drain_right.t13 1.6505
R1195 drain_right.n14 drain_right.t16 1.6505
R1196 drain_right.n14 drain_right.t4 1.6505
R1197 drain_right.n16 drain_right.t17 1.6505
R1198 drain_right.n16 drain_right.t3 1.6505
R1199 drain_right.n18 drain_right.t15 1.6505
R1200 drain_right.n18 drain_right.t2 1.6505
R1201 drain_right.n20 drain_right.t10 1.6505
R1202 drain_right.n20 drain_right.t21 1.6505
R1203 drain_right.n9 drain_right.n7 0.5005
R1204 drain_right.n4 drain_right.n2 0.5005
R1205 drain_right.n21 drain_right.n19 0.5005
R1206 drain_right.n19 drain_right.n17 0.5005
R1207 drain_right.n17 drain_right.n15 0.5005
R1208 drain_right.n15 drain_right.n13 0.5005
R1209 drain_right.n10 drain_right.n9 0.195154
R1210 drain_right.n10 drain_right.n4 0.195154
C0 plus minus 5.93414f
C1 drain_left minus 0.172313f
C2 plus source 7.11409f
C3 drain_left source 48.549397f
C4 drain_right plus 0.374075f
C5 drain_left drain_right 1.19771f
C6 minus source 7.10006f
C7 drain_left plus 7.57399f
C8 drain_right minus 7.35532f
C9 drain_right source 48.5498f
C10 drain_right a_n2224_n3288# 7.39055f
C11 drain_left a_n2224_n3288# 7.72916f
C12 source a_n2224_n3288# 8.828288f
C13 minus a_n2224_n3288# 8.72191f
C14 plus a_n2224_n3288# 10.796109f
C15 drain_right.t0 a_n2224_n3288# 0.344517f
C16 drain_right.t20 a_n2224_n3288# 0.344517f
C17 drain_right.n0 a_n2224_n3288# 3.0693f
C18 drain_right.t6 a_n2224_n3288# 0.344517f
C19 drain_right.t11 a_n2224_n3288# 0.344517f
C20 drain_right.n1 a_n2224_n3288# 3.06567f
C21 drain_right.n2 a_n2224_n3288# 0.854948f
C22 drain_right.t18 a_n2224_n3288# 0.344517f
C23 drain_right.t1 a_n2224_n3288# 0.344517f
C24 drain_right.n3 a_n2224_n3288# 3.06567f
C25 drain_right.n4 a_n2224_n3288# 0.390556f
C26 drain_right.t5 a_n2224_n3288# 0.344517f
C27 drain_right.t9 a_n2224_n3288# 0.344517f
C28 drain_right.n5 a_n2224_n3288# 3.0693f
C29 drain_right.t14 a_n2224_n3288# 0.344517f
C30 drain_right.t19 a_n2224_n3288# 0.344517f
C31 drain_right.n6 a_n2224_n3288# 3.06567f
C32 drain_right.n7 a_n2224_n3288# 0.854948f
C33 drain_right.t7 a_n2224_n3288# 0.344517f
C34 drain_right.t8 a_n2224_n3288# 0.344517f
C35 drain_right.n8 a_n2224_n3288# 3.06567f
C36 drain_right.n9 a_n2224_n3288# 0.390556f
C37 drain_right.n10 a_n2224_n3288# 1.84247f
C38 drain_right.t22 a_n2224_n3288# 0.344517f
C39 drain_right.t12 a_n2224_n3288# 0.344517f
C40 drain_right.n11 a_n2224_n3288# 3.0693f
C41 drain_right.t23 a_n2224_n3288# 0.344517f
C42 drain_right.t13 a_n2224_n3288# 0.344517f
C43 drain_right.n12 a_n2224_n3288# 3.06568f
C44 drain_right.n13 a_n2224_n3288# 0.854935f
C45 drain_right.t16 a_n2224_n3288# 0.344517f
C46 drain_right.t4 a_n2224_n3288# 0.344517f
C47 drain_right.n14 a_n2224_n3288# 3.06568f
C48 drain_right.n15 a_n2224_n3288# 0.421962f
C49 drain_right.t17 a_n2224_n3288# 0.344517f
C50 drain_right.t3 a_n2224_n3288# 0.344517f
C51 drain_right.n16 a_n2224_n3288# 3.06568f
C52 drain_right.n17 a_n2224_n3288# 0.421962f
C53 drain_right.t15 a_n2224_n3288# 0.344517f
C54 drain_right.t2 a_n2224_n3288# 0.344517f
C55 drain_right.n18 a_n2224_n3288# 3.06568f
C56 drain_right.n19 a_n2224_n3288# 0.421962f
C57 drain_right.t10 a_n2224_n3288# 0.344517f
C58 drain_right.t21 a_n2224_n3288# 0.344517f
C59 drain_right.n20 a_n2224_n3288# 3.06568f
C60 drain_right.n21 a_n2224_n3288# 0.721849f
C61 minus.n0 a_n2224_n3288# 0.049933f
C62 minus.t13 a_n2224_n3288# 0.426875f
C63 minus.t2 a_n2224_n3288# 0.423302f
C64 minus.t8 a_n2224_n3288# 0.423302f
C65 minus.n1 a_n2224_n3288# 0.018104f
C66 minus.n2 a_n2224_n3288# 0.049933f
C67 minus.t21 a_n2224_n3288# 0.423302f
C68 minus.n3 a_n2224_n3288# 0.170487f
C69 minus.t6 a_n2224_n3288# 0.423302f
C70 minus.t20 a_n2224_n3288# 0.423302f
C71 minus.t7 a_n2224_n3288# 0.423302f
C72 minus.n4 a_n2224_n3288# 0.170487f
C73 minus.n5 a_n2224_n3288# 0.049933f
C74 minus.t19 a_n2224_n3288# 0.423302f
C75 minus.t0 a_n2224_n3288# 0.423302f
C76 minus.n6 a_n2224_n3288# 0.017488f
C77 minus.t11 a_n2224_n3288# 0.426875f
C78 minus.n7 a_n2224_n3288# 0.184158f
C79 minus.t10 a_n2224_n3288# 0.423302f
C80 minus.n8 a_n2224_n3288# 0.170487f
C81 minus.t1 a_n2224_n3288# 0.423302f
C82 minus.n9 a_n2224_n3288# 0.170487f
C83 minus.n10 a_n2224_n3288# 0.019027f
C84 minus.n11 a_n2224_n3288# 0.103804f
C85 minus.n12 a_n2224_n3288# 0.049933f
C86 minus.n13 a_n2224_n3288# 0.049933f
C87 minus.n14 a_n2224_n3288# 0.018104f
C88 minus.n15 a_n2224_n3288# 0.170487f
C89 minus.n16 a_n2224_n3288# 0.019027f
C90 minus.n17 a_n2224_n3288# 0.170487f
C91 minus.n18 a_n2224_n3288# 0.019027f
C92 minus.n19 a_n2224_n3288# 0.049933f
C93 minus.n20 a_n2224_n3288# 0.049933f
C94 minus.n21 a_n2224_n3288# 0.019027f
C95 minus.n22 a_n2224_n3288# 0.170487f
C96 minus.n23 a_n2224_n3288# 0.019027f
C97 minus.n24 a_n2224_n3288# 0.170487f
C98 minus.n25 a_n2224_n3288# 0.019027f
C99 minus.n26 a_n2224_n3288# 0.049933f
C100 minus.n27 a_n2224_n3288# 0.049933f
C101 minus.n28 a_n2224_n3288# 0.049933f
C102 minus.n29 a_n2224_n3288# 0.017488f
C103 minus.n30 a_n2224_n3288# 0.170487f
C104 minus.n31 a_n2224_n3288# 0.019027f
C105 minus.n32 a_n2224_n3288# 0.170487f
C106 minus.n33 a_n2224_n3288# 0.184094f
C107 minus.n34 a_n2224_n3288# 1.86026f
C108 minus.n35 a_n2224_n3288# 0.049933f
C109 minus.t18 a_n2224_n3288# 0.423302f
C110 minus.t4 a_n2224_n3288# 0.423302f
C111 minus.n36 a_n2224_n3288# 0.018104f
C112 minus.n37 a_n2224_n3288# 0.049933f
C113 minus.t15 a_n2224_n3288# 0.423302f
C114 minus.t16 a_n2224_n3288# 0.423302f
C115 minus.t22 a_n2224_n3288# 0.423302f
C116 minus.n38 a_n2224_n3288# 0.170487f
C117 minus.n39 a_n2224_n3288# 0.049933f
C118 minus.t5 a_n2224_n3288# 0.423302f
C119 minus.t12 a_n2224_n3288# 0.423302f
C120 minus.n40 a_n2224_n3288# 0.017488f
C121 minus.t23 a_n2224_n3288# 0.426875f
C122 minus.n41 a_n2224_n3288# 0.184158f
C123 minus.t3 a_n2224_n3288# 0.423302f
C124 minus.n42 a_n2224_n3288# 0.170487f
C125 minus.t17 a_n2224_n3288# 0.423302f
C126 minus.n43 a_n2224_n3288# 0.170487f
C127 minus.n44 a_n2224_n3288# 0.019027f
C128 minus.n45 a_n2224_n3288# 0.103804f
C129 minus.n46 a_n2224_n3288# 0.049933f
C130 minus.n47 a_n2224_n3288# 0.049933f
C131 minus.n48 a_n2224_n3288# 0.018104f
C132 minus.n49 a_n2224_n3288# 0.170487f
C133 minus.n50 a_n2224_n3288# 0.019027f
C134 minus.n51 a_n2224_n3288# 0.170487f
C135 minus.n52 a_n2224_n3288# 0.019027f
C136 minus.n53 a_n2224_n3288# 0.049933f
C137 minus.n54 a_n2224_n3288# 0.049933f
C138 minus.n55 a_n2224_n3288# 0.019027f
C139 minus.n56 a_n2224_n3288# 0.170487f
C140 minus.n57 a_n2224_n3288# 0.019027f
C141 minus.n58 a_n2224_n3288# 0.170487f
C142 minus.t9 a_n2224_n3288# 0.423302f
C143 minus.n59 a_n2224_n3288# 0.170487f
C144 minus.n60 a_n2224_n3288# 0.019027f
C145 minus.n61 a_n2224_n3288# 0.049933f
C146 minus.n62 a_n2224_n3288# 0.049933f
C147 minus.n63 a_n2224_n3288# 0.049933f
C148 minus.n64 a_n2224_n3288# 0.017488f
C149 minus.n65 a_n2224_n3288# 0.170487f
C150 minus.n66 a_n2224_n3288# 0.019027f
C151 minus.n67 a_n2224_n3288# 0.170487f
C152 minus.t14 a_n2224_n3288# 0.426875f
C153 minus.n68 a_n2224_n3288# 0.184094f
C154 minus.n69 a_n2224_n3288# 0.318459f
C155 minus.n70 a_n2224_n3288# 2.25368f
C156 drain_left.t14 a_n2224_n3288# 0.344873f
C157 drain_left.t10 a_n2224_n3288# 0.344873f
C158 drain_left.n0 a_n2224_n3288# 3.07247f
C159 drain_left.t8 a_n2224_n3288# 0.344873f
C160 drain_left.t4 a_n2224_n3288# 0.344873f
C161 drain_left.n1 a_n2224_n3288# 3.06883f
C162 drain_left.n2 a_n2224_n3288# 0.855831f
C163 drain_left.t16 a_n2224_n3288# 0.344873f
C164 drain_left.t6 a_n2224_n3288# 0.344873f
C165 drain_left.n3 a_n2224_n3288# 3.06883f
C166 drain_left.n4 a_n2224_n3288# 0.39096f
C167 drain_left.t5 a_n2224_n3288# 0.344873f
C168 drain_left.t2 a_n2224_n3288# 0.344873f
C169 drain_left.n5 a_n2224_n3288# 3.07247f
C170 drain_left.t0 a_n2224_n3288# 0.344873f
C171 drain_left.t15 a_n2224_n3288# 0.344873f
C172 drain_left.n6 a_n2224_n3288# 3.06883f
C173 drain_left.n7 a_n2224_n3288# 0.855831f
C174 drain_left.t3 a_n2224_n3288# 0.344873f
C175 drain_left.t18 a_n2224_n3288# 0.344873f
C176 drain_left.n8 a_n2224_n3288# 3.06883f
C177 drain_left.n9 a_n2224_n3288# 0.39096f
C178 drain_left.n10 a_n2224_n3288# 1.9193f
C179 drain_left.t17 a_n2224_n3288# 0.344873f
C180 drain_left.t22 a_n2224_n3288# 0.344873f
C181 drain_left.n11 a_n2224_n3288# 3.07249f
C182 drain_left.t11 a_n2224_n3288# 0.344873f
C183 drain_left.t23 a_n2224_n3288# 0.344873f
C184 drain_left.n12 a_n2224_n3288# 3.06885f
C185 drain_left.n13 a_n2224_n3288# 0.855806f
C186 drain_left.t12 a_n2224_n3288# 0.344873f
C187 drain_left.t1 a_n2224_n3288# 0.344873f
C188 drain_left.n14 a_n2224_n3288# 3.06885f
C189 drain_left.n15 a_n2224_n3288# 0.422398f
C190 drain_left.t13 a_n2224_n3288# 0.344873f
C191 drain_left.t19 a_n2224_n3288# 0.344873f
C192 drain_left.n16 a_n2224_n3288# 3.06885f
C193 drain_left.n17 a_n2224_n3288# 0.422398f
C194 drain_left.t7 a_n2224_n3288# 0.344873f
C195 drain_left.t20 a_n2224_n3288# 0.344873f
C196 drain_left.n18 a_n2224_n3288# 3.06885f
C197 drain_left.n19 a_n2224_n3288# 0.422398f
C198 drain_left.t9 a_n2224_n3288# 0.344873f
C199 drain_left.t21 a_n2224_n3288# 0.344873f
C200 drain_left.n20 a_n2224_n3288# 3.06883f
C201 drain_left.n21 a_n2224_n3288# 0.722607f
C202 source.n0 a_n2224_n3288# 0.042758f
C203 source.n1 a_n2224_n3288# 0.03228f
C204 source.n2 a_n2224_n3288# 0.017346f
C205 source.n3 a_n2224_n3288# 0.040999f
C206 source.n4 a_n2224_n3288# 0.018366f
C207 source.n5 a_n2224_n3288# 0.03228f
C208 source.n6 a_n2224_n3288# 0.017346f
C209 source.n7 a_n2224_n3288# 0.040999f
C210 source.n8 a_n2224_n3288# 0.018366f
C211 source.n9 a_n2224_n3288# 0.03228f
C212 source.n10 a_n2224_n3288# 0.017856f
C213 source.n11 a_n2224_n3288# 0.040999f
C214 source.n12 a_n2224_n3288# 0.017346f
C215 source.n13 a_n2224_n3288# 0.018366f
C216 source.n14 a_n2224_n3288# 0.03228f
C217 source.n15 a_n2224_n3288# 0.017346f
C218 source.n16 a_n2224_n3288# 0.040999f
C219 source.n17 a_n2224_n3288# 0.018366f
C220 source.n18 a_n2224_n3288# 0.03228f
C221 source.n19 a_n2224_n3288# 0.017346f
C222 source.n20 a_n2224_n3288# 0.030749f
C223 source.n21 a_n2224_n3288# 0.028983f
C224 source.t24 a_n2224_n3288# 0.069244f
C225 source.n22 a_n2224_n3288# 0.232733f
C226 source.n23 a_n2224_n3288# 1.62845f
C227 source.n24 a_n2224_n3288# 0.017346f
C228 source.n25 a_n2224_n3288# 0.018366f
C229 source.n26 a_n2224_n3288# 0.040999f
C230 source.n27 a_n2224_n3288# 0.040999f
C231 source.n28 a_n2224_n3288# 0.018366f
C232 source.n29 a_n2224_n3288# 0.017346f
C233 source.n30 a_n2224_n3288# 0.03228f
C234 source.n31 a_n2224_n3288# 0.03228f
C235 source.n32 a_n2224_n3288# 0.017346f
C236 source.n33 a_n2224_n3288# 0.018366f
C237 source.n34 a_n2224_n3288# 0.040999f
C238 source.n35 a_n2224_n3288# 0.040999f
C239 source.n36 a_n2224_n3288# 0.018366f
C240 source.n37 a_n2224_n3288# 0.017346f
C241 source.n38 a_n2224_n3288# 0.03228f
C242 source.n39 a_n2224_n3288# 0.03228f
C243 source.n40 a_n2224_n3288# 0.017346f
C244 source.n41 a_n2224_n3288# 0.018366f
C245 source.n42 a_n2224_n3288# 0.040999f
C246 source.n43 a_n2224_n3288# 0.040999f
C247 source.n44 a_n2224_n3288# 0.040999f
C248 source.n45 a_n2224_n3288# 0.017856f
C249 source.n46 a_n2224_n3288# 0.017346f
C250 source.n47 a_n2224_n3288# 0.03228f
C251 source.n48 a_n2224_n3288# 0.03228f
C252 source.n49 a_n2224_n3288# 0.017346f
C253 source.n50 a_n2224_n3288# 0.018366f
C254 source.n51 a_n2224_n3288# 0.040999f
C255 source.n52 a_n2224_n3288# 0.040999f
C256 source.n53 a_n2224_n3288# 0.018366f
C257 source.n54 a_n2224_n3288# 0.017346f
C258 source.n55 a_n2224_n3288# 0.03228f
C259 source.n56 a_n2224_n3288# 0.03228f
C260 source.n57 a_n2224_n3288# 0.017346f
C261 source.n58 a_n2224_n3288# 0.018366f
C262 source.n59 a_n2224_n3288# 0.040999f
C263 source.n60 a_n2224_n3288# 0.084134f
C264 source.n61 a_n2224_n3288# 0.018366f
C265 source.n62 a_n2224_n3288# 0.017346f
C266 source.n63 a_n2224_n3288# 0.069321f
C267 source.n64 a_n2224_n3288# 0.046433f
C268 source.n65 a_n2224_n3288# 1.29174f
C269 source.t47 a_n2224_n3288# 0.3061f
C270 source.t43 a_n2224_n3288# 0.3061f
C271 source.n66 a_n2224_n3288# 2.62084f
C272 source.n67 a_n2224_n3288# 0.43403f
C273 source.t36 a_n2224_n3288# 0.3061f
C274 source.t37 a_n2224_n3288# 0.3061f
C275 source.n68 a_n2224_n3288# 2.62084f
C276 source.n69 a_n2224_n3288# 0.43403f
C277 source.t35 a_n2224_n3288# 0.3061f
C278 source.t27 a_n2224_n3288# 0.3061f
C279 source.n70 a_n2224_n3288# 2.62084f
C280 source.n71 a_n2224_n3288# 0.43403f
C281 source.t31 a_n2224_n3288# 0.3061f
C282 source.t29 a_n2224_n3288# 0.3061f
C283 source.n72 a_n2224_n3288# 2.62084f
C284 source.n73 a_n2224_n3288# 0.43403f
C285 source.t39 a_n2224_n3288# 0.3061f
C286 source.t42 a_n2224_n3288# 0.3061f
C287 source.n74 a_n2224_n3288# 2.62084f
C288 source.n75 a_n2224_n3288# 0.43403f
C289 source.n76 a_n2224_n3288# 0.042758f
C290 source.n77 a_n2224_n3288# 0.03228f
C291 source.n78 a_n2224_n3288# 0.017346f
C292 source.n79 a_n2224_n3288# 0.040999f
C293 source.n80 a_n2224_n3288# 0.018366f
C294 source.n81 a_n2224_n3288# 0.03228f
C295 source.n82 a_n2224_n3288# 0.017346f
C296 source.n83 a_n2224_n3288# 0.040999f
C297 source.n84 a_n2224_n3288# 0.018366f
C298 source.n85 a_n2224_n3288# 0.03228f
C299 source.n86 a_n2224_n3288# 0.017856f
C300 source.n87 a_n2224_n3288# 0.040999f
C301 source.n88 a_n2224_n3288# 0.017346f
C302 source.n89 a_n2224_n3288# 0.018366f
C303 source.n90 a_n2224_n3288# 0.03228f
C304 source.n91 a_n2224_n3288# 0.017346f
C305 source.n92 a_n2224_n3288# 0.040999f
C306 source.n93 a_n2224_n3288# 0.018366f
C307 source.n94 a_n2224_n3288# 0.03228f
C308 source.n95 a_n2224_n3288# 0.017346f
C309 source.n96 a_n2224_n3288# 0.030749f
C310 source.n97 a_n2224_n3288# 0.028983f
C311 source.t45 a_n2224_n3288# 0.069244f
C312 source.n98 a_n2224_n3288# 0.232733f
C313 source.n99 a_n2224_n3288# 1.62845f
C314 source.n100 a_n2224_n3288# 0.017346f
C315 source.n101 a_n2224_n3288# 0.018366f
C316 source.n102 a_n2224_n3288# 0.040999f
C317 source.n103 a_n2224_n3288# 0.040999f
C318 source.n104 a_n2224_n3288# 0.018366f
C319 source.n105 a_n2224_n3288# 0.017346f
C320 source.n106 a_n2224_n3288# 0.03228f
C321 source.n107 a_n2224_n3288# 0.03228f
C322 source.n108 a_n2224_n3288# 0.017346f
C323 source.n109 a_n2224_n3288# 0.018366f
C324 source.n110 a_n2224_n3288# 0.040999f
C325 source.n111 a_n2224_n3288# 0.040999f
C326 source.n112 a_n2224_n3288# 0.018366f
C327 source.n113 a_n2224_n3288# 0.017346f
C328 source.n114 a_n2224_n3288# 0.03228f
C329 source.n115 a_n2224_n3288# 0.03228f
C330 source.n116 a_n2224_n3288# 0.017346f
C331 source.n117 a_n2224_n3288# 0.018366f
C332 source.n118 a_n2224_n3288# 0.040999f
C333 source.n119 a_n2224_n3288# 0.040999f
C334 source.n120 a_n2224_n3288# 0.040999f
C335 source.n121 a_n2224_n3288# 0.017856f
C336 source.n122 a_n2224_n3288# 0.017346f
C337 source.n123 a_n2224_n3288# 0.03228f
C338 source.n124 a_n2224_n3288# 0.03228f
C339 source.n125 a_n2224_n3288# 0.017346f
C340 source.n126 a_n2224_n3288# 0.018366f
C341 source.n127 a_n2224_n3288# 0.040999f
C342 source.n128 a_n2224_n3288# 0.040999f
C343 source.n129 a_n2224_n3288# 0.018366f
C344 source.n130 a_n2224_n3288# 0.017346f
C345 source.n131 a_n2224_n3288# 0.03228f
C346 source.n132 a_n2224_n3288# 0.03228f
C347 source.n133 a_n2224_n3288# 0.017346f
C348 source.n134 a_n2224_n3288# 0.018366f
C349 source.n135 a_n2224_n3288# 0.040999f
C350 source.n136 a_n2224_n3288# 0.084134f
C351 source.n137 a_n2224_n3288# 0.018366f
C352 source.n138 a_n2224_n3288# 0.017346f
C353 source.n139 a_n2224_n3288# 0.069321f
C354 source.n140 a_n2224_n3288# 0.046433f
C355 source.n141 a_n2224_n3288# 0.125462f
C356 source.n142 a_n2224_n3288# 0.042758f
C357 source.n143 a_n2224_n3288# 0.03228f
C358 source.n144 a_n2224_n3288# 0.017346f
C359 source.n145 a_n2224_n3288# 0.040999f
C360 source.n146 a_n2224_n3288# 0.018366f
C361 source.n147 a_n2224_n3288# 0.03228f
C362 source.n148 a_n2224_n3288# 0.017346f
C363 source.n149 a_n2224_n3288# 0.040999f
C364 source.n150 a_n2224_n3288# 0.018366f
C365 source.n151 a_n2224_n3288# 0.03228f
C366 source.n152 a_n2224_n3288# 0.017856f
C367 source.n153 a_n2224_n3288# 0.040999f
C368 source.n154 a_n2224_n3288# 0.017346f
C369 source.n155 a_n2224_n3288# 0.018366f
C370 source.n156 a_n2224_n3288# 0.03228f
C371 source.n157 a_n2224_n3288# 0.017346f
C372 source.n158 a_n2224_n3288# 0.040999f
C373 source.n159 a_n2224_n3288# 0.018366f
C374 source.n160 a_n2224_n3288# 0.03228f
C375 source.n161 a_n2224_n3288# 0.017346f
C376 source.n162 a_n2224_n3288# 0.030749f
C377 source.n163 a_n2224_n3288# 0.028983f
C378 source.t23 a_n2224_n3288# 0.069244f
C379 source.n164 a_n2224_n3288# 0.232733f
C380 source.n165 a_n2224_n3288# 1.62845f
C381 source.n166 a_n2224_n3288# 0.017346f
C382 source.n167 a_n2224_n3288# 0.018366f
C383 source.n168 a_n2224_n3288# 0.040999f
C384 source.n169 a_n2224_n3288# 0.040999f
C385 source.n170 a_n2224_n3288# 0.018366f
C386 source.n171 a_n2224_n3288# 0.017346f
C387 source.n172 a_n2224_n3288# 0.03228f
C388 source.n173 a_n2224_n3288# 0.03228f
C389 source.n174 a_n2224_n3288# 0.017346f
C390 source.n175 a_n2224_n3288# 0.018366f
C391 source.n176 a_n2224_n3288# 0.040999f
C392 source.n177 a_n2224_n3288# 0.040999f
C393 source.n178 a_n2224_n3288# 0.018366f
C394 source.n179 a_n2224_n3288# 0.017346f
C395 source.n180 a_n2224_n3288# 0.03228f
C396 source.n181 a_n2224_n3288# 0.03228f
C397 source.n182 a_n2224_n3288# 0.017346f
C398 source.n183 a_n2224_n3288# 0.018366f
C399 source.n184 a_n2224_n3288# 0.040999f
C400 source.n185 a_n2224_n3288# 0.040999f
C401 source.n186 a_n2224_n3288# 0.040999f
C402 source.n187 a_n2224_n3288# 0.017856f
C403 source.n188 a_n2224_n3288# 0.017346f
C404 source.n189 a_n2224_n3288# 0.03228f
C405 source.n190 a_n2224_n3288# 0.03228f
C406 source.n191 a_n2224_n3288# 0.017346f
C407 source.n192 a_n2224_n3288# 0.018366f
C408 source.n193 a_n2224_n3288# 0.040999f
C409 source.n194 a_n2224_n3288# 0.040999f
C410 source.n195 a_n2224_n3288# 0.018366f
C411 source.n196 a_n2224_n3288# 0.017346f
C412 source.n197 a_n2224_n3288# 0.03228f
C413 source.n198 a_n2224_n3288# 0.03228f
C414 source.n199 a_n2224_n3288# 0.017346f
C415 source.n200 a_n2224_n3288# 0.018366f
C416 source.n201 a_n2224_n3288# 0.040999f
C417 source.n202 a_n2224_n3288# 0.084134f
C418 source.n203 a_n2224_n3288# 0.018366f
C419 source.n204 a_n2224_n3288# 0.017346f
C420 source.n205 a_n2224_n3288# 0.069321f
C421 source.n206 a_n2224_n3288# 0.046433f
C422 source.n207 a_n2224_n3288# 0.125462f
C423 source.t20 a_n2224_n3288# 0.3061f
C424 source.t15 a_n2224_n3288# 0.3061f
C425 source.n208 a_n2224_n3288# 2.62084f
C426 source.n209 a_n2224_n3288# 0.43403f
C427 source.t10 a_n2224_n3288# 0.3061f
C428 source.t11 a_n2224_n3288# 0.3061f
C429 source.n210 a_n2224_n3288# 2.62084f
C430 source.n211 a_n2224_n3288# 0.43403f
C431 source.t13 a_n2224_n3288# 0.3061f
C432 source.t12 a_n2224_n3288# 0.3061f
C433 source.n212 a_n2224_n3288# 2.62084f
C434 source.n213 a_n2224_n3288# 0.43403f
C435 source.t5 a_n2224_n3288# 0.3061f
C436 source.t21 a_n2224_n3288# 0.3061f
C437 source.n214 a_n2224_n3288# 2.62084f
C438 source.n215 a_n2224_n3288# 0.43403f
C439 source.t0 a_n2224_n3288# 0.3061f
C440 source.t17 a_n2224_n3288# 0.3061f
C441 source.n216 a_n2224_n3288# 2.62084f
C442 source.n217 a_n2224_n3288# 0.43403f
C443 source.n218 a_n2224_n3288# 0.042758f
C444 source.n219 a_n2224_n3288# 0.03228f
C445 source.n220 a_n2224_n3288# 0.017346f
C446 source.n221 a_n2224_n3288# 0.040999f
C447 source.n222 a_n2224_n3288# 0.018366f
C448 source.n223 a_n2224_n3288# 0.03228f
C449 source.n224 a_n2224_n3288# 0.017346f
C450 source.n225 a_n2224_n3288# 0.040999f
C451 source.n226 a_n2224_n3288# 0.018366f
C452 source.n227 a_n2224_n3288# 0.03228f
C453 source.n228 a_n2224_n3288# 0.017856f
C454 source.n229 a_n2224_n3288# 0.040999f
C455 source.n230 a_n2224_n3288# 0.017346f
C456 source.n231 a_n2224_n3288# 0.018366f
C457 source.n232 a_n2224_n3288# 0.03228f
C458 source.n233 a_n2224_n3288# 0.017346f
C459 source.n234 a_n2224_n3288# 0.040999f
C460 source.n235 a_n2224_n3288# 0.018366f
C461 source.n236 a_n2224_n3288# 0.03228f
C462 source.n237 a_n2224_n3288# 0.017346f
C463 source.n238 a_n2224_n3288# 0.030749f
C464 source.n239 a_n2224_n3288# 0.028983f
C465 source.t18 a_n2224_n3288# 0.069244f
C466 source.n240 a_n2224_n3288# 0.232733f
C467 source.n241 a_n2224_n3288# 1.62845f
C468 source.n242 a_n2224_n3288# 0.017346f
C469 source.n243 a_n2224_n3288# 0.018366f
C470 source.n244 a_n2224_n3288# 0.040999f
C471 source.n245 a_n2224_n3288# 0.040999f
C472 source.n246 a_n2224_n3288# 0.018366f
C473 source.n247 a_n2224_n3288# 0.017346f
C474 source.n248 a_n2224_n3288# 0.03228f
C475 source.n249 a_n2224_n3288# 0.03228f
C476 source.n250 a_n2224_n3288# 0.017346f
C477 source.n251 a_n2224_n3288# 0.018366f
C478 source.n252 a_n2224_n3288# 0.040999f
C479 source.n253 a_n2224_n3288# 0.040999f
C480 source.n254 a_n2224_n3288# 0.018366f
C481 source.n255 a_n2224_n3288# 0.017346f
C482 source.n256 a_n2224_n3288# 0.03228f
C483 source.n257 a_n2224_n3288# 0.03228f
C484 source.n258 a_n2224_n3288# 0.017346f
C485 source.n259 a_n2224_n3288# 0.018366f
C486 source.n260 a_n2224_n3288# 0.040999f
C487 source.n261 a_n2224_n3288# 0.040999f
C488 source.n262 a_n2224_n3288# 0.040999f
C489 source.n263 a_n2224_n3288# 0.017856f
C490 source.n264 a_n2224_n3288# 0.017346f
C491 source.n265 a_n2224_n3288# 0.03228f
C492 source.n266 a_n2224_n3288# 0.03228f
C493 source.n267 a_n2224_n3288# 0.017346f
C494 source.n268 a_n2224_n3288# 0.018366f
C495 source.n269 a_n2224_n3288# 0.040999f
C496 source.n270 a_n2224_n3288# 0.040999f
C497 source.n271 a_n2224_n3288# 0.018366f
C498 source.n272 a_n2224_n3288# 0.017346f
C499 source.n273 a_n2224_n3288# 0.03228f
C500 source.n274 a_n2224_n3288# 0.03228f
C501 source.n275 a_n2224_n3288# 0.017346f
C502 source.n276 a_n2224_n3288# 0.018366f
C503 source.n277 a_n2224_n3288# 0.040999f
C504 source.n278 a_n2224_n3288# 0.084134f
C505 source.n279 a_n2224_n3288# 0.018366f
C506 source.n280 a_n2224_n3288# 0.017346f
C507 source.n281 a_n2224_n3288# 0.069321f
C508 source.n282 a_n2224_n3288# 0.046433f
C509 source.n283 a_n2224_n3288# 1.7977f
C510 source.n284 a_n2224_n3288# 0.042758f
C511 source.n285 a_n2224_n3288# 0.03228f
C512 source.n286 a_n2224_n3288# 0.017346f
C513 source.n287 a_n2224_n3288# 0.040999f
C514 source.n288 a_n2224_n3288# 0.018366f
C515 source.n289 a_n2224_n3288# 0.03228f
C516 source.n290 a_n2224_n3288# 0.017346f
C517 source.n291 a_n2224_n3288# 0.040999f
C518 source.n292 a_n2224_n3288# 0.018366f
C519 source.n293 a_n2224_n3288# 0.03228f
C520 source.n294 a_n2224_n3288# 0.017856f
C521 source.n295 a_n2224_n3288# 0.040999f
C522 source.n296 a_n2224_n3288# 0.018366f
C523 source.n297 a_n2224_n3288# 0.03228f
C524 source.n298 a_n2224_n3288# 0.017346f
C525 source.n299 a_n2224_n3288# 0.040999f
C526 source.n300 a_n2224_n3288# 0.018366f
C527 source.n301 a_n2224_n3288# 0.03228f
C528 source.n302 a_n2224_n3288# 0.017346f
C529 source.n303 a_n2224_n3288# 0.030749f
C530 source.n304 a_n2224_n3288# 0.028983f
C531 source.t40 a_n2224_n3288# 0.069244f
C532 source.n305 a_n2224_n3288# 0.232733f
C533 source.n306 a_n2224_n3288# 1.62845f
C534 source.n307 a_n2224_n3288# 0.017346f
C535 source.n308 a_n2224_n3288# 0.018366f
C536 source.n309 a_n2224_n3288# 0.040999f
C537 source.n310 a_n2224_n3288# 0.040999f
C538 source.n311 a_n2224_n3288# 0.018366f
C539 source.n312 a_n2224_n3288# 0.017346f
C540 source.n313 a_n2224_n3288# 0.03228f
C541 source.n314 a_n2224_n3288# 0.03228f
C542 source.n315 a_n2224_n3288# 0.017346f
C543 source.n316 a_n2224_n3288# 0.018366f
C544 source.n317 a_n2224_n3288# 0.040999f
C545 source.n318 a_n2224_n3288# 0.040999f
C546 source.n319 a_n2224_n3288# 0.018366f
C547 source.n320 a_n2224_n3288# 0.017346f
C548 source.n321 a_n2224_n3288# 0.03228f
C549 source.n322 a_n2224_n3288# 0.03228f
C550 source.n323 a_n2224_n3288# 0.017346f
C551 source.n324 a_n2224_n3288# 0.017346f
C552 source.n325 a_n2224_n3288# 0.018366f
C553 source.n326 a_n2224_n3288# 0.040999f
C554 source.n327 a_n2224_n3288# 0.040999f
C555 source.n328 a_n2224_n3288# 0.040999f
C556 source.n329 a_n2224_n3288# 0.017856f
C557 source.n330 a_n2224_n3288# 0.017346f
C558 source.n331 a_n2224_n3288# 0.03228f
C559 source.n332 a_n2224_n3288# 0.03228f
C560 source.n333 a_n2224_n3288# 0.017346f
C561 source.n334 a_n2224_n3288# 0.018366f
C562 source.n335 a_n2224_n3288# 0.040999f
C563 source.n336 a_n2224_n3288# 0.040999f
C564 source.n337 a_n2224_n3288# 0.018366f
C565 source.n338 a_n2224_n3288# 0.017346f
C566 source.n339 a_n2224_n3288# 0.03228f
C567 source.n340 a_n2224_n3288# 0.03228f
C568 source.n341 a_n2224_n3288# 0.017346f
C569 source.n342 a_n2224_n3288# 0.018366f
C570 source.n343 a_n2224_n3288# 0.040999f
C571 source.n344 a_n2224_n3288# 0.084134f
C572 source.n345 a_n2224_n3288# 0.018366f
C573 source.n346 a_n2224_n3288# 0.017346f
C574 source.n347 a_n2224_n3288# 0.069321f
C575 source.n348 a_n2224_n3288# 0.046433f
C576 source.n349 a_n2224_n3288# 1.7977f
C577 source.t41 a_n2224_n3288# 0.3061f
C578 source.t25 a_n2224_n3288# 0.3061f
C579 source.n350 a_n2224_n3288# 2.62082f
C580 source.n351 a_n2224_n3288# 0.434046f
C581 source.t28 a_n2224_n3288# 0.3061f
C582 source.t33 a_n2224_n3288# 0.3061f
C583 source.n352 a_n2224_n3288# 2.62082f
C584 source.n353 a_n2224_n3288# 0.434046f
C585 source.t38 a_n2224_n3288# 0.3061f
C586 source.t26 a_n2224_n3288# 0.3061f
C587 source.n354 a_n2224_n3288# 2.62082f
C588 source.n355 a_n2224_n3288# 0.434046f
C589 source.t46 a_n2224_n3288# 0.3061f
C590 source.t34 a_n2224_n3288# 0.3061f
C591 source.n356 a_n2224_n3288# 2.62082f
C592 source.n357 a_n2224_n3288# 0.434046f
C593 source.t32 a_n2224_n3288# 0.3061f
C594 source.t30 a_n2224_n3288# 0.3061f
C595 source.n358 a_n2224_n3288# 2.62082f
C596 source.n359 a_n2224_n3288# 0.434046f
C597 source.n360 a_n2224_n3288# 0.042758f
C598 source.n361 a_n2224_n3288# 0.03228f
C599 source.n362 a_n2224_n3288# 0.017346f
C600 source.n363 a_n2224_n3288# 0.040999f
C601 source.n364 a_n2224_n3288# 0.018366f
C602 source.n365 a_n2224_n3288# 0.03228f
C603 source.n366 a_n2224_n3288# 0.017346f
C604 source.n367 a_n2224_n3288# 0.040999f
C605 source.n368 a_n2224_n3288# 0.018366f
C606 source.n369 a_n2224_n3288# 0.03228f
C607 source.n370 a_n2224_n3288# 0.017856f
C608 source.n371 a_n2224_n3288# 0.040999f
C609 source.n372 a_n2224_n3288# 0.018366f
C610 source.n373 a_n2224_n3288# 0.03228f
C611 source.n374 a_n2224_n3288# 0.017346f
C612 source.n375 a_n2224_n3288# 0.040999f
C613 source.n376 a_n2224_n3288# 0.018366f
C614 source.n377 a_n2224_n3288# 0.03228f
C615 source.n378 a_n2224_n3288# 0.017346f
C616 source.n379 a_n2224_n3288# 0.030749f
C617 source.n380 a_n2224_n3288# 0.028983f
C618 source.t44 a_n2224_n3288# 0.069244f
C619 source.n381 a_n2224_n3288# 0.232733f
C620 source.n382 a_n2224_n3288# 1.62845f
C621 source.n383 a_n2224_n3288# 0.017346f
C622 source.n384 a_n2224_n3288# 0.018366f
C623 source.n385 a_n2224_n3288# 0.040999f
C624 source.n386 a_n2224_n3288# 0.040999f
C625 source.n387 a_n2224_n3288# 0.018366f
C626 source.n388 a_n2224_n3288# 0.017346f
C627 source.n389 a_n2224_n3288# 0.03228f
C628 source.n390 a_n2224_n3288# 0.03228f
C629 source.n391 a_n2224_n3288# 0.017346f
C630 source.n392 a_n2224_n3288# 0.018366f
C631 source.n393 a_n2224_n3288# 0.040999f
C632 source.n394 a_n2224_n3288# 0.040999f
C633 source.n395 a_n2224_n3288# 0.018366f
C634 source.n396 a_n2224_n3288# 0.017346f
C635 source.n397 a_n2224_n3288# 0.03228f
C636 source.n398 a_n2224_n3288# 0.03228f
C637 source.n399 a_n2224_n3288# 0.017346f
C638 source.n400 a_n2224_n3288# 0.017346f
C639 source.n401 a_n2224_n3288# 0.018366f
C640 source.n402 a_n2224_n3288# 0.040999f
C641 source.n403 a_n2224_n3288# 0.040999f
C642 source.n404 a_n2224_n3288# 0.040999f
C643 source.n405 a_n2224_n3288# 0.017856f
C644 source.n406 a_n2224_n3288# 0.017346f
C645 source.n407 a_n2224_n3288# 0.03228f
C646 source.n408 a_n2224_n3288# 0.03228f
C647 source.n409 a_n2224_n3288# 0.017346f
C648 source.n410 a_n2224_n3288# 0.018366f
C649 source.n411 a_n2224_n3288# 0.040999f
C650 source.n412 a_n2224_n3288# 0.040999f
C651 source.n413 a_n2224_n3288# 0.018366f
C652 source.n414 a_n2224_n3288# 0.017346f
C653 source.n415 a_n2224_n3288# 0.03228f
C654 source.n416 a_n2224_n3288# 0.03228f
C655 source.n417 a_n2224_n3288# 0.017346f
C656 source.n418 a_n2224_n3288# 0.018366f
C657 source.n419 a_n2224_n3288# 0.040999f
C658 source.n420 a_n2224_n3288# 0.084134f
C659 source.n421 a_n2224_n3288# 0.018366f
C660 source.n422 a_n2224_n3288# 0.017346f
C661 source.n423 a_n2224_n3288# 0.069321f
C662 source.n424 a_n2224_n3288# 0.046433f
C663 source.n425 a_n2224_n3288# 0.125462f
C664 source.n426 a_n2224_n3288# 0.042758f
C665 source.n427 a_n2224_n3288# 0.03228f
C666 source.n428 a_n2224_n3288# 0.017346f
C667 source.n429 a_n2224_n3288# 0.040999f
C668 source.n430 a_n2224_n3288# 0.018366f
C669 source.n431 a_n2224_n3288# 0.03228f
C670 source.n432 a_n2224_n3288# 0.017346f
C671 source.n433 a_n2224_n3288# 0.040999f
C672 source.n434 a_n2224_n3288# 0.018366f
C673 source.n435 a_n2224_n3288# 0.03228f
C674 source.n436 a_n2224_n3288# 0.017856f
C675 source.n437 a_n2224_n3288# 0.040999f
C676 source.n438 a_n2224_n3288# 0.018366f
C677 source.n439 a_n2224_n3288# 0.03228f
C678 source.n440 a_n2224_n3288# 0.017346f
C679 source.n441 a_n2224_n3288# 0.040999f
C680 source.n442 a_n2224_n3288# 0.018366f
C681 source.n443 a_n2224_n3288# 0.03228f
C682 source.n444 a_n2224_n3288# 0.017346f
C683 source.n445 a_n2224_n3288# 0.030749f
C684 source.n446 a_n2224_n3288# 0.028983f
C685 source.t6 a_n2224_n3288# 0.069244f
C686 source.n447 a_n2224_n3288# 0.232733f
C687 source.n448 a_n2224_n3288# 1.62845f
C688 source.n449 a_n2224_n3288# 0.017346f
C689 source.n450 a_n2224_n3288# 0.018366f
C690 source.n451 a_n2224_n3288# 0.040999f
C691 source.n452 a_n2224_n3288# 0.040999f
C692 source.n453 a_n2224_n3288# 0.018366f
C693 source.n454 a_n2224_n3288# 0.017346f
C694 source.n455 a_n2224_n3288# 0.03228f
C695 source.n456 a_n2224_n3288# 0.03228f
C696 source.n457 a_n2224_n3288# 0.017346f
C697 source.n458 a_n2224_n3288# 0.018366f
C698 source.n459 a_n2224_n3288# 0.040999f
C699 source.n460 a_n2224_n3288# 0.040999f
C700 source.n461 a_n2224_n3288# 0.018366f
C701 source.n462 a_n2224_n3288# 0.017346f
C702 source.n463 a_n2224_n3288# 0.03228f
C703 source.n464 a_n2224_n3288# 0.03228f
C704 source.n465 a_n2224_n3288# 0.017346f
C705 source.n466 a_n2224_n3288# 0.017346f
C706 source.n467 a_n2224_n3288# 0.018366f
C707 source.n468 a_n2224_n3288# 0.040999f
C708 source.n469 a_n2224_n3288# 0.040999f
C709 source.n470 a_n2224_n3288# 0.040999f
C710 source.n471 a_n2224_n3288# 0.017856f
C711 source.n472 a_n2224_n3288# 0.017346f
C712 source.n473 a_n2224_n3288# 0.03228f
C713 source.n474 a_n2224_n3288# 0.03228f
C714 source.n475 a_n2224_n3288# 0.017346f
C715 source.n476 a_n2224_n3288# 0.018366f
C716 source.n477 a_n2224_n3288# 0.040999f
C717 source.n478 a_n2224_n3288# 0.040999f
C718 source.n479 a_n2224_n3288# 0.018366f
C719 source.n480 a_n2224_n3288# 0.017346f
C720 source.n481 a_n2224_n3288# 0.03228f
C721 source.n482 a_n2224_n3288# 0.03228f
C722 source.n483 a_n2224_n3288# 0.017346f
C723 source.n484 a_n2224_n3288# 0.018366f
C724 source.n485 a_n2224_n3288# 0.040999f
C725 source.n486 a_n2224_n3288# 0.084134f
C726 source.n487 a_n2224_n3288# 0.018366f
C727 source.n488 a_n2224_n3288# 0.017346f
C728 source.n489 a_n2224_n3288# 0.069321f
C729 source.n490 a_n2224_n3288# 0.046433f
C730 source.n491 a_n2224_n3288# 0.125462f
C731 source.t1 a_n2224_n3288# 0.3061f
C732 source.t22 a_n2224_n3288# 0.3061f
C733 source.n492 a_n2224_n3288# 2.62082f
C734 source.n493 a_n2224_n3288# 0.434046f
C735 source.t16 a_n2224_n3288# 0.3061f
C736 source.t2 a_n2224_n3288# 0.3061f
C737 source.n494 a_n2224_n3288# 2.62082f
C738 source.n495 a_n2224_n3288# 0.434046f
C739 source.t3 a_n2224_n3288# 0.3061f
C740 source.t19 a_n2224_n3288# 0.3061f
C741 source.n496 a_n2224_n3288# 2.62082f
C742 source.n497 a_n2224_n3288# 0.434046f
C743 source.t14 a_n2224_n3288# 0.3061f
C744 source.t9 a_n2224_n3288# 0.3061f
C745 source.n498 a_n2224_n3288# 2.62082f
C746 source.n499 a_n2224_n3288# 0.434046f
C747 source.t7 a_n2224_n3288# 0.3061f
C748 source.t4 a_n2224_n3288# 0.3061f
C749 source.n500 a_n2224_n3288# 2.62082f
C750 source.n501 a_n2224_n3288# 0.434046f
C751 source.n502 a_n2224_n3288# 0.042758f
C752 source.n503 a_n2224_n3288# 0.03228f
C753 source.n504 a_n2224_n3288# 0.017346f
C754 source.n505 a_n2224_n3288# 0.040999f
C755 source.n506 a_n2224_n3288# 0.018366f
C756 source.n507 a_n2224_n3288# 0.03228f
C757 source.n508 a_n2224_n3288# 0.017346f
C758 source.n509 a_n2224_n3288# 0.040999f
C759 source.n510 a_n2224_n3288# 0.018366f
C760 source.n511 a_n2224_n3288# 0.03228f
C761 source.n512 a_n2224_n3288# 0.017856f
C762 source.n513 a_n2224_n3288# 0.040999f
C763 source.n514 a_n2224_n3288# 0.018366f
C764 source.n515 a_n2224_n3288# 0.03228f
C765 source.n516 a_n2224_n3288# 0.017346f
C766 source.n517 a_n2224_n3288# 0.040999f
C767 source.n518 a_n2224_n3288# 0.018366f
C768 source.n519 a_n2224_n3288# 0.03228f
C769 source.n520 a_n2224_n3288# 0.017346f
C770 source.n521 a_n2224_n3288# 0.030749f
C771 source.n522 a_n2224_n3288# 0.028983f
C772 source.t8 a_n2224_n3288# 0.069244f
C773 source.n523 a_n2224_n3288# 0.232733f
C774 source.n524 a_n2224_n3288# 1.62845f
C775 source.n525 a_n2224_n3288# 0.017346f
C776 source.n526 a_n2224_n3288# 0.018366f
C777 source.n527 a_n2224_n3288# 0.040999f
C778 source.n528 a_n2224_n3288# 0.040999f
C779 source.n529 a_n2224_n3288# 0.018366f
C780 source.n530 a_n2224_n3288# 0.017346f
C781 source.n531 a_n2224_n3288# 0.03228f
C782 source.n532 a_n2224_n3288# 0.03228f
C783 source.n533 a_n2224_n3288# 0.017346f
C784 source.n534 a_n2224_n3288# 0.018366f
C785 source.n535 a_n2224_n3288# 0.040999f
C786 source.n536 a_n2224_n3288# 0.040999f
C787 source.n537 a_n2224_n3288# 0.018366f
C788 source.n538 a_n2224_n3288# 0.017346f
C789 source.n539 a_n2224_n3288# 0.03228f
C790 source.n540 a_n2224_n3288# 0.03228f
C791 source.n541 a_n2224_n3288# 0.017346f
C792 source.n542 a_n2224_n3288# 0.017346f
C793 source.n543 a_n2224_n3288# 0.018366f
C794 source.n544 a_n2224_n3288# 0.040999f
C795 source.n545 a_n2224_n3288# 0.040999f
C796 source.n546 a_n2224_n3288# 0.040999f
C797 source.n547 a_n2224_n3288# 0.017856f
C798 source.n548 a_n2224_n3288# 0.017346f
C799 source.n549 a_n2224_n3288# 0.03228f
C800 source.n550 a_n2224_n3288# 0.03228f
C801 source.n551 a_n2224_n3288# 0.017346f
C802 source.n552 a_n2224_n3288# 0.018366f
C803 source.n553 a_n2224_n3288# 0.040999f
C804 source.n554 a_n2224_n3288# 0.040999f
C805 source.n555 a_n2224_n3288# 0.018366f
C806 source.n556 a_n2224_n3288# 0.017346f
C807 source.n557 a_n2224_n3288# 0.03228f
C808 source.n558 a_n2224_n3288# 0.03228f
C809 source.n559 a_n2224_n3288# 0.017346f
C810 source.n560 a_n2224_n3288# 0.018366f
C811 source.n561 a_n2224_n3288# 0.040999f
C812 source.n562 a_n2224_n3288# 0.084134f
C813 source.n563 a_n2224_n3288# 0.018366f
C814 source.n564 a_n2224_n3288# 0.017346f
C815 source.n565 a_n2224_n3288# 0.069321f
C816 source.n566 a_n2224_n3288# 0.046433f
C817 source.n567 a_n2224_n3288# 0.304092f
C818 source.n568 a_n2224_n3288# 2.02253f
C819 plus.n0 a_n2224_n3288# 0.050673f
C820 plus.t14 a_n2224_n3288# 0.429579f
C821 plus.t3 a_n2224_n3288# 0.429579f
C822 plus.n1 a_n2224_n3288# 0.018372f
C823 plus.n2 a_n2224_n3288# 0.050673f
C824 plus.t4 a_n2224_n3288# 0.429579f
C825 plus.t10 a_n2224_n3288# 0.429579f
C826 plus.t22 a_n2224_n3288# 0.429579f
C827 plus.n3 a_n2224_n3288# 0.173015f
C828 plus.n4 a_n2224_n3288# 0.050673f
C829 plus.t11 a_n2224_n3288# 0.429579f
C830 plus.t0 a_n2224_n3288# 0.429579f
C831 plus.n5 a_n2224_n3288# 0.017747f
C832 plus.t6 a_n2224_n3288# 0.433205f
C833 plus.n6 a_n2224_n3288# 0.186888f
C834 plus.t1 a_n2224_n3288# 0.429579f
C835 plus.n7 a_n2224_n3288# 0.173015f
C836 plus.t12 a_n2224_n3288# 0.429579f
C837 plus.n8 a_n2224_n3288# 0.173015f
C838 plus.n9 a_n2224_n3288# 0.019309f
C839 plus.n10 a_n2224_n3288# 0.105343f
C840 plus.n11 a_n2224_n3288# 0.050673f
C841 plus.n12 a_n2224_n3288# 0.050673f
C842 plus.n13 a_n2224_n3288# 0.018372f
C843 plus.n14 a_n2224_n3288# 0.173015f
C844 plus.n15 a_n2224_n3288# 0.019309f
C845 plus.n16 a_n2224_n3288# 0.173015f
C846 plus.n17 a_n2224_n3288# 0.019309f
C847 plus.n18 a_n2224_n3288# 0.050673f
C848 plus.n19 a_n2224_n3288# 0.050673f
C849 plus.n20 a_n2224_n3288# 0.019309f
C850 plus.n21 a_n2224_n3288# 0.173015f
C851 plus.n22 a_n2224_n3288# 0.019309f
C852 plus.n23 a_n2224_n3288# 0.173015f
C853 plus.t16 a_n2224_n3288# 0.429579f
C854 plus.n24 a_n2224_n3288# 0.173015f
C855 plus.n25 a_n2224_n3288# 0.019309f
C856 plus.n26 a_n2224_n3288# 0.050673f
C857 plus.n27 a_n2224_n3288# 0.050673f
C858 plus.n28 a_n2224_n3288# 0.050673f
C859 plus.n29 a_n2224_n3288# 0.017747f
C860 plus.n30 a_n2224_n3288# 0.173015f
C861 plus.n31 a_n2224_n3288# 0.019309f
C862 plus.n32 a_n2224_n3288# 0.173015f
C863 plus.t2 a_n2224_n3288# 0.433205f
C864 plus.n33 a_n2224_n3288# 0.186824f
C865 plus.n34 a_n2224_n3288# 0.558739f
C866 plus.n35 a_n2224_n3288# 0.050673f
C867 plus.t9 a_n2224_n3288# 0.433205f
C868 plus.t13 a_n2224_n3288# 0.429579f
C869 plus.t15 a_n2224_n3288# 0.429579f
C870 plus.n36 a_n2224_n3288# 0.018372f
C871 plus.n37 a_n2224_n3288# 0.050673f
C872 plus.t19 a_n2224_n3288# 0.429579f
C873 plus.n38 a_n2224_n3288# 0.173015f
C874 plus.t7 a_n2224_n3288# 0.429579f
C875 plus.t17 a_n2224_n3288# 0.429579f
C876 plus.t20 a_n2224_n3288# 0.429579f
C877 plus.n39 a_n2224_n3288# 0.173015f
C878 plus.n40 a_n2224_n3288# 0.050673f
C879 plus.t5 a_n2224_n3288# 0.429579f
C880 plus.t23 a_n2224_n3288# 0.429579f
C881 plus.n41 a_n2224_n3288# 0.017747f
C882 plus.t21 a_n2224_n3288# 0.433205f
C883 plus.n42 a_n2224_n3288# 0.186888f
C884 plus.t8 a_n2224_n3288# 0.429579f
C885 plus.n43 a_n2224_n3288# 0.173015f
C886 plus.t18 a_n2224_n3288# 0.429579f
C887 plus.n44 a_n2224_n3288# 0.173015f
C888 plus.n45 a_n2224_n3288# 0.019309f
C889 plus.n46 a_n2224_n3288# 0.105343f
C890 plus.n47 a_n2224_n3288# 0.050673f
C891 plus.n48 a_n2224_n3288# 0.050673f
C892 plus.n49 a_n2224_n3288# 0.018372f
C893 plus.n50 a_n2224_n3288# 0.173015f
C894 plus.n51 a_n2224_n3288# 0.019309f
C895 plus.n52 a_n2224_n3288# 0.173015f
C896 plus.n53 a_n2224_n3288# 0.019309f
C897 plus.n54 a_n2224_n3288# 0.050673f
C898 plus.n55 a_n2224_n3288# 0.050673f
C899 plus.n56 a_n2224_n3288# 0.019309f
C900 plus.n57 a_n2224_n3288# 0.173015f
C901 plus.n58 a_n2224_n3288# 0.019309f
C902 plus.n59 a_n2224_n3288# 0.173015f
C903 plus.n60 a_n2224_n3288# 0.019309f
C904 plus.n61 a_n2224_n3288# 0.050673f
C905 plus.n62 a_n2224_n3288# 0.050673f
C906 plus.n63 a_n2224_n3288# 0.050673f
C907 plus.n64 a_n2224_n3288# 0.017747f
C908 plus.n65 a_n2224_n3288# 0.173015f
C909 plus.n66 a_n2224_n3288# 0.019309f
C910 plus.n67 a_n2224_n3288# 0.173015f
C911 plus.n68 a_n2224_n3288# 0.186824f
C912 plus.n69 a_n2224_n3288# 1.60047f
.ends

