* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t35 minus.t0 drain_right.t7 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X1 drain_right.t13 minus.t1 source.t34 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X2 drain_right.t5 minus.t2 source.t33 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X3 drain_right.t19 minus.t3 source.t32 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X4 source.t1 plus.t0 drain_left.t19 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X5 source.t31 minus.t4 drain_right.t17 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X6 drain_left.t18 plus.t1 source.t0 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X7 source.t9 plus.t2 drain_left.t17 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X8 drain_left.t16 plus.t3 source.t15 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X9 a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.2
X10 source.t30 minus.t5 drain_right.t4 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X11 source.t29 minus.t6 drain_right.t18 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X12 source.t28 minus.t7 drain_right.t0 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X13 drain_left.t15 plus.t4 source.t8 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X14 drain_right.t16 minus.t8 source.t27 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X15 source.t14 plus.t5 drain_left.t14 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X16 source.t26 minus.t9 drain_right.t12 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X17 a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X18 drain_left.t13 plus.t6 source.t7 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X19 source.t6 plus.t7 drain_left.t12 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X20 source.t25 minus.t10 drain_right.t6 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X21 drain_left.t11 plus.t8 source.t5 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X22 drain_right.t3 minus.t11 source.t24 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X23 drain_right.t1 minus.t12 source.t23 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X24 drain_left.t10 plus.t9 source.t13 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X25 drain_right.t2 minus.t13 source.t22 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X26 drain_right.t10 minus.t14 source.t21 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X27 drain_left.t9 plus.t10 source.t11 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X28 source.t20 minus.t15 drain_right.t8 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X29 source.t10 plus.t11 drain_left.t8 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X30 a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X31 drain_right.t14 minus.t16 source.t19 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X32 source.t12 plus.t12 drain_left.t7 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X33 source.t4 plus.t13 drain_left.t6 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X34 drain_left.t5 plus.t14 source.t3 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X35 source.t2 plus.t15 drain_left.t4 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X36 source.t37 plus.t16 drain_left.t3 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X37 drain_right.t11 minus.t17 source.t18 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X38 source.t17 minus.t18 drain_right.t9 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X39 source.t16 minus.t19 drain_right.t15 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X40 drain_left.t2 plus.t17 source.t39 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X41 drain_left.t1 plus.t18 source.t38 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X42 source.t36 plus.t19 drain_left.t0 a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X43 a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# a_n1882_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
R0 minus.n23 minus.t9 333.384
R1 minus.n5 minus.t13 333.384
R2 minus.n48 minus.t12 333.384
R3 minus.n30 minus.t10 333.384
R4 minus.n22 minus.t11 277.151
R5 minus.n20 minus.t19 277.151
R6 minus.n1 minus.t2 277.151
R7 minus.n15 minus.t5 277.151
R8 minus.n13 minus.t14 277.151
R9 minus.n3 minus.t18 277.151
R10 minus.n8 minus.t1 277.151
R11 minus.n6 minus.t7 277.151
R12 minus.n47 minus.t0 277.151
R13 minus.n45 minus.t17 277.151
R14 minus.n26 minus.t6 277.151
R15 minus.n40 minus.t3 277.151
R16 minus.n38 minus.t15 277.151
R17 minus.n28 minus.t8 277.151
R18 minus.n33 minus.t4 277.151
R19 minus.n31 minus.t16 277.151
R20 minus.n5 minus.n4 161.489
R21 minus.n30 minus.n29 161.489
R22 minus.n24 minus.n23 161.3
R23 minus.n21 minus.n0 161.3
R24 minus.n19 minus.n18 161.3
R25 minus.n17 minus.n16 161.3
R26 minus.n14 minus.n2 161.3
R27 minus.n12 minus.n11 161.3
R28 minus.n10 minus.n9 161.3
R29 minus.n7 minus.n4 161.3
R30 minus.n49 minus.n48 161.3
R31 minus.n46 minus.n25 161.3
R32 minus.n44 minus.n43 161.3
R33 minus.n42 minus.n41 161.3
R34 minus.n39 minus.n27 161.3
R35 minus.n37 minus.n36 161.3
R36 minus.n35 minus.n34 161.3
R37 minus.n32 minus.n29 161.3
R38 minus.n22 minus.n21 51.852
R39 minus.n7 minus.n6 51.852
R40 minus.n32 minus.n31 51.852
R41 minus.n47 minus.n46 51.852
R42 minus.n20 minus.n19 47.4702
R43 minus.n9 minus.n8 47.4702
R44 minus.n34 minus.n33 47.4702
R45 minus.n45 minus.n44 47.4702
R46 minus.n16 minus.n1 43.0884
R47 minus.n12 minus.n3 43.0884
R48 minus.n37 minus.n28 43.0884
R49 minus.n41 minus.n26 43.0884
R50 minus.n15 minus.n14 38.7066
R51 minus.n14 minus.n13 38.7066
R52 minus.n39 minus.n38 38.7066
R53 minus.n40 minus.n39 38.7066
R54 minus.n16 minus.n15 34.3247
R55 minus.n13 minus.n12 34.3247
R56 minus.n38 minus.n37 34.3247
R57 minus.n41 minus.n40 34.3247
R58 minus.n19 minus.n1 29.9429
R59 minus.n9 minus.n3 29.9429
R60 minus.n34 minus.n28 29.9429
R61 minus.n44 minus.n26 29.9429
R62 minus.n50 minus.n24 27.8944
R63 minus.n21 minus.n20 25.5611
R64 minus.n8 minus.n7 25.5611
R65 minus.n33 minus.n32 25.5611
R66 minus.n46 minus.n45 25.5611
R67 minus.n23 minus.n22 21.1793
R68 minus.n6 minus.n5 21.1793
R69 minus.n31 minus.n30 21.1793
R70 minus.n48 minus.n47 21.1793
R71 minus.n50 minus.n49 6.47777
R72 minus.n24 minus.n0 0.189894
R73 minus.n18 minus.n0 0.189894
R74 minus.n18 minus.n17 0.189894
R75 minus.n17 minus.n2 0.189894
R76 minus.n11 minus.n2 0.189894
R77 minus.n11 minus.n10 0.189894
R78 minus.n10 minus.n4 0.189894
R79 minus.n35 minus.n29 0.189894
R80 minus.n36 minus.n35 0.189894
R81 minus.n36 minus.n27 0.189894
R82 minus.n42 minus.n27 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n25 0.189894
R85 minus.n49 minus.n25 0.189894
R86 minus minus.n50 0.188
R87 drain_right.n10 drain_right.n8 240.589
R88 drain_right.n6 drain_right.n4 240.589
R89 drain_right.n2 drain_right.n0 240.589
R90 drain_right.n10 drain_right.n9 240.132
R91 drain_right.n12 drain_right.n11 240.132
R92 drain_right.n14 drain_right.n13 240.132
R93 drain_right.n16 drain_right.n15 240.132
R94 drain_right.n7 drain_right.n3 240.131
R95 drain_right.n6 drain_right.n5 240.131
R96 drain_right.n2 drain_right.n1 240.131
R97 drain_right drain_right.n7 22.1357
R98 drain_right.n3 drain_right.t8 19.8005
R99 drain_right.n3 drain_right.t19 19.8005
R100 drain_right.n4 drain_right.t7 19.8005
R101 drain_right.n4 drain_right.t1 19.8005
R102 drain_right.n5 drain_right.t18 19.8005
R103 drain_right.n5 drain_right.t11 19.8005
R104 drain_right.n1 drain_right.t17 19.8005
R105 drain_right.n1 drain_right.t16 19.8005
R106 drain_right.n0 drain_right.t6 19.8005
R107 drain_right.n0 drain_right.t14 19.8005
R108 drain_right.n8 drain_right.t0 19.8005
R109 drain_right.n8 drain_right.t2 19.8005
R110 drain_right.n9 drain_right.t9 19.8005
R111 drain_right.n9 drain_right.t13 19.8005
R112 drain_right.n11 drain_right.t4 19.8005
R113 drain_right.n11 drain_right.t10 19.8005
R114 drain_right.n13 drain_right.t15 19.8005
R115 drain_right.n13 drain_right.t5 19.8005
R116 drain_right.n15 drain_right.t12 19.8005
R117 drain_right.n15 drain_right.t3 19.8005
R118 drain_right drain_right.n16 6.11011
R119 drain_right.n16 drain_right.n14 0.457397
R120 drain_right.n14 drain_right.n12 0.457397
R121 drain_right.n12 drain_right.n10 0.457397
R122 drain_right.n7 drain_right.n6 0.402051
R123 drain_right.n7 drain_right.n2 0.402051
R124 source.n0 source.t8 243.255
R125 source.n9 source.t6 243.255
R126 source.n10 source.t22 243.255
R127 source.n19 source.t26 243.255
R128 source.n39 source.t23 243.254
R129 source.n30 source.t25 243.254
R130 source.n29 source.t5 243.254
R131 source.n20 source.t37 243.254
R132 source.n2 source.n1 223.454
R133 source.n4 source.n3 223.454
R134 source.n6 source.n5 223.454
R135 source.n8 source.n7 223.454
R136 source.n12 source.n11 223.454
R137 source.n14 source.n13 223.454
R138 source.n16 source.n15 223.454
R139 source.n18 source.n17 223.454
R140 source.n38 source.n37 223.453
R141 source.n36 source.n35 223.453
R142 source.n34 source.n33 223.453
R143 source.n32 source.n31 223.453
R144 source.n28 source.n27 223.453
R145 source.n26 source.n25 223.453
R146 source.n24 source.n23 223.453
R147 source.n22 source.n21 223.453
R148 source.n37 source.t18 19.8005
R149 source.n37 source.t35 19.8005
R150 source.n35 source.t32 19.8005
R151 source.n35 source.t29 19.8005
R152 source.n33 source.t27 19.8005
R153 source.n33 source.t20 19.8005
R154 source.n31 source.t19 19.8005
R155 source.n31 source.t31 19.8005
R156 source.n27 source.t0 19.8005
R157 source.n27 source.t2 19.8005
R158 source.n25 source.t39 19.8005
R159 source.n25 source.t12 19.8005
R160 source.n23 source.t11 19.8005
R161 source.n23 source.t14 19.8005
R162 source.n21 source.t13 19.8005
R163 source.n21 source.t1 19.8005
R164 source.n1 source.t38 19.8005
R165 source.n1 source.t10 19.8005
R166 source.n3 source.t7 19.8005
R167 source.n3 source.t9 19.8005
R168 source.n5 source.t3 19.8005
R169 source.n5 source.t4 19.8005
R170 source.n7 source.t15 19.8005
R171 source.n7 source.t36 19.8005
R172 source.n11 source.t34 19.8005
R173 source.n11 source.t28 19.8005
R174 source.n13 source.t21 19.8005
R175 source.n13 source.t17 19.8005
R176 source.n15 source.t33 19.8005
R177 source.n15 source.t30 19.8005
R178 source.n17 source.t24 19.8005
R179 source.n17 source.t16 19.8005
R180 source.n20 source.n19 13.4113
R181 source.n40 source.n0 7.91991
R182 source.n40 source.n39 5.49188
R183 source.n10 source.n9 0.470328
R184 source.n30 source.n29 0.470328
R185 source.n19 source.n18 0.457397
R186 source.n18 source.n16 0.457397
R187 source.n16 source.n14 0.457397
R188 source.n14 source.n12 0.457397
R189 source.n12 source.n10 0.457397
R190 source.n9 source.n8 0.457397
R191 source.n8 source.n6 0.457397
R192 source.n6 source.n4 0.457397
R193 source.n4 source.n2 0.457397
R194 source.n2 source.n0 0.457397
R195 source.n22 source.n20 0.457397
R196 source.n24 source.n22 0.457397
R197 source.n26 source.n24 0.457397
R198 source.n28 source.n26 0.457397
R199 source.n29 source.n28 0.457397
R200 source.n32 source.n30 0.457397
R201 source.n34 source.n32 0.457397
R202 source.n36 source.n34 0.457397
R203 source.n38 source.n36 0.457397
R204 source.n39 source.n38 0.457397
R205 source source.n40 0.188
R206 plus.n5 plus.t7 333.384
R207 plus.n23 plus.t4 333.384
R208 plus.n30 plus.t8 333.384
R209 plus.n48 plus.t16 333.384
R210 plus.n6 plus.t3 277.151
R211 plus.n8 plus.t19 277.151
R212 plus.n3 plus.t14 277.151
R213 plus.n13 plus.t13 277.151
R214 plus.n15 plus.t6 277.151
R215 plus.n1 plus.t2 277.151
R216 plus.n20 plus.t18 277.151
R217 plus.n22 plus.t11 277.151
R218 plus.n31 plus.t15 277.151
R219 plus.n33 plus.t1 277.151
R220 plus.n28 plus.t12 277.151
R221 plus.n38 plus.t17 277.151
R222 plus.n40 plus.t5 277.151
R223 plus.n26 plus.t10 277.151
R224 plus.n45 plus.t0 277.151
R225 plus.n47 plus.t9 277.151
R226 plus.n5 plus.n4 161.489
R227 plus.n30 plus.n29 161.489
R228 plus.n7 plus.n4 161.3
R229 plus.n10 plus.n9 161.3
R230 plus.n12 plus.n11 161.3
R231 plus.n14 plus.n2 161.3
R232 plus.n17 plus.n16 161.3
R233 plus.n19 plus.n18 161.3
R234 plus.n21 plus.n0 161.3
R235 plus.n24 plus.n23 161.3
R236 plus.n32 plus.n29 161.3
R237 plus.n35 plus.n34 161.3
R238 plus.n37 plus.n36 161.3
R239 plus.n39 plus.n27 161.3
R240 plus.n42 plus.n41 161.3
R241 plus.n44 plus.n43 161.3
R242 plus.n46 plus.n25 161.3
R243 plus.n49 plus.n48 161.3
R244 plus.n7 plus.n6 51.852
R245 plus.n22 plus.n21 51.852
R246 plus.n47 plus.n46 51.852
R247 plus.n32 plus.n31 51.852
R248 plus.n9 plus.n8 47.4702
R249 plus.n20 plus.n19 47.4702
R250 plus.n45 plus.n44 47.4702
R251 plus.n34 plus.n33 47.4702
R252 plus.n12 plus.n3 43.0884
R253 plus.n16 plus.n1 43.0884
R254 plus.n41 plus.n26 43.0884
R255 plus.n37 plus.n28 43.0884
R256 plus.n14 plus.n13 38.7066
R257 plus.n15 plus.n14 38.7066
R258 plus.n40 plus.n39 38.7066
R259 plus.n39 plus.n38 38.7066
R260 plus.n13 plus.n12 34.3247
R261 plus.n16 plus.n15 34.3247
R262 plus.n41 plus.n40 34.3247
R263 plus.n38 plus.n37 34.3247
R264 plus.n9 plus.n3 29.9429
R265 plus.n19 plus.n1 29.9429
R266 plus.n44 plus.n26 29.9429
R267 plus.n34 plus.n28 29.9429
R268 plus plus.n49 25.9422
R269 plus.n8 plus.n7 25.5611
R270 plus.n21 plus.n20 25.5611
R271 plus.n46 plus.n45 25.5611
R272 plus.n33 plus.n32 25.5611
R273 plus.n6 plus.n5 21.1793
R274 plus.n23 plus.n22 21.1793
R275 plus.n48 plus.n47 21.1793
R276 plus.n31 plus.n30 21.1793
R277 plus plus.n24 7.95505
R278 plus.n10 plus.n4 0.189894
R279 plus.n11 plus.n10 0.189894
R280 plus.n11 plus.n2 0.189894
R281 plus.n17 plus.n2 0.189894
R282 plus.n18 plus.n17 0.189894
R283 plus.n18 plus.n0 0.189894
R284 plus.n24 plus.n0 0.189894
R285 plus.n49 plus.n25 0.189894
R286 plus.n43 plus.n25 0.189894
R287 plus.n43 plus.n42 0.189894
R288 plus.n42 plus.n27 0.189894
R289 plus.n36 plus.n27 0.189894
R290 plus.n36 plus.n35 0.189894
R291 plus.n35 plus.n29 0.189894
R292 drain_left.n10 drain_left.n8 240.589
R293 drain_left.n6 drain_left.n4 240.589
R294 drain_left.n2 drain_left.n0 240.589
R295 drain_left.n16 drain_left.n15 240.132
R296 drain_left.n14 drain_left.n13 240.132
R297 drain_left.n12 drain_left.n11 240.132
R298 drain_left.n10 drain_left.n9 240.132
R299 drain_left.n7 drain_left.n3 240.131
R300 drain_left.n6 drain_left.n5 240.131
R301 drain_left.n2 drain_left.n1 240.131
R302 drain_left drain_left.n7 22.6889
R303 drain_left.n3 drain_left.t14 19.8005
R304 drain_left.n3 drain_left.t2 19.8005
R305 drain_left.n4 drain_left.t4 19.8005
R306 drain_left.n4 drain_left.t11 19.8005
R307 drain_left.n5 drain_left.t7 19.8005
R308 drain_left.n5 drain_left.t18 19.8005
R309 drain_left.n1 drain_left.t19 19.8005
R310 drain_left.n1 drain_left.t9 19.8005
R311 drain_left.n0 drain_left.t3 19.8005
R312 drain_left.n0 drain_left.t10 19.8005
R313 drain_left.n15 drain_left.t8 19.8005
R314 drain_left.n15 drain_left.t15 19.8005
R315 drain_left.n13 drain_left.t17 19.8005
R316 drain_left.n13 drain_left.t1 19.8005
R317 drain_left.n11 drain_left.t6 19.8005
R318 drain_left.n11 drain_left.t13 19.8005
R319 drain_left.n9 drain_left.t0 19.8005
R320 drain_left.n9 drain_left.t5 19.8005
R321 drain_left.n8 drain_left.t12 19.8005
R322 drain_left.n8 drain_left.t16 19.8005
R323 drain_left drain_left.n16 6.11011
R324 drain_left.n12 drain_left.n10 0.457397
R325 drain_left.n14 drain_left.n12 0.457397
R326 drain_left.n16 drain_left.n14 0.457397
R327 drain_left.n7 drain_left.n6 0.402051
R328 drain_left.n7 drain_left.n2 0.402051
C0 plus minus 3.47445f
C1 source drain_right 6.67852f
C2 drain_left minus 0.178609f
C3 drain_left plus 1.15323f
C4 drain_right minus 0.970184f
C5 drain_right plus 0.345653f
C6 source minus 1.22118f
C7 source plus 1.23504f
C8 drain_left drain_right 0.982528f
C9 source drain_left 6.67855f
C10 drain_right a_n1882_n1088# 3.95975f
C11 drain_left a_n1882_n1088# 4.21953f
C12 source a_n1882_n1088# 2.571512f
C13 minus a_n1882_n1088# 6.407832f
C14 plus a_n1882_n1088# 7.11281f
C15 drain_left.t3 a_n1882_n1088# 0.022806f
C16 drain_left.t10 a_n1882_n1088# 0.022806f
C17 drain_left.n0 a_n1882_n1088# 0.089185f
C18 drain_left.t19 a_n1882_n1088# 0.022806f
C19 drain_left.t9 a_n1882_n1088# 0.022806f
C20 drain_left.n1 a_n1882_n1088# 0.088618f
C21 drain_left.n2 a_n1882_n1088# 0.581177f
C22 drain_left.t14 a_n1882_n1088# 0.022806f
C23 drain_left.t2 a_n1882_n1088# 0.022806f
C24 drain_left.n3 a_n1882_n1088# 0.088618f
C25 drain_left.t4 a_n1882_n1088# 0.022806f
C26 drain_left.t11 a_n1882_n1088# 0.022806f
C27 drain_left.n4 a_n1882_n1088# 0.089185f
C28 drain_left.t7 a_n1882_n1088# 0.022806f
C29 drain_left.t18 a_n1882_n1088# 0.022806f
C30 drain_left.n5 a_n1882_n1088# 0.088618f
C31 drain_left.n6 a_n1882_n1088# 0.581177f
C32 drain_left.n7 a_n1882_n1088# 1.02744f
C33 drain_left.t12 a_n1882_n1088# 0.022806f
C34 drain_left.t16 a_n1882_n1088# 0.022806f
C35 drain_left.n8 a_n1882_n1088# 0.089185f
C36 drain_left.t0 a_n1882_n1088# 0.022806f
C37 drain_left.t5 a_n1882_n1088# 0.022806f
C38 drain_left.n9 a_n1882_n1088# 0.088618f
C39 drain_left.n10 a_n1882_n1088# 0.584657f
C40 drain_left.t6 a_n1882_n1088# 0.022806f
C41 drain_left.t13 a_n1882_n1088# 0.022806f
C42 drain_left.n11 a_n1882_n1088# 0.088618f
C43 drain_left.n12 a_n1882_n1088# 0.2868f
C44 drain_left.t17 a_n1882_n1088# 0.022806f
C45 drain_left.t1 a_n1882_n1088# 0.022806f
C46 drain_left.n13 a_n1882_n1088# 0.088618f
C47 drain_left.n14 a_n1882_n1088# 0.2868f
C48 drain_left.t8 a_n1882_n1088# 0.022806f
C49 drain_left.t15 a_n1882_n1088# 0.022806f
C50 drain_left.n15 a_n1882_n1088# 0.088618f
C51 drain_left.n16 a_n1882_n1088# 0.522994f
C52 plus.n0 a_n1882_n1088# 0.032853f
C53 plus.t11 a_n1882_n1088# 0.020255f
C54 plus.t18 a_n1882_n1088# 0.020255f
C55 plus.t2 a_n1882_n1088# 0.020255f
C56 plus.n1 a_n1882_n1088# 0.024245f
C57 plus.n2 a_n1882_n1088# 0.032853f
C58 plus.t6 a_n1882_n1088# 0.020255f
C59 plus.t13 a_n1882_n1088# 0.020255f
C60 plus.t14 a_n1882_n1088# 0.020255f
C61 plus.n3 a_n1882_n1088# 0.024245f
C62 plus.n4 a_n1882_n1088# 0.075175f
C63 plus.t19 a_n1882_n1088# 0.020255f
C64 plus.t3 a_n1882_n1088# 0.020255f
C65 plus.t7 a_n1882_n1088# 0.024635f
C66 plus.n5 a_n1882_n1088# 0.033142f
C67 plus.n6 a_n1882_n1088# 0.024245f
C68 plus.n7 a_n1882_n1088# 0.011506f
C69 plus.n8 a_n1882_n1088# 0.024245f
C70 plus.n9 a_n1882_n1088# 0.011506f
C71 plus.n10 a_n1882_n1088# 0.032853f
C72 plus.n11 a_n1882_n1088# 0.032853f
C73 plus.n12 a_n1882_n1088# 0.011506f
C74 plus.n13 a_n1882_n1088# 0.024245f
C75 plus.n14 a_n1882_n1088# 0.011506f
C76 plus.n15 a_n1882_n1088# 0.024245f
C77 plus.n16 a_n1882_n1088# 0.011506f
C78 plus.n17 a_n1882_n1088# 0.032853f
C79 plus.n18 a_n1882_n1088# 0.032853f
C80 plus.n19 a_n1882_n1088# 0.011506f
C81 plus.n20 a_n1882_n1088# 0.024245f
C82 plus.n21 a_n1882_n1088# 0.011506f
C83 plus.n22 a_n1882_n1088# 0.024245f
C84 plus.t4 a_n1882_n1088# 0.024635f
C85 plus.n23 a_n1882_n1088# 0.033092f
C86 plus.n24 a_n1882_n1088# 0.223422f
C87 plus.n25 a_n1882_n1088# 0.032853f
C88 plus.t16 a_n1882_n1088# 0.024635f
C89 plus.t9 a_n1882_n1088# 0.020255f
C90 plus.t0 a_n1882_n1088# 0.020255f
C91 plus.t10 a_n1882_n1088# 0.020255f
C92 plus.n26 a_n1882_n1088# 0.024245f
C93 plus.n27 a_n1882_n1088# 0.032853f
C94 plus.t5 a_n1882_n1088# 0.020255f
C95 plus.t17 a_n1882_n1088# 0.020255f
C96 plus.t12 a_n1882_n1088# 0.020255f
C97 plus.n28 a_n1882_n1088# 0.024245f
C98 plus.n29 a_n1882_n1088# 0.075175f
C99 plus.t1 a_n1882_n1088# 0.020255f
C100 plus.t15 a_n1882_n1088# 0.020255f
C101 plus.t8 a_n1882_n1088# 0.024635f
C102 plus.n30 a_n1882_n1088# 0.033142f
C103 plus.n31 a_n1882_n1088# 0.024245f
C104 plus.n32 a_n1882_n1088# 0.011506f
C105 plus.n33 a_n1882_n1088# 0.024245f
C106 plus.n34 a_n1882_n1088# 0.011506f
C107 plus.n35 a_n1882_n1088# 0.032853f
C108 plus.n36 a_n1882_n1088# 0.032853f
C109 plus.n37 a_n1882_n1088# 0.011506f
C110 plus.n38 a_n1882_n1088# 0.024245f
C111 plus.n39 a_n1882_n1088# 0.011506f
C112 plus.n40 a_n1882_n1088# 0.024245f
C113 plus.n41 a_n1882_n1088# 0.011506f
C114 plus.n42 a_n1882_n1088# 0.032853f
C115 plus.n43 a_n1882_n1088# 0.032853f
C116 plus.n44 a_n1882_n1088# 0.011506f
C117 plus.n45 a_n1882_n1088# 0.024245f
C118 plus.n46 a_n1882_n1088# 0.011506f
C119 plus.n47 a_n1882_n1088# 0.024245f
C120 plus.n48 a_n1882_n1088# 0.033092f
C121 plus.n49 a_n1882_n1088# 0.729213f
C122 source.t8 a_n1882_n1088# 0.150192f
C123 source.n0 a_n1882_n1088# 0.627887f
C124 source.t38 a_n1882_n1088# 0.026985f
C125 source.t10 a_n1882_n1088# 0.026985f
C126 source.n1 a_n1882_n1088# 0.087515f
C127 source.n2 a_n1882_n1088# 0.310269f
C128 source.t7 a_n1882_n1088# 0.026985f
C129 source.t9 a_n1882_n1088# 0.026985f
C130 source.n3 a_n1882_n1088# 0.087515f
C131 source.n4 a_n1882_n1088# 0.310269f
C132 source.t3 a_n1882_n1088# 0.026985f
C133 source.t4 a_n1882_n1088# 0.026985f
C134 source.n5 a_n1882_n1088# 0.087515f
C135 source.n6 a_n1882_n1088# 0.310269f
C136 source.t15 a_n1882_n1088# 0.026985f
C137 source.t36 a_n1882_n1088# 0.026985f
C138 source.n7 a_n1882_n1088# 0.087515f
C139 source.n8 a_n1882_n1088# 0.310269f
C140 source.t6 a_n1882_n1088# 0.150192f
C141 source.n9 a_n1882_n1088# 0.322609f
C142 source.t22 a_n1882_n1088# 0.150192f
C143 source.n10 a_n1882_n1088# 0.322609f
C144 source.t34 a_n1882_n1088# 0.026985f
C145 source.t28 a_n1882_n1088# 0.026985f
C146 source.n11 a_n1882_n1088# 0.087515f
C147 source.n12 a_n1882_n1088# 0.310269f
C148 source.t21 a_n1882_n1088# 0.026985f
C149 source.t17 a_n1882_n1088# 0.026985f
C150 source.n13 a_n1882_n1088# 0.087515f
C151 source.n14 a_n1882_n1088# 0.310269f
C152 source.t33 a_n1882_n1088# 0.026985f
C153 source.t30 a_n1882_n1088# 0.026985f
C154 source.n15 a_n1882_n1088# 0.087515f
C155 source.n16 a_n1882_n1088# 0.310269f
C156 source.t24 a_n1882_n1088# 0.026985f
C157 source.t16 a_n1882_n1088# 0.026985f
C158 source.n17 a_n1882_n1088# 0.087515f
C159 source.n18 a_n1882_n1088# 0.310269f
C160 source.t26 a_n1882_n1088# 0.150192f
C161 source.n19 a_n1882_n1088# 0.899553f
C162 source.t37 a_n1882_n1088# 0.150192f
C163 source.n20 a_n1882_n1088# 0.899554f
C164 source.t13 a_n1882_n1088# 0.026985f
C165 source.t1 a_n1882_n1088# 0.026985f
C166 source.n21 a_n1882_n1088# 0.087515f
C167 source.n22 a_n1882_n1088# 0.310269f
C168 source.t11 a_n1882_n1088# 0.026985f
C169 source.t14 a_n1882_n1088# 0.026985f
C170 source.n23 a_n1882_n1088# 0.087515f
C171 source.n24 a_n1882_n1088# 0.310269f
C172 source.t39 a_n1882_n1088# 0.026985f
C173 source.t12 a_n1882_n1088# 0.026985f
C174 source.n25 a_n1882_n1088# 0.087515f
C175 source.n26 a_n1882_n1088# 0.310269f
C176 source.t0 a_n1882_n1088# 0.026985f
C177 source.t2 a_n1882_n1088# 0.026985f
C178 source.n27 a_n1882_n1088# 0.087515f
C179 source.n28 a_n1882_n1088# 0.310269f
C180 source.t5 a_n1882_n1088# 0.150192f
C181 source.n29 a_n1882_n1088# 0.322609f
C182 source.t25 a_n1882_n1088# 0.150192f
C183 source.n30 a_n1882_n1088# 0.322609f
C184 source.t19 a_n1882_n1088# 0.026985f
C185 source.t31 a_n1882_n1088# 0.026985f
C186 source.n31 a_n1882_n1088# 0.087515f
C187 source.n32 a_n1882_n1088# 0.310269f
C188 source.t27 a_n1882_n1088# 0.026985f
C189 source.t20 a_n1882_n1088# 0.026985f
C190 source.n33 a_n1882_n1088# 0.087515f
C191 source.n34 a_n1882_n1088# 0.310269f
C192 source.t32 a_n1882_n1088# 0.026985f
C193 source.t29 a_n1882_n1088# 0.026985f
C194 source.n35 a_n1882_n1088# 0.087515f
C195 source.n36 a_n1882_n1088# 0.310269f
C196 source.t18 a_n1882_n1088# 0.026985f
C197 source.t35 a_n1882_n1088# 0.026985f
C198 source.n37 a_n1882_n1088# 0.087515f
C199 source.n38 a_n1882_n1088# 0.310269f
C200 source.t23 a_n1882_n1088# 0.150192f
C201 source.n39 a_n1882_n1088# 0.507768f
C202 source.n40 a_n1882_n1088# 0.687741f
C203 drain_right.t6 a_n1882_n1088# 0.023197f
C204 drain_right.t14 a_n1882_n1088# 0.023197f
C205 drain_right.n0 a_n1882_n1088# 0.090714f
C206 drain_right.t17 a_n1882_n1088# 0.023197f
C207 drain_right.t16 a_n1882_n1088# 0.023197f
C208 drain_right.n1 a_n1882_n1088# 0.090137f
C209 drain_right.n2 a_n1882_n1088# 0.591138f
C210 drain_right.t8 a_n1882_n1088# 0.023197f
C211 drain_right.t19 a_n1882_n1088# 0.023197f
C212 drain_right.n3 a_n1882_n1088# 0.090137f
C213 drain_right.t7 a_n1882_n1088# 0.023197f
C214 drain_right.t1 a_n1882_n1088# 0.023197f
C215 drain_right.n4 a_n1882_n1088# 0.090714f
C216 drain_right.t18 a_n1882_n1088# 0.023197f
C217 drain_right.t11 a_n1882_n1088# 0.023197f
C218 drain_right.n5 a_n1882_n1088# 0.090137f
C219 drain_right.n6 a_n1882_n1088# 0.591138f
C220 drain_right.n7 a_n1882_n1088# 0.988327f
C221 drain_right.t0 a_n1882_n1088# 0.023197f
C222 drain_right.t2 a_n1882_n1088# 0.023197f
C223 drain_right.n8 a_n1882_n1088# 0.090714f
C224 drain_right.t9 a_n1882_n1088# 0.023197f
C225 drain_right.t13 a_n1882_n1088# 0.023197f
C226 drain_right.n9 a_n1882_n1088# 0.090137f
C227 drain_right.n10 a_n1882_n1088# 0.594678f
C228 drain_right.t4 a_n1882_n1088# 0.023197f
C229 drain_right.t10 a_n1882_n1088# 0.023197f
C230 drain_right.n11 a_n1882_n1088# 0.090137f
C231 drain_right.n12 a_n1882_n1088# 0.291715f
C232 drain_right.t15 a_n1882_n1088# 0.023197f
C233 drain_right.t5 a_n1882_n1088# 0.023197f
C234 drain_right.n13 a_n1882_n1088# 0.090137f
C235 drain_right.n14 a_n1882_n1088# 0.291715f
C236 drain_right.t12 a_n1882_n1088# 0.023197f
C237 drain_right.t3 a_n1882_n1088# 0.023197f
C238 drain_right.n15 a_n1882_n1088# 0.090137f
C239 drain_right.n16 a_n1882_n1088# 0.531957f
C240 minus.n0 a_n1882_n1088# 0.032241f
C241 minus.t9 a_n1882_n1088# 0.024176f
C242 minus.t11 a_n1882_n1088# 0.019878f
C243 minus.t19 a_n1882_n1088# 0.019878f
C244 minus.t2 a_n1882_n1088# 0.019878f
C245 minus.n1 a_n1882_n1088# 0.023793f
C246 minus.n2 a_n1882_n1088# 0.032241f
C247 minus.t5 a_n1882_n1088# 0.019878f
C248 minus.t14 a_n1882_n1088# 0.019878f
C249 minus.t18 a_n1882_n1088# 0.019878f
C250 minus.n3 a_n1882_n1088# 0.023793f
C251 minus.n4 a_n1882_n1088# 0.073775f
C252 minus.t1 a_n1882_n1088# 0.019878f
C253 minus.t7 a_n1882_n1088# 0.019878f
C254 minus.t13 a_n1882_n1088# 0.024176f
C255 minus.n5 a_n1882_n1088# 0.032525f
C256 minus.n6 a_n1882_n1088# 0.023793f
C257 minus.n7 a_n1882_n1088# 0.011292f
C258 minus.n8 a_n1882_n1088# 0.023793f
C259 minus.n9 a_n1882_n1088# 0.011292f
C260 minus.n10 a_n1882_n1088# 0.032241f
C261 minus.n11 a_n1882_n1088# 0.032241f
C262 minus.n12 a_n1882_n1088# 0.011292f
C263 minus.n13 a_n1882_n1088# 0.023793f
C264 minus.n14 a_n1882_n1088# 0.011292f
C265 minus.n15 a_n1882_n1088# 0.023793f
C266 minus.n16 a_n1882_n1088# 0.011292f
C267 minus.n17 a_n1882_n1088# 0.032241f
C268 minus.n18 a_n1882_n1088# 0.032241f
C269 minus.n19 a_n1882_n1088# 0.011292f
C270 minus.n20 a_n1882_n1088# 0.023793f
C271 minus.n21 a_n1882_n1088# 0.011292f
C272 minus.n22 a_n1882_n1088# 0.023793f
C273 minus.n23 a_n1882_n1088# 0.032476f
C274 minus.n24 a_n1882_n1088# 0.738232f
C275 minus.n25 a_n1882_n1088# 0.032241f
C276 minus.t0 a_n1882_n1088# 0.019878f
C277 minus.t17 a_n1882_n1088# 0.019878f
C278 minus.t6 a_n1882_n1088# 0.019878f
C279 minus.n26 a_n1882_n1088# 0.023793f
C280 minus.n27 a_n1882_n1088# 0.032241f
C281 minus.t3 a_n1882_n1088# 0.019878f
C282 minus.t15 a_n1882_n1088# 0.019878f
C283 minus.t8 a_n1882_n1088# 0.019878f
C284 minus.n28 a_n1882_n1088# 0.023793f
C285 minus.n29 a_n1882_n1088# 0.073775f
C286 minus.t4 a_n1882_n1088# 0.019878f
C287 minus.t16 a_n1882_n1088# 0.019878f
C288 minus.t10 a_n1882_n1088# 0.024176f
C289 minus.n30 a_n1882_n1088# 0.032525f
C290 minus.n31 a_n1882_n1088# 0.023793f
C291 minus.n32 a_n1882_n1088# 0.011292f
C292 minus.n33 a_n1882_n1088# 0.023793f
C293 minus.n34 a_n1882_n1088# 0.011292f
C294 minus.n35 a_n1882_n1088# 0.032241f
C295 minus.n36 a_n1882_n1088# 0.032241f
C296 minus.n37 a_n1882_n1088# 0.011292f
C297 minus.n38 a_n1882_n1088# 0.023793f
C298 minus.n39 a_n1882_n1088# 0.011292f
C299 minus.n40 a_n1882_n1088# 0.023793f
C300 minus.n41 a_n1882_n1088# 0.011292f
C301 minus.n42 a_n1882_n1088# 0.032241f
C302 minus.n43 a_n1882_n1088# 0.032241f
C303 minus.n44 a_n1882_n1088# 0.011292f
C304 minus.n45 a_n1882_n1088# 0.023793f
C305 minus.n46 a_n1882_n1088# 0.011292f
C306 minus.n47 a_n1882_n1088# 0.023793f
C307 minus.t12 a_n1882_n1088# 0.024176f
C308 minus.n48 a_n1882_n1088# 0.032476f
C309 minus.n49 a_n1882_n1088# 0.20909f
C310 minus.n50 a_n1882_n1088# 0.913553f
.ends

