* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t10 plus.t0 drain_left.t0 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_left.t5 plus.t1 source.t9 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X2 a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X3 source.t11 minus.t0 drain_right.t5 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 drain_left.t4 plus.t2 source.t8 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X5 source.t1 minus.t1 drain_right.t4 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 drain_right.t3 minus.t2 source.t4 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X7 drain_left.t3 plus.t3 source.t7 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X8 a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X9 drain_right.t2 minus.t3 source.t0 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X10 drain_right.t1 minus.t4 source.t3 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X11 drain_right.t0 minus.t5 source.t2 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X12 a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X13 source.t6 plus.t4 drain_left.t2 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X14 a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X15 drain_left.t1 plus.t5 source.t5 a_n1180_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
R0 plus.n0 plus.t2 366.32
R1 plus.n2 plus.t3 366.32
R2 plus.n4 plus.t5 366.32
R3 plus.n6 plus.t1 366.32
R4 plus.n1 plus.t0 318.12
R5 plus.n5 plus.t4 318.12
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 23.6695
R15 plus plus.n3 8.34141
R16 drain_left.n2 drain_left.n0 289.615
R17 drain_left.n11 drain_left.n9 289.615
R18 drain_left.n3 drain_left.n2 185
R19 drain_left.n12 drain_left.n11 185
R20 drain_left.t5 drain_left.n1 167.117
R21 drain_left.t4 drain_left.n10 167.117
R22 drain_left.n8 drain_left.n7 100.865
R23 drain_left.n17 drain_left.n16 100.796
R24 drain_left.n2 drain_left.t5 52.3082
R25 drain_left.n11 drain_left.t4 52.3082
R26 drain_left.n17 drain_left.n15 48.5884
R27 drain_left.n8 drain_left.n6 48.408
R28 drain_left drain_left.n8 21.1663
R29 drain_left.n7 drain_left.t2 9.9005
R30 drain_left.n7 drain_left.t1 9.9005
R31 drain_left.n16 drain_left.t0 9.9005
R32 drain_left.n16 drain_left.t3 9.9005
R33 drain_left.n3 drain_left.n1 9.71174
R34 drain_left.n12 drain_left.n10 9.71174
R35 drain_left.n6 drain_left.n5 9.45567
R36 drain_left.n15 drain_left.n14 9.45567
R37 drain_left.n5 drain_left.n4 9.3005
R38 drain_left.n14 drain_left.n13 9.3005
R39 drain_left.n6 drain_left.n0 8.14595
R40 drain_left.n15 drain_left.n9 8.14595
R41 drain_left.n4 drain_left.n3 7.3702
R42 drain_left.n13 drain_left.n12 7.3702
R43 drain_left drain_left.n17 6.15322
R44 drain_left.n4 drain_left.n0 5.81868
R45 drain_left.n13 drain_left.n9 5.81868
R46 drain_left.n5 drain_left.n1 3.44771
R47 drain_left.n14 drain_left.n10 3.44771
R48 source.n34 source.n32 289.615
R49 source.n24 source.n22 289.615
R50 source.n2 source.n0 289.615
R51 source.n12 source.n10 289.615
R52 source.n35 source.n34 185
R53 source.n25 source.n24 185
R54 source.n3 source.n2 185
R55 source.n13 source.n12 185
R56 source.t4 source.n33 167.117
R57 source.t5 source.n23 167.117
R58 source.t7 source.n1 167.117
R59 source.t2 source.n11 167.117
R60 source.n9 source.n8 84.1169
R61 source.n19 source.n18 84.1169
R62 source.n31 source.n30 84.1168
R63 source.n21 source.n20 84.1168
R64 source.n34 source.t4 52.3082
R65 source.n24 source.t5 52.3082
R66 source.n2 source.t7 52.3082
R67 source.n12 source.t2 52.3082
R68 source.n39 source.n38 31.4096
R69 source.n29 source.n28 31.4096
R70 source.n7 source.n6 31.4096
R71 source.n17 source.n16 31.4096
R72 source.n21 source.n19 14.712
R73 source.n30 source.t0 9.9005
R74 source.n30 source.t1 9.9005
R75 source.n20 source.t9 9.9005
R76 source.n20 source.t6 9.9005
R77 source.n8 source.t8 9.9005
R78 source.n8 source.t10 9.9005
R79 source.n18 source.t3 9.9005
R80 source.n18 source.t11 9.9005
R81 source.n35 source.n33 9.71174
R82 source.n25 source.n23 9.71174
R83 source.n3 source.n1 9.71174
R84 source.n13 source.n11 9.71174
R85 source.n38 source.n37 9.45567
R86 source.n28 source.n27 9.45567
R87 source.n6 source.n5 9.45567
R88 source.n16 source.n15 9.45567
R89 source.n37 source.n36 9.3005
R90 source.n27 source.n26 9.3005
R91 source.n5 source.n4 9.3005
R92 source.n15 source.n14 9.3005
R93 source.n40 source.n7 8.69904
R94 source.n38 source.n32 8.14595
R95 source.n28 source.n22 8.14595
R96 source.n6 source.n0 8.14595
R97 source.n16 source.n10 8.14595
R98 source.n36 source.n35 7.3702
R99 source.n26 source.n25 7.3702
R100 source.n4 source.n3 7.3702
R101 source.n14 source.n13 7.3702
R102 source.n36 source.n32 5.81868
R103 source.n26 source.n22 5.81868
R104 source.n4 source.n0 5.81868
R105 source.n14 source.n10 5.81868
R106 source.n40 source.n39 5.51343
R107 source.n37 source.n33 3.44771
R108 source.n27 source.n23 3.44771
R109 source.n5 source.n1 3.44771
R110 source.n15 source.n11 3.44771
R111 source.n17 source.n9 0.720328
R112 source.n31 source.n29 0.720328
R113 source.n19 source.n17 0.5005
R114 source.n9 source.n7 0.5005
R115 source.n29 source.n21 0.5005
R116 source.n39 source.n31 0.5005
R117 source source.n40 0.188
R118 minus.n2 minus.t4 366.32
R119 minus.n0 minus.t5 366.32
R120 minus.n6 minus.t2 366.32
R121 minus.n4 minus.t3 366.32
R122 minus.n1 minus.t0 318.12
R123 minus.n5 minus.t1 318.12
R124 minus.n3 minus.n0 161.489
R125 minus.n7 minus.n4 161.489
R126 minus.n3 minus.n2 161.3
R127 minus.n7 minus.n6 161.3
R128 minus.n2 minus.n1 36.5157
R129 minus.n1 minus.n0 36.5157
R130 minus.n5 minus.n4 36.5157
R131 minus.n6 minus.n5 36.5157
R132 minus.n8 minus.n3 26.0005
R133 minus.n8 minus.n7 6.48535
R134 minus minus.n8 0.188
R135 drain_right.n2 drain_right.n0 289.615
R136 drain_right.n12 drain_right.n10 289.615
R137 drain_right.n3 drain_right.n2 185
R138 drain_right.n13 drain_right.n12 185
R139 drain_right.t2 drain_right.n1 167.117
R140 drain_right.t1 drain_right.n11 167.117
R141 drain_right.n17 drain_right.n9 101.296
R142 drain_right.n8 drain_right.n7 100.865
R143 drain_right.n2 drain_right.t2 52.3082
R144 drain_right.n12 drain_right.t1 52.3082
R145 drain_right.n8 drain_right.n6 48.408
R146 drain_right.n17 drain_right.n16 48.0884
R147 drain_right drain_right.n8 20.6131
R148 drain_right.n7 drain_right.t4 9.9005
R149 drain_right.n7 drain_right.t3 9.9005
R150 drain_right.n9 drain_right.t5 9.9005
R151 drain_right.n9 drain_right.t0 9.9005
R152 drain_right.n3 drain_right.n1 9.71174
R153 drain_right.n13 drain_right.n11 9.71174
R154 drain_right.n6 drain_right.n5 9.45567
R155 drain_right.n16 drain_right.n15 9.45567
R156 drain_right.n5 drain_right.n4 9.3005
R157 drain_right.n15 drain_right.n14 9.3005
R158 drain_right.n6 drain_right.n0 8.14595
R159 drain_right.n16 drain_right.n10 8.14595
R160 drain_right.n4 drain_right.n3 7.3702
R161 drain_right.n14 drain_right.n13 7.3702
R162 drain_right drain_right.n17 5.90322
R163 drain_right.n4 drain_right.n0 5.81868
R164 drain_right.n14 drain_right.n10 5.81868
R165 drain_right.n5 drain_right.n1 3.44771
R166 drain_right.n15 drain_right.n11 3.44771
C0 drain_left drain_right 0.547725f
C1 minus source 0.698843f
C2 drain_left minus 0.176775f
C3 drain_left source 3.87172f
C4 plus drain_right 0.270474f
C5 plus minus 2.77789f
C6 plus source 0.712919f
C7 plus drain_left 0.776988f
C8 drain_right minus 0.667487f
C9 drain_right source 3.8678f
C10 drain_right a_n1180_n1288# 3.07623f
C11 drain_left a_n1180_n1288# 3.22681f
C12 source a_n1180_n1288# 2.308679f
C13 minus a_n1180_n1288# 3.727622f
C14 plus a_n1180_n1288# 4.499111f
C15 drain_right.n0 a_n1180_n1288# 0.03367f
C16 drain_right.n1 a_n1180_n1288# 0.074499f
C17 drain_right.t2 a_n1180_n1288# 0.055907f
C18 drain_right.n2 a_n1180_n1288# 0.058306f
C19 drain_right.n3 a_n1180_n1288# 0.018796f
C20 drain_right.n4 a_n1180_n1288# 0.012396f
C21 drain_right.n5 a_n1180_n1288# 0.164213f
C22 drain_right.n6 a_n1180_n1288# 0.053305f
C23 drain_right.t4 a_n1180_n1288# 0.036459f
C24 drain_right.t3 a_n1180_n1288# 0.036459f
C25 drain_right.n7 a_n1180_n1288# 0.229208f
C26 drain_right.n8 a_n1180_n1288# 0.760102f
C27 drain_right.t5 a_n1180_n1288# 0.036459f
C28 drain_right.t0 a_n1180_n1288# 0.036459f
C29 drain_right.n9 a_n1180_n1288# 0.23033f
C30 drain_right.n10 a_n1180_n1288# 0.03367f
C31 drain_right.n11 a_n1180_n1288# 0.074499f
C32 drain_right.t1 a_n1180_n1288# 0.055907f
C33 drain_right.n12 a_n1180_n1288# 0.058306f
C34 drain_right.n13 a_n1180_n1288# 0.018796f
C35 drain_right.n14 a_n1180_n1288# 0.012396f
C36 drain_right.n15 a_n1180_n1288# 0.164213f
C37 drain_right.n16 a_n1180_n1288# 0.052848f
C38 drain_right.n17 a_n1180_n1288# 0.52974f
C39 minus.t5 a_n1180_n1288# 0.063198f
C40 minus.n0 a_n1180_n1288# 0.053155f
C41 minus.t4 a_n1180_n1288# 0.063198f
C42 minus.t0 a_n1180_n1288# 0.057406f
C43 minus.n1 a_n1180_n1288# 0.042098f
C44 minus.n2 a_n1180_n1288# 0.053098f
C45 minus.n3 a_n1180_n1288# 0.835681f
C46 minus.t3 a_n1180_n1288# 0.063198f
C47 minus.n4 a_n1180_n1288# 0.053155f
C48 minus.t1 a_n1180_n1288# 0.057406f
C49 minus.n5 a_n1180_n1288# 0.042098f
C50 minus.t2 a_n1180_n1288# 0.063198f
C51 minus.n6 a_n1180_n1288# 0.053098f
C52 minus.n7 a_n1180_n1288# 0.30256f
C53 minus.n8 a_n1180_n1288# 0.97183f
C54 source.n0 a_n1180_n1288# 0.041505f
C55 source.n1 a_n1180_n1288# 0.091835f
C56 source.t7 a_n1180_n1288# 0.068917f
C57 source.n2 a_n1180_n1288# 0.071874f
C58 source.n3 a_n1180_n1288# 0.023169f
C59 source.n4 a_n1180_n1288# 0.015281f
C60 source.n5 a_n1180_n1288# 0.202426f
C61 source.n6 a_n1180_n1288# 0.045499f
C62 source.n7 a_n1180_n1288# 0.422325f
C63 source.t8 a_n1180_n1288# 0.044943f
C64 source.t10 a_n1180_n1288# 0.044943f
C65 source.n8 a_n1180_n1288# 0.240263f
C66 source.n9 a_n1180_n1288# 0.332853f
C67 source.n10 a_n1180_n1288# 0.041505f
C68 source.n11 a_n1180_n1288# 0.091835f
C69 source.t2 a_n1180_n1288# 0.068917f
C70 source.n12 a_n1180_n1288# 0.071874f
C71 source.n13 a_n1180_n1288# 0.023169f
C72 source.n14 a_n1180_n1288# 0.015281f
C73 source.n15 a_n1180_n1288# 0.202426f
C74 source.n16 a_n1180_n1288# 0.045499f
C75 source.n17 a_n1180_n1288# 0.135182f
C76 source.t3 a_n1180_n1288# 0.044943f
C77 source.t11 a_n1180_n1288# 0.044943f
C78 source.n18 a_n1180_n1288# 0.240263f
C79 source.n19 a_n1180_n1288# 0.930047f
C80 source.t9 a_n1180_n1288# 0.044943f
C81 source.t6 a_n1180_n1288# 0.044943f
C82 source.n20 a_n1180_n1288# 0.240262f
C83 source.n21 a_n1180_n1288# 0.930049f
C84 source.n22 a_n1180_n1288# 0.041505f
C85 source.n23 a_n1180_n1288# 0.091835f
C86 source.t5 a_n1180_n1288# 0.068917f
C87 source.n24 a_n1180_n1288# 0.071874f
C88 source.n25 a_n1180_n1288# 0.023169f
C89 source.n26 a_n1180_n1288# 0.015281f
C90 source.n27 a_n1180_n1288# 0.202426f
C91 source.n28 a_n1180_n1288# 0.045499f
C92 source.n29 a_n1180_n1288# 0.135182f
C93 source.t0 a_n1180_n1288# 0.044943f
C94 source.t1 a_n1180_n1288# 0.044943f
C95 source.n30 a_n1180_n1288# 0.240262f
C96 source.n31 a_n1180_n1288# 0.332854f
C97 source.n32 a_n1180_n1288# 0.041505f
C98 source.n33 a_n1180_n1288# 0.091835f
C99 source.t4 a_n1180_n1288# 0.068917f
C100 source.n34 a_n1180_n1288# 0.071874f
C101 source.n35 a_n1180_n1288# 0.023169f
C102 source.n36 a_n1180_n1288# 0.015281f
C103 source.n37 a_n1180_n1288# 0.202426f
C104 source.n38 a_n1180_n1288# 0.045499f
C105 source.n39 a_n1180_n1288# 0.269637f
C106 source.n40 a_n1180_n1288# 0.701388f
C107 drain_left.n0 a_n1180_n1288# 0.032908f
C108 drain_left.n1 a_n1180_n1288# 0.072814f
C109 drain_left.t5 a_n1180_n1288# 0.054643f
C110 drain_left.n2 a_n1180_n1288# 0.056987f
C111 drain_left.n3 a_n1180_n1288# 0.01837f
C112 drain_left.n4 a_n1180_n1288# 0.012116f
C113 drain_left.n5 a_n1180_n1288# 0.160499f
C114 drain_left.n6 a_n1180_n1288# 0.052099f
C115 drain_left.t2 a_n1180_n1288# 0.035634f
C116 drain_left.t1 a_n1180_n1288# 0.035634f
C117 drain_left.n7 a_n1180_n1288# 0.224024f
C118 drain_left.n8 a_n1180_n1288# 0.787383f
C119 drain_left.n9 a_n1180_n1288# 0.032908f
C120 drain_left.n10 a_n1180_n1288# 0.072814f
C121 drain_left.t4 a_n1180_n1288# 0.054643f
C122 drain_left.n11 a_n1180_n1288# 0.056987f
C123 drain_left.n12 a_n1180_n1288# 0.01837f
C124 drain_left.n13 a_n1180_n1288# 0.012116f
C125 drain_left.n14 a_n1180_n1288# 0.160499f
C126 drain_left.n15 a_n1180_n1288# 0.052467f
C127 drain_left.t0 a_n1180_n1288# 0.035634f
C128 drain_left.t3 a_n1180_n1288# 0.035634f
C129 drain_left.n16 a_n1180_n1288# 0.223866f
C130 drain_left.n17 a_n1180_n1288# 0.50955f
C131 plus.t2 a_n1180_n1288# 0.065031f
C132 plus.n0 a_n1180_n1288# 0.054696f
C133 plus.t0 a_n1180_n1288# 0.059071f
C134 plus.n1 a_n1180_n1288# 0.043318f
C135 plus.t3 a_n1180_n1288# 0.065031f
C136 plus.n2 a_n1180_n1288# 0.054637f
C137 plus.n3 a_n1180_n1288# 0.335797f
C138 plus.t5 a_n1180_n1288# 0.065031f
C139 plus.n4 a_n1180_n1288# 0.054696f
C140 plus.t1 a_n1180_n1288# 0.065031f
C141 plus.t4 a_n1180_n1288# 0.059071f
C142 plus.n5 a_n1180_n1288# 0.043318f
C143 plus.n6 a_n1180_n1288# 0.054637f
C144 plus.n7 a_n1180_n1288# 0.829953f
.ends

