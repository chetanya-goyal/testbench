* NGSPICE file created from diffpair493.ext - technology: sky130A

.subckt diffpair493 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t10 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t6 plus.t1 source.t7 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X2 drain_right.t7 minus.t0 source.t4 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X3 a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X4 source.t11 plus.t2 drain_left.t5 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 drain_left.t4 plus.t3 source.t8 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X7 source.t0 minus.t1 drain_right.t6 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 source.t15 minus.t2 drain_right.t5 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 source.t2 minus.t3 drain_right.t4 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X10 source.t9 plus.t4 drain_left.t3 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X11 drain_right.t3 minus.t4 source.t1 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X12 drain_right.t2 minus.t5 source.t5 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X13 a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X14 drain_right.t1 minus.t6 source.t6 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X15 drain_left.t2 plus.t5 source.t13 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X16 source.t3 minus.t7 drain_right.t0 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X17 source.t12 plus.t6 drain_left.t1 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X18 a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X19 source.t14 plus.t7 drain_left.t0 a_n1246_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n1 plus.t4 2007.24
R1 plus.n5 plus.t5 2007.24
R2 plus.n8 plus.t1 2007.24
R3 plus.n12 plus.t6 2007.24
R4 plus.n2 plus.t3 1964.15
R5 plus.n4 plus.t7 1964.15
R6 plus.n9 plus.t2 1964.15
R7 plus.n11 plus.t0 1964.15
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 38.7066
R15 plus.n4 plus.n3 38.7066
R16 plus.n11 plus.n10 38.7066
R17 plus.n10 plus.n9 38.7066
R18 plus.n2 plus.n1 34.3247
R19 plus.n5 plus.n4 34.3247
R20 plus.n12 plus.n11 34.3247
R21 plus.n9 plus.n8 34.3247
R22 plus plus.n13 28.802
R23 plus plus.n6 13.224
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n3 source.t9 45.521
R27 source.n4 source.t6 45.521
R28 source.n7 source.t3 45.521
R29 source.n15 source.t1 45.5208
R30 source.n12 source.t2 45.5208
R31 source.n11 source.t7 45.5208
R32 source.n8 source.t12 45.5208
R33 source.n0 source.t13 45.5208
R34 source.n2 source.n1 44.201
R35 source.n6 source.n5 44.201
R36 source.n14 source.n13 44.2008
R37 source.n10 source.n9 44.2008
R38 source.n8 source.n7 24.0173
R39 source.n16 source.n0 18.526
R40 source.n16 source.n15 5.49188
R41 source.n13 source.t5 1.3205
R42 source.n13 source.t0 1.3205
R43 source.n9 source.t10 1.3205
R44 source.n9 source.t11 1.3205
R45 source.n1 source.t8 1.3205
R46 source.n1 source.t14 1.3205
R47 source.n5 source.t4 1.3205
R48 source.n5 source.t15 1.3205
R49 source.n4 source.n3 0.470328
R50 source.n12 source.n11 0.470328
R51 source.n7 source.n6 0.457397
R52 source.n6 source.n4 0.457397
R53 source.n3 source.n2 0.457397
R54 source.n2 source.n0 0.457397
R55 source.n10 source.n8 0.457397
R56 source.n11 source.n10 0.457397
R57 source.n14 source.n12 0.457397
R58 source.n15 source.n14 0.457397
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 61.3367
R61 drain_left.n2 drain_left.n1 61.0527
R62 drain_left.n2 drain_left.n0 61.0527
R63 drain_left.n5 drain_left.n4 60.8796
R64 drain_left drain_left.n2 31.2389
R65 drain_left drain_left.n5 6.11011
R66 drain_left.n1 drain_left.t5 1.3205
R67 drain_left.n1 drain_left.t6 1.3205
R68 drain_left.n0 drain_left.t1 1.3205
R69 drain_left.n0 drain_left.t7 1.3205
R70 drain_left.n4 drain_left.t0 1.3205
R71 drain_left.n4 drain_left.t2 1.3205
R72 drain_left.n3 drain_left.t3 1.3205
R73 drain_left.n3 drain_left.t4 1.3205
R74 minus.n5 minus.t7 2007.24
R75 minus.n1 minus.t6 2007.24
R76 minus.n12 minus.t4 2007.24
R77 minus.n8 minus.t3 2007.24
R78 minus.n4 minus.t0 1964.15
R79 minus.n2 minus.t2 1964.15
R80 minus.n11 minus.t1 1964.15
R81 minus.n9 minus.t5 1964.15
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 38.7066
R89 minus.n3 minus.n2 38.7066
R90 minus.n10 minus.n9 38.7066
R91 minus.n11 minus.n10 38.7066
R92 minus.n14 minus.n6 36.0573
R93 minus.n5 minus.n4 34.3247
R94 minus.n2 minus.n1 34.3247
R95 minus.n9 minus.n8 34.3247
R96 minus.n12 minus.n11 34.3247
R97 minus.n14 minus.n13 6.44368
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 61.3365
R102 drain_right.n2 drain_right.n1 61.0527
R103 drain_right.n2 drain_right.n0 61.0527
R104 drain_right.n5 drain_right.n4 60.8798
R105 drain_right drain_right.n2 30.6857
R106 drain_right drain_right.n5 6.11011
R107 drain_right.n1 drain_right.t6 1.3205
R108 drain_right.n1 drain_right.t3 1.3205
R109 drain_right.n0 drain_right.t4 1.3205
R110 drain_right.n0 drain_right.t2 1.3205
R111 drain_right.n3 drain_right.t5 1.3205
R112 drain_right.n3 drain_right.t1 1.3205
R113 drain_right.n4 drain_right.t0 1.3205
R114 drain_right.n4 drain_right.t7 1.3205
C0 source plus 2.57597f
C1 source minus 2.56193f
C2 minus plus 5.2639f
C3 drain_right drain_left 0.58123f
C4 drain_right source 24.1286f
C5 drain_right plus 0.269775f
C6 drain_right minus 3.19682f
C7 source drain_left 24.130001f
C8 drain_left plus 3.31361f
C9 drain_left minus 0.17017f
C10 drain_right a_n1246_n3888# 6.71892f
C11 drain_left a_n1246_n3888# 6.91115f
C12 source a_n1246_n3888# 10.01166f
C13 minus a_n1246_n3888# 4.995718f
C14 plus a_n1246_n3888# 7.36227f
C15 drain_right.t4 a_n1246_n3888# 0.446009f
C16 drain_right.t2 a_n1246_n3888# 0.446009f
C17 drain_right.n0 a_n1246_n3888# 4.03255f
C18 drain_right.t6 a_n1246_n3888# 0.446009f
C19 drain_right.t3 a_n1246_n3888# 0.446009f
C20 drain_right.n1 a_n1246_n3888# 4.03255f
C21 drain_right.n2 a_n1246_n3888# 2.59417f
C22 drain_right.t5 a_n1246_n3888# 0.446009f
C23 drain_right.t1 a_n1246_n3888# 0.446009f
C24 drain_right.n3 a_n1246_n3888# 4.03462f
C25 drain_right.t0 a_n1246_n3888# 0.446009f
C26 drain_right.t7 a_n1246_n3888# 0.446009f
C27 drain_right.n4 a_n1246_n3888# 4.0314f
C28 drain_right.n5 a_n1246_n3888# 1.15783f
C29 minus.n0 a_n1246_n3888# 0.130068f
C30 minus.t7 a_n1246_n3888# 0.509862f
C31 minus.t0 a_n1246_n3888# 0.505565f
C32 minus.t2 a_n1246_n3888# 0.505565f
C33 minus.t6 a_n1246_n3888# 0.509862f
C34 minus.n1 a_n1246_n3888# 0.216852f
C35 minus.n2 a_n1246_n3888# 0.200329f
C36 minus.n3 a_n1246_n3888# 0.020921f
C37 minus.n4 a_n1246_n3888# 0.200329f
C38 minus.n5 a_n1246_n3888# 0.216769f
C39 minus.n6 a_n1246_n3888# 2.09606f
C40 minus.n7 a_n1246_n3888# 0.130068f
C41 minus.t1 a_n1246_n3888# 0.505565f
C42 minus.t5 a_n1246_n3888# 0.505565f
C43 minus.t3 a_n1246_n3888# 0.509862f
C44 minus.n8 a_n1246_n3888# 0.216852f
C45 minus.n9 a_n1246_n3888# 0.200329f
C46 minus.n10 a_n1246_n3888# 0.020921f
C47 minus.n11 a_n1246_n3888# 0.200329f
C48 minus.t4 a_n1246_n3888# 0.509862f
C49 minus.n12 a_n1246_n3888# 0.216769f
C50 minus.n13 a_n1246_n3888# 0.382586f
C51 minus.n14 a_n1246_n3888# 2.54989f
C52 drain_left.t1 a_n1246_n3888# 0.445242f
C53 drain_left.t7 a_n1246_n3888# 0.445242f
C54 drain_left.n0 a_n1246_n3888# 4.02561f
C55 drain_left.t5 a_n1246_n3888# 0.445242f
C56 drain_left.t6 a_n1246_n3888# 0.445242f
C57 drain_left.n1 a_n1246_n3888# 4.02561f
C58 drain_left.n2 a_n1246_n3888# 2.66872f
C59 drain_left.t3 a_n1246_n3888# 0.445242f
C60 drain_left.t4 a_n1246_n3888# 0.445242f
C61 drain_left.n3 a_n1246_n3888# 4.0277f
C62 drain_left.t0 a_n1246_n3888# 0.445242f
C63 drain_left.t2 a_n1246_n3888# 0.445242f
C64 drain_left.n4 a_n1246_n3888# 4.02446f
C65 drain_left.n5 a_n1246_n3888# 1.15583f
C66 source.t13 a_n1246_n3888# 3.54006f
C67 source.n0 a_n1246_n3888# 1.62775f
C68 source.t8 a_n1246_n3888# 0.315891f
C69 source.t14 a_n1246_n3888# 0.315891f
C70 source.n1 a_n1246_n3888# 2.77483f
C71 source.n2 a_n1246_n3888# 0.340971f
C72 source.t9 a_n1246_n3888# 3.54007f
C73 source.n3 a_n1246_n3888# 0.438368f
C74 source.t6 a_n1246_n3888# 3.54007f
C75 source.n4 a_n1246_n3888# 0.438368f
C76 source.t4 a_n1246_n3888# 0.315891f
C77 source.t15 a_n1246_n3888# 0.315891f
C78 source.n5 a_n1246_n3888# 2.77483f
C79 source.n6 a_n1246_n3888# 0.340971f
C80 source.t3 a_n1246_n3888# 3.54007f
C81 source.n7 a_n1246_n3888# 2.06796f
C82 source.t12 a_n1246_n3888# 3.54006f
C83 source.n8 a_n1246_n3888# 2.06796f
C84 source.t10 a_n1246_n3888# 0.315891f
C85 source.t11 a_n1246_n3888# 0.315891f
C86 source.n9 a_n1246_n3888# 2.77483f
C87 source.n10 a_n1246_n3888# 0.340975f
C88 source.t7 a_n1246_n3888# 3.54006f
C89 source.n11 a_n1246_n3888# 0.438372f
C90 source.t2 a_n1246_n3888# 3.54006f
C91 source.n12 a_n1246_n3888# 0.438372f
C92 source.t5 a_n1246_n3888# 0.315891f
C93 source.t0 a_n1246_n3888# 0.315891f
C94 source.n13 a_n1246_n3888# 2.77483f
C95 source.n14 a_n1246_n3888# 0.340975f
C96 source.t1 a_n1246_n3888# 3.54006f
C97 source.n15 a_n1246_n3888# 0.582875f
C98 source.n16 a_n1246_n3888# 1.94425f
C99 plus.n0 a_n1246_n3888# 0.132684f
C100 plus.t7 a_n1246_n3888# 0.515732f
C101 plus.t3 a_n1246_n3888# 0.515732f
C102 plus.t4 a_n1246_n3888# 0.520115f
C103 plus.n1 a_n1246_n3888# 0.221213f
C104 plus.n2 a_n1246_n3888# 0.204358f
C105 plus.n3 a_n1246_n3888# 0.021342f
C106 plus.n4 a_n1246_n3888# 0.204358f
C107 plus.t5 a_n1246_n3888# 0.520115f
C108 plus.n5 a_n1246_n3888# 0.221129f
C109 plus.n6 a_n1246_n3888# 0.761948f
C110 plus.n7 a_n1246_n3888# 0.132684f
C111 plus.t6 a_n1246_n3888# 0.520115f
C112 plus.t0 a_n1246_n3888# 0.515732f
C113 plus.t2 a_n1246_n3888# 0.515732f
C114 plus.t1 a_n1246_n3888# 0.520115f
C115 plus.n8 a_n1246_n3888# 0.221213f
C116 plus.n9 a_n1246_n3888# 0.204358f
C117 plus.n10 a_n1246_n3888# 0.021342f
C118 plus.n11 a_n1246_n3888# 0.204358f
C119 plus.n12 a_n1246_n3888# 0.221129f
C120 plus.n13 a_n1246_n3888# 1.74728f
.ends

