* NGSPICE file created from diffpair499.ext - technology: sky130A

.subckt diffpair499 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t26 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t22 plus.t1 source.t43 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X2 drain_left.t21 plus.t2 source.t41 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X3 source.t24 plus.t3 drain_left.t20 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X4 drain_right.t23 minus.t0 source.t15 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 drain_right.t22 minus.t1 source.t21 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 source.t39 plus.t4 drain_left.t19 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X7 a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X8 source.t19 minus.t2 drain_right.t21 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X9 a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X10 source.t31 plus.t5 drain_left.t18 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X11 drain_left.t17 plus.t6 source.t40 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X12 source.t18 minus.t3 drain_right.t20 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X13 source.t17 minus.t4 drain_right.t19 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X14 source.t22 minus.t5 drain_right.t18 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X15 source.t2 minus.t6 drain_right.t17 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X16 source.t5 minus.t7 drain_right.t16 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X17 drain_left.t16 plus.t7 source.t32 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X18 source.t8 minus.t8 drain_right.t15 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X19 drain_right.t14 minus.t9 source.t11 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X20 drain_right.t13 minus.t10 source.t16 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X21 drain_left.t15 plus.t8 source.t38 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X22 source.t36 plus.t9 drain_left.t14 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X23 a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X24 drain_right.t12 minus.t11 source.t0 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X25 drain_right.t11 minus.t12 source.t14 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X26 drain_right.t10 minus.t13 source.t1 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X27 drain_right.t9 minus.t14 source.t23 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X28 drain_right.t8 minus.t15 source.t13 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X29 drain_right.t7 minus.t16 source.t3 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X30 source.t4 minus.t17 drain_right.t6 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X31 drain_right.t5 minus.t18 source.t6 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X32 drain_right.t4 minus.t19 source.t9 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X33 source.t12 minus.t20 drain_right.t3 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X34 source.t28 plus.t10 drain_left.t13 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X35 source.t20 minus.t21 drain_right.t2 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X36 source.t33 plus.t11 drain_left.t12 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X37 drain_left.t11 plus.t12 source.t45 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X38 source.t35 plus.t13 drain_left.t10 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X39 drain_left.t9 plus.t14 source.t30 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X40 a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X41 source.t7 minus.t22 drain_right.t1 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X42 source.t10 minus.t23 drain_right.t0 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X43 source.t37 plus.t15 drain_left.t8 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X44 drain_left.t7 plus.t16 source.t42 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X45 source.t47 plus.t17 drain_left.t6 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X46 source.t34 plus.t18 drain_left.t5 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X47 drain_left.t4 plus.t19 source.t44 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X48 source.t46 plus.t20 drain_left.t3 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X49 drain_left.t2 plus.t21 source.t25 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X50 source.t27 plus.t22 drain_left.t1 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X51 drain_left.t0 plus.t23 source.t29 a_n2094_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n6 plus.t9 2024.77
R1 plus.n29 plus.t19 2024.77
R2 plus.n37 plus.t2 2024.77
R3 plus.n60 plus.t20 2024.77
R4 plus.n7 plus.t6 1964.15
R5 plus.n5 plus.t22 1964.15
R6 plus.n12 plus.t14 1964.15
R7 plus.n14 plus.t13 1964.15
R8 plus.n3 plus.t8 1964.15
R9 plus.n19 plus.t5 1964.15
R10 plus.n21 plus.t21 1964.15
R11 plus.n1 plus.t11 1964.15
R12 plus.n26 plus.t7 1964.15
R13 plus.n28 plus.t3 1964.15
R14 plus.n38 plus.t4 1964.15
R15 plus.n36 plus.t1 1964.15
R16 plus.n43 plus.t17 1964.15
R17 plus.n45 plus.t0 1964.15
R18 plus.n34 plus.t18 1964.15
R19 plus.n50 plus.t23 1964.15
R20 plus.n52 plus.t15 1964.15
R21 plus.n32 plus.t12 1964.15
R22 plus.n57 plus.t10 1964.15
R23 plus.n59 plus.t16 1964.15
R24 plus.n9 plus.n6 161.489
R25 plus.n40 plus.n37 161.489
R26 plus.n9 plus.n8 161.3
R27 plus.n11 plus.n10 161.3
R28 plus.n13 plus.n4 161.3
R29 plus.n16 plus.n15 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n2 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n0 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n40 plus.n39 161.3
R37 plus.n42 plus.n41 161.3
R38 plus.n44 plus.n35 161.3
R39 plus.n47 plus.n46 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n33 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n31 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n8 plus.n7 56.2338
R47 plus.n28 plus.n27 56.2338
R48 plus.n59 plus.n58 56.2338
R49 plus.n39 plus.n38 56.2338
R50 plus.n11 plus.n5 51.852
R51 plus.n26 plus.n25 51.852
R52 plus.n57 plus.n56 51.852
R53 plus.n42 plus.n36 51.852
R54 plus.n13 plus.n12 47.4702
R55 plus.n22 plus.n1 47.4702
R56 plus.n53 plus.n32 47.4702
R57 plus.n44 plus.n43 47.4702
R58 plus.n15 plus.n14 43.0884
R59 plus.n21 plus.n20 43.0884
R60 plus.n52 plus.n51 43.0884
R61 plus.n46 plus.n45 43.0884
R62 plus.n18 plus.n3 38.7066
R63 plus.n19 plus.n18 38.7066
R64 plus.n50 plus.n49 38.7066
R65 plus.n49 plus.n34 38.7066
R66 plus.n15 plus.n3 34.3247
R67 plus.n20 plus.n19 34.3247
R68 plus.n51 plus.n50 34.3247
R69 plus.n46 plus.n34 34.3247
R70 plus plus.n61 32.0596
R71 plus.n14 plus.n13 29.9429
R72 plus.n22 plus.n21 29.9429
R73 plus.n53 plus.n52 29.9429
R74 plus.n45 plus.n44 29.9429
R75 plus.n12 plus.n11 25.5611
R76 plus.n25 plus.n1 25.5611
R77 plus.n56 plus.n32 25.5611
R78 plus.n43 plus.n42 25.5611
R79 plus.n8 plus.n5 21.1793
R80 plus.n27 plus.n26 21.1793
R81 plus.n58 plus.n57 21.1793
R82 plus.n39 plus.n36 21.1793
R83 plus.n7 plus.n6 16.7975
R84 plus.n29 plus.n28 16.7975
R85 plus.n60 plus.n59 16.7975
R86 plus.n38 plus.n37 16.7975
R87 plus plus.n30 13.2694
R88 plus.n10 plus.n9 0.189894
R89 plus.n10 plus.n4 0.189894
R90 plus.n16 plus.n4 0.189894
R91 plus.n17 plus.n16 0.189894
R92 plus.n17 plus.n2 0.189894
R93 plus.n23 plus.n2 0.189894
R94 plus.n24 plus.n23 0.189894
R95 plus.n24 plus.n0 0.189894
R96 plus.n30 plus.n0 0.189894
R97 plus.n61 plus.n31 0.189894
R98 plus.n55 plus.n31 0.189894
R99 plus.n55 plus.n54 0.189894
R100 plus.n54 plus.n33 0.189894
R101 plus.n48 plus.n33 0.189894
R102 plus.n48 plus.n47 0.189894
R103 plus.n47 plus.n35 0.189894
R104 plus.n41 plus.n35 0.189894
R105 plus.n41 plus.n40 0.189894
R106 source.n11 source.t36 45.521
R107 source.n12 source.t6 45.521
R108 source.n23 source.t19 45.521
R109 source.n47 source.t16 45.5208
R110 source.n36 source.t5 45.5208
R111 source.n35 source.t41 45.5208
R112 source.n24 source.t46 45.5208
R113 source.n0 source.t44 45.5208
R114 source.n2 source.n1 44.201
R115 source.n4 source.n3 44.201
R116 source.n6 source.n5 44.201
R117 source.n8 source.n7 44.201
R118 source.n10 source.n9 44.201
R119 source.n14 source.n13 44.201
R120 source.n16 source.n15 44.201
R121 source.n18 source.n17 44.201
R122 source.n20 source.n19 44.201
R123 source.n22 source.n21 44.201
R124 source.n46 source.n45 44.2008
R125 source.n44 source.n43 44.2008
R126 source.n42 source.n41 44.2008
R127 source.n40 source.n39 44.2008
R128 source.n38 source.n37 44.2008
R129 source.n34 source.n33 44.2008
R130 source.n32 source.n31 44.2008
R131 source.n30 source.n29 44.2008
R132 source.n28 source.n27 44.2008
R133 source.n26 source.n25 44.2008
R134 source.n24 source.n23 24.0173
R135 source.n48 source.n0 18.526
R136 source.n48 source.n47 5.49188
R137 source.n45 source.t0 1.3205
R138 source.n45 source.t18 1.3205
R139 source.n43 source.t23 1.3205
R140 source.n43 source.t4 1.3205
R141 source.n41 source.t13 1.3205
R142 source.n41 source.t12 1.3205
R143 source.n39 source.t14 1.3205
R144 source.n39 source.t20 1.3205
R145 source.n37 source.t1 1.3205
R146 source.n37 source.t22 1.3205
R147 source.n33 source.t43 1.3205
R148 source.n33 source.t39 1.3205
R149 source.n31 source.t26 1.3205
R150 source.n31 source.t47 1.3205
R151 source.n29 source.t29 1.3205
R152 source.n29 source.t34 1.3205
R153 source.n27 source.t45 1.3205
R154 source.n27 source.t37 1.3205
R155 source.n25 source.t42 1.3205
R156 source.n25 source.t28 1.3205
R157 source.n1 source.t32 1.3205
R158 source.n1 source.t24 1.3205
R159 source.n3 source.t25 1.3205
R160 source.n3 source.t33 1.3205
R161 source.n5 source.t38 1.3205
R162 source.n5 source.t31 1.3205
R163 source.n7 source.t30 1.3205
R164 source.n7 source.t35 1.3205
R165 source.n9 source.t40 1.3205
R166 source.n9 source.t27 1.3205
R167 source.n13 source.t15 1.3205
R168 source.n13 source.t2 1.3205
R169 source.n15 source.t9 1.3205
R170 source.n15 source.t7 1.3205
R171 source.n17 source.t21 1.3205
R172 source.n17 source.t17 1.3205
R173 source.n19 source.t3 1.3205
R174 source.n19 source.t10 1.3205
R175 source.n21 source.t11 1.3205
R176 source.n21 source.t8 1.3205
R177 source.n12 source.n11 0.470328
R178 source.n36 source.n35 0.470328
R179 source.n23 source.n22 0.457397
R180 source.n22 source.n20 0.457397
R181 source.n20 source.n18 0.457397
R182 source.n18 source.n16 0.457397
R183 source.n16 source.n14 0.457397
R184 source.n14 source.n12 0.457397
R185 source.n11 source.n10 0.457397
R186 source.n10 source.n8 0.457397
R187 source.n8 source.n6 0.457397
R188 source.n6 source.n4 0.457397
R189 source.n4 source.n2 0.457397
R190 source.n2 source.n0 0.457397
R191 source.n26 source.n24 0.457397
R192 source.n28 source.n26 0.457397
R193 source.n30 source.n28 0.457397
R194 source.n32 source.n30 0.457397
R195 source.n34 source.n32 0.457397
R196 source.n35 source.n34 0.457397
R197 source.n38 source.n36 0.457397
R198 source.n40 source.n38 0.457397
R199 source.n42 source.n40 0.457397
R200 source.n44 source.n42 0.457397
R201 source.n46 source.n44 0.457397
R202 source.n47 source.n46 0.457397
R203 source source.n48 0.188
R204 drain_left.n13 drain_left.n11 61.3367
R205 drain_left.n7 drain_left.n5 61.3365
R206 drain_left.n2 drain_left.n0 61.3365
R207 drain_left.n19 drain_left.n18 60.8798
R208 drain_left.n17 drain_left.n16 60.8798
R209 drain_left.n15 drain_left.n14 60.8798
R210 drain_left.n13 drain_left.n12 60.8798
R211 drain_left.n21 drain_left.n20 60.8796
R212 drain_left.n7 drain_left.n6 60.8796
R213 drain_left.n9 drain_left.n8 60.8796
R214 drain_left.n4 drain_left.n3 60.8796
R215 drain_left.n2 drain_left.n1 60.8796
R216 drain_left drain_left.n10 33.9803
R217 drain_left drain_left.n21 6.11011
R218 drain_left.n5 drain_left.t19 1.3205
R219 drain_left.n5 drain_left.t21 1.3205
R220 drain_left.n6 drain_left.t6 1.3205
R221 drain_left.n6 drain_left.t22 1.3205
R222 drain_left.n8 drain_left.t5 1.3205
R223 drain_left.n8 drain_left.t23 1.3205
R224 drain_left.n3 drain_left.t8 1.3205
R225 drain_left.n3 drain_left.t0 1.3205
R226 drain_left.n1 drain_left.t13 1.3205
R227 drain_left.n1 drain_left.t11 1.3205
R228 drain_left.n0 drain_left.t3 1.3205
R229 drain_left.n0 drain_left.t7 1.3205
R230 drain_left.n20 drain_left.t20 1.3205
R231 drain_left.n20 drain_left.t4 1.3205
R232 drain_left.n18 drain_left.t12 1.3205
R233 drain_left.n18 drain_left.t16 1.3205
R234 drain_left.n16 drain_left.t18 1.3205
R235 drain_left.n16 drain_left.t2 1.3205
R236 drain_left.n14 drain_left.t10 1.3205
R237 drain_left.n14 drain_left.t15 1.3205
R238 drain_left.n12 drain_left.t1 1.3205
R239 drain_left.n12 drain_left.t9 1.3205
R240 drain_left.n11 drain_left.t14 1.3205
R241 drain_left.n11 drain_left.t17 1.3205
R242 drain_left.n9 drain_left.n7 0.457397
R243 drain_left.n4 drain_left.n2 0.457397
R244 drain_left.n15 drain_left.n13 0.457397
R245 drain_left.n17 drain_left.n15 0.457397
R246 drain_left.n19 drain_left.n17 0.457397
R247 drain_left.n21 drain_left.n19 0.457397
R248 drain_left.n10 drain_left.n9 0.173602
R249 drain_left.n10 drain_left.n4 0.173602
R250 minus.n29 minus.t2 2024.77
R251 minus.n6 minus.t18 2024.77
R252 minus.n60 minus.t10 2024.77
R253 minus.n37 minus.t7 2024.77
R254 minus.n28 minus.t9 1964.15
R255 minus.n26 minus.t8 1964.15
R256 minus.n1 minus.t16 1964.15
R257 minus.n21 minus.t23 1964.15
R258 minus.n19 minus.t1 1964.15
R259 minus.n3 minus.t4 1964.15
R260 minus.n14 minus.t19 1964.15
R261 minus.n12 minus.t22 1964.15
R262 minus.n5 minus.t0 1964.15
R263 minus.n7 minus.t6 1964.15
R264 minus.n59 minus.t3 1964.15
R265 minus.n57 minus.t11 1964.15
R266 minus.n32 minus.t17 1964.15
R267 minus.n52 minus.t14 1964.15
R268 minus.n50 minus.t20 1964.15
R269 minus.n34 minus.t15 1964.15
R270 minus.n45 minus.t21 1964.15
R271 minus.n43 minus.t12 1964.15
R272 minus.n36 minus.t5 1964.15
R273 minus.n38 minus.t13 1964.15
R274 minus.n9 minus.n6 161.489
R275 minus.n40 minus.n37 161.489
R276 minus.n30 minus.n29 161.3
R277 minus.n27 minus.n0 161.3
R278 minus.n25 minus.n24 161.3
R279 minus.n23 minus.n22 161.3
R280 minus.n20 minus.n2 161.3
R281 minus.n18 minus.n17 161.3
R282 minus.n16 minus.n15 161.3
R283 minus.n13 minus.n4 161.3
R284 minus.n11 minus.n10 161.3
R285 minus.n9 minus.n8 161.3
R286 minus.n61 minus.n60 161.3
R287 minus.n58 minus.n31 161.3
R288 minus.n56 minus.n55 161.3
R289 minus.n54 minus.n53 161.3
R290 minus.n51 minus.n33 161.3
R291 minus.n49 minus.n48 161.3
R292 minus.n47 minus.n46 161.3
R293 minus.n44 minus.n35 161.3
R294 minus.n42 minus.n41 161.3
R295 minus.n40 minus.n39 161.3
R296 minus.n28 minus.n27 56.2338
R297 minus.n8 minus.n7 56.2338
R298 minus.n39 minus.n38 56.2338
R299 minus.n59 minus.n58 56.2338
R300 minus.n26 minus.n25 51.852
R301 minus.n11 minus.n5 51.852
R302 minus.n42 minus.n36 51.852
R303 minus.n57 minus.n56 51.852
R304 minus.n22 minus.n1 47.4702
R305 minus.n13 minus.n12 47.4702
R306 minus.n44 minus.n43 47.4702
R307 minus.n53 minus.n32 47.4702
R308 minus.n21 minus.n20 43.0884
R309 minus.n15 minus.n14 43.0884
R310 minus.n46 minus.n45 43.0884
R311 minus.n52 minus.n51 43.0884
R312 minus.n62 minus.n30 39.3149
R313 minus.n19 minus.n18 38.7066
R314 minus.n18 minus.n3 38.7066
R315 minus.n49 minus.n34 38.7066
R316 minus.n50 minus.n49 38.7066
R317 minus.n20 minus.n19 34.3247
R318 minus.n15 minus.n3 34.3247
R319 minus.n46 minus.n34 34.3247
R320 minus.n51 minus.n50 34.3247
R321 minus.n22 minus.n21 29.9429
R322 minus.n14 minus.n13 29.9429
R323 minus.n45 minus.n44 29.9429
R324 minus.n53 minus.n52 29.9429
R325 minus.n25 minus.n1 25.5611
R326 minus.n12 minus.n11 25.5611
R327 minus.n43 minus.n42 25.5611
R328 minus.n56 minus.n32 25.5611
R329 minus.n27 minus.n26 21.1793
R330 minus.n8 minus.n5 21.1793
R331 minus.n39 minus.n36 21.1793
R332 minus.n58 minus.n57 21.1793
R333 minus.n29 minus.n28 16.7975
R334 minus.n7 minus.n6 16.7975
R335 minus.n38 minus.n37 16.7975
R336 minus.n60 minus.n59 16.7975
R337 minus.n62 minus.n61 6.48914
R338 minus.n30 minus.n0 0.189894
R339 minus.n24 minus.n0 0.189894
R340 minus.n24 minus.n23 0.189894
R341 minus.n23 minus.n2 0.189894
R342 minus.n17 minus.n2 0.189894
R343 minus.n17 minus.n16 0.189894
R344 minus.n16 minus.n4 0.189894
R345 minus.n10 minus.n4 0.189894
R346 minus.n10 minus.n9 0.189894
R347 minus.n41 minus.n40 0.189894
R348 minus.n41 minus.n35 0.189894
R349 minus.n47 minus.n35 0.189894
R350 minus.n48 minus.n47 0.189894
R351 minus.n48 minus.n33 0.189894
R352 minus.n54 minus.n33 0.189894
R353 minus.n55 minus.n54 0.189894
R354 minus.n55 minus.n31 0.189894
R355 minus.n61 minus.n31 0.189894
R356 minus minus.n62 0.188
R357 drain_right.n13 drain_right.n11 61.3365
R358 drain_right.n7 drain_right.n5 61.3365
R359 drain_right.n2 drain_right.n0 61.3365
R360 drain_right.n13 drain_right.n12 60.8798
R361 drain_right.n15 drain_right.n14 60.8798
R362 drain_right.n17 drain_right.n16 60.8798
R363 drain_right.n19 drain_right.n18 60.8798
R364 drain_right.n21 drain_right.n20 60.8798
R365 drain_right.n7 drain_right.n6 60.8796
R366 drain_right.n9 drain_right.n8 60.8796
R367 drain_right.n4 drain_right.n3 60.8796
R368 drain_right.n2 drain_right.n1 60.8796
R369 drain_right drain_right.n10 33.4271
R370 drain_right drain_right.n21 6.11011
R371 drain_right.n5 drain_right.t20 1.3205
R372 drain_right.n5 drain_right.t13 1.3205
R373 drain_right.n6 drain_right.t6 1.3205
R374 drain_right.n6 drain_right.t12 1.3205
R375 drain_right.n8 drain_right.t3 1.3205
R376 drain_right.n8 drain_right.t9 1.3205
R377 drain_right.n3 drain_right.t2 1.3205
R378 drain_right.n3 drain_right.t8 1.3205
R379 drain_right.n1 drain_right.t18 1.3205
R380 drain_right.n1 drain_right.t11 1.3205
R381 drain_right.n0 drain_right.t16 1.3205
R382 drain_right.n0 drain_right.t10 1.3205
R383 drain_right.n11 drain_right.t17 1.3205
R384 drain_right.n11 drain_right.t5 1.3205
R385 drain_right.n12 drain_right.t1 1.3205
R386 drain_right.n12 drain_right.t23 1.3205
R387 drain_right.n14 drain_right.t19 1.3205
R388 drain_right.n14 drain_right.t4 1.3205
R389 drain_right.n16 drain_right.t0 1.3205
R390 drain_right.n16 drain_right.t22 1.3205
R391 drain_right.n18 drain_right.t15 1.3205
R392 drain_right.n18 drain_right.t7 1.3205
R393 drain_right.n20 drain_right.t21 1.3205
R394 drain_right.n20 drain_right.t14 1.3205
R395 drain_right.n9 drain_right.n7 0.457397
R396 drain_right.n4 drain_right.n2 0.457397
R397 drain_right.n21 drain_right.n19 0.457397
R398 drain_right.n19 drain_right.n17 0.457397
R399 drain_right.n17 drain_right.n15 0.457397
R400 drain_right.n15 drain_right.n13 0.457397
R401 drain_right.n10 drain_right.n9 0.173602
R402 drain_right.n10 drain_right.n4 0.173602
C0 drain_left plus 7.81812f
C1 drain_right drain_left 1.11966f
C2 source minus 7.16396f
C3 drain_right plus 0.359911f
C4 source drain_left 66.239204f
C5 minus drain_left 0.171754f
C6 source plus 7.178f
C7 minus plus 6.32167f
C8 source drain_right 66.2395f
C9 drain_right minus 7.61297f
C10 drain_right a_n2094_n3888# 8.19267f
C11 drain_left a_n2094_n3888# 8.52024f
C12 source a_n2094_n3888# 10.276295f
C13 minus a_n2094_n3888# 8.352074f
C14 plus a_n2094_n3888# 10.67135f
C15 drain_right.t16 a_n2094_n3888# 0.465539f
C16 drain_right.t10 a_n2094_n3888# 0.465539f
C17 drain_right.n0 a_n2094_n3888# 4.21131f
C18 drain_right.t18 a_n2094_n3888# 0.465539f
C19 drain_right.t11 a_n2094_n3888# 0.465539f
C20 drain_right.n1 a_n2094_n3888# 4.20793f
C21 drain_right.n2 a_n2094_n3888# 0.887092f
C22 drain_right.t2 a_n2094_n3888# 0.465539f
C23 drain_right.t8 a_n2094_n3888# 0.465539f
C24 drain_right.n3 a_n2094_n3888# 4.20793f
C25 drain_right.n4 a_n2094_n3888# 0.40667f
C26 drain_right.t20 a_n2094_n3888# 0.465539f
C27 drain_right.t13 a_n2094_n3888# 0.465539f
C28 drain_right.n5 a_n2094_n3888# 4.21131f
C29 drain_right.t6 a_n2094_n3888# 0.465539f
C30 drain_right.t12 a_n2094_n3888# 0.465539f
C31 drain_right.n6 a_n2094_n3888# 4.20793f
C32 drain_right.n7 a_n2094_n3888# 0.887092f
C33 drain_right.t3 a_n2094_n3888# 0.465539f
C34 drain_right.t9 a_n2094_n3888# 0.465539f
C35 drain_right.n8 a_n2094_n3888# 4.20793f
C36 drain_right.n9 a_n2094_n3888# 0.40667f
C37 drain_right.n10 a_n2094_n3888# 2.21312f
C38 drain_right.t17 a_n2094_n3888# 0.465539f
C39 drain_right.t5 a_n2094_n3888# 0.465539f
C40 drain_right.n11 a_n2094_n3888# 4.2113f
C41 drain_right.t1 a_n2094_n3888# 0.465539f
C42 drain_right.t23 a_n2094_n3888# 0.465539f
C43 drain_right.n12 a_n2094_n3888# 4.20794f
C44 drain_right.n13 a_n2094_n3888# 0.8871f
C45 drain_right.t19 a_n2094_n3888# 0.465539f
C46 drain_right.t4 a_n2094_n3888# 0.465539f
C47 drain_right.n14 a_n2094_n3888# 4.20794f
C48 drain_right.n15 a_n2094_n3888# 0.437321f
C49 drain_right.t0 a_n2094_n3888# 0.465539f
C50 drain_right.t22 a_n2094_n3888# 0.465539f
C51 drain_right.n16 a_n2094_n3888# 4.20794f
C52 drain_right.n17 a_n2094_n3888# 0.437321f
C53 drain_right.t15 a_n2094_n3888# 0.465539f
C54 drain_right.t7 a_n2094_n3888# 0.465539f
C55 drain_right.n18 a_n2094_n3888# 4.20794f
C56 drain_right.n19 a_n2094_n3888# 0.437321f
C57 drain_right.t21 a_n2094_n3888# 0.465539f
C58 drain_right.t14 a_n2094_n3888# 0.465539f
C59 drain_right.n20 a_n2094_n3888# 4.20794f
C60 drain_right.n21 a_n2094_n3888# 0.758746f
C61 minus.n0 a_n2094_n3888# 0.051736f
C62 minus.t2 a_n2094_n3888# 0.443167f
C63 minus.t9 a_n2094_n3888# 0.437863f
C64 minus.t8 a_n2094_n3888# 0.437863f
C65 minus.t16 a_n2094_n3888# 0.437863f
C66 minus.n1 a_n2094_n3888# 0.173502f
C67 minus.n2 a_n2094_n3888# 0.051736f
C68 minus.t23 a_n2094_n3888# 0.437863f
C69 minus.t1 a_n2094_n3888# 0.437863f
C70 minus.t4 a_n2094_n3888# 0.437863f
C71 minus.n3 a_n2094_n3888# 0.173502f
C72 minus.n4 a_n2094_n3888# 0.051736f
C73 minus.t19 a_n2094_n3888# 0.437863f
C74 minus.t22 a_n2094_n3888# 0.437863f
C75 minus.t0 a_n2094_n3888# 0.437863f
C76 minus.n5 a_n2094_n3888# 0.173502f
C77 minus.t18 a_n2094_n3888# 0.443167f
C78 minus.n6 a_n2094_n3888# 0.190066f
C79 minus.t6 a_n2094_n3888# 0.437863f
C80 minus.n7 a_n2094_n3888# 0.173502f
C81 minus.n8 a_n2094_n3888# 0.018119f
C82 minus.n9 a_n2094_n3888# 0.120297f
C83 minus.n10 a_n2094_n3888# 0.051736f
C84 minus.n11 a_n2094_n3888# 0.018119f
C85 minus.n12 a_n2094_n3888# 0.173502f
C86 minus.n13 a_n2094_n3888# 0.018119f
C87 minus.n14 a_n2094_n3888# 0.173502f
C88 minus.n15 a_n2094_n3888# 0.018119f
C89 minus.n16 a_n2094_n3888# 0.051736f
C90 minus.n17 a_n2094_n3888# 0.051736f
C91 minus.n18 a_n2094_n3888# 0.018119f
C92 minus.n19 a_n2094_n3888# 0.173502f
C93 minus.n20 a_n2094_n3888# 0.018119f
C94 minus.n21 a_n2094_n3888# 0.173502f
C95 minus.n22 a_n2094_n3888# 0.018119f
C96 minus.n23 a_n2094_n3888# 0.051736f
C97 minus.n24 a_n2094_n3888# 0.051736f
C98 minus.n25 a_n2094_n3888# 0.018119f
C99 minus.n26 a_n2094_n3888# 0.173502f
C100 minus.n27 a_n2094_n3888# 0.018119f
C101 minus.n28 a_n2094_n3888# 0.173502f
C102 minus.n29 a_n2094_n3888# 0.189986f
C103 minus.n30 a_n2094_n3888# 2.07581f
C104 minus.n31 a_n2094_n3888# 0.051736f
C105 minus.t3 a_n2094_n3888# 0.437863f
C106 minus.t11 a_n2094_n3888# 0.437863f
C107 minus.t17 a_n2094_n3888# 0.437863f
C108 minus.n32 a_n2094_n3888# 0.173502f
C109 minus.n33 a_n2094_n3888# 0.051736f
C110 minus.t14 a_n2094_n3888# 0.437863f
C111 minus.t20 a_n2094_n3888# 0.437863f
C112 minus.t15 a_n2094_n3888# 0.437863f
C113 minus.n34 a_n2094_n3888# 0.173502f
C114 minus.n35 a_n2094_n3888# 0.051736f
C115 minus.t21 a_n2094_n3888# 0.437863f
C116 minus.t12 a_n2094_n3888# 0.437863f
C117 minus.t5 a_n2094_n3888# 0.437863f
C118 minus.n36 a_n2094_n3888# 0.173502f
C119 minus.t7 a_n2094_n3888# 0.443167f
C120 minus.n37 a_n2094_n3888# 0.190066f
C121 minus.t13 a_n2094_n3888# 0.437863f
C122 minus.n38 a_n2094_n3888# 0.173502f
C123 minus.n39 a_n2094_n3888# 0.018119f
C124 minus.n40 a_n2094_n3888# 0.120297f
C125 minus.n41 a_n2094_n3888# 0.051736f
C126 minus.n42 a_n2094_n3888# 0.018119f
C127 minus.n43 a_n2094_n3888# 0.173502f
C128 minus.n44 a_n2094_n3888# 0.018119f
C129 minus.n45 a_n2094_n3888# 0.173502f
C130 minus.n46 a_n2094_n3888# 0.018119f
C131 minus.n47 a_n2094_n3888# 0.051736f
C132 minus.n48 a_n2094_n3888# 0.051736f
C133 minus.n49 a_n2094_n3888# 0.018119f
C134 minus.n50 a_n2094_n3888# 0.173502f
C135 minus.n51 a_n2094_n3888# 0.018119f
C136 minus.n52 a_n2094_n3888# 0.173502f
C137 minus.n53 a_n2094_n3888# 0.018119f
C138 minus.n54 a_n2094_n3888# 0.051736f
C139 minus.n55 a_n2094_n3888# 0.051736f
C140 minus.n56 a_n2094_n3888# 0.018119f
C141 minus.n57 a_n2094_n3888# 0.173502f
C142 minus.n58 a_n2094_n3888# 0.018119f
C143 minus.n59 a_n2094_n3888# 0.173502f
C144 minus.t10 a_n2094_n3888# 0.443167f
C145 minus.n60 a_n2094_n3888# 0.189986f
C146 minus.n61 a_n2094_n3888# 0.33691f
C147 minus.n62 a_n2094_n3888# 2.49871f
C148 drain_left.t3 a_n2094_n3888# 0.465831f
C149 drain_left.t7 a_n2094_n3888# 0.465831f
C150 drain_left.n0 a_n2094_n3888# 4.21395f
C151 drain_left.t13 a_n2094_n3888# 0.465831f
C152 drain_left.t11 a_n2094_n3888# 0.465831f
C153 drain_left.n1 a_n2094_n3888# 4.21057f
C154 drain_left.n2 a_n2094_n3888# 0.887649f
C155 drain_left.t8 a_n2094_n3888# 0.465831f
C156 drain_left.t0 a_n2094_n3888# 0.465831f
C157 drain_left.n3 a_n2094_n3888# 4.21057f
C158 drain_left.n4 a_n2094_n3888# 0.406925f
C159 drain_left.t19 a_n2094_n3888# 0.465831f
C160 drain_left.t21 a_n2094_n3888# 0.465831f
C161 drain_left.n5 a_n2094_n3888# 4.21395f
C162 drain_left.t6 a_n2094_n3888# 0.465831f
C163 drain_left.t22 a_n2094_n3888# 0.465831f
C164 drain_left.n6 a_n2094_n3888# 4.21057f
C165 drain_left.n7 a_n2094_n3888# 0.887649f
C166 drain_left.t5 a_n2094_n3888# 0.465831f
C167 drain_left.t23 a_n2094_n3888# 0.465831f
C168 drain_left.n8 a_n2094_n3888# 4.21057f
C169 drain_left.n9 a_n2094_n3888# 0.406925f
C170 drain_left.n10 a_n2094_n3888# 2.29594f
C171 drain_left.t14 a_n2094_n3888# 0.465831f
C172 drain_left.t17 a_n2094_n3888# 0.465831f
C173 drain_left.n11 a_n2094_n3888# 4.21395f
C174 drain_left.t1 a_n2094_n3888# 0.465831f
C175 drain_left.t9 a_n2094_n3888# 0.465831f
C176 drain_left.n12 a_n2094_n3888# 4.21057f
C177 drain_left.n13 a_n2094_n3888# 0.887642f
C178 drain_left.t10 a_n2094_n3888# 0.465831f
C179 drain_left.t15 a_n2094_n3888# 0.465831f
C180 drain_left.n14 a_n2094_n3888# 4.21057f
C181 drain_left.n15 a_n2094_n3888# 0.437595f
C182 drain_left.t18 a_n2094_n3888# 0.465831f
C183 drain_left.t2 a_n2094_n3888# 0.465831f
C184 drain_left.n16 a_n2094_n3888# 4.21057f
C185 drain_left.n17 a_n2094_n3888# 0.437595f
C186 drain_left.t12 a_n2094_n3888# 0.465831f
C187 drain_left.t16 a_n2094_n3888# 0.465831f
C188 drain_left.n18 a_n2094_n3888# 4.21057f
C189 drain_left.n19 a_n2094_n3888# 0.437595f
C190 drain_left.t20 a_n2094_n3888# 0.465831f
C191 drain_left.t4 a_n2094_n3888# 0.465831f
C192 drain_left.n20 a_n2094_n3888# 4.21056f
C193 drain_left.n21 a_n2094_n3888# 0.759237f
C194 source.t44 a_n2094_n3888# 4.58429f
C195 source.n0 a_n2094_n3888# 2.10789f
C196 source.t32 a_n2094_n3888# 0.40907f
C197 source.t24 a_n2094_n3888# 0.40907f
C198 source.n1 a_n2094_n3888# 3.59334f
C199 source.n2 a_n2094_n3888# 0.441548f
C200 source.t25 a_n2094_n3888# 0.40907f
C201 source.t33 a_n2094_n3888# 0.40907f
C202 source.n3 a_n2094_n3888# 3.59334f
C203 source.n4 a_n2094_n3888# 0.441548f
C204 source.t38 a_n2094_n3888# 0.40907f
C205 source.t31 a_n2094_n3888# 0.40907f
C206 source.n5 a_n2094_n3888# 3.59334f
C207 source.n6 a_n2094_n3888# 0.441548f
C208 source.t30 a_n2094_n3888# 0.40907f
C209 source.t35 a_n2094_n3888# 0.40907f
C210 source.n7 a_n2094_n3888# 3.59334f
C211 source.n8 a_n2094_n3888# 0.441548f
C212 source.t40 a_n2094_n3888# 0.40907f
C213 source.t27 a_n2094_n3888# 0.40907f
C214 source.n9 a_n2094_n3888# 3.59334f
C215 source.n10 a_n2094_n3888# 0.441548f
C216 source.t36 a_n2094_n3888# 4.58429f
C217 source.n11 a_n2094_n3888# 0.567675f
C218 source.t6 a_n2094_n3888# 4.58429f
C219 source.n12 a_n2094_n3888# 0.567675f
C220 source.t15 a_n2094_n3888# 0.40907f
C221 source.t2 a_n2094_n3888# 0.40907f
C222 source.n13 a_n2094_n3888# 3.59334f
C223 source.n14 a_n2094_n3888# 0.441548f
C224 source.t9 a_n2094_n3888# 0.40907f
C225 source.t7 a_n2094_n3888# 0.40907f
C226 source.n15 a_n2094_n3888# 3.59334f
C227 source.n16 a_n2094_n3888# 0.441548f
C228 source.t21 a_n2094_n3888# 0.40907f
C229 source.t17 a_n2094_n3888# 0.40907f
C230 source.n17 a_n2094_n3888# 3.59334f
C231 source.n18 a_n2094_n3888# 0.441548f
C232 source.t3 a_n2094_n3888# 0.40907f
C233 source.t10 a_n2094_n3888# 0.40907f
C234 source.n19 a_n2094_n3888# 3.59334f
C235 source.n20 a_n2094_n3888# 0.441548f
C236 source.t11 a_n2094_n3888# 0.40907f
C237 source.t8 a_n2094_n3888# 0.40907f
C238 source.n21 a_n2094_n3888# 3.59334f
C239 source.n22 a_n2094_n3888# 0.441548f
C240 source.t19 a_n2094_n3888# 4.58429f
C241 source.n23 a_n2094_n3888# 2.67795f
C242 source.t46 a_n2094_n3888# 4.58429f
C243 source.n24 a_n2094_n3888# 2.67795f
C244 source.t42 a_n2094_n3888# 0.40907f
C245 source.t28 a_n2094_n3888# 0.40907f
C246 source.n25 a_n2094_n3888# 3.59333f
C247 source.n26 a_n2094_n3888# 0.441553f
C248 source.t45 a_n2094_n3888# 0.40907f
C249 source.t37 a_n2094_n3888# 0.40907f
C250 source.n27 a_n2094_n3888# 3.59333f
C251 source.n28 a_n2094_n3888# 0.441553f
C252 source.t29 a_n2094_n3888# 0.40907f
C253 source.t34 a_n2094_n3888# 0.40907f
C254 source.n29 a_n2094_n3888# 3.59333f
C255 source.n30 a_n2094_n3888# 0.441553f
C256 source.t26 a_n2094_n3888# 0.40907f
C257 source.t47 a_n2094_n3888# 0.40907f
C258 source.n31 a_n2094_n3888# 3.59333f
C259 source.n32 a_n2094_n3888# 0.441553f
C260 source.t43 a_n2094_n3888# 0.40907f
C261 source.t39 a_n2094_n3888# 0.40907f
C262 source.n33 a_n2094_n3888# 3.59333f
C263 source.n34 a_n2094_n3888# 0.441553f
C264 source.t41 a_n2094_n3888# 4.58429f
C265 source.n35 a_n2094_n3888# 0.56768f
C266 source.t5 a_n2094_n3888# 4.58429f
C267 source.n36 a_n2094_n3888# 0.56768f
C268 source.t1 a_n2094_n3888# 0.40907f
C269 source.t22 a_n2094_n3888# 0.40907f
C270 source.n37 a_n2094_n3888# 3.59333f
C271 source.n38 a_n2094_n3888# 0.441553f
C272 source.t14 a_n2094_n3888# 0.40907f
C273 source.t20 a_n2094_n3888# 0.40907f
C274 source.n39 a_n2094_n3888# 3.59333f
C275 source.n40 a_n2094_n3888# 0.441553f
C276 source.t13 a_n2094_n3888# 0.40907f
C277 source.t12 a_n2094_n3888# 0.40907f
C278 source.n41 a_n2094_n3888# 3.59333f
C279 source.n42 a_n2094_n3888# 0.441553f
C280 source.t23 a_n2094_n3888# 0.40907f
C281 source.t4 a_n2094_n3888# 0.40907f
C282 source.n43 a_n2094_n3888# 3.59333f
C283 source.n44 a_n2094_n3888# 0.441553f
C284 source.t0 a_n2094_n3888# 0.40907f
C285 source.t18 a_n2094_n3888# 0.40907f
C286 source.n45 a_n2094_n3888# 3.59333f
C287 source.n46 a_n2094_n3888# 0.441553f
C288 source.t16 a_n2094_n3888# 4.58429f
C289 source.n47 a_n2094_n3888# 0.754808f
C290 source.n48 a_n2094_n3888# 2.51776f
C291 plus.n0 a_n2094_n3888# 0.052486f
C292 plus.t3 a_n2094_n3888# 0.444216f
C293 plus.t7 a_n2094_n3888# 0.444216f
C294 plus.t11 a_n2094_n3888# 0.444216f
C295 plus.n1 a_n2094_n3888# 0.176019f
C296 plus.n2 a_n2094_n3888# 0.052486f
C297 plus.t21 a_n2094_n3888# 0.444216f
C298 plus.t5 a_n2094_n3888# 0.444216f
C299 plus.t8 a_n2094_n3888# 0.444216f
C300 plus.n3 a_n2094_n3888# 0.176019f
C301 plus.n4 a_n2094_n3888# 0.052486f
C302 plus.t13 a_n2094_n3888# 0.444216f
C303 plus.t14 a_n2094_n3888# 0.444216f
C304 plus.t22 a_n2094_n3888# 0.444216f
C305 plus.n5 a_n2094_n3888# 0.176019f
C306 plus.t9 a_n2094_n3888# 0.449597f
C307 plus.n6 a_n2094_n3888# 0.192824f
C308 plus.t6 a_n2094_n3888# 0.444216f
C309 plus.n7 a_n2094_n3888# 0.176019f
C310 plus.n8 a_n2094_n3888# 0.018382f
C311 plus.n9 a_n2094_n3888# 0.122042f
C312 plus.n10 a_n2094_n3888# 0.052486f
C313 plus.n11 a_n2094_n3888# 0.018382f
C314 plus.n12 a_n2094_n3888# 0.176019f
C315 plus.n13 a_n2094_n3888# 0.018382f
C316 plus.n14 a_n2094_n3888# 0.176019f
C317 plus.n15 a_n2094_n3888# 0.018382f
C318 plus.n16 a_n2094_n3888# 0.052486f
C319 plus.n17 a_n2094_n3888# 0.052486f
C320 plus.n18 a_n2094_n3888# 0.018382f
C321 plus.n19 a_n2094_n3888# 0.176019f
C322 plus.n20 a_n2094_n3888# 0.018382f
C323 plus.n21 a_n2094_n3888# 0.176019f
C324 plus.n22 a_n2094_n3888# 0.018382f
C325 plus.n23 a_n2094_n3888# 0.052486f
C326 plus.n24 a_n2094_n3888# 0.052486f
C327 plus.n25 a_n2094_n3888# 0.018382f
C328 plus.n26 a_n2094_n3888# 0.176019f
C329 plus.n27 a_n2094_n3888# 0.018382f
C330 plus.n28 a_n2094_n3888# 0.176019f
C331 plus.t19 a_n2094_n3888# 0.449597f
C332 plus.n29 a_n2094_n3888# 0.192742f
C333 plus.n30 a_n2094_n3888# 0.661918f
C334 plus.n31 a_n2094_n3888# 0.052486f
C335 plus.t20 a_n2094_n3888# 0.449597f
C336 plus.t16 a_n2094_n3888# 0.444216f
C337 plus.t10 a_n2094_n3888# 0.444216f
C338 plus.t12 a_n2094_n3888# 0.444216f
C339 plus.n32 a_n2094_n3888# 0.176019f
C340 plus.n33 a_n2094_n3888# 0.052486f
C341 plus.t15 a_n2094_n3888# 0.444216f
C342 plus.t23 a_n2094_n3888# 0.444216f
C343 plus.t18 a_n2094_n3888# 0.444216f
C344 plus.n34 a_n2094_n3888# 0.176019f
C345 plus.n35 a_n2094_n3888# 0.052486f
C346 plus.t0 a_n2094_n3888# 0.444216f
C347 plus.t17 a_n2094_n3888# 0.444216f
C348 plus.t1 a_n2094_n3888# 0.444216f
C349 plus.n36 a_n2094_n3888# 0.176019f
C350 plus.t2 a_n2094_n3888# 0.449597f
C351 plus.n37 a_n2094_n3888# 0.192824f
C352 plus.t4 a_n2094_n3888# 0.444216f
C353 plus.n38 a_n2094_n3888# 0.176019f
C354 plus.n39 a_n2094_n3888# 0.018382f
C355 plus.n40 a_n2094_n3888# 0.122042f
C356 plus.n41 a_n2094_n3888# 0.052486f
C357 plus.n42 a_n2094_n3888# 0.018382f
C358 plus.n43 a_n2094_n3888# 0.176019f
C359 plus.n44 a_n2094_n3888# 0.018382f
C360 plus.n45 a_n2094_n3888# 0.176019f
C361 plus.n46 a_n2094_n3888# 0.018382f
C362 plus.n47 a_n2094_n3888# 0.052486f
C363 plus.n48 a_n2094_n3888# 0.052486f
C364 plus.n49 a_n2094_n3888# 0.018382f
C365 plus.n50 a_n2094_n3888# 0.176019f
C366 plus.n51 a_n2094_n3888# 0.018382f
C367 plus.n52 a_n2094_n3888# 0.176019f
C368 plus.n53 a_n2094_n3888# 0.018382f
C369 plus.n54 a_n2094_n3888# 0.052486f
C370 plus.n55 a_n2094_n3888# 0.052486f
C371 plus.n56 a_n2094_n3888# 0.018382f
C372 plus.n57 a_n2094_n3888# 0.176019f
C373 plus.n58 a_n2094_n3888# 0.018382f
C374 plus.n59 a_n2094_n3888# 0.176019f
C375 plus.n60 a_n2094_n3888# 0.192742f
C376 plus.n61 a_n2094_n3888# 1.73726f
.ends

