* NGSPICE file created from diffpair71.ext - technology: sky130A

.subckt diffpair71 minus drain_right drain_left source plus
X0 a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 source.t4 minus.t0 drain_right.t2 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X3 drain_left.t3 plus.t0 source.t0 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X4 source.t3 minus.t1 drain_right.t1 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X5 drain_right.t0 minus.t2 source.t2 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X6 a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X7 drain_right.t3 minus.t3 source.t1 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X8 a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X9 drain_left.t2 plus.t1 source.t7 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X10 source.t6 plus.t2 drain_left.t1 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X11 source.t5 plus.t3 drain_left.t0 a_n1394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n0 minus.t2 100.225
R1 minus.n1 minus.t0 100.225
R2 minus.n0 minus.t1 100.175
R3 minus.n1 minus.t3 100.175
R4 minus.n2 minus.n0 70.9272
R5 minus.n2 minus.n1 51.3591
R6 minus minus.n2 0.188
R7 drain_right drain_right.n0 260.56
R8 drain_right drain_right.n1 246.76
R9 drain_right.n0 drain_right.t2 19.8005
R10 drain_right.n0 drain_right.t3 19.8005
R11 drain_right.n1 drain_right.t1 19.8005
R12 drain_right.n1 drain_right.t0 19.8005
R13 source.n0 source.t7 243.255
R14 source.n1 source.t5 243.255
R15 source.n2 source.t2 243.255
R16 source.n3 source.t3 243.255
R17 source.n7 source.t1 243.254
R18 source.n6 source.t4 243.254
R19 source.n5 source.t0 243.254
R20 source.n4 source.t6 243.254
R21 source.n4 source.n3 13.9285
R22 source.n8 source.n0 8.17853
R23 source.n8 source.n7 5.7505
R24 source.n3 source.n2 0.974638
R25 source.n1 source.n0 0.974638
R26 source.n5 source.n4 0.974638
R27 source.n7 source.n6 0.974638
R28 source.n2 source.n1 0.470328
R29 source.n6 source.n5 0.470328
R30 source source.n8 0.188
R31 plus.n0 plus.t3 100.225
R32 plus.n1 plus.t0 100.225
R33 plus.n0 plus.t1 100.175
R34 plus.n1 plus.t2 100.175
R35 plus plus.n1 68.975
R36 plus plus.n0 52.8363
R37 drain_left drain_left.n0 261.113
R38 drain_left drain_left.n1 246.76
R39 drain_left.n0 drain_left.t1 19.8005
R40 drain_left.n0 drain_left.t3 19.8005
R41 drain_left.n1 drain_left.t0 19.8005
R42 drain_left.n1 drain_left.t2 19.8005
C0 drain_left drain_right 0.588954f
C1 drain_left source 1.99498f
C2 drain_left minus 0.177361f
C3 source drain_right 1.99659f
C4 minus drain_right 0.557449f
C5 source minus 0.777238f
C6 plus drain_left 0.689622f
C7 plus drain_right 0.293504f
C8 plus source 0.791101f
C9 plus minus 2.84471f
C10 drain_right a_n1394_n1088# 1.78962f
C11 drain_left a_n1394_n1088# 1.92686f
C12 source a_n1394_n1088# 2.28974f
C13 minus a_n1394_n1088# 4.309216f
C14 plus a_n1394_n1088# 5.8127f
C15 plus.t1 a_n1394_n1088# 0.117413f
C16 plus.t3 a_n1394_n1088# 0.117482f
C17 plus.n0 a_n1394_n1088# 0.207458f
C18 plus.t0 a_n1394_n1088# 0.117482f
C19 plus.t2 a_n1394_n1088# 0.117413f
C20 plus.n1 a_n1394_n1088# 0.439512f
C21 minus.t2 a_n1394_n1088# 0.114511f
C22 minus.t1 a_n1394_n1088# 0.114444f
C23 minus.n0 a_n1394_n1088# 0.448854f
C24 minus.t0 a_n1394_n1088# 0.114511f
C25 minus.t3 a_n1394_n1088# 0.114444f
C26 minus.n1 a_n1394_n1088# 0.192469f
C27 minus.n2 a_n1394_n1088# 1.67777f
.ends

