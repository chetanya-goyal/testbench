* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.25
X1 a_n948_n1092# a_n948_n1092# a_n948_n1092# a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X2 a_n948_n1092# a_n948_n1092# a_n948_n1092# a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X3 drain_right.t0 minus.t1 source.t3 a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.25
X4 drain_left.t1 plus.t0 source.t0 a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.25
X5 a_n948_n1092# a_n948_n1092# a_n948_n1092# a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X6 a_n948_n1092# a_n948_n1092# a_n948_n1092# a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X7 drain_left.t0 plus.t1 source.t1 a_n948_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.25
R0 minus.n0 minus.t0 431.375
R1 minus.n0 minus.t1 413.481
R2 minus minus.n0 0.188
R3 source.n0 source.t0 243.255
R4 source.n1 source.t2 243.255
R5 source.n3 source.t3 243.254
R6 source.n2 source.t1 243.254
R7 source.n2 source.n1 13.9695
R8 source.n4 source.n0 7.95661
R9 source.n4 source.n3 5.51343
R10 source.n1 source.n0 0.720328
R11 source.n3 source.n2 0.720328
R12 source source.n4 0.188
R13 drain_right drain_right.t0 279.122
R14 drain_right drain_right.t1 265.836
R15 plus plus.t1 429.423
R16 plus plus.t0 414.957
R17 drain_left drain_left.t0 279.675
R18 drain_left drain_left.t1 266.086
C0 source drain_left 1.66641f
C1 source minus 0.375063f
C2 drain_left minus 0.179109f
C3 source plus 0.388982f
C4 drain_right source 1.6659f
C5 drain_left plus 0.414836f
C6 drain_right drain_left 0.417552f
C7 minus plus 2.31518f
C8 drain_right minus 0.329251f
C9 drain_right plus 0.248763f
C10 drain_right a_n948_n1092# 1.54446f
C11 drain_left a_n948_n1092# 1.63914f
C12 source a_n948_n1092# 1.63858f
C13 minus a_n948_n1092# 2.760308f
C14 plus a_n948_n1092# 4.72024f
C15 plus.t0 a_n948_n1092# 0.064216f
C16 plus.t1 a_n948_n1092# 0.102589f
C17 minus.t0 a_n948_n1092# 0.102533f
C18 minus.t1 a_n948_n1092# 0.060239f
C19 minus.n0 a_n948_n1092# 2.10666f
.ends

