* NGSPICE file created from diffpair496.ext - technology: sky130A

.subckt diffpair496 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t25 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t12 plus.t1 source.t14 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X2 drain_left.t11 plus.t2 source.t18 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X3 drain_right.t13 minus.t0 source.t8 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X4 drain_right.t12 minus.t1 source.t4 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X5 source.t17 plus.t3 drain_left.t10 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 drain_left.t9 plus.t4 source.t21 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X7 source.t24 plus.t5 drain_left.t8 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 source.t11 minus.t2 drain_right.t11 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 drain_right.t10 minus.t3 source.t5 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X10 source.t7 minus.t4 drain_right.t9 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X11 drain_right.t8 minus.t5 source.t9 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X12 a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X13 a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X14 source.t20 plus.t6 drain_left.t7 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X15 drain_left.t6 plus.t7 source.t26 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X16 source.t2 minus.t6 drain_right.t7 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X17 source.t0 minus.t7 drain_right.t6 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X18 source.t1 minus.t8 drain_right.t5 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X19 drain_right.t4 minus.t9 source.t3 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X20 drain_right.t3 minus.t10 source.t10 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X21 drain_right.t2 minus.t11 source.t6 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X22 drain_right.t1 minus.t12 source.t12 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X23 a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X24 drain_left.t5 plus.t8 source.t16 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X25 source.t23 plus.t9 drain_left.t4 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X26 source.t13 minus.t13 drain_right.t0 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X27 source.t27 plus.t10 drain_left.t3 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X28 source.t15 plus.t11 drain_left.t2 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X29 a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X30 drain_left.t1 plus.t12 source.t22 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X31 drain_left.t0 plus.t13 source.t19 a_n1564_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n3 plus.t7 2013.81
R1 plus.n14 plus.t4 2013.81
R2 plus.n19 plus.t2 2013.81
R3 plus.n30 plus.t13 2013.81
R4 plus.n4 plus.t5 1964.15
R5 plus.n6 plus.t12 1964.15
R6 plus.n1 plus.t9 1964.15
R7 plus.n11 plus.t8 1964.15
R8 plus.n13 plus.t6 1964.15
R9 plus.n20 plus.t3 1964.15
R10 plus.n22 plus.t1 1964.15
R11 plus.n17 plus.t10 1964.15
R12 plus.n27 plus.t0 1964.15
R13 plus.n29 plus.t11 1964.15
R14 plus.n3 plus.n2 161.489
R15 plus.n19 plus.n18 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n10 plus.n9 161.3
R19 plus.n12 plus.n0 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n21 plus.n18 161.3
R22 plus.n24 plus.n23 161.3
R23 plus.n26 plus.n25 161.3
R24 plus.n28 plus.n16 161.3
R25 plus.n31 plus.n30 161.3
R26 plus.n5 plus.n4 45.2793
R27 plus.n13 plus.n12 45.2793
R28 plus.n29 plus.n28 45.2793
R29 plus.n21 plus.n20 45.2793
R30 plus.n7 plus.n6 40.8975
R31 plus.n11 plus.n10 40.8975
R32 plus.n27 plus.n26 40.8975
R33 plus.n23 plus.n22 40.8975
R34 plus.n7 plus.n1 36.5157
R35 plus.n10 plus.n1 36.5157
R36 plus.n26 plus.n17 36.5157
R37 plus.n23 plus.n17 36.5157
R38 plus.n6 plus.n5 32.1338
R39 plus.n12 plus.n11 32.1338
R40 plus.n28 plus.n27 32.1338
R41 plus.n22 plus.n21 32.1338
R42 plus plus.n31 30.0236
R43 plus.n4 plus.n3 27.752
R44 plus.n14 plus.n13 27.752
R45 plus.n30 plus.n29 27.752
R46 plus.n20 plus.n19 27.752
R47 plus plus.n15 13.241
R48 plus.n8 plus.n2 0.189894
R49 plus.n9 plus.n8 0.189894
R50 plus.n9 plus.n0 0.189894
R51 plus.n15 plus.n0 0.189894
R52 plus.n31 plus.n16 0.189894
R53 plus.n25 plus.n16 0.189894
R54 plus.n25 plus.n24 0.189894
R55 plus.n24 plus.n18 0.189894
R56 source.n7 source.t3 45.521
R57 source.n27 source.t6 45.5208
R58 source.n20 source.t18 45.5208
R59 source.n0 source.t21 45.5208
R60 source.n2 source.n1 44.201
R61 source.n4 source.n3 44.201
R62 source.n6 source.n5 44.201
R63 source.n9 source.n8 44.201
R64 source.n11 source.n10 44.201
R65 source.n13 source.n12 44.201
R66 source.n26 source.n25 44.2008
R67 source.n24 source.n23 44.2008
R68 source.n22 source.n21 44.2008
R69 source.n19 source.n18 44.2008
R70 source.n17 source.n16 44.2008
R71 source.n15 source.n14 44.2008
R72 source.n15 source.n13 24.4742
R73 source.n28 source.n0 18.526
R74 source.n28 source.n27 5.49188
R75 source.n25 source.t12 1.3205
R76 source.n25 source.t1 1.3205
R77 source.n23 source.t5 1.3205
R78 source.n23 source.t2 1.3205
R79 source.n21 source.t9 1.3205
R80 source.n21 source.t0 1.3205
R81 source.n18 source.t14 1.3205
R82 source.n18 source.t17 1.3205
R83 source.n16 source.t25 1.3205
R84 source.n16 source.t27 1.3205
R85 source.n14 source.t19 1.3205
R86 source.n14 source.t15 1.3205
R87 source.n1 source.t16 1.3205
R88 source.n1 source.t20 1.3205
R89 source.n3 source.t22 1.3205
R90 source.n3 source.t23 1.3205
R91 source.n5 source.t26 1.3205
R92 source.n5 source.t24 1.3205
R93 source.n8 source.t8 1.3205
R94 source.n8 source.t7 1.3205
R95 source.n10 source.t10 1.3205
R96 source.n10 source.t13 1.3205
R97 source.n12 source.t4 1.3205
R98 source.n12 source.t11 1.3205
R99 source.n7 source.n6 0.698776
R100 source.n22 source.n20 0.698776
R101 source.n13 source.n11 0.457397
R102 source.n11 source.n9 0.457397
R103 source.n9 source.n7 0.457397
R104 source.n6 source.n4 0.457397
R105 source.n4 source.n2 0.457397
R106 source.n2 source.n0 0.457397
R107 source.n17 source.n15 0.457397
R108 source.n19 source.n17 0.457397
R109 source.n20 source.n19 0.457397
R110 source.n24 source.n22 0.457397
R111 source.n26 source.n24 0.457397
R112 source.n27 source.n26 0.457397
R113 source source.n28 0.188
R114 drain_left.n7 drain_left.t6 62.6567
R115 drain_left.n1 drain_left.t0 62.6565
R116 drain_left.n4 drain_left.n2 61.3365
R117 drain_left.n9 drain_left.n8 60.8798
R118 drain_left.n7 drain_left.n6 60.8798
R119 drain_left.n11 drain_left.n10 60.8796
R120 drain_left.n4 drain_left.n3 60.8796
R121 drain_left.n1 drain_left.n0 60.8796
R122 drain_left drain_left.n5 32.267
R123 drain_left drain_left.n11 6.11011
R124 drain_left.n2 drain_left.t10 1.3205
R125 drain_left.n2 drain_left.t11 1.3205
R126 drain_left.n3 drain_left.t3 1.3205
R127 drain_left.n3 drain_left.t12 1.3205
R128 drain_left.n0 drain_left.t2 1.3205
R129 drain_left.n0 drain_left.t13 1.3205
R130 drain_left.n10 drain_left.t7 1.3205
R131 drain_left.n10 drain_left.t9 1.3205
R132 drain_left.n8 drain_left.t4 1.3205
R133 drain_left.n8 drain_left.t5 1.3205
R134 drain_left.n6 drain_left.t8 1.3205
R135 drain_left.n6 drain_left.t1 1.3205
R136 drain_left.n9 drain_left.n7 0.457397
R137 drain_left.n11 drain_left.n9 0.457397
R138 drain_left.n5 drain_left.n1 0.287826
R139 drain_left.n5 drain_left.n4 0.0593781
R140 minus.n14 minus.t1 2013.81
R141 minus.n3 minus.t9 2013.81
R142 minus.n30 minus.t11 2013.81
R143 minus.n19 minus.t5 2013.81
R144 minus.n13 minus.t2 1964.15
R145 minus.n11 minus.t10 1964.15
R146 minus.n1 minus.t13 1964.15
R147 minus.n6 minus.t0 1964.15
R148 minus.n4 minus.t4 1964.15
R149 minus.n29 minus.t8 1964.15
R150 minus.n27 minus.t12 1964.15
R151 minus.n17 minus.t6 1964.15
R152 minus.n22 minus.t3 1964.15
R153 minus.n20 minus.t7 1964.15
R154 minus.n3 minus.n2 161.489
R155 minus.n19 minus.n18 161.489
R156 minus.n15 minus.n14 161.3
R157 minus.n12 minus.n0 161.3
R158 minus.n10 minus.n9 161.3
R159 minus.n8 minus.n7 161.3
R160 minus.n5 minus.n2 161.3
R161 minus.n31 minus.n30 161.3
R162 minus.n28 minus.n16 161.3
R163 minus.n26 minus.n25 161.3
R164 minus.n24 minus.n23 161.3
R165 minus.n21 minus.n18 161.3
R166 minus.n13 minus.n12 45.2793
R167 minus.n5 minus.n4 45.2793
R168 minus.n21 minus.n20 45.2793
R169 minus.n29 minus.n28 45.2793
R170 minus.n11 minus.n10 40.8975
R171 minus.n7 minus.n6 40.8975
R172 minus.n23 minus.n22 40.8975
R173 minus.n27 minus.n26 40.8975
R174 minus.n32 minus.n15 37.2789
R175 minus.n10 minus.n1 36.5157
R176 minus.n7 minus.n1 36.5157
R177 minus.n23 minus.n17 36.5157
R178 minus.n26 minus.n17 36.5157
R179 minus.n12 minus.n11 32.1338
R180 minus.n6 minus.n5 32.1338
R181 minus.n22 minus.n21 32.1338
R182 minus.n28 minus.n27 32.1338
R183 minus.n14 minus.n13 27.752
R184 minus.n4 minus.n3 27.752
R185 minus.n20 minus.n19 27.752
R186 minus.n30 minus.n29 27.752
R187 minus.n32 minus.n31 6.46073
R188 minus.n15 minus.n0 0.189894
R189 minus.n9 minus.n0 0.189894
R190 minus.n9 minus.n8 0.189894
R191 minus.n8 minus.n2 0.189894
R192 minus.n24 minus.n18 0.189894
R193 minus.n25 minus.n24 0.189894
R194 minus.n25 minus.n16 0.189894
R195 minus.n31 minus.n16 0.189894
R196 minus minus.n32 0.188
R197 drain_right.n1 drain_right.t8 62.6565
R198 drain_right.n11 drain_right.t12 62.1998
R199 drain_right.n8 drain_right.n6 61.3365
R200 drain_right.n4 drain_right.n2 61.3365
R201 drain_right.n8 drain_right.n7 60.8798
R202 drain_right.n10 drain_right.n9 60.8798
R203 drain_right.n4 drain_right.n3 60.8796
R204 drain_right.n1 drain_right.n0 60.8796
R205 drain_right drain_right.n5 31.7137
R206 drain_right drain_right.n11 5.88166
R207 drain_right.n2 drain_right.t5 1.3205
R208 drain_right.n2 drain_right.t2 1.3205
R209 drain_right.n3 drain_right.t7 1.3205
R210 drain_right.n3 drain_right.t1 1.3205
R211 drain_right.n0 drain_right.t6 1.3205
R212 drain_right.n0 drain_right.t10 1.3205
R213 drain_right.n6 drain_right.t9 1.3205
R214 drain_right.n6 drain_right.t4 1.3205
R215 drain_right.n7 drain_right.t0 1.3205
R216 drain_right.n7 drain_right.t13 1.3205
R217 drain_right.n9 drain_right.t11 1.3205
R218 drain_right.n9 drain_right.t3 1.3205
R219 drain_right.n11 drain_right.n10 0.457397
R220 drain_right.n10 drain_right.n8 0.457397
R221 drain_right.n5 drain_right.n1 0.287826
R222 drain_right.n5 drain_right.n4 0.0593781
C0 drain_right drain_left 0.796704f
C1 drain_right minus 4.85576f
C2 drain_left minus 0.171065f
C3 drain_right source 41.1429f
C4 drain_left source 41.1573f
C5 source minus 4.29847f
C6 drain_right plus 0.306693f
C7 drain_left plus 5.002069f
C8 plus minus 5.66056f
C9 plus source 4.31338f
C10 drain_right a_n1564_n3888# 8.49991f
C11 drain_left a_n1564_n3888# 8.76831f
C12 source a_n1564_n3888# 7.048458f
C13 minus a_n1564_n3888# 6.255233f
C14 plus a_n1564_n3888# 8.54813f
C15 drain_right.t8 a_n1564_n3888# 4.78947f
C16 drain_right.t6 a_n1564_n3888# 0.414835f
C17 drain_right.t10 a_n1564_n3888# 0.414835f
C18 drain_right.n0 a_n1564_n3888# 3.74962f
C19 drain_right.n1 a_n1564_n3888# 0.817182f
C20 drain_right.t5 a_n1564_n3888# 0.414835f
C21 drain_right.t2 a_n1564_n3888# 0.414835f
C22 drain_right.n2 a_n1564_n3888# 3.75263f
C23 drain_right.t7 a_n1564_n3888# 0.414835f
C24 drain_right.t1 a_n1564_n3888# 0.414835f
C25 drain_right.n3 a_n1564_n3888# 3.74962f
C26 drain_right.n4 a_n1564_n3888# 0.759371f
C27 drain_right.n5 a_n1564_n3888# 1.77109f
C28 drain_right.t9 a_n1564_n3888# 0.414835f
C29 drain_right.t4 a_n1564_n3888# 0.414835f
C30 drain_right.n6 a_n1564_n3888# 3.75262f
C31 drain_right.t0 a_n1564_n3888# 0.414835f
C32 drain_right.t13 a_n1564_n3888# 0.414835f
C33 drain_right.n7 a_n1564_n3888# 3.74963f
C34 drain_right.n8 a_n1564_n3888# 0.790481f
C35 drain_right.t11 a_n1564_n3888# 0.414835f
C36 drain_right.t3 a_n1564_n3888# 0.414835f
C37 drain_right.n9 a_n1564_n3888# 3.74963f
C38 drain_right.n10 a_n1564_n3888# 0.38969f
C39 drain_right.t12 a_n1564_n3888# 4.78621f
C40 drain_right.n11 a_n1564_n3888# 0.731491f
C41 minus.n0 a_n1564_n3888# 0.055374f
C42 minus.t1 a_n1564_n3888# 0.47327f
C43 minus.t2 a_n1564_n3888# 0.468657f
C44 minus.t10 a_n1564_n3888# 0.468657f
C45 minus.t13 a_n1564_n3888# 0.468657f
C46 minus.n1 a_n1564_n3888# 0.185704f
C47 minus.n2 a_n1564_n3888# 0.123642f
C48 minus.t0 a_n1564_n3888# 0.468657f
C49 minus.t4 a_n1564_n3888# 0.468657f
C50 minus.t9 a_n1564_n3888# 0.47327f
C51 minus.n3 a_n1564_n3888# 0.20193f
C52 minus.n4 a_n1564_n3888# 0.185704f
C53 minus.n5 a_n1564_n3888# 0.019394f
C54 minus.n6 a_n1564_n3888# 0.185704f
C55 minus.n7 a_n1564_n3888# 0.019394f
C56 minus.n8 a_n1564_n3888# 0.055374f
C57 minus.n9 a_n1564_n3888# 0.055374f
C58 minus.n10 a_n1564_n3888# 0.019394f
C59 minus.n11 a_n1564_n3888# 0.185704f
C60 minus.n12 a_n1564_n3888# 0.019394f
C61 minus.n13 a_n1564_n3888# 0.185704f
C62 minus.n14 a_n1564_n3888# 0.20185f
C63 minus.n15 a_n1564_n3888# 2.04727f
C64 minus.n16 a_n1564_n3888# 0.055374f
C65 minus.t8 a_n1564_n3888# 0.468657f
C66 minus.t12 a_n1564_n3888# 0.468657f
C67 minus.t6 a_n1564_n3888# 0.468657f
C68 minus.n17 a_n1564_n3888# 0.185704f
C69 minus.n18 a_n1564_n3888# 0.123642f
C70 minus.t3 a_n1564_n3888# 0.468657f
C71 minus.t7 a_n1564_n3888# 0.468657f
C72 minus.t5 a_n1564_n3888# 0.47327f
C73 minus.n19 a_n1564_n3888# 0.20193f
C74 minus.n20 a_n1564_n3888# 0.185704f
C75 minus.n21 a_n1564_n3888# 0.019394f
C76 minus.n22 a_n1564_n3888# 0.185704f
C77 minus.n23 a_n1564_n3888# 0.019394f
C78 minus.n24 a_n1564_n3888# 0.055374f
C79 minus.n25 a_n1564_n3888# 0.055374f
C80 minus.n26 a_n1564_n3888# 0.019394f
C81 minus.n27 a_n1564_n3888# 0.185704f
C82 minus.n28 a_n1564_n3888# 0.019394f
C83 minus.n29 a_n1564_n3888# 0.185704f
C84 minus.t11 a_n1564_n3888# 0.47327f
C85 minus.n30 a_n1564_n3888# 0.20185f
C86 minus.n31 a_n1564_n3888# 0.356889f
C87 minus.n32 a_n1564_n3888# 2.48055f
C88 drain_left.t0 a_n1564_n3888# 4.79602f
C89 drain_left.t2 a_n1564_n3888# 0.415402f
C90 drain_left.t13 a_n1564_n3888# 0.415402f
C91 drain_left.n0 a_n1564_n3888# 3.75475f
C92 drain_left.n1 a_n1564_n3888# 0.8183f
C93 drain_left.t10 a_n1564_n3888# 0.415402f
C94 drain_left.t11 a_n1564_n3888# 0.415402f
C95 drain_left.n2 a_n1564_n3888# 3.75776f
C96 drain_left.t3 a_n1564_n3888# 0.415402f
C97 drain_left.t12 a_n1564_n3888# 0.415402f
C98 drain_left.n3 a_n1564_n3888# 3.75475f
C99 drain_left.n4 a_n1564_n3888# 0.760409f
C100 drain_left.n5 a_n1564_n3888# 1.8468f
C101 drain_left.t6 a_n1564_n3888# 4.79602f
C102 drain_left.t8 a_n1564_n3888# 0.415402f
C103 drain_left.t1 a_n1564_n3888# 0.415402f
C104 drain_left.n6 a_n1564_n3888# 3.75475f
C105 drain_left.n7 a_n1564_n3888# 0.834614f
C106 drain_left.t4 a_n1564_n3888# 0.415402f
C107 drain_left.t5 a_n1564_n3888# 0.415402f
C108 drain_left.n8 a_n1564_n3888# 3.75475f
C109 drain_left.n9 a_n1564_n3888# 0.390223f
C110 drain_left.t7 a_n1564_n3888# 0.415402f
C111 drain_left.t9 a_n1564_n3888# 0.415402f
C112 drain_left.n10 a_n1564_n3888# 3.75474f
C113 drain_left.n11 a_n1564_n3888# 0.677045f
C114 source.t21 a_n1564_n3888# 4.75824f
C115 source.n0 a_n1564_n3888# 2.18787f
C116 source.t16 a_n1564_n3888# 0.424592f
C117 source.t20 a_n1564_n3888# 0.424592f
C118 source.n1 a_n1564_n3888# 3.72969f
C119 source.n2 a_n1564_n3888# 0.458303f
C120 source.t22 a_n1564_n3888# 0.424592f
C121 source.t23 a_n1564_n3888# 0.424592f
C122 source.n3 a_n1564_n3888# 3.72969f
C123 source.n4 a_n1564_n3888# 0.458303f
C124 source.t26 a_n1564_n3888# 0.424592f
C125 source.t24 a_n1564_n3888# 0.424592f
C126 source.n5 a_n1564_n3888# 3.72969f
C127 source.n6 a_n1564_n3888# 0.486163f
C128 source.t3 a_n1564_n3888# 4.75824f
C129 source.n7 a_n1564_n3888# 0.615583f
C130 source.t8 a_n1564_n3888# 0.424592f
C131 source.t7 a_n1564_n3888# 0.424592f
C132 source.n8 a_n1564_n3888# 3.72969f
C133 source.n9 a_n1564_n3888# 0.458303f
C134 source.t10 a_n1564_n3888# 0.424592f
C135 source.t13 a_n1564_n3888# 0.424592f
C136 source.n10 a_n1564_n3888# 3.72969f
C137 source.n11 a_n1564_n3888# 0.458303f
C138 source.t4 a_n1564_n3888# 0.424592f
C139 source.t11 a_n1564_n3888# 0.424592f
C140 source.n12 a_n1564_n3888# 3.72969f
C141 source.n13 a_n1564_n3888# 2.70288f
C142 source.t19 a_n1564_n3888# 0.424592f
C143 source.t15 a_n1564_n3888# 0.424592f
C144 source.n14 a_n1564_n3888# 3.72968f
C145 source.n15 a_n1564_n3888# 2.70288f
C146 source.t25 a_n1564_n3888# 0.424592f
C147 source.t27 a_n1564_n3888# 0.424592f
C148 source.n16 a_n1564_n3888# 3.72968f
C149 source.n17 a_n1564_n3888# 0.458308f
C150 source.t14 a_n1564_n3888# 0.424592f
C151 source.t17 a_n1564_n3888# 0.424592f
C152 source.n18 a_n1564_n3888# 3.72968f
C153 source.n19 a_n1564_n3888# 0.458308f
C154 source.t18 a_n1564_n3888# 4.75824f
C155 source.n20 a_n1564_n3888# 0.615588f
C156 source.t9 a_n1564_n3888# 0.424592f
C157 source.t0 a_n1564_n3888# 0.424592f
C158 source.n21 a_n1564_n3888# 3.72968f
C159 source.n22 a_n1564_n3888# 0.486168f
C160 source.t5 a_n1564_n3888# 0.424592f
C161 source.t2 a_n1564_n3888# 0.424592f
C162 source.n23 a_n1564_n3888# 3.72968f
C163 source.n24 a_n1564_n3888# 0.458308f
C164 source.t12 a_n1564_n3888# 0.424592f
C165 source.t1 a_n1564_n3888# 0.424592f
C166 source.n25 a_n1564_n3888# 3.72968f
C167 source.n26 a_n1564_n3888# 0.458308f
C168 source.t6 a_n1564_n3888# 4.75824f
C169 source.n27 a_n1564_n3888# 0.783449f
C170 source.n28 a_n1564_n3888# 2.61329f
C171 plus.n0 a_n1564_n3888# 0.056168f
C172 plus.t6 a_n1564_n3888# 0.475375f
C173 plus.t8 a_n1564_n3888# 0.475375f
C174 plus.t9 a_n1564_n3888# 0.475375f
C175 plus.n1 a_n1564_n3888# 0.188366f
C176 plus.n2 a_n1564_n3888# 0.125414f
C177 plus.t12 a_n1564_n3888# 0.475375f
C178 plus.t5 a_n1564_n3888# 0.475375f
C179 plus.t7 a_n1564_n3888# 0.480054f
C180 plus.n3 a_n1564_n3888# 0.204825f
C181 plus.n4 a_n1564_n3888# 0.188366f
C182 plus.n5 a_n1564_n3888# 0.019672f
C183 plus.n6 a_n1564_n3888# 0.188366f
C184 plus.n7 a_n1564_n3888# 0.019672f
C185 plus.n8 a_n1564_n3888# 0.056168f
C186 plus.n9 a_n1564_n3888# 0.056168f
C187 plus.n10 a_n1564_n3888# 0.019672f
C188 plus.n11 a_n1564_n3888# 0.188366f
C189 plus.n12 a_n1564_n3888# 0.019672f
C190 plus.n13 a_n1564_n3888# 0.188366f
C191 plus.t4 a_n1564_n3888# 0.480054f
C192 plus.n14 a_n1564_n3888# 0.204744f
C193 plus.n15 a_n1564_n3888# 0.704584f
C194 plus.n16 a_n1564_n3888# 0.056168f
C195 plus.t13 a_n1564_n3888# 0.480054f
C196 plus.t11 a_n1564_n3888# 0.475375f
C197 plus.t0 a_n1564_n3888# 0.475375f
C198 plus.t10 a_n1564_n3888# 0.475375f
C199 plus.n17 a_n1564_n3888# 0.188366f
C200 plus.n18 a_n1564_n3888# 0.125414f
C201 plus.t1 a_n1564_n3888# 0.475375f
C202 plus.t3 a_n1564_n3888# 0.475375f
C203 plus.t2 a_n1564_n3888# 0.480054f
C204 plus.n19 a_n1564_n3888# 0.204825f
C205 plus.n20 a_n1564_n3888# 0.188366f
C206 plus.n21 a_n1564_n3888# 0.019672f
C207 plus.n22 a_n1564_n3888# 0.188366f
C208 plus.n23 a_n1564_n3888# 0.019672f
C209 plus.n24 a_n1564_n3888# 0.056168f
C210 plus.n25 a_n1564_n3888# 0.056168f
C211 plus.n26 a_n1564_n3888# 0.019672f
C212 plus.n27 a_n1564_n3888# 0.188366f
C213 plus.n28 a_n1564_n3888# 0.019672f
C214 plus.n29 a_n1564_n3888# 0.188366f
C215 plus.n30 a_n1564_n3888# 0.204744f
C216 plus.n31 a_n1564_n3888# 1.70251f
.ends

