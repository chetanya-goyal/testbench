* NGSPICE file created from diffpair347.ext - technology: sky130A

.subckt diffpair347 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t17 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 drain_left.t14 plus.t1 source.t31 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 drain_right.t15 minus.t0 source.t3 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_left.t13 plus.t2 source.t26 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 source.t8 minus.t1 drain_right.t14 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 source.t1 minus.t2 drain_right.t13 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X6 drain_left.t12 plus.t3 source.t27 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X7 source.t10 minus.t3 drain_right.t12 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 source.t18 plus.t4 drain_left.t11 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X9 a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X10 drain_left.t10 plus.t5 source.t20 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X11 source.t24 plus.t6 drain_left.t9 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X12 source.t13 minus.t4 drain_right.t11 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X13 a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X14 source.t7 minus.t5 drain_right.t10 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X15 source.t22 plus.t7 drain_left.t8 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X16 source.t21 plus.t8 drain_left.t7 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 source.t16 plus.t9 drain_left.t6 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X18 a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X19 drain_right.t9 minus.t6 source.t9 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X20 drain_left.t5 plus.t10 source.t30 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X21 drain_right.t8 minus.t7 source.t12 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X22 source.t25 plus.t11 drain_left.t4 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X23 drain_right.t7 minus.t8 source.t6 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X24 source.t15 minus.t9 drain_right.t6 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X25 source.t4 minus.t10 drain_right.t5 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X26 drain_right.t4 minus.t11 source.t0 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X27 source.t23 plus.t12 drain_left.t3 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X28 drain_left.t2 plus.t13 source.t29 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X29 drain_right.t3 minus.t12 source.t2 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X30 a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X31 source.t5 minus.t13 drain_right.t2 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X32 source.t28 plus.t14 drain_left.t1 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X33 drain_right.t1 minus.t14 source.t11 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X34 drain_right.t0 minus.t15 source.t14 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X35 drain_left.t0 plus.t15 source.t19 a_n1760_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
R0 plus.n4 plus.t6 1033.82
R1 plus.n19 plus.t3 1033.82
R2 plus.n25 plus.t13 1033.82
R3 plus.n40 plus.t4 1033.82
R4 plus.n5 plus.t1 992.92
R5 plus.n3 plus.t9 992.92
R6 plus.n10 plus.t0 992.92
R7 plus.n1 plus.t8 992.92
R8 plus.n16 plus.t15 992.92
R9 plus.n18 plus.t7 992.92
R10 plus.n26 plus.t11 992.92
R11 plus.n24 plus.t5 992.92
R12 plus.n31 plus.t14 992.92
R13 plus.n22 plus.t2 992.92
R14 plus.n37 plus.t12 992.92
R15 plus.n39 plus.t10 992.92
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus.n6 plus.n5 29.2126
R47 plus.n18 plus.n17 29.2126
R48 plus.n39 plus.n38 29.2126
R49 plus.n27 plus.n26 29.2126
R50 plus plus.n41 28.499
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 10.974
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n7 source.t24 51.0588
R73 source.n8 source.t0 51.0588
R74 source.n15 source.t13 51.0588
R75 source.n31 source.t12 51.0586
R76 source.n24 source.t5 51.0586
R77 source.n23 source.t29 51.0586
R78 source.n16 source.t18 51.0586
R79 source.n0 source.t27 51.0586
R80 source.n2 source.n1 48.8588
R81 source.n4 source.n3 48.8588
R82 source.n6 source.n5 48.8588
R83 source.n10 source.n9 48.8588
R84 source.n12 source.n11 48.8588
R85 source.n14 source.n13 48.8588
R86 source.n30 source.n29 48.8586
R87 source.n28 source.n27 48.8586
R88 source.n26 source.n25 48.8586
R89 source.n22 source.n21 48.8586
R90 source.n20 source.n19 48.8586
R91 source.n18 source.n17 48.8586
R92 source.n16 source.n15 19.515
R93 source.n32 source.n0 14.0021
R94 source.n32 source.n31 5.51343
R95 source.n29 source.t2 2.2005
R96 source.n29 source.t15 2.2005
R97 source.n27 source.t9 2.2005
R98 source.n27 source.t1 2.2005
R99 source.n25 source.t3 2.2005
R100 source.n25 source.t4 2.2005
R101 source.n21 source.t20 2.2005
R102 source.n21 source.t25 2.2005
R103 source.n19 source.t26 2.2005
R104 source.n19 source.t28 2.2005
R105 source.n17 source.t30 2.2005
R106 source.n17 source.t23 2.2005
R107 source.n1 source.t19 2.2005
R108 source.n1 source.t22 2.2005
R109 source.n3 source.t17 2.2005
R110 source.n3 source.t21 2.2005
R111 source.n5 source.t31 2.2005
R112 source.n5 source.t16 2.2005
R113 source.n9 source.t6 2.2005
R114 source.n9 source.t10 2.2005
R115 source.n11 source.t11 2.2005
R116 source.n11 source.t8 2.2005
R117 source.n13 source.t14 2.2005
R118 source.n13 source.t7 2.2005
R119 source.n15 source.n14 0.5005
R120 source.n14 source.n12 0.5005
R121 source.n12 source.n10 0.5005
R122 source.n10 source.n8 0.5005
R123 source.n7 source.n6 0.5005
R124 source.n6 source.n4 0.5005
R125 source.n4 source.n2 0.5005
R126 source.n2 source.n0 0.5005
R127 source.n18 source.n16 0.5005
R128 source.n20 source.n18 0.5005
R129 source.n22 source.n20 0.5005
R130 source.n23 source.n22 0.5005
R131 source.n26 source.n24 0.5005
R132 source.n28 source.n26 0.5005
R133 source.n30 source.n28 0.5005
R134 source.n31 source.n30 0.5005
R135 source.n8 source.n7 0.470328
R136 source.n24 source.n23 0.470328
R137 source source.n32 0.188
R138 drain_left.n9 drain_left.n7 66.0376
R139 drain_left.n5 drain_left.n3 66.0373
R140 drain_left.n2 drain_left.n0 66.0373
R141 drain_left.n11 drain_left.n10 65.5376
R142 drain_left.n9 drain_left.n8 65.5376
R143 drain_left.n13 drain_left.n12 65.5374
R144 drain_left.n5 drain_left.n4 65.5373
R145 drain_left.n2 drain_left.n1 65.5373
R146 drain_left drain_left.n6 28.3443
R147 drain_left drain_left.n13 6.15322
R148 drain_left.n3 drain_left.t4 2.2005
R149 drain_left.n3 drain_left.t2 2.2005
R150 drain_left.n4 drain_left.t1 2.2005
R151 drain_left.n4 drain_left.t10 2.2005
R152 drain_left.n1 drain_left.t3 2.2005
R153 drain_left.n1 drain_left.t13 2.2005
R154 drain_left.n0 drain_left.t11 2.2005
R155 drain_left.n0 drain_left.t5 2.2005
R156 drain_left.n12 drain_left.t8 2.2005
R157 drain_left.n12 drain_left.t12 2.2005
R158 drain_left.n10 drain_left.t7 2.2005
R159 drain_left.n10 drain_left.t0 2.2005
R160 drain_left.n8 drain_left.t6 2.2005
R161 drain_left.n8 drain_left.t15 2.2005
R162 drain_left.n7 drain_left.t9 2.2005
R163 drain_left.n7 drain_left.t14 2.2005
R164 drain_left.n11 drain_left.n9 0.5005
R165 drain_left.n13 drain_left.n11 0.5005
R166 drain_left.n6 drain_left.n5 0.195154
R167 drain_left.n6 drain_left.n2 0.195154
R168 minus.n19 minus.t4 1033.82
R169 minus.n4 minus.t11 1033.82
R170 minus.n40 minus.t7 1033.82
R171 minus.n25 minus.t13 1033.82
R172 minus.n18 minus.t15 992.92
R173 minus.n16 minus.t5 992.92
R174 minus.n1 minus.t14 992.92
R175 minus.n10 minus.t1 992.92
R176 minus.n3 minus.t8 992.92
R177 minus.n5 minus.t3 992.92
R178 minus.n39 minus.t9 992.92
R179 minus.n37 minus.t12 992.92
R180 minus.n22 minus.t2 992.92
R181 minus.n31 minus.t6 992.92
R182 minus.n24 minus.t10 992.92
R183 minus.n26 minus.t0 992.92
R184 minus.n7 minus.n4 161.489
R185 minus.n28 minus.n25 161.489
R186 minus.n20 minus.n19 161.3
R187 minus.n17 minus.n0 161.3
R188 minus.n15 minus.n14 161.3
R189 minus.n13 minus.n12 161.3
R190 minus.n11 minus.n2 161.3
R191 minus.n9 minus.n8 161.3
R192 minus.n7 minus.n6 161.3
R193 minus.n41 minus.n40 161.3
R194 minus.n38 minus.n21 161.3
R195 minus.n36 minus.n35 161.3
R196 minus.n34 minus.n33 161.3
R197 minus.n32 minus.n23 161.3
R198 minus.n30 minus.n29 161.3
R199 minus.n28 minus.n27 161.3
R200 minus.n12 minus.n11 73.0308
R201 minus.n33 minus.n32 73.0308
R202 minus.n15 minus.n1 67.1884
R203 minus.n10 minus.n9 67.1884
R204 minus.n31 minus.n30 67.1884
R205 minus.n36 minus.n22 67.1884
R206 minus.n17 minus.n16 55.5035
R207 minus.n6 minus.n3 55.5035
R208 minus.n27 minus.n24 55.5035
R209 minus.n38 minus.n37 55.5035
R210 minus.n19 minus.n18 43.8187
R211 minus.n5 minus.n4 43.8187
R212 minus.n26 minus.n25 43.8187
R213 minus.n40 minus.n39 43.8187
R214 minus.n42 minus.n20 33.4816
R215 minus.n18 minus.n17 29.2126
R216 minus.n6 minus.n5 29.2126
R217 minus.n27 minus.n26 29.2126
R218 minus.n39 minus.n38 29.2126
R219 minus.n16 minus.n15 17.5278
R220 minus.n9 minus.n3 17.5278
R221 minus.n30 minus.n24 17.5278
R222 minus.n37 minus.n36 17.5278
R223 minus.n42 minus.n41 6.46641
R224 minus.n12 minus.n1 5.84292
R225 minus.n11 minus.n10 5.84292
R226 minus.n32 minus.n31 5.84292
R227 minus.n33 minus.n22 5.84292
R228 minus.n20 minus.n0 0.189894
R229 minus.n14 minus.n0 0.189894
R230 minus.n14 minus.n13 0.189894
R231 minus.n13 minus.n2 0.189894
R232 minus.n8 minus.n2 0.189894
R233 minus.n8 minus.n7 0.189894
R234 minus.n29 minus.n28 0.189894
R235 minus.n29 minus.n23 0.189894
R236 minus.n34 minus.n23 0.189894
R237 minus.n35 minus.n34 0.189894
R238 minus.n35 minus.n21 0.189894
R239 minus.n41 minus.n21 0.189894
R240 minus minus.n42 0.188
R241 drain_right.n9 drain_right.n7 66.0374
R242 drain_right.n5 drain_right.n3 66.0373
R243 drain_right.n2 drain_right.n0 66.0373
R244 drain_right.n9 drain_right.n8 65.5376
R245 drain_right.n11 drain_right.n10 65.5376
R246 drain_right.n13 drain_right.n12 65.5376
R247 drain_right.n5 drain_right.n4 65.5373
R248 drain_right.n2 drain_right.n1 65.5373
R249 drain_right drain_right.n6 27.7911
R250 drain_right drain_right.n13 6.15322
R251 drain_right.n3 drain_right.t6 2.2005
R252 drain_right.n3 drain_right.t8 2.2005
R253 drain_right.n4 drain_right.t13 2.2005
R254 drain_right.n4 drain_right.t3 2.2005
R255 drain_right.n1 drain_right.t5 2.2005
R256 drain_right.n1 drain_right.t9 2.2005
R257 drain_right.n0 drain_right.t2 2.2005
R258 drain_right.n0 drain_right.t15 2.2005
R259 drain_right.n7 drain_right.t12 2.2005
R260 drain_right.n7 drain_right.t4 2.2005
R261 drain_right.n8 drain_right.t14 2.2005
R262 drain_right.n8 drain_right.t7 2.2005
R263 drain_right.n10 drain_right.t10 2.2005
R264 drain_right.n10 drain_right.t1 2.2005
R265 drain_right.n12 drain_right.t11 2.2005
R266 drain_right.n12 drain_right.t0 2.2005
R267 drain_right.n13 drain_right.n11 0.5005
R268 drain_right.n11 drain_right.n9 0.5005
R269 drain_right.n6 drain_right.n5 0.195154
R270 drain_right.n6 drain_right.n2 0.195154
C0 source drain_left 25.6219f
C1 drain_right minus 4.01194f
C2 source plus 3.79189f
C3 drain_right drain_left 0.897273f
C4 drain_left minus 0.171252f
C5 drain_right plus 0.324551f
C6 minus plus 4.79461f
C7 drain_left plus 4.18228f
C8 drain_right source 25.6219f
C9 source minus 3.77786f
C10 drain_right a_n1760_n2688# 5.95423f
C11 drain_left a_n1760_n2688# 6.23622f
C12 source a_n1760_n2688# 7.031454f
C13 minus a_n1760_n2688# 6.648073f
C14 plus a_n1760_n2688# 8.466929f
C15 drain_right.t2 a_n1760_n2688# 0.253097f
C16 drain_right.t15 a_n1760_n2688# 0.253097f
C17 drain_right.n0 a_n1760_n2688# 2.21689f
C18 drain_right.t5 a_n1760_n2688# 0.253097f
C19 drain_right.t9 a_n1760_n2688# 0.253097f
C20 drain_right.n1 a_n1760_n2688# 2.21376f
C21 drain_right.n2 a_n1760_n2688# 0.779873f
C22 drain_right.t6 a_n1760_n2688# 0.253097f
C23 drain_right.t8 a_n1760_n2688# 0.253097f
C24 drain_right.n3 a_n1760_n2688# 2.21689f
C25 drain_right.t13 a_n1760_n2688# 0.253097f
C26 drain_right.t3 a_n1760_n2688# 0.253097f
C27 drain_right.n4 a_n1760_n2688# 2.21376f
C28 drain_right.n5 a_n1760_n2688# 0.779873f
C29 drain_right.n6 a_n1760_n2688# 1.393f
C30 drain_right.t12 a_n1760_n2688# 0.253097f
C31 drain_right.t4 a_n1760_n2688# 0.253097f
C32 drain_right.n7 a_n1760_n2688# 2.21689f
C33 drain_right.t14 a_n1760_n2688# 0.253097f
C34 drain_right.t7 a_n1760_n2688# 0.253097f
C35 drain_right.n8 a_n1760_n2688# 2.21376f
C36 drain_right.n9 a_n1760_n2688# 0.810649f
C37 drain_right.t10 a_n1760_n2688# 0.253097f
C38 drain_right.t1 a_n1760_n2688# 0.253097f
C39 drain_right.n10 a_n1760_n2688# 2.21376f
C40 drain_right.n11 a_n1760_n2688# 0.399721f
C41 drain_right.t11 a_n1760_n2688# 0.253097f
C42 drain_right.t0 a_n1760_n2688# 0.253097f
C43 drain_right.n12 a_n1760_n2688# 2.21376f
C44 drain_right.n13 a_n1760_n2688# 0.693467f
C45 minus.n0 a_n1760_n2688# 0.051978f
C46 minus.t4 a_n1760_n2688# 0.33701f
C47 minus.t15 a_n1760_n2688# 0.331392f
C48 minus.t5 a_n1760_n2688# 0.331392f
C49 minus.t14 a_n1760_n2688# 0.331392f
C50 minus.n1 a_n1760_n2688# 0.141054f
C51 minus.n2 a_n1760_n2688# 0.051978f
C52 minus.t1 a_n1760_n2688# 0.331392f
C53 minus.t8 a_n1760_n2688# 0.331392f
C54 minus.n3 a_n1760_n2688# 0.141054f
C55 minus.t11 a_n1760_n2688# 0.33701f
C56 minus.n4 a_n1760_n2688# 0.156277f
C57 minus.t3 a_n1760_n2688# 0.331392f
C58 minus.n5 a_n1760_n2688# 0.141054f
C59 minus.n6 a_n1760_n2688# 0.019807f
C60 minus.n7 a_n1760_n2688# 0.113818f
C61 minus.n8 a_n1760_n2688# 0.051978f
C62 minus.n9 a_n1760_n2688# 0.019807f
C63 minus.n10 a_n1760_n2688# 0.141054f
C64 minus.n11 a_n1760_n2688# 0.018525f
C65 minus.n12 a_n1760_n2688# 0.018525f
C66 minus.n13 a_n1760_n2688# 0.051978f
C67 minus.n14 a_n1760_n2688# 0.051978f
C68 minus.n15 a_n1760_n2688# 0.019807f
C69 minus.n16 a_n1760_n2688# 0.141054f
C70 minus.n17 a_n1760_n2688# 0.019807f
C71 minus.n18 a_n1760_n2688# 0.141054f
C72 minus.n19 a_n1760_n2688# 0.156204f
C73 minus.n20 a_n1760_n2688# 1.62143f
C74 minus.n21 a_n1760_n2688# 0.051978f
C75 minus.t9 a_n1760_n2688# 0.331392f
C76 minus.t12 a_n1760_n2688# 0.331392f
C77 minus.t2 a_n1760_n2688# 0.331392f
C78 minus.n22 a_n1760_n2688# 0.141054f
C79 minus.n23 a_n1760_n2688# 0.051978f
C80 minus.t6 a_n1760_n2688# 0.331392f
C81 minus.t10 a_n1760_n2688# 0.331392f
C82 minus.n24 a_n1760_n2688# 0.141054f
C83 minus.t13 a_n1760_n2688# 0.33701f
C84 minus.n25 a_n1760_n2688# 0.156277f
C85 minus.t0 a_n1760_n2688# 0.331392f
C86 minus.n26 a_n1760_n2688# 0.141054f
C87 minus.n27 a_n1760_n2688# 0.019807f
C88 minus.n28 a_n1760_n2688# 0.113818f
C89 minus.n29 a_n1760_n2688# 0.051978f
C90 minus.n30 a_n1760_n2688# 0.019807f
C91 minus.n31 a_n1760_n2688# 0.141054f
C92 minus.n32 a_n1760_n2688# 0.018525f
C93 minus.n33 a_n1760_n2688# 0.018525f
C94 minus.n34 a_n1760_n2688# 0.051978f
C95 minus.n35 a_n1760_n2688# 0.051978f
C96 minus.n36 a_n1760_n2688# 0.019807f
C97 minus.n37 a_n1760_n2688# 0.141054f
C98 minus.n38 a_n1760_n2688# 0.019807f
C99 minus.n39 a_n1760_n2688# 0.141054f
C100 minus.t7 a_n1760_n2688# 0.33701f
C101 minus.n40 a_n1760_n2688# 0.156204f
C102 minus.n41 a_n1760_n2688# 0.335699f
C103 minus.n42 a_n1760_n2688# 1.98642f
C104 drain_left.t11 a_n1760_n2688# 0.253615f
C105 drain_left.t5 a_n1760_n2688# 0.253615f
C106 drain_left.n0 a_n1760_n2688# 2.22142f
C107 drain_left.t3 a_n1760_n2688# 0.253615f
C108 drain_left.t13 a_n1760_n2688# 0.253615f
C109 drain_left.n1 a_n1760_n2688# 2.21828f
C110 drain_left.n2 a_n1760_n2688# 0.781467f
C111 drain_left.t4 a_n1760_n2688# 0.253615f
C112 drain_left.t2 a_n1760_n2688# 0.253615f
C113 drain_left.n3 a_n1760_n2688# 2.22142f
C114 drain_left.t1 a_n1760_n2688# 0.253615f
C115 drain_left.t10 a_n1760_n2688# 0.253615f
C116 drain_left.n4 a_n1760_n2688# 2.21828f
C117 drain_left.n5 a_n1760_n2688# 0.781467f
C118 drain_left.n6 a_n1760_n2688# 1.46935f
C119 drain_left.t9 a_n1760_n2688# 0.253615f
C120 drain_left.t14 a_n1760_n2688# 0.253615f
C121 drain_left.n7 a_n1760_n2688# 2.22143f
C122 drain_left.t6 a_n1760_n2688# 0.253615f
C123 drain_left.t15 a_n1760_n2688# 0.253615f
C124 drain_left.n8 a_n1760_n2688# 2.21828f
C125 drain_left.n9 a_n1760_n2688# 0.812297f
C126 drain_left.t7 a_n1760_n2688# 0.253615f
C127 drain_left.t0 a_n1760_n2688# 0.253615f
C128 drain_left.n10 a_n1760_n2688# 2.21828f
C129 drain_left.n11 a_n1760_n2688# 0.400538f
C130 drain_left.t8 a_n1760_n2688# 0.253615f
C131 drain_left.t12 a_n1760_n2688# 0.253615f
C132 drain_left.n12 a_n1760_n2688# 2.21828f
C133 drain_left.n13 a_n1760_n2688# 0.694894f
C134 source.t27 a_n1760_n2688# 2.30057f
C135 source.n0 a_n1760_n2688# 1.31584f
C136 source.t19 a_n1760_n2688# 0.215743f
C137 source.t22 a_n1760_n2688# 0.215743f
C138 source.n1 a_n1760_n2688# 1.80606f
C139 source.n2 a_n1760_n2688# 0.380471f
C140 source.t17 a_n1760_n2688# 0.215743f
C141 source.t21 a_n1760_n2688# 0.215743f
C142 source.n3 a_n1760_n2688# 1.80606f
C143 source.n4 a_n1760_n2688# 0.380471f
C144 source.t31 a_n1760_n2688# 0.215743f
C145 source.t16 a_n1760_n2688# 0.215743f
C146 source.n5 a_n1760_n2688# 1.80606f
C147 source.n6 a_n1760_n2688# 0.380471f
C148 source.t24 a_n1760_n2688# 2.30058f
C149 source.n7 a_n1760_n2688# 0.471398f
C150 source.t0 a_n1760_n2688# 2.30058f
C151 source.n8 a_n1760_n2688# 0.471398f
C152 source.t6 a_n1760_n2688# 0.215743f
C153 source.t10 a_n1760_n2688# 0.215743f
C154 source.n9 a_n1760_n2688# 1.80606f
C155 source.n10 a_n1760_n2688# 0.380471f
C156 source.t11 a_n1760_n2688# 0.215743f
C157 source.t8 a_n1760_n2688# 0.215743f
C158 source.n11 a_n1760_n2688# 1.80606f
C159 source.n12 a_n1760_n2688# 0.380471f
C160 source.t14 a_n1760_n2688# 0.215743f
C161 source.t7 a_n1760_n2688# 0.215743f
C162 source.n13 a_n1760_n2688# 1.80606f
C163 source.n14 a_n1760_n2688# 0.380471f
C164 source.t13 a_n1760_n2688# 2.30058f
C165 source.n15 a_n1760_n2688# 1.75522f
C166 source.t18 a_n1760_n2688# 2.30057f
C167 source.n16 a_n1760_n2688# 1.75523f
C168 source.t30 a_n1760_n2688# 0.215743f
C169 source.t23 a_n1760_n2688# 0.215743f
C170 source.n17 a_n1760_n2688# 1.80606f
C171 source.n18 a_n1760_n2688# 0.380477f
C172 source.t26 a_n1760_n2688# 0.215743f
C173 source.t28 a_n1760_n2688# 0.215743f
C174 source.n19 a_n1760_n2688# 1.80606f
C175 source.n20 a_n1760_n2688# 0.380477f
C176 source.t20 a_n1760_n2688# 0.215743f
C177 source.t25 a_n1760_n2688# 0.215743f
C178 source.n21 a_n1760_n2688# 1.80606f
C179 source.n22 a_n1760_n2688# 0.380477f
C180 source.t29 a_n1760_n2688# 2.30057f
C181 source.n23 a_n1760_n2688# 0.471404f
C182 source.t5 a_n1760_n2688# 2.30057f
C183 source.n24 a_n1760_n2688# 0.471404f
C184 source.t3 a_n1760_n2688# 0.215743f
C185 source.t4 a_n1760_n2688# 0.215743f
C186 source.n25 a_n1760_n2688# 1.80606f
C187 source.n26 a_n1760_n2688# 0.380477f
C188 source.t9 a_n1760_n2688# 0.215743f
C189 source.t1 a_n1760_n2688# 0.215743f
C190 source.n27 a_n1760_n2688# 1.80606f
C191 source.n28 a_n1760_n2688# 0.380477f
C192 source.t2 a_n1760_n2688# 0.215743f
C193 source.t15 a_n1760_n2688# 0.215743f
C194 source.n29 a_n1760_n2688# 1.80606f
C195 source.n30 a_n1760_n2688# 0.380477f
C196 source.t12 a_n1760_n2688# 2.30057f
C197 source.n31 a_n1760_n2688# 0.639271f
C198 source.n32 a_n1760_n2688# 1.57693f
C199 plus.n0 a_n1760_n2688# 0.053247f
C200 plus.t7 a_n1760_n2688# 0.339484f
C201 plus.t15 a_n1760_n2688# 0.339484f
C202 plus.t8 a_n1760_n2688# 0.339484f
C203 plus.n1 a_n1760_n2688# 0.144498f
C204 plus.n2 a_n1760_n2688# 0.053247f
C205 plus.t0 a_n1760_n2688# 0.339484f
C206 plus.t9 a_n1760_n2688# 0.339484f
C207 plus.n3 a_n1760_n2688# 0.144498f
C208 plus.t6 a_n1760_n2688# 0.345239f
C209 plus.n4 a_n1760_n2688# 0.160093f
C210 plus.t1 a_n1760_n2688# 0.339484f
C211 plus.n5 a_n1760_n2688# 0.144498f
C212 plus.n6 a_n1760_n2688# 0.02029f
C213 plus.n7 a_n1760_n2688# 0.116597f
C214 plus.n8 a_n1760_n2688# 0.053247f
C215 plus.n9 a_n1760_n2688# 0.02029f
C216 plus.n10 a_n1760_n2688# 0.144498f
C217 plus.n11 a_n1760_n2688# 0.018977f
C218 plus.n12 a_n1760_n2688# 0.018977f
C219 plus.n13 a_n1760_n2688# 0.053247f
C220 plus.n14 a_n1760_n2688# 0.053247f
C221 plus.n15 a_n1760_n2688# 0.02029f
C222 plus.n16 a_n1760_n2688# 0.144498f
C223 plus.n17 a_n1760_n2688# 0.02029f
C224 plus.n18 a_n1760_n2688# 0.144498f
C225 plus.t3 a_n1760_n2688# 0.345239f
C226 plus.n19 a_n1760_n2688# 0.160018f
C227 plus.n20 a_n1760_n2688# 0.518704f
C228 plus.n21 a_n1760_n2688# 0.053247f
C229 plus.t4 a_n1760_n2688# 0.345239f
C230 plus.t10 a_n1760_n2688# 0.339484f
C231 plus.t12 a_n1760_n2688# 0.339484f
C232 plus.t2 a_n1760_n2688# 0.339484f
C233 plus.n22 a_n1760_n2688# 0.144498f
C234 plus.n23 a_n1760_n2688# 0.053247f
C235 plus.t14 a_n1760_n2688# 0.339484f
C236 plus.t5 a_n1760_n2688# 0.339484f
C237 plus.n24 a_n1760_n2688# 0.144498f
C238 plus.t13 a_n1760_n2688# 0.345239f
C239 plus.n25 a_n1760_n2688# 0.160093f
C240 plus.t11 a_n1760_n2688# 0.339484f
C241 plus.n26 a_n1760_n2688# 0.144498f
C242 plus.n27 a_n1760_n2688# 0.02029f
C243 plus.n28 a_n1760_n2688# 0.116597f
C244 plus.n29 a_n1760_n2688# 0.053247f
C245 plus.n30 a_n1760_n2688# 0.02029f
C246 plus.n31 a_n1760_n2688# 0.144498f
C247 plus.n32 a_n1760_n2688# 0.018977f
C248 plus.n33 a_n1760_n2688# 0.018977f
C249 plus.n34 a_n1760_n2688# 0.053247f
C250 plus.n35 a_n1760_n2688# 0.053247f
C251 plus.n36 a_n1760_n2688# 0.02029f
C252 plus.n37 a_n1760_n2688# 0.144498f
C253 plus.n38 a_n1760_n2688# 0.02029f
C254 plus.n39 a_n1760_n2688# 0.144498f
C255 plus.n40 a_n1760_n2688# 0.160018f
C256 plus.n41 a_n1760_n2688# 1.44756f
.ends

