* NGSPICE file created from diffpair712.ext - technology: sky130A

.subckt diffpair712 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t7 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.8
X1 a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.8
X2 a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.8
X3 a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.8
X4 a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.8
X5 drain_right.t4 minus.t1 source.t11 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.8
X6 source.t4 plus.t0 drain_left.t5 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.8
X7 source.t6 minus.t2 drain_right.t3 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.8
X8 source.t9 minus.t3 drain_right.t2 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.8
X9 drain_right.t1 minus.t4 source.t8 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.8
X10 drain_left.t4 plus.t1 source.t3 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.8
X11 drain_left.t3 plus.t2 source.t0 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.8
X12 source.t1 plus.t3 drain_left.t2 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.8
X13 drain_right.t0 minus.t5 source.t10 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.8
X14 drain_left.t1 plus.t4 source.t2 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.8
X15 drain_left.t0 plus.t5 source.t5 a_n1620_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.8
R0 minus.n1 minus.t4 825.716
R1 minus.n7 minus.t0 825.716
R2 minus.n2 minus.t2 802.23
R3 minus.n4 minus.t1 802.23
R4 minus.n8 minus.t3 802.23
R5 minus.n10 minus.t5 802.23
R6 minus.n5 minus.n4 161.3
R7 minus.n3 minus.n0 161.3
R8 minus.n11 minus.n10 161.3
R9 minus.n9 minus.n6 161.3
R10 minus.n12 minus.n5 45.3282
R11 minus.n1 minus.n0 44.8973
R12 minus.n7 minus.n6 44.8973
R13 minus.n4 minus.n3 33.5944
R14 minus.n10 minus.n9 33.5944
R15 minus.n2 minus.n1 18.1882
R16 minus.n8 minus.n7 18.1882
R17 minus.n3 minus.n2 14.6066
R18 minus.n9 minus.n8 14.6066
R19 minus.n12 minus.n11 6.72209
R20 minus.n5 minus.n0 0.189894
R21 minus.n11 minus.n6 0.189894
R22 minus minus.n12 0.188
R23 source.n562 source.n428 289.615
R24 source.n420 source.n286 289.615
R25 source.n134 source.n0 289.615
R26 source.n276 source.n142 289.615
R27 source.n472 source.n471 185
R28 source.n477 source.n476 185
R29 source.n479 source.n478 185
R30 source.n468 source.n467 185
R31 source.n485 source.n484 185
R32 source.n487 source.n486 185
R33 source.n464 source.n463 185
R34 source.n494 source.n493 185
R35 source.n495 source.n462 185
R36 source.n497 source.n496 185
R37 source.n460 source.n459 185
R38 source.n503 source.n502 185
R39 source.n505 source.n504 185
R40 source.n456 source.n455 185
R41 source.n511 source.n510 185
R42 source.n513 source.n512 185
R43 source.n452 source.n451 185
R44 source.n519 source.n518 185
R45 source.n521 source.n520 185
R46 source.n448 source.n447 185
R47 source.n527 source.n526 185
R48 source.n529 source.n528 185
R49 source.n444 source.n443 185
R50 source.n535 source.n534 185
R51 source.n538 source.n537 185
R52 source.n536 source.n440 185
R53 source.n543 source.n439 185
R54 source.n545 source.n544 185
R55 source.n547 source.n546 185
R56 source.n436 source.n435 185
R57 source.n553 source.n552 185
R58 source.n555 source.n554 185
R59 source.n432 source.n431 185
R60 source.n561 source.n560 185
R61 source.n563 source.n562 185
R62 source.n330 source.n329 185
R63 source.n335 source.n334 185
R64 source.n337 source.n336 185
R65 source.n326 source.n325 185
R66 source.n343 source.n342 185
R67 source.n345 source.n344 185
R68 source.n322 source.n321 185
R69 source.n352 source.n351 185
R70 source.n353 source.n320 185
R71 source.n355 source.n354 185
R72 source.n318 source.n317 185
R73 source.n361 source.n360 185
R74 source.n363 source.n362 185
R75 source.n314 source.n313 185
R76 source.n369 source.n368 185
R77 source.n371 source.n370 185
R78 source.n310 source.n309 185
R79 source.n377 source.n376 185
R80 source.n379 source.n378 185
R81 source.n306 source.n305 185
R82 source.n385 source.n384 185
R83 source.n387 source.n386 185
R84 source.n302 source.n301 185
R85 source.n393 source.n392 185
R86 source.n396 source.n395 185
R87 source.n394 source.n298 185
R88 source.n401 source.n297 185
R89 source.n403 source.n402 185
R90 source.n405 source.n404 185
R91 source.n294 source.n293 185
R92 source.n411 source.n410 185
R93 source.n413 source.n412 185
R94 source.n290 source.n289 185
R95 source.n419 source.n418 185
R96 source.n421 source.n420 185
R97 source.n135 source.n134 185
R98 source.n133 source.n132 185
R99 source.n4 source.n3 185
R100 source.n127 source.n126 185
R101 source.n125 source.n124 185
R102 source.n8 source.n7 185
R103 source.n119 source.n118 185
R104 source.n117 source.n116 185
R105 source.n115 source.n11 185
R106 source.n15 source.n12 185
R107 source.n110 source.n109 185
R108 source.n108 source.n107 185
R109 source.n17 source.n16 185
R110 source.n102 source.n101 185
R111 source.n100 source.n99 185
R112 source.n21 source.n20 185
R113 source.n94 source.n93 185
R114 source.n92 source.n91 185
R115 source.n25 source.n24 185
R116 source.n86 source.n85 185
R117 source.n84 source.n83 185
R118 source.n29 source.n28 185
R119 source.n78 source.n77 185
R120 source.n76 source.n75 185
R121 source.n33 source.n32 185
R122 source.n70 source.n69 185
R123 source.n68 source.n35 185
R124 source.n67 source.n66 185
R125 source.n38 source.n36 185
R126 source.n61 source.n60 185
R127 source.n59 source.n58 185
R128 source.n42 source.n41 185
R129 source.n53 source.n52 185
R130 source.n51 source.n50 185
R131 source.n46 source.n45 185
R132 source.n277 source.n276 185
R133 source.n275 source.n274 185
R134 source.n146 source.n145 185
R135 source.n269 source.n268 185
R136 source.n267 source.n266 185
R137 source.n150 source.n149 185
R138 source.n261 source.n260 185
R139 source.n259 source.n258 185
R140 source.n257 source.n153 185
R141 source.n157 source.n154 185
R142 source.n252 source.n251 185
R143 source.n250 source.n249 185
R144 source.n159 source.n158 185
R145 source.n244 source.n243 185
R146 source.n242 source.n241 185
R147 source.n163 source.n162 185
R148 source.n236 source.n235 185
R149 source.n234 source.n233 185
R150 source.n167 source.n166 185
R151 source.n228 source.n227 185
R152 source.n226 source.n225 185
R153 source.n171 source.n170 185
R154 source.n220 source.n219 185
R155 source.n218 source.n217 185
R156 source.n175 source.n174 185
R157 source.n212 source.n211 185
R158 source.n210 source.n177 185
R159 source.n209 source.n208 185
R160 source.n180 source.n178 185
R161 source.n203 source.n202 185
R162 source.n201 source.n200 185
R163 source.n184 source.n183 185
R164 source.n195 source.n194 185
R165 source.n193 source.n192 185
R166 source.n188 source.n187 185
R167 source.n473 source.t10 149.524
R168 source.n331 source.t5 149.524
R169 source.n47 source.t3 149.524
R170 source.n189 source.t8 149.524
R171 source.n477 source.n471 104.615
R172 source.n478 source.n477 104.615
R173 source.n478 source.n467 104.615
R174 source.n485 source.n467 104.615
R175 source.n486 source.n485 104.615
R176 source.n486 source.n463 104.615
R177 source.n494 source.n463 104.615
R178 source.n495 source.n494 104.615
R179 source.n496 source.n495 104.615
R180 source.n496 source.n459 104.615
R181 source.n503 source.n459 104.615
R182 source.n504 source.n503 104.615
R183 source.n504 source.n455 104.615
R184 source.n511 source.n455 104.615
R185 source.n512 source.n511 104.615
R186 source.n512 source.n451 104.615
R187 source.n519 source.n451 104.615
R188 source.n520 source.n519 104.615
R189 source.n520 source.n447 104.615
R190 source.n527 source.n447 104.615
R191 source.n528 source.n527 104.615
R192 source.n528 source.n443 104.615
R193 source.n535 source.n443 104.615
R194 source.n537 source.n535 104.615
R195 source.n537 source.n536 104.615
R196 source.n536 source.n439 104.615
R197 source.n545 source.n439 104.615
R198 source.n546 source.n545 104.615
R199 source.n546 source.n435 104.615
R200 source.n553 source.n435 104.615
R201 source.n554 source.n553 104.615
R202 source.n554 source.n431 104.615
R203 source.n561 source.n431 104.615
R204 source.n562 source.n561 104.615
R205 source.n335 source.n329 104.615
R206 source.n336 source.n335 104.615
R207 source.n336 source.n325 104.615
R208 source.n343 source.n325 104.615
R209 source.n344 source.n343 104.615
R210 source.n344 source.n321 104.615
R211 source.n352 source.n321 104.615
R212 source.n353 source.n352 104.615
R213 source.n354 source.n353 104.615
R214 source.n354 source.n317 104.615
R215 source.n361 source.n317 104.615
R216 source.n362 source.n361 104.615
R217 source.n362 source.n313 104.615
R218 source.n369 source.n313 104.615
R219 source.n370 source.n369 104.615
R220 source.n370 source.n309 104.615
R221 source.n377 source.n309 104.615
R222 source.n378 source.n377 104.615
R223 source.n378 source.n305 104.615
R224 source.n385 source.n305 104.615
R225 source.n386 source.n385 104.615
R226 source.n386 source.n301 104.615
R227 source.n393 source.n301 104.615
R228 source.n395 source.n393 104.615
R229 source.n395 source.n394 104.615
R230 source.n394 source.n297 104.615
R231 source.n403 source.n297 104.615
R232 source.n404 source.n403 104.615
R233 source.n404 source.n293 104.615
R234 source.n411 source.n293 104.615
R235 source.n412 source.n411 104.615
R236 source.n412 source.n289 104.615
R237 source.n419 source.n289 104.615
R238 source.n420 source.n419 104.615
R239 source.n134 source.n133 104.615
R240 source.n133 source.n3 104.615
R241 source.n126 source.n3 104.615
R242 source.n126 source.n125 104.615
R243 source.n125 source.n7 104.615
R244 source.n118 source.n7 104.615
R245 source.n118 source.n117 104.615
R246 source.n117 source.n11 104.615
R247 source.n15 source.n11 104.615
R248 source.n109 source.n15 104.615
R249 source.n109 source.n108 104.615
R250 source.n108 source.n16 104.615
R251 source.n101 source.n16 104.615
R252 source.n101 source.n100 104.615
R253 source.n100 source.n20 104.615
R254 source.n93 source.n20 104.615
R255 source.n93 source.n92 104.615
R256 source.n92 source.n24 104.615
R257 source.n85 source.n24 104.615
R258 source.n85 source.n84 104.615
R259 source.n84 source.n28 104.615
R260 source.n77 source.n28 104.615
R261 source.n77 source.n76 104.615
R262 source.n76 source.n32 104.615
R263 source.n69 source.n32 104.615
R264 source.n69 source.n68 104.615
R265 source.n68 source.n67 104.615
R266 source.n67 source.n36 104.615
R267 source.n60 source.n36 104.615
R268 source.n60 source.n59 104.615
R269 source.n59 source.n41 104.615
R270 source.n52 source.n41 104.615
R271 source.n52 source.n51 104.615
R272 source.n51 source.n45 104.615
R273 source.n276 source.n275 104.615
R274 source.n275 source.n145 104.615
R275 source.n268 source.n145 104.615
R276 source.n268 source.n267 104.615
R277 source.n267 source.n149 104.615
R278 source.n260 source.n149 104.615
R279 source.n260 source.n259 104.615
R280 source.n259 source.n153 104.615
R281 source.n157 source.n153 104.615
R282 source.n251 source.n157 104.615
R283 source.n251 source.n250 104.615
R284 source.n250 source.n158 104.615
R285 source.n243 source.n158 104.615
R286 source.n243 source.n242 104.615
R287 source.n242 source.n162 104.615
R288 source.n235 source.n162 104.615
R289 source.n235 source.n234 104.615
R290 source.n234 source.n166 104.615
R291 source.n227 source.n166 104.615
R292 source.n227 source.n226 104.615
R293 source.n226 source.n170 104.615
R294 source.n219 source.n170 104.615
R295 source.n219 source.n218 104.615
R296 source.n218 source.n174 104.615
R297 source.n211 source.n174 104.615
R298 source.n211 source.n210 104.615
R299 source.n210 source.n209 104.615
R300 source.n209 source.n178 104.615
R301 source.n202 source.n178 104.615
R302 source.n202 source.n201 104.615
R303 source.n201 source.n183 104.615
R304 source.n194 source.n183 104.615
R305 source.n194 source.n193 104.615
R306 source.n193 source.n187 104.615
R307 source.t10 source.n471 52.3082
R308 source.t5 source.n329 52.3082
R309 source.t3 source.n45 52.3082
R310 source.t8 source.n187 52.3082
R311 source.n427 source.n426 42.0366
R312 source.n285 source.n284 42.0366
R313 source.n141 source.n140 42.0366
R314 source.n283 source.n282 42.0366
R315 source.n285 source.n283 33.0845
R316 source.n567 source.n566 30.6338
R317 source.n425 source.n424 30.6338
R318 source.n139 source.n138 30.6338
R319 source.n281 source.n280 30.6338
R320 source.n568 source.n139 26.3603
R321 source.n497 source.n462 13.1884
R322 source.n544 source.n543 13.1884
R323 source.n355 source.n320 13.1884
R324 source.n402 source.n401 13.1884
R325 source.n116 source.n115 13.1884
R326 source.n70 source.n35 13.1884
R327 source.n258 source.n257 13.1884
R328 source.n212 source.n177 13.1884
R329 source.n493 source.n492 12.8005
R330 source.n498 source.n460 12.8005
R331 source.n542 source.n440 12.8005
R332 source.n547 source.n438 12.8005
R333 source.n351 source.n350 12.8005
R334 source.n356 source.n318 12.8005
R335 source.n400 source.n298 12.8005
R336 source.n405 source.n296 12.8005
R337 source.n119 source.n10 12.8005
R338 source.n114 source.n12 12.8005
R339 source.n71 source.n33 12.8005
R340 source.n66 source.n37 12.8005
R341 source.n261 source.n152 12.8005
R342 source.n256 source.n154 12.8005
R343 source.n213 source.n175 12.8005
R344 source.n208 source.n179 12.8005
R345 source.n491 source.n464 12.0247
R346 source.n502 source.n501 12.0247
R347 source.n539 source.n538 12.0247
R348 source.n548 source.n436 12.0247
R349 source.n349 source.n322 12.0247
R350 source.n360 source.n359 12.0247
R351 source.n397 source.n396 12.0247
R352 source.n406 source.n294 12.0247
R353 source.n120 source.n8 12.0247
R354 source.n111 source.n110 12.0247
R355 source.n75 source.n74 12.0247
R356 source.n65 source.n38 12.0247
R357 source.n262 source.n150 12.0247
R358 source.n253 source.n252 12.0247
R359 source.n217 source.n216 12.0247
R360 source.n207 source.n180 12.0247
R361 source.n488 source.n487 11.249
R362 source.n505 source.n458 11.249
R363 source.n534 source.n442 11.249
R364 source.n552 source.n551 11.249
R365 source.n346 source.n345 11.249
R366 source.n363 source.n316 11.249
R367 source.n392 source.n300 11.249
R368 source.n410 source.n409 11.249
R369 source.n124 source.n123 11.249
R370 source.n107 source.n14 11.249
R371 source.n78 source.n31 11.249
R372 source.n62 source.n61 11.249
R373 source.n266 source.n265 11.249
R374 source.n249 source.n156 11.249
R375 source.n220 source.n173 11.249
R376 source.n204 source.n203 11.249
R377 source.n484 source.n466 10.4732
R378 source.n506 source.n456 10.4732
R379 source.n533 source.n444 10.4732
R380 source.n555 source.n434 10.4732
R381 source.n342 source.n324 10.4732
R382 source.n364 source.n314 10.4732
R383 source.n391 source.n302 10.4732
R384 source.n413 source.n292 10.4732
R385 source.n127 source.n6 10.4732
R386 source.n106 source.n17 10.4732
R387 source.n79 source.n29 10.4732
R388 source.n58 source.n40 10.4732
R389 source.n269 source.n148 10.4732
R390 source.n248 source.n159 10.4732
R391 source.n221 source.n171 10.4732
R392 source.n200 source.n182 10.4732
R393 source.n473 source.n472 10.2747
R394 source.n331 source.n330 10.2747
R395 source.n47 source.n46 10.2747
R396 source.n189 source.n188 10.2747
R397 source.n483 source.n468 9.69747
R398 source.n510 source.n509 9.69747
R399 source.n530 source.n529 9.69747
R400 source.n556 source.n432 9.69747
R401 source.n341 source.n326 9.69747
R402 source.n368 source.n367 9.69747
R403 source.n388 source.n387 9.69747
R404 source.n414 source.n290 9.69747
R405 source.n128 source.n4 9.69747
R406 source.n103 source.n102 9.69747
R407 source.n83 source.n82 9.69747
R408 source.n57 source.n42 9.69747
R409 source.n270 source.n146 9.69747
R410 source.n245 source.n244 9.69747
R411 source.n225 source.n224 9.69747
R412 source.n199 source.n184 9.69747
R413 source.n566 source.n565 9.45567
R414 source.n424 source.n423 9.45567
R415 source.n138 source.n137 9.45567
R416 source.n280 source.n279 9.45567
R417 source.n430 source.n429 9.3005
R418 source.n559 source.n558 9.3005
R419 source.n557 source.n556 9.3005
R420 source.n434 source.n433 9.3005
R421 source.n551 source.n550 9.3005
R422 source.n549 source.n548 9.3005
R423 source.n438 source.n437 9.3005
R424 source.n517 source.n516 9.3005
R425 source.n515 source.n514 9.3005
R426 source.n454 source.n453 9.3005
R427 source.n509 source.n508 9.3005
R428 source.n507 source.n506 9.3005
R429 source.n458 source.n457 9.3005
R430 source.n501 source.n500 9.3005
R431 source.n499 source.n498 9.3005
R432 source.n475 source.n474 9.3005
R433 source.n470 source.n469 9.3005
R434 source.n481 source.n480 9.3005
R435 source.n483 source.n482 9.3005
R436 source.n466 source.n465 9.3005
R437 source.n489 source.n488 9.3005
R438 source.n491 source.n490 9.3005
R439 source.n492 source.n461 9.3005
R440 source.n450 source.n449 9.3005
R441 source.n523 source.n522 9.3005
R442 source.n525 source.n524 9.3005
R443 source.n446 source.n445 9.3005
R444 source.n531 source.n530 9.3005
R445 source.n533 source.n532 9.3005
R446 source.n442 source.n441 9.3005
R447 source.n540 source.n539 9.3005
R448 source.n542 source.n541 9.3005
R449 source.n565 source.n564 9.3005
R450 source.n288 source.n287 9.3005
R451 source.n417 source.n416 9.3005
R452 source.n415 source.n414 9.3005
R453 source.n292 source.n291 9.3005
R454 source.n409 source.n408 9.3005
R455 source.n407 source.n406 9.3005
R456 source.n296 source.n295 9.3005
R457 source.n375 source.n374 9.3005
R458 source.n373 source.n372 9.3005
R459 source.n312 source.n311 9.3005
R460 source.n367 source.n366 9.3005
R461 source.n365 source.n364 9.3005
R462 source.n316 source.n315 9.3005
R463 source.n359 source.n358 9.3005
R464 source.n357 source.n356 9.3005
R465 source.n333 source.n332 9.3005
R466 source.n328 source.n327 9.3005
R467 source.n339 source.n338 9.3005
R468 source.n341 source.n340 9.3005
R469 source.n324 source.n323 9.3005
R470 source.n347 source.n346 9.3005
R471 source.n349 source.n348 9.3005
R472 source.n350 source.n319 9.3005
R473 source.n308 source.n307 9.3005
R474 source.n381 source.n380 9.3005
R475 source.n383 source.n382 9.3005
R476 source.n304 source.n303 9.3005
R477 source.n389 source.n388 9.3005
R478 source.n391 source.n390 9.3005
R479 source.n300 source.n299 9.3005
R480 source.n398 source.n397 9.3005
R481 source.n400 source.n399 9.3005
R482 source.n423 source.n422 9.3005
R483 source.n49 source.n48 9.3005
R484 source.n44 source.n43 9.3005
R485 source.n55 source.n54 9.3005
R486 source.n57 source.n56 9.3005
R487 source.n40 source.n39 9.3005
R488 source.n63 source.n62 9.3005
R489 source.n65 source.n64 9.3005
R490 source.n37 source.n34 9.3005
R491 source.n96 source.n95 9.3005
R492 source.n98 source.n97 9.3005
R493 source.n19 source.n18 9.3005
R494 source.n104 source.n103 9.3005
R495 source.n106 source.n105 9.3005
R496 source.n14 source.n13 9.3005
R497 source.n112 source.n111 9.3005
R498 source.n114 source.n113 9.3005
R499 source.n137 source.n136 9.3005
R500 source.n2 source.n1 9.3005
R501 source.n131 source.n130 9.3005
R502 source.n129 source.n128 9.3005
R503 source.n6 source.n5 9.3005
R504 source.n123 source.n122 9.3005
R505 source.n121 source.n120 9.3005
R506 source.n10 source.n9 9.3005
R507 source.n23 source.n22 9.3005
R508 source.n90 source.n89 9.3005
R509 source.n88 source.n87 9.3005
R510 source.n27 source.n26 9.3005
R511 source.n82 source.n81 9.3005
R512 source.n80 source.n79 9.3005
R513 source.n31 source.n30 9.3005
R514 source.n74 source.n73 9.3005
R515 source.n72 source.n71 9.3005
R516 source.n191 source.n190 9.3005
R517 source.n186 source.n185 9.3005
R518 source.n197 source.n196 9.3005
R519 source.n199 source.n198 9.3005
R520 source.n182 source.n181 9.3005
R521 source.n205 source.n204 9.3005
R522 source.n207 source.n206 9.3005
R523 source.n179 source.n176 9.3005
R524 source.n238 source.n237 9.3005
R525 source.n240 source.n239 9.3005
R526 source.n161 source.n160 9.3005
R527 source.n246 source.n245 9.3005
R528 source.n248 source.n247 9.3005
R529 source.n156 source.n155 9.3005
R530 source.n254 source.n253 9.3005
R531 source.n256 source.n255 9.3005
R532 source.n279 source.n278 9.3005
R533 source.n144 source.n143 9.3005
R534 source.n273 source.n272 9.3005
R535 source.n271 source.n270 9.3005
R536 source.n148 source.n147 9.3005
R537 source.n265 source.n264 9.3005
R538 source.n263 source.n262 9.3005
R539 source.n152 source.n151 9.3005
R540 source.n165 source.n164 9.3005
R541 source.n232 source.n231 9.3005
R542 source.n230 source.n229 9.3005
R543 source.n169 source.n168 9.3005
R544 source.n224 source.n223 9.3005
R545 source.n222 source.n221 9.3005
R546 source.n173 source.n172 9.3005
R547 source.n216 source.n215 9.3005
R548 source.n214 source.n213 9.3005
R549 source.n480 source.n479 8.92171
R550 source.n513 source.n454 8.92171
R551 source.n526 source.n446 8.92171
R552 source.n560 source.n559 8.92171
R553 source.n338 source.n337 8.92171
R554 source.n371 source.n312 8.92171
R555 source.n384 source.n304 8.92171
R556 source.n418 source.n417 8.92171
R557 source.n132 source.n131 8.92171
R558 source.n99 source.n19 8.92171
R559 source.n86 source.n27 8.92171
R560 source.n54 source.n53 8.92171
R561 source.n274 source.n273 8.92171
R562 source.n241 source.n161 8.92171
R563 source.n228 source.n169 8.92171
R564 source.n196 source.n195 8.92171
R565 source.n476 source.n470 8.14595
R566 source.n514 source.n452 8.14595
R567 source.n525 source.n448 8.14595
R568 source.n563 source.n430 8.14595
R569 source.n334 source.n328 8.14595
R570 source.n372 source.n310 8.14595
R571 source.n383 source.n306 8.14595
R572 source.n421 source.n288 8.14595
R573 source.n135 source.n2 8.14595
R574 source.n98 source.n21 8.14595
R575 source.n87 source.n25 8.14595
R576 source.n50 source.n44 8.14595
R577 source.n277 source.n144 8.14595
R578 source.n240 source.n163 8.14595
R579 source.n229 source.n167 8.14595
R580 source.n192 source.n186 8.14595
R581 source.n475 source.n472 7.3702
R582 source.n518 source.n517 7.3702
R583 source.n522 source.n521 7.3702
R584 source.n564 source.n428 7.3702
R585 source.n333 source.n330 7.3702
R586 source.n376 source.n375 7.3702
R587 source.n380 source.n379 7.3702
R588 source.n422 source.n286 7.3702
R589 source.n136 source.n0 7.3702
R590 source.n95 source.n94 7.3702
R591 source.n91 source.n90 7.3702
R592 source.n49 source.n46 7.3702
R593 source.n278 source.n142 7.3702
R594 source.n237 source.n236 7.3702
R595 source.n233 source.n232 7.3702
R596 source.n191 source.n188 7.3702
R597 source.n518 source.n450 6.59444
R598 source.n521 source.n450 6.59444
R599 source.n566 source.n428 6.59444
R600 source.n376 source.n308 6.59444
R601 source.n379 source.n308 6.59444
R602 source.n424 source.n286 6.59444
R603 source.n138 source.n0 6.59444
R604 source.n94 source.n23 6.59444
R605 source.n91 source.n23 6.59444
R606 source.n280 source.n142 6.59444
R607 source.n236 source.n165 6.59444
R608 source.n233 source.n165 6.59444
R609 source.n476 source.n475 5.81868
R610 source.n517 source.n452 5.81868
R611 source.n522 source.n448 5.81868
R612 source.n564 source.n563 5.81868
R613 source.n334 source.n333 5.81868
R614 source.n375 source.n310 5.81868
R615 source.n380 source.n306 5.81868
R616 source.n422 source.n421 5.81868
R617 source.n136 source.n135 5.81868
R618 source.n95 source.n21 5.81868
R619 source.n90 source.n25 5.81868
R620 source.n50 source.n49 5.81868
R621 source.n278 source.n277 5.81868
R622 source.n237 source.n163 5.81868
R623 source.n232 source.n167 5.81868
R624 source.n192 source.n191 5.81868
R625 source.n568 source.n567 5.7505
R626 source.n479 source.n470 5.04292
R627 source.n514 source.n513 5.04292
R628 source.n526 source.n525 5.04292
R629 source.n560 source.n430 5.04292
R630 source.n337 source.n328 5.04292
R631 source.n372 source.n371 5.04292
R632 source.n384 source.n383 5.04292
R633 source.n418 source.n288 5.04292
R634 source.n132 source.n2 5.04292
R635 source.n99 source.n98 5.04292
R636 source.n87 source.n86 5.04292
R637 source.n53 source.n44 5.04292
R638 source.n274 source.n144 5.04292
R639 source.n241 source.n240 5.04292
R640 source.n229 source.n228 5.04292
R641 source.n195 source.n186 5.04292
R642 source.n480 source.n468 4.26717
R643 source.n510 source.n454 4.26717
R644 source.n529 source.n446 4.26717
R645 source.n559 source.n432 4.26717
R646 source.n338 source.n326 4.26717
R647 source.n368 source.n312 4.26717
R648 source.n387 source.n304 4.26717
R649 source.n417 source.n290 4.26717
R650 source.n131 source.n4 4.26717
R651 source.n102 source.n19 4.26717
R652 source.n83 source.n27 4.26717
R653 source.n54 source.n42 4.26717
R654 source.n273 source.n146 4.26717
R655 source.n244 source.n161 4.26717
R656 source.n225 source.n169 4.26717
R657 source.n196 source.n184 4.26717
R658 source.n484 source.n483 3.49141
R659 source.n509 source.n456 3.49141
R660 source.n530 source.n444 3.49141
R661 source.n556 source.n555 3.49141
R662 source.n342 source.n341 3.49141
R663 source.n367 source.n314 3.49141
R664 source.n388 source.n302 3.49141
R665 source.n414 source.n413 3.49141
R666 source.n128 source.n127 3.49141
R667 source.n103 source.n17 3.49141
R668 source.n82 source.n29 3.49141
R669 source.n58 source.n57 3.49141
R670 source.n270 source.n269 3.49141
R671 source.n245 source.n159 3.49141
R672 source.n224 source.n171 3.49141
R673 source.n200 source.n199 3.49141
R674 source.n48 source.n47 2.84303
R675 source.n190 source.n189 2.84303
R676 source.n474 source.n473 2.84303
R677 source.n332 source.n331 2.84303
R678 source.n487 source.n466 2.71565
R679 source.n506 source.n505 2.71565
R680 source.n534 source.n533 2.71565
R681 source.n552 source.n434 2.71565
R682 source.n345 source.n324 2.71565
R683 source.n364 source.n363 2.71565
R684 source.n392 source.n391 2.71565
R685 source.n410 source.n292 2.71565
R686 source.n124 source.n6 2.71565
R687 source.n107 source.n106 2.71565
R688 source.n79 source.n78 2.71565
R689 source.n61 source.n40 2.71565
R690 source.n266 source.n148 2.71565
R691 source.n249 source.n248 2.71565
R692 source.n221 source.n220 2.71565
R693 source.n203 source.n182 2.71565
R694 source.n488 source.n464 1.93989
R695 source.n502 source.n458 1.93989
R696 source.n538 source.n442 1.93989
R697 source.n551 source.n436 1.93989
R698 source.n346 source.n322 1.93989
R699 source.n360 source.n316 1.93989
R700 source.n396 source.n300 1.93989
R701 source.n409 source.n294 1.93989
R702 source.n123 source.n8 1.93989
R703 source.n110 source.n14 1.93989
R704 source.n75 source.n31 1.93989
R705 source.n62 source.n38 1.93989
R706 source.n265 source.n150 1.93989
R707 source.n252 source.n156 1.93989
R708 source.n217 source.n173 1.93989
R709 source.n204 source.n180 1.93989
R710 source.n493 source.n491 1.16414
R711 source.n501 source.n460 1.16414
R712 source.n539 source.n440 1.16414
R713 source.n548 source.n547 1.16414
R714 source.n351 source.n349 1.16414
R715 source.n359 source.n318 1.16414
R716 source.n397 source.n298 1.16414
R717 source.n406 source.n405 1.16414
R718 source.n120 source.n119 1.16414
R719 source.n111 source.n12 1.16414
R720 source.n74 source.n33 1.16414
R721 source.n66 source.n65 1.16414
R722 source.n262 source.n261 1.16414
R723 source.n253 source.n154 1.16414
R724 source.n216 source.n175 1.16414
R725 source.n208 source.n207 1.16414
R726 source.n283 source.n281 0.974638
R727 source.n141 source.n139 0.974638
R728 source.n425 source.n285 0.974638
R729 source.n567 source.n427 0.974638
R730 source.n281 source.n141 0.957397
R731 source.n427 source.n425 0.957397
R732 source.n426 source.t7 0.7925
R733 source.n426 source.t9 0.7925
R734 source.n284 source.t0 0.7925
R735 source.n284 source.t4 0.7925
R736 source.n140 source.t2 0.7925
R737 source.n140 source.t1 0.7925
R738 source.n282 source.t11 0.7925
R739 source.n282 source.t6 0.7925
R740 source.n492 source.n462 0.388379
R741 source.n498 source.n497 0.388379
R742 source.n543 source.n542 0.388379
R743 source.n544 source.n438 0.388379
R744 source.n350 source.n320 0.388379
R745 source.n356 source.n355 0.388379
R746 source.n401 source.n400 0.388379
R747 source.n402 source.n296 0.388379
R748 source.n116 source.n10 0.388379
R749 source.n115 source.n114 0.388379
R750 source.n71 source.n70 0.388379
R751 source.n37 source.n35 0.388379
R752 source.n258 source.n152 0.388379
R753 source.n257 source.n256 0.388379
R754 source.n213 source.n212 0.388379
R755 source.n179 source.n177 0.388379
R756 source source.n568 0.188
R757 source.n474 source.n469 0.155672
R758 source.n481 source.n469 0.155672
R759 source.n482 source.n481 0.155672
R760 source.n482 source.n465 0.155672
R761 source.n489 source.n465 0.155672
R762 source.n490 source.n489 0.155672
R763 source.n490 source.n461 0.155672
R764 source.n499 source.n461 0.155672
R765 source.n500 source.n499 0.155672
R766 source.n500 source.n457 0.155672
R767 source.n507 source.n457 0.155672
R768 source.n508 source.n507 0.155672
R769 source.n508 source.n453 0.155672
R770 source.n515 source.n453 0.155672
R771 source.n516 source.n515 0.155672
R772 source.n516 source.n449 0.155672
R773 source.n523 source.n449 0.155672
R774 source.n524 source.n523 0.155672
R775 source.n524 source.n445 0.155672
R776 source.n531 source.n445 0.155672
R777 source.n532 source.n531 0.155672
R778 source.n532 source.n441 0.155672
R779 source.n540 source.n441 0.155672
R780 source.n541 source.n540 0.155672
R781 source.n541 source.n437 0.155672
R782 source.n549 source.n437 0.155672
R783 source.n550 source.n549 0.155672
R784 source.n550 source.n433 0.155672
R785 source.n557 source.n433 0.155672
R786 source.n558 source.n557 0.155672
R787 source.n558 source.n429 0.155672
R788 source.n565 source.n429 0.155672
R789 source.n332 source.n327 0.155672
R790 source.n339 source.n327 0.155672
R791 source.n340 source.n339 0.155672
R792 source.n340 source.n323 0.155672
R793 source.n347 source.n323 0.155672
R794 source.n348 source.n347 0.155672
R795 source.n348 source.n319 0.155672
R796 source.n357 source.n319 0.155672
R797 source.n358 source.n357 0.155672
R798 source.n358 source.n315 0.155672
R799 source.n365 source.n315 0.155672
R800 source.n366 source.n365 0.155672
R801 source.n366 source.n311 0.155672
R802 source.n373 source.n311 0.155672
R803 source.n374 source.n373 0.155672
R804 source.n374 source.n307 0.155672
R805 source.n381 source.n307 0.155672
R806 source.n382 source.n381 0.155672
R807 source.n382 source.n303 0.155672
R808 source.n389 source.n303 0.155672
R809 source.n390 source.n389 0.155672
R810 source.n390 source.n299 0.155672
R811 source.n398 source.n299 0.155672
R812 source.n399 source.n398 0.155672
R813 source.n399 source.n295 0.155672
R814 source.n407 source.n295 0.155672
R815 source.n408 source.n407 0.155672
R816 source.n408 source.n291 0.155672
R817 source.n415 source.n291 0.155672
R818 source.n416 source.n415 0.155672
R819 source.n416 source.n287 0.155672
R820 source.n423 source.n287 0.155672
R821 source.n137 source.n1 0.155672
R822 source.n130 source.n1 0.155672
R823 source.n130 source.n129 0.155672
R824 source.n129 source.n5 0.155672
R825 source.n122 source.n5 0.155672
R826 source.n122 source.n121 0.155672
R827 source.n121 source.n9 0.155672
R828 source.n113 source.n9 0.155672
R829 source.n113 source.n112 0.155672
R830 source.n112 source.n13 0.155672
R831 source.n105 source.n13 0.155672
R832 source.n105 source.n104 0.155672
R833 source.n104 source.n18 0.155672
R834 source.n97 source.n18 0.155672
R835 source.n97 source.n96 0.155672
R836 source.n96 source.n22 0.155672
R837 source.n89 source.n22 0.155672
R838 source.n89 source.n88 0.155672
R839 source.n88 source.n26 0.155672
R840 source.n81 source.n26 0.155672
R841 source.n81 source.n80 0.155672
R842 source.n80 source.n30 0.155672
R843 source.n73 source.n30 0.155672
R844 source.n73 source.n72 0.155672
R845 source.n72 source.n34 0.155672
R846 source.n64 source.n34 0.155672
R847 source.n64 source.n63 0.155672
R848 source.n63 source.n39 0.155672
R849 source.n56 source.n39 0.155672
R850 source.n56 source.n55 0.155672
R851 source.n55 source.n43 0.155672
R852 source.n48 source.n43 0.155672
R853 source.n279 source.n143 0.155672
R854 source.n272 source.n143 0.155672
R855 source.n272 source.n271 0.155672
R856 source.n271 source.n147 0.155672
R857 source.n264 source.n147 0.155672
R858 source.n264 source.n263 0.155672
R859 source.n263 source.n151 0.155672
R860 source.n255 source.n151 0.155672
R861 source.n255 source.n254 0.155672
R862 source.n254 source.n155 0.155672
R863 source.n247 source.n155 0.155672
R864 source.n247 source.n246 0.155672
R865 source.n246 source.n160 0.155672
R866 source.n239 source.n160 0.155672
R867 source.n239 source.n238 0.155672
R868 source.n238 source.n164 0.155672
R869 source.n231 source.n164 0.155672
R870 source.n231 source.n230 0.155672
R871 source.n230 source.n168 0.155672
R872 source.n223 source.n168 0.155672
R873 source.n223 source.n222 0.155672
R874 source.n222 source.n172 0.155672
R875 source.n215 source.n172 0.155672
R876 source.n215 source.n214 0.155672
R877 source.n214 source.n176 0.155672
R878 source.n206 source.n176 0.155672
R879 source.n206 source.n205 0.155672
R880 source.n205 source.n181 0.155672
R881 source.n198 source.n181 0.155672
R882 source.n198 source.n197 0.155672
R883 source.n197 source.n185 0.155672
R884 source.n190 source.n185 0.155672
R885 drain_right.n134 drain_right.n0 289.615
R886 drain_right.n276 drain_right.n142 289.615
R887 drain_right.n44 drain_right.n43 185
R888 drain_right.n49 drain_right.n48 185
R889 drain_right.n51 drain_right.n50 185
R890 drain_right.n40 drain_right.n39 185
R891 drain_right.n57 drain_right.n56 185
R892 drain_right.n59 drain_right.n58 185
R893 drain_right.n36 drain_right.n35 185
R894 drain_right.n66 drain_right.n65 185
R895 drain_right.n67 drain_right.n34 185
R896 drain_right.n69 drain_right.n68 185
R897 drain_right.n32 drain_right.n31 185
R898 drain_right.n75 drain_right.n74 185
R899 drain_right.n77 drain_right.n76 185
R900 drain_right.n28 drain_right.n27 185
R901 drain_right.n83 drain_right.n82 185
R902 drain_right.n85 drain_right.n84 185
R903 drain_right.n24 drain_right.n23 185
R904 drain_right.n91 drain_right.n90 185
R905 drain_right.n93 drain_right.n92 185
R906 drain_right.n20 drain_right.n19 185
R907 drain_right.n99 drain_right.n98 185
R908 drain_right.n101 drain_right.n100 185
R909 drain_right.n16 drain_right.n15 185
R910 drain_right.n107 drain_right.n106 185
R911 drain_right.n110 drain_right.n109 185
R912 drain_right.n108 drain_right.n12 185
R913 drain_right.n115 drain_right.n11 185
R914 drain_right.n117 drain_right.n116 185
R915 drain_right.n119 drain_right.n118 185
R916 drain_right.n8 drain_right.n7 185
R917 drain_right.n125 drain_right.n124 185
R918 drain_right.n127 drain_right.n126 185
R919 drain_right.n4 drain_right.n3 185
R920 drain_right.n133 drain_right.n132 185
R921 drain_right.n135 drain_right.n134 185
R922 drain_right.n277 drain_right.n276 185
R923 drain_right.n275 drain_right.n274 185
R924 drain_right.n146 drain_right.n145 185
R925 drain_right.n269 drain_right.n268 185
R926 drain_right.n267 drain_right.n266 185
R927 drain_right.n150 drain_right.n149 185
R928 drain_right.n261 drain_right.n260 185
R929 drain_right.n259 drain_right.n258 185
R930 drain_right.n257 drain_right.n153 185
R931 drain_right.n157 drain_right.n154 185
R932 drain_right.n252 drain_right.n251 185
R933 drain_right.n250 drain_right.n249 185
R934 drain_right.n159 drain_right.n158 185
R935 drain_right.n244 drain_right.n243 185
R936 drain_right.n242 drain_right.n241 185
R937 drain_right.n163 drain_right.n162 185
R938 drain_right.n236 drain_right.n235 185
R939 drain_right.n234 drain_right.n233 185
R940 drain_right.n167 drain_right.n166 185
R941 drain_right.n228 drain_right.n227 185
R942 drain_right.n226 drain_right.n225 185
R943 drain_right.n171 drain_right.n170 185
R944 drain_right.n220 drain_right.n219 185
R945 drain_right.n218 drain_right.n217 185
R946 drain_right.n175 drain_right.n174 185
R947 drain_right.n212 drain_right.n211 185
R948 drain_right.n210 drain_right.n177 185
R949 drain_right.n209 drain_right.n208 185
R950 drain_right.n180 drain_right.n178 185
R951 drain_right.n203 drain_right.n202 185
R952 drain_right.n201 drain_right.n200 185
R953 drain_right.n184 drain_right.n183 185
R954 drain_right.n195 drain_right.n194 185
R955 drain_right.n193 drain_right.n192 185
R956 drain_right.n188 drain_right.n187 185
R957 drain_right.n45 drain_right.t5 149.524
R958 drain_right.n189 drain_right.t4 149.524
R959 drain_right.n49 drain_right.n43 104.615
R960 drain_right.n50 drain_right.n49 104.615
R961 drain_right.n50 drain_right.n39 104.615
R962 drain_right.n57 drain_right.n39 104.615
R963 drain_right.n58 drain_right.n57 104.615
R964 drain_right.n58 drain_right.n35 104.615
R965 drain_right.n66 drain_right.n35 104.615
R966 drain_right.n67 drain_right.n66 104.615
R967 drain_right.n68 drain_right.n67 104.615
R968 drain_right.n68 drain_right.n31 104.615
R969 drain_right.n75 drain_right.n31 104.615
R970 drain_right.n76 drain_right.n75 104.615
R971 drain_right.n76 drain_right.n27 104.615
R972 drain_right.n83 drain_right.n27 104.615
R973 drain_right.n84 drain_right.n83 104.615
R974 drain_right.n84 drain_right.n23 104.615
R975 drain_right.n91 drain_right.n23 104.615
R976 drain_right.n92 drain_right.n91 104.615
R977 drain_right.n92 drain_right.n19 104.615
R978 drain_right.n99 drain_right.n19 104.615
R979 drain_right.n100 drain_right.n99 104.615
R980 drain_right.n100 drain_right.n15 104.615
R981 drain_right.n107 drain_right.n15 104.615
R982 drain_right.n109 drain_right.n107 104.615
R983 drain_right.n109 drain_right.n108 104.615
R984 drain_right.n108 drain_right.n11 104.615
R985 drain_right.n117 drain_right.n11 104.615
R986 drain_right.n118 drain_right.n117 104.615
R987 drain_right.n118 drain_right.n7 104.615
R988 drain_right.n125 drain_right.n7 104.615
R989 drain_right.n126 drain_right.n125 104.615
R990 drain_right.n126 drain_right.n3 104.615
R991 drain_right.n133 drain_right.n3 104.615
R992 drain_right.n134 drain_right.n133 104.615
R993 drain_right.n276 drain_right.n275 104.615
R994 drain_right.n275 drain_right.n145 104.615
R995 drain_right.n268 drain_right.n145 104.615
R996 drain_right.n268 drain_right.n267 104.615
R997 drain_right.n267 drain_right.n149 104.615
R998 drain_right.n260 drain_right.n149 104.615
R999 drain_right.n260 drain_right.n259 104.615
R1000 drain_right.n259 drain_right.n153 104.615
R1001 drain_right.n157 drain_right.n153 104.615
R1002 drain_right.n251 drain_right.n157 104.615
R1003 drain_right.n251 drain_right.n250 104.615
R1004 drain_right.n250 drain_right.n158 104.615
R1005 drain_right.n243 drain_right.n158 104.615
R1006 drain_right.n243 drain_right.n242 104.615
R1007 drain_right.n242 drain_right.n162 104.615
R1008 drain_right.n235 drain_right.n162 104.615
R1009 drain_right.n235 drain_right.n234 104.615
R1010 drain_right.n234 drain_right.n166 104.615
R1011 drain_right.n227 drain_right.n166 104.615
R1012 drain_right.n227 drain_right.n226 104.615
R1013 drain_right.n226 drain_right.n170 104.615
R1014 drain_right.n219 drain_right.n170 104.615
R1015 drain_right.n219 drain_right.n218 104.615
R1016 drain_right.n218 drain_right.n174 104.615
R1017 drain_right.n211 drain_right.n174 104.615
R1018 drain_right.n211 drain_right.n210 104.615
R1019 drain_right.n210 drain_right.n209 104.615
R1020 drain_right.n209 drain_right.n178 104.615
R1021 drain_right.n202 drain_right.n178 104.615
R1022 drain_right.n202 drain_right.n201 104.615
R1023 drain_right.n201 drain_right.n183 104.615
R1024 drain_right.n194 drain_right.n183 104.615
R1025 drain_right.n194 drain_right.n193 104.615
R1026 drain_right.n193 drain_right.n187 104.615
R1027 drain_right.n281 drain_right.n141 59.6894
R1028 drain_right.n140 drain_right.n139 58.9036
R1029 drain_right.t5 drain_right.n43 52.3082
R1030 drain_right.t4 drain_right.n187 52.3082
R1031 drain_right.n140 drain_right.n138 47.9879
R1032 drain_right.n281 drain_right.n280 47.3126
R1033 drain_right drain_right.n140 39.3412
R1034 drain_right.n69 drain_right.n34 13.1884
R1035 drain_right.n116 drain_right.n115 13.1884
R1036 drain_right.n258 drain_right.n257 13.1884
R1037 drain_right.n212 drain_right.n177 13.1884
R1038 drain_right.n65 drain_right.n64 12.8005
R1039 drain_right.n70 drain_right.n32 12.8005
R1040 drain_right.n114 drain_right.n12 12.8005
R1041 drain_right.n119 drain_right.n10 12.8005
R1042 drain_right.n261 drain_right.n152 12.8005
R1043 drain_right.n256 drain_right.n154 12.8005
R1044 drain_right.n213 drain_right.n175 12.8005
R1045 drain_right.n208 drain_right.n179 12.8005
R1046 drain_right.n63 drain_right.n36 12.0247
R1047 drain_right.n74 drain_right.n73 12.0247
R1048 drain_right.n111 drain_right.n110 12.0247
R1049 drain_right.n120 drain_right.n8 12.0247
R1050 drain_right.n262 drain_right.n150 12.0247
R1051 drain_right.n253 drain_right.n252 12.0247
R1052 drain_right.n217 drain_right.n216 12.0247
R1053 drain_right.n207 drain_right.n180 12.0247
R1054 drain_right.n60 drain_right.n59 11.249
R1055 drain_right.n77 drain_right.n30 11.249
R1056 drain_right.n106 drain_right.n14 11.249
R1057 drain_right.n124 drain_right.n123 11.249
R1058 drain_right.n266 drain_right.n265 11.249
R1059 drain_right.n249 drain_right.n156 11.249
R1060 drain_right.n220 drain_right.n173 11.249
R1061 drain_right.n204 drain_right.n203 11.249
R1062 drain_right.n56 drain_right.n38 10.4732
R1063 drain_right.n78 drain_right.n28 10.4732
R1064 drain_right.n105 drain_right.n16 10.4732
R1065 drain_right.n127 drain_right.n6 10.4732
R1066 drain_right.n269 drain_right.n148 10.4732
R1067 drain_right.n248 drain_right.n159 10.4732
R1068 drain_right.n221 drain_right.n171 10.4732
R1069 drain_right.n200 drain_right.n182 10.4732
R1070 drain_right.n45 drain_right.n44 10.2747
R1071 drain_right.n189 drain_right.n188 10.2747
R1072 drain_right.n55 drain_right.n40 9.69747
R1073 drain_right.n82 drain_right.n81 9.69747
R1074 drain_right.n102 drain_right.n101 9.69747
R1075 drain_right.n128 drain_right.n4 9.69747
R1076 drain_right.n270 drain_right.n146 9.69747
R1077 drain_right.n245 drain_right.n244 9.69747
R1078 drain_right.n225 drain_right.n224 9.69747
R1079 drain_right.n199 drain_right.n184 9.69747
R1080 drain_right.n138 drain_right.n137 9.45567
R1081 drain_right.n280 drain_right.n279 9.45567
R1082 drain_right.n2 drain_right.n1 9.3005
R1083 drain_right.n131 drain_right.n130 9.3005
R1084 drain_right.n129 drain_right.n128 9.3005
R1085 drain_right.n6 drain_right.n5 9.3005
R1086 drain_right.n123 drain_right.n122 9.3005
R1087 drain_right.n121 drain_right.n120 9.3005
R1088 drain_right.n10 drain_right.n9 9.3005
R1089 drain_right.n89 drain_right.n88 9.3005
R1090 drain_right.n87 drain_right.n86 9.3005
R1091 drain_right.n26 drain_right.n25 9.3005
R1092 drain_right.n81 drain_right.n80 9.3005
R1093 drain_right.n79 drain_right.n78 9.3005
R1094 drain_right.n30 drain_right.n29 9.3005
R1095 drain_right.n73 drain_right.n72 9.3005
R1096 drain_right.n71 drain_right.n70 9.3005
R1097 drain_right.n47 drain_right.n46 9.3005
R1098 drain_right.n42 drain_right.n41 9.3005
R1099 drain_right.n53 drain_right.n52 9.3005
R1100 drain_right.n55 drain_right.n54 9.3005
R1101 drain_right.n38 drain_right.n37 9.3005
R1102 drain_right.n61 drain_right.n60 9.3005
R1103 drain_right.n63 drain_right.n62 9.3005
R1104 drain_right.n64 drain_right.n33 9.3005
R1105 drain_right.n22 drain_right.n21 9.3005
R1106 drain_right.n95 drain_right.n94 9.3005
R1107 drain_right.n97 drain_right.n96 9.3005
R1108 drain_right.n18 drain_right.n17 9.3005
R1109 drain_right.n103 drain_right.n102 9.3005
R1110 drain_right.n105 drain_right.n104 9.3005
R1111 drain_right.n14 drain_right.n13 9.3005
R1112 drain_right.n112 drain_right.n111 9.3005
R1113 drain_right.n114 drain_right.n113 9.3005
R1114 drain_right.n137 drain_right.n136 9.3005
R1115 drain_right.n191 drain_right.n190 9.3005
R1116 drain_right.n186 drain_right.n185 9.3005
R1117 drain_right.n197 drain_right.n196 9.3005
R1118 drain_right.n199 drain_right.n198 9.3005
R1119 drain_right.n182 drain_right.n181 9.3005
R1120 drain_right.n205 drain_right.n204 9.3005
R1121 drain_right.n207 drain_right.n206 9.3005
R1122 drain_right.n179 drain_right.n176 9.3005
R1123 drain_right.n238 drain_right.n237 9.3005
R1124 drain_right.n240 drain_right.n239 9.3005
R1125 drain_right.n161 drain_right.n160 9.3005
R1126 drain_right.n246 drain_right.n245 9.3005
R1127 drain_right.n248 drain_right.n247 9.3005
R1128 drain_right.n156 drain_right.n155 9.3005
R1129 drain_right.n254 drain_right.n253 9.3005
R1130 drain_right.n256 drain_right.n255 9.3005
R1131 drain_right.n279 drain_right.n278 9.3005
R1132 drain_right.n144 drain_right.n143 9.3005
R1133 drain_right.n273 drain_right.n272 9.3005
R1134 drain_right.n271 drain_right.n270 9.3005
R1135 drain_right.n148 drain_right.n147 9.3005
R1136 drain_right.n265 drain_right.n264 9.3005
R1137 drain_right.n263 drain_right.n262 9.3005
R1138 drain_right.n152 drain_right.n151 9.3005
R1139 drain_right.n165 drain_right.n164 9.3005
R1140 drain_right.n232 drain_right.n231 9.3005
R1141 drain_right.n230 drain_right.n229 9.3005
R1142 drain_right.n169 drain_right.n168 9.3005
R1143 drain_right.n224 drain_right.n223 9.3005
R1144 drain_right.n222 drain_right.n221 9.3005
R1145 drain_right.n173 drain_right.n172 9.3005
R1146 drain_right.n216 drain_right.n215 9.3005
R1147 drain_right.n214 drain_right.n213 9.3005
R1148 drain_right.n52 drain_right.n51 8.92171
R1149 drain_right.n85 drain_right.n26 8.92171
R1150 drain_right.n98 drain_right.n18 8.92171
R1151 drain_right.n132 drain_right.n131 8.92171
R1152 drain_right.n274 drain_right.n273 8.92171
R1153 drain_right.n241 drain_right.n161 8.92171
R1154 drain_right.n228 drain_right.n169 8.92171
R1155 drain_right.n196 drain_right.n195 8.92171
R1156 drain_right.n48 drain_right.n42 8.14595
R1157 drain_right.n86 drain_right.n24 8.14595
R1158 drain_right.n97 drain_right.n20 8.14595
R1159 drain_right.n135 drain_right.n2 8.14595
R1160 drain_right.n277 drain_right.n144 8.14595
R1161 drain_right.n240 drain_right.n163 8.14595
R1162 drain_right.n229 drain_right.n167 8.14595
R1163 drain_right.n192 drain_right.n186 8.14595
R1164 drain_right.n47 drain_right.n44 7.3702
R1165 drain_right.n90 drain_right.n89 7.3702
R1166 drain_right.n94 drain_right.n93 7.3702
R1167 drain_right.n136 drain_right.n0 7.3702
R1168 drain_right.n278 drain_right.n142 7.3702
R1169 drain_right.n237 drain_right.n236 7.3702
R1170 drain_right.n233 drain_right.n232 7.3702
R1171 drain_right.n191 drain_right.n188 7.3702
R1172 drain_right.n90 drain_right.n22 6.59444
R1173 drain_right.n93 drain_right.n22 6.59444
R1174 drain_right.n138 drain_right.n0 6.59444
R1175 drain_right.n280 drain_right.n142 6.59444
R1176 drain_right.n236 drain_right.n165 6.59444
R1177 drain_right.n233 drain_right.n165 6.59444
R1178 drain_right drain_right.n281 6.14028
R1179 drain_right.n48 drain_right.n47 5.81868
R1180 drain_right.n89 drain_right.n24 5.81868
R1181 drain_right.n94 drain_right.n20 5.81868
R1182 drain_right.n136 drain_right.n135 5.81868
R1183 drain_right.n278 drain_right.n277 5.81868
R1184 drain_right.n237 drain_right.n163 5.81868
R1185 drain_right.n232 drain_right.n167 5.81868
R1186 drain_right.n192 drain_right.n191 5.81868
R1187 drain_right.n51 drain_right.n42 5.04292
R1188 drain_right.n86 drain_right.n85 5.04292
R1189 drain_right.n98 drain_right.n97 5.04292
R1190 drain_right.n132 drain_right.n2 5.04292
R1191 drain_right.n274 drain_right.n144 5.04292
R1192 drain_right.n241 drain_right.n240 5.04292
R1193 drain_right.n229 drain_right.n228 5.04292
R1194 drain_right.n195 drain_right.n186 5.04292
R1195 drain_right.n52 drain_right.n40 4.26717
R1196 drain_right.n82 drain_right.n26 4.26717
R1197 drain_right.n101 drain_right.n18 4.26717
R1198 drain_right.n131 drain_right.n4 4.26717
R1199 drain_right.n273 drain_right.n146 4.26717
R1200 drain_right.n244 drain_right.n161 4.26717
R1201 drain_right.n225 drain_right.n169 4.26717
R1202 drain_right.n196 drain_right.n184 4.26717
R1203 drain_right.n56 drain_right.n55 3.49141
R1204 drain_right.n81 drain_right.n28 3.49141
R1205 drain_right.n102 drain_right.n16 3.49141
R1206 drain_right.n128 drain_right.n127 3.49141
R1207 drain_right.n270 drain_right.n269 3.49141
R1208 drain_right.n245 drain_right.n159 3.49141
R1209 drain_right.n224 drain_right.n171 3.49141
R1210 drain_right.n200 drain_right.n199 3.49141
R1211 drain_right.n190 drain_right.n189 2.84303
R1212 drain_right.n46 drain_right.n45 2.84303
R1213 drain_right.n59 drain_right.n38 2.71565
R1214 drain_right.n78 drain_right.n77 2.71565
R1215 drain_right.n106 drain_right.n105 2.71565
R1216 drain_right.n124 drain_right.n6 2.71565
R1217 drain_right.n266 drain_right.n148 2.71565
R1218 drain_right.n249 drain_right.n248 2.71565
R1219 drain_right.n221 drain_right.n220 2.71565
R1220 drain_right.n203 drain_right.n182 2.71565
R1221 drain_right.n60 drain_right.n36 1.93989
R1222 drain_right.n74 drain_right.n30 1.93989
R1223 drain_right.n110 drain_right.n14 1.93989
R1224 drain_right.n123 drain_right.n8 1.93989
R1225 drain_right.n265 drain_right.n150 1.93989
R1226 drain_right.n252 drain_right.n156 1.93989
R1227 drain_right.n217 drain_right.n173 1.93989
R1228 drain_right.n204 drain_right.n180 1.93989
R1229 drain_right.n65 drain_right.n63 1.16414
R1230 drain_right.n73 drain_right.n32 1.16414
R1231 drain_right.n111 drain_right.n12 1.16414
R1232 drain_right.n120 drain_right.n119 1.16414
R1233 drain_right.n262 drain_right.n261 1.16414
R1234 drain_right.n253 drain_right.n154 1.16414
R1235 drain_right.n216 drain_right.n175 1.16414
R1236 drain_right.n208 drain_right.n207 1.16414
R1237 drain_right.n139 drain_right.t2 0.7925
R1238 drain_right.n139 drain_right.t0 0.7925
R1239 drain_right.n141 drain_right.t3 0.7925
R1240 drain_right.n141 drain_right.t1 0.7925
R1241 drain_right.n64 drain_right.n34 0.388379
R1242 drain_right.n70 drain_right.n69 0.388379
R1243 drain_right.n115 drain_right.n114 0.388379
R1244 drain_right.n116 drain_right.n10 0.388379
R1245 drain_right.n258 drain_right.n152 0.388379
R1246 drain_right.n257 drain_right.n256 0.388379
R1247 drain_right.n213 drain_right.n212 0.388379
R1248 drain_right.n179 drain_right.n177 0.388379
R1249 drain_right.n46 drain_right.n41 0.155672
R1250 drain_right.n53 drain_right.n41 0.155672
R1251 drain_right.n54 drain_right.n53 0.155672
R1252 drain_right.n54 drain_right.n37 0.155672
R1253 drain_right.n61 drain_right.n37 0.155672
R1254 drain_right.n62 drain_right.n61 0.155672
R1255 drain_right.n62 drain_right.n33 0.155672
R1256 drain_right.n71 drain_right.n33 0.155672
R1257 drain_right.n72 drain_right.n71 0.155672
R1258 drain_right.n72 drain_right.n29 0.155672
R1259 drain_right.n79 drain_right.n29 0.155672
R1260 drain_right.n80 drain_right.n79 0.155672
R1261 drain_right.n80 drain_right.n25 0.155672
R1262 drain_right.n87 drain_right.n25 0.155672
R1263 drain_right.n88 drain_right.n87 0.155672
R1264 drain_right.n88 drain_right.n21 0.155672
R1265 drain_right.n95 drain_right.n21 0.155672
R1266 drain_right.n96 drain_right.n95 0.155672
R1267 drain_right.n96 drain_right.n17 0.155672
R1268 drain_right.n103 drain_right.n17 0.155672
R1269 drain_right.n104 drain_right.n103 0.155672
R1270 drain_right.n104 drain_right.n13 0.155672
R1271 drain_right.n112 drain_right.n13 0.155672
R1272 drain_right.n113 drain_right.n112 0.155672
R1273 drain_right.n113 drain_right.n9 0.155672
R1274 drain_right.n121 drain_right.n9 0.155672
R1275 drain_right.n122 drain_right.n121 0.155672
R1276 drain_right.n122 drain_right.n5 0.155672
R1277 drain_right.n129 drain_right.n5 0.155672
R1278 drain_right.n130 drain_right.n129 0.155672
R1279 drain_right.n130 drain_right.n1 0.155672
R1280 drain_right.n137 drain_right.n1 0.155672
R1281 drain_right.n279 drain_right.n143 0.155672
R1282 drain_right.n272 drain_right.n143 0.155672
R1283 drain_right.n272 drain_right.n271 0.155672
R1284 drain_right.n271 drain_right.n147 0.155672
R1285 drain_right.n264 drain_right.n147 0.155672
R1286 drain_right.n264 drain_right.n263 0.155672
R1287 drain_right.n263 drain_right.n151 0.155672
R1288 drain_right.n255 drain_right.n151 0.155672
R1289 drain_right.n255 drain_right.n254 0.155672
R1290 drain_right.n254 drain_right.n155 0.155672
R1291 drain_right.n247 drain_right.n155 0.155672
R1292 drain_right.n247 drain_right.n246 0.155672
R1293 drain_right.n246 drain_right.n160 0.155672
R1294 drain_right.n239 drain_right.n160 0.155672
R1295 drain_right.n239 drain_right.n238 0.155672
R1296 drain_right.n238 drain_right.n164 0.155672
R1297 drain_right.n231 drain_right.n164 0.155672
R1298 drain_right.n231 drain_right.n230 0.155672
R1299 drain_right.n230 drain_right.n168 0.155672
R1300 drain_right.n223 drain_right.n168 0.155672
R1301 drain_right.n223 drain_right.n222 0.155672
R1302 drain_right.n222 drain_right.n172 0.155672
R1303 drain_right.n215 drain_right.n172 0.155672
R1304 drain_right.n215 drain_right.n214 0.155672
R1305 drain_right.n214 drain_right.n176 0.155672
R1306 drain_right.n206 drain_right.n176 0.155672
R1307 drain_right.n206 drain_right.n205 0.155672
R1308 drain_right.n205 drain_right.n181 0.155672
R1309 drain_right.n198 drain_right.n181 0.155672
R1310 drain_right.n198 drain_right.n197 0.155672
R1311 drain_right.n197 drain_right.n185 0.155672
R1312 drain_right.n190 drain_right.n185 0.155672
R1313 plus.n1 plus.t4 825.716
R1314 plus.n7 plus.t5 825.716
R1315 plus.n4 plus.t1 802.23
R1316 plus.n2 plus.t3 802.23
R1317 plus.n10 plus.t2 802.23
R1318 plus.n8 plus.t0 802.23
R1319 plus.n3 plus.n0 161.3
R1320 plus.n5 plus.n4 161.3
R1321 plus.n9 plus.n6 161.3
R1322 plus.n11 plus.n10 161.3
R1323 plus.n7 plus.n6 44.8973
R1324 plus.n1 plus.n0 44.8973
R1325 plus plus.n11 34.285
R1326 plus.n4 plus.n3 33.5944
R1327 plus.n10 plus.n9 33.5944
R1328 plus.n8 plus.n7 18.1882
R1329 plus.n2 plus.n1 18.1882
R1330 plus plus.n5 17.2903
R1331 plus.n3 plus.n2 14.6066
R1332 plus.n9 plus.n8 14.6066
R1333 plus.n5 plus.n0 0.189894
R1334 plus.n11 plus.n6 0.189894
R1335 drain_left.n134 drain_left.n0 289.615
R1336 drain_left.n275 drain_left.n141 289.615
R1337 drain_left.n44 drain_left.n43 185
R1338 drain_left.n49 drain_left.n48 185
R1339 drain_left.n51 drain_left.n50 185
R1340 drain_left.n40 drain_left.n39 185
R1341 drain_left.n57 drain_left.n56 185
R1342 drain_left.n59 drain_left.n58 185
R1343 drain_left.n36 drain_left.n35 185
R1344 drain_left.n66 drain_left.n65 185
R1345 drain_left.n67 drain_left.n34 185
R1346 drain_left.n69 drain_left.n68 185
R1347 drain_left.n32 drain_left.n31 185
R1348 drain_left.n75 drain_left.n74 185
R1349 drain_left.n77 drain_left.n76 185
R1350 drain_left.n28 drain_left.n27 185
R1351 drain_left.n83 drain_left.n82 185
R1352 drain_left.n85 drain_left.n84 185
R1353 drain_left.n24 drain_left.n23 185
R1354 drain_left.n91 drain_left.n90 185
R1355 drain_left.n93 drain_left.n92 185
R1356 drain_left.n20 drain_left.n19 185
R1357 drain_left.n99 drain_left.n98 185
R1358 drain_left.n101 drain_left.n100 185
R1359 drain_left.n16 drain_left.n15 185
R1360 drain_left.n107 drain_left.n106 185
R1361 drain_left.n110 drain_left.n109 185
R1362 drain_left.n108 drain_left.n12 185
R1363 drain_left.n115 drain_left.n11 185
R1364 drain_left.n117 drain_left.n116 185
R1365 drain_left.n119 drain_left.n118 185
R1366 drain_left.n8 drain_left.n7 185
R1367 drain_left.n125 drain_left.n124 185
R1368 drain_left.n127 drain_left.n126 185
R1369 drain_left.n4 drain_left.n3 185
R1370 drain_left.n133 drain_left.n132 185
R1371 drain_left.n135 drain_left.n134 185
R1372 drain_left.n276 drain_left.n275 185
R1373 drain_left.n274 drain_left.n273 185
R1374 drain_left.n145 drain_left.n144 185
R1375 drain_left.n268 drain_left.n267 185
R1376 drain_left.n266 drain_left.n265 185
R1377 drain_left.n149 drain_left.n148 185
R1378 drain_left.n260 drain_left.n259 185
R1379 drain_left.n258 drain_left.n257 185
R1380 drain_left.n256 drain_left.n152 185
R1381 drain_left.n156 drain_left.n153 185
R1382 drain_left.n251 drain_left.n250 185
R1383 drain_left.n249 drain_left.n248 185
R1384 drain_left.n158 drain_left.n157 185
R1385 drain_left.n243 drain_left.n242 185
R1386 drain_left.n241 drain_left.n240 185
R1387 drain_left.n162 drain_left.n161 185
R1388 drain_left.n235 drain_left.n234 185
R1389 drain_left.n233 drain_left.n232 185
R1390 drain_left.n166 drain_left.n165 185
R1391 drain_left.n227 drain_left.n226 185
R1392 drain_left.n225 drain_left.n224 185
R1393 drain_left.n170 drain_left.n169 185
R1394 drain_left.n219 drain_left.n218 185
R1395 drain_left.n217 drain_left.n216 185
R1396 drain_left.n174 drain_left.n173 185
R1397 drain_left.n211 drain_left.n210 185
R1398 drain_left.n209 drain_left.n176 185
R1399 drain_left.n208 drain_left.n207 185
R1400 drain_left.n179 drain_left.n177 185
R1401 drain_left.n202 drain_left.n201 185
R1402 drain_left.n200 drain_left.n199 185
R1403 drain_left.n183 drain_left.n182 185
R1404 drain_left.n194 drain_left.n193 185
R1405 drain_left.n192 drain_left.n191 185
R1406 drain_left.n187 drain_left.n186 185
R1407 drain_left.n45 drain_left.t3 149.524
R1408 drain_left.n188 drain_left.t1 149.524
R1409 drain_left.n49 drain_left.n43 104.615
R1410 drain_left.n50 drain_left.n49 104.615
R1411 drain_left.n50 drain_left.n39 104.615
R1412 drain_left.n57 drain_left.n39 104.615
R1413 drain_left.n58 drain_left.n57 104.615
R1414 drain_left.n58 drain_left.n35 104.615
R1415 drain_left.n66 drain_left.n35 104.615
R1416 drain_left.n67 drain_left.n66 104.615
R1417 drain_left.n68 drain_left.n67 104.615
R1418 drain_left.n68 drain_left.n31 104.615
R1419 drain_left.n75 drain_left.n31 104.615
R1420 drain_left.n76 drain_left.n75 104.615
R1421 drain_left.n76 drain_left.n27 104.615
R1422 drain_left.n83 drain_left.n27 104.615
R1423 drain_left.n84 drain_left.n83 104.615
R1424 drain_left.n84 drain_left.n23 104.615
R1425 drain_left.n91 drain_left.n23 104.615
R1426 drain_left.n92 drain_left.n91 104.615
R1427 drain_left.n92 drain_left.n19 104.615
R1428 drain_left.n99 drain_left.n19 104.615
R1429 drain_left.n100 drain_left.n99 104.615
R1430 drain_left.n100 drain_left.n15 104.615
R1431 drain_left.n107 drain_left.n15 104.615
R1432 drain_left.n109 drain_left.n107 104.615
R1433 drain_left.n109 drain_left.n108 104.615
R1434 drain_left.n108 drain_left.n11 104.615
R1435 drain_left.n117 drain_left.n11 104.615
R1436 drain_left.n118 drain_left.n117 104.615
R1437 drain_left.n118 drain_left.n7 104.615
R1438 drain_left.n125 drain_left.n7 104.615
R1439 drain_left.n126 drain_left.n125 104.615
R1440 drain_left.n126 drain_left.n3 104.615
R1441 drain_left.n133 drain_left.n3 104.615
R1442 drain_left.n134 drain_left.n133 104.615
R1443 drain_left.n275 drain_left.n274 104.615
R1444 drain_left.n274 drain_left.n144 104.615
R1445 drain_left.n267 drain_left.n144 104.615
R1446 drain_left.n267 drain_left.n266 104.615
R1447 drain_left.n266 drain_left.n148 104.615
R1448 drain_left.n259 drain_left.n148 104.615
R1449 drain_left.n259 drain_left.n258 104.615
R1450 drain_left.n258 drain_left.n152 104.615
R1451 drain_left.n156 drain_left.n152 104.615
R1452 drain_left.n250 drain_left.n156 104.615
R1453 drain_left.n250 drain_left.n249 104.615
R1454 drain_left.n249 drain_left.n157 104.615
R1455 drain_left.n242 drain_left.n157 104.615
R1456 drain_left.n242 drain_left.n241 104.615
R1457 drain_left.n241 drain_left.n161 104.615
R1458 drain_left.n234 drain_left.n161 104.615
R1459 drain_left.n234 drain_left.n233 104.615
R1460 drain_left.n233 drain_left.n165 104.615
R1461 drain_left.n226 drain_left.n165 104.615
R1462 drain_left.n226 drain_left.n225 104.615
R1463 drain_left.n225 drain_left.n169 104.615
R1464 drain_left.n218 drain_left.n169 104.615
R1465 drain_left.n218 drain_left.n217 104.615
R1466 drain_left.n217 drain_left.n173 104.615
R1467 drain_left.n210 drain_left.n173 104.615
R1468 drain_left.n210 drain_left.n209 104.615
R1469 drain_left.n209 drain_left.n208 104.615
R1470 drain_left.n208 drain_left.n177 104.615
R1471 drain_left.n201 drain_left.n177 104.615
R1472 drain_left.n201 drain_left.n200 104.615
R1473 drain_left.n200 drain_left.n182 104.615
R1474 drain_left.n193 drain_left.n182 104.615
R1475 drain_left.n193 drain_left.n192 104.615
R1476 drain_left.n192 drain_left.n186 104.615
R1477 drain_left.n140 drain_left.n139 58.9036
R1478 drain_left.n281 drain_left.n280 58.7153
R1479 drain_left.t3 drain_left.n43 52.3082
R1480 drain_left.t1 drain_left.n186 52.3082
R1481 drain_left.n281 drain_left.n279 48.2868
R1482 drain_left.n140 drain_left.n138 47.9879
R1483 drain_left drain_left.n140 39.8944
R1484 drain_left.n69 drain_left.n34 13.1884
R1485 drain_left.n116 drain_left.n115 13.1884
R1486 drain_left.n257 drain_left.n256 13.1884
R1487 drain_left.n211 drain_left.n176 13.1884
R1488 drain_left.n65 drain_left.n64 12.8005
R1489 drain_left.n70 drain_left.n32 12.8005
R1490 drain_left.n114 drain_left.n12 12.8005
R1491 drain_left.n119 drain_left.n10 12.8005
R1492 drain_left.n260 drain_left.n151 12.8005
R1493 drain_left.n255 drain_left.n153 12.8005
R1494 drain_left.n212 drain_left.n174 12.8005
R1495 drain_left.n207 drain_left.n178 12.8005
R1496 drain_left.n63 drain_left.n36 12.0247
R1497 drain_left.n74 drain_left.n73 12.0247
R1498 drain_left.n111 drain_left.n110 12.0247
R1499 drain_left.n120 drain_left.n8 12.0247
R1500 drain_left.n261 drain_left.n149 12.0247
R1501 drain_left.n252 drain_left.n251 12.0247
R1502 drain_left.n216 drain_left.n215 12.0247
R1503 drain_left.n206 drain_left.n179 12.0247
R1504 drain_left.n60 drain_left.n59 11.249
R1505 drain_left.n77 drain_left.n30 11.249
R1506 drain_left.n106 drain_left.n14 11.249
R1507 drain_left.n124 drain_left.n123 11.249
R1508 drain_left.n265 drain_left.n264 11.249
R1509 drain_left.n248 drain_left.n155 11.249
R1510 drain_left.n219 drain_left.n172 11.249
R1511 drain_left.n203 drain_left.n202 11.249
R1512 drain_left.n56 drain_left.n38 10.4732
R1513 drain_left.n78 drain_left.n28 10.4732
R1514 drain_left.n105 drain_left.n16 10.4732
R1515 drain_left.n127 drain_left.n6 10.4732
R1516 drain_left.n268 drain_left.n147 10.4732
R1517 drain_left.n247 drain_left.n158 10.4732
R1518 drain_left.n220 drain_left.n170 10.4732
R1519 drain_left.n199 drain_left.n181 10.4732
R1520 drain_left.n45 drain_left.n44 10.2747
R1521 drain_left.n188 drain_left.n187 10.2747
R1522 drain_left.n55 drain_left.n40 9.69747
R1523 drain_left.n82 drain_left.n81 9.69747
R1524 drain_left.n102 drain_left.n101 9.69747
R1525 drain_left.n128 drain_left.n4 9.69747
R1526 drain_left.n269 drain_left.n145 9.69747
R1527 drain_left.n244 drain_left.n243 9.69747
R1528 drain_left.n224 drain_left.n223 9.69747
R1529 drain_left.n198 drain_left.n183 9.69747
R1530 drain_left.n138 drain_left.n137 9.45567
R1531 drain_left.n279 drain_left.n278 9.45567
R1532 drain_left.n2 drain_left.n1 9.3005
R1533 drain_left.n131 drain_left.n130 9.3005
R1534 drain_left.n129 drain_left.n128 9.3005
R1535 drain_left.n6 drain_left.n5 9.3005
R1536 drain_left.n123 drain_left.n122 9.3005
R1537 drain_left.n121 drain_left.n120 9.3005
R1538 drain_left.n10 drain_left.n9 9.3005
R1539 drain_left.n89 drain_left.n88 9.3005
R1540 drain_left.n87 drain_left.n86 9.3005
R1541 drain_left.n26 drain_left.n25 9.3005
R1542 drain_left.n81 drain_left.n80 9.3005
R1543 drain_left.n79 drain_left.n78 9.3005
R1544 drain_left.n30 drain_left.n29 9.3005
R1545 drain_left.n73 drain_left.n72 9.3005
R1546 drain_left.n71 drain_left.n70 9.3005
R1547 drain_left.n47 drain_left.n46 9.3005
R1548 drain_left.n42 drain_left.n41 9.3005
R1549 drain_left.n53 drain_left.n52 9.3005
R1550 drain_left.n55 drain_left.n54 9.3005
R1551 drain_left.n38 drain_left.n37 9.3005
R1552 drain_left.n61 drain_left.n60 9.3005
R1553 drain_left.n63 drain_left.n62 9.3005
R1554 drain_left.n64 drain_left.n33 9.3005
R1555 drain_left.n22 drain_left.n21 9.3005
R1556 drain_left.n95 drain_left.n94 9.3005
R1557 drain_left.n97 drain_left.n96 9.3005
R1558 drain_left.n18 drain_left.n17 9.3005
R1559 drain_left.n103 drain_left.n102 9.3005
R1560 drain_left.n105 drain_left.n104 9.3005
R1561 drain_left.n14 drain_left.n13 9.3005
R1562 drain_left.n112 drain_left.n111 9.3005
R1563 drain_left.n114 drain_left.n113 9.3005
R1564 drain_left.n137 drain_left.n136 9.3005
R1565 drain_left.n190 drain_left.n189 9.3005
R1566 drain_left.n185 drain_left.n184 9.3005
R1567 drain_left.n196 drain_left.n195 9.3005
R1568 drain_left.n198 drain_left.n197 9.3005
R1569 drain_left.n181 drain_left.n180 9.3005
R1570 drain_left.n204 drain_left.n203 9.3005
R1571 drain_left.n206 drain_left.n205 9.3005
R1572 drain_left.n178 drain_left.n175 9.3005
R1573 drain_left.n237 drain_left.n236 9.3005
R1574 drain_left.n239 drain_left.n238 9.3005
R1575 drain_left.n160 drain_left.n159 9.3005
R1576 drain_left.n245 drain_left.n244 9.3005
R1577 drain_left.n247 drain_left.n246 9.3005
R1578 drain_left.n155 drain_left.n154 9.3005
R1579 drain_left.n253 drain_left.n252 9.3005
R1580 drain_left.n255 drain_left.n254 9.3005
R1581 drain_left.n278 drain_left.n277 9.3005
R1582 drain_left.n143 drain_left.n142 9.3005
R1583 drain_left.n272 drain_left.n271 9.3005
R1584 drain_left.n270 drain_left.n269 9.3005
R1585 drain_left.n147 drain_left.n146 9.3005
R1586 drain_left.n264 drain_left.n263 9.3005
R1587 drain_left.n262 drain_left.n261 9.3005
R1588 drain_left.n151 drain_left.n150 9.3005
R1589 drain_left.n164 drain_left.n163 9.3005
R1590 drain_left.n231 drain_left.n230 9.3005
R1591 drain_left.n229 drain_left.n228 9.3005
R1592 drain_left.n168 drain_left.n167 9.3005
R1593 drain_left.n223 drain_left.n222 9.3005
R1594 drain_left.n221 drain_left.n220 9.3005
R1595 drain_left.n172 drain_left.n171 9.3005
R1596 drain_left.n215 drain_left.n214 9.3005
R1597 drain_left.n213 drain_left.n212 9.3005
R1598 drain_left.n52 drain_left.n51 8.92171
R1599 drain_left.n85 drain_left.n26 8.92171
R1600 drain_left.n98 drain_left.n18 8.92171
R1601 drain_left.n132 drain_left.n131 8.92171
R1602 drain_left.n273 drain_left.n272 8.92171
R1603 drain_left.n240 drain_left.n160 8.92171
R1604 drain_left.n227 drain_left.n168 8.92171
R1605 drain_left.n195 drain_left.n194 8.92171
R1606 drain_left.n48 drain_left.n42 8.14595
R1607 drain_left.n86 drain_left.n24 8.14595
R1608 drain_left.n97 drain_left.n20 8.14595
R1609 drain_left.n135 drain_left.n2 8.14595
R1610 drain_left.n276 drain_left.n143 8.14595
R1611 drain_left.n239 drain_left.n162 8.14595
R1612 drain_left.n228 drain_left.n166 8.14595
R1613 drain_left.n191 drain_left.n185 8.14595
R1614 drain_left.n47 drain_left.n44 7.3702
R1615 drain_left.n90 drain_left.n89 7.3702
R1616 drain_left.n94 drain_left.n93 7.3702
R1617 drain_left.n136 drain_left.n0 7.3702
R1618 drain_left.n277 drain_left.n141 7.3702
R1619 drain_left.n236 drain_left.n235 7.3702
R1620 drain_left.n232 drain_left.n231 7.3702
R1621 drain_left.n190 drain_left.n187 7.3702
R1622 drain_left drain_left.n281 6.62735
R1623 drain_left.n90 drain_left.n22 6.59444
R1624 drain_left.n93 drain_left.n22 6.59444
R1625 drain_left.n138 drain_left.n0 6.59444
R1626 drain_left.n279 drain_left.n141 6.59444
R1627 drain_left.n235 drain_left.n164 6.59444
R1628 drain_left.n232 drain_left.n164 6.59444
R1629 drain_left.n48 drain_left.n47 5.81868
R1630 drain_left.n89 drain_left.n24 5.81868
R1631 drain_left.n94 drain_left.n20 5.81868
R1632 drain_left.n136 drain_left.n135 5.81868
R1633 drain_left.n277 drain_left.n276 5.81868
R1634 drain_left.n236 drain_left.n162 5.81868
R1635 drain_left.n231 drain_left.n166 5.81868
R1636 drain_left.n191 drain_left.n190 5.81868
R1637 drain_left.n51 drain_left.n42 5.04292
R1638 drain_left.n86 drain_left.n85 5.04292
R1639 drain_left.n98 drain_left.n97 5.04292
R1640 drain_left.n132 drain_left.n2 5.04292
R1641 drain_left.n273 drain_left.n143 5.04292
R1642 drain_left.n240 drain_left.n239 5.04292
R1643 drain_left.n228 drain_left.n227 5.04292
R1644 drain_left.n194 drain_left.n185 5.04292
R1645 drain_left.n52 drain_left.n40 4.26717
R1646 drain_left.n82 drain_left.n26 4.26717
R1647 drain_left.n101 drain_left.n18 4.26717
R1648 drain_left.n131 drain_left.n4 4.26717
R1649 drain_left.n272 drain_left.n145 4.26717
R1650 drain_left.n243 drain_left.n160 4.26717
R1651 drain_left.n224 drain_left.n168 4.26717
R1652 drain_left.n195 drain_left.n183 4.26717
R1653 drain_left.n56 drain_left.n55 3.49141
R1654 drain_left.n81 drain_left.n28 3.49141
R1655 drain_left.n102 drain_left.n16 3.49141
R1656 drain_left.n128 drain_left.n127 3.49141
R1657 drain_left.n269 drain_left.n268 3.49141
R1658 drain_left.n244 drain_left.n158 3.49141
R1659 drain_left.n223 drain_left.n170 3.49141
R1660 drain_left.n199 drain_left.n198 3.49141
R1661 drain_left.n189 drain_left.n188 2.84303
R1662 drain_left.n46 drain_left.n45 2.84303
R1663 drain_left.n59 drain_left.n38 2.71565
R1664 drain_left.n78 drain_left.n77 2.71565
R1665 drain_left.n106 drain_left.n105 2.71565
R1666 drain_left.n124 drain_left.n6 2.71565
R1667 drain_left.n265 drain_left.n147 2.71565
R1668 drain_left.n248 drain_left.n247 2.71565
R1669 drain_left.n220 drain_left.n219 2.71565
R1670 drain_left.n202 drain_left.n181 2.71565
R1671 drain_left.n60 drain_left.n36 1.93989
R1672 drain_left.n74 drain_left.n30 1.93989
R1673 drain_left.n110 drain_left.n14 1.93989
R1674 drain_left.n123 drain_left.n8 1.93989
R1675 drain_left.n264 drain_left.n149 1.93989
R1676 drain_left.n251 drain_left.n155 1.93989
R1677 drain_left.n216 drain_left.n172 1.93989
R1678 drain_left.n203 drain_left.n179 1.93989
R1679 drain_left.n65 drain_left.n63 1.16414
R1680 drain_left.n73 drain_left.n32 1.16414
R1681 drain_left.n111 drain_left.n12 1.16414
R1682 drain_left.n120 drain_left.n119 1.16414
R1683 drain_left.n261 drain_left.n260 1.16414
R1684 drain_left.n252 drain_left.n153 1.16414
R1685 drain_left.n215 drain_left.n174 1.16414
R1686 drain_left.n207 drain_left.n206 1.16414
R1687 drain_left.n139 drain_left.t5 0.7925
R1688 drain_left.n139 drain_left.t0 0.7925
R1689 drain_left.n280 drain_left.t2 0.7925
R1690 drain_left.n280 drain_left.t4 0.7925
R1691 drain_left.n64 drain_left.n34 0.388379
R1692 drain_left.n70 drain_left.n69 0.388379
R1693 drain_left.n115 drain_left.n114 0.388379
R1694 drain_left.n116 drain_left.n10 0.388379
R1695 drain_left.n257 drain_left.n151 0.388379
R1696 drain_left.n256 drain_left.n255 0.388379
R1697 drain_left.n212 drain_left.n211 0.388379
R1698 drain_left.n178 drain_left.n176 0.388379
R1699 drain_left.n46 drain_left.n41 0.155672
R1700 drain_left.n53 drain_left.n41 0.155672
R1701 drain_left.n54 drain_left.n53 0.155672
R1702 drain_left.n54 drain_left.n37 0.155672
R1703 drain_left.n61 drain_left.n37 0.155672
R1704 drain_left.n62 drain_left.n61 0.155672
R1705 drain_left.n62 drain_left.n33 0.155672
R1706 drain_left.n71 drain_left.n33 0.155672
R1707 drain_left.n72 drain_left.n71 0.155672
R1708 drain_left.n72 drain_left.n29 0.155672
R1709 drain_left.n79 drain_left.n29 0.155672
R1710 drain_left.n80 drain_left.n79 0.155672
R1711 drain_left.n80 drain_left.n25 0.155672
R1712 drain_left.n87 drain_left.n25 0.155672
R1713 drain_left.n88 drain_left.n87 0.155672
R1714 drain_left.n88 drain_left.n21 0.155672
R1715 drain_left.n95 drain_left.n21 0.155672
R1716 drain_left.n96 drain_left.n95 0.155672
R1717 drain_left.n96 drain_left.n17 0.155672
R1718 drain_left.n103 drain_left.n17 0.155672
R1719 drain_left.n104 drain_left.n103 0.155672
R1720 drain_left.n104 drain_left.n13 0.155672
R1721 drain_left.n112 drain_left.n13 0.155672
R1722 drain_left.n113 drain_left.n112 0.155672
R1723 drain_left.n113 drain_left.n9 0.155672
R1724 drain_left.n121 drain_left.n9 0.155672
R1725 drain_left.n122 drain_left.n121 0.155672
R1726 drain_left.n122 drain_left.n5 0.155672
R1727 drain_left.n129 drain_left.n5 0.155672
R1728 drain_left.n130 drain_left.n129 0.155672
R1729 drain_left.n130 drain_left.n1 0.155672
R1730 drain_left.n137 drain_left.n1 0.155672
R1731 drain_left.n278 drain_left.n142 0.155672
R1732 drain_left.n271 drain_left.n142 0.155672
R1733 drain_left.n271 drain_left.n270 0.155672
R1734 drain_left.n270 drain_left.n146 0.155672
R1735 drain_left.n263 drain_left.n146 0.155672
R1736 drain_left.n263 drain_left.n262 0.155672
R1737 drain_left.n262 drain_left.n150 0.155672
R1738 drain_left.n254 drain_left.n150 0.155672
R1739 drain_left.n254 drain_left.n253 0.155672
R1740 drain_left.n253 drain_left.n154 0.155672
R1741 drain_left.n246 drain_left.n154 0.155672
R1742 drain_left.n246 drain_left.n245 0.155672
R1743 drain_left.n245 drain_left.n159 0.155672
R1744 drain_left.n238 drain_left.n159 0.155672
R1745 drain_left.n238 drain_left.n237 0.155672
R1746 drain_left.n237 drain_left.n163 0.155672
R1747 drain_left.n230 drain_left.n163 0.155672
R1748 drain_left.n230 drain_left.n229 0.155672
R1749 drain_left.n229 drain_left.n167 0.155672
R1750 drain_left.n222 drain_left.n167 0.155672
R1751 drain_left.n222 drain_left.n221 0.155672
R1752 drain_left.n221 drain_left.n171 0.155672
R1753 drain_left.n214 drain_left.n171 0.155672
R1754 drain_left.n214 drain_left.n213 0.155672
R1755 drain_left.n213 drain_left.n175 0.155672
R1756 drain_left.n205 drain_left.n175 0.155672
R1757 drain_left.n205 drain_left.n204 0.155672
R1758 drain_left.n204 drain_left.n180 0.155672
R1759 drain_left.n197 drain_left.n180 0.155672
R1760 drain_left.n197 drain_left.n196 0.155672
R1761 drain_left.n196 drain_left.n184 0.155672
R1762 drain_left.n189 drain_left.n184 0.155672
C0 minus plus 7.56129f
C1 source minus 8.47654f
C2 drain_left plus 9.44831f
C3 drain_right minus 9.29725f
C4 drain_left source 17.870802f
C5 drain_right drain_left 0.749358f
C6 source plus 8.49156f
C7 drain_right plus 0.313788f
C8 drain_left minus 0.171398f
C9 drain_right source 17.8571f
C10 drain_right a_n1620_n5888# 9.83215f
C11 drain_left a_n1620_n5888# 10.074979f
C12 source a_n1620_n5888# 11.374064f
C13 minus a_n1620_n5888# 7.053319f
C14 plus a_n1620_n5888# 9.38962f
C15 drain_left.n0 a_n1620_n5888# 0.031335f
C16 drain_left.n1 a_n1620_n5888# 0.02273f
C17 drain_left.n2 a_n1620_n5888# 0.012214f
C18 drain_left.n3 a_n1620_n5888# 0.028869f
C19 drain_left.n4 a_n1620_n5888# 0.012932f
C20 drain_left.n5 a_n1620_n5888# 0.02273f
C21 drain_left.n6 a_n1620_n5888# 0.012214f
C22 drain_left.n7 a_n1620_n5888# 0.028869f
C23 drain_left.n8 a_n1620_n5888# 0.012932f
C24 drain_left.n9 a_n1620_n5888# 0.02273f
C25 drain_left.n10 a_n1620_n5888# 0.012214f
C26 drain_left.n11 a_n1620_n5888# 0.028869f
C27 drain_left.n12 a_n1620_n5888# 0.012932f
C28 drain_left.n13 a_n1620_n5888# 0.02273f
C29 drain_left.n14 a_n1620_n5888# 0.012214f
C30 drain_left.n15 a_n1620_n5888# 0.028869f
C31 drain_left.n16 a_n1620_n5888# 0.012932f
C32 drain_left.n17 a_n1620_n5888# 0.02273f
C33 drain_left.n18 a_n1620_n5888# 0.012214f
C34 drain_left.n19 a_n1620_n5888# 0.028869f
C35 drain_left.n20 a_n1620_n5888# 0.012932f
C36 drain_left.n21 a_n1620_n5888# 0.02273f
C37 drain_left.n22 a_n1620_n5888# 0.012214f
C38 drain_left.n23 a_n1620_n5888# 0.028869f
C39 drain_left.n24 a_n1620_n5888# 0.012932f
C40 drain_left.n25 a_n1620_n5888# 0.02273f
C41 drain_left.n26 a_n1620_n5888# 0.012214f
C42 drain_left.n27 a_n1620_n5888# 0.028869f
C43 drain_left.n28 a_n1620_n5888# 0.012932f
C44 drain_left.n29 a_n1620_n5888# 0.02273f
C45 drain_left.n30 a_n1620_n5888# 0.012214f
C46 drain_left.n31 a_n1620_n5888# 0.028869f
C47 drain_left.n32 a_n1620_n5888# 0.012932f
C48 drain_left.n33 a_n1620_n5888# 0.02273f
C49 drain_left.n34 a_n1620_n5888# 0.012573f
C50 drain_left.n35 a_n1620_n5888# 0.028869f
C51 drain_left.n36 a_n1620_n5888# 0.012932f
C52 drain_left.n37 a_n1620_n5888# 0.02273f
C53 drain_left.n38 a_n1620_n5888# 0.012214f
C54 drain_left.n39 a_n1620_n5888# 0.028869f
C55 drain_left.n40 a_n1620_n5888# 0.012932f
C56 drain_left.n41 a_n1620_n5888# 0.02273f
C57 drain_left.n42 a_n1620_n5888# 0.012214f
C58 drain_left.n43 a_n1620_n5888# 0.021652f
C59 drain_left.n44 a_n1620_n5888# 0.020408f
C60 drain_left.t3 a_n1620_n5888# 0.05035f
C61 drain_left.n45 a_n1620_n5888# 0.27732f
C62 drain_left.n46 a_n1620_n5888# 2.46095f
C63 drain_left.n47 a_n1620_n5888# 0.012214f
C64 drain_left.n48 a_n1620_n5888# 0.012932f
C65 drain_left.n49 a_n1620_n5888# 0.028869f
C66 drain_left.n50 a_n1620_n5888# 0.028869f
C67 drain_left.n51 a_n1620_n5888# 0.012932f
C68 drain_left.n52 a_n1620_n5888# 0.012214f
C69 drain_left.n53 a_n1620_n5888# 0.02273f
C70 drain_left.n54 a_n1620_n5888# 0.02273f
C71 drain_left.n55 a_n1620_n5888# 0.012214f
C72 drain_left.n56 a_n1620_n5888# 0.012932f
C73 drain_left.n57 a_n1620_n5888# 0.028869f
C74 drain_left.n58 a_n1620_n5888# 0.028869f
C75 drain_left.n59 a_n1620_n5888# 0.012932f
C76 drain_left.n60 a_n1620_n5888# 0.012214f
C77 drain_left.n61 a_n1620_n5888# 0.02273f
C78 drain_left.n62 a_n1620_n5888# 0.02273f
C79 drain_left.n63 a_n1620_n5888# 0.012214f
C80 drain_left.n64 a_n1620_n5888# 0.012214f
C81 drain_left.n65 a_n1620_n5888# 0.012932f
C82 drain_left.n66 a_n1620_n5888# 0.028869f
C83 drain_left.n67 a_n1620_n5888# 0.028869f
C84 drain_left.n68 a_n1620_n5888# 0.028869f
C85 drain_left.n69 a_n1620_n5888# 0.012573f
C86 drain_left.n70 a_n1620_n5888# 0.012214f
C87 drain_left.n71 a_n1620_n5888# 0.02273f
C88 drain_left.n72 a_n1620_n5888# 0.02273f
C89 drain_left.n73 a_n1620_n5888# 0.012214f
C90 drain_left.n74 a_n1620_n5888# 0.012932f
C91 drain_left.n75 a_n1620_n5888# 0.028869f
C92 drain_left.n76 a_n1620_n5888# 0.028869f
C93 drain_left.n77 a_n1620_n5888# 0.012932f
C94 drain_left.n78 a_n1620_n5888# 0.012214f
C95 drain_left.n79 a_n1620_n5888# 0.02273f
C96 drain_left.n80 a_n1620_n5888# 0.02273f
C97 drain_left.n81 a_n1620_n5888# 0.012214f
C98 drain_left.n82 a_n1620_n5888# 0.012932f
C99 drain_left.n83 a_n1620_n5888# 0.028869f
C100 drain_left.n84 a_n1620_n5888# 0.028869f
C101 drain_left.n85 a_n1620_n5888# 0.012932f
C102 drain_left.n86 a_n1620_n5888# 0.012214f
C103 drain_left.n87 a_n1620_n5888# 0.02273f
C104 drain_left.n88 a_n1620_n5888# 0.02273f
C105 drain_left.n89 a_n1620_n5888# 0.012214f
C106 drain_left.n90 a_n1620_n5888# 0.012932f
C107 drain_left.n91 a_n1620_n5888# 0.028869f
C108 drain_left.n92 a_n1620_n5888# 0.028869f
C109 drain_left.n93 a_n1620_n5888# 0.012932f
C110 drain_left.n94 a_n1620_n5888# 0.012214f
C111 drain_left.n95 a_n1620_n5888# 0.02273f
C112 drain_left.n96 a_n1620_n5888# 0.02273f
C113 drain_left.n97 a_n1620_n5888# 0.012214f
C114 drain_left.n98 a_n1620_n5888# 0.012932f
C115 drain_left.n99 a_n1620_n5888# 0.028869f
C116 drain_left.n100 a_n1620_n5888# 0.028869f
C117 drain_left.n101 a_n1620_n5888# 0.012932f
C118 drain_left.n102 a_n1620_n5888# 0.012214f
C119 drain_left.n103 a_n1620_n5888# 0.02273f
C120 drain_left.n104 a_n1620_n5888# 0.02273f
C121 drain_left.n105 a_n1620_n5888# 0.012214f
C122 drain_left.n106 a_n1620_n5888# 0.012932f
C123 drain_left.n107 a_n1620_n5888# 0.028869f
C124 drain_left.n108 a_n1620_n5888# 0.028869f
C125 drain_left.n109 a_n1620_n5888# 0.028869f
C126 drain_left.n110 a_n1620_n5888# 0.012932f
C127 drain_left.n111 a_n1620_n5888# 0.012214f
C128 drain_left.n112 a_n1620_n5888# 0.02273f
C129 drain_left.n113 a_n1620_n5888# 0.02273f
C130 drain_left.n114 a_n1620_n5888# 0.012214f
C131 drain_left.n115 a_n1620_n5888# 0.012573f
C132 drain_left.n116 a_n1620_n5888# 0.012573f
C133 drain_left.n117 a_n1620_n5888# 0.028869f
C134 drain_left.n118 a_n1620_n5888# 0.028869f
C135 drain_left.n119 a_n1620_n5888# 0.012932f
C136 drain_left.n120 a_n1620_n5888# 0.012214f
C137 drain_left.n121 a_n1620_n5888# 0.02273f
C138 drain_left.n122 a_n1620_n5888# 0.02273f
C139 drain_left.n123 a_n1620_n5888# 0.012214f
C140 drain_left.n124 a_n1620_n5888# 0.012932f
C141 drain_left.n125 a_n1620_n5888# 0.028869f
C142 drain_left.n126 a_n1620_n5888# 0.028869f
C143 drain_left.n127 a_n1620_n5888# 0.012932f
C144 drain_left.n128 a_n1620_n5888# 0.012214f
C145 drain_left.n129 a_n1620_n5888# 0.02273f
C146 drain_left.n130 a_n1620_n5888# 0.02273f
C147 drain_left.n131 a_n1620_n5888# 0.012214f
C148 drain_left.n132 a_n1620_n5888# 0.012932f
C149 drain_left.n133 a_n1620_n5888# 0.028869f
C150 drain_left.n134 a_n1620_n5888# 0.061412f
C151 drain_left.n135 a_n1620_n5888# 0.012932f
C152 drain_left.n136 a_n1620_n5888# 0.012214f
C153 drain_left.n137 a_n1620_n5888# 0.050054f
C154 drain_left.n138 a_n1620_n5888# 0.051191f
C155 drain_left.t5 a_n1620_n5888# 0.449041f
C156 drain_left.t0 a_n1620_n5888# 0.449041f
C157 drain_left.n139 a_n1620_n5888# 4.13932f
C158 drain_left.n140 a_n1620_n5888# 2.21002f
C159 drain_left.n141 a_n1620_n5888# 0.031335f
C160 drain_left.n142 a_n1620_n5888# 0.02273f
C161 drain_left.n143 a_n1620_n5888# 0.012214f
C162 drain_left.n144 a_n1620_n5888# 0.028869f
C163 drain_left.n145 a_n1620_n5888# 0.012932f
C164 drain_left.n146 a_n1620_n5888# 0.02273f
C165 drain_left.n147 a_n1620_n5888# 0.012214f
C166 drain_left.n148 a_n1620_n5888# 0.028869f
C167 drain_left.n149 a_n1620_n5888# 0.012932f
C168 drain_left.n150 a_n1620_n5888# 0.02273f
C169 drain_left.n151 a_n1620_n5888# 0.012214f
C170 drain_left.n152 a_n1620_n5888# 0.028869f
C171 drain_left.n153 a_n1620_n5888# 0.012932f
C172 drain_left.n154 a_n1620_n5888# 0.02273f
C173 drain_left.n155 a_n1620_n5888# 0.012214f
C174 drain_left.n156 a_n1620_n5888# 0.028869f
C175 drain_left.n157 a_n1620_n5888# 0.028869f
C176 drain_left.n158 a_n1620_n5888# 0.012932f
C177 drain_left.n159 a_n1620_n5888# 0.02273f
C178 drain_left.n160 a_n1620_n5888# 0.012214f
C179 drain_left.n161 a_n1620_n5888# 0.028869f
C180 drain_left.n162 a_n1620_n5888# 0.012932f
C181 drain_left.n163 a_n1620_n5888# 0.02273f
C182 drain_left.n164 a_n1620_n5888# 0.012214f
C183 drain_left.n165 a_n1620_n5888# 0.028869f
C184 drain_left.n166 a_n1620_n5888# 0.012932f
C185 drain_left.n167 a_n1620_n5888# 0.02273f
C186 drain_left.n168 a_n1620_n5888# 0.012214f
C187 drain_left.n169 a_n1620_n5888# 0.028869f
C188 drain_left.n170 a_n1620_n5888# 0.012932f
C189 drain_left.n171 a_n1620_n5888# 0.02273f
C190 drain_left.n172 a_n1620_n5888# 0.012214f
C191 drain_left.n173 a_n1620_n5888# 0.028869f
C192 drain_left.n174 a_n1620_n5888# 0.012932f
C193 drain_left.n175 a_n1620_n5888# 0.02273f
C194 drain_left.n176 a_n1620_n5888# 0.012573f
C195 drain_left.n177 a_n1620_n5888# 0.028869f
C196 drain_left.n178 a_n1620_n5888# 0.012214f
C197 drain_left.n179 a_n1620_n5888# 0.012932f
C198 drain_left.n180 a_n1620_n5888# 0.02273f
C199 drain_left.n181 a_n1620_n5888# 0.012214f
C200 drain_left.n182 a_n1620_n5888# 0.028869f
C201 drain_left.n183 a_n1620_n5888# 0.012932f
C202 drain_left.n184 a_n1620_n5888# 0.02273f
C203 drain_left.n185 a_n1620_n5888# 0.012214f
C204 drain_left.n186 a_n1620_n5888# 0.021652f
C205 drain_left.n187 a_n1620_n5888# 0.020408f
C206 drain_left.t1 a_n1620_n5888# 0.05035f
C207 drain_left.n188 a_n1620_n5888# 0.27732f
C208 drain_left.n189 a_n1620_n5888# 2.46095f
C209 drain_left.n190 a_n1620_n5888# 0.012214f
C210 drain_left.n191 a_n1620_n5888# 0.012932f
C211 drain_left.n192 a_n1620_n5888# 0.028869f
C212 drain_left.n193 a_n1620_n5888# 0.028869f
C213 drain_left.n194 a_n1620_n5888# 0.012932f
C214 drain_left.n195 a_n1620_n5888# 0.012214f
C215 drain_left.n196 a_n1620_n5888# 0.02273f
C216 drain_left.n197 a_n1620_n5888# 0.02273f
C217 drain_left.n198 a_n1620_n5888# 0.012214f
C218 drain_left.n199 a_n1620_n5888# 0.012932f
C219 drain_left.n200 a_n1620_n5888# 0.028869f
C220 drain_left.n201 a_n1620_n5888# 0.028869f
C221 drain_left.n202 a_n1620_n5888# 0.012932f
C222 drain_left.n203 a_n1620_n5888# 0.012214f
C223 drain_left.n204 a_n1620_n5888# 0.02273f
C224 drain_left.n205 a_n1620_n5888# 0.02273f
C225 drain_left.n206 a_n1620_n5888# 0.012214f
C226 drain_left.n207 a_n1620_n5888# 0.012932f
C227 drain_left.n208 a_n1620_n5888# 0.028869f
C228 drain_left.n209 a_n1620_n5888# 0.028869f
C229 drain_left.n210 a_n1620_n5888# 0.028869f
C230 drain_left.n211 a_n1620_n5888# 0.012573f
C231 drain_left.n212 a_n1620_n5888# 0.012214f
C232 drain_left.n213 a_n1620_n5888# 0.02273f
C233 drain_left.n214 a_n1620_n5888# 0.02273f
C234 drain_left.n215 a_n1620_n5888# 0.012214f
C235 drain_left.n216 a_n1620_n5888# 0.012932f
C236 drain_left.n217 a_n1620_n5888# 0.028869f
C237 drain_left.n218 a_n1620_n5888# 0.028869f
C238 drain_left.n219 a_n1620_n5888# 0.012932f
C239 drain_left.n220 a_n1620_n5888# 0.012214f
C240 drain_left.n221 a_n1620_n5888# 0.02273f
C241 drain_left.n222 a_n1620_n5888# 0.02273f
C242 drain_left.n223 a_n1620_n5888# 0.012214f
C243 drain_left.n224 a_n1620_n5888# 0.012932f
C244 drain_left.n225 a_n1620_n5888# 0.028869f
C245 drain_left.n226 a_n1620_n5888# 0.028869f
C246 drain_left.n227 a_n1620_n5888# 0.012932f
C247 drain_left.n228 a_n1620_n5888# 0.012214f
C248 drain_left.n229 a_n1620_n5888# 0.02273f
C249 drain_left.n230 a_n1620_n5888# 0.02273f
C250 drain_left.n231 a_n1620_n5888# 0.012214f
C251 drain_left.n232 a_n1620_n5888# 0.012932f
C252 drain_left.n233 a_n1620_n5888# 0.028869f
C253 drain_left.n234 a_n1620_n5888# 0.028869f
C254 drain_left.n235 a_n1620_n5888# 0.012932f
C255 drain_left.n236 a_n1620_n5888# 0.012214f
C256 drain_left.n237 a_n1620_n5888# 0.02273f
C257 drain_left.n238 a_n1620_n5888# 0.02273f
C258 drain_left.n239 a_n1620_n5888# 0.012214f
C259 drain_left.n240 a_n1620_n5888# 0.012932f
C260 drain_left.n241 a_n1620_n5888# 0.028869f
C261 drain_left.n242 a_n1620_n5888# 0.028869f
C262 drain_left.n243 a_n1620_n5888# 0.012932f
C263 drain_left.n244 a_n1620_n5888# 0.012214f
C264 drain_left.n245 a_n1620_n5888# 0.02273f
C265 drain_left.n246 a_n1620_n5888# 0.02273f
C266 drain_left.n247 a_n1620_n5888# 0.012214f
C267 drain_left.n248 a_n1620_n5888# 0.012932f
C268 drain_left.n249 a_n1620_n5888# 0.028869f
C269 drain_left.n250 a_n1620_n5888# 0.028869f
C270 drain_left.n251 a_n1620_n5888# 0.012932f
C271 drain_left.n252 a_n1620_n5888# 0.012214f
C272 drain_left.n253 a_n1620_n5888# 0.02273f
C273 drain_left.n254 a_n1620_n5888# 0.02273f
C274 drain_left.n255 a_n1620_n5888# 0.012214f
C275 drain_left.n256 a_n1620_n5888# 0.012573f
C276 drain_left.n257 a_n1620_n5888# 0.012573f
C277 drain_left.n258 a_n1620_n5888# 0.028869f
C278 drain_left.n259 a_n1620_n5888# 0.028869f
C279 drain_left.n260 a_n1620_n5888# 0.012932f
C280 drain_left.n261 a_n1620_n5888# 0.012214f
C281 drain_left.n262 a_n1620_n5888# 0.02273f
C282 drain_left.n263 a_n1620_n5888# 0.02273f
C283 drain_left.n264 a_n1620_n5888# 0.012214f
C284 drain_left.n265 a_n1620_n5888# 0.012932f
C285 drain_left.n266 a_n1620_n5888# 0.028869f
C286 drain_left.n267 a_n1620_n5888# 0.028869f
C287 drain_left.n268 a_n1620_n5888# 0.012932f
C288 drain_left.n269 a_n1620_n5888# 0.012214f
C289 drain_left.n270 a_n1620_n5888# 0.02273f
C290 drain_left.n271 a_n1620_n5888# 0.02273f
C291 drain_left.n272 a_n1620_n5888# 0.012214f
C292 drain_left.n273 a_n1620_n5888# 0.012932f
C293 drain_left.n274 a_n1620_n5888# 0.028869f
C294 drain_left.n275 a_n1620_n5888# 0.061412f
C295 drain_left.n276 a_n1620_n5888# 0.012932f
C296 drain_left.n277 a_n1620_n5888# 0.012214f
C297 drain_left.n278 a_n1620_n5888# 0.050054f
C298 drain_left.n279 a_n1620_n5888# 0.052182f
C299 drain_left.t2 a_n1620_n5888# 0.449041f
C300 drain_left.t4 a_n1620_n5888# 0.449041f
C301 drain_left.n280 a_n1620_n5888# 4.13839f
C302 drain_left.n281 a_n1620_n5888# 0.650046f
C303 plus.n0 a_n1620_n5888# 0.188159f
C304 plus.t1 a_n1620_n5888# 2.45974f
C305 plus.t3 a_n1620_n5888# 2.45974f
C306 plus.t4 a_n1620_n5888# 2.48524f
C307 plus.n1 a_n1620_n5888# 0.875035f
C308 plus.n2 a_n1620_n5888# 0.898986f
C309 plus.n3 a_n1620_n5888# 0.009876f
C310 plus.n4 a_n1620_n5888# 0.894754f
C311 plus.n5 a_n1620_n5888# 0.798522f
C312 plus.n6 a_n1620_n5888# 0.188159f
C313 plus.t2 a_n1620_n5888# 2.45974f
C314 plus.t5 a_n1620_n5888# 2.48524f
C315 plus.n7 a_n1620_n5888# 0.875035f
C316 plus.t0 a_n1620_n5888# 2.45974f
C317 plus.n8 a_n1620_n5888# 0.898986f
C318 plus.n9 a_n1620_n5888# 0.009876f
C319 plus.n10 a_n1620_n5888# 0.894754f
C320 plus.n11 a_n1620_n5888# 1.65048f
C321 drain_right.n0 a_n1620_n5888# 0.031322f
C322 drain_right.n1 a_n1620_n5888# 0.02272f
C323 drain_right.n2 a_n1620_n5888# 0.012209f
C324 drain_right.n3 a_n1620_n5888# 0.028857f
C325 drain_right.n4 a_n1620_n5888# 0.012927f
C326 drain_right.n5 a_n1620_n5888# 0.02272f
C327 drain_right.n6 a_n1620_n5888# 0.012209f
C328 drain_right.n7 a_n1620_n5888# 0.028857f
C329 drain_right.n8 a_n1620_n5888# 0.012927f
C330 drain_right.n9 a_n1620_n5888# 0.02272f
C331 drain_right.n10 a_n1620_n5888# 0.012209f
C332 drain_right.n11 a_n1620_n5888# 0.028857f
C333 drain_right.n12 a_n1620_n5888# 0.012927f
C334 drain_right.n13 a_n1620_n5888# 0.02272f
C335 drain_right.n14 a_n1620_n5888# 0.012209f
C336 drain_right.n15 a_n1620_n5888# 0.028857f
C337 drain_right.n16 a_n1620_n5888# 0.012927f
C338 drain_right.n17 a_n1620_n5888# 0.02272f
C339 drain_right.n18 a_n1620_n5888# 0.012209f
C340 drain_right.n19 a_n1620_n5888# 0.028857f
C341 drain_right.n20 a_n1620_n5888# 0.012927f
C342 drain_right.n21 a_n1620_n5888# 0.02272f
C343 drain_right.n22 a_n1620_n5888# 0.012209f
C344 drain_right.n23 a_n1620_n5888# 0.028857f
C345 drain_right.n24 a_n1620_n5888# 0.012927f
C346 drain_right.n25 a_n1620_n5888# 0.02272f
C347 drain_right.n26 a_n1620_n5888# 0.012209f
C348 drain_right.n27 a_n1620_n5888# 0.028857f
C349 drain_right.n28 a_n1620_n5888# 0.012927f
C350 drain_right.n29 a_n1620_n5888# 0.02272f
C351 drain_right.n30 a_n1620_n5888# 0.012209f
C352 drain_right.n31 a_n1620_n5888# 0.028857f
C353 drain_right.n32 a_n1620_n5888# 0.012927f
C354 drain_right.n33 a_n1620_n5888# 0.02272f
C355 drain_right.n34 a_n1620_n5888# 0.012568f
C356 drain_right.n35 a_n1620_n5888# 0.028857f
C357 drain_right.n36 a_n1620_n5888# 0.012927f
C358 drain_right.n37 a_n1620_n5888# 0.02272f
C359 drain_right.n38 a_n1620_n5888# 0.012209f
C360 drain_right.n39 a_n1620_n5888# 0.028857f
C361 drain_right.n40 a_n1620_n5888# 0.012927f
C362 drain_right.n41 a_n1620_n5888# 0.02272f
C363 drain_right.n42 a_n1620_n5888# 0.012209f
C364 drain_right.n43 a_n1620_n5888# 0.021643f
C365 drain_right.n44 a_n1620_n5888# 0.0204f
C366 drain_right.t5 a_n1620_n5888# 0.050329f
C367 drain_right.n45 a_n1620_n5888# 0.277207f
C368 drain_right.n46 a_n1620_n5888# 2.45995f
C369 drain_right.n47 a_n1620_n5888# 0.012209f
C370 drain_right.n48 a_n1620_n5888# 0.012927f
C371 drain_right.n49 a_n1620_n5888# 0.028857f
C372 drain_right.n50 a_n1620_n5888# 0.028857f
C373 drain_right.n51 a_n1620_n5888# 0.012927f
C374 drain_right.n52 a_n1620_n5888# 0.012209f
C375 drain_right.n53 a_n1620_n5888# 0.02272f
C376 drain_right.n54 a_n1620_n5888# 0.02272f
C377 drain_right.n55 a_n1620_n5888# 0.012209f
C378 drain_right.n56 a_n1620_n5888# 0.012927f
C379 drain_right.n57 a_n1620_n5888# 0.028857f
C380 drain_right.n58 a_n1620_n5888# 0.028857f
C381 drain_right.n59 a_n1620_n5888# 0.012927f
C382 drain_right.n60 a_n1620_n5888# 0.012209f
C383 drain_right.n61 a_n1620_n5888# 0.02272f
C384 drain_right.n62 a_n1620_n5888# 0.02272f
C385 drain_right.n63 a_n1620_n5888# 0.012209f
C386 drain_right.n64 a_n1620_n5888# 0.012209f
C387 drain_right.n65 a_n1620_n5888# 0.012927f
C388 drain_right.n66 a_n1620_n5888# 0.028857f
C389 drain_right.n67 a_n1620_n5888# 0.028857f
C390 drain_right.n68 a_n1620_n5888# 0.028857f
C391 drain_right.n69 a_n1620_n5888# 0.012568f
C392 drain_right.n70 a_n1620_n5888# 0.012209f
C393 drain_right.n71 a_n1620_n5888# 0.02272f
C394 drain_right.n72 a_n1620_n5888# 0.02272f
C395 drain_right.n73 a_n1620_n5888# 0.012209f
C396 drain_right.n74 a_n1620_n5888# 0.012927f
C397 drain_right.n75 a_n1620_n5888# 0.028857f
C398 drain_right.n76 a_n1620_n5888# 0.028857f
C399 drain_right.n77 a_n1620_n5888# 0.012927f
C400 drain_right.n78 a_n1620_n5888# 0.012209f
C401 drain_right.n79 a_n1620_n5888# 0.02272f
C402 drain_right.n80 a_n1620_n5888# 0.02272f
C403 drain_right.n81 a_n1620_n5888# 0.012209f
C404 drain_right.n82 a_n1620_n5888# 0.012927f
C405 drain_right.n83 a_n1620_n5888# 0.028857f
C406 drain_right.n84 a_n1620_n5888# 0.028857f
C407 drain_right.n85 a_n1620_n5888# 0.012927f
C408 drain_right.n86 a_n1620_n5888# 0.012209f
C409 drain_right.n87 a_n1620_n5888# 0.02272f
C410 drain_right.n88 a_n1620_n5888# 0.02272f
C411 drain_right.n89 a_n1620_n5888# 0.012209f
C412 drain_right.n90 a_n1620_n5888# 0.012927f
C413 drain_right.n91 a_n1620_n5888# 0.028857f
C414 drain_right.n92 a_n1620_n5888# 0.028857f
C415 drain_right.n93 a_n1620_n5888# 0.012927f
C416 drain_right.n94 a_n1620_n5888# 0.012209f
C417 drain_right.n95 a_n1620_n5888# 0.02272f
C418 drain_right.n96 a_n1620_n5888# 0.02272f
C419 drain_right.n97 a_n1620_n5888# 0.012209f
C420 drain_right.n98 a_n1620_n5888# 0.012927f
C421 drain_right.n99 a_n1620_n5888# 0.028857f
C422 drain_right.n100 a_n1620_n5888# 0.028857f
C423 drain_right.n101 a_n1620_n5888# 0.012927f
C424 drain_right.n102 a_n1620_n5888# 0.012209f
C425 drain_right.n103 a_n1620_n5888# 0.02272f
C426 drain_right.n104 a_n1620_n5888# 0.02272f
C427 drain_right.n105 a_n1620_n5888# 0.012209f
C428 drain_right.n106 a_n1620_n5888# 0.012927f
C429 drain_right.n107 a_n1620_n5888# 0.028857f
C430 drain_right.n108 a_n1620_n5888# 0.028857f
C431 drain_right.n109 a_n1620_n5888# 0.028857f
C432 drain_right.n110 a_n1620_n5888# 0.012927f
C433 drain_right.n111 a_n1620_n5888# 0.012209f
C434 drain_right.n112 a_n1620_n5888# 0.02272f
C435 drain_right.n113 a_n1620_n5888# 0.02272f
C436 drain_right.n114 a_n1620_n5888# 0.012209f
C437 drain_right.n115 a_n1620_n5888# 0.012568f
C438 drain_right.n116 a_n1620_n5888# 0.012568f
C439 drain_right.n117 a_n1620_n5888# 0.028857f
C440 drain_right.n118 a_n1620_n5888# 0.028857f
C441 drain_right.n119 a_n1620_n5888# 0.012927f
C442 drain_right.n120 a_n1620_n5888# 0.012209f
C443 drain_right.n121 a_n1620_n5888# 0.02272f
C444 drain_right.n122 a_n1620_n5888# 0.02272f
C445 drain_right.n123 a_n1620_n5888# 0.012209f
C446 drain_right.n124 a_n1620_n5888# 0.012927f
C447 drain_right.n125 a_n1620_n5888# 0.028857f
C448 drain_right.n126 a_n1620_n5888# 0.028857f
C449 drain_right.n127 a_n1620_n5888# 0.012927f
C450 drain_right.n128 a_n1620_n5888# 0.012209f
C451 drain_right.n129 a_n1620_n5888# 0.02272f
C452 drain_right.n130 a_n1620_n5888# 0.02272f
C453 drain_right.n131 a_n1620_n5888# 0.012209f
C454 drain_right.n132 a_n1620_n5888# 0.012927f
C455 drain_right.n133 a_n1620_n5888# 0.028857f
C456 drain_right.n134 a_n1620_n5888# 0.061387f
C457 drain_right.n135 a_n1620_n5888# 0.012927f
C458 drain_right.n136 a_n1620_n5888# 0.012209f
C459 drain_right.n137 a_n1620_n5888# 0.050034f
C460 drain_right.n138 a_n1620_n5888# 0.05117f
C461 drain_right.t2 a_n1620_n5888# 0.448858f
C462 drain_right.t0 a_n1620_n5888# 0.448858f
C463 drain_right.n139 a_n1620_n5888# 4.13764f
C464 drain_right.n140 a_n1620_n5888# 2.16186f
C465 drain_right.t3 a_n1620_n5888# 0.448858f
C466 drain_right.t1 a_n1620_n5888# 0.448858f
C467 drain_right.n141 a_n1620_n5888# 4.14231f
C468 drain_right.n142 a_n1620_n5888# 0.031322f
C469 drain_right.n143 a_n1620_n5888# 0.02272f
C470 drain_right.n144 a_n1620_n5888# 0.012209f
C471 drain_right.n145 a_n1620_n5888# 0.028857f
C472 drain_right.n146 a_n1620_n5888# 0.012927f
C473 drain_right.n147 a_n1620_n5888# 0.02272f
C474 drain_right.n148 a_n1620_n5888# 0.012209f
C475 drain_right.n149 a_n1620_n5888# 0.028857f
C476 drain_right.n150 a_n1620_n5888# 0.012927f
C477 drain_right.n151 a_n1620_n5888# 0.02272f
C478 drain_right.n152 a_n1620_n5888# 0.012209f
C479 drain_right.n153 a_n1620_n5888# 0.028857f
C480 drain_right.n154 a_n1620_n5888# 0.012927f
C481 drain_right.n155 a_n1620_n5888# 0.02272f
C482 drain_right.n156 a_n1620_n5888# 0.012209f
C483 drain_right.n157 a_n1620_n5888# 0.028857f
C484 drain_right.n158 a_n1620_n5888# 0.028857f
C485 drain_right.n159 a_n1620_n5888# 0.012927f
C486 drain_right.n160 a_n1620_n5888# 0.02272f
C487 drain_right.n161 a_n1620_n5888# 0.012209f
C488 drain_right.n162 a_n1620_n5888# 0.028857f
C489 drain_right.n163 a_n1620_n5888# 0.012927f
C490 drain_right.n164 a_n1620_n5888# 0.02272f
C491 drain_right.n165 a_n1620_n5888# 0.012209f
C492 drain_right.n166 a_n1620_n5888# 0.028857f
C493 drain_right.n167 a_n1620_n5888# 0.012927f
C494 drain_right.n168 a_n1620_n5888# 0.02272f
C495 drain_right.n169 a_n1620_n5888# 0.012209f
C496 drain_right.n170 a_n1620_n5888# 0.028857f
C497 drain_right.n171 a_n1620_n5888# 0.012927f
C498 drain_right.n172 a_n1620_n5888# 0.02272f
C499 drain_right.n173 a_n1620_n5888# 0.012209f
C500 drain_right.n174 a_n1620_n5888# 0.028857f
C501 drain_right.n175 a_n1620_n5888# 0.012927f
C502 drain_right.n176 a_n1620_n5888# 0.02272f
C503 drain_right.n177 a_n1620_n5888# 0.012568f
C504 drain_right.n178 a_n1620_n5888# 0.028857f
C505 drain_right.n179 a_n1620_n5888# 0.012209f
C506 drain_right.n180 a_n1620_n5888# 0.012927f
C507 drain_right.n181 a_n1620_n5888# 0.02272f
C508 drain_right.n182 a_n1620_n5888# 0.012209f
C509 drain_right.n183 a_n1620_n5888# 0.028857f
C510 drain_right.n184 a_n1620_n5888# 0.012927f
C511 drain_right.n185 a_n1620_n5888# 0.02272f
C512 drain_right.n186 a_n1620_n5888# 0.012209f
C513 drain_right.n187 a_n1620_n5888# 0.021643f
C514 drain_right.n188 a_n1620_n5888# 0.0204f
C515 drain_right.t4 a_n1620_n5888# 0.050329f
C516 drain_right.n189 a_n1620_n5888# 0.277207f
C517 drain_right.n190 a_n1620_n5888# 2.45995f
C518 drain_right.n191 a_n1620_n5888# 0.012209f
C519 drain_right.n192 a_n1620_n5888# 0.012927f
C520 drain_right.n193 a_n1620_n5888# 0.028857f
C521 drain_right.n194 a_n1620_n5888# 0.028857f
C522 drain_right.n195 a_n1620_n5888# 0.012927f
C523 drain_right.n196 a_n1620_n5888# 0.012209f
C524 drain_right.n197 a_n1620_n5888# 0.02272f
C525 drain_right.n198 a_n1620_n5888# 0.02272f
C526 drain_right.n199 a_n1620_n5888# 0.012209f
C527 drain_right.n200 a_n1620_n5888# 0.012927f
C528 drain_right.n201 a_n1620_n5888# 0.028857f
C529 drain_right.n202 a_n1620_n5888# 0.028857f
C530 drain_right.n203 a_n1620_n5888# 0.012927f
C531 drain_right.n204 a_n1620_n5888# 0.012209f
C532 drain_right.n205 a_n1620_n5888# 0.02272f
C533 drain_right.n206 a_n1620_n5888# 0.02272f
C534 drain_right.n207 a_n1620_n5888# 0.012209f
C535 drain_right.n208 a_n1620_n5888# 0.012927f
C536 drain_right.n209 a_n1620_n5888# 0.028857f
C537 drain_right.n210 a_n1620_n5888# 0.028857f
C538 drain_right.n211 a_n1620_n5888# 0.028857f
C539 drain_right.n212 a_n1620_n5888# 0.012568f
C540 drain_right.n213 a_n1620_n5888# 0.012209f
C541 drain_right.n214 a_n1620_n5888# 0.02272f
C542 drain_right.n215 a_n1620_n5888# 0.02272f
C543 drain_right.n216 a_n1620_n5888# 0.012209f
C544 drain_right.n217 a_n1620_n5888# 0.012927f
C545 drain_right.n218 a_n1620_n5888# 0.028857f
C546 drain_right.n219 a_n1620_n5888# 0.028857f
C547 drain_right.n220 a_n1620_n5888# 0.012927f
C548 drain_right.n221 a_n1620_n5888# 0.012209f
C549 drain_right.n222 a_n1620_n5888# 0.02272f
C550 drain_right.n223 a_n1620_n5888# 0.02272f
C551 drain_right.n224 a_n1620_n5888# 0.012209f
C552 drain_right.n225 a_n1620_n5888# 0.012927f
C553 drain_right.n226 a_n1620_n5888# 0.028857f
C554 drain_right.n227 a_n1620_n5888# 0.028857f
C555 drain_right.n228 a_n1620_n5888# 0.012927f
C556 drain_right.n229 a_n1620_n5888# 0.012209f
C557 drain_right.n230 a_n1620_n5888# 0.02272f
C558 drain_right.n231 a_n1620_n5888# 0.02272f
C559 drain_right.n232 a_n1620_n5888# 0.012209f
C560 drain_right.n233 a_n1620_n5888# 0.012927f
C561 drain_right.n234 a_n1620_n5888# 0.028857f
C562 drain_right.n235 a_n1620_n5888# 0.028857f
C563 drain_right.n236 a_n1620_n5888# 0.012927f
C564 drain_right.n237 a_n1620_n5888# 0.012209f
C565 drain_right.n238 a_n1620_n5888# 0.02272f
C566 drain_right.n239 a_n1620_n5888# 0.02272f
C567 drain_right.n240 a_n1620_n5888# 0.012209f
C568 drain_right.n241 a_n1620_n5888# 0.012927f
C569 drain_right.n242 a_n1620_n5888# 0.028857f
C570 drain_right.n243 a_n1620_n5888# 0.028857f
C571 drain_right.n244 a_n1620_n5888# 0.012927f
C572 drain_right.n245 a_n1620_n5888# 0.012209f
C573 drain_right.n246 a_n1620_n5888# 0.02272f
C574 drain_right.n247 a_n1620_n5888# 0.02272f
C575 drain_right.n248 a_n1620_n5888# 0.012209f
C576 drain_right.n249 a_n1620_n5888# 0.012927f
C577 drain_right.n250 a_n1620_n5888# 0.028857f
C578 drain_right.n251 a_n1620_n5888# 0.028857f
C579 drain_right.n252 a_n1620_n5888# 0.012927f
C580 drain_right.n253 a_n1620_n5888# 0.012209f
C581 drain_right.n254 a_n1620_n5888# 0.02272f
C582 drain_right.n255 a_n1620_n5888# 0.02272f
C583 drain_right.n256 a_n1620_n5888# 0.012209f
C584 drain_right.n257 a_n1620_n5888# 0.012568f
C585 drain_right.n258 a_n1620_n5888# 0.012568f
C586 drain_right.n259 a_n1620_n5888# 0.028857f
C587 drain_right.n260 a_n1620_n5888# 0.028857f
C588 drain_right.n261 a_n1620_n5888# 0.012927f
C589 drain_right.n262 a_n1620_n5888# 0.012209f
C590 drain_right.n263 a_n1620_n5888# 0.02272f
C591 drain_right.n264 a_n1620_n5888# 0.02272f
C592 drain_right.n265 a_n1620_n5888# 0.012209f
C593 drain_right.n266 a_n1620_n5888# 0.012927f
C594 drain_right.n267 a_n1620_n5888# 0.028857f
C595 drain_right.n268 a_n1620_n5888# 0.028857f
C596 drain_right.n269 a_n1620_n5888# 0.012927f
C597 drain_right.n270 a_n1620_n5888# 0.012209f
C598 drain_right.n271 a_n1620_n5888# 0.02272f
C599 drain_right.n272 a_n1620_n5888# 0.02272f
C600 drain_right.n273 a_n1620_n5888# 0.012209f
C601 drain_right.n274 a_n1620_n5888# 0.012927f
C602 drain_right.n275 a_n1620_n5888# 0.028857f
C603 drain_right.n276 a_n1620_n5888# 0.061387f
C604 drain_right.n277 a_n1620_n5888# 0.012927f
C605 drain_right.n278 a_n1620_n5888# 0.012209f
C606 drain_right.n279 a_n1620_n5888# 0.050034f
C607 drain_right.n280 a_n1620_n5888# 0.049868f
C608 drain_right.n281 a_n1620_n5888# 0.665453f
C609 source.n0 a_n1620_n5888# 0.031419f
C610 source.n1 a_n1620_n5888# 0.022791f
C611 source.n2 a_n1620_n5888# 0.012247f
C612 source.n3 a_n1620_n5888# 0.028947f
C613 source.n4 a_n1620_n5888# 0.012967f
C614 source.n5 a_n1620_n5888# 0.022791f
C615 source.n6 a_n1620_n5888# 0.012247f
C616 source.n7 a_n1620_n5888# 0.028947f
C617 source.n8 a_n1620_n5888# 0.012967f
C618 source.n9 a_n1620_n5888# 0.022791f
C619 source.n10 a_n1620_n5888# 0.012247f
C620 source.n11 a_n1620_n5888# 0.028947f
C621 source.n12 a_n1620_n5888# 0.012967f
C622 source.n13 a_n1620_n5888# 0.022791f
C623 source.n14 a_n1620_n5888# 0.012247f
C624 source.n15 a_n1620_n5888# 0.028947f
C625 source.n16 a_n1620_n5888# 0.028947f
C626 source.n17 a_n1620_n5888# 0.012967f
C627 source.n18 a_n1620_n5888# 0.022791f
C628 source.n19 a_n1620_n5888# 0.012247f
C629 source.n20 a_n1620_n5888# 0.028947f
C630 source.n21 a_n1620_n5888# 0.012967f
C631 source.n22 a_n1620_n5888# 0.022791f
C632 source.n23 a_n1620_n5888# 0.012247f
C633 source.n24 a_n1620_n5888# 0.028947f
C634 source.n25 a_n1620_n5888# 0.012967f
C635 source.n26 a_n1620_n5888# 0.022791f
C636 source.n27 a_n1620_n5888# 0.012247f
C637 source.n28 a_n1620_n5888# 0.028947f
C638 source.n29 a_n1620_n5888# 0.012967f
C639 source.n30 a_n1620_n5888# 0.022791f
C640 source.n31 a_n1620_n5888# 0.012247f
C641 source.n32 a_n1620_n5888# 0.028947f
C642 source.n33 a_n1620_n5888# 0.012967f
C643 source.n34 a_n1620_n5888# 0.022791f
C644 source.n35 a_n1620_n5888# 0.012607f
C645 source.n36 a_n1620_n5888# 0.028947f
C646 source.n37 a_n1620_n5888# 0.012247f
C647 source.n38 a_n1620_n5888# 0.012967f
C648 source.n39 a_n1620_n5888# 0.022791f
C649 source.n40 a_n1620_n5888# 0.012247f
C650 source.n41 a_n1620_n5888# 0.028947f
C651 source.n42 a_n1620_n5888# 0.012967f
C652 source.n43 a_n1620_n5888# 0.022791f
C653 source.n44 a_n1620_n5888# 0.012247f
C654 source.n45 a_n1620_n5888# 0.02171f
C655 source.n46 a_n1620_n5888# 0.020463f
C656 source.t3 a_n1620_n5888# 0.050485f
C657 source.n47 a_n1620_n5888# 0.278064f
C658 source.n48 a_n1620_n5888# 2.46755f
C659 source.n49 a_n1620_n5888# 0.012247f
C660 source.n50 a_n1620_n5888# 0.012967f
C661 source.n51 a_n1620_n5888# 0.028947f
C662 source.n52 a_n1620_n5888# 0.028947f
C663 source.n53 a_n1620_n5888# 0.012967f
C664 source.n54 a_n1620_n5888# 0.012247f
C665 source.n55 a_n1620_n5888# 0.022791f
C666 source.n56 a_n1620_n5888# 0.022791f
C667 source.n57 a_n1620_n5888# 0.012247f
C668 source.n58 a_n1620_n5888# 0.012967f
C669 source.n59 a_n1620_n5888# 0.028947f
C670 source.n60 a_n1620_n5888# 0.028947f
C671 source.n61 a_n1620_n5888# 0.012967f
C672 source.n62 a_n1620_n5888# 0.012247f
C673 source.n63 a_n1620_n5888# 0.022791f
C674 source.n64 a_n1620_n5888# 0.022791f
C675 source.n65 a_n1620_n5888# 0.012247f
C676 source.n66 a_n1620_n5888# 0.012967f
C677 source.n67 a_n1620_n5888# 0.028947f
C678 source.n68 a_n1620_n5888# 0.028947f
C679 source.n69 a_n1620_n5888# 0.028947f
C680 source.n70 a_n1620_n5888# 0.012607f
C681 source.n71 a_n1620_n5888# 0.012247f
C682 source.n72 a_n1620_n5888# 0.022791f
C683 source.n73 a_n1620_n5888# 0.022791f
C684 source.n74 a_n1620_n5888# 0.012247f
C685 source.n75 a_n1620_n5888# 0.012967f
C686 source.n76 a_n1620_n5888# 0.028947f
C687 source.n77 a_n1620_n5888# 0.028947f
C688 source.n78 a_n1620_n5888# 0.012967f
C689 source.n79 a_n1620_n5888# 0.012247f
C690 source.n80 a_n1620_n5888# 0.022791f
C691 source.n81 a_n1620_n5888# 0.022791f
C692 source.n82 a_n1620_n5888# 0.012247f
C693 source.n83 a_n1620_n5888# 0.012967f
C694 source.n84 a_n1620_n5888# 0.028947f
C695 source.n85 a_n1620_n5888# 0.028947f
C696 source.n86 a_n1620_n5888# 0.012967f
C697 source.n87 a_n1620_n5888# 0.012247f
C698 source.n88 a_n1620_n5888# 0.022791f
C699 source.n89 a_n1620_n5888# 0.022791f
C700 source.n90 a_n1620_n5888# 0.012247f
C701 source.n91 a_n1620_n5888# 0.012967f
C702 source.n92 a_n1620_n5888# 0.028947f
C703 source.n93 a_n1620_n5888# 0.028947f
C704 source.n94 a_n1620_n5888# 0.012967f
C705 source.n95 a_n1620_n5888# 0.012247f
C706 source.n96 a_n1620_n5888# 0.022791f
C707 source.n97 a_n1620_n5888# 0.022791f
C708 source.n98 a_n1620_n5888# 0.012247f
C709 source.n99 a_n1620_n5888# 0.012967f
C710 source.n100 a_n1620_n5888# 0.028947f
C711 source.n101 a_n1620_n5888# 0.028947f
C712 source.n102 a_n1620_n5888# 0.012967f
C713 source.n103 a_n1620_n5888# 0.012247f
C714 source.n104 a_n1620_n5888# 0.022791f
C715 source.n105 a_n1620_n5888# 0.022791f
C716 source.n106 a_n1620_n5888# 0.012247f
C717 source.n107 a_n1620_n5888# 0.012967f
C718 source.n108 a_n1620_n5888# 0.028947f
C719 source.n109 a_n1620_n5888# 0.028947f
C720 source.n110 a_n1620_n5888# 0.012967f
C721 source.n111 a_n1620_n5888# 0.012247f
C722 source.n112 a_n1620_n5888# 0.022791f
C723 source.n113 a_n1620_n5888# 0.022791f
C724 source.n114 a_n1620_n5888# 0.012247f
C725 source.n115 a_n1620_n5888# 0.012607f
C726 source.n116 a_n1620_n5888# 0.012607f
C727 source.n117 a_n1620_n5888# 0.028947f
C728 source.n118 a_n1620_n5888# 0.028947f
C729 source.n119 a_n1620_n5888# 0.012967f
C730 source.n120 a_n1620_n5888# 0.012247f
C731 source.n121 a_n1620_n5888# 0.022791f
C732 source.n122 a_n1620_n5888# 0.022791f
C733 source.n123 a_n1620_n5888# 0.012247f
C734 source.n124 a_n1620_n5888# 0.012967f
C735 source.n125 a_n1620_n5888# 0.028947f
C736 source.n126 a_n1620_n5888# 0.028947f
C737 source.n127 a_n1620_n5888# 0.012967f
C738 source.n128 a_n1620_n5888# 0.012247f
C739 source.n129 a_n1620_n5888# 0.022791f
C740 source.n130 a_n1620_n5888# 0.022791f
C741 source.n131 a_n1620_n5888# 0.012247f
C742 source.n132 a_n1620_n5888# 0.012967f
C743 source.n133 a_n1620_n5888# 0.028947f
C744 source.n134 a_n1620_n5888# 0.061577f
C745 source.n135 a_n1620_n5888# 0.012967f
C746 source.n136 a_n1620_n5888# 0.012247f
C747 source.n137 a_n1620_n5888# 0.050189f
C748 source.n138 a_n1620_n5888# 0.034265f
C749 source.n139 a_n1620_n5888# 1.84017f
C750 source.t2 a_n1620_n5888# 0.450245f
C751 source.t1 a_n1620_n5888# 0.450245f
C752 source.n140 a_n1620_n5888# 4.07478f
C753 source.n141 a_n1620_n5888# 0.378191f
C754 source.n142 a_n1620_n5888# 0.031419f
C755 source.n143 a_n1620_n5888# 0.022791f
C756 source.n144 a_n1620_n5888# 0.012247f
C757 source.n145 a_n1620_n5888# 0.028947f
C758 source.n146 a_n1620_n5888# 0.012967f
C759 source.n147 a_n1620_n5888# 0.022791f
C760 source.n148 a_n1620_n5888# 0.012247f
C761 source.n149 a_n1620_n5888# 0.028947f
C762 source.n150 a_n1620_n5888# 0.012967f
C763 source.n151 a_n1620_n5888# 0.022791f
C764 source.n152 a_n1620_n5888# 0.012247f
C765 source.n153 a_n1620_n5888# 0.028947f
C766 source.n154 a_n1620_n5888# 0.012967f
C767 source.n155 a_n1620_n5888# 0.022791f
C768 source.n156 a_n1620_n5888# 0.012247f
C769 source.n157 a_n1620_n5888# 0.028947f
C770 source.n158 a_n1620_n5888# 0.028947f
C771 source.n159 a_n1620_n5888# 0.012967f
C772 source.n160 a_n1620_n5888# 0.022791f
C773 source.n161 a_n1620_n5888# 0.012247f
C774 source.n162 a_n1620_n5888# 0.028947f
C775 source.n163 a_n1620_n5888# 0.012967f
C776 source.n164 a_n1620_n5888# 0.022791f
C777 source.n165 a_n1620_n5888# 0.012247f
C778 source.n166 a_n1620_n5888# 0.028947f
C779 source.n167 a_n1620_n5888# 0.012967f
C780 source.n168 a_n1620_n5888# 0.022791f
C781 source.n169 a_n1620_n5888# 0.012247f
C782 source.n170 a_n1620_n5888# 0.028947f
C783 source.n171 a_n1620_n5888# 0.012967f
C784 source.n172 a_n1620_n5888# 0.022791f
C785 source.n173 a_n1620_n5888# 0.012247f
C786 source.n174 a_n1620_n5888# 0.028947f
C787 source.n175 a_n1620_n5888# 0.012967f
C788 source.n176 a_n1620_n5888# 0.022791f
C789 source.n177 a_n1620_n5888# 0.012607f
C790 source.n178 a_n1620_n5888# 0.028947f
C791 source.n179 a_n1620_n5888# 0.012247f
C792 source.n180 a_n1620_n5888# 0.012967f
C793 source.n181 a_n1620_n5888# 0.022791f
C794 source.n182 a_n1620_n5888# 0.012247f
C795 source.n183 a_n1620_n5888# 0.028947f
C796 source.n184 a_n1620_n5888# 0.012967f
C797 source.n185 a_n1620_n5888# 0.022791f
C798 source.n186 a_n1620_n5888# 0.012247f
C799 source.n187 a_n1620_n5888# 0.02171f
C800 source.n188 a_n1620_n5888# 0.020463f
C801 source.t8 a_n1620_n5888# 0.050485f
C802 source.n189 a_n1620_n5888# 0.278064f
C803 source.n190 a_n1620_n5888# 2.46755f
C804 source.n191 a_n1620_n5888# 0.012247f
C805 source.n192 a_n1620_n5888# 0.012967f
C806 source.n193 a_n1620_n5888# 0.028947f
C807 source.n194 a_n1620_n5888# 0.028947f
C808 source.n195 a_n1620_n5888# 0.012967f
C809 source.n196 a_n1620_n5888# 0.012247f
C810 source.n197 a_n1620_n5888# 0.022791f
C811 source.n198 a_n1620_n5888# 0.022791f
C812 source.n199 a_n1620_n5888# 0.012247f
C813 source.n200 a_n1620_n5888# 0.012967f
C814 source.n201 a_n1620_n5888# 0.028947f
C815 source.n202 a_n1620_n5888# 0.028947f
C816 source.n203 a_n1620_n5888# 0.012967f
C817 source.n204 a_n1620_n5888# 0.012247f
C818 source.n205 a_n1620_n5888# 0.022791f
C819 source.n206 a_n1620_n5888# 0.022791f
C820 source.n207 a_n1620_n5888# 0.012247f
C821 source.n208 a_n1620_n5888# 0.012967f
C822 source.n209 a_n1620_n5888# 0.028947f
C823 source.n210 a_n1620_n5888# 0.028947f
C824 source.n211 a_n1620_n5888# 0.028947f
C825 source.n212 a_n1620_n5888# 0.012607f
C826 source.n213 a_n1620_n5888# 0.012247f
C827 source.n214 a_n1620_n5888# 0.022791f
C828 source.n215 a_n1620_n5888# 0.022791f
C829 source.n216 a_n1620_n5888# 0.012247f
C830 source.n217 a_n1620_n5888# 0.012967f
C831 source.n218 a_n1620_n5888# 0.028947f
C832 source.n219 a_n1620_n5888# 0.028947f
C833 source.n220 a_n1620_n5888# 0.012967f
C834 source.n221 a_n1620_n5888# 0.012247f
C835 source.n222 a_n1620_n5888# 0.022791f
C836 source.n223 a_n1620_n5888# 0.022791f
C837 source.n224 a_n1620_n5888# 0.012247f
C838 source.n225 a_n1620_n5888# 0.012967f
C839 source.n226 a_n1620_n5888# 0.028947f
C840 source.n227 a_n1620_n5888# 0.028947f
C841 source.n228 a_n1620_n5888# 0.012967f
C842 source.n229 a_n1620_n5888# 0.012247f
C843 source.n230 a_n1620_n5888# 0.022791f
C844 source.n231 a_n1620_n5888# 0.022791f
C845 source.n232 a_n1620_n5888# 0.012247f
C846 source.n233 a_n1620_n5888# 0.012967f
C847 source.n234 a_n1620_n5888# 0.028947f
C848 source.n235 a_n1620_n5888# 0.028947f
C849 source.n236 a_n1620_n5888# 0.012967f
C850 source.n237 a_n1620_n5888# 0.012247f
C851 source.n238 a_n1620_n5888# 0.022791f
C852 source.n239 a_n1620_n5888# 0.022791f
C853 source.n240 a_n1620_n5888# 0.012247f
C854 source.n241 a_n1620_n5888# 0.012967f
C855 source.n242 a_n1620_n5888# 0.028947f
C856 source.n243 a_n1620_n5888# 0.028947f
C857 source.n244 a_n1620_n5888# 0.012967f
C858 source.n245 a_n1620_n5888# 0.012247f
C859 source.n246 a_n1620_n5888# 0.022791f
C860 source.n247 a_n1620_n5888# 0.022791f
C861 source.n248 a_n1620_n5888# 0.012247f
C862 source.n249 a_n1620_n5888# 0.012967f
C863 source.n250 a_n1620_n5888# 0.028947f
C864 source.n251 a_n1620_n5888# 0.028947f
C865 source.n252 a_n1620_n5888# 0.012967f
C866 source.n253 a_n1620_n5888# 0.012247f
C867 source.n254 a_n1620_n5888# 0.022791f
C868 source.n255 a_n1620_n5888# 0.022791f
C869 source.n256 a_n1620_n5888# 0.012247f
C870 source.n257 a_n1620_n5888# 0.012607f
C871 source.n258 a_n1620_n5888# 0.012607f
C872 source.n259 a_n1620_n5888# 0.028947f
C873 source.n260 a_n1620_n5888# 0.028947f
C874 source.n261 a_n1620_n5888# 0.012967f
C875 source.n262 a_n1620_n5888# 0.012247f
C876 source.n263 a_n1620_n5888# 0.022791f
C877 source.n264 a_n1620_n5888# 0.022791f
C878 source.n265 a_n1620_n5888# 0.012247f
C879 source.n266 a_n1620_n5888# 0.012967f
C880 source.n267 a_n1620_n5888# 0.028947f
C881 source.n268 a_n1620_n5888# 0.028947f
C882 source.n269 a_n1620_n5888# 0.012967f
C883 source.n270 a_n1620_n5888# 0.012247f
C884 source.n271 a_n1620_n5888# 0.022791f
C885 source.n272 a_n1620_n5888# 0.022791f
C886 source.n273 a_n1620_n5888# 0.012247f
C887 source.n274 a_n1620_n5888# 0.012967f
C888 source.n275 a_n1620_n5888# 0.028947f
C889 source.n276 a_n1620_n5888# 0.061577f
C890 source.n277 a_n1620_n5888# 0.012967f
C891 source.n278 a_n1620_n5888# 0.012247f
C892 source.n279 a_n1620_n5888# 0.050189f
C893 source.n280 a_n1620_n5888# 0.034265f
C894 source.n281 a_n1620_n5888# 0.159869f
C895 source.t11 a_n1620_n5888# 0.450245f
C896 source.t6 a_n1620_n5888# 0.450245f
C897 source.n282 a_n1620_n5888# 4.07478f
C898 source.n283 a_n1620_n5888# 2.56594f
C899 source.t0 a_n1620_n5888# 0.450245f
C900 source.t4 a_n1620_n5888# 0.450245f
C901 source.n284 a_n1620_n5888# 4.07478f
C902 source.n285 a_n1620_n5888# 2.56595f
C903 source.n286 a_n1620_n5888# 0.031419f
C904 source.n287 a_n1620_n5888# 0.022791f
C905 source.n288 a_n1620_n5888# 0.012247f
C906 source.n289 a_n1620_n5888# 0.028947f
C907 source.n290 a_n1620_n5888# 0.012967f
C908 source.n291 a_n1620_n5888# 0.022791f
C909 source.n292 a_n1620_n5888# 0.012247f
C910 source.n293 a_n1620_n5888# 0.028947f
C911 source.n294 a_n1620_n5888# 0.012967f
C912 source.n295 a_n1620_n5888# 0.022791f
C913 source.n296 a_n1620_n5888# 0.012247f
C914 source.n297 a_n1620_n5888# 0.028947f
C915 source.n298 a_n1620_n5888# 0.012967f
C916 source.n299 a_n1620_n5888# 0.022791f
C917 source.n300 a_n1620_n5888# 0.012247f
C918 source.n301 a_n1620_n5888# 0.028947f
C919 source.n302 a_n1620_n5888# 0.012967f
C920 source.n303 a_n1620_n5888# 0.022791f
C921 source.n304 a_n1620_n5888# 0.012247f
C922 source.n305 a_n1620_n5888# 0.028947f
C923 source.n306 a_n1620_n5888# 0.012967f
C924 source.n307 a_n1620_n5888# 0.022791f
C925 source.n308 a_n1620_n5888# 0.012247f
C926 source.n309 a_n1620_n5888# 0.028947f
C927 source.n310 a_n1620_n5888# 0.012967f
C928 source.n311 a_n1620_n5888# 0.022791f
C929 source.n312 a_n1620_n5888# 0.012247f
C930 source.n313 a_n1620_n5888# 0.028947f
C931 source.n314 a_n1620_n5888# 0.012967f
C932 source.n315 a_n1620_n5888# 0.022791f
C933 source.n316 a_n1620_n5888# 0.012247f
C934 source.n317 a_n1620_n5888# 0.028947f
C935 source.n318 a_n1620_n5888# 0.012967f
C936 source.n319 a_n1620_n5888# 0.022791f
C937 source.n320 a_n1620_n5888# 0.012607f
C938 source.n321 a_n1620_n5888# 0.028947f
C939 source.n322 a_n1620_n5888# 0.012967f
C940 source.n323 a_n1620_n5888# 0.022791f
C941 source.n324 a_n1620_n5888# 0.012247f
C942 source.n325 a_n1620_n5888# 0.028947f
C943 source.n326 a_n1620_n5888# 0.012967f
C944 source.n327 a_n1620_n5888# 0.022791f
C945 source.n328 a_n1620_n5888# 0.012247f
C946 source.n329 a_n1620_n5888# 0.02171f
C947 source.n330 a_n1620_n5888# 0.020463f
C948 source.t5 a_n1620_n5888# 0.050485f
C949 source.n331 a_n1620_n5888# 0.278064f
C950 source.n332 a_n1620_n5888# 2.46755f
C951 source.n333 a_n1620_n5888# 0.012247f
C952 source.n334 a_n1620_n5888# 0.012967f
C953 source.n335 a_n1620_n5888# 0.028947f
C954 source.n336 a_n1620_n5888# 0.028947f
C955 source.n337 a_n1620_n5888# 0.012967f
C956 source.n338 a_n1620_n5888# 0.012247f
C957 source.n339 a_n1620_n5888# 0.022791f
C958 source.n340 a_n1620_n5888# 0.022791f
C959 source.n341 a_n1620_n5888# 0.012247f
C960 source.n342 a_n1620_n5888# 0.012967f
C961 source.n343 a_n1620_n5888# 0.028947f
C962 source.n344 a_n1620_n5888# 0.028947f
C963 source.n345 a_n1620_n5888# 0.012967f
C964 source.n346 a_n1620_n5888# 0.012247f
C965 source.n347 a_n1620_n5888# 0.022791f
C966 source.n348 a_n1620_n5888# 0.022791f
C967 source.n349 a_n1620_n5888# 0.012247f
C968 source.n350 a_n1620_n5888# 0.012247f
C969 source.n351 a_n1620_n5888# 0.012967f
C970 source.n352 a_n1620_n5888# 0.028947f
C971 source.n353 a_n1620_n5888# 0.028947f
C972 source.n354 a_n1620_n5888# 0.028947f
C973 source.n355 a_n1620_n5888# 0.012607f
C974 source.n356 a_n1620_n5888# 0.012247f
C975 source.n357 a_n1620_n5888# 0.022791f
C976 source.n358 a_n1620_n5888# 0.022791f
C977 source.n359 a_n1620_n5888# 0.012247f
C978 source.n360 a_n1620_n5888# 0.012967f
C979 source.n361 a_n1620_n5888# 0.028947f
C980 source.n362 a_n1620_n5888# 0.028947f
C981 source.n363 a_n1620_n5888# 0.012967f
C982 source.n364 a_n1620_n5888# 0.012247f
C983 source.n365 a_n1620_n5888# 0.022791f
C984 source.n366 a_n1620_n5888# 0.022791f
C985 source.n367 a_n1620_n5888# 0.012247f
C986 source.n368 a_n1620_n5888# 0.012967f
C987 source.n369 a_n1620_n5888# 0.028947f
C988 source.n370 a_n1620_n5888# 0.028947f
C989 source.n371 a_n1620_n5888# 0.012967f
C990 source.n372 a_n1620_n5888# 0.012247f
C991 source.n373 a_n1620_n5888# 0.022791f
C992 source.n374 a_n1620_n5888# 0.022791f
C993 source.n375 a_n1620_n5888# 0.012247f
C994 source.n376 a_n1620_n5888# 0.012967f
C995 source.n377 a_n1620_n5888# 0.028947f
C996 source.n378 a_n1620_n5888# 0.028947f
C997 source.n379 a_n1620_n5888# 0.012967f
C998 source.n380 a_n1620_n5888# 0.012247f
C999 source.n381 a_n1620_n5888# 0.022791f
C1000 source.n382 a_n1620_n5888# 0.022791f
C1001 source.n383 a_n1620_n5888# 0.012247f
C1002 source.n384 a_n1620_n5888# 0.012967f
C1003 source.n385 a_n1620_n5888# 0.028947f
C1004 source.n386 a_n1620_n5888# 0.028947f
C1005 source.n387 a_n1620_n5888# 0.012967f
C1006 source.n388 a_n1620_n5888# 0.012247f
C1007 source.n389 a_n1620_n5888# 0.022791f
C1008 source.n390 a_n1620_n5888# 0.022791f
C1009 source.n391 a_n1620_n5888# 0.012247f
C1010 source.n392 a_n1620_n5888# 0.012967f
C1011 source.n393 a_n1620_n5888# 0.028947f
C1012 source.n394 a_n1620_n5888# 0.028947f
C1013 source.n395 a_n1620_n5888# 0.028947f
C1014 source.n396 a_n1620_n5888# 0.012967f
C1015 source.n397 a_n1620_n5888# 0.012247f
C1016 source.n398 a_n1620_n5888# 0.022791f
C1017 source.n399 a_n1620_n5888# 0.022791f
C1018 source.n400 a_n1620_n5888# 0.012247f
C1019 source.n401 a_n1620_n5888# 0.012607f
C1020 source.n402 a_n1620_n5888# 0.012607f
C1021 source.n403 a_n1620_n5888# 0.028947f
C1022 source.n404 a_n1620_n5888# 0.028947f
C1023 source.n405 a_n1620_n5888# 0.012967f
C1024 source.n406 a_n1620_n5888# 0.012247f
C1025 source.n407 a_n1620_n5888# 0.022791f
C1026 source.n408 a_n1620_n5888# 0.022791f
C1027 source.n409 a_n1620_n5888# 0.012247f
C1028 source.n410 a_n1620_n5888# 0.012967f
C1029 source.n411 a_n1620_n5888# 0.028947f
C1030 source.n412 a_n1620_n5888# 0.028947f
C1031 source.n413 a_n1620_n5888# 0.012967f
C1032 source.n414 a_n1620_n5888# 0.012247f
C1033 source.n415 a_n1620_n5888# 0.022791f
C1034 source.n416 a_n1620_n5888# 0.022791f
C1035 source.n417 a_n1620_n5888# 0.012247f
C1036 source.n418 a_n1620_n5888# 0.012967f
C1037 source.n419 a_n1620_n5888# 0.028947f
C1038 source.n420 a_n1620_n5888# 0.061577f
C1039 source.n421 a_n1620_n5888# 0.012967f
C1040 source.n422 a_n1620_n5888# 0.012247f
C1041 source.n423 a_n1620_n5888# 0.050189f
C1042 source.n424 a_n1620_n5888# 0.034265f
C1043 source.n425 a_n1620_n5888# 0.159869f
C1044 source.t7 a_n1620_n5888# 0.450245f
C1045 source.t9 a_n1620_n5888# 0.450245f
C1046 source.n426 a_n1620_n5888# 4.07478f
C1047 source.n427 a_n1620_n5888# 0.378193f
C1048 source.n428 a_n1620_n5888# 0.031419f
C1049 source.n429 a_n1620_n5888# 0.022791f
C1050 source.n430 a_n1620_n5888# 0.012247f
C1051 source.n431 a_n1620_n5888# 0.028947f
C1052 source.n432 a_n1620_n5888# 0.012967f
C1053 source.n433 a_n1620_n5888# 0.022791f
C1054 source.n434 a_n1620_n5888# 0.012247f
C1055 source.n435 a_n1620_n5888# 0.028947f
C1056 source.n436 a_n1620_n5888# 0.012967f
C1057 source.n437 a_n1620_n5888# 0.022791f
C1058 source.n438 a_n1620_n5888# 0.012247f
C1059 source.n439 a_n1620_n5888# 0.028947f
C1060 source.n440 a_n1620_n5888# 0.012967f
C1061 source.n441 a_n1620_n5888# 0.022791f
C1062 source.n442 a_n1620_n5888# 0.012247f
C1063 source.n443 a_n1620_n5888# 0.028947f
C1064 source.n444 a_n1620_n5888# 0.012967f
C1065 source.n445 a_n1620_n5888# 0.022791f
C1066 source.n446 a_n1620_n5888# 0.012247f
C1067 source.n447 a_n1620_n5888# 0.028947f
C1068 source.n448 a_n1620_n5888# 0.012967f
C1069 source.n449 a_n1620_n5888# 0.022791f
C1070 source.n450 a_n1620_n5888# 0.012247f
C1071 source.n451 a_n1620_n5888# 0.028947f
C1072 source.n452 a_n1620_n5888# 0.012967f
C1073 source.n453 a_n1620_n5888# 0.022791f
C1074 source.n454 a_n1620_n5888# 0.012247f
C1075 source.n455 a_n1620_n5888# 0.028947f
C1076 source.n456 a_n1620_n5888# 0.012967f
C1077 source.n457 a_n1620_n5888# 0.022791f
C1078 source.n458 a_n1620_n5888# 0.012247f
C1079 source.n459 a_n1620_n5888# 0.028947f
C1080 source.n460 a_n1620_n5888# 0.012967f
C1081 source.n461 a_n1620_n5888# 0.022791f
C1082 source.n462 a_n1620_n5888# 0.012607f
C1083 source.n463 a_n1620_n5888# 0.028947f
C1084 source.n464 a_n1620_n5888# 0.012967f
C1085 source.n465 a_n1620_n5888# 0.022791f
C1086 source.n466 a_n1620_n5888# 0.012247f
C1087 source.n467 a_n1620_n5888# 0.028947f
C1088 source.n468 a_n1620_n5888# 0.012967f
C1089 source.n469 a_n1620_n5888# 0.022791f
C1090 source.n470 a_n1620_n5888# 0.012247f
C1091 source.n471 a_n1620_n5888# 0.02171f
C1092 source.n472 a_n1620_n5888# 0.020463f
C1093 source.t10 a_n1620_n5888# 0.050485f
C1094 source.n473 a_n1620_n5888# 0.278064f
C1095 source.n474 a_n1620_n5888# 2.46755f
C1096 source.n475 a_n1620_n5888# 0.012247f
C1097 source.n476 a_n1620_n5888# 0.012967f
C1098 source.n477 a_n1620_n5888# 0.028947f
C1099 source.n478 a_n1620_n5888# 0.028947f
C1100 source.n479 a_n1620_n5888# 0.012967f
C1101 source.n480 a_n1620_n5888# 0.012247f
C1102 source.n481 a_n1620_n5888# 0.022791f
C1103 source.n482 a_n1620_n5888# 0.022791f
C1104 source.n483 a_n1620_n5888# 0.012247f
C1105 source.n484 a_n1620_n5888# 0.012967f
C1106 source.n485 a_n1620_n5888# 0.028947f
C1107 source.n486 a_n1620_n5888# 0.028947f
C1108 source.n487 a_n1620_n5888# 0.012967f
C1109 source.n488 a_n1620_n5888# 0.012247f
C1110 source.n489 a_n1620_n5888# 0.022791f
C1111 source.n490 a_n1620_n5888# 0.022791f
C1112 source.n491 a_n1620_n5888# 0.012247f
C1113 source.n492 a_n1620_n5888# 0.012247f
C1114 source.n493 a_n1620_n5888# 0.012967f
C1115 source.n494 a_n1620_n5888# 0.028947f
C1116 source.n495 a_n1620_n5888# 0.028947f
C1117 source.n496 a_n1620_n5888# 0.028947f
C1118 source.n497 a_n1620_n5888# 0.012607f
C1119 source.n498 a_n1620_n5888# 0.012247f
C1120 source.n499 a_n1620_n5888# 0.022791f
C1121 source.n500 a_n1620_n5888# 0.022791f
C1122 source.n501 a_n1620_n5888# 0.012247f
C1123 source.n502 a_n1620_n5888# 0.012967f
C1124 source.n503 a_n1620_n5888# 0.028947f
C1125 source.n504 a_n1620_n5888# 0.028947f
C1126 source.n505 a_n1620_n5888# 0.012967f
C1127 source.n506 a_n1620_n5888# 0.012247f
C1128 source.n507 a_n1620_n5888# 0.022791f
C1129 source.n508 a_n1620_n5888# 0.022791f
C1130 source.n509 a_n1620_n5888# 0.012247f
C1131 source.n510 a_n1620_n5888# 0.012967f
C1132 source.n511 a_n1620_n5888# 0.028947f
C1133 source.n512 a_n1620_n5888# 0.028947f
C1134 source.n513 a_n1620_n5888# 0.012967f
C1135 source.n514 a_n1620_n5888# 0.012247f
C1136 source.n515 a_n1620_n5888# 0.022791f
C1137 source.n516 a_n1620_n5888# 0.022791f
C1138 source.n517 a_n1620_n5888# 0.012247f
C1139 source.n518 a_n1620_n5888# 0.012967f
C1140 source.n519 a_n1620_n5888# 0.028947f
C1141 source.n520 a_n1620_n5888# 0.028947f
C1142 source.n521 a_n1620_n5888# 0.012967f
C1143 source.n522 a_n1620_n5888# 0.012247f
C1144 source.n523 a_n1620_n5888# 0.022791f
C1145 source.n524 a_n1620_n5888# 0.022791f
C1146 source.n525 a_n1620_n5888# 0.012247f
C1147 source.n526 a_n1620_n5888# 0.012967f
C1148 source.n527 a_n1620_n5888# 0.028947f
C1149 source.n528 a_n1620_n5888# 0.028947f
C1150 source.n529 a_n1620_n5888# 0.012967f
C1151 source.n530 a_n1620_n5888# 0.012247f
C1152 source.n531 a_n1620_n5888# 0.022791f
C1153 source.n532 a_n1620_n5888# 0.022791f
C1154 source.n533 a_n1620_n5888# 0.012247f
C1155 source.n534 a_n1620_n5888# 0.012967f
C1156 source.n535 a_n1620_n5888# 0.028947f
C1157 source.n536 a_n1620_n5888# 0.028947f
C1158 source.n537 a_n1620_n5888# 0.028947f
C1159 source.n538 a_n1620_n5888# 0.012967f
C1160 source.n539 a_n1620_n5888# 0.012247f
C1161 source.n540 a_n1620_n5888# 0.022791f
C1162 source.n541 a_n1620_n5888# 0.022791f
C1163 source.n542 a_n1620_n5888# 0.012247f
C1164 source.n543 a_n1620_n5888# 0.012607f
C1165 source.n544 a_n1620_n5888# 0.012607f
C1166 source.n545 a_n1620_n5888# 0.028947f
C1167 source.n546 a_n1620_n5888# 0.028947f
C1168 source.n547 a_n1620_n5888# 0.012967f
C1169 source.n548 a_n1620_n5888# 0.012247f
C1170 source.n549 a_n1620_n5888# 0.022791f
C1171 source.n550 a_n1620_n5888# 0.022791f
C1172 source.n551 a_n1620_n5888# 0.012247f
C1173 source.n552 a_n1620_n5888# 0.012967f
C1174 source.n553 a_n1620_n5888# 0.028947f
C1175 source.n554 a_n1620_n5888# 0.028947f
C1176 source.n555 a_n1620_n5888# 0.012967f
C1177 source.n556 a_n1620_n5888# 0.012247f
C1178 source.n557 a_n1620_n5888# 0.022791f
C1179 source.n558 a_n1620_n5888# 0.022791f
C1180 source.n559 a_n1620_n5888# 0.012247f
C1181 source.n560 a_n1620_n5888# 0.012967f
C1182 source.n561 a_n1620_n5888# 0.028947f
C1183 source.n562 a_n1620_n5888# 0.061577f
C1184 source.n563 a_n1620_n5888# 0.012967f
C1185 source.n564 a_n1620_n5888# 0.012247f
C1186 source.n565 a_n1620_n5888# 0.050189f
C1187 source.n566 a_n1620_n5888# 0.034265f
C1188 source.n567 a_n1620_n5888# 0.277698f
C1189 source.n568 a_n1620_n5888# 2.45052f
C1190 minus.n0 a_n1620_n5888# 0.186777f
C1191 minus.t4 a_n1620_n5888# 2.46698f
C1192 minus.n1 a_n1620_n5888# 0.868605f
C1193 minus.t2 a_n1620_n5888# 2.44167f
C1194 minus.n2 a_n1620_n5888# 0.892381f
C1195 minus.n3 a_n1620_n5888# 0.009803f
C1196 minus.t1 a_n1620_n5888# 2.44167f
C1197 minus.n4 a_n1620_n5888# 0.88818f
C1198 minus.n5 a_n1620_n5888# 2.14311f
C1199 minus.n6 a_n1620_n5888# 0.186777f
C1200 minus.t0 a_n1620_n5888# 2.46698f
C1201 minus.n7 a_n1620_n5888# 0.868605f
C1202 minus.t3 a_n1620_n5888# 2.44167f
C1203 minus.n8 a_n1620_n5888# 0.892381f
C1204 minus.n9 a_n1620_n5888# 0.009803f
C1205 minus.t5 a_n1620_n5888# 2.44167f
C1206 minus.n10 a_n1620_n5888# 0.88818f
C1207 minus.n11 a_n1620_n5888# 0.304802f
C1208 minus.n12 a_n1620_n5888# 2.5316f
.ends

