* NGSPICE file created from diffpair482.ext - technology: sky130A

.subckt diffpair482 minus drain_right drain_left source plus
X0 a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X1 a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X2 drain_right.t5 minus.t0 source.t11 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X3 a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X4 drain_left.t5 plus.t0 source.t2 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X5 source.t10 minus.t1 drain_right.t4 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X6 a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X7 drain_right.t3 minus.t2 source.t6 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X8 drain_left.t4 plus.t1 source.t3 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X9 drain_right.t2 minus.t3 source.t9 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X10 drain_left.t3 plus.t2 source.t1 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X11 source.t7 minus.t4 drain_right.t1 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X12 drain_left.t2 plus.t3 source.t0 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X13 source.t5 plus.t4 drain_left.t1 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X14 source.t4 plus.t5 drain_left.t0 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X15 drain_right.t0 minus.t5 source.t8 a_n1236_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
R0 minus.n2 minus.t3 2677.29
R1 minus.n0 minus.t2 2677.29
R2 minus.n6 minus.t5 2677.29
R3 minus.n4 minus.t0 2677.29
R4 minus.n1 minus.t1 2618.87
R5 minus.n5 minus.t4 2618.87
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 36.1274
R15 minus.n8 minus.n7 6.55164
R16 minus minus.n8 0.188
R17 source.n3 source.t6 46.201
R18 source.n11 source.t8 46.2008
R19 source.n8 source.t1 46.2008
R20 source.n0 source.t0 46.2008
R21 source.n2 source.n1 44.201
R22 source.n5 source.n4 44.201
R23 source.n10 source.n9 44.2008
R24 source.n7 source.n6 44.2008
R25 source.n7 source.n5 24.6811
R26 source.n12 source.n0 18.5777
R27 source.n12 source.n11 5.5436
R28 source.n9 source.t11 2.0005
R29 source.n9 source.t7 2.0005
R30 source.n6 source.t2 2.0005
R31 source.n6 source.t4 2.0005
R32 source.n1 source.t3 2.0005
R33 source.n1 source.t5 2.0005
R34 source.n4 source.t9 2.0005
R35 source.n4 source.t10 2.0005
R36 source.n3 source.n2 0.7505
R37 source.n10 source.n8 0.7505
R38 source.n5 source.n3 0.560845
R39 source.n2 source.n0 0.560845
R40 source.n8 source.n7 0.560845
R41 source.n11 source.n10 0.560845
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t5 63.2445
R44 drain_right.n3 drain_right.t2 62.8798
R45 drain_right.n3 drain_right.n2 61.44
R46 drain_right.n1 drain_right.n0 60.9643
R47 drain_right drain_right.n1 30.6275
R48 drain_right drain_right.n3 5.93339
R49 drain_right.n0 drain_right.t1 2.0005
R50 drain_right.n0 drain_right.t0 2.0005
R51 drain_right.n2 drain_right.t4 2.0005
R52 drain_right.n2 drain_right.t3 2.0005
R53 plus.n0 plus.t1 2677.29
R54 plus.n2 plus.t3 2677.29
R55 plus.n4 plus.t2 2677.29
R56 plus.n6 plus.t0 2677.29
R57 plus.n1 plus.t4 2618.87
R58 plus.n5 plus.t5 2618.87
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 28.8721
R68 plus plus.n3 13.3319
R69 drain_left.n3 drain_left.t4 63.4402
R70 drain_left.n1 drain_left.t5 63.2445
R71 drain_left.n1 drain_left.n0 60.9643
R72 drain_left.n3 drain_left.n2 60.8796
R73 drain_left drain_left.n1 31.1808
R74 drain_left drain_left.n3 6.21356
R75 drain_left.n0 drain_left.t0 2.0005
R76 drain_left.n0 drain_left.t3 2.0005
R77 drain_left.n2 drain_left.t1 2.0005
R78 drain_left.n2 drain_left.t2 2.0005
C0 minus drain_left 0.170478f
C1 source plus 1.5196f
C2 minus plus 5.23042f
C3 source drain_right 17.4975f
C4 minus drain_right 2.21909f
C5 minus source 1.50475f
C6 drain_left plus 2.33147f
C7 drain_left drain_right 0.57706f
C8 drain_left source 17.5113f
C9 drain_right plus 0.271684f
C10 drain_right a_n1236_n3888# 6.89656f
C11 drain_left a_n1236_n3888# 7.07905f
C12 source a_n1236_n3888# 7.146767f
C13 minus a_n1236_n3888# 4.71124f
C14 plus a_n1236_n3888# 6.76134f
C15 drain_left.t5 a_n1236_n3888# 3.56622f
C16 drain_left.t0 a_n1236_n3888# 0.434199f
C17 drain_left.t3 a_n1236_n3888# 0.434199f
C18 drain_left.n0 a_n1236_n3888# 2.88589f
C19 drain_left.n1 a_n1236_n3888# 1.8037f
C20 drain_left.t4 a_n1236_n3888# 3.56739f
C21 drain_left.t1 a_n1236_n3888# 0.434199f
C22 drain_left.t2 a_n1236_n3888# 0.434199f
C23 drain_left.n2 a_n1236_n3888# 2.88552f
C24 drain_left.n3 a_n1236_n3888# 0.838329f
C25 plus.t1 a_n1236_n3888# 0.339698f
C26 plus.n0 a_n1236_n3888# 0.158667f
C27 plus.t4 a_n1236_n3888# 0.336662f
C28 plus.n1 a_n1236_n3888# 0.137489f
C29 plus.t3 a_n1236_n3888# 0.339698f
C30 plus.n2 a_n1236_n3888# 0.158587f
C31 plus.n3 a_n1236_n3888# 0.744346f
C32 plus.t2 a_n1236_n3888# 0.339698f
C33 plus.n4 a_n1236_n3888# 0.158667f
C34 plus.t0 a_n1236_n3888# 0.339698f
C35 plus.t5 a_n1236_n3888# 0.336662f
C36 plus.n5 a_n1236_n3888# 0.137489f
C37 plus.n6 a_n1236_n3888# 0.158587f
C38 plus.n7 a_n1236_n3888# 1.59889f
C39 drain_right.t5 a_n1236_n3888# 3.56524f
C40 drain_right.t1 a_n1236_n3888# 0.43408f
C41 drain_right.t0 a_n1236_n3888# 0.43408f
C42 drain_right.n0 a_n1236_n3888# 2.8851f
C43 drain_right.n1 a_n1236_n3888# 1.75234f
C44 drain_right.t4 a_n1236_n3888# 0.43408f
C45 drain_right.t3 a_n1236_n3888# 0.43408f
C46 drain_right.n2 a_n1236_n3888# 2.88741f
C47 drain_right.t2 a_n1236_n3888# 3.56328f
C48 drain_right.n3 a_n1236_n3888# 0.849098f
C49 source.t0 a_n1236_n3888# 3.19906f
C50 source.n0 a_n1236_n3888# 1.42414f
C51 source.t3 a_n1236_n3888# 0.401766f
C52 source.t5 a_n1236_n3888# 0.401766f
C53 source.n1 a_n1236_n3888# 2.60246f
C54 source.n2 a_n1236_n3888# 0.314803f
C55 source.t6 a_n1236_n3888# 3.19907f
C56 source.n3 a_n1236_n3888# 0.441376f
C57 source.t9 a_n1236_n3888# 0.401766f
C58 source.t10 a_n1236_n3888# 0.401766f
C59 source.n4 a_n1236_n3888# 2.60246f
C60 source.n5 a_n1236_n3888# 1.71037f
C61 source.t2 a_n1236_n3888# 0.401766f
C62 source.t4 a_n1236_n3888# 0.401766f
C63 source.n6 a_n1236_n3888# 2.60246f
C64 source.n7 a_n1236_n3888# 1.71037f
C65 source.t1 a_n1236_n3888# 3.19906f
C66 source.n8 a_n1236_n3888# 0.44138f
C67 source.t11 a_n1236_n3888# 0.401766f
C68 source.t7 a_n1236_n3888# 0.401766f
C69 source.n9 a_n1236_n3888# 2.60246f
C70 source.n10 a_n1236_n3888# 0.314806f
C71 source.t8 a_n1236_n3888# 3.19906f
C72 source.n11 a_n1236_n3888# 0.548458f
C73 source.n12 a_n1236_n3888# 1.63642f
C74 minus.t2 a_n1236_n3888# 0.330443f
C75 minus.n0 a_n1236_n3888# 0.154344f
C76 minus.t3 a_n1236_n3888# 0.330443f
C77 minus.t1 a_n1236_n3888# 0.32749f
C78 minus.n1 a_n1236_n3888# 0.133743f
C79 minus.n2 a_n1236_n3888# 0.154267f
C80 minus.n3 a_n1236_n3888# 1.886f
C81 minus.t0 a_n1236_n3888# 0.330443f
C82 minus.n4 a_n1236_n3888# 0.154344f
C83 minus.t4 a_n1236_n3888# 0.32749f
C84 minus.n5 a_n1236_n3888# 0.133743f
C85 minus.t5 a_n1236_n3888# 0.330443f
C86 minus.n6 a_n1236_n3888# 0.154267f
C87 minus.n7 a_n1236_n3888# 0.40939f
C88 minus.n8 a_n1236_n3888# 2.20927f
.ends

