* NGSPICE file created from diffpair109.ext - technology: sky130A

.subckt diffpair109 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t42 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_left.t22 plus.t1 source.t25 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t21 plus.t2 source.t41 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t35 plus.t3 drain_left.t20 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 drain_left.t19 plus.t4 source.t28 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X5 drain_left.t18 plus.t5 source.t46 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 source.t0 minus.t0 drain_right.t23 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X7 source.t47 plus.t6 drain_left.t17 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X8 drain_left.t16 plus.t7 source.t38 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X9 source.t17 minus.t1 drain_right.t22 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X10 drain_right.t21 minus.t2 source.t22 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X11 source.t27 plus.t8 drain_left.t15 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 drain_left.t14 plus.t9 source.t39 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X13 a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X14 source.t44 plus.t10 drain_left.t13 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X15 source.t40 plus.t11 drain_left.t12 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X16 source.t45 plus.t12 drain_left.t11 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X17 drain_right.t20 minus.t3 source.t21 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X18 source.t18 minus.t4 drain_right.t19 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X19 drain_left.t10 plus.t13 source.t34 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X20 source.t9 minus.t5 drain_right.t18 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X21 drain_right.t17 minus.t6 source.t4 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X22 a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X23 source.t6 minus.t7 drain_right.t16 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X24 source.t10 minus.t8 drain_right.t15 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X25 source.t36 plus.t14 drain_left.t9 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X26 source.t26 plus.t15 drain_left.t8 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X27 source.t24 plus.t16 drain_left.t7 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X28 source.t13 minus.t9 drain_right.t14 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X29 source.t1 minus.t10 drain_right.t13 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X30 source.t2 minus.t11 drain_right.t12 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X31 source.t29 plus.t17 drain_left.t6 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X32 drain_right.t11 minus.t12 source.t5 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X33 source.t33 plus.t18 drain_left.t5 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X34 drain_right.t10 minus.t13 source.t3 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X35 drain_right.t9 minus.t14 source.t20 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X36 source.t11 minus.t15 drain_right.t8 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X37 source.t15 minus.t16 drain_right.t7 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X38 a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X39 a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X40 drain_right.t6 minus.t17 source.t8 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X41 drain_right.t5 minus.t18 source.t19 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X42 source.t43 plus.t19 drain_left.t4 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X43 drain_right.t4 minus.t19 source.t23 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X44 drain_right.t3 minus.t20 source.t14 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X45 drain_right.t2 minus.t21 source.t16 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X46 drain_right.t1 minus.t22 source.t7 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X47 drain_left.t3 plus.t20 source.t30 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X48 source.t12 minus.t23 drain_right.t0 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X49 drain_left.t2 plus.t21 source.t37 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X50 drain_left.t1 plus.t22 source.t32 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X51 drain_left.t0 plus.t23 source.t31 a_n2224_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
R0 plus.n6 plus.t11 345.872
R1 plus.n33 plus.t4 345.872
R2 plus.n42 plus.t21 345.872
R3 plus.n68 plus.t6 345.872
R4 plus.n7 plus.t1 318.12
R5 plus.n8 plus.t16 318.12
R6 plus.n14 plus.t0 318.12
R7 plus.n16 plus.t15 318.12
R8 plus.n3 plus.t22 318.12
R9 plus.n21 plus.t14 318.12
R10 plus.n23 plus.t7 318.12
R11 plus.n24 plus.t18 318.12
R12 plus.n30 plus.t5 318.12
R13 plus.n32 plus.t17 318.12
R14 plus.n44 plus.t19 318.12
R15 plus.n43 plus.t2 318.12
R16 plus.n50 plus.t10 318.12
R17 plus.n52 plus.t20 318.12
R18 plus.n39 plus.t3 318.12
R19 plus.n57 plus.t23 318.12
R20 plus.n59 plus.t8 318.12
R21 plus.n38 plus.t13 318.12
R22 plus.n65 plus.t12 318.12
R23 plus.n67 plus.t9 318.12
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus.n17 plus.n3 30.6732
R75 plus.n22 plus.n21 30.6732
R76 plus.n58 plus.n57 30.6732
R77 plus.n53 plus.n39 30.6732
R78 plus plus.n69 27.571
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 8.28838
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n98 source.n96 289.615
R119 source.n80 source.n78 289.615
R120 source.n72 source.n70 289.615
R121 source.n54 source.n52 289.615
R122 source.n2 source.n0 289.615
R123 source.n20 source.n18 289.615
R124 source.n28 source.n26 289.615
R125 source.n46 source.n44 289.615
R126 source.n99 source.n98 185
R127 source.n81 source.n80 185
R128 source.n73 source.n72 185
R129 source.n55 source.n54 185
R130 source.n3 source.n2 185
R131 source.n21 source.n20 185
R132 source.n29 source.n28 185
R133 source.n47 source.n46 185
R134 source.t16 source.n97 167.117
R135 source.t2 source.n79 167.117
R136 source.t37 source.n71 167.117
R137 source.t47 source.n53 167.117
R138 source.t28 source.n1 167.117
R139 source.t40 source.n19 167.117
R140 source.t3 source.n27 167.117
R141 source.t15 source.n45 167.117
R142 source.n9 source.n8 84.1169
R143 source.n11 source.n10 84.1169
R144 source.n13 source.n12 84.1169
R145 source.n15 source.n14 84.1169
R146 source.n17 source.n16 84.1169
R147 source.n35 source.n34 84.1169
R148 source.n37 source.n36 84.1169
R149 source.n39 source.n38 84.1169
R150 source.n41 source.n40 84.1169
R151 source.n43 source.n42 84.1169
R152 source.n95 source.n94 84.1168
R153 source.n93 source.n92 84.1168
R154 source.n91 source.n90 84.1168
R155 source.n89 source.n88 84.1168
R156 source.n87 source.n86 84.1168
R157 source.n69 source.n68 84.1168
R158 source.n67 source.n66 84.1168
R159 source.n65 source.n64 84.1168
R160 source.n63 source.n62 84.1168
R161 source.n61 source.n60 84.1168
R162 source.n98 source.t16 52.3082
R163 source.n80 source.t2 52.3082
R164 source.n72 source.t37 52.3082
R165 source.n54 source.t47 52.3082
R166 source.n2 source.t28 52.3082
R167 source.n20 source.t40 52.3082
R168 source.n28 source.t3 52.3082
R169 source.n46 source.t15 52.3082
R170 source.n103 source.n102 31.4096
R171 source.n85 source.n84 31.4096
R172 source.n77 source.n76 31.4096
R173 source.n59 source.n58 31.4096
R174 source.n7 source.n6 31.4096
R175 source.n25 source.n24 31.4096
R176 source.n33 source.n32 31.4096
R177 source.n51 source.n50 31.4096
R178 source.n59 source.n51 14.212
R179 source.n94 source.t8 9.9005
R180 source.n94 source.t12 9.9005
R181 source.n92 source.t20 9.9005
R182 source.n92 source.t13 9.9005
R183 source.n90 source.t19 9.9005
R184 source.n90 source.t11 9.9005
R185 source.n88 source.t4 9.9005
R186 source.n88 source.t1 9.9005
R187 source.n86 source.t21 9.9005
R188 source.n86 source.t10 9.9005
R189 source.n68 source.t41 9.9005
R190 source.n68 source.t43 9.9005
R191 source.n66 source.t30 9.9005
R192 source.n66 source.t44 9.9005
R193 source.n64 source.t31 9.9005
R194 source.n64 source.t35 9.9005
R195 source.n62 source.t34 9.9005
R196 source.n62 source.t27 9.9005
R197 source.n60 source.t39 9.9005
R198 source.n60 source.t45 9.9005
R199 source.n8 source.t46 9.9005
R200 source.n8 source.t29 9.9005
R201 source.n10 source.t38 9.9005
R202 source.n10 source.t33 9.9005
R203 source.n12 source.t32 9.9005
R204 source.n12 source.t36 9.9005
R205 source.n14 source.t42 9.9005
R206 source.n14 source.t26 9.9005
R207 source.n16 source.t25 9.9005
R208 source.n16 source.t24 9.9005
R209 source.n34 source.t5 9.9005
R210 source.n34 source.t17 9.9005
R211 source.n36 source.t23 9.9005
R212 source.n36 source.t0 9.9005
R213 source.n38 source.t14 9.9005
R214 source.n38 source.t9 9.9005
R215 source.n40 source.t7 9.9005
R216 source.n40 source.t18 9.9005
R217 source.n42 source.t22 9.9005
R218 source.n42 source.t6 9.9005
R219 source.n99 source.n97 9.71174
R220 source.n81 source.n79 9.71174
R221 source.n73 source.n71 9.71174
R222 source.n55 source.n53 9.71174
R223 source.n3 source.n1 9.71174
R224 source.n21 source.n19 9.71174
R225 source.n29 source.n27 9.71174
R226 source.n47 source.n45 9.71174
R227 source.n102 source.n101 9.45567
R228 source.n84 source.n83 9.45567
R229 source.n76 source.n75 9.45567
R230 source.n58 source.n57 9.45567
R231 source.n6 source.n5 9.45567
R232 source.n24 source.n23 9.45567
R233 source.n32 source.n31 9.45567
R234 source.n50 source.n49 9.45567
R235 source.n101 source.n100 9.3005
R236 source.n83 source.n82 9.3005
R237 source.n75 source.n74 9.3005
R238 source.n57 source.n56 9.3005
R239 source.n5 source.n4 9.3005
R240 source.n23 source.n22 9.3005
R241 source.n31 source.n30 9.3005
R242 source.n49 source.n48 9.3005
R243 source.n104 source.n7 8.69904
R244 source.n102 source.n96 8.14595
R245 source.n84 source.n78 8.14595
R246 source.n76 source.n70 8.14595
R247 source.n58 source.n52 8.14595
R248 source.n6 source.n0 8.14595
R249 source.n24 source.n18 8.14595
R250 source.n32 source.n26 8.14595
R251 source.n50 source.n44 8.14595
R252 source.n100 source.n99 7.3702
R253 source.n82 source.n81 7.3702
R254 source.n74 source.n73 7.3702
R255 source.n56 source.n55 7.3702
R256 source.n4 source.n3 7.3702
R257 source.n22 source.n21 7.3702
R258 source.n30 source.n29 7.3702
R259 source.n48 source.n47 7.3702
R260 source.n100 source.n96 5.81868
R261 source.n82 source.n78 5.81868
R262 source.n74 source.n70 5.81868
R263 source.n56 source.n52 5.81868
R264 source.n4 source.n0 5.81868
R265 source.n22 source.n18 5.81868
R266 source.n30 source.n26 5.81868
R267 source.n48 source.n44 5.81868
R268 source.n104 source.n103 5.51343
R269 source.n101 source.n97 3.44771
R270 source.n83 source.n79 3.44771
R271 source.n75 source.n71 3.44771
R272 source.n57 source.n53 3.44771
R273 source.n5 source.n1 3.44771
R274 source.n23 source.n19 3.44771
R275 source.n31 source.n27 3.44771
R276 source.n49 source.n45 3.44771
R277 source.n51 source.n43 0.5005
R278 source.n43 source.n41 0.5005
R279 source.n41 source.n39 0.5005
R280 source.n39 source.n37 0.5005
R281 source.n37 source.n35 0.5005
R282 source.n35 source.n33 0.5005
R283 source.n25 source.n17 0.5005
R284 source.n17 source.n15 0.5005
R285 source.n15 source.n13 0.5005
R286 source.n13 source.n11 0.5005
R287 source.n11 source.n9 0.5005
R288 source.n9 source.n7 0.5005
R289 source.n61 source.n59 0.5005
R290 source.n63 source.n61 0.5005
R291 source.n65 source.n63 0.5005
R292 source.n67 source.n65 0.5005
R293 source.n69 source.n67 0.5005
R294 source.n77 source.n69 0.5005
R295 source.n87 source.n85 0.5005
R296 source.n89 source.n87 0.5005
R297 source.n91 source.n89 0.5005
R298 source.n93 source.n91 0.5005
R299 source.n95 source.n93 0.5005
R300 source.n103 source.n95 0.5005
R301 source.n33 source.n25 0.470328
R302 source.n85 source.n77 0.470328
R303 source source.n104 0.188
R304 drain_left.n13 drain_left.n11 101.296
R305 drain_left.n7 drain_left.n5 101.296
R306 drain_left.n2 drain_left.n0 101.296
R307 drain_left.n21 drain_left.n20 100.796
R308 drain_left.n19 drain_left.n18 100.796
R309 drain_left.n17 drain_left.n16 100.796
R310 drain_left.n15 drain_left.n14 100.796
R311 drain_left.n13 drain_left.n12 100.796
R312 drain_left.n7 drain_left.n6 100.796
R313 drain_left.n9 drain_left.n8 100.796
R314 drain_left.n4 drain_left.n3 100.796
R315 drain_left.n2 drain_left.n1 100.796
R316 drain_left drain_left.n10 24.5413
R317 drain_left.n5 drain_left.t4 9.9005
R318 drain_left.n5 drain_left.t2 9.9005
R319 drain_left.n6 drain_left.t13 9.9005
R320 drain_left.n6 drain_left.t21 9.9005
R321 drain_left.n8 drain_left.t20 9.9005
R322 drain_left.n8 drain_left.t3 9.9005
R323 drain_left.n3 drain_left.t15 9.9005
R324 drain_left.n3 drain_left.t0 9.9005
R325 drain_left.n1 drain_left.t11 9.9005
R326 drain_left.n1 drain_left.t10 9.9005
R327 drain_left.n0 drain_left.t17 9.9005
R328 drain_left.n0 drain_left.t14 9.9005
R329 drain_left.n20 drain_left.t6 9.9005
R330 drain_left.n20 drain_left.t19 9.9005
R331 drain_left.n18 drain_left.t5 9.9005
R332 drain_left.n18 drain_left.t18 9.9005
R333 drain_left.n16 drain_left.t9 9.9005
R334 drain_left.n16 drain_left.t16 9.9005
R335 drain_left.n14 drain_left.t8 9.9005
R336 drain_left.n14 drain_left.t1 9.9005
R337 drain_left.n12 drain_left.t7 9.9005
R338 drain_left.n12 drain_left.t23 9.9005
R339 drain_left.n11 drain_left.t12 9.9005
R340 drain_left.n11 drain_left.t22 9.9005
R341 drain_left drain_left.n21 6.15322
R342 drain_left.n9 drain_left.n7 0.5005
R343 drain_left.n4 drain_left.n2 0.5005
R344 drain_left.n15 drain_left.n13 0.5005
R345 drain_left.n17 drain_left.n15 0.5005
R346 drain_left.n19 drain_left.n17 0.5005
R347 drain_left.n21 drain_left.n19 0.5005
R348 drain_left.n10 drain_left.n9 0.195154
R349 drain_left.n10 drain_left.n4 0.195154
R350 minus.n33 minus.t16 345.872
R351 minus.n7 minus.t13 345.872
R352 minus.n68 minus.t21 345.872
R353 minus.n41 minus.t11 345.872
R354 minus.n32 minus.t2 318.12
R355 minus.n30 minus.t7 318.12
R356 minus.n3 minus.t22 318.12
R357 minus.n24 minus.t4 318.12
R358 minus.n22 minus.t20 318.12
R359 minus.n4 minus.t5 318.12
R360 minus.n17 minus.t19 318.12
R361 minus.n15 minus.t0 318.12
R362 minus.n8 minus.t12 318.12
R363 minus.n9 minus.t1 318.12
R364 minus.n67 minus.t23 318.12
R365 minus.n65 minus.t17 318.12
R366 minus.n59 minus.t9 318.12
R367 minus.n58 minus.t14 318.12
R368 minus.n56 minus.t15 318.12
R369 minus.n38 minus.t18 318.12
R370 minus.n51 minus.t10 318.12
R371 minus.n49 minus.t6 318.12
R372 minus.n43 minus.t8 318.12
R373 minus.n42 minus.t3 318.12
R374 minus.n11 minus.n7 161.489
R375 minus.n45 minus.n41 161.489
R376 minus.n34 minus.n33 161.3
R377 minus.n31 minus.n0 161.3
R378 minus.n29 minus.n28 161.3
R379 minus.n27 minus.n1 161.3
R380 minus.n26 minus.n25 161.3
R381 minus.n23 minus.n2 161.3
R382 minus.n21 minus.n20 161.3
R383 minus.n19 minus.n18 161.3
R384 minus.n16 minus.n5 161.3
R385 minus.n14 minus.n13 161.3
R386 minus.n12 minus.n6 161.3
R387 minus.n11 minus.n10 161.3
R388 minus.n69 minus.n68 161.3
R389 minus.n66 minus.n35 161.3
R390 minus.n64 minus.n63 161.3
R391 minus.n62 minus.n36 161.3
R392 minus.n61 minus.n60 161.3
R393 minus.n57 minus.n37 161.3
R394 minus.n55 minus.n54 161.3
R395 minus.n53 minus.n52 161.3
R396 minus.n50 minus.n39 161.3
R397 minus.n48 minus.n47 161.3
R398 minus.n46 minus.n40 161.3
R399 minus.n45 minus.n44 161.3
R400 minus.n29 minus.n1 73.0308
R401 minus.n14 minus.n6 73.0308
R402 minus.n48 minus.n40 73.0308
R403 minus.n64 minus.n36 73.0308
R404 minus.n31 minus.n30 68.649
R405 minus.n10 minus.n8 68.649
R406 minus.n44 minus.n43 68.649
R407 minus.n66 minus.n65 68.649
R408 minus.n25 minus.n3 65.7278
R409 minus.n16 minus.n15 65.7278
R410 minus.n50 minus.n49 65.7278
R411 minus.n60 minus.n59 65.7278
R412 minus.n33 minus.n32 56.9641
R413 minus.n9 minus.n7 56.9641
R414 minus.n42 minus.n41 56.9641
R415 minus.n68 minus.n67 56.9641
R416 minus.n24 minus.n23 54.0429
R417 minus.n18 minus.n17 54.0429
R418 minus.n52 minus.n51 54.0429
R419 minus.n58 minus.n57 54.0429
R420 minus.n22 minus.n21 42.3581
R421 minus.n21 minus.n4 42.3581
R422 minus.n55 minus.n38 42.3581
R423 minus.n56 minus.n55 42.3581
R424 minus.n23 minus.n22 30.6732
R425 minus.n18 minus.n4 30.6732
R426 minus.n52 minus.n38 30.6732
R427 minus.n57 minus.n56 30.6732
R428 minus.n70 minus.n34 29.902
R429 minus.n25 minus.n24 18.9884
R430 minus.n17 minus.n16 18.9884
R431 minus.n51 minus.n50 18.9884
R432 minus.n60 minus.n58 18.9884
R433 minus.n32 minus.n31 16.0672
R434 minus.n10 minus.n9 16.0672
R435 minus.n44 minus.n42 16.0672
R436 minus.n67 minus.n66 16.0672
R437 minus.n3 minus.n1 7.30353
R438 minus.n15 minus.n14 7.30353
R439 minus.n49 minus.n48 7.30353
R440 minus.n59 minus.n36 7.30353
R441 minus.n70 minus.n69 6.43232
R442 minus.n30 minus.n29 4.38232
R443 minus.n8 minus.n6 4.38232
R444 minus.n43 minus.n40 4.38232
R445 minus.n65 minus.n64 4.38232
R446 minus.n34 minus.n0 0.189894
R447 minus.n28 minus.n0 0.189894
R448 minus.n28 minus.n27 0.189894
R449 minus.n27 minus.n26 0.189894
R450 minus.n26 minus.n2 0.189894
R451 minus.n20 minus.n2 0.189894
R452 minus.n20 minus.n19 0.189894
R453 minus.n19 minus.n5 0.189894
R454 minus.n13 minus.n5 0.189894
R455 minus.n13 minus.n12 0.189894
R456 minus.n12 minus.n11 0.189894
R457 minus.n46 minus.n45 0.189894
R458 minus.n47 minus.n46 0.189894
R459 minus.n47 minus.n39 0.189894
R460 minus.n53 minus.n39 0.189894
R461 minus.n54 minus.n53 0.189894
R462 minus.n54 minus.n37 0.189894
R463 minus.n61 minus.n37 0.189894
R464 minus.n62 minus.n61 0.189894
R465 minus.n63 minus.n62 0.189894
R466 minus.n63 minus.n35 0.189894
R467 minus.n69 minus.n35 0.189894
R468 minus minus.n70 0.188
R469 drain_right.n13 drain_right.n11 101.296
R470 drain_right.n7 drain_right.n5 101.296
R471 drain_right.n2 drain_right.n0 101.296
R472 drain_right.n13 drain_right.n12 100.796
R473 drain_right.n15 drain_right.n14 100.796
R474 drain_right.n17 drain_right.n16 100.796
R475 drain_right.n19 drain_right.n18 100.796
R476 drain_right.n21 drain_right.n20 100.796
R477 drain_right.n7 drain_right.n6 100.796
R478 drain_right.n9 drain_right.n8 100.796
R479 drain_right.n4 drain_right.n3 100.796
R480 drain_right.n2 drain_right.n1 100.796
R481 drain_right drain_right.n10 23.9881
R482 drain_right.n5 drain_right.t0 9.9005
R483 drain_right.n5 drain_right.t2 9.9005
R484 drain_right.n6 drain_right.t14 9.9005
R485 drain_right.n6 drain_right.t6 9.9005
R486 drain_right.n8 drain_right.t8 9.9005
R487 drain_right.n8 drain_right.t9 9.9005
R488 drain_right.n3 drain_right.t13 9.9005
R489 drain_right.n3 drain_right.t5 9.9005
R490 drain_right.n1 drain_right.t15 9.9005
R491 drain_right.n1 drain_right.t17 9.9005
R492 drain_right.n0 drain_right.t12 9.9005
R493 drain_right.n0 drain_right.t20 9.9005
R494 drain_right.n11 drain_right.t22 9.9005
R495 drain_right.n11 drain_right.t10 9.9005
R496 drain_right.n12 drain_right.t23 9.9005
R497 drain_right.n12 drain_right.t11 9.9005
R498 drain_right.n14 drain_right.t18 9.9005
R499 drain_right.n14 drain_right.t4 9.9005
R500 drain_right.n16 drain_right.t19 9.9005
R501 drain_right.n16 drain_right.t3 9.9005
R502 drain_right.n18 drain_right.t16 9.9005
R503 drain_right.n18 drain_right.t1 9.9005
R504 drain_right.n20 drain_right.t7 9.9005
R505 drain_right.n20 drain_right.t21 9.9005
R506 drain_right drain_right.n21 6.15322
R507 drain_right.n9 drain_right.n7 0.5005
R508 drain_right.n4 drain_right.n2 0.5005
R509 drain_right.n21 drain_right.n19 0.5005
R510 drain_right.n19 drain_right.n17 0.5005
R511 drain_right.n17 drain_right.n15 0.5005
R512 drain_right.n15 drain_right.n13 0.5005
R513 drain_right.n10 drain_right.n9 0.195154
R514 drain_right.n10 drain_right.n4 0.195154
C0 drain_left minus 0.178374f
C1 source plus 2.06795f
C2 plus minus 4.09048f
C3 drain_left plus 1.99342f
C4 drain_right source 11.197701f
C5 drain_right minus 1.77479f
C6 drain_right drain_left 1.19771f
C7 drain_right plus 0.380894f
C8 source minus 2.05399f
C9 drain_left source 11.1973f
C10 drain_right a_n2224_n1288# 4.66756f
C11 drain_left a_n2224_n1288# 4.97523f
C12 source a_n2224_n1288# 3.322397f
C13 minus a_n2224_n1288# 7.920766f
C14 plus a_n2224_n1288# 8.934879f
C15 drain_right.t12 a_n2224_n1288# 0.046161f
C16 drain_right.t20 a_n2224_n1288# 0.046161f
C17 drain_right.n0 a_n2224_n1288# 0.291625f
C18 drain_right.t15 a_n2224_n1288# 0.046161f
C19 drain_right.t17 a_n2224_n1288# 0.046161f
C20 drain_right.n1 a_n2224_n1288# 0.289999f
C21 drain_right.n2 a_n2224_n1288# 0.645467f
C22 drain_right.t13 a_n2224_n1288# 0.046161f
C23 drain_right.t5 a_n2224_n1288# 0.046161f
C24 drain_right.n3 a_n2224_n1288# 0.289999f
C25 drain_right.n4 a_n2224_n1288# 0.292406f
C26 drain_right.t0 a_n2224_n1288# 0.046161f
C27 drain_right.t2 a_n2224_n1288# 0.046161f
C28 drain_right.n5 a_n2224_n1288# 0.291625f
C29 drain_right.t14 a_n2224_n1288# 0.046161f
C30 drain_right.t6 a_n2224_n1288# 0.046161f
C31 drain_right.n6 a_n2224_n1288# 0.289999f
C32 drain_right.n7 a_n2224_n1288# 0.645467f
C33 drain_right.t8 a_n2224_n1288# 0.046161f
C34 drain_right.t9 a_n2224_n1288# 0.046161f
C35 drain_right.n8 a_n2224_n1288# 0.289999f
C36 drain_right.n9 a_n2224_n1288# 0.292406f
C37 drain_right.n10 a_n2224_n1288# 0.8814f
C38 drain_right.t22 a_n2224_n1288# 0.046161f
C39 drain_right.t10 a_n2224_n1288# 0.046161f
C40 drain_right.n11 a_n2224_n1288# 0.291626f
C41 drain_right.t23 a_n2224_n1288# 0.046161f
C42 drain_right.t11 a_n2224_n1288# 0.046161f
C43 drain_right.n12 a_n2224_n1288# 0.29f
C44 drain_right.n13 a_n2224_n1288# 0.645464f
C45 drain_right.t18 a_n2224_n1288# 0.046161f
C46 drain_right.t4 a_n2224_n1288# 0.046161f
C47 drain_right.n14 a_n2224_n1288# 0.29f
C48 drain_right.n15 a_n2224_n1288# 0.317663f
C49 drain_right.t19 a_n2224_n1288# 0.046161f
C50 drain_right.t3 a_n2224_n1288# 0.046161f
C51 drain_right.n16 a_n2224_n1288# 0.29f
C52 drain_right.n17 a_n2224_n1288# 0.317663f
C53 drain_right.t16 a_n2224_n1288# 0.046161f
C54 drain_right.t1 a_n2224_n1288# 0.046161f
C55 drain_right.n18 a_n2224_n1288# 0.29f
C56 drain_right.n19 a_n2224_n1288# 0.317663f
C57 drain_right.t7 a_n2224_n1288# 0.046161f
C58 drain_right.t21 a_n2224_n1288# 0.046161f
C59 drain_right.n20 a_n2224_n1288# 0.29f
C60 drain_right.n21 a_n2224_n1288# 0.558751f
C61 minus.n0 a_n2224_n1288# 0.038825f
C62 minus.t16 a_n2224_n1288# 0.060369f
C63 minus.t2 a_n2224_n1288# 0.057123f
C64 minus.t7 a_n2224_n1288# 0.057123f
C65 minus.n1 a_n2224_n1288# 0.014076f
C66 minus.n2 a_n2224_n1288# 0.038825f
C67 minus.t22 a_n2224_n1288# 0.057123f
C68 minus.n3 a_n2224_n1288# 0.04189f
C69 minus.t4 a_n2224_n1288# 0.057123f
C70 minus.t20 a_n2224_n1288# 0.057123f
C71 minus.t5 a_n2224_n1288# 0.057123f
C72 minus.n4 a_n2224_n1288# 0.04189f
C73 minus.n5 a_n2224_n1288# 0.038825f
C74 minus.t19 a_n2224_n1288# 0.057123f
C75 minus.t0 a_n2224_n1288# 0.057123f
C76 minus.n6 a_n2224_n1288# 0.013598f
C77 minus.t13 a_n2224_n1288# 0.060369f
C78 minus.n7 a_n2224_n1288# 0.052052f
C79 minus.t12 a_n2224_n1288# 0.057123f
C80 minus.n8 a_n2224_n1288# 0.04189f
C81 minus.t1 a_n2224_n1288# 0.057123f
C82 minus.n9 a_n2224_n1288# 0.04189f
C83 minus.n10 a_n2224_n1288# 0.014795f
C84 minus.n11 a_n2224_n1288# 0.080713f
C85 minus.n12 a_n2224_n1288# 0.038825f
C86 minus.n13 a_n2224_n1288# 0.038825f
C87 minus.n14 a_n2224_n1288# 0.014076f
C88 minus.n15 a_n2224_n1288# 0.04189f
C89 minus.n16 a_n2224_n1288# 0.014795f
C90 minus.n17 a_n2224_n1288# 0.04189f
C91 minus.n18 a_n2224_n1288# 0.014795f
C92 minus.n19 a_n2224_n1288# 0.038825f
C93 minus.n20 a_n2224_n1288# 0.038825f
C94 minus.n21 a_n2224_n1288# 0.014795f
C95 minus.n22 a_n2224_n1288# 0.04189f
C96 minus.n23 a_n2224_n1288# 0.014795f
C97 minus.n24 a_n2224_n1288# 0.04189f
C98 minus.n25 a_n2224_n1288# 0.014795f
C99 minus.n26 a_n2224_n1288# 0.038825f
C100 minus.n27 a_n2224_n1288# 0.038825f
C101 minus.n28 a_n2224_n1288# 0.038825f
C102 minus.n29 a_n2224_n1288# 0.013598f
C103 minus.n30 a_n2224_n1288# 0.04189f
C104 minus.n31 a_n2224_n1288# 0.014795f
C105 minus.n32 a_n2224_n1288# 0.04189f
C106 minus.n33 a_n2224_n1288# 0.052003f
C107 minus.n34 a_n2224_n1288# 1.00192f
C108 minus.n35 a_n2224_n1288# 0.038825f
C109 minus.t23 a_n2224_n1288# 0.057123f
C110 minus.t17 a_n2224_n1288# 0.057123f
C111 minus.n36 a_n2224_n1288# 0.014076f
C112 minus.n37 a_n2224_n1288# 0.038825f
C113 minus.t14 a_n2224_n1288# 0.057123f
C114 minus.t15 a_n2224_n1288# 0.057123f
C115 minus.t18 a_n2224_n1288# 0.057123f
C116 minus.n38 a_n2224_n1288# 0.04189f
C117 minus.n39 a_n2224_n1288# 0.038825f
C118 minus.t10 a_n2224_n1288# 0.057123f
C119 minus.t6 a_n2224_n1288# 0.057123f
C120 minus.n40 a_n2224_n1288# 0.013598f
C121 minus.t11 a_n2224_n1288# 0.060369f
C122 minus.n41 a_n2224_n1288# 0.052052f
C123 minus.t3 a_n2224_n1288# 0.057123f
C124 minus.n42 a_n2224_n1288# 0.04189f
C125 minus.t8 a_n2224_n1288# 0.057123f
C126 minus.n43 a_n2224_n1288# 0.04189f
C127 minus.n44 a_n2224_n1288# 0.014795f
C128 minus.n45 a_n2224_n1288# 0.080713f
C129 minus.n46 a_n2224_n1288# 0.038825f
C130 minus.n47 a_n2224_n1288# 0.038825f
C131 minus.n48 a_n2224_n1288# 0.014076f
C132 minus.n49 a_n2224_n1288# 0.04189f
C133 minus.n50 a_n2224_n1288# 0.014795f
C134 minus.n51 a_n2224_n1288# 0.04189f
C135 minus.n52 a_n2224_n1288# 0.014795f
C136 minus.n53 a_n2224_n1288# 0.038825f
C137 minus.n54 a_n2224_n1288# 0.038825f
C138 minus.n55 a_n2224_n1288# 0.014795f
C139 minus.n56 a_n2224_n1288# 0.04189f
C140 minus.n57 a_n2224_n1288# 0.014795f
C141 minus.n58 a_n2224_n1288# 0.04189f
C142 minus.t9 a_n2224_n1288# 0.057123f
C143 minus.n59 a_n2224_n1288# 0.04189f
C144 minus.n60 a_n2224_n1288# 0.014795f
C145 minus.n61 a_n2224_n1288# 0.038825f
C146 minus.n62 a_n2224_n1288# 0.038825f
C147 minus.n63 a_n2224_n1288# 0.038825f
C148 minus.n64 a_n2224_n1288# 0.013598f
C149 minus.n65 a_n2224_n1288# 0.04189f
C150 minus.n66 a_n2224_n1288# 0.014795f
C151 minus.n67 a_n2224_n1288# 0.04189f
C152 minus.t21 a_n2224_n1288# 0.060369f
C153 minus.n68 a_n2224_n1288# 0.052003f
C154 minus.n69 a_n2224_n1288# 0.247617f
C155 minus.n70 a_n2224_n1288# 1.23938f
C156 drain_left.t17 a_n2224_n1288# 0.045695f
C157 drain_left.t14 a_n2224_n1288# 0.045695f
C158 drain_left.n0 a_n2224_n1288# 0.28868f
C159 drain_left.t11 a_n2224_n1288# 0.045695f
C160 drain_left.t10 a_n2224_n1288# 0.045695f
C161 drain_left.n1 a_n2224_n1288# 0.287071f
C162 drain_left.n2 a_n2224_n1288# 0.638949f
C163 drain_left.t15 a_n2224_n1288# 0.045695f
C164 drain_left.t0 a_n2224_n1288# 0.045695f
C165 drain_left.n3 a_n2224_n1288# 0.287071f
C166 drain_left.n4 a_n2224_n1288# 0.289453f
C167 drain_left.t4 a_n2224_n1288# 0.045695f
C168 drain_left.t2 a_n2224_n1288# 0.045695f
C169 drain_left.n5 a_n2224_n1288# 0.28868f
C170 drain_left.t13 a_n2224_n1288# 0.045695f
C171 drain_left.t21 a_n2224_n1288# 0.045695f
C172 drain_left.n6 a_n2224_n1288# 0.287071f
C173 drain_left.n7 a_n2224_n1288# 0.638949f
C174 drain_left.t20 a_n2224_n1288# 0.045695f
C175 drain_left.t3 a_n2224_n1288# 0.045695f
C176 drain_left.n8 a_n2224_n1288# 0.287071f
C177 drain_left.n9 a_n2224_n1288# 0.289453f
C178 drain_left.n10 a_n2224_n1288# 0.928922f
C179 drain_left.t12 a_n2224_n1288# 0.045695f
C180 drain_left.t22 a_n2224_n1288# 0.045695f
C181 drain_left.n11 a_n2224_n1288# 0.288682f
C182 drain_left.t7 a_n2224_n1288# 0.045695f
C183 drain_left.t23 a_n2224_n1288# 0.045695f
C184 drain_left.n12 a_n2224_n1288# 0.287072f
C185 drain_left.n13 a_n2224_n1288# 0.638946f
C186 drain_left.t8 a_n2224_n1288# 0.045695f
C187 drain_left.t1 a_n2224_n1288# 0.045695f
C188 drain_left.n14 a_n2224_n1288# 0.287072f
C189 drain_left.n15 a_n2224_n1288# 0.314455f
C190 drain_left.t9 a_n2224_n1288# 0.045695f
C191 drain_left.t16 a_n2224_n1288# 0.045695f
C192 drain_left.n16 a_n2224_n1288# 0.287072f
C193 drain_left.n17 a_n2224_n1288# 0.314455f
C194 drain_left.t5 a_n2224_n1288# 0.045695f
C195 drain_left.t18 a_n2224_n1288# 0.045695f
C196 drain_left.n18 a_n2224_n1288# 0.287072f
C197 drain_left.n19 a_n2224_n1288# 0.314455f
C198 drain_left.t6 a_n2224_n1288# 0.045695f
C199 drain_left.t19 a_n2224_n1288# 0.045695f
C200 drain_left.n20 a_n2224_n1288# 0.287072f
C201 drain_left.n21 a_n2224_n1288# 0.553108f
C202 source.n0 a_n2224_n1288# 0.053582f
C203 source.n1 a_n2224_n1288# 0.118556f
C204 source.t28 a_n2224_n1288# 0.08897f
C205 source.n2 a_n2224_n1288# 0.092786f
C206 source.n3 a_n2224_n1288# 0.029911f
C207 source.n4 a_n2224_n1288# 0.019727f
C208 source.n5 a_n2224_n1288# 0.261326f
C209 source.n6 a_n2224_n1288# 0.058738f
C210 source.n7 a_n2224_n1288# 0.545208f
C211 source.t46 a_n2224_n1288# 0.05802f
C212 source.t29 a_n2224_n1288# 0.05802f
C213 source.n8 a_n2224_n1288# 0.310173f
C214 source.n9 a_n2224_n1288# 0.403699f
C215 source.t38 a_n2224_n1288# 0.05802f
C216 source.t33 a_n2224_n1288# 0.05802f
C217 source.n10 a_n2224_n1288# 0.310173f
C218 source.n11 a_n2224_n1288# 0.403699f
C219 source.t32 a_n2224_n1288# 0.05802f
C220 source.t36 a_n2224_n1288# 0.05802f
C221 source.n12 a_n2224_n1288# 0.310173f
C222 source.n13 a_n2224_n1288# 0.403699f
C223 source.t42 a_n2224_n1288# 0.05802f
C224 source.t26 a_n2224_n1288# 0.05802f
C225 source.n14 a_n2224_n1288# 0.310173f
C226 source.n15 a_n2224_n1288# 0.403699f
C227 source.t25 a_n2224_n1288# 0.05802f
C228 source.t24 a_n2224_n1288# 0.05802f
C229 source.n16 a_n2224_n1288# 0.310173f
C230 source.n17 a_n2224_n1288# 0.403699f
C231 source.n18 a_n2224_n1288# 0.053582f
C232 source.n19 a_n2224_n1288# 0.118556f
C233 source.t40 a_n2224_n1288# 0.08897f
C234 source.n20 a_n2224_n1288# 0.092786f
C235 source.n21 a_n2224_n1288# 0.029911f
C236 source.n22 a_n2224_n1288# 0.019727f
C237 source.n23 a_n2224_n1288# 0.261326f
C238 source.n24 a_n2224_n1288# 0.058738f
C239 source.n25 a_n2224_n1288# 0.144943f
C240 source.n26 a_n2224_n1288# 0.053582f
C241 source.n27 a_n2224_n1288# 0.118556f
C242 source.t3 a_n2224_n1288# 0.08897f
C243 source.n28 a_n2224_n1288# 0.092786f
C244 source.n29 a_n2224_n1288# 0.029911f
C245 source.n30 a_n2224_n1288# 0.019727f
C246 source.n31 a_n2224_n1288# 0.261326f
C247 source.n32 a_n2224_n1288# 0.058738f
C248 source.n33 a_n2224_n1288# 0.144943f
C249 source.t5 a_n2224_n1288# 0.05802f
C250 source.t17 a_n2224_n1288# 0.05802f
C251 source.n34 a_n2224_n1288# 0.310173f
C252 source.n35 a_n2224_n1288# 0.403699f
C253 source.t23 a_n2224_n1288# 0.05802f
C254 source.t0 a_n2224_n1288# 0.05802f
C255 source.n36 a_n2224_n1288# 0.310173f
C256 source.n37 a_n2224_n1288# 0.403699f
C257 source.t14 a_n2224_n1288# 0.05802f
C258 source.t9 a_n2224_n1288# 0.05802f
C259 source.n38 a_n2224_n1288# 0.310173f
C260 source.n39 a_n2224_n1288# 0.403699f
C261 source.t7 a_n2224_n1288# 0.05802f
C262 source.t18 a_n2224_n1288# 0.05802f
C263 source.n40 a_n2224_n1288# 0.310173f
C264 source.n41 a_n2224_n1288# 0.403699f
C265 source.t22 a_n2224_n1288# 0.05802f
C266 source.t6 a_n2224_n1288# 0.05802f
C267 source.n42 a_n2224_n1288# 0.310173f
C268 source.n43 a_n2224_n1288# 0.403699f
C269 source.n44 a_n2224_n1288# 0.053582f
C270 source.n45 a_n2224_n1288# 0.118556f
C271 source.t15 a_n2224_n1288# 0.08897f
C272 source.n46 a_n2224_n1288# 0.092786f
C273 source.n47 a_n2224_n1288# 0.029911f
C274 source.n48 a_n2224_n1288# 0.019727f
C275 source.n49 a_n2224_n1288# 0.261326f
C276 source.n50 a_n2224_n1288# 0.058738f
C277 source.n51 a_n2224_n1288# 0.88633f
C278 source.n52 a_n2224_n1288# 0.053582f
C279 source.n53 a_n2224_n1288# 0.118556f
C280 source.t47 a_n2224_n1288# 0.08897f
C281 source.n54 a_n2224_n1288# 0.092786f
C282 source.n55 a_n2224_n1288# 0.029911f
C283 source.n56 a_n2224_n1288# 0.019727f
C284 source.n57 a_n2224_n1288# 0.261326f
C285 source.n58 a_n2224_n1288# 0.058738f
C286 source.n59 a_n2224_n1288# 0.88633f
C287 source.t39 a_n2224_n1288# 0.05802f
C288 source.t45 a_n2224_n1288# 0.05802f
C289 source.n60 a_n2224_n1288# 0.310171f
C290 source.n61 a_n2224_n1288# 0.403701f
C291 source.t34 a_n2224_n1288# 0.05802f
C292 source.t27 a_n2224_n1288# 0.05802f
C293 source.n62 a_n2224_n1288# 0.310171f
C294 source.n63 a_n2224_n1288# 0.403701f
C295 source.t31 a_n2224_n1288# 0.05802f
C296 source.t35 a_n2224_n1288# 0.05802f
C297 source.n64 a_n2224_n1288# 0.310171f
C298 source.n65 a_n2224_n1288# 0.403701f
C299 source.t30 a_n2224_n1288# 0.05802f
C300 source.t44 a_n2224_n1288# 0.05802f
C301 source.n66 a_n2224_n1288# 0.310171f
C302 source.n67 a_n2224_n1288# 0.403701f
C303 source.t41 a_n2224_n1288# 0.05802f
C304 source.t43 a_n2224_n1288# 0.05802f
C305 source.n68 a_n2224_n1288# 0.310171f
C306 source.n69 a_n2224_n1288# 0.403701f
C307 source.n70 a_n2224_n1288# 0.053582f
C308 source.n71 a_n2224_n1288# 0.118556f
C309 source.t37 a_n2224_n1288# 0.08897f
C310 source.n72 a_n2224_n1288# 0.092786f
C311 source.n73 a_n2224_n1288# 0.029911f
C312 source.n74 a_n2224_n1288# 0.019727f
C313 source.n75 a_n2224_n1288# 0.261326f
C314 source.n76 a_n2224_n1288# 0.058738f
C315 source.n77 a_n2224_n1288# 0.144943f
C316 source.n78 a_n2224_n1288# 0.053582f
C317 source.n79 a_n2224_n1288# 0.118556f
C318 source.t2 a_n2224_n1288# 0.08897f
C319 source.n80 a_n2224_n1288# 0.092786f
C320 source.n81 a_n2224_n1288# 0.029911f
C321 source.n82 a_n2224_n1288# 0.019727f
C322 source.n83 a_n2224_n1288# 0.261326f
C323 source.n84 a_n2224_n1288# 0.058738f
C324 source.n85 a_n2224_n1288# 0.144943f
C325 source.t21 a_n2224_n1288# 0.05802f
C326 source.t10 a_n2224_n1288# 0.05802f
C327 source.n86 a_n2224_n1288# 0.310171f
C328 source.n87 a_n2224_n1288# 0.403701f
C329 source.t4 a_n2224_n1288# 0.05802f
C330 source.t1 a_n2224_n1288# 0.05802f
C331 source.n88 a_n2224_n1288# 0.310171f
C332 source.n89 a_n2224_n1288# 0.403701f
C333 source.t19 a_n2224_n1288# 0.05802f
C334 source.t11 a_n2224_n1288# 0.05802f
C335 source.n90 a_n2224_n1288# 0.310171f
C336 source.n91 a_n2224_n1288# 0.403701f
C337 source.t20 a_n2224_n1288# 0.05802f
C338 source.t13 a_n2224_n1288# 0.05802f
C339 source.n92 a_n2224_n1288# 0.310171f
C340 source.n93 a_n2224_n1288# 0.403701f
C341 source.t8 a_n2224_n1288# 0.05802f
C342 source.t12 a_n2224_n1288# 0.05802f
C343 source.n94 a_n2224_n1288# 0.310171f
C344 source.n95 a_n2224_n1288# 0.403701f
C345 source.n96 a_n2224_n1288# 0.053582f
C346 source.n97 a_n2224_n1288# 0.118556f
C347 source.t16 a_n2224_n1288# 0.08897f
C348 source.n98 a_n2224_n1288# 0.092786f
C349 source.n99 a_n2224_n1288# 0.029911f
C350 source.n100 a_n2224_n1288# 0.019727f
C351 source.n101 a_n2224_n1288# 0.261326f
C352 source.n102 a_n2224_n1288# 0.058738f
C353 source.n103 a_n2224_n1288# 0.348093f
C354 source.n104 a_n2224_n1288# 0.905471f
C355 plus.n0 a_n2224_n1288# 0.039323f
C356 plus.t17 a_n2224_n1288# 0.057856f
C357 plus.t5 a_n2224_n1288# 0.057856f
C358 plus.n1 a_n2224_n1288# 0.014257f
C359 plus.n2 a_n2224_n1288# 0.039323f
C360 plus.t7 a_n2224_n1288# 0.057856f
C361 plus.t14 a_n2224_n1288# 0.057856f
C362 plus.t22 a_n2224_n1288# 0.057856f
C363 plus.n3 a_n2224_n1288# 0.042428f
C364 plus.n4 a_n2224_n1288# 0.039323f
C365 plus.t15 a_n2224_n1288# 0.057856f
C366 plus.t0 a_n2224_n1288# 0.057856f
C367 plus.n5 a_n2224_n1288# 0.013772f
C368 plus.t11 a_n2224_n1288# 0.061143f
C369 plus.n6 a_n2224_n1288# 0.052719f
C370 plus.t1 a_n2224_n1288# 0.057856f
C371 plus.n7 a_n2224_n1288# 0.042428f
C372 plus.t16 a_n2224_n1288# 0.057856f
C373 plus.n8 a_n2224_n1288# 0.042428f
C374 plus.n9 a_n2224_n1288# 0.014984f
C375 plus.n10 a_n2224_n1288# 0.081748f
C376 plus.n11 a_n2224_n1288# 0.039323f
C377 plus.n12 a_n2224_n1288# 0.039323f
C378 plus.n13 a_n2224_n1288# 0.014257f
C379 plus.n14 a_n2224_n1288# 0.042428f
C380 plus.n15 a_n2224_n1288# 0.014984f
C381 plus.n16 a_n2224_n1288# 0.042428f
C382 plus.n17 a_n2224_n1288# 0.014984f
C383 plus.n18 a_n2224_n1288# 0.039323f
C384 plus.n19 a_n2224_n1288# 0.039323f
C385 plus.n20 a_n2224_n1288# 0.014984f
C386 plus.n21 a_n2224_n1288# 0.042428f
C387 plus.n22 a_n2224_n1288# 0.014984f
C388 plus.n23 a_n2224_n1288# 0.042428f
C389 plus.t18 a_n2224_n1288# 0.057856f
C390 plus.n24 a_n2224_n1288# 0.042428f
C391 plus.n25 a_n2224_n1288# 0.014984f
C392 plus.n26 a_n2224_n1288# 0.039323f
C393 plus.n27 a_n2224_n1288# 0.039323f
C394 plus.n28 a_n2224_n1288# 0.039323f
C395 plus.n29 a_n2224_n1288# 0.013772f
C396 plus.n30 a_n2224_n1288# 0.042428f
C397 plus.n31 a_n2224_n1288# 0.014984f
C398 plus.n32 a_n2224_n1288# 0.042428f
C399 plus.t4 a_n2224_n1288# 0.061143f
C400 plus.n33 a_n2224_n1288# 0.05267f
C401 plus.n34 a_n2224_n1288# 0.27449f
C402 plus.n35 a_n2224_n1288# 0.039323f
C403 plus.t6 a_n2224_n1288# 0.061143f
C404 plus.t9 a_n2224_n1288# 0.057856f
C405 plus.t12 a_n2224_n1288# 0.057856f
C406 plus.n36 a_n2224_n1288# 0.014257f
C407 plus.n37 a_n2224_n1288# 0.039323f
C408 plus.t13 a_n2224_n1288# 0.057856f
C409 plus.n38 a_n2224_n1288# 0.042428f
C410 plus.t8 a_n2224_n1288# 0.057856f
C411 plus.t23 a_n2224_n1288# 0.057856f
C412 plus.t3 a_n2224_n1288# 0.057856f
C413 plus.n39 a_n2224_n1288# 0.042428f
C414 plus.n40 a_n2224_n1288# 0.039323f
C415 plus.t20 a_n2224_n1288# 0.057856f
C416 plus.t10 a_n2224_n1288# 0.057856f
C417 plus.n41 a_n2224_n1288# 0.013772f
C418 plus.t21 a_n2224_n1288# 0.061143f
C419 plus.n42 a_n2224_n1288# 0.052719f
C420 plus.t2 a_n2224_n1288# 0.057856f
C421 plus.n43 a_n2224_n1288# 0.042428f
C422 plus.t19 a_n2224_n1288# 0.057856f
C423 plus.n44 a_n2224_n1288# 0.042428f
C424 plus.n45 a_n2224_n1288# 0.014984f
C425 plus.n46 a_n2224_n1288# 0.081748f
C426 plus.n47 a_n2224_n1288# 0.039323f
C427 plus.n48 a_n2224_n1288# 0.039323f
C428 plus.n49 a_n2224_n1288# 0.014257f
C429 plus.n50 a_n2224_n1288# 0.042428f
C430 plus.n51 a_n2224_n1288# 0.014984f
C431 plus.n52 a_n2224_n1288# 0.042428f
C432 plus.n53 a_n2224_n1288# 0.014984f
C433 plus.n54 a_n2224_n1288# 0.039323f
C434 plus.n55 a_n2224_n1288# 0.039323f
C435 plus.n56 a_n2224_n1288# 0.014984f
C436 plus.n57 a_n2224_n1288# 0.042428f
C437 plus.n58 a_n2224_n1288# 0.014984f
C438 plus.n59 a_n2224_n1288# 0.042428f
C439 plus.n60 a_n2224_n1288# 0.014984f
C440 plus.n61 a_n2224_n1288# 0.039323f
C441 plus.n62 a_n2224_n1288# 0.039323f
C442 plus.n63 a_n2224_n1288# 0.039323f
C443 plus.n64 a_n2224_n1288# 0.013772f
C444 plus.n65 a_n2224_n1288# 0.042428f
C445 plus.n66 a_n2224_n1288# 0.014984f
C446 plus.n67 a_n2224_n1288# 0.042428f
C447 plus.n68 a_n2224_n1288# 0.05267f
C448 plus.n69 a_n2224_n1288# 0.966098f
.ends

