* NGSPICE file created from diffpair107.ext - technology: sky130A

.subckt diffpair107 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t22 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_left.t14 plus.t1 source.t31 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t13 plus.t2 source.t28 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t23 plus.t3 drain_left.t12 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 source.t8 minus.t0 drain_right.t15 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X5 drain_left.t11 plus.t4 source.t25 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X6 source.t13 minus.t1 drain_right.t14 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X7 a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X8 source.t30 plus.t5 drain_left.t10 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X9 source.t19 plus.t6 drain_left.t9 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X10 source.t17 plus.t7 drain_left.t8 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X11 drain_right.t13 minus.t2 source.t3 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 source.t1 minus.t3 drain_right.t12 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X13 source.t2 minus.t4 drain_right.t11 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X14 drain_right.t10 minus.t5 source.t5 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X15 source.t9 minus.t6 drain_right.t9 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X16 source.t16 plus.t8 drain_left.t7 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X17 source.t18 plus.t9 drain_left.t6 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X18 source.t27 plus.t10 drain_left.t5 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X19 a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X20 a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X21 source.t10 minus.t7 drain_right.t8 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X22 source.t0 minus.t8 drain_right.t7 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X23 drain_right.t6 minus.t9 source.t11 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X24 drain_right.t5 minus.t10 source.t7 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X25 drain_right.t4 minus.t11 source.t12 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X26 source.t15 minus.t12 drain_right.t3 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X27 drain_right.t2 minus.t13 source.t4 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X28 source.t24 plus.t11 drain_left.t4 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X29 drain_right.t1 minus.t14 source.t14 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X30 drain_right.t0 minus.t15 source.t6 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X31 drain_left.t3 plus.t12 source.t21 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X32 drain_left.t2 plus.t13 source.t29 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X33 drain_left.t1 plus.t14 source.t20 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X34 a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X35 drain_left.t0 plus.t15 source.t26 a_n1760_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
R0 plus.n4 plus.t7 359.017
R1 plus.n19 plus.t4 359.017
R2 plus.n25 plus.t13 359.017
R3 plus.n40 plus.t5 359.017
R4 plus.n5 plus.t1 318.12
R5 plus.n3 plus.t10 318.12
R6 plus.n10 plus.t0 318.12
R7 plus.n1 plus.t9 318.12
R8 plus.n16 plus.t14 318.12
R9 plus.n18 plus.t8 318.12
R10 plus.n26 plus.t11 318.12
R11 plus.n24 plus.t2 318.12
R12 plus.n31 plus.t6 318.12
R13 plus.n22 plus.t12 318.12
R14 plus.n37 plus.t3 318.12
R15 plus.n39 plus.t15 318.12
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus.n6 plus.n5 29.2126
R47 plus.n18 plus.n17 29.2126
R48 plus.n39 plus.n38 29.2126
R49 plus.n27 plus.n26 29.2126
R50 plus plus.n41 25.8475
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 8.32247
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n82 source.n80 289.615
R73 source.n68 source.n66 289.615
R74 source.n60 source.n58 289.615
R75 source.n46 source.n44 289.615
R76 source.n2 source.n0 289.615
R77 source.n16 source.n14 289.615
R78 source.n24 source.n22 289.615
R79 source.n38 source.n36 289.615
R80 source.n83 source.n82 185
R81 source.n69 source.n68 185
R82 source.n61 source.n60 185
R83 source.n47 source.n46 185
R84 source.n3 source.n2 185
R85 source.n17 source.n16 185
R86 source.n25 source.n24 185
R87 source.n39 source.n38 185
R88 source.t12 source.n81 167.117
R89 source.t0 source.n67 167.117
R90 source.t29 source.n59 167.117
R91 source.t30 source.n45 167.117
R92 source.t25 source.n1 167.117
R93 source.t17 source.n15 167.117
R94 source.t7 source.n23 167.117
R95 source.t1 source.n37 167.117
R96 source.n9 source.n8 84.1169
R97 source.n11 source.n10 84.1169
R98 source.n13 source.n12 84.1169
R99 source.n31 source.n30 84.1169
R100 source.n33 source.n32 84.1169
R101 source.n35 source.n34 84.1169
R102 source.n79 source.n78 84.1168
R103 source.n77 source.n76 84.1168
R104 source.n75 source.n74 84.1168
R105 source.n57 source.n56 84.1168
R106 source.n55 source.n54 84.1168
R107 source.n53 source.n52 84.1168
R108 source.n82 source.t12 52.3082
R109 source.n68 source.t0 52.3082
R110 source.n60 source.t29 52.3082
R111 source.n46 source.t30 52.3082
R112 source.n2 source.t25 52.3082
R113 source.n16 source.t17 52.3082
R114 source.n24 source.t7 52.3082
R115 source.n38 source.t1 52.3082
R116 source.n87 source.n86 31.4096
R117 source.n73 source.n72 31.4096
R118 source.n65 source.n64 31.4096
R119 source.n51 source.n50 31.4096
R120 source.n7 source.n6 31.4096
R121 source.n21 source.n20 31.4096
R122 source.n29 source.n28 31.4096
R123 source.n43 source.n42 31.4096
R124 source.n51 source.n43 14.212
R125 source.n78 source.t4 9.9005
R126 source.n78 source.t15 9.9005
R127 source.n76 source.t5 9.9005
R128 source.n76 source.t10 9.9005
R129 source.n74 source.t3 9.9005
R130 source.n74 source.t9 9.9005
R131 source.n56 source.t28 9.9005
R132 source.n56 source.t24 9.9005
R133 source.n54 source.t21 9.9005
R134 source.n54 source.t19 9.9005
R135 source.n52 source.t26 9.9005
R136 source.n52 source.t23 9.9005
R137 source.n8 source.t20 9.9005
R138 source.n8 source.t16 9.9005
R139 source.n10 source.t22 9.9005
R140 source.n10 source.t18 9.9005
R141 source.n12 source.t31 9.9005
R142 source.n12 source.t27 9.9005
R143 source.n30 source.t11 9.9005
R144 source.n30 source.t13 9.9005
R145 source.n32 source.t14 9.9005
R146 source.n32 source.t8 9.9005
R147 source.n34 source.t6 9.9005
R148 source.n34 source.t2 9.9005
R149 source.n83 source.n81 9.71174
R150 source.n69 source.n67 9.71174
R151 source.n61 source.n59 9.71174
R152 source.n47 source.n45 9.71174
R153 source.n3 source.n1 9.71174
R154 source.n17 source.n15 9.71174
R155 source.n25 source.n23 9.71174
R156 source.n39 source.n37 9.71174
R157 source.n86 source.n85 9.45567
R158 source.n72 source.n71 9.45567
R159 source.n64 source.n63 9.45567
R160 source.n50 source.n49 9.45567
R161 source.n6 source.n5 9.45567
R162 source.n20 source.n19 9.45567
R163 source.n28 source.n27 9.45567
R164 source.n42 source.n41 9.45567
R165 source.n85 source.n84 9.3005
R166 source.n71 source.n70 9.3005
R167 source.n63 source.n62 9.3005
R168 source.n49 source.n48 9.3005
R169 source.n5 source.n4 9.3005
R170 source.n19 source.n18 9.3005
R171 source.n27 source.n26 9.3005
R172 source.n41 source.n40 9.3005
R173 source.n88 source.n7 8.69904
R174 source.n86 source.n80 8.14595
R175 source.n72 source.n66 8.14595
R176 source.n64 source.n58 8.14595
R177 source.n50 source.n44 8.14595
R178 source.n6 source.n0 8.14595
R179 source.n20 source.n14 8.14595
R180 source.n28 source.n22 8.14595
R181 source.n42 source.n36 8.14595
R182 source.n84 source.n83 7.3702
R183 source.n70 source.n69 7.3702
R184 source.n62 source.n61 7.3702
R185 source.n48 source.n47 7.3702
R186 source.n4 source.n3 7.3702
R187 source.n18 source.n17 7.3702
R188 source.n26 source.n25 7.3702
R189 source.n40 source.n39 7.3702
R190 source.n84 source.n80 5.81868
R191 source.n70 source.n66 5.81868
R192 source.n62 source.n58 5.81868
R193 source.n48 source.n44 5.81868
R194 source.n4 source.n0 5.81868
R195 source.n18 source.n14 5.81868
R196 source.n26 source.n22 5.81868
R197 source.n40 source.n36 5.81868
R198 source.n88 source.n87 5.51343
R199 source.n85 source.n81 3.44771
R200 source.n71 source.n67 3.44771
R201 source.n63 source.n59 3.44771
R202 source.n49 source.n45 3.44771
R203 source.n5 source.n1 3.44771
R204 source.n19 source.n15 3.44771
R205 source.n27 source.n23 3.44771
R206 source.n41 source.n37 3.44771
R207 source.n43 source.n35 0.5005
R208 source.n35 source.n33 0.5005
R209 source.n33 source.n31 0.5005
R210 source.n31 source.n29 0.5005
R211 source.n21 source.n13 0.5005
R212 source.n13 source.n11 0.5005
R213 source.n11 source.n9 0.5005
R214 source.n9 source.n7 0.5005
R215 source.n53 source.n51 0.5005
R216 source.n55 source.n53 0.5005
R217 source.n57 source.n55 0.5005
R218 source.n65 source.n57 0.5005
R219 source.n75 source.n73 0.5005
R220 source.n77 source.n75 0.5005
R221 source.n79 source.n77 0.5005
R222 source.n87 source.n79 0.5005
R223 source.n29 source.n21 0.470328
R224 source.n73 source.n65 0.470328
R225 source source.n88 0.188
R226 drain_left.n9 drain_left.n7 101.296
R227 drain_left.n5 drain_left.n3 101.296
R228 drain_left.n2 drain_left.n0 101.296
R229 drain_left.n13 drain_left.n12 100.796
R230 drain_left.n11 drain_left.n10 100.796
R231 drain_left.n9 drain_left.n8 100.796
R232 drain_left.n5 drain_left.n4 100.796
R233 drain_left.n2 drain_left.n1 100.796
R234 drain_left drain_left.n6 23.0413
R235 drain_left.n3 drain_left.t4 9.9005
R236 drain_left.n3 drain_left.t2 9.9005
R237 drain_left.n4 drain_left.t9 9.9005
R238 drain_left.n4 drain_left.t13 9.9005
R239 drain_left.n1 drain_left.t12 9.9005
R240 drain_left.n1 drain_left.t3 9.9005
R241 drain_left.n0 drain_left.t10 9.9005
R242 drain_left.n0 drain_left.t0 9.9005
R243 drain_left.n12 drain_left.t7 9.9005
R244 drain_left.n12 drain_left.t11 9.9005
R245 drain_left.n10 drain_left.t6 9.9005
R246 drain_left.n10 drain_left.t1 9.9005
R247 drain_left.n8 drain_left.t5 9.9005
R248 drain_left.n8 drain_left.t15 9.9005
R249 drain_left.n7 drain_left.t8 9.9005
R250 drain_left.n7 drain_left.t14 9.9005
R251 drain_left drain_left.n13 6.15322
R252 drain_left.n11 drain_left.n9 0.5005
R253 drain_left.n13 drain_left.n11 0.5005
R254 drain_left.n6 drain_left.n5 0.195154
R255 drain_left.n6 drain_left.n2 0.195154
R256 minus.n19 minus.t3 359.017
R257 minus.n4 minus.t10 359.017
R258 minus.n40 minus.t11 359.017
R259 minus.n25 minus.t8 359.017
R260 minus.n18 minus.t15 318.12
R261 minus.n16 minus.t4 318.12
R262 minus.n1 minus.t14 318.12
R263 minus.n10 minus.t0 318.12
R264 minus.n3 minus.t9 318.12
R265 minus.n5 minus.t1 318.12
R266 minus.n39 minus.t12 318.12
R267 minus.n37 minus.t13 318.12
R268 minus.n22 minus.t7 318.12
R269 minus.n31 minus.t5 318.12
R270 minus.n24 minus.t6 318.12
R271 minus.n26 minus.t2 318.12
R272 minus.n7 minus.n4 161.489
R273 minus.n28 minus.n25 161.489
R274 minus.n20 minus.n19 161.3
R275 minus.n17 minus.n0 161.3
R276 minus.n15 minus.n14 161.3
R277 minus.n13 minus.n12 161.3
R278 minus.n11 minus.n2 161.3
R279 minus.n9 minus.n8 161.3
R280 minus.n7 minus.n6 161.3
R281 minus.n41 minus.n40 161.3
R282 minus.n38 minus.n21 161.3
R283 minus.n36 minus.n35 161.3
R284 minus.n34 minus.n33 161.3
R285 minus.n32 minus.n23 161.3
R286 minus.n30 minus.n29 161.3
R287 minus.n28 minus.n27 161.3
R288 minus.n12 minus.n11 73.0308
R289 minus.n33 minus.n32 73.0308
R290 minus.n15 minus.n1 67.1884
R291 minus.n10 minus.n9 67.1884
R292 minus.n31 minus.n30 67.1884
R293 minus.n36 minus.n22 67.1884
R294 minus.n17 minus.n16 55.5035
R295 minus.n6 minus.n3 55.5035
R296 minus.n27 minus.n24 55.5035
R297 minus.n38 minus.n37 55.5035
R298 minus.n19 minus.n18 43.8187
R299 minus.n5 minus.n4 43.8187
R300 minus.n26 minus.n25 43.8187
R301 minus.n40 minus.n39 43.8187
R302 minus.n18 minus.n17 29.2126
R303 minus.n6 minus.n5 29.2126
R304 minus.n27 minus.n26 29.2126
R305 minus.n39 minus.n38 29.2126
R306 minus.n42 minus.n20 28.1785
R307 minus.n16 minus.n15 17.5278
R308 minus.n9 minus.n3 17.5278
R309 minus.n30 minus.n24 17.5278
R310 minus.n37 minus.n36 17.5278
R311 minus.n42 minus.n41 6.46641
R312 minus.n12 minus.n1 5.84292
R313 minus.n11 minus.n10 5.84292
R314 minus.n32 minus.n31 5.84292
R315 minus.n33 minus.n22 5.84292
R316 minus.n20 minus.n0 0.189894
R317 minus.n14 minus.n0 0.189894
R318 minus.n14 minus.n13 0.189894
R319 minus.n13 minus.n2 0.189894
R320 minus.n8 minus.n2 0.189894
R321 minus.n8 minus.n7 0.189894
R322 minus.n29 minus.n28 0.189894
R323 minus.n29 minus.n23 0.189894
R324 minus.n34 minus.n23 0.189894
R325 minus.n35 minus.n34 0.189894
R326 minus.n35 minus.n21 0.189894
R327 minus.n41 minus.n21 0.189894
R328 minus minus.n42 0.188
R329 drain_right.n9 drain_right.n7 101.296
R330 drain_right.n5 drain_right.n3 101.296
R331 drain_right.n2 drain_right.n0 101.296
R332 drain_right.n9 drain_right.n8 100.796
R333 drain_right.n11 drain_right.n10 100.796
R334 drain_right.n13 drain_right.n12 100.796
R335 drain_right.n5 drain_right.n4 100.796
R336 drain_right.n2 drain_right.n1 100.796
R337 drain_right drain_right.n6 22.4881
R338 drain_right.n3 drain_right.t3 9.9005
R339 drain_right.n3 drain_right.t4 9.9005
R340 drain_right.n4 drain_right.t8 9.9005
R341 drain_right.n4 drain_right.t2 9.9005
R342 drain_right.n1 drain_right.t9 9.9005
R343 drain_right.n1 drain_right.t10 9.9005
R344 drain_right.n0 drain_right.t7 9.9005
R345 drain_right.n0 drain_right.t13 9.9005
R346 drain_right.n7 drain_right.t14 9.9005
R347 drain_right.n7 drain_right.t5 9.9005
R348 drain_right.n8 drain_right.t15 9.9005
R349 drain_right.n8 drain_right.t6 9.9005
R350 drain_right.n10 drain_right.t11 9.9005
R351 drain_right.n10 drain_right.t1 9.9005
R352 drain_right.n12 drain_right.t12 9.9005
R353 drain_right.n12 drain_right.t0 9.9005
R354 drain_right drain_right.n13 6.15322
R355 drain_right.n13 drain_right.n11 0.5005
R356 drain_right.n11 drain_right.n9 0.5005
R357 drain_right.n6 drain_right.n5 0.195154
R358 drain_right.n6 drain_right.n2 0.195154
C0 source drain_right 7.83877f
C1 source minus 1.44997f
C2 drain_left drain_right 0.897273f
C3 drain_left minus 0.177171f
C4 source plus 1.46394f
C5 drain_left plus 1.45741f
C6 drain_right minus 1.2871f
C7 plus drain_right 0.331152f
C8 plus minus 3.50621f
C9 source drain_left 7.83879f
C10 drain_right a_n1760_n1288# 3.91233f
C11 drain_left a_n1760_n1288# 4.15624f
C12 source a_n1760_n1288# 3.084316f
C13 minus a_n1760_n1288# 6.04853f
C14 plus a_n1760_n1288# 6.681848f
C15 drain_right.t7 a_n1760_n1288# 0.044354f
C16 drain_right.t13 a_n1760_n1288# 0.044354f
C17 drain_right.n0 a_n1760_n1288# 0.280211f
C18 drain_right.t9 a_n1760_n1288# 0.044354f
C19 drain_right.t10 a_n1760_n1288# 0.044354f
C20 drain_right.n1 a_n1760_n1288# 0.278649f
C21 drain_right.n2 a_n1760_n1288# 0.595934f
C22 drain_right.t3 a_n1760_n1288# 0.044354f
C23 drain_right.t4 a_n1760_n1288# 0.044354f
C24 drain_right.n3 a_n1760_n1288# 0.280211f
C25 drain_right.t8 a_n1760_n1288# 0.044354f
C26 drain_right.t2 a_n1760_n1288# 0.044354f
C27 drain_right.n4 a_n1760_n1288# 0.278649f
C28 drain_right.n5 a_n1760_n1288# 0.595934f
C29 drain_right.n6 a_n1760_n1288# 0.718345f
C30 drain_right.t14 a_n1760_n1288# 0.044354f
C31 drain_right.t5 a_n1760_n1288# 0.044354f
C32 drain_right.n7 a_n1760_n1288# 0.280213f
C33 drain_right.t15 a_n1760_n1288# 0.044354f
C34 drain_right.t6 a_n1760_n1288# 0.044354f
C35 drain_right.n8 a_n1760_n1288# 0.27865f
C36 drain_right.n9 a_n1760_n1288# 0.620202f
C37 drain_right.t11 a_n1760_n1288# 0.044354f
C38 drain_right.t1 a_n1760_n1288# 0.044354f
C39 drain_right.n10 a_n1760_n1288# 0.27865f
C40 drain_right.n11 a_n1760_n1288# 0.30523f
C41 drain_right.t12 a_n1760_n1288# 0.044354f
C42 drain_right.t0 a_n1760_n1288# 0.044354f
C43 drain_right.n12 a_n1760_n1288# 0.27865f
C44 drain_right.n13 a_n1760_n1288# 0.536882f
C45 minus.n0 a_n1760_n1288# 0.029041f
C46 minus.t3 a_n1760_n1288# 0.046358f
C47 minus.t15 a_n1760_n1288# 0.042727f
C48 minus.t4 a_n1760_n1288# 0.042727f
C49 minus.t14 a_n1760_n1288# 0.042727f
C50 minus.n1 a_n1760_n1288# 0.031333f
C51 minus.n2 a_n1760_n1288# 0.029041f
C52 minus.t0 a_n1760_n1288# 0.042727f
C53 minus.t9 a_n1760_n1288# 0.042727f
C54 minus.n3 a_n1760_n1288# 0.031333f
C55 minus.t10 a_n1760_n1288# 0.046358f
C56 minus.n4 a_n1760_n1288# 0.039347f
C57 minus.t1 a_n1760_n1288# 0.042727f
C58 minus.n5 a_n1760_n1288# 0.031333f
C59 minus.n6 a_n1760_n1288# 0.011066f
C60 minus.n7 a_n1760_n1288# 0.063591f
C61 minus.n8 a_n1760_n1288# 0.029041f
C62 minus.n9 a_n1760_n1288# 0.011066f
C63 minus.n10 a_n1760_n1288# 0.031333f
C64 minus.n11 a_n1760_n1288# 0.01035f
C65 minus.n12 a_n1760_n1288# 0.01035f
C66 minus.n13 a_n1760_n1288# 0.029041f
C67 minus.n14 a_n1760_n1288# 0.029041f
C68 minus.n15 a_n1760_n1288# 0.011066f
C69 minus.n16 a_n1760_n1288# 0.031333f
C70 minus.n17 a_n1760_n1288# 0.011066f
C71 minus.n18 a_n1760_n1288# 0.031333f
C72 minus.n19 a_n1760_n1288# 0.039306f
C73 minus.n20 a_n1760_n1288# 0.676678f
C74 minus.n21 a_n1760_n1288# 0.029041f
C75 minus.t12 a_n1760_n1288# 0.042727f
C76 minus.t13 a_n1760_n1288# 0.042727f
C77 minus.t7 a_n1760_n1288# 0.042727f
C78 minus.n22 a_n1760_n1288# 0.031333f
C79 minus.n23 a_n1760_n1288# 0.029041f
C80 minus.t5 a_n1760_n1288# 0.042727f
C81 minus.t6 a_n1760_n1288# 0.042727f
C82 minus.n24 a_n1760_n1288# 0.031333f
C83 minus.t8 a_n1760_n1288# 0.046358f
C84 minus.n25 a_n1760_n1288# 0.039347f
C85 minus.t2 a_n1760_n1288# 0.042727f
C86 minus.n26 a_n1760_n1288# 0.031333f
C87 minus.n27 a_n1760_n1288# 0.011066f
C88 minus.n28 a_n1760_n1288# 0.063591f
C89 minus.n29 a_n1760_n1288# 0.029041f
C90 minus.n30 a_n1760_n1288# 0.011066f
C91 minus.n31 a_n1760_n1288# 0.031333f
C92 minus.n32 a_n1760_n1288# 0.01035f
C93 minus.n33 a_n1760_n1288# 0.01035f
C94 minus.n34 a_n1760_n1288# 0.029041f
C95 minus.n35 a_n1760_n1288# 0.029041f
C96 minus.n36 a_n1760_n1288# 0.011066f
C97 minus.n37 a_n1760_n1288# 0.031333f
C98 minus.n38 a_n1760_n1288# 0.011066f
C99 minus.n39 a_n1760_n1288# 0.031333f
C100 minus.t11 a_n1760_n1288# 0.046358f
C101 minus.n40 a_n1760_n1288# 0.039306f
C102 minus.n41 a_n1760_n1288# 0.187557f
C103 minus.n42 a_n1760_n1288# 0.83772f
C104 drain_left.t10 a_n1760_n1288# 0.043739f
C105 drain_left.t0 a_n1760_n1288# 0.043739f
C106 drain_left.n0 a_n1760_n1288# 0.276322f
C107 drain_left.t12 a_n1760_n1288# 0.043739f
C108 drain_left.t3 a_n1760_n1288# 0.043739f
C109 drain_left.n1 a_n1760_n1288# 0.274781f
C110 drain_left.n2 a_n1760_n1288# 0.587663f
C111 drain_left.t4 a_n1760_n1288# 0.043739f
C112 drain_left.t2 a_n1760_n1288# 0.043739f
C113 drain_left.n3 a_n1760_n1288# 0.276322f
C114 drain_left.t9 a_n1760_n1288# 0.043739f
C115 drain_left.t13 a_n1760_n1288# 0.043739f
C116 drain_left.n4 a_n1760_n1288# 0.274781f
C117 drain_left.n5 a_n1760_n1288# 0.587663f
C118 drain_left.n6 a_n1760_n1288# 0.762633f
C119 drain_left.t8 a_n1760_n1288# 0.043739f
C120 drain_left.t14 a_n1760_n1288# 0.043739f
C121 drain_left.n7 a_n1760_n1288# 0.276323f
C122 drain_left.t5 a_n1760_n1288# 0.043739f
C123 drain_left.t15 a_n1760_n1288# 0.043739f
C124 drain_left.n8 a_n1760_n1288# 0.274783f
C125 drain_left.n9 a_n1760_n1288# 0.611594f
C126 drain_left.t6 a_n1760_n1288# 0.043739f
C127 drain_left.t1 a_n1760_n1288# 0.043739f
C128 drain_left.n10 a_n1760_n1288# 0.274783f
C129 drain_left.n11 a_n1760_n1288# 0.300994f
C130 drain_left.t7 a_n1760_n1288# 0.043739f
C131 drain_left.t11 a_n1760_n1288# 0.043739f
C132 drain_left.n12 a_n1760_n1288# 0.274783f
C133 drain_left.n13 a_n1760_n1288# 0.52943f
C134 source.n0 a_n1760_n1288# 0.041876f
C135 source.n1 a_n1760_n1288# 0.092656f
C136 source.t25 a_n1760_n1288# 0.069533f
C137 source.n2 a_n1760_n1288# 0.072516f
C138 source.n3 a_n1760_n1288# 0.023376f
C139 source.n4 a_n1760_n1288# 0.015417f
C140 source.n5 a_n1760_n1288# 0.204236f
C141 source.n6 a_n1760_n1288# 0.045906f
C142 source.n7 a_n1760_n1288# 0.426099f
C143 source.t20 a_n1760_n1288# 0.045345f
C144 source.t16 a_n1760_n1288# 0.045345f
C145 source.n8 a_n1760_n1288# 0.242411f
C146 source.n9 a_n1760_n1288# 0.315505f
C147 source.t22 a_n1760_n1288# 0.045345f
C148 source.t18 a_n1760_n1288# 0.045345f
C149 source.n10 a_n1760_n1288# 0.242411f
C150 source.n11 a_n1760_n1288# 0.315505f
C151 source.t31 a_n1760_n1288# 0.045345f
C152 source.t27 a_n1760_n1288# 0.045345f
C153 source.n12 a_n1760_n1288# 0.242411f
C154 source.n13 a_n1760_n1288# 0.315505f
C155 source.n14 a_n1760_n1288# 0.041876f
C156 source.n15 a_n1760_n1288# 0.092656f
C157 source.t17 a_n1760_n1288# 0.069533f
C158 source.n16 a_n1760_n1288# 0.072516f
C159 source.n17 a_n1760_n1288# 0.023376f
C160 source.n18 a_n1760_n1288# 0.015417f
C161 source.n19 a_n1760_n1288# 0.204236f
C162 source.n20 a_n1760_n1288# 0.045906f
C163 source.n21 a_n1760_n1288# 0.113278f
C164 source.n22 a_n1760_n1288# 0.041876f
C165 source.n23 a_n1760_n1288# 0.092656f
C166 source.t7 a_n1760_n1288# 0.069533f
C167 source.n24 a_n1760_n1288# 0.072516f
C168 source.n25 a_n1760_n1288# 0.023376f
C169 source.n26 a_n1760_n1288# 0.015417f
C170 source.n27 a_n1760_n1288# 0.204236f
C171 source.n28 a_n1760_n1288# 0.045906f
C172 source.n29 a_n1760_n1288# 0.113278f
C173 source.t11 a_n1760_n1288# 0.045345f
C174 source.t13 a_n1760_n1288# 0.045345f
C175 source.n30 a_n1760_n1288# 0.242411f
C176 source.n31 a_n1760_n1288# 0.315505f
C177 source.t14 a_n1760_n1288# 0.045345f
C178 source.t8 a_n1760_n1288# 0.045345f
C179 source.n32 a_n1760_n1288# 0.242411f
C180 source.n33 a_n1760_n1288# 0.315505f
C181 source.t6 a_n1760_n1288# 0.045345f
C182 source.t2 a_n1760_n1288# 0.045345f
C183 source.n34 a_n1760_n1288# 0.242411f
C184 source.n35 a_n1760_n1288# 0.315505f
C185 source.n36 a_n1760_n1288# 0.041876f
C186 source.n37 a_n1760_n1288# 0.092656f
C187 source.t1 a_n1760_n1288# 0.069533f
C188 source.n38 a_n1760_n1288# 0.072516f
C189 source.n39 a_n1760_n1288# 0.023376f
C190 source.n40 a_n1760_n1288# 0.015417f
C191 source.n41 a_n1760_n1288# 0.204236f
C192 source.n42 a_n1760_n1288# 0.045906f
C193 source.n43 a_n1760_n1288# 0.692699f
C194 source.n44 a_n1760_n1288# 0.041876f
C195 source.n45 a_n1760_n1288# 0.092656f
C196 source.t30 a_n1760_n1288# 0.069533f
C197 source.n46 a_n1760_n1288# 0.072516f
C198 source.n47 a_n1760_n1288# 0.023376f
C199 source.n48 a_n1760_n1288# 0.015417f
C200 source.n49 a_n1760_n1288# 0.204236f
C201 source.n50 a_n1760_n1288# 0.045906f
C202 source.n51 a_n1760_n1288# 0.692699f
C203 source.t26 a_n1760_n1288# 0.045345f
C204 source.t23 a_n1760_n1288# 0.045345f
C205 source.n52 a_n1760_n1288# 0.242409f
C206 source.n53 a_n1760_n1288# 0.315507f
C207 source.t21 a_n1760_n1288# 0.045345f
C208 source.t19 a_n1760_n1288# 0.045345f
C209 source.n54 a_n1760_n1288# 0.242409f
C210 source.n55 a_n1760_n1288# 0.315507f
C211 source.t28 a_n1760_n1288# 0.045345f
C212 source.t24 a_n1760_n1288# 0.045345f
C213 source.n56 a_n1760_n1288# 0.242409f
C214 source.n57 a_n1760_n1288# 0.315507f
C215 source.n58 a_n1760_n1288# 0.041876f
C216 source.n59 a_n1760_n1288# 0.092656f
C217 source.t29 a_n1760_n1288# 0.069533f
C218 source.n60 a_n1760_n1288# 0.072516f
C219 source.n61 a_n1760_n1288# 0.023376f
C220 source.n62 a_n1760_n1288# 0.015417f
C221 source.n63 a_n1760_n1288# 0.204236f
C222 source.n64 a_n1760_n1288# 0.045906f
C223 source.n65 a_n1760_n1288# 0.113278f
C224 source.n66 a_n1760_n1288# 0.041876f
C225 source.n67 a_n1760_n1288# 0.092656f
C226 source.t0 a_n1760_n1288# 0.069533f
C227 source.n68 a_n1760_n1288# 0.072516f
C228 source.n69 a_n1760_n1288# 0.023376f
C229 source.n70 a_n1760_n1288# 0.015417f
C230 source.n71 a_n1760_n1288# 0.204236f
C231 source.n72 a_n1760_n1288# 0.045906f
C232 source.n73 a_n1760_n1288# 0.113278f
C233 source.t3 a_n1760_n1288# 0.045345f
C234 source.t9 a_n1760_n1288# 0.045345f
C235 source.n74 a_n1760_n1288# 0.242409f
C236 source.n75 a_n1760_n1288# 0.315507f
C237 source.t5 a_n1760_n1288# 0.045345f
C238 source.t10 a_n1760_n1288# 0.045345f
C239 source.n76 a_n1760_n1288# 0.242409f
C240 source.n77 a_n1760_n1288# 0.315507f
C241 source.t4 a_n1760_n1288# 0.045345f
C242 source.t15 a_n1760_n1288# 0.045345f
C243 source.n78 a_n1760_n1288# 0.242409f
C244 source.n79 a_n1760_n1288# 0.315507f
C245 source.n80 a_n1760_n1288# 0.041876f
C246 source.n81 a_n1760_n1288# 0.092656f
C247 source.t12 a_n1760_n1288# 0.069533f
C248 source.n82 a_n1760_n1288# 0.072516f
C249 source.n83 a_n1760_n1288# 0.023376f
C250 source.n84 a_n1760_n1288# 0.015417f
C251 source.n85 a_n1760_n1288# 0.204236f
C252 source.n86 a_n1760_n1288# 0.045906f
C253 source.n87 a_n1760_n1288# 0.272047f
C254 source.n88 a_n1760_n1288# 0.707658f
C255 plus.n0 a_n1760_n1288# 0.029536f
C256 plus.t8 a_n1760_n1288# 0.043456f
C257 plus.t14 a_n1760_n1288# 0.043456f
C258 plus.t9 a_n1760_n1288# 0.043456f
C259 plus.n1 a_n1760_n1288# 0.031868f
C260 plus.n2 a_n1760_n1288# 0.029536f
C261 plus.t0 a_n1760_n1288# 0.043456f
C262 plus.t10 a_n1760_n1288# 0.043456f
C263 plus.n3 a_n1760_n1288# 0.031868f
C264 plus.t7 a_n1760_n1288# 0.047149f
C265 plus.n4 a_n1760_n1288# 0.040018f
C266 plus.t1 a_n1760_n1288# 0.043456f
C267 plus.n5 a_n1760_n1288# 0.031868f
C268 plus.n6 a_n1760_n1288# 0.011255f
C269 plus.n7 a_n1760_n1288# 0.064676f
C270 plus.n8 a_n1760_n1288# 0.029536f
C271 plus.n9 a_n1760_n1288# 0.011255f
C272 plus.n10 a_n1760_n1288# 0.031868f
C273 plus.n11 a_n1760_n1288# 0.010526f
C274 plus.n12 a_n1760_n1288# 0.010526f
C275 plus.n13 a_n1760_n1288# 0.029536f
C276 plus.n14 a_n1760_n1288# 0.029536f
C277 plus.n15 a_n1760_n1288# 0.011255f
C278 plus.n16 a_n1760_n1288# 0.031868f
C279 plus.n17 a_n1760_n1288# 0.011255f
C280 plus.n18 a_n1760_n1288# 0.031868f
C281 plus.t4 a_n1760_n1288# 0.047149f
C282 plus.n19 a_n1760_n1288# 0.039977f
C283 plus.n20 a_n1760_n1288# 0.208684f
C284 plus.n21 a_n1760_n1288# 0.029536f
C285 plus.t5 a_n1760_n1288# 0.047149f
C286 plus.t15 a_n1760_n1288# 0.043456f
C287 plus.t3 a_n1760_n1288# 0.043456f
C288 plus.t12 a_n1760_n1288# 0.043456f
C289 plus.n22 a_n1760_n1288# 0.031868f
C290 plus.n23 a_n1760_n1288# 0.029536f
C291 plus.t6 a_n1760_n1288# 0.043456f
C292 plus.t2 a_n1760_n1288# 0.043456f
C293 plus.n24 a_n1760_n1288# 0.031868f
C294 plus.t13 a_n1760_n1288# 0.047149f
C295 plus.n25 a_n1760_n1288# 0.040018f
C296 plus.t11 a_n1760_n1288# 0.043456f
C297 plus.n26 a_n1760_n1288# 0.031868f
C298 plus.n27 a_n1760_n1288# 0.011255f
C299 plus.n28 a_n1760_n1288# 0.064676f
C300 plus.n29 a_n1760_n1288# 0.029536f
C301 plus.n30 a_n1760_n1288# 0.011255f
C302 plus.n31 a_n1760_n1288# 0.031868f
C303 plus.n32 a_n1760_n1288# 0.010526f
C304 plus.n33 a_n1760_n1288# 0.010526f
C305 plus.n34 a_n1760_n1288# 0.029536f
C306 plus.n35 a_n1760_n1288# 0.029536f
C307 plus.n36 a_n1760_n1288# 0.011255f
C308 plus.n37 a_n1760_n1288# 0.031868f
C309 plus.n38 a_n1760_n1288# 0.011255f
C310 plus.n39 a_n1760_n1288# 0.031868f
C311 plus.n40 a_n1760_n1288# 0.039977f
C312 plus.n41 a_n1760_n1288# 0.657505f
.ends

