* NGSPICE file created from diffpair323.ext - technology: sky130A

.subckt diffpair323 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t7 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X2 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X3 source.t8 plus.t1 drain_left.t6 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X4 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X5 drain_left.t5 plus.t2 source.t6 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X6 drain_right.t7 minus.t0 source.t0 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X8 source.t15 minus.t1 drain_right.t6 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 source.t13 plus.t3 drain_left.t4 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 drain_right.t5 minus.t2 source.t2 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X11 source.t1 minus.t3 drain_right.t4 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X12 source.t14 minus.t4 drain_right.t3 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X13 source.t9 plus.t4 drain_left.t3 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X14 drain_right.t2 minus.t5 source.t3 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X15 drain_left.t2 plus.t5 source.t10 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X16 drain_right.t1 minus.t6 source.t4 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X17 source.t11 plus.t6 drain_left.t1 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 drain_left.t0 plus.t7 source.t12 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t5 minus.t7 drain_right.t0 a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n1 plus.t4 1724.25
R1 plus.n5 plus.t5 1724.25
R2 plus.n8 plus.t2 1724.25
R3 plus.n12 plus.t1 1724.25
R4 plus.n2 plus.t7 1654.87
R5 plus.n4 plus.t6 1654.87
R6 plus.n9 plus.t3 1654.87
R7 plus.n11 plus.t0 1654.87
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 47.4702
R15 plus.n4 plus.n3 47.4702
R16 plus.n11 plus.n10 47.4702
R17 plus.n10 plus.n9 47.4702
R18 plus plus.n13 27.1202
R19 plus.n2 plus.n1 25.5611
R20 plus.n5 plus.n4 25.5611
R21 plus.n12 plus.n11 25.5611
R22 plus.n9 plus.n8 25.5611
R23 plus plus.n6 11.0876
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n3 source.t9 52.1921
R27 source.n4 source.t2 52.1921
R28 source.n7 source.t14 52.1921
R29 source.n15 source.t4 52.1919
R30 source.n12 source.t5 52.1919
R31 source.n11 source.t6 52.1919
R32 source.n8 source.t8 52.1919
R33 source.n0 source.t10 52.1919
R34 source.n2 source.n1 48.8588
R35 source.n6 source.n5 48.8588
R36 source.n14 source.n13 48.8586
R37 source.n10 source.n9 48.8586
R38 source.n8 source.n7 19.5753
R39 source.n16 source.n0 14.0322
R40 source.n16 source.n15 5.5436
R41 source.n13 source.t0 3.33383
R42 source.n13 source.t1 3.33383
R43 source.n9 source.t7 3.33383
R44 source.n9 source.t13 3.33383
R45 source.n1 source.t12 3.33383
R46 source.n1 source.t11 3.33383
R47 source.n5 source.t3 3.33383
R48 source.n5 source.t15 3.33383
R49 source.n7 source.n6 0.560845
R50 source.n6 source.n4 0.560845
R51 source.n3 source.n2 0.560845
R52 source.n2 source.n0 0.560845
R53 source.n10 source.n8 0.560845
R54 source.n11 source.n10 0.560845
R55 source.n14 source.n12 0.560845
R56 source.n15 source.n14 0.560845
R57 source.n4 source.n3 0.470328
R58 source.n12 source.n11 0.470328
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 66.0979
R61 drain_left.n2 drain_left.n1 65.7622
R62 drain_left.n2 drain_left.n0 65.7622
R63 drain_left.n5 drain_left.n4 65.5374
R64 drain_left drain_left.n2 27.0556
R65 drain_left drain_left.n5 6.21356
R66 drain_left.n1 drain_left.t4 3.33383
R67 drain_left.n1 drain_left.t5 3.33383
R68 drain_left.n0 drain_left.t6 3.33383
R69 drain_left.n0 drain_left.t7 3.33383
R70 drain_left.n4 drain_left.t1 3.33383
R71 drain_left.n4 drain_left.t2 3.33383
R72 drain_left.n3 drain_left.t3 3.33383
R73 drain_left.n3 drain_left.t0 3.33383
R74 minus.n5 minus.t4 1724.25
R75 minus.n1 minus.t2 1724.25
R76 minus.n12 minus.t6 1724.25
R77 minus.n8 minus.t7 1724.25
R78 minus.n4 minus.t5 1654.87
R79 minus.n2 minus.t1 1654.87
R80 minus.n11 minus.t3 1654.87
R81 minus.n9 minus.t0 1654.87
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 47.4702
R89 minus.n3 minus.n2 47.4702
R90 minus.n10 minus.n9 47.4702
R91 minus.n11 minus.n10 47.4702
R92 minus.n14 minus.n6 32.1028
R93 minus.n5 minus.n4 25.5611
R94 minus.n2 minus.n1 25.5611
R95 minus.n9 minus.n8 25.5611
R96 minus.n12 minus.n11 25.5611
R97 minus.n14 minus.n13 6.58005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 66.0978
R102 drain_right.n2 drain_right.n1 65.7622
R103 drain_right.n2 drain_right.n0 65.7622
R104 drain_right.n5 drain_right.n4 65.5376
R105 drain_right drain_right.n2 26.5023
R106 drain_right drain_right.n5 6.21356
R107 drain_right.n1 drain_right.t4 3.33383
R108 drain_right.n1 drain_right.t1 3.33383
R109 drain_right.n0 drain_right.t0 3.33383
R110 drain_right.n0 drain_right.t7 3.33383
R111 drain_right.n3 drain_right.t6 3.33383
R112 drain_right.n3 drain_right.t5 3.33383
R113 drain_right.n4 drain_right.t3 3.33383
R114 drain_right.n4 drain_right.t2 3.33383
C0 source minus 1.30448f
C1 minus plus 4.27952f
C2 drain_right drain_left 0.640281f
C3 drain_right source 13.1429f
C4 drain_right plus 0.282599f
C5 drain_right minus 1.71899f
C6 source drain_left 13.1436f
C7 drain_left plus 1.84839f
C8 drain_left minus 0.170499f
C9 source plus 1.31852f
C10 drain_right a_n1366_n2688# 4.47982f
C11 drain_left a_n1366_n2688# 4.654f
C12 source a_n1366_n2688# 6.914804f
C13 minus a_n1366_n2688# 4.774579f
C14 plus a_n1366_n2688# 5.84083f
C15 drain_right.t0 a_n1366_n2688# 0.26476f
C16 drain_right.t7 a_n1366_n2688# 0.26476f
C17 drain_right.n0 a_n1366_n2688# 1.70937f
C18 drain_right.t4 a_n1366_n2688# 0.26476f
C19 drain_right.t1 a_n1366_n2688# 0.26476f
C20 drain_right.n1 a_n1366_n2688# 1.70937f
C21 drain_right.n2 a_n1366_n2688# 1.40681f
C22 drain_right.t6 a_n1366_n2688# 0.26476f
C23 drain_right.t5 a_n1366_n2688# 0.26476f
C24 drain_right.n3 a_n1366_n2688# 1.71094f
C25 drain_right.t3 a_n1366_n2688# 0.26476f
C26 drain_right.t2 a_n1366_n2688# 0.26476f
C27 drain_right.n4 a_n1366_n2688# 1.70845f
C28 drain_right.n5 a_n1366_n2688# 0.783636f
C29 minus.n0 a_n1366_n2688# 0.081721f
C30 minus.t4 a_n1366_n2688# 0.134537f
C31 minus.t5 a_n1366_n2688# 0.131998f
C32 minus.t1 a_n1366_n2688# 0.131998f
C33 minus.t2 a_n1366_n2688# 0.134537f
C34 minus.n1 a_n1366_n2688# 0.075252f
C35 minus.n2 a_n1366_n2688# 0.060438f
C36 minus.n3 a_n1366_n2688# 0.014638f
C37 minus.n4 a_n1366_n2688# 0.060438f
C38 minus.n5 a_n1366_n2688# 0.075197f
C39 minus.n6 a_n1366_n2688# 1.00818f
C40 minus.n7 a_n1366_n2688# 0.081721f
C41 minus.t3 a_n1366_n2688# 0.131998f
C42 minus.t0 a_n1366_n2688# 0.131998f
C43 minus.t7 a_n1366_n2688# 0.134537f
C44 minus.n8 a_n1366_n2688# 0.075252f
C45 minus.n9 a_n1366_n2688# 0.060438f
C46 minus.n10 a_n1366_n2688# 0.014638f
C47 minus.n11 a_n1366_n2688# 0.060438f
C48 minus.t6 a_n1366_n2688# 0.134537f
C49 minus.n12 a_n1366_n2688# 0.075197f
C50 minus.n13 a_n1366_n2688# 0.232073f
C51 minus.n14 a_n1366_n2688# 1.23558f
C52 drain_left.t6 a_n1366_n2688# 0.262832f
C53 drain_left.t7 a_n1366_n2688# 0.262832f
C54 drain_left.n0 a_n1366_n2688# 1.69692f
C55 drain_left.t4 a_n1366_n2688# 0.262832f
C56 drain_left.t5 a_n1366_n2688# 0.262832f
C57 drain_left.n1 a_n1366_n2688# 1.69692f
C58 drain_left.n2 a_n1366_n2688# 1.44722f
C59 drain_left.t3 a_n1366_n2688# 0.262832f
C60 drain_left.t0 a_n1366_n2688# 0.262832f
C61 drain_left.n3 a_n1366_n2688# 1.69849f
C62 drain_left.t1 a_n1366_n2688# 0.262832f
C63 drain_left.t2 a_n1366_n2688# 0.262832f
C64 drain_left.n4 a_n1366_n2688# 1.696f
C65 drain_left.n5 a_n1366_n2688# 0.777928f
C66 source.t10 a_n1366_n2688# 1.55854f
C67 source.n0 a_n1366_n2688# 0.869383f
C68 source.t12 a_n1366_n2688# 0.20622f
C69 source.t11 a_n1366_n2688# 0.20622f
C70 source.n1 a_n1366_n2688# 1.27961f
C71 source.n2 a_n1366_n2688# 0.247468f
C72 source.t9 a_n1366_n2688# 1.55854f
C73 source.n3 a_n1366_n2688# 0.334148f
C74 source.t2 a_n1366_n2688# 1.55854f
C75 source.n4 a_n1366_n2688# 0.334148f
C76 source.t3 a_n1366_n2688# 0.20622f
C77 source.t15 a_n1366_n2688# 0.20622f
C78 source.n5 a_n1366_n2688# 1.27961f
C79 source.n6 a_n1366_n2688# 0.247468f
C80 source.t14 a_n1366_n2688# 1.55854f
C81 source.n7 a_n1366_n2688# 1.14779f
C82 source.t8 a_n1366_n2688# 1.55854f
C83 source.n8 a_n1366_n2688# 1.14779f
C84 source.t7 a_n1366_n2688# 0.20622f
C85 source.t13 a_n1366_n2688# 0.20622f
C86 source.n9 a_n1366_n2688# 1.27961f
C87 source.n10 a_n1366_n2688# 0.247471f
C88 source.t6 a_n1366_n2688# 1.55854f
C89 source.n11 a_n1366_n2688# 0.334152f
C90 source.t5 a_n1366_n2688# 1.55854f
C91 source.n12 a_n1366_n2688# 0.334152f
C92 source.t0 a_n1366_n2688# 0.20622f
C93 source.t1 a_n1366_n2688# 0.20622f
C94 source.n13 a_n1366_n2688# 1.27961f
C95 source.n14 a_n1366_n2688# 0.247471f
C96 source.t4 a_n1366_n2688# 1.55854f
C97 source.n15 a_n1366_n2688# 0.44303f
C98 source.n16 a_n1366_n2688# 0.996785f
C99 plus.n0 a_n1366_n2688# 0.083069f
C100 plus.t6 a_n1366_n2688# 0.134175f
C101 plus.t7 a_n1366_n2688# 0.134175f
C102 plus.t4 a_n1366_n2688# 0.136756f
C103 plus.n1 a_n1366_n2688# 0.076494f
C104 plus.n2 a_n1366_n2688# 0.061435f
C105 plus.n3 a_n1366_n2688# 0.014879f
C106 plus.n4 a_n1366_n2688# 0.061435f
C107 plus.t5 a_n1366_n2688# 0.136756f
C108 plus.n5 a_n1366_n2688# 0.076437f
C109 plus.n6 a_n1366_n2688# 0.351336f
C110 plus.n7 a_n1366_n2688# 0.083069f
C111 plus.t1 a_n1366_n2688# 0.136756f
C112 plus.t0 a_n1366_n2688# 0.134175f
C113 plus.t3 a_n1366_n2688# 0.134175f
C114 plus.t2 a_n1366_n2688# 0.136756f
C115 plus.n8 a_n1366_n2688# 0.076494f
C116 plus.n9 a_n1366_n2688# 0.061435f
C117 plus.n10 a_n1366_n2688# 0.014879f
C118 plus.n11 a_n1366_n2688# 0.061435f
C119 plus.n12 a_n1366_n2688# 0.076437f
C120 plus.n13 a_n1366_n2688# 0.893235f
.ends

