* NGSPICE file created from diffpair423.ext - technology: sky130A

.subckt diffpair423 minus drain_right drain_left source plus
X0 a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X1 drain_left.t7 plus.t0 source.t4 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X2 drain_left.t6 plus.t1 source.t10 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X3 source.t1 minus.t0 drain_right.t7 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X4 a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X5 source.t12 minus.t1 drain_right.t6 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 drain_right.t5 minus.t2 source.t13 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X7 a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X8 source.t9 plus.t2 drain_left.t5 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X9 drain_left.t4 plus.t3 source.t8 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X11 source.t7 plus.t4 drain_left.t3 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X12 drain_right.t4 minus.t3 source.t14 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X13 drain_right.t3 minus.t4 source.t15 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X14 drain_right.t2 minus.t5 source.t0 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X15 source.t5 plus.t5 drain_left.t2 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X16 source.t3 minus.t6 drain_right.t1 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X17 drain_left.t1 plus.t6 source.t6 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X18 source.t2 minus.t7 drain_right.t0 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X19 source.t11 plus.t7 drain_left.t0 a_n1296_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n1 plus.t2 1336.16
R1 plus.n5 plus.t0 1336.16
R2 plus.n8 plus.t6 1336.16
R3 plus.n12 plus.t7 1336.16
R4 plus.n2 plus.t1 1282.12
R5 plus.n4 plus.t4 1282.12
R6 plus.n9 plus.t5 1282.12
R7 plus.n11 plus.t3 1282.12
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 27.9119
R23 plus plus.n6 12.1444
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n530 source.n470 289.615
R27 source.n462 source.n402 289.615
R28 source.n396 source.n336 289.615
R29 source.n328 source.n268 289.615
R30 source.n60 source.n0 289.615
R31 source.n128 source.n68 289.615
R32 source.n194 source.n134 289.615
R33 source.n262 source.n202 289.615
R34 source.n490 source.n489 185
R35 source.n495 source.n494 185
R36 source.n497 source.n496 185
R37 source.n486 source.n485 185
R38 source.n503 source.n502 185
R39 source.n505 source.n504 185
R40 source.n482 source.n481 185
R41 source.n512 source.n511 185
R42 source.n513 source.n480 185
R43 source.n515 source.n514 185
R44 source.n478 source.n477 185
R45 source.n521 source.n520 185
R46 source.n523 source.n522 185
R47 source.n474 source.n473 185
R48 source.n529 source.n528 185
R49 source.n531 source.n530 185
R50 source.n422 source.n421 185
R51 source.n427 source.n426 185
R52 source.n429 source.n428 185
R53 source.n418 source.n417 185
R54 source.n435 source.n434 185
R55 source.n437 source.n436 185
R56 source.n414 source.n413 185
R57 source.n444 source.n443 185
R58 source.n445 source.n412 185
R59 source.n447 source.n446 185
R60 source.n410 source.n409 185
R61 source.n453 source.n452 185
R62 source.n455 source.n454 185
R63 source.n406 source.n405 185
R64 source.n461 source.n460 185
R65 source.n463 source.n462 185
R66 source.n356 source.n355 185
R67 source.n361 source.n360 185
R68 source.n363 source.n362 185
R69 source.n352 source.n351 185
R70 source.n369 source.n368 185
R71 source.n371 source.n370 185
R72 source.n348 source.n347 185
R73 source.n378 source.n377 185
R74 source.n379 source.n346 185
R75 source.n381 source.n380 185
R76 source.n344 source.n343 185
R77 source.n387 source.n386 185
R78 source.n389 source.n388 185
R79 source.n340 source.n339 185
R80 source.n395 source.n394 185
R81 source.n397 source.n396 185
R82 source.n288 source.n287 185
R83 source.n293 source.n292 185
R84 source.n295 source.n294 185
R85 source.n284 source.n283 185
R86 source.n301 source.n300 185
R87 source.n303 source.n302 185
R88 source.n280 source.n279 185
R89 source.n310 source.n309 185
R90 source.n311 source.n278 185
R91 source.n313 source.n312 185
R92 source.n276 source.n275 185
R93 source.n319 source.n318 185
R94 source.n321 source.n320 185
R95 source.n272 source.n271 185
R96 source.n327 source.n326 185
R97 source.n329 source.n328 185
R98 source.n61 source.n60 185
R99 source.n59 source.n58 185
R100 source.n4 source.n3 185
R101 source.n53 source.n52 185
R102 source.n51 source.n50 185
R103 source.n8 source.n7 185
R104 source.n45 source.n44 185
R105 source.n43 source.n10 185
R106 source.n42 source.n41 185
R107 source.n13 source.n11 185
R108 source.n36 source.n35 185
R109 source.n34 source.n33 185
R110 source.n17 source.n16 185
R111 source.n28 source.n27 185
R112 source.n26 source.n25 185
R113 source.n21 source.n20 185
R114 source.n129 source.n128 185
R115 source.n127 source.n126 185
R116 source.n72 source.n71 185
R117 source.n121 source.n120 185
R118 source.n119 source.n118 185
R119 source.n76 source.n75 185
R120 source.n113 source.n112 185
R121 source.n111 source.n78 185
R122 source.n110 source.n109 185
R123 source.n81 source.n79 185
R124 source.n104 source.n103 185
R125 source.n102 source.n101 185
R126 source.n85 source.n84 185
R127 source.n96 source.n95 185
R128 source.n94 source.n93 185
R129 source.n89 source.n88 185
R130 source.n195 source.n194 185
R131 source.n193 source.n192 185
R132 source.n138 source.n137 185
R133 source.n187 source.n186 185
R134 source.n185 source.n184 185
R135 source.n142 source.n141 185
R136 source.n179 source.n178 185
R137 source.n177 source.n144 185
R138 source.n176 source.n175 185
R139 source.n147 source.n145 185
R140 source.n170 source.n169 185
R141 source.n168 source.n167 185
R142 source.n151 source.n150 185
R143 source.n162 source.n161 185
R144 source.n160 source.n159 185
R145 source.n155 source.n154 185
R146 source.n263 source.n262 185
R147 source.n261 source.n260 185
R148 source.n206 source.n205 185
R149 source.n255 source.n254 185
R150 source.n253 source.n252 185
R151 source.n210 source.n209 185
R152 source.n247 source.n246 185
R153 source.n245 source.n212 185
R154 source.n244 source.n243 185
R155 source.n215 source.n213 185
R156 source.n238 source.n237 185
R157 source.n236 source.n235 185
R158 source.n219 source.n218 185
R159 source.n230 source.n229 185
R160 source.n228 source.n227 185
R161 source.n223 source.n222 185
R162 source.n491 source.t0 149.524
R163 source.n423 source.t2 149.524
R164 source.n357 source.t6 149.524
R165 source.n289 source.t11 149.524
R166 source.n22 source.t4 149.524
R167 source.n90 source.t9 149.524
R168 source.n156 source.t15 149.524
R169 source.n224 source.t1 149.524
R170 source.n495 source.n489 104.615
R171 source.n496 source.n495 104.615
R172 source.n496 source.n485 104.615
R173 source.n503 source.n485 104.615
R174 source.n504 source.n503 104.615
R175 source.n504 source.n481 104.615
R176 source.n512 source.n481 104.615
R177 source.n513 source.n512 104.615
R178 source.n514 source.n513 104.615
R179 source.n514 source.n477 104.615
R180 source.n521 source.n477 104.615
R181 source.n522 source.n521 104.615
R182 source.n522 source.n473 104.615
R183 source.n529 source.n473 104.615
R184 source.n530 source.n529 104.615
R185 source.n427 source.n421 104.615
R186 source.n428 source.n427 104.615
R187 source.n428 source.n417 104.615
R188 source.n435 source.n417 104.615
R189 source.n436 source.n435 104.615
R190 source.n436 source.n413 104.615
R191 source.n444 source.n413 104.615
R192 source.n445 source.n444 104.615
R193 source.n446 source.n445 104.615
R194 source.n446 source.n409 104.615
R195 source.n453 source.n409 104.615
R196 source.n454 source.n453 104.615
R197 source.n454 source.n405 104.615
R198 source.n461 source.n405 104.615
R199 source.n462 source.n461 104.615
R200 source.n361 source.n355 104.615
R201 source.n362 source.n361 104.615
R202 source.n362 source.n351 104.615
R203 source.n369 source.n351 104.615
R204 source.n370 source.n369 104.615
R205 source.n370 source.n347 104.615
R206 source.n378 source.n347 104.615
R207 source.n379 source.n378 104.615
R208 source.n380 source.n379 104.615
R209 source.n380 source.n343 104.615
R210 source.n387 source.n343 104.615
R211 source.n388 source.n387 104.615
R212 source.n388 source.n339 104.615
R213 source.n395 source.n339 104.615
R214 source.n396 source.n395 104.615
R215 source.n293 source.n287 104.615
R216 source.n294 source.n293 104.615
R217 source.n294 source.n283 104.615
R218 source.n301 source.n283 104.615
R219 source.n302 source.n301 104.615
R220 source.n302 source.n279 104.615
R221 source.n310 source.n279 104.615
R222 source.n311 source.n310 104.615
R223 source.n312 source.n311 104.615
R224 source.n312 source.n275 104.615
R225 source.n319 source.n275 104.615
R226 source.n320 source.n319 104.615
R227 source.n320 source.n271 104.615
R228 source.n327 source.n271 104.615
R229 source.n328 source.n327 104.615
R230 source.n60 source.n59 104.615
R231 source.n59 source.n3 104.615
R232 source.n52 source.n3 104.615
R233 source.n52 source.n51 104.615
R234 source.n51 source.n7 104.615
R235 source.n44 source.n7 104.615
R236 source.n44 source.n43 104.615
R237 source.n43 source.n42 104.615
R238 source.n42 source.n11 104.615
R239 source.n35 source.n11 104.615
R240 source.n35 source.n34 104.615
R241 source.n34 source.n16 104.615
R242 source.n27 source.n16 104.615
R243 source.n27 source.n26 104.615
R244 source.n26 source.n20 104.615
R245 source.n128 source.n127 104.615
R246 source.n127 source.n71 104.615
R247 source.n120 source.n71 104.615
R248 source.n120 source.n119 104.615
R249 source.n119 source.n75 104.615
R250 source.n112 source.n75 104.615
R251 source.n112 source.n111 104.615
R252 source.n111 source.n110 104.615
R253 source.n110 source.n79 104.615
R254 source.n103 source.n79 104.615
R255 source.n103 source.n102 104.615
R256 source.n102 source.n84 104.615
R257 source.n95 source.n84 104.615
R258 source.n95 source.n94 104.615
R259 source.n94 source.n88 104.615
R260 source.n194 source.n193 104.615
R261 source.n193 source.n137 104.615
R262 source.n186 source.n137 104.615
R263 source.n186 source.n185 104.615
R264 source.n185 source.n141 104.615
R265 source.n178 source.n141 104.615
R266 source.n178 source.n177 104.615
R267 source.n177 source.n176 104.615
R268 source.n176 source.n145 104.615
R269 source.n169 source.n145 104.615
R270 source.n169 source.n168 104.615
R271 source.n168 source.n150 104.615
R272 source.n161 source.n150 104.615
R273 source.n161 source.n160 104.615
R274 source.n160 source.n154 104.615
R275 source.n262 source.n261 104.615
R276 source.n261 source.n205 104.615
R277 source.n254 source.n205 104.615
R278 source.n254 source.n253 104.615
R279 source.n253 source.n209 104.615
R280 source.n246 source.n209 104.615
R281 source.n246 source.n245 104.615
R282 source.n245 source.n244 104.615
R283 source.n244 source.n213 104.615
R284 source.n237 source.n213 104.615
R285 source.n237 source.n236 104.615
R286 source.n236 source.n218 104.615
R287 source.n229 source.n218 104.615
R288 source.n229 source.n228 104.615
R289 source.n228 source.n222 104.615
R290 source.t0 source.n489 52.3082
R291 source.t2 source.n421 52.3082
R292 source.t6 source.n355 52.3082
R293 source.t11 source.n287 52.3082
R294 source.t4 source.n20 52.3082
R295 source.t9 source.n88 52.3082
R296 source.t15 source.n154 52.3082
R297 source.t1 source.n222 52.3082
R298 source.n67 source.n66 42.8739
R299 source.n201 source.n200 42.8739
R300 source.n469 source.n468 42.8737
R301 source.n335 source.n334 42.8737
R302 source.n535 source.n534 29.8581
R303 source.n467 source.n466 29.8581
R304 source.n401 source.n400 29.8581
R305 source.n333 source.n332 29.8581
R306 source.n65 source.n64 29.8581
R307 source.n133 source.n132 29.8581
R308 source.n199 source.n198 29.8581
R309 source.n267 source.n266 29.8581
R310 source.n333 source.n267 21.7877
R311 source.n536 source.n65 16.2748
R312 source.n515 source.n480 13.1884
R313 source.n447 source.n412 13.1884
R314 source.n381 source.n346 13.1884
R315 source.n313 source.n278 13.1884
R316 source.n45 source.n10 13.1884
R317 source.n113 source.n78 13.1884
R318 source.n179 source.n144 13.1884
R319 source.n247 source.n212 13.1884
R320 source.n511 source.n510 12.8005
R321 source.n516 source.n478 12.8005
R322 source.n443 source.n442 12.8005
R323 source.n448 source.n410 12.8005
R324 source.n377 source.n376 12.8005
R325 source.n382 source.n344 12.8005
R326 source.n309 source.n308 12.8005
R327 source.n314 source.n276 12.8005
R328 source.n46 source.n8 12.8005
R329 source.n41 source.n12 12.8005
R330 source.n114 source.n76 12.8005
R331 source.n109 source.n80 12.8005
R332 source.n180 source.n142 12.8005
R333 source.n175 source.n146 12.8005
R334 source.n248 source.n210 12.8005
R335 source.n243 source.n214 12.8005
R336 source.n509 source.n482 12.0247
R337 source.n520 source.n519 12.0247
R338 source.n441 source.n414 12.0247
R339 source.n452 source.n451 12.0247
R340 source.n375 source.n348 12.0247
R341 source.n386 source.n385 12.0247
R342 source.n307 source.n280 12.0247
R343 source.n318 source.n317 12.0247
R344 source.n50 source.n49 12.0247
R345 source.n40 source.n13 12.0247
R346 source.n118 source.n117 12.0247
R347 source.n108 source.n81 12.0247
R348 source.n184 source.n183 12.0247
R349 source.n174 source.n147 12.0247
R350 source.n252 source.n251 12.0247
R351 source.n242 source.n215 12.0247
R352 source.n506 source.n505 11.249
R353 source.n523 source.n476 11.249
R354 source.n438 source.n437 11.249
R355 source.n455 source.n408 11.249
R356 source.n372 source.n371 11.249
R357 source.n389 source.n342 11.249
R358 source.n304 source.n303 11.249
R359 source.n321 source.n274 11.249
R360 source.n53 source.n6 11.249
R361 source.n37 source.n36 11.249
R362 source.n121 source.n74 11.249
R363 source.n105 source.n104 11.249
R364 source.n187 source.n140 11.249
R365 source.n171 source.n170 11.249
R366 source.n255 source.n208 11.249
R367 source.n239 source.n238 11.249
R368 source.n502 source.n484 10.4732
R369 source.n524 source.n474 10.4732
R370 source.n434 source.n416 10.4732
R371 source.n456 source.n406 10.4732
R372 source.n368 source.n350 10.4732
R373 source.n390 source.n340 10.4732
R374 source.n300 source.n282 10.4732
R375 source.n322 source.n272 10.4732
R376 source.n54 source.n4 10.4732
R377 source.n33 source.n15 10.4732
R378 source.n122 source.n72 10.4732
R379 source.n101 source.n83 10.4732
R380 source.n188 source.n138 10.4732
R381 source.n167 source.n149 10.4732
R382 source.n256 source.n206 10.4732
R383 source.n235 source.n217 10.4732
R384 source.n491 source.n490 10.2747
R385 source.n423 source.n422 10.2747
R386 source.n357 source.n356 10.2747
R387 source.n289 source.n288 10.2747
R388 source.n22 source.n21 10.2747
R389 source.n90 source.n89 10.2747
R390 source.n156 source.n155 10.2747
R391 source.n224 source.n223 10.2747
R392 source.n501 source.n486 9.69747
R393 source.n528 source.n527 9.69747
R394 source.n433 source.n418 9.69747
R395 source.n460 source.n459 9.69747
R396 source.n367 source.n352 9.69747
R397 source.n394 source.n393 9.69747
R398 source.n299 source.n284 9.69747
R399 source.n326 source.n325 9.69747
R400 source.n58 source.n57 9.69747
R401 source.n32 source.n17 9.69747
R402 source.n126 source.n125 9.69747
R403 source.n100 source.n85 9.69747
R404 source.n192 source.n191 9.69747
R405 source.n166 source.n151 9.69747
R406 source.n260 source.n259 9.69747
R407 source.n234 source.n219 9.69747
R408 source.n534 source.n533 9.45567
R409 source.n466 source.n465 9.45567
R410 source.n400 source.n399 9.45567
R411 source.n332 source.n331 9.45567
R412 source.n64 source.n63 9.45567
R413 source.n132 source.n131 9.45567
R414 source.n198 source.n197 9.45567
R415 source.n266 source.n265 9.45567
R416 source.n533 source.n532 9.3005
R417 source.n472 source.n471 9.3005
R418 source.n527 source.n526 9.3005
R419 source.n525 source.n524 9.3005
R420 source.n476 source.n475 9.3005
R421 source.n519 source.n518 9.3005
R422 source.n517 source.n516 9.3005
R423 source.n493 source.n492 9.3005
R424 source.n488 source.n487 9.3005
R425 source.n499 source.n498 9.3005
R426 source.n501 source.n500 9.3005
R427 source.n484 source.n483 9.3005
R428 source.n507 source.n506 9.3005
R429 source.n509 source.n508 9.3005
R430 source.n510 source.n479 9.3005
R431 source.n465 source.n464 9.3005
R432 source.n404 source.n403 9.3005
R433 source.n459 source.n458 9.3005
R434 source.n457 source.n456 9.3005
R435 source.n408 source.n407 9.3005
R436 source.n451 source.n450 9.3005
R437 source.n449 source.n448 9.3005
R438 source.n425 source.n424 9.3005
R439 source.n420 source.n419 9.3005
R440 source.n431 source.n430 9.3005
R441 source.n433 source.n432 9.3005
R442 source.n416 source.n415 9.3005
R443 source.n439 source.n438 9.3005
R444 source.n441 source.n440 9.3005
R445 source.n442 source.n411 9.3005
R446 source.n399 source.n398 9.3005
R447 source.n338 source.n337 9.3005
R448 source.n393 source.n392 9.3005
R449 source.n391 source.n390 9.3005
R450 source.n342 source.n341 9.3005
R451 source.n385 source.n384 9.3005
R452 source.n383 source.n382 9.3005
R453 source.n359 source.n358 9.3005
R454 source.n354 source.n353 9.3005
R455 source.n365 source.n364 9.3005
R456 source.n367 source.n366 9.3005
R457 source.n350 source.n349 9.3005
R458 source.n373 source.n372 9.3005
R459 source.n375 source.n374 9.3005
R460 source.n376 source.n345 9.3005
R461 source.n331 source.n330 9.3005
R462 source.n270 source.n269 9.3005
R463 source.n325 source.n324 9.3005
R464 source.n323 source.n322 9.3005
R465 source.n274 source.n273 9.3005
R466 source.n317 source.n316 9.3005
R467 source.n315 source.n314 9.3005
R468 source.n291 source.n290 9.3005
R469 source.n286 source.n285 9.3005
R470 source.n297 source.n296 9.3005
R471 source.n299 source.n298 9.3005
R472 source.n282 source.n281 9.3005
R473 source.n305 source.n304 9.3005
R474 source.n307 source.n306 9.3005
R475 source.n308 source.n277 9.3005
R476 source.n24 source.n23 9.3005
R477 source.n19 source.n18 9.3005
R478 source.n30 source.n29 9.3005
R479 source.n32 source.n31 9.3005
R480 source.n15 source.n14 9.3005
R481 source.n38 source.n37 9.3005
R482 source.n40 source.n39 9.3005
R483 source.n12 source.n9 9.3005
R484 source.n63 source.n62 9.3005
R485 source.n2 source.n1 9.3005
R486 source.n57 source.n56 9.3005
R487 source.n55 source.n54 9.3005
R488 source.n6 source.n5 9.3005
R489 source.n49 source.n48 9.3005
R490 source.n47 source.n46 9.3005
R491 source.n92 source.n91 9.3005
R492 source.n87 source.n86 9.3005
R493 source.n98 source.n97 9.3005
R494 source.n100 source.n99 9.3005
R495 source.n83 source.n82 9.3005
R496 source.n106 source.n105 9.3005
R497 source.n108 source.n107 9.3005
R498 source.n80 source.n77 9.3005
R499 source.n131 source.n130 9.3005
R500 source.n70 source.n69 9.3005
R501 source.n125 source.n124 9.3005
R502 source.n123 source.n122 9.3005
R503 source.n74 source.n73 9.3005
R504 source.n117 source.n116 9.3005
R505 source.n115 source.n114 9.3005
R506 source.n158 source.n157 9.3005
R507 source.n153 source.n152 9.3005
R508 source.n164 source.n163 9.3005
R509 source.n166 source.n165 9.3005
R510 source.n149 source.n148 9.3005
R511 source.n172 source.n171 9.3005
R512 source.n174 source.n173 9.3005
R513 source.n146 source.n143 9.3005
R514 source.n197 source.n196 9.3005
R515 source.n136 source.n135 9.3005
R516 source.n191 source.n190 9.3005
R517 source.n189 source.n188 9.3005
R518 source.n140 source.n139 9.3005
R519 source.n183 source.n182 9.3005
R520 source.n181 source.n180 9.3005
R521 source.n226 source.n225 9.3005
R522 source.n221 source.n220 9.3005
R523 source.n232 source.n231 9.3005
R524 source.n234 source.n233 9.3005
R525 source.n217 source.n216 9.3005
R526 source.n240 source.n239 9.3005
R527 source.n242 source.n241 9.3005
R528 source.n214 source.n211 9.3005
R529 source.n265 source.n264 9.3005
R530 source.n204 source.n203 9.3005
R531 source.n259 source.n258 9.3005
R532 source.n257 source.n256 9.3005
R533 source.n208 source.n207 9.3005
R534 source.n251 source.n250 9.3005
R535 source.n249 source.n248 9.3005
R536 source.n498 source.n497 8.92171
R537 source.n531 source.n472 8.92171
R538 source.n430 source.n429 8.92171
R539 source.n463 source.n404 8.92171
R540 source.n364 source.n363 8.92171
R541 source.n397 source.n338 8.92171
R542 source.n296 source.n295 8.92171
R543 source.n329 source.n270 8.92171
R544 source.n61 source.n2 8.92171
R545 source.n29 source.n28 8.92171
R546 source.n129 source.n70 8.92171
R547 source.n97 source.n96 8.92171
R548 source.n195 source.n136 8.92171
R549 source.n163 source.n162 8.92171
R550 source.n263 source.n204 8.92171
R551 source.n231 source.n230 8.92171
R552 source.n494 source.n488 8.14595
R553 source.n532 source.n470 8.14595
R554 source.n426 source.n420 8.14595
R555 source.n464 source.n402 8.14595
R556 source.n360 source.n354 8.14595
R557 source.n398 source.n336 8.14595
R558 source.n292 source.n286 8.14595
R559 source.n330 source.n268 8.14595
R560 source.n62 source.n0 8.14595
R561 source.n25 source.n19 8.14595
R562 source.n130 source.n68 8.14595
R563 source.n93 source.n87 8.14595
R564 source.n196 source.n134 8.14595
R565 source.n159 source.n153 8.14595
R566 source.n264 source.n202 8.14595
R567 source.n227 source.n221 8.14595
R568 source.n493 source.n490 7.3702
R569 source.n425 source.n422 7.3702
R570 source.n359 source.n356 7.3702
R571 source.n291 source.n288 7.3702
R572 source.n24 source.n21 7.3702
R573 source.n92 source.n89 7.3702
R574 source.n158 source.n155 7.3702
R575 source.n226 source.n223 7.3702
R576 source.n494 source.n493 5.81868
R577 source.n534 source.n470 5.81868
R578 source.n426 source.n425 5.81868
R579 source.n466 source.n402 5.81868
R580 source.n360 source.n359 5.81868
R581 source.n400 source.n336 5.81868
R582 source.n292 source.n291 5.81868
R583 source.n332 source.n268 5.81868
R584 source.n64 source.n0 5.81868
R585 source.n25 source.n24 5.81868
R586 source.n132 source.n68 5.81868
R587 source.n93 source.n92 5.81868
R588 source.n198 source.n134 5.81868
R589 source.n159 source.n158 5.81868
R590 source.n266 source.n202 5.81868
R591 source.n227 source.n226 5.81868
R592 source.n536 source.n535 5.51343
R593 source.n497 source.n488 5.04292
R594 source.n532 source.n531 5.04292
R595 source.n429 source.n420 5.04292
R596 source.n464 source.n463 5.04292
R597 source.n363 source.n354 5.04292
R598 source.n398 source.n397 5.04292
R599 source.n295 source.n286 5.04292
R600 source.n330 source.n329 5.04292
R601 source.n62 source.n61 5.04292
R602 source.n28 source.n19 5.04292
R603 source.n130 source.n129 5.04292
R604 source.n96 source.n87 5.04292
R605 source.n196 source.n195 5.04292
R606 source.n162 source.n153 5.04292
R607 source.n264 source.n263 5.04292
R608 source.n230 source.n221 5.04292
R609 source.n498 source.n486 4.26717
R610 source.n528 source.n472 4.26717
R611 source.n430 source.n418 4.26717
R612 source.n460 source.n404 4.26717
R613 source.n364 source.n352 4.26717
R614 source.n394 source.n338 4.26717
R615 source.n296 source.n284 4.26717
R616 source.n326 source.n270 4.26717
R617 source.n58 source.n2 4.26717
R618 source.n29 source.n17 4.26717
R619 source.n126 source.n70 4.26717
R620 source.n97 source.n85 4.26717
R621 source.n192 source.n136 4.26717
R622 source.n163 source.n151 4.26717
R623 source.n260 source.n204 4.26717
R624 source.n231 source.n219 4.26717
R625 source.n502 source.n501 3.49141
R626 source.n527 source.n474 3.49141
R627 source.n434 source.n433 3.49141
R628 source.n459 source.n406 3.49141
R629 source.n368 source.n367 3.49141
R630 source.n393 source.n340 3.49141
R631 source.n300 source.n299 3.49141
R632 source.n325 source.n272 3.49141
R633 source.n57 source.n4 3.49141
R634 source.n33 source.n32 3.49141
R635 source.n125 source.n72 3.49141
R636 source.n101 source.n100 3.49141
R637 source.n191 source.n138 3.49141
R638 source.n167 source.n166 3.49141
R639 source.n259 source.n206 3.49141
R640 source.n235 source.n234 3.49141
R641 source.n492 source.n491 2.84303
R642 source.n424 source.n423 2.84303
R643 source.n358 source.n357 2.84303
R644 source.n290 source.n289 2.84303
R645 source.n23 source.n22 2.84303
R646 source.n91 source.n90 2.84303
R647 source.n157 source.n156 2.84303
R648 source.n225 source.n224 2.84303
R649 source.n505 source.n484 2.71565
R650 source.n524 source.n523 2.71565
R651 source.n437 source.n416 2.71565
R652 source.n456 source.n455 2.71565
R653 source.n371 source.n350 2.71565
R654 source.n390 source.n389 2.71565
R655 source.n303 source.n282 2.71565
R656 source.n322 source.n321 2.71565
R657 source.n54 source.n53 2.71565
R658 source.n36 source.n15 2.71565
R659 source.n122 source.n121 2.71565
R660 source.n104 source.n83 2.71565
R661 source.n188 source.n187 2.71565
R662 source.n170 source.n149 2.71565
R663 source.n256 source.n255 2.71565
R664 source.n238 source.n217 2.71565
R665 source.n506 source.n482 1.93989
R666 source.n520 source.n476 1.93989
R667 source.n438 source.n414 1.93989
R668 source.n452 source.n408 1.93989
R669 source.n372 source.n348 1.93989
R670 source.n386 source.n342 1.93989
R671 source.n304 source.n280 1.93989
R672 source.n318 source.n274 1.93989
R673 source.n50 source.n6 1.93989
R674 source.n37 source.n13 1.93989
R675 source.n118 source.n74 1.93989
R676 source.n105 source.n81 1.93989
R677 source.n184 source.n140 1.93989
R678 source.n171 source.n147 1.93989
R679 source.n252 source.n208 1.93989
R680 source.n239 source.n215 1.93989
R681 source.n468 source.t13 1.6505
R682 source.n468 source.t3 1.6505
R683 source.n334 source.t8 1.6505
R684 source.n334 source.t5 1.6505
R685 source.n66 source.t10 1.6505
R686 source.n66 source.t7 1.6505
R687 source.n200 source.t14 1.6505
R688 source.n200 source.t12 1.6505
R689 source.n511 source.n509 1.16414
R690 source.n519 source.n478 1.16414
R691 source.n443 source.n441 1.16414
R692 source.n451 source.n410 1.16414
R693 source.n377 source.n375 1.16414
R694 source.n385 source.n344 1.16414
R695 source.n309 source.n307 1.16414
R696 source.n317 source.n276 1.16414
R697 source.n49 source.n8 1.16414
R698 source.n41 source.n40 1.16414
R699 source.n117 source.n76 1.16414
R700 source.n109 source.n108 1.16414
R701 source.n183 source.n142 1.16414
R702 source.n175 source.n174 1.16414
R703 source.n251 source.n210 1.16414
R704 source.n243 source.n242 1.16414
R705 source.n267 source.n201 0.5005
R706 source.n201 source.n199 0.5005
R707 source.n133 source.n67 0.5005
R708 source.n67 source.n65 0.5005
R709 source.n335 source.n333 0.5005
R710 source.n401 source.n335 0.5005
R711 source.n469 source.n467 0.5005
R712 source.n535 source.n469 0.5005
R713 source.n199 source.n133 0.470328
R714 source.n467 source.n401 0.470328
R715 source.n510 source.n480 0.388379
R716 source.n516 source.n515 0.388379
R717 source.n442 source.n412 0.388379
R718 source.n448 source.n447 0.388379
R719 source.n376 source.n346 0.388379
R720 source.n382 source.n381 0.388379
R721 source.n308 source.n278 0.388379
R722 source.n314 source.n313 0.388379
R723 source.n46 source.n45 0.388379
R724 source.n12 source.n10 0.388379
R725 source.n114 source.n113 0.388379
R726 source.n80 source.n78 0.388379
R727 source.n180 source.n179 0.388379
R728 source.n146 source.n144 0.388379
R729 source.n248 source.n247 0.388379
R730 source.n214 source.n212 0.388379
R731 source source.n536 0.188
R732 source.n492 source.n487 0.155672
R733 source.n499 source.n487 0.155672
R734 source.n500 source.n499 0.155672
R735 source.n500 source.n483 0.155672
R736 source.n507 source.n483 0.155672
R737 source.n508 source.n507 0.155672
R738 source.n508 source.n479 0.155672
R739 source.n517 source.n479 0.155672
R740 source.n518 source.n517 0.155672
R741 source.n518 source.n475 0.155672
R742 source.n525 source.n475 0.155672
R743 source.n526 source.n525 0.155672
R744 source.n526 source.n471 0.155672
R745 source.n533 source.n471 0.155672
R746 source.n424 source.n419 0.155672
R747 source.n431 source.n419 0.155672
R748 source.n432 source.n431 0.155672
R749 source.n432 source.n415 0.155672
R750 source.n439 source.n415 0.155672
R751 source.n440 source.n439 0.155672
R752 source.n440 source.n411 0.155672
R753 source.n449 source.n411 0.155672
R754 source.n450 source.n449 0.155672
R755 source.n450 source.n407 0.155672
R756 source.n457 source.n407 0.155672
R757 source.n458 source.n457 0.155672
R758 source.n458 source.n403 0.155672
R759 source.n465 source.n403 0.155672
R760 source.n358 source.n353 0.155672
R761 source.n365 source.n353 0.155672
R762 source.n366 source.n365 0.155672
R763 source.n366 source.n349 0.155672
R764 source.n373 source.n349 0.155672
R765 source.n374 source.n373 0.155672
R766 source.n374 source.n345 0.155672
R767 source.n383 source.n345 0.155672
R768 source.n384 source.n383 0.155672
R769 source.n384 source.n341 0.155672
R770 source.n391 source.n341 0.155672
R771 source.n392 source.n391 0.155672
R772 source.n392 source.n337 0.155672
R773 source.n399 source.n337 0.155672
R774 source.n290 source.n285 0.155672
R775 source.n297 source.n285 0.155672
R776 source.n298 source.n297 0.155672
R777 source.n298 source.n281 0.155672
R778 source.n305 source.n281 0.155672
R779 source.n306 source.n305 0.155672
R780 source.n306 source.n277 0.155672
R781 source.n315 source.n277 0.155672
R782 source.n316 source.n315 0.155672
R783 source.n316 source.n273 0.155672
R784 source.n323 source.n273 0.155672
R785 source.n324 source.n323 0.155672
R786 source.n324 source.n269 0.155672
R787 source.n331 source.n269 0.155672
R788 source.n63 source.n1 0.155672
R789 source.n56 source.n1 0.155672
R790 source.n56 source.n55 0.155672
R791 source.n55 source.n5 0.155672
R792 source.n48 source.n5 0.155672
R793 source.n48 source.n47 0.155672
R794 source.n47 source.n9 0.155672
R795 source.n39 source.n9 0.155672
R796 source.n39 source.n38 0.155672
R797 source.n38 source.n14 0.155672
R798 source.n31 source.n14 0.155672
R799 source.n31 source.n30 0.155672
R800 source.n30 source.n18 0.155672
R801 source.n23 source.n18 0.155672
R802 source.n131 source.n69 0.155672
R803 source.n124 source.n69 0.155672
R804 source.n124 source.n123 0.155672
R805 source.n123 source.n73 0.155672
R806 source.n116 source.n73 0.155672
R807 source.n116 source.n115 0.155672
R808 source.n115 source.n77 0.155672
R809 source.n107 source.n77 0.155672
R810 source.n107 source.n106 0.155672
R811 source.n106 source.n82 0.155672
R812 source.n99 source.n82 0.155672
R813 source.n99 source.n98 0.155672
R814 source.n98 source.n86 0.155672
R815 source.n91 source.n86 0.155672
R816 source.n197 source.n135 0.155672
R817 source.n190 source.n135 0.155672
R818 source.n190 source.n189 0.155672
R819 source.n189 source.n139 0.155672
R820 source.n182 source.n139 0.155672
R821 source.n182 source.n181 0.155672
R822 source.n181 source.n143 0.155672
R823 source.n173 source.n143 0.155672
R824 source.n173 source.n172 0.155672
R825 source.n172 source.n148 0.155672
R826 source.n165 source.n148 0.155672
R827 source.n165 source.n164 0.155672
R828 source.n164 source.n152 0.155672
R829 source.n157 source.n152 0.155672
R830 source.n265 source.n203 0.155672
R831 source.n258 source.n203 0.155672
R832 source.n258 source.n257 0.155672
R833 source.n257 source.n207 0.155672
R834 source.n250 source.n207 0.155672
R835 source.n250 source.n249 0.155672
R836 source.n249 source.n211 0.155672
R837 source.n241 source.n211 0.155672
R838 source.n241 source.n240 0.155672
R839 source.n240 source.n216 0.155672
R840 source.n233 source.n216 0.155672
R841 source.n233 source.n232 0.155672
R842 source.n232 source.n220 0.155672
R843 source.n225 source.n220 0.155672
R844 drain_left.n5 drain_left.n3 60.0527
R845 drain_left.n2 drain_left.n1 59.7472
R846 drain_left.n2 drain_left.n0 59.7472
R847 drain_left.n5 drain_left.n4 59.5525
R848 drain_left drain_left.n2 29.1171
R849 drain_left drain_left.n5 6.15322
R850 drain_left.n1 drain_left.t2 1.6505
R851 drain_left.n1 drain_left.t1 1.6505
R852 drain_left.n0 drain_left.t0 1.6505
R853 drain_left.n0 drain_left.t4 1.6505
R854 drain_left.n4 drain_left.t3 1.6505
R855 drain_left.n4 drain_left.t7 1.6505
R856 drain_left.n3 drain_left.t5 1.6505
R857 drain_left.n3 drain_left.t6 1.6505
R858 minus.n5 minus.t0 1336.16
R859 minus.n1 minus.t4 1336.16
R860 minus.n12 minus.t5 1336.16
R861 minus.n8 minus.t7 1336.16
R862 minus.n4 minus.t3 1282.12
R863 minus.n2 minus.t1 1282.12
R864 minus.n11 minus.t6 1282.12
R865 minus.n9 minus.t2 1282.12
R866 minus.n1 minus.n0 161.489
R867 minus.n8 minus.n7 161.489
R868 minus.n6 minus.n5 161.3
R869 minus.n3 minus.n0 161.3
R870 minus.n13 minus.n12 161.3
R871 minus.n10 minus.n7 161.3
R872 minus.n4 minus.n3 42.3581
R873 minus.n3 minus.n2 42.3581
R874 minus.n10 minus.n9 42.3581
R875 minus.n11 minus.n10 42.3581
R876 minus.n14 minus.n6 34.0308
R877 minus.n5 minus.n4 30.6732
R878 minus.n2 minus.n1 30.6732
R879 minus.n9 minus.n8 30.6732
R880 minus.n12 minus.n11 30.6732
R881 minus.n14 minus.n13 6.5005
R882 minus.n6 minus.n0 0.189894
R883 minus.n13 minus.n7 0.189894
R884 minus minus.n14 0.188
R885 drain_right.n5 drain_right.n3 60.0525
R886 drain_right.n2 drain_right.n1 59.7472
R887 drain_right.n2 drain_right.n0 59.7472
R888 drain_right.n5 drain_right.n4 59.5527
R889 drain_right drain_right.n2 28.5638
R890 drain_right drain_right.n5 6.15322
R891 drain_right.n1 drain_right.t1 1.6505
R892 drain_right.n1 drain_right.t2 1.6505
R893 drain_right.n0 drain_right.t0 1.6505
R894 drain_right.n0 drain_right.t5 1.6505
R895 drain_right.n3 drain_right.t6 1.6505
R896 drain_right.n3 drain_right.t3 1.6505
R897 drain_right.n4 drain_right.t7 1.6505
R898 drain_right.n4 drain_right.t4 1.6505
C0 plus source 2.55647f
C1 plus minus 4.76613f
C2 drain_right drain_left 0.605638f
C3 drain_left source 17.9349f
C4 minus drain_left 0.170438f
C5 drain_right source 17.9337f
C6 minus drain_right 3.00247f
C7 plus drain_left 3.12447f
C8 minus source 2.54243f
C9 plus drain_right 0.275273f
C10 drain_right a_n1296_n3288# 5.85451f
C11 drain_left a_n1296_n3288# 6.04844f
C12 source a_n1296_n3288# 8.449471f
C13 minus a_n1296_n3288# 4.978832f
C14 plus a_n1296_n3288# 7.05333f
C15 drain_right.t0 a_n1296_n3288# 0.330533f
C16 drain_right.t5 a_n1296_n3288# 0.330533f
C17 drain_right.n0 a_n1296_n3288# 2.9425f
C18 drain_right.t1 a_n1296_n3288# 0.330533f
C19 drain_right.t2 a_n1296_n3288# 0.330533f
C20 drain_right.n1 a_n1296_n3288# 2.9425f
C21 drain_right.n2 a_n1296_n3288# 2.20537f
C22 drain_right.t6 a_n1296_n3288# 0.330533f
C23 drain_right.t3 a_n1296_n3288# 0.330533f
C24 drain_right.n3 a_n1296_n3288# 2.94472f
C25 drain_right.t7 a_n1296_n3288# 0.330533f
C26 drain_right.t4 a_n1296_n3288# 0.330533f
C27 drain_right.n4 a_n1296_n3288# 2.94125f
C28 drain_right.n5 a_n1296_n3288# 1.10795f
C29 minus.n0 a_n1296_n3288# 0.131101f
C30 minus.t0 a_n1296_n3288# 0.491137f
C31 minus.t3 a_n1296_n3288# 0.483097f
C32 minus.t1 a_n1296_n3288# 0.483097f
C33 minus.t4 a_n1296_n3288# 0.491137f
C34 minus.n1 a_n1296_n3288# 0.212548f
C35 minus.n2 a_n1296_n3288# 0.19457f
C36 minus.n3 a_n1296_n3288# 0.021715f
C37 minus.n4 a_n1296_n3288# 0.19457f
C38 minus.n5 a_n1296_n3288# 0.212461f
C39 minus.n6 a_n1296_n3288# 1.82658f
C40 minus.n7 a_n1296_n3288# 0.131101f
C41 minus.t6 a_n1296_n3288# 0.483097f
C42 minus.t2 a_n1296_n3288# 0.483097f
C43 minus.t7 a_n1296_n3288# 0.491137f
C44 minus.n8 a_n1296_n3288# 0.212548f
C45 minus.n9 a_n1296_n3288# 0.19457f
C46 minus.n10 a_n1296_n3288# 0.021715f
C47 minus.n11 a_n1296_n3288# 0.19457f
C48 minus.t5 a_n1296_n3288# 0.491137f
C49 minus.n12 a_n1296_n3288# 0.212461f
C50 minus.n13 a_n1296_n3288# 0.372627f
C51 minus.n14 a_n1296_n3288# 2.23251f
C52 drain_left.t0 a_n1296_n3288# 0.329962f
C53 drain_left.t4 a_n1296_n3288# 0.329962f
C54 drain_left.n0 a_n1296_n3288# 2.93742f
C55 drain_left.t2 a_n1296_n3288# 0.329962f
C56 drain_left.t1 a_n1296_n3288# 0.329962f
C57 drain_left.n1 a_n1296_n3288# 2.93742f
C58 drain_left.n2 a_n1296_n3288# 2.27447f
C59 drain_left.t5 a_n1296_n3288# 0.329962f
C60 drain_left.t6 a_n1296_n3288# 0.329962f
C61 drain_left.n3 a_n1296_n3288# 2.93965f
C62 drain_left.t3 a_n1296_n3288# 0.329962f
C63 drain_left.t7 a_n1296_n3288# 0.329962f
C64 drain_left.n4 a_n1296_n3288# 2.93615f
C65 drain_left.n5 a_n1296_n3288# 1.10603f
C66 source.n0 a_n1296_n3288# 0.033294f
C67 source.n1 a_n1296_n3288# 0.025135f
C68 source.n2 a_n1296_n3288# 0.013506f
C69 source.n3 a_n1296_n3288# 0.031924f
C70 source.n4 a_n1296_n3288# 0.014301f
C71 source.n5 a_n1296_n3288# 0.025135f
C72 source.n6 a_n1296_n3288# 0.013506f
C73 source.n7 a_n1296_n3288# 0.031924f
C74 source.n8 a_n1296_n3288# 0.014301f
C75 source.n9 a_n1296_n3288# 0.025135f
C76 source.n10 a_n1296_n3288# 0.013903f
C77 source.n11 a_n1296_n3288# 0.031924f
C78 source.n12 a_n1296_n3288# 0.013506f
C79 source.n13 a_n1296_n3288# 0.014301f
C80 source.n14 a_n1296_n3288# 0.025135f
C81 source.n15 a_n1296_n3288# 0.013506f
C82 source.n16 a_n1296_n3288# 0.031924f
C83 source.n17 a_n1296_n3288# 0.014301f
C84 source.n18 a_n1296_n3288# 0.025135f
C85 source.n19 a_n1296_n3288# 0.013506f
C86 source.n20 a_n1296_n3288# 0.023943f
C87 source.n21 a_n1296_n3288# 0.022568f
C88 source.t4 a_n1296_n3288# 0.053917f
C89 source.n22 a_n1296_n3288# 0.181217f
C90 source.n23 a_n1296_n3288# 1.26799f
C91 source.n24 a_n1296_n3288# 0.013506f
C92 source.n25 a_n1296_n3288# 0.014301f
C93 source.n26 a_n1296_n3288# 0.031924f
C94 source.n27 a_n1296_n3288# 0.031924f
C95 source.n28 a_n1296_n3288# 0.014301f
C96 source.n29 a_n1296_n3288# 0.013506f
C97 source.n30 a_n1296_n3288# 0.025135f
C98 source.n31 a_n1296_n3288# 0.025135f
C99 source.n32 a_n1296_n3288# 0.013506f
C100 source.n33 a_n1296_n3288# 0.014301f
C101 source.n34 a_n1296_n3288# 0.031924f
C102 source.n35 a_n1296_n3288# 0.031924f
C103 source.n36 a_n1296_n3288# 0.014301f
C104 source.n37 a_n1296_n3288# 0.013506f
C105 source.n38 a_n1296_n3288# 0.025135f
C106 source.n39 a_n1296_n3288# 0.025135f
C107 source.n40 a_n1296_n3288# 0.013506f
C108 source.n41 a_n1296_n3288# 0.014301f
C109 source.n42 a_n1296_n3288# 0.031924f
C110 source.n43 a_n1296_n3288# 0.031924f
C111 source.n44 a_n1296_n3288# 0.031924f
C112 source.n45 a_n1296_n3288# 0.013903f
C113 source.n46 a_n1296_n3288# 0.013506f
C114 source.n47 a_n1296_n3288# 0.025135f
C115 source.n48 a_n1296_n3288# 0.025135f
C116 source.n49 a_n1296_n3288# 0.013506f
C117 source.n50 a_n1296_n3288# 0.014301f
C118 source.n51 a_n1296_n3288# 0.031924f
C119 source.n52 a_n1296_n3288# 0.031924f
C120 source.n53 a_n1296_n3288# 0.014301f
C121 source.n54 a_n1296_n3288# 0.013506f
C122 source.n55 a_n1296_n3288# 0.025135f
C123 source.n56 a_n1296_n3288# 0.025135f
C124 source.n57 a_n1296_n3288# 0.013506f
C125 source.n58 a_n1296_n3288# 0.014301f
C126 source.n59 a_n1296_n3288# 0.031924f
C127 source.n60 a_n1296_n3288# 0.065511f
C128 source.n61 a_n1296_n3288# 0.014301f
C129 source.n62 a_n1296_n3288# 0.013506f
C130 source.n63 a_n1296_n3288# 0.053977f
C131 source.n64 a_n1296_n3288# 0.036155f
C132 source.n65 a_n1296_n3288# 1.00581f
C133 source.t10 a_n1296_n3288# 0.238345f
C134 source.t7 a_n1296_n3288# 0.238345f
C135 source.n66 a_n1296_n3288# 2.04071f
C136 source.n67 a_n1296_n3288# 0.337957f
C137 source.n68 a_n1296_n3288# 0.033294f
C138 source.n69 a_n1296_n3288# 0.025135f
C139 source.n70 a_n1296_n3288# 0.013506f
C140 source.n71 a_n1296_n3288# 0.031924f
C141 source.n72 a_n1296_n3288# 0.014301f
C142 source.n73 a_n1296_n3288# 0.025135f
C143 source.n74 a_n1296_n3288# 0.013506f
C144 source.n75 a_n1296_n3288# 0.031924f
C145 source.n76 a_n1296_n3288# 0.014301f
C146 source.n77 a_n1296_n3288# 0.025135f
C147 source.n78 a_n1296_n3288# 0.013903f
C148 source.n79 a_n1296_n3288# 0.031924f
C149 source.n80 a_n1296_n3288# 0.013506f
C150 source.n81 a_n1296_n3288# 0.014301f
C151 source.n82 a_n1296_n3288# 0.025135f
C152 source.n83 a_n1296_n3288# 0.013506f
C153 source.n84 a_n1296_n3288# 0.031924f
C154 source.n85 a_n1296_n3288# 0.014301f
C155 source.n86 a_n1296_n3288# 0.025135f
C156 source.n87 a_n1296_n3288# 0.013506f
C157 source.n88 a_n1296_n3288# 0.023943f
C158 source.n89 a_n1296_n3288# 0.022568f
C159 source.t9 a_n1296_n3288# 0.053917f
C160 source.n90 a_n1296_n3288# 0.181217f
C161 source.n91 a_n1296_n3288# 1.26799f
C162 source.n92 a_n1296_n3288# 0.013506f
C163 source.n93 a_n1296_n3288# 0.014301f
C164 source.n94 a_n1296_n3288# 0.031924f
C165 source.n95 a_n1296_n3288# 0.031924f
C166 source.n96 a_n1296_n3288# 0.014301f
C167 source.n97 a_n1296_n3288# 0.013506f
C168 source.n98 a_n1296_n3288# 0.025135f
C169 source.n99 a_n1296_n3288# 0.025135f
C170 source.n100 a_n1296_n3288# 0.013506f
C171 source.n101 a_n1296_n3288# 0.014301f
C172 source.n102 a_n1296_n3288# 0.031924f
C173 source.n103 a_n1296_n3288# 0.031924f
C174 source.n104 a_n1296_n3288# 0.014301f
C175 source.n105 a_n1296_n3288# 0.013506f
C176 source.n106 a_n1296_n3288# 0.025135f
C177 source.n107 a_n1296_n3288# 0.025135f
C178 source.n108 a_n1296_n3288# 0.013506f
C179 source.n109 a_n1296_n3288# 0.014301f
C180 source.n110 a_n1296_n3288# 0.031924f
C181 source.n111 a_n1296_n3288# 0.031924f
C182 source.n112 a_n1296_n3288# 0.031924f
C183 source.n113 a_n1296_n3288# 0.013903f
C184 source.n114 a_n1296_n3288# 0.013506f
C185 source.n115 a_n1296_n3288# 0.025135f
C186 source.n116 a_n1296_n3288# 0.025135f
C187 source.n117 a_n1296_n3288# 0.013506f
C188 source.n118 a_n1296_n3288# 0.014301f
C189 source.n119 a_n1296_n3288# 0.031924f
C190 source.n120 a_n1296_n3288# 0.031924f
C191 source.n121 a_n1296_n3288# 0.014301f
C192 source.n122 a_n1296_n3288# 0.013506f
C193 source.n123 a_n1296_n3288# 0.025135f
C194 source.n124 a_n1296_n3288# 0.025135f
C195 source.n125 a_n1296_n3288# 0.013506f
C196 source.n126 a_n1296_n3288# 0.014301f
C197 source.n127 a_n1296_n3288# 0.031924f
C198 source.n128 a_n1296_n3288# 0.065511f
C199 source.n129 a_n1296_n3288# 0.014301f
C200 source.n130 a_n1296_n3288# 0.013506f
C201 source.n131 a_n1296_n3288# 0.053977f
C202 source.n132 a_n1296_n3288# 0.036155f
C203 source.n133 a_n1296_n3288# 0.097691f
C204 source.n134 a_n1296_n3288# 0.033294f
C205 source.n135 a_n1296_n3288# 0.025135f
C206 source.n136 a_n1296_n3288# 0.013506f
C207 source.n137 a_n1296_n3288# 0.031924f
C208 source.n138 a_n1296_n3288# 0.014301f
C209 source.n139 a_n1296_n3288# 0.025135f
C210 source.n140 a_n1296_n3288# 0.013506f
C211 source.n141 a_n1296_n3288# 0.031924f
C212 source.n142 a_n1296_n3288# 0.014301f
C213 source.n143 a_n1296_n3288# 0.025135f
C214 source.n144 a_n1296_n3288# 0.013903f
C215 source.n145 a_n1296_n3288# 0.031924f
C216 source.n146 a_n1296_n3288# 0.013506f
C217 source.n147 a_n1296_n3288# 0.014301f
C218 source.n148 a_n1296_n3288# 0.025135f
C219 source.n149 a_n1296_n3288# 0.013506f
C220 source.n150 a_n1296_n3288# 0.031924f
C221 source.n151 a_n1296_n3288# 0.014301f
C222 source.n152 a_n1296_n3288# 0.025135f
C223 source.n153 a_n1296_n3288# 0.013506f
C224 source.n154 a_n1296_n3288# 0.023943f
C225 source.n155 a_n1296_n3288# 0.022568f
C226 source.t15 a_n1296_n3288# 0.053917f
C227 source.n156 a_n1296_n3288# 0.181217f
C228 source.n157 a_n1296_n3288# 1.26799f
C229 source.n158 a_n1296_n3288# 0.013506f
C230 source.n159 a_n1296_n3288# 0.014301f
C231 source.n160 a_n1296_n3288# 0.031924f
C232 source.n161 a_n1296_n3288# 0.031924f
C233 source.n162 a_n1296_n3288# 0.014301f
C234 source.n163 a_n1296_n3288# 0.013506f
C235 source.n164 a_n1296_n3288# 0.025135f
C236 source.n165 a_n1296_n3288# 0.025135f
C237 source.n166 a_n1296_n3288# 0.013506f
C238 source.n167 a_n1296_n3288# 0.014301f
C239 source.n168 a_n1296_n3288# 0.031924f
C240 source.n169 a_n1296_n3288# 0.031924f
C241 source.n170 a_n1296_n3288# 0.014301f
C242 source.n171 a_n1296_n3288# 0.013506f
C243 source.n172 a_n1296_n3288# 0.025135f
C244 source.n173 a_n1296_n3288# 0.025135f
C245 source.n174 a_n1296_n3288# 0.013506f
C246 source.n175 a_n1296_n3288# 0.014301f
C247 source.n176 a_n1296_n3288# 0.031924f
C248 source.n177 a_n1296_n3288# 0.031924f
C249 source.n178 a_n1296_n3288# 0.031924f
C250 source.n179 a_n1296_n3288# 0.013903f
C251 source.n180 a_n1296_n3288# 0.013506f
C252 source.n181 a_n1296_n3288# 0.025135f
C253 source.n182 a_n1296_n3288# 0.025135f
C254 source.n183 a_n1296_n3288# 0.013506f
C255 source.n184 a_n1296_n3288# 0.014301f
C256 source.n185 a_n1296_n3288# 0.031924f
C257 source.n186 a_n1296_n3288# 0.031924f
C258 source.n187 a_n1296_n3288# 0.014301f
C259 source.n188 a_n1296_n3288# 0.013506f
C260 source.n189 a_n1296_n3288# 0.025135f
C261 source.n190 a_n1296_n3288# 0.025135f
C262 source.n191 a_n1296_n3288# 0.013506f
C263 source.n192 a_n1296_n3288# 0.014301f
C264 source.n193 a_n1296_n3288# 0.031924f
C265 source.n194 a_n1296_n3288# 0.065511f
C266 source.n195 a_n1296_n3288# 0.014301f
C267 source.n196 a_n1296_n3288# 0.013506f
C268 source.n197 a_n1296_n3288# 0.053977f
C269 source.n198 a_n1296_n3288# 0.036155f
C270 source.n199 a_n1296_n3288# 0.097691f
C271 source.t14 a_n1296_n3288# 0.238345f
C272 source.t12 a_n1296_n3288# 0.238345f
C273 source.n200 a_n1296_n3288# 2.04071f
C274 source.n201 a_n1296_n3288# 0.337957f
C275 source.n202 a_n1296_n3288# 0.033294f
C276 source.n203 a_n1296_n3288# 0.025135f
C277 source.n204 a_n1296_n3288# 0.013506f
C278 source.n205 a_n1296_n3288# 0.031924f
C279 source.n206 a_n1296_n3288# 0.014301f
C280 source.n207 a_n1296_n3288# 0.025135f
C281 source.n208 a_n1296_n3288# 0.013506f
C282 source.n209 a_n1296_n3288# 0.031924f
C283 source.n210 a_n1296_n3288# 0.014301f
C284 source.n211 a_n1296_n3288# 0.025135f
C285 source.n212 a_n1296_n3288# 0.013903f
C286 source.n213 a_n1296_n3288# 0.031924f
C287 source.n214 a_n1296_n3288# 0.013506f
C288 source.n215 a_n1296_n3288# 0.014301f
C289 source.n216 a_n1296_n3288# 0.025135f
C290 source.n217 a_n1296_n3288# 0.013506f
C291 source.n218 a_n1296_n3288# 0.031924f
C292 source.n219 a_n1296_n3288# 0.014301f
C293 source.n220 a_n1296_n3288# 0.025135f
C294 source.n221 a_n1296_n3288# 0.013506f
C295 source.n222 a_n1296_n3288# 0.023943f
C296 source.n223 a_n1296_n3288# 0.022568f
C297 source.t1 a_n1296_n3288# 0.053917f
C298 source.n224 a_n1296_n3288# 0.181217f
C299 source.n225 a_n1296_n3288# 1.26799f
C300 source.n226 a_n1296_n3288# 0.013506f
C301 source.n227 a_n1296_n3288# 0.014301f
C302 source.n228 a_n1296_n3288# 0.031924f
C303 source.n229 a_n1296_n3288# 0.031924f
C304 source.n230 a_n1296_n3288# 0.014301f
C305 source.n231 a_n1296_n3288# 0.013506f
C306 source.n232 a_n1296_n3288# 0.025135f
C307 source.n233 a_n1296_n3288# 0.025135f
C308 source.n234 a_n1296_n3288# 0.013506f
C309 source.n235 a_n1296_n3288# 0.014301f
C310 source.n236 a_n1296_n3288# 0.031924f
C311 source.n237 a_n1296_n3288# 0.031924f
C312 source.n238 a_n1296_n3288# 0.014301f
C313 source.n239 a_n1296_n3288# 0.013506f
C314 source.n240 a_n1296_n3288# 0.025135f
C315 source.n241 a_n1296_n3288# 0.025135f
C316 source.n242 a_n1296_n3288# 0.013506f
C317 source.n243 a_n1296_n3288# 0.014301f
C318 source.n244 a_n1296_n3288# 0.031924f
C319 source.n245 a_n1296_n3288# 0.031924f
C320 source.n246 a_n1296_n3288# 0.031924f
C321 source.n247 a_n1296_n3288# 0.013903f
C322 source.n248 a_n1296_n3288# 0.013506f
C323 source.n249 a_n1296_n3288# 0.025135f
C324 source.n250 a_n1296_n3288# 0.025135f
C325 source.n251 a_n1296_n3288# 0.013506f
C326 source.n252 a_n1296_n3288# 0.014301f
C327 source.n253 a_n1296_n3288# 0.031924f
C328 source.n254 a_n1296_n3288# 0.031924f
C329 source.n255 a_n1296_n3288# 0.014301f
C330 source.n256 a_n1296_n3288# 0.013506f
C331 source.n257 a_n1296_n3288# 0.025135f
C332 source.n258 a_n1296_n3288# 0.025135f
C333 source.n259 a_n1296_n3288# 0.013506f
C334 source.n260 a_n1296_n3288# 0.014301f
C335 source.n261 a_n1296_n3288# 0.031924f
C336 source.n262 a_n1296_n3288# 0.065511f
C337 source.n263 a_n1296_n3288# 0.014301f
C338 source.n264 a_n1296_n3288# 0.013506f
C339 source.n265 a_n1296_n3288# 0.053977f
C340 source.n266 a_n1296_n3288# 0.036155f
C341 source.n267 a_n1296_n3288# 1.39978f
C342 source.n268 a_n1296_n3288# 0.033294f
C343 source.n269 a_n1296_n3288# 0.025135f
C344 source.n270 a_n1296_n3288# 0.013506f
C345 source.n271 a_n1296_n3288# 0.031924f
C346 source.n272 a_n1296_n3288# 0.014301f
C347 source.n273 a_n1296_n3288# 0.025135f
C348 source.n274 a_n1296_n3288# 0.013506f
C349 source.n275 a_n1296_n3288# 0.031924f
C350 source.n276 a_n1296_n3288# 0.014301f
C351 source.n277 a_n1296_n3288# 0.025135f
C352 source.n278 a_n1296_n3288# 0.013903f
C353 source.n279 a_n1296_n3288# 0.031924f
C354 source.n280 a_n1296_n3288# 0.014301f
C355 source.n281 a_n1296_n3288# 0.025135f
C356 source.n282 a_n1296_n3288# 0.013506f
C357 source.n283 a_n1296_n3288# 0.031924f
C358 source.n284 a_n1296_n3288# 0.014301f
C359 source.n285 a_n1296_n3288# 0.025135f
C360 source.n286 a_n1296_n3288# 0.013506f
C361 source.n287 a_n1296_n3288# 0.023943f
C362 source.n288 a_n1296_n3288# 0.022568f
C363 source.t11 a_n1296_n3288# 0.053917f
C364 source.n289 a_n1296_n3288# 0.181217f
C365 source.n290 a_n1296_n3288# 1.26799f
C366 source.n291 a_n1296_n3288# 0.013506f
C367 source.n292 a_n1296_n3288# 0.014301f
C368 source.n293 a_n1296_n3288# 0.031924f
C369 source.n294 a_n1296_n3288# 0.031924f
C370 source.n295 a_n1296_n3288# 0.014301f
C371 source.n296 a_n1296_n3288# 0.013506f
C372 source.n297 a_n1296_n3288# 0.025135f
C373 source.n298 a_n1296_n3288# 0.025135f
C374 source.n299 a_n1296_n3288# 0.013506f
C375 source.n300 a_n1296_n3288# 0.014301f
C376 source.n301 a_n1296_n3288# 0.031924f
C377 source.n302 a_n1296_n3288# 0.031924f
C378 source.n303 a_n1296_n3288# 0.014301f
C379 source.n304 a_n1296_n3288# 0.013506f
C380 source.n305 a_n1296_n3288# 0.025135f
C381 source.n306 a_n1296_n3288# 0.025135f
C382 source.n307 a_n1296_n3288# 0.013506f
C383 source.n308 a_n1296_n3288# 0.013506f
C384 source.n309 a_n1296_n3288# 0.014301f
C385 source.n310 a_n1296_n3288# 0.031924f
C386 source.n311 a_n1296_n3288# 0.031924f
C387 source.n312 a_n1296_n3288# 0.031924f
C388 source.n313 a_n1296_n3288# 0.013903f
C389 source.n314 a_n1296_n3288# 0.013506f
C390 source.n315 a_n1296_n3288# 0.025135f
C391 source.n316 a_n1296_n3288# 0.025135f
C392 source.n317 a_n1296_n3288# 0.013506f
C393 source.n318 a_n1296_n3288# 0.014301f
C394 source.n319 a_n1296_n3288# 0.031924f
C395 source.n320 a_n1296_n3288# 0.031924f
C396 source.n321 a_n1296_n3288# 0.014301f
C397 source.n322 a_n1296_n3288# 0.013506f
C398 source.n323 a_n1296_n3288# 0.025135f
C399 source.n324 a_n1296_n3288# 0.025135f
C400 source.n325 a_n1296_n3288# 0.013506f
C401 source.n326 a_n1296_n3288# 0.014301f
C402 source.n327 a_n1296_n3288# 0.031924f
C403 source.n328 a_n1296_n3288# 0.065511f
C404 source.n329 a_n1296_n3288# 0.014301f
C405 source.n330 a_n1296_n3288# 0.013506f
C406 source.n331 a_n1296_n3288# 0.053977f
C407 source.n332 a_n1296_n3288# 0.036155f
C408 source.n333 a_n1296_n3288# 1.39978f
C409 source.t8 a_n1296_n3288# 0.238345f
C410 source.t5 a_n1296_n3288# 0.238345f
C411 source.n334 a_n1296_n3288# 2.0407f
C412 source.n335 a_n1296_n3288# 0.33797f
C413 source.n336 a_n1296_n3288# 0.033294f
C414 source.n337 a_n1296_n3288# 0.025135f
C415 source.n338 a_n1296_n3288# 0.013506f
C416 source.n339 a_n1296_n3288# 0.031924f
C417 source.n340 a_n1296_n3288# 0.014301f
C418 source.n341 a_n1296_n3288# 0.025135f
C419 source.n342 a_n1296_n3288# 0.013506f
C420 source.n343 a_n1296_n3288# 0.031924f
C421 source.n344 a_n1296_n3288# 0.014301f
C422 source.n345 a_n1296_n3288# 0.025135f
C423 source.n346 a_n1296_n3288# 0.013903f
C424 source.n347 a_n1296_n3288# 0.031924f
C425 source.n348 a_n1296_n3288# 0.014301f
C426 source.n349 a_n1296_n3288# 0.025135f
C427 source.n350 a_n1296_n3288# 0.013506f
C428 source.n351 a_n1296_n3288# 0.031924f
C429 source.n352 a_n1296_n3288# 0.014301f
C430 source.n353 a_n1296_n3288# 0.025135f
C431 source.n354 a_n1296_n3288# 0.013506f
C432 source.n355 a_n1296_n3288# 0.023943f
C433 source.n356 a_n1296_n3288# 0.022568f
C434 source.t6 a_n1296_n3288# 0.053917f
C435 source.n357 a_n1296_n3288# 0.181217f
C436 source.n358 a_n1296_n3288# 1.26799f
C437 source.n359 a_n1296_n3288# 0.013506f
C438 source.n360 a_n1296_n3288# 0.014301f
C439 source.n361 a_n1296_n3288# 0.031924f
C440 source.n362 a_n1296_n3288# 0.031924f
C441 source.n363 a_n1296_n3288# 0.014301f
C442 source.n364 a_n1296_n3288# 0.013506f
C443 source.n365 a_n1296_n3288# 0.025135f
C444 source.n366 a_n1296_n3288# 0.025135f
C445 source.n367 a_n1296_n3288# 0.013506f
C446 source.n368 a_n1296_n3288# 0.014301f
C447 source.n369 a_n1296_n3288# 0.031924f
C448 source.n370 a_n1296_n3288# 0.031924f
C449 source.n371 a_n1296_n3288# 0.014301f
C450 source.n372 a_n1296_n3288# 0.013506f
C451 source.n373 a_n1296_n3288# 0.025135f
C452 source.n374 a_n1296_n3288# 0.025135f
C453 source.n375 a_n1296_n3288# 0.013506f
C454 source.n376 a_n1296_n3288# 0.013506f
C455 source.n377 a_n1296_n3288# 0.014301f
C456 source.n378 a_n1296_n3288# 0.031924f
C457 source.n379 a_n1296_n3288# 0.031924f
C458 source.n380 a_n1296_n3288# 0.031924f
C459 source.n381 a_n1296_n3288# 0.013903f
C460 source.n382 a_n1296_n3288# 0.013506f
C461 source.n383 a_n1296_n3288# 0.025135f
C462 source.n384 a_n1296_n3288# 0.025135f
C463 source.n385 a_n1296_n3288# 0.013506f
C464 source.n386 a_n1296_n3288# 0.014301f
C465 source.n387 a_n1296_n3288# 0.031924f
C466 source.n388 a_n1296_n3288# 0.031924f
C467 source.n389 a_n1296_n3288# 0.014301f
C468 source.n390 a_n1296_n3288# 0.013506f
C469 source.n391 a_n1296_n3288# 0.025135f
C470 source.n392 a_n1296_n3288# 0.025135f
C471 source.n393 a_n1296_n3288# 0.013506f
C472 source.n394 a_n1296_n3288# 0.014301f
C473 source.n395 a_n1296_n3288# 0.031924f
C474 source.n396 a_n1296_n3288# 0.065511f
C475 source.n397 a_n1296_n3288# 0.014301f
C476 source.n398 a_n1296_n3288# 0.013506f
C477 source.n399 a_n1296_n3288# 0.053977f
C478 source.n400 a_n1296_n3288# 0.036155f
C479 source.n401 a_n1296_n3288# 0.097691f
C480 source.n402 a_n1296_n3288# 0.033294f
C481 source.n403 a_n1296_n3288# 0.025135f
C482 source.n404 a_n1296_n3288# 0.013506f
C483 source.n405 a_n1296_n3288# 0.031924f
C484 source.n406 a_n1296_n3288# 0.014301f
C485 source.n407 a_n1296_n3288# 0.025135f
C486 source.n408 a_n1296_n3288# 0.013506f
C487 source.n409 a_n1296_n3288# 0.031924f
C488 source.n410 a_n1296_n3288# 0.014301f
C489 source.n411 a_n1296_n3288# 0.025135f
C490 source.n412 a_n1296_n3288# 0.013903f
C491 source.n413 a_n1296_n3288# 0.031924f
C492 source.n414 a_n1296_n3288# 0.014301f
C493 source.n415 a_n1296_n3288# 0.025135f
C494 source.n416 a_n1296_n3288# 0.013506f
C495 source.n417 a_n1296_n3288# 0.031924f
C496 source.n418 a_n1296_n3288# 0.014301f
C497 source.n419 a_n1296_n3288# 0.025135f
C498 source.n420 a_n1296_n3288# 0.013506f
C499 source.n421 a_n1296_n3288# 0.023943f
C500 source.n422 a_n1296_n3288# 0.022568f
C501 source.t2 a_n1296_n3288# 0.053917f
C502 source.n423 a_n1296_n3288# 0.181217f
C503 source.n424 a_n1296_n3288# 1.26799f
C504 source.n425 a_n1296_n3288# 0.013506f
C505 source.n426 a_n1296_n3288# 0.014301f
C506 source.n427 a_n1296_n3288# 0.031924f
C507 source.n428 a_n1296_n3288# 0.031924f
C508 source.n429 a_n1296_n3288# 0.014301f
C509 source.n430 a_n1296_n3288# 0.013506f
C510 source.n431 a_n1296_n3288# 0.025135f
C511 source.n432 a_n1296_n3288# 0.025135f
C512 source.n433 a_n1296_n3288# 0.013506f
C513 source.n434 a_n1296_n3288# 0.014301f
C514 source.n435 a_n1296_n3288# 0.031924f
C515 source.n436 a_n1296_n3288# 0.031924f
C516 source.n437 a_n1296_n3288# 0.014301f
C517 source.n438 a_n1296_n3288# 0.013506f
C518 source.n439 a_n1296_n3288# 0.025135f
C519 source.n440 a_n1296_n3288# 0.025135f
C520 source.n441 a_n1296_n3288# 0.013506f
C521 source.n442 a_n1296_n3288# 0.013506f
C522 source.n443 a_n1296_n3288# 0.014301f
C523 source.n444 a_n1296_n3288# 0.031924f
C524 source.n445 a_n1296_n3288# 0.031924f
C525 source.n446 a_n1296_n3288# 0.031924f
C526 source.n447 a_n1296_n3288# 0.013903f
C527 source.n448 a_n1296_n3288# 0.013506f
C528 source.n449 a_n1296_n3288# 0.025135f
C529 source.n450 a_n1296_n3288# 0.025135f
C530 source.n451 a_n1296_n3288# 0.013506f
C531 source.n452 a_n1296_n3288# 0.014301f
C532 source.n453 a_n1296_n3288# 0.031924f
C533 source.n454 a_n1296_n3288# 0.031924f
C534 source.n455 a_n1296_n3288# 0.014301f
C535 source.n456 a_n1296_n3288# 0.013506f
C536 source.n457 a_n1296_n3288# 0.025135f
C537 source.n458 a_n1296_n3288# 0.025135f
C538 source.n459 a_n1296_n3288# 0.013506f
C539 source.n460 a_n1296_n3288# 0.014301f
C540 source.n461 a_n1296_n3288# 0.031924f
C541 source.n462 a_n1296_n3288# 0.065511f
C542 source.n463 a_n1296_n3288# 0.014301f
C543 source.n464 a_n1296_n3288# 0.013506f
C544 source.n465 a_n1296_n3288# 0.053977f
C545 source.n466 a_n1296_n3288# 0.036155f
C546 source.n467 a_n1296_n3288# 0.097691f
C547 source.t13 a_n1296_n3288# 0.238345f
C548 source.t3 a_n1296_n3288# 0.238345f
C549 source.n468 a_n1296_n3288# 2.0407f
C550 source.n469 a_n1296_n3288# 0.33797f
C551 source.n470 a_n1296_n3288# 0.033294f
C552 source.n471 a_n1296_n3288# 0.025135f
C553 source.n472 a_n1296_n3288# 0.013506f
C554 source.n473 a_n1296_n3288# 0.031924f
C555 source.n474 a_n1296_n3288# 0.014301f
C556 source.n475 a_n1296_n3288# 0.025135f
C557 source.n476 a_n1296_n3288# 0.013506f
C558 source.n477 a_n1296_n3288# 0.031924f
C559 source.n478 a_n1296_n3288# 0.014301f
C560 source.n479 a_n1296_n3288# 0.025135f
C561 source.n480 a_n1296_n3288# 0.013903f
C562 source.n481 a_n1296_n3288# 0.031924f
C563 source.n482 a_n1296_n3288# 0.014301f
C564 source.n483 a_n1296_n3288# 0.025135f
C565 source.n484 a_n1296_n3288# 0.013506f
C566 source.n485 a_n1296_n3288# 0.031924f
C567 source.n486 a_n1296_n3288# 0.014301f
C568 source.n487 a_n1296_n3288# 0.025135f
C569 source.n488 a_n1296_n3288# 0.013506f
C570 source.n489 a_n1296_n3288# 0.023943f
C571 source.n490 a_n1296_n3288# 0.022568f
C572 source.t0 a_n1296_n3288# 0.053917f
C573 source.n491 a_n1296_n3288# 0.181217f
C574 source.n492 a_n1296_n3288# 1.26799f
C575 source.n493 a_n1296_n3288# 0.013506f
C576 source.n494 a_n1296_n3288# 0.014301f
C577 source.n495 a_n1296_n3288# 0.031924f
C578 source.n496 a_n1296_n3288# 0.031924f
C579 source.n497 a_n1296_n3288# 0.014301f
C580 source.n498 a_n1296_n3288# 0.013506f
C581 source.n499 a_n1296_n3288# 0.025135f
C582 source.n500 a_n1296_n3288# 0.025135f
C583 source.n501 a_n1296_n3288# 0.013506f
C584 source.n502 a_n1296_n3288# 0.014301f
C585 source.n503 a_n1296_n3288# 0.031924f
C586 source.n504 a_n1296_n3288# 0.031924f
C587 source.n505 a_n1296_n3288# 0.014301f
C588 source.n506 a_n1296_n3288# 0.013506f
C589 source.n507 a_n1296_n3288# 0.025135f
C590 source.n508 a_n1296_n3288# 0.025135f
C591 source.n509 a_n1296_n3288# 0.013506f
C592 source.n510 a_n1296_n3288# 0.013506f
C593 source.n511 a_n1296_n3288# 0.014301f
C594 source.n512 a_n1296_n3288# 0.031924f
C595 source.n513 a_n1296_n3288# 0.031924f
C596 source.n514 a_n1296_n3288# 0.031924f
C597 source.n515 a_n1296_n3288# 0.013903f
C598 source.n516 a_n1296_n3288# 0.013506f
C599 source.n517 a_n1296_n3288# 0.025135f
C600 source.n518 a_n1296_n3288# 0.025135f
C601 source.n519 a_n1296_n3288# 0.013506f
C602 source.n520 a_n1296_n3288# 0.014301f
C603 source.n521 a_n1296_n3288# 0.031924f
C604 source.n522 a_n1296_n3288# 0.031924f
C605 source.n523 a_n1296_n3288# 0.014301f
C606 source.n524 a_n1296_n3288# 0.013506f
C607 source.n525 a_n1296_n3288# 0.025135f
C608 source.n526 a_n1296_n3288# 0.025135f
C609 source.n527 a_n1296_n3288# 0.013506f
C610 source.n528 a_n1296_n3288# 0.014301f
C611 source.n529 a_n1296_n3288# 0.031924f
C612 source.n530 a_n1296_n3288# 0.065511f
C613 source.n531 a_n1296_n3288# 0.014301f
C614 source.n532 a_n1296_n3288# 0.013506f
C615 source.n533 a_n1296_n3288# 0.053977f
C616 source.n534 a_n1296_n3288# 0.036155f
C617 source.n535 a_n1296_n3288# 0.236781f
C618 source.n536 a_n1296_n3288# 1.57484f
C619 plus.n0 a_n1296_n3288# 0.135159f
C620 plus.t4 a_n1296_n3288# 0.49805f
C621 plus.t1 a_n1296_n3288# 0.49805f
C622 plus.t2 a_n1296_n3288# 0.506339f
C623 plus.n1 a_n1296_n3288# 0.219126f
C624 plus.n2 a_n1296_n3288# 0.200592f
C625 plus.n3 a_n1296_n3288# 0.022387f
C626 plus.n4 a_n1296_n3288# 0.200592f
C627 plus.t0 a_n1296_n3288# 0.506339f
C628 plus.n5 a_n1296_n3288# 0.219037f
C629 plus.n6 a_n1296_n3288# 0.657392f
C630 plus.n7 a_n1296_n3288# 0.135159f
C631 plus.t7 a_n1296_n3288# 0.506339f
C632 plus.t3 a_n1296_n3288# 0.49805f
C633 plus.t5 a_n1296_n3288# 0.49805f
C634 plus.t6 a_n1296_n3288# 0.506339f
C635 plus.n8 a_n1296_n3288# 0.219126f
C636 plus.n9 a_n1296_n3288# 0.200592f
C637 plus.n10 a_n1296_n3288# 0.022387f
C638 plus.n11 a_n1296_n3288# 0.200592f
C639 plus.n12 a_n1296_n3288# 0.219037f
C640 plus.n13 a_n1296_n3288# 1.58632f
.ends

