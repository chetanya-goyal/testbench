* NGSPICE file created from diffpair283.ext - technology: sky130A

.subckt diffpair283 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t11 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X1 source.t14 minus.t1 drain_right.t6 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X2 source.t12 minus.t2 drain_right.t5 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X3 source.t4 plus.t0 drain_left.t7 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X4 a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X5 drain_right.t4 minus.t3 source.t13 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X6 drain_left.t6 plus.t1 source.t7 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X7 a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X8 drain_left.t5 plus.t2 source.t5 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X9 source.t6 plus.t3 drain_left.t4 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X10 drain_right.t3 minus.t4 source.t9 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X11 source.t2 plus.t4 drain_left.t3 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X12 drain_left.t2 plus.t5 source.t3 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X13 drain_right.t2 minus.t5 source.t8 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X14 source.t10 minus.t6 drain_right.t1 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X15 source.t15 minus.t7 drain_right.t0 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X16 a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X17 a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X18 source.t1 plus.t6 drain_left.t1 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X19 drain_left.t0 plus.t7 source.t0 a_n1546_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
R0 minus.n2 minus.t4 388.748
R1 minus.n10 minus.t6 388.748
R2 minus.n1 minus.t2 367.767
R3 minus.n5 minus.t3 367.767
R4 minus.n6 minus.t7 367.767
R5 minus.n9 minus.t5 367.767
R6 minus.n13 minus.t1 367.767
R7 minus.n14 minus.t0 367.767
R8 minus.n7 minus.n6 161.3
R9 minus.n5 minus.n0 161.3
R10 minus.n4 minus.n3 161.3
R11 minus.n15 minus.n14 161.3
R12 minus.n13 minus.n8 161.3
R13 minus.n12 minus.n11 161.3
R14 minus.n3 minus.n2 70.4033
R15 minus.n11 minus.n10 70.4033
R16 minus.n6 minus.n5 48.2005
R17 minus.n14 minus.n13 48.2005
R18 minus.n16 minus.n7 30.527
R19 minus.n5 minus.n4 24.1005
R20 minus.n4 minus.n1 24.1005
R21 minus.n12 minus.n9 24.1005
R22 minus.n13 minus.n12 24.1005
R23 minus.n2 minus.n1 20.9576
R24 minus.n10 minus.n9 20.9576
R25 minus.n16 minus.n15 6.5952
R26 minus.n7 minus.n0 0.189894
R27 minus.n3 minus.n0 0.189894
R28 minus.n11 minus.n8 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 source.n258 source.n232 289.615
R32 source.n224 source.n198 289.615
R33 source.n192 source.n166 289.615
R34 source.n158 source.n132 289.615
R35 source.n26 source.n0 289.615
R36 source.n60 source.n34 289.615
R37 source.n92 source.n66 289.615
R38 source.n126 source.n100 289.615
R39 source.n243 source.n242 185
R40 source.n240 source.n239 185
R41 source.n249 source.n248 185
R42 source.n251 source.n250 185
R43 source.n236 source.n235 185
R44 source.n257 source.n256 185
R45 source.n259 source.n258 185
R46 source.n209 source.n208 185
R47 source.n206 source.n205 185
R48 source.n215 source.n214 185
R49 source.n217 source.n216 185
R50 source.n202 source.n201 185
R51 source.n223 source.n222 185
R52 source.n225 source.n224 185
R53 source.n177 source.n176 185
R54 source.n174 source.n173 185
R55 source.n183 source.n182 185
R56 source.n185 source.n184 185
R57 source.n170 source.n169 185
R58 source.n191 source.n190 185
R59 source.n193 source.n192 185
R60 source.n143 source.n142 185
R61 source.n140 source.n139 185
R62 source.n149 source.n148 185
R63 source.n151 source.n150 185
R64 source.n136 source.n135 185
R65 source.n157 source.n156 185
R66 source.n159 source.n158 185
R67 source.n27 source.n26 185
R68 source.n25 source.n24 185
R69 source.n4 source.n3 185
R70 source.n19 source.n18 185
R71 source.n17 source.n16 185
R72 source.n8 source.n7 185
R73 source.n11 source.n10 185
R74 source.n61 source.n60 185
R75 source.n59 source.n58 185
R76 source.n38 source.n37 185
R77 source.n53 source.n52 185
R78 source.n51 source.n50 185
R79 source.n42 source.n41 185
R80 source.n45 source.n44 185
R81 source.n93 source.n92 185
R82 source.n91 source.n90 185
R83 source.n70 source.n69 185
R84 source.n85 source.n84 185
R85 source.n83 source.n82 185
R86 source.n74 source.n73 185
R87 source.n77 source.n76 185
R88 source.n127 source.n126 185
R89 source.n125 source.n124 185
R90 source.n104 source.n103 185
R91 source.n119 source.n118 185
R92 source.n117 source.n116 185
R93 source.n108 source.n107 185
R94 source.n111 source.n110 185
R95 source.t11 source.n241 147.661
R96 source.t10 source.n207 147.661
R97 source.t5 source.n175 147.661
R98 source.t2 source.n141 147.661
R99 source.t7 source.n9 147.661
R100 source.t4 source.n43 147.661
R101 source.t9 source.n75 147.661
R102 source.t15 source.n109 147.661
R103 source.n242 source.n239 104.615
R104 source.n249 source.n239 104.615
R105 source.n250 source.n249 104.615
R106 source.n250 source.n235 104.615
R107 source.n257 source.n235 104.615
R108 source.n258 source.n257 104.615
R109 source.n208 source.n205 104.615
R110 source.n215 source.n205 104.615
R111 source.n216 source.n215 104.615
R112 source.n216 source.n201 104.615
R113 source.n223 source.n201 104.615
R114 source.n224 source.n223 104.615
R115 source.n176 source.n173 104.615
R116 source.n183 source.n173 104.615
R117 source.n184 source.n183 104.615
R118 source.n184 source.n169 104.615
R119 source.n191 source.n169 104.615
R120 source.n192 source.n191 104.615
R121 source.n142 source.n139 104.615
R122 source.n149 source.n139 104.615
R123 source.n150 source.n149 104.615
R124 source.n150 source.n135 104.615
R125 source.n157 source.n135 104.615
R126 source.n158 source.n157 104.615
R127 source.n26 source.n25 104.615
R128 source.n25 source.n3 104.615
R129 source.n18 source.n3 104.615
R130 source.n18 source.n17 104.615
R131 source.n17 source.n7 104.615
R132 source.n10 source.n7 104.615
R133 source.n60 source.n59 104.615
R134 source.n59 source.n37 104.615
R135 source.n52 source.n37 104.615
R136 source.n52 source.n51 104.615
R137 source.n51 source.n41 104.615
R138 source.n44 source.n41 104.615
R139 source.n92 source.n91 104.615
R140 source.n91 source.n69 104.615
R141 source.n84 source.n69 104.615
R142 source.n84 source.n83 104.615
R143 source.n83 source.n73 104.615
R144 source.n76 source.n73 104.615
R145 source.n126 source.n125 104.615
R146 source.n125 source.n103 104.615
R147 source.n118 source.n103 104.615
R148 source.n118 source.n117 104.615
R149 source.n117 source.n107 104.615
R150 source.n110 source.n107 104.615
R151 source.n242 source.t11 52.3082
R152 source.n208 source.t10 52.3082
R153 source.n176 source.t5 52.3082
R154 source.n142 source.t2 52.3082
R155 source.n10 source.t7 52.3082
R156 source.n44 source.t4 52.3082
R157 source.n76 source.t9 52.3082
R158 source.n110 source.t15 52.3082
R159 source.n33 source.n32 50.512
R160 source.n99 source.n98 50.512
R161 source.n231 source.n230 50.5119
R162 source.n165 source.n164 50.5119
R163 source.n263 source.n262 32.1853
R164 source.n229 source.n228 32.1853
R165 source.n197 source.n196 32.1853
R166 source.n163 source.n162 32.1853
R167 source.n31 source.n30 32.1853
R168 source.n65 source.n64 32.1853
R169 source.n97 source.n96 32.1853
R170 source.n131 source.n130 32.1853
R171 source.n163 source.n131 17.4578
R172 source.n243 source.n241 15.6674
R173 source.n209 source.n207 15.6674
R174 source.n177 source.n175 15.6674
R175 source.n143 source.n141 15.6674
R176 source.n11 source.n9 15.6674
R177 source.n45 source.n43 15.6674
R178 source.n77 source.n75 15.6674
R179 source.n111 source.n109 15.6674
R180 source.n244 source.n240 12.8005
R181 source.n210 source.n206 12.8005
R182 source.n178 source.n174 12.8005
R183 source.n144 source.n140 12.8005
R184 source.n12 source.n8 12.8005
R185 source.n46 source.n42 12.8005
R186 source.n78 source.n74 12.8005
R187 source.n112 source.n108 12.8005
R188 source.n248 source.n247 12.0247
R189 source.n214 source.n213 12.0247
R190 source.n182 source.n181 12.0247
R191 source.n148 source.n147 12.0247
R192 source.n16 source.n15 12.0247
R193 source.n50 source.n49 12.0247
R194 source.n82 source.n81 12.0247
R195 source.n116 source.n115 12.0247
R196 source.n264 source.n31 11.8371
R197 source.n251 source.n238 11.249
R198 source.n217 source.n204 11.249
R199 source.n185 source.n172 11.249
R200 source.n151 source.n138 11.249
R201 source.n19 source.n6 11.249
R202 source.n53 source.n40 11.249
R203 source.n85 source.n72 11.249
R204 source.n119 source.n106 11.249
R205 source.n252 source.n236 10.4732
R206 source.n218 source.n202 10.4732
R207 source.n186 source.n170 10.4732
R208 source.n152 source.n136 10.4732
R209 source.n20 source.n4 10.4732
R210 source.n54 source.n38 10.4732
R211 source.n86 source.n70 10.4732
R212 source.n120 source.n104 10.4732
R213 source.n256 source.n255 9.69747
R214 source.n222 source.n221 9.69747
R215 source.n190 source.n189 9.69747
R216 source.n156 source.n155 9.69747
R217 source.n24 source.n23 9.69747
R218 source.n58 source.n57 9.69747
R219 source.n90 source.n89 9.69747
R220 source.n124 source.n123 9.69747
R221 source.n262 source.n261 9.45567
R222 source.n228 source.n227 9.45567
R223 source.n196 source.n195 9.45567
R224 source.n162 source.n161 9.45567
R225 source.n30 source.n29 9.45567
R226 source.n64 source.n63 9.45567
R227 source.n96 source.n95 9.45567
R228 source.n130 source.n129 9.45567
R229 source.n261 source.n260 9.3005
R230 source.n234 source.n233 9.3005
R231 source.n255 source.n254 9.3005
R232 source.n253 source.n252 9.3005
R233 source.n238 source.n237 9.3005
R234 source.n247 source.n246 9.3005
R235 source.n245 source.n244 9.3005
R236 source.n227 source.n226 9.3005
R237 source.n200 source.n199 9.3005
R238 source.n221 source.n220 9.3005
R239 source.n219 source.n218 9.3005
R240 source.n204 source.n203 9.3005
R241 source.n213 source.n212 9.3005
R242 source.n211 source.n210 9.3005
R243 source.n195 source.n194 9.3005
R244 source.n168 source.n167 9.3005
R245 source.n189 source.n188 9.3005
R246 source.n187 source.n186 9.3005
R247 source.n172 source.n171 9.3005
R248 source.n181 source.n180 9.3005
R249 source.n179 source.n178 9.3005
R250 source.n161 source.n160 9.3005
R251 source.n134 source.n133 9.3005
R252 source.n155 source.n154 9.3005
R253 source.n153 source.n152 9.3005
R254 source.n138 source.n137 9.3005
R255 source.n147 source.n146 9.3005
R256 source.n145 source.n144 9.3005
R257 source.n29 source.n28 9.3005
R258 source.n2 source.n1 9.3005
R259 source.n23 source.n22 9.3005
R260 source.n21 source.n20 9.3005
R261 source.n6 source.n5 9.3005
R262 source.n15 source.n14 9.3005
R263 source.n13 source.n12 9.3005
R264 source.n63 source.n62 9.3005
R265 source.n36 source.n35 9.3005
R266 source.n57 source.n56 9.3005
R267 source.n55 source.n54 9.3005
R268 source.n40 source.n39 9.3005
R269 source.n49 source.n48 9.3005
R270 source.n47 source.n46 9.3005
R271 source.n95 source.n94 9.3005
R272 source.n68 source.n67 9.3005
R273 source.n89 source.n88 9.3005
R274 source.n87 source.n86 9.3005
R275 source.n72 source.n71 9.3005
R276 source.n81 source.n80 9.3005
R277 source.n79 source.n78 9.3005
R278 source.n129 source.n128 9.3005
R279 source.n102 source.n101 9.3005
R280 source.n123 source.n122 9.3005
R281 source.n121 source.n120 9.3005
R282 source.n106 source.n105 9.3005
R283 source.n115 source.n114 9.3005
R284 source.n113 source.n112 9.3005
R285 source.n259 source.n234 8.92171
R286 source.n225 source.n200 8.92171
R287 source.n193 source.n168 8.92171
R288 source.n159 source.n134 8.92171
R289 source.n27 source.n2 8.92171
R290 source.n61 source.n36 8.92171
R291 source.n93 source.n68 8.92171
R292 source.n127 source.n102 8.92171
R293 source.n260 source.n232 8.14595
R294 source.n226 source.n198 8.14595
R295 source.n194 source.n166 8.14595
R296 source.n160 source.n132 8.14595
R297 source.n28 source.n0 8.14595
R298 source.n62 source.n34 8.14595
R299 source.n94 source.n66 8.14595
R300 source.n128 source.n100 8.14595
R301 source.n262 source.n232 5.81868
R302 source.n228 source.n198 5.81868
R303 source.n196 source.n166 5.81868
R304 source.n162 source.n132 5.81868
R305 source.n30 source.n0 5.81868
R306 source.n64 source.n34 5.81868
R307 source.n96 source.n66 5.81868
R308 source.n130 source.n100 5.81868
R309 source.n264 source.n263 5.62119
R310 source.n260 source.n259 5.04292
R311 source.n226 source.n225 5.04292
R312 source.n194 source.n193 5.04292
R313 source.n160 source.n159 5.04292
R314 source.n28 source.n27 5.04292
R315 source.n62 source.n61 5.04292
R316 source.n94 source.n93 5.04292
R317 source.n128 source.n127 5.04292
R318 source.n245 source.n241 4.38594
R319 source.n211 source.n207 4.38594
R320 source.n179 source.n175 4.38594
R321 source.n145 source.n141 4.38594
R322 source.n13 source.n9 4.38594
R323 source.n47 source.n43 4.38594
R324 source.n79 source.n75 4.38594
R325 source.n113 source.n109 4.38594
R326 source.n256 source.n234 4.26717
R327 source.n222 source.n200 4.26717
R328 source.n190 source.n168 4.26717
R329 source.n156 source.n134 4.26717
R330 source.n24 source.n2 4.26717
R331 source.n58 source.n36 4.26717
R332 source.n90 source.n68 4.26717
R333 source.n124 source.n102 4.26717
R334 source.n255 source.n236 3.49141
R335 source.n221 source.n202 3.49141
R336 source.n189 source.n170 3.49141
R337 source.n155 source.n136 3.49141
R338 source.n23 source.n4 3.49141
R339 source.n57 source.n38 3.49141
R340 source.n89 source.n70 3.49141
R341 source.n123 source.n104 3.49141
R342 source.n230 source.t8 3.3005
R343 source.n230 source.t14 3.3005
R344 source.n164 source.t0 3.3005
R345 source.n164 source.t6 3.3005
R346 source.n32 source.t3 3.3005
R347 source.n32 source.t1 3.3005
R348 source.n98 source.t13 3.3005
R349 source.n98 source.t12 3.3005
R350 source.n252 source.n251 2.71565
R351 source.n218 source.n217 2.71565
R352 source.n186 source.n185 2.71565
R353 source.n152 source.n151 2.71565
R354 source.n20 source.n19 2.71565
R355 source.n54 source.n53 2.71565
R356 source.n86 source.n85 2.71565
R357 source.n120 source.n119 2.71565
R358 source.n248 source.n238 1.93989
R359 source.n214 source.n204 1.93989
R360 source.n182 source.n172 1.93989
R361 source.n148 source.n138 1.93989
R362 source.n16 source.n6 1.93989
R363 source.n50 source.n40 1.93989
R364 source.n82 source.n72 1.93989
R365 source.n116 source.n106 1.93989
R366 source.n247 source.n240 1.16414
R367 source.n213 source.n206 1.16414
R368 source.n181 source.n174 1.16414
R369 source.n147 source.n140 1.16414
R370 source.n15 source.n8 1.16414
R371 source.n49 source.n42 1.16414
R372 source.n81 source.n74 1.16414
R373 source.n115 source.n108 1.16414
R374 source.n131 source.n99 0.716017
R375 source.n99 source.n97 0.716017
R376 source.n65 source.n33 0.716017
R377 source.n33 source.n31 0.716017
R378 source.n165 source.n163 0.716017
R379 source.n197 source.n165 0.716017
R380 source.n231 source.n229 0.716017
R381 source.n263 source.n231 0.716017
R382 source.n97 source.n65 0.470328
R383 source.n229 source.n197 0.470328
R384 source.n244 source.n243 0.388379
R385 source.n210 source.n209 0.388379
R386 source.n178 source.n177 0.388379
R387 source.n144 source.n143 0.388379
R388 source.n12 source.n11 0.388379
R389 source.n46 source.n45 0.388379
R390 source.n78 source.n77 0.388379
R391 source.n112 source.n111 0.388379
R392 source source.n264 0.188
R393 source.n246 source.n245 0.155672
R394 source.n246 source.n237 0.155672
R395 source.n253 source.n237 0.155672
R396 source.n254 source.n253 0.155672
R397 source.n254 source.n233 0.155672
R398 source.n261 source.n233 0.155672
R399 source.n212 source.n211 0.155672
R400 source.n212 source.n203 0.155672
R401 source.n219 source.n203 0.155672
R402 source.n220 source.n219 0.155672
R403 source.n220 source.n199 0.155672
R404 source.n227 source.n199 0.155672
R405 source.n180 source.n179 0.155672
R406 source.n180 source.n171 0.155672
R407 source.n187 source.n171 0.155672
R408 source.n188 source.n187 0.155672
R409 source.n188 source.n167 0.155672
R410 source.n195 source.n167 0.155672
R411 source.n146 source.n145 0.155672
R412 source.n146 source.n137 0.155672
R413 source.n153 source.n137 0.155672
R414 source.n154 source.n153 0.155672
R415 source.n154 source.n133 0.155672
R416 source.n161 source.n133 0.155672
R417 source.n29 source.n1 0.155672
R418 source.n22 source.n1 0.155672
R419 source.n22 source.n21 0.155672
R420 source.n21 source.n5 0.155672
R421 source.n14 source.n5 0.155672
R422 source.n14 source.n13 0.155672
R423 source.n63 source.n35 0.155672
R424 source.n56 source.n35 0.155672
R425 source.n56 source.n55 0.155672
R426 source.n55 source.n39 0.155672
R427 source.n48 source.n39 0.155672
R428 source.n48 source.n47 0.155672
R429 source.n95 source.n67 0.155672
R430 source.n88 source.n67 0.155672
R431 source.n88 source.n87 0.155672
R432 source.n87 source.n71 0.155672
R433 source.n80 source.n71 0.155672
R434 source.n80 source.n79 0.155672
R435 source.n129 source.n101 0.155672
R436 source.n122 source.n101 0.155672
R437 source.n122 source.n121 0.155672
R438 source.n121 source.n105 0.155672
R439 source.n114 source.n105 0.155672
R440 source.n114 source.n113 0.155672
R441 drain_right.n5 drain_right.n3 67.9062
R442 drain_right.n2 drain_right.n1 67.4931
R443 drain_right.n2 drain_right.n0 67.4931
R444 drain_right.n5 drain_right.n4 67.1908
R445 drain_right drain_right.n2 24.7727
R446 drain_right drain_right.n5 6.36873
R447 drain_right.n1 drain_right.t6 3.3005
R448 drain_right.n1 drain_right.t7 3.3005
R449 drain_right.n0 drain_right.t1 3.3005
R450 drain_right.n0 drain_right.t2 3.3005
R451 drain_right.n3 drain_right.t5 3.3005
R452 drain_right.n3 drain_right.t3 3.3005
R453 drain_right.n4 drain_right.t0 3.3005
R454 drain_right.n4 drain_right.t4 3.3005
R455 plus.n2 plus.t0 388.748
R456 plus.n10 plus.t2 388.748
R457 plus.n6 plus.t1 367.767
R458 plus.n5 plus.t6 367.767
R459 plus.n1 plus.t5 367.767
R460 plus.n14 plus.t4 367.767
R461 plus.n13 plus.t7 367.767
R462 plus.n9 plus.t3 367.767
R463 plus.n4 plus.n3 161.3
R464 plus.n5 plus.n0 161.3
R465 plus.n7 plus.n6 161.3
R466 plus.n12 plus.n11 161.3
R467 plus.n13 plus.n8 161.3
R468 plus.n15 plus.n14 161.3
R469 plus.n3 plus.n2 70.4033
R470 plus.n11 plus.n10 70.4033
R471 plus.n6 plus.n5 48.2005
R472 plus.n14 plus.n13 48.2005
R473 plus plus.n15 26.6808
R474 plus.n4 plus.n1 24.1005
R475 plus.n5 plus.n4 24.1005
R476 plus.n13 plus.n12 24.1005
R477 plus.n12 plus.n9 24.1005
R478 plus.n2 plus.n1 20.9576
R479 plus.n10 plus.n9 20.9576
R480 plus plus.n7 9.96641
R481 plus.n3 plus.n0 0.189894
R482 plus.n7 plus.n0 0.189894
R483 plus.n15 plus.n8 0.189894
R484 plus.n11 plus.n8 0.189894
R485 drain_left.n5 drain_left.n3 67.9063
R486 drain_left.n2 drain_left.n1 67.4931
R487 drain_left.n2 drain_left.n0 67.4931
R488 drain_left.n5 drain_left.n4 67.1907
R489 drain_left drain_left.n2 25.3259
R490 drain_left drain_left.n5 6.36873
R491 drain_left.n1 drain_left.t4 3.3005
R492 drain_left.n1 drain_left.t5 3.3005
R493 drain_left.n0 drain_left.t3 3.3005
R494 drain_left.n0 drain_left.t0 3.3005
R495 drain_left.n4 drain_left.t1 3.3005
R496 drain_left.n4 drain_left.t6 3.3005
R497 drain_left.n3 drain_left.t7 3.3005
R498 drain_left.n3 drain_left.t2 3.3005
C0 minus source 2.45219f
C1 drain_right minus 2.47803f
C2 source plus 2.46621f
C3 drain_right plus 0.302201f
C4 minus plus 3.96056f
C5 drain_left source 7.538579f
C6 drain_right drain_left 0.727126f
C7 drain_left minus 0.171215f
C8 drain_right source 7.53907f
C9 drain_left plus 2.62605f
C10 drain_right a_n1546_n2088# 4.37594f
C11 drain_left a_n1546_n2088# 4.60434f
C12 source a_n1546_n2088# 5.280389f
C13 minus a_n1546_n2088# 5.489971f
C14 plus a_n1546_n2088# 6.96934f
C15 drain_left.t3 a_n1546_n2088# 0.133651f
C16 drain_left.t0 a_n1546_n2088# 0.133651f
C17 drain_left.n0 a_n1546_n2088# 1.11615f
C18 drain_left.t4 a_n1546_n2088# 0.133651f
C19 drain_left.t5 a_n1546_n2088# 0.133651f
C20 drain_left.n1 a_n1546_n2088# 1.11615f
C21 drain_left.n2 a_n1546_n2088# 1.60702f
C22 drain_left.t7 a_n1546_n2088# 0.133651f
C23 drain_left.t2 a_n1546_n2088# 0.133651f
C24 drain_left.n3 a_n1546_n2088# 1.11855f
C25 drain_left.t1 a_n1546_n2088# 0.133651f
C26 drain_left.t6 a_n1546_n2088# 0.133651f
C27 drain_left.n4 a_n1546_n2088# 1.11465f
C28 drain_left.n5 a_n1546_n2088# 0.967151f
C29 plus.n0 a_n1546_n2088# 0.051362f
C30 plus.t1 a_n1546_n2088# 0.446931f
C31 plus.t6 a_n1546_n2088# 0.446931f
C32 plus.t5 a_n1546_n2088# 0.446931f
C33 plus.n1 a_n1546_n2088# 0.215756f
C34 plus.t0 a_n1546_n2088# 0.458298f
C35 plus.n2 a_n1546_n2088# 0.19956f
C36 plus.n3 a_n1546_n2088# 0.169205f
C37 plus.n4 a_n1546_n2088# 0.011655f
C38 plus.n5 a_n1546_n2088# 0.215756f
C39 plus.n6 a_n1546_n2088# 0.210531f
C40 plus.n7 a_n1546_n2088# 0.45209f
C41 plus.n8 a_n1546_n2088# 0.051362f
C42 plus.t4 a_n1546_n2088# 0.446931f
C43 plus.t7 a_n1546_n2088# 0.446931f
C44 plus.t3 a_n1546_n2088# 0.446931f
C45 plus.n9 a_n1546_n2088# 0.215756f
C46 plus.t2 a_n1546_n2088# 0.458298f
C47 plus.n10 a_n1546_n2088# 0.19956f
C48 plus.n11 a_n1546_n2088# 0.169205f
C49 plus.n12 a_n1546_n2088# 0.011655f
C50 plus.n13 a_n1546_n2088# 0.215756f
C51 plus.n14 a_n1546_n2088# 0.210531f
C52 plus.n15 a_n1546_n2088# 1.24877f
C53 drain_right.t1 a_n1546_n2088# 0.133788f
C54 drain_right.t2 a_n1546_n2088# 0.133788f
C55 drain_right.n0 a_n1546_n2088# 1.1173f
C56 drain_right.t6 a_n1546_n2088# 0.133788f
C57 drain_right.t7 a_n1546_n2088# 0.133788f
C58 drain_right.n1 a_n1546_n2088# 1.1173f
C59 drain_right.n2 a_n1546_n2088# 1.5511f
C60 drain_right.t5 a_n1546_n2088# 0.133788f
C61 drain_right.t3 a_n1546_n2088# 0.133788f
C62 drain_right.n3 a_n1546_n2088# 1.1197f
C63 drain_right.t0 a_n1546_n2088# 0.133788f
C64 drain_right.t4 a_n1546_n2088# 0.133788f
C65 drain_right.n4 a_n1546_n2088# 1.1158f
C66 drain_right.n5 a_n1546_n2088# 0.968145f
C67 source.n0 a_n1546_n2088# 0.031854f
C68 source.n1 a_n1546_n2088# 0.022663f
C69 source.n2 a_n1546_n2088# 0.012178f
C70 source.n3 a_n1546_n2088# 0.028784f
C71 source.n4 a_n1546_n2088# 0.012894f
C72 source.n5 a_n1546_n2088# 0.022663f
C73 source.n6 a_n1546_n2088# 0.012178f
C74 source.n7 a_n1546_n2088# 0.028784f
C75 source.n8 a_n1546_n2088# 0.012894f
C76 source.n9 a_n1546_n2088# 0.09698f
C77 source.t7 a_n1546_n2088# 0.046914f
C78 source.n10 a_n1546_n2088# 0.021588f
C79 source.n11 a_n1546_n2088# 0.017003f
C80 source.n12 a_n1546_n2088# 0.012178f
C81 source.n13 a_n1546_n2088# 0.539234f
C82 source.n14 a_n1546_n2088# 0.022663f
C83 source.n15 a_n1546_n2088# 0.012178f
C84 source.n16 a_n1546_n2088# 0.012894f
C85 source.n17 a_n1546_n2088# 0.028784f
C86 source.n18 a_n1546_n2088# 0.028784f
C87 source.n19 a_n1546_n2088# 0.012894f
C88 source.n20 a_n1546_n2088# 0.012178f
C89 source.n21 a_n1546_n2088# 0.022663f
C90 source.n22 a_n1546_n2088# 0.022663f
C91 source.n23 a_n1546_n2088# 0.012178f
C92 source.n24 a_n1546_n2088# 0.012894f
C93 source.n25 a_n1546_n2088# 0.028784f
C94 source.n26 a_n1546_n2088# 0.062313f
C95 source.n27 a_n1546_n2088# 0.012894f
C96 source.n28 a_n1546_n2088# 0.012178f
C97 source.n29 a_n1546_n2088# 0.052383f
C98 source.n30 a_n1546_n2088# 0.034866f
C99 source.n31 a_n1546_n2088# 0.5705f
C100 source.t3 a_n1546_n2088# 0.107452f
C101 source.t1 a_n1546_n2088# 0.107452f
C102 source.n32 a_n1546_n2088# 0.836845f
C103 source.n33 a_n1546_n2088# 0.31694f
C104 source.n34 a_n1546_n2088# 0.031854f
C105 source.n35 a_n1546_n2088# 0.022663f
C106 source.n36 a_n1546_n2088# 0.012178f
C107 source.n37 a_n1546_n2088# 0.028784f
C108 source.n38 a_n1546_n2088# 0.012894f
C109 source.n39 a_n1546_n2088# 0.022663f
C110 source.n40 a_n1546_n2088# 0.012178f
C111 source.n41 a_n1546_n2088# 0.028784f
C112 source.n42 a_n1546_n2088# 0.012894f
C113 source.n43 a_n1546_n2088# 0.09698f
C114 source.t4 a_n1546_n2088# 0.046914f
C115 source.n44 a_n1546_n2088# 0.021588f
C116 source.n45 a_n1546_n2088# 0.017003f
C117 source.n46 a_n1546_n2088# 0.012178f
C118 source.n47 a_n1546_n2088# 0.539234f
C119 source.n48 a_n1546_n2088# 0.022663f
C120 source.n49 a_n1546_n2088# 0.012178f
C121 source.n50 a_n1546_n2088# 0.012894f
C122 source.n51 a_n1546_n2088# 0.028784f
C123 source.n52 a_n1546_n2088# 0.028784f
C124 source.n53 a_n1546_n2088# 0.012894f
C125 source.n54 a_n1546_n2088# 0.012178f
C126 source.n55 a_n1546_n2088# 0.022663f
C127 source.n56 a_n1546_n2088# 0.022663f
C128 source.n57 a_n1546_n2088# 0.012178f
C129 source.n58 a_n1546_n2088# 0.012894f
C130 source.n59 a_n1546_n2088# 0.028784f
C131 source.n60 a_n1546_n2088# 0.062313f
C132 source.n61 a_n1546_n2088# 0.012894f
C133 source.n62 a_n1546_n2088# 0.012178f
C134 source.n63 a_n1546_n2088# 0.052383f
C135 source.n64 a_n1546_n2088# 0.034866f
C136 source.n65 a_n1546_n2088# 0.105914f
C137 source.n66 a_n1546_n2088# 0.031854f
C138 source.n67 a_n1546_n2088# 0.022663f
C139 source.n68 a_n1546_n2088# 0.012178f
C140 source.n69 a_n1546_n2088# 0.028784f
C141 source.n70 a_n1546_n2088# 0.012894f
C142 source.n71 a_n1546_n2088# 0.022663f
C143 source.n72 a_n1546_n2088# 0.012178f
C144 source.n73 a_n1546_n2088# 0.028784f
C145 source.n74 a_n1546_n2088# 0.012894f
C146 source.n75 a_n1546_n2088# 0.09698f
C147 source.t9 a_n1546_n2088# 0.046914f
C148 source.n76 a_n1546_n2088# 0.021588f
C149 source.n77 a_n1546_n2088# 0.017003f
C150 source.n78 a_n1546_n2088# 0.012178f
C151 source.n79 a_n1546_n2088# 0.539234f
C152 source.n80 a_n1546_n2088# 0.022663f
C153 source.n81 a_n1546_n2088# 0.012178f
C154 source.n82 a_n1546_n2088# 0.012894f
C155 source.n83 a_n1546_n2088# 0.028784f
C156 source.n84 a_n1546_n2088# 0.028784f
C157 source.n85 a_n1546_n2088# 0.012894f
C158 source.n86 a_n1546_n2088# 0.012178f
C159 source.n87 a_n1546_n2088# 0.022663f
C160 source.n88 a_n1546_n2088# 0.022663f
C161 source.n89 a_n1546_n2088# 0.012178f
C162 source.n90 a_n1546_n2088# 0.012894f
C163 source.n91 a_n1546_n2088# 0.028784f
C164 source.n92 a_n1546_n2088# 0.062313f
C165 source.n93 a_n1546_n2088# 0.012894f
C166 source.n94 a_n1546_n2088# 0.012178f
C167 source.n95 a_n1546_n2088# 0.052383f
C168 source.n96 a_n1546_n2088# 0.034866f
C169 source.n97 a_n1546_n2088# 0.105914f
C170 source.t13 a_n1546_n2088# 0.107452f
C171 source.t12 a_n1546_n2088# 0.107452f
C172 source.n98 a_n1546_n2088# 0.836845f
C173 source.n99 a_n1546_n2088# 0.31694f
C174 source.n100 a_n1546_n2088# 0.031854f
C175 source.n101 a_n1546_n2088# 0.022663f
C176 source.n102 a_n1546_n2088# 0.012178f
C177 source.n103 a_n1546_n2088# 0.028784f
C178 source.n104 a_n1546_n2088# 0.012894f
C179 source.n105 a_n1546_n2088# 0.022663f
C180 source.n106 a_n1546_n2088# 0.012178f
C181 source.n107 a_n1546_n2088# 0.028784f
C182 source.n108 a_n1546_n2088# 0.012894f
C183 source.n109 a_n1546_n2088# 0.09698f
C184 source.t15 a_n1546_n2088# 0.046914f
C185 source.n110 a_n1546_n2088# 0.021588f
C186 source.n111 a_n1546_n2088# 0.017003f
C187 source.n112 a_n1546_n2088# 0.012178f
C188 source.n113 a_n1546_n2088# 0.539234f
C189 source.n114 a_n1546_n2088# 0.022663f
C190 source.n115 a_n1546_n2088# 0.012178f
C191 source.n116 a_n1546_n2088# 0.012894f
C192 source.n117 a_n1546_n2088# 0.028784f
C193 source.n118 a_n1546_n2088# 0.028784f
C194 source.n119 a_n1546_n2088# 0.012894f
C195 source.n120 a_n1546_n2088# 0.012178f
C196 source.n121 a_n1546_n2088# 0.022663f
C197 source.n122 a_n1546_n2088# 0.022663f
C198 source.n123 a_n1546_n2088# 0.012178f
C199 source.n124 a_n1546_n2088# 0.012894f
C200 source.n125 a_n1546_n2088# 0.028784f
C201 source.n126 a_n1546_n2088# 0.062313f
C202 source.n127 a_n1546_n2088# 0.012894f
C203 source.n128 a_n1546_n2088# 0.012178f
C204 source.n129 a_n1546_n2088# 0.052383f
C205 source.n130 a_n1546_n2088# 0.034866f
C206 source.n131 a_n1546_n2088# 0.865871f
C207 source.n132 a_n1546_n2088# 0.031854f
C208 source.n133 a_n1546_n2088# 0.022663f
C209 source.n134 a_n1546_n2088# 0.012178f
C210 source.n135 a_n1546_n2088# 0.028784f
C211 source.n136 a_n1546_n2088# 0.012894f
C212 source.n137 a_n1546_n2088# 0.022663f
C213 source.n138 a_n1546_n2088# 0.012178f
C214 source.n139 a_n1546_n2088# 0.028784f
C215 source.n140 a_n1546_n2088# 0.012894f
C216 source.n141 a_n1546_n2088# 0.09698f
C217 source.t2 a_n1546_n2088# 0.046914f
C218 source.n142 a_n1546_n2088# 0.021588f
C219 source.n143 a_n1546_n2088# 0.017003f
C220 source.n144 a_n1546_n2088# 0.012178f
C221 source.n145 a_n1546_n2088# 0.539234f
C222 source.n146 a_n1546_n2088# 0.022663f
C223 source.n147 a_n1546_n2088# 0.012178f
C224 source.n148 a_n1546_n2088# 0.012894f
C225 source.n149 a_n1546_n2088# 0.028784f
C226 source.n150 a_n1546_n2088# 0.028784f
C227 source.n151 a_n1546_n2088# 0.012894f
C228 source.n152 a_n1546_n2088# 0.012178f
C229 source.n153 a_n1546_n2088# 0.022663f
C230 source.n154 a_n1546_n2088# 0.022663f
C231 source.n155 a_n1546_n2088# 0.012178f
C232 source.n156 a_n1546_n2088# 0.012894f
C233 source.n157 a_n1546_n2088# 0.028784f
C234 source.n158 a_n1546_n2088# 0.062313f
C235 source.n159 a_n1546_n2088# 0.012894f
C236 source.n160 a_n1546_n2088# 0.012178f
C237 source.n161 a_n1546_n2088# 0.052383f
C238 source.n162 a_n1546_n2088# 0.034866f
C239 source.n163 a_n1546_n2088# 0.865871f
C240 source.t0 a_n1546_n2088# 0.107452f
C241 source.t6 a_n1546_n2088# 0.107452f
C242 source.n164 a_n1546_n2088# 0.836839f
C243 source.n165 a_n1546_n2088# 0.316946f
C244 source.n166 a_n1546_n2088# 0.031854f
C245 source.n167 a_n1546_n2088# 0.022663f
C246 source.n168 a_n1546_n2088# 0.012178f
C247 source.n169 a_n1546_n2088# 0.028784f
C248 source.n170 a_n1546_n2088# 0.012894f
C249 source.n171 a_n1546_n2088# 0.022663f
C250 source.n172 a_n1546_n2088# 0.012178f
C251 source.n173 a_n1546_n2088# 0.028784f
C252 source.n174 a_n1546_n2088# 0.012894f
C253 source.n175 a_n1546_n2088# 0.09698f
C254 source.t5 a_n1546_n2088# 0.046914f
C255 source.n176 a_n1546_n2088# 0.021588f
C256 source.n177 a_n1546_n2088# 0.017003f
C257 source.n178 a_n1546_n2088# 0.012178f
C258 source.n179 a_n1546_n2088# 0.539234f
C259 source.n180 a_n1546_n2088# 0.022663f
C260 source.n181 a_n1546_n2088# 0.012178f
C261 source.n182 a_n1546_n2088# 0.012894f
C262 source.n183 a_n1546_n2088# 0.028784f
C263 source.n184 a_n1546_n2088# 0.028784f
C264 source.n185 a_n1546_n2088# 0.012894f
C265 source.n186 a_n1546_n2088# 0.012178f
C266 source.n187 a_n1546_n2088# 0.022663f
C267 source.n188 a_n1546_n2088# 0.022663f
C268 source.n189 a_n1546_n2088# 0.012178f
C269 source.n190 a_n1546_n2088# 0.012894f
C270 source.n191 a_n1546_n2088# 0.028784f
C271 source.n192 a_n1546_n2088# 0.062313f
C272 source.n193 a_n1546_n2088# 0.012894f
C273 source.n194 a_n1546_n2088# 0.012178f
C274 source.n195 a_n1546_n2088# 0.052383f
C275 source.n196 a_n1546_n2088# 0.034866f
C276 source.n197 a_n1546_n2088# 0.105914f
C277 source.n198 a_n1546_n2088# 0.031854f
C278 source.n199 a_n1546_n2088# 0.022663f
C279 source.n200 a_n1546_n2088# 0.012178f
C280 source.n201 a_n1546_n2088# 0.028784f
C281 source.n202 a_n1546_n2088# 0.012894f
C282 source.n203 a_n1546_n2088# 0.022663f
C283 source.n204 a_n1546_n2088# 0.012178f
C284 source.n205 a_n1546_n2088# 0.028784f
C285 source.n206 a_n1546_n2088# 0.012894f
C286 source.n207 a_n1546_n2088# 0.09698f
C287 source.t10 a_n1546_n2088# 0.046914f
C288 source.n208 a_n1546_n2088# 0.021588f
C289 source.n209 a_n1546_n2088# 0.017003f
C290 source.n210 a_n1546_n2088# 0.012178f
C291 source.n211 a_n1546_n2088# 0.539234f
C292 source.n212 a_n1546_n2088# 0.022663f
C293 source.n213 a_n1546_n2088# 0.012178f
C294 source.n214 a_n1546_n2088# 0.012894f
C295 source.n215 a_n1546_n2088# 0.028784f
C296 source.n216 a_n1546_n2088# 0.028784f
C297 source.n217 a_n1546_n2088# 0.012894f
C298 source.n218 a_n1546_n2088# 0.012178f
C299 source.n219 a_n1546_n2088# 0.022663f
C300 source.n220 a_n1546_n2088# 0.022663f
C301 source.n221 a_n1546_n2088# 0.012178f
C302 source.n222 a_n1546_n2088# 0.012894f
C303 source.n223 a_n1546_n2088# 0.028784f
C304 source.n224 a_n1546_n2088# 0.062313f
C305 source.n225 a_n1546_n2088# 0.012894f
C306 source.n226 a_n1546_n2088# 0.012178f
C307 source.n227 a_n1546_n2088# 0.052383f
C308 source.n228 a_n1546_n2088# 0.034866f
C309 source.n229 a_n1546_n2088# 0.105914f
C310 source.t8 a_n1546_n2088# 0.107452f
C311 source.t14 a_n1546_n2088# 0.107452f
C312 source.n230 a_n1546_n2088# 0.836839f
C313 source.n231 a_n1546_n2088# 0.316946f
C314 source.n232 a_n1546_n2088# 0.031854f
C315 source.n233 a_n1546_n2088# 0.022663f
C316 source.n234 a_n1546_n2088# 0.012178f
C317 source.n235 a_n1546_n2088# 0.028784f
C318 source.n236 a_n1546_n2088# 0.012894f
C319 source.n237 a_n1546_n2088# 0.022663f
C320 source.n238 a_n1546_n2088# 0.012178f
C321 source.n239 a_n1546_n2088# 0.028784f
C322 source.n240 a_n1546_n2088# 0.012894f
C323 source.n241 a_n1546_n2088# 0.09698f
C324 source.t11 a_n1546_n2088# 0.046914f
C325 source.n242 a_n1546_n2088# 0.021588f
C326 source.n243 a_n1546_n2088# 0.017003f
C327 source.n244 a_n1546_n2088# 0.012178f
C328 source.n245 a_n1546_n2088# 0.539234f
C329 source.n246 a_n1546_n2088# 0.022663f
C330 source.n247 a_n1546_n2088# 0.012178f
C331 source.n248 a_n1546_n2088# 0.012894f
C332 source.n249 a_n1546_n2088# 0.028784f
C333 source.n250 a_n1546_n2088# 0.028784f
C334 source.n251 a_n1546_n2088# 0.012894f
C335 source.n252 a_n1546_n2088# 0.012178f
C336 source.n253 a_n1546_n2088# 0.022663f
C337 source.n254 a_n1546_n2088# 0.022663f
C338 source.n255 a_n1546_n2088# 0.012178f
C339 source.n256 a_n1546_n2088# 0.012894f
C340 source.n257 a_n1546_n2088# 0.028784f
C341 source.n258 a_n1546_n2088# 0.062313f
C342 source.n259 a_n1546_n2088# 0.012894f
C343 source.n260 a_n1546_n2088# 0.012178f
C344 source.n261 a_n1546_n2088# 0.052383f
C345 source.n262 a_n1546_n2088# 0.034866f
C346 source.n263 a_n1546_n2088# 0.24385f
C347 source.n264 a_n1546_n2088# 0.933512f
C348 minus.n0 a_n1546_n2088# 0.050224f
C349 minus.t2 a_n1546_n2088# 0.437031f
C350 minus.n1 a_n1546_n2088# 0.210977f
C351 minus.t4 a_n1546_n2088# 0.448147f
C352 minus.n2 a_n1546_n2088# 0.19514f
C353 minus.n3 a_n1546_n2088# 0.165457f
C354 minus.n4 a_n1546_n2088# 0.011397f
C355 minus.t3 a_n1546_n2088# 0.437031f
C356 minus.n5 a_n1546_n2088# 0.210977f
C357 minus.t7 a_n1546_n2088# 0.437031f
C358 minus.n6 a_n1546_n2088# 0.205868f
C359 minus.n7 a_n1546_n2088# 1.35017f
C360 minus.n8 a_n1546_n2088# 0.050224f
C361 minus.t5 a_n1546_n2088# 0.437031f
C362 minus.n9 a_n1546_n2088# 0.210977f
C363 minus.t6 a_n1546_n2088# 0.448147f
C364 minus.n10 a_n1546_n2088# 0.19514f
C365 minus.n11 a_n1546_n2088# 0.165457f
C366 minus.n12 a_n1546_n2088# 0.011397f
C367 minus.t1 a_n1546_n2088# 0.437031f
C368 minus.n13 a_n1546_n2088# 0.210977f
C369 minus.t0 a_n1546_n2088# 0.437031f
C370 minus.n14 a_n1546_n2088# 0.205868f
C371 minus.n15 a_n1546_n2088# 0.339564f
C372 minus.n16 a_n1546_n2088# 1.65873f
.ends

