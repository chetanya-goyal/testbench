* NGSPICE file created from diffpair190.ext - technology: sky130A

.subckt diffpair190 minus drain_right drain_left source plus
X0 drain_right minus source a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.3
X1 a_n968_n1492# a_n968_n1492# a_n968_n1492# a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X2 a_n968_n1492# a_n968_n1492# a_n968_n1492# a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X3 a_n968_n1492# a_n968_n1492# a_n968_n1492# a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X4 drain_left plus source a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.3
X5 drain_left plus source a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.3
X6 a_n968_n1492# a_n968_n1492# a_n968_n1492# a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X7 drain_right minus source a_n968_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.3
.ends

