* NGSPICE file created from diffpair534.ext - technology: sky130A

.subckt diffpair534 minus drain_right drain_left source plus
X0 a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.6
X1 source.t14 minus.t0 drain_right.t7 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X2 drain_left.t9 plus.t0 source.t19 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X3 source.t0 plus.t1 drain_left.t8 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X4 drain_right.t4 minus.t1 source.t13 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X5 drain_left.t7 plus.t2 source.t3 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X6 a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X7 drain_right.t9 minus.t2 source.t12 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X8 source.t11 minus.t3 drain_right.t6 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X9 drain_left.t6 plus.t3 source.t17 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X10 source.t10 minus.t4 drain_right.t0 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X11 drain_right.t1 minus.t5 source.t9 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X12 drain_right.t5 minus.t6 source.t8 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X13 source.t4 plus.t4 drain_left.t5 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X14 source.t16 plus.t5 drain_left.t4 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X15 source.t7 minus.t7 drain_right.t3 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X16 drain_left.t3 plus.t6 source.t1 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X17 drain_right.t8 minus.t8 source.t6 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X18 source.t2 plus.t7 drain_left.t2 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X19 drain_left.t1 plus.t8 source.t15 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X20 a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X21 drain_right.t2 minus.t9 source.t5 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X22 a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X23 drain_left.t0 plus.t9 source.t18 a_n1832_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
R0 minus.n3 minus.t8 694.173
R1 minus.n13 minus.t9 694.173
R2 minus.n2 minus.t7 667.972
R3 minus.n1 minus.t5 667.972
R4 minus.n6 minus.t4 667.972
R5 minus.n8 minus.t1 667.972
R6 minus.n12 minus.t3 667.972
R7 minus.n11 minus.t6 667.972
R8 minus.n16 minus.t0 667.972
R9 minus.n18 minus.t2 667.972
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n6 minus.n5 161.3
R13 minus.n19 minus.n18 161.3
R14 minus.n17 minus.n10 161.3
R15 minus.n16 minus.n15 161.3
R16 minus.n4 minus.n1 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n8 minus.n7 45.2793
R23 minus.n18 minus.n17 45.2793
R24 minus.n4 minus.n3 45.1669
R25 minus.n14 minus.n13 45.1669
R26 minus.n20 minus.n9 38.4342
R27 minus.n3 minus.n2 14.3992
R28 minus.n13 minus.n12 14.3992
R29 minus.n20 minus.n19 6.60088
R30 minus.n7 minus.n6 2.92171
R31 minus.n17 minus.n16 2.92171
R32 minus.n5 minus.n4 0.285035
R33 minus.n15 minus.n14 0.285035
R34 minus.n9 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n15 minus.n10 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 drain_right.n1 drain_right.t2 63.0013
R40 drain_right.n7 drain_right.t4 62.1998
R41 drain_right.n6 drain_right.n4 61.6814
R42 drain_right.n3 drain_right.n2 61.4255
R43 drain_right.n6 drain_right.n5 60.8798
R44 drain_right.n1 drain_right.n0 60.8796
R45 drain_right drain_right.n3 32.4939
R46 drain_right drain_right.n7 6.05408
R47 drain_right.n2 drain_right.t7 1.3205
R48 drain_right.n2 drain_right.t9 1.3205
R49 drain_right.n0 drain_right.t6 1.3205
R50 drain_right.n0 drain_right.t5 1.3205
R51 drain_right.n4 drain_right.t3 1.3205
R52 drain_right.n4 drain_right.t8 1.3205
R53 drain_right.n5 drain_right.t0 1.3205
R54 drain_right.n5 drain_right.t1 1.3205
R55 drain_right.n7 drain_right.n6 0.802224
R56 drain_right.n3 drain_right.n1 0.145585
R57 source.n5 source.t6 45.521
R58 source.n19 source.t12 45.5208
R59 source.n14 source.t19 45.5208
R60 source.n0 source.t17 45.5208
R61 source.n2 source.n1 44.201
R62 source.n4 source.n3 44.201
R63 source.n7 source.n6 44.201
R64 source.n9 source.n8 44.201
R65 source.n18 source.n17 44.2008
R66 source.n16 source.n15 44.2008
R67 source.n13 source.n12 44.2008
R68 source.n11 source.n10 44.2008
R69 source.n11 source.n9 25.1639
R70 source.n20 source.n0 18.6984
R71 source.n20 source.n19 5.66429
R72 source.n17 source.t8 1.3205
R73 source.n17 source.t14 1.3205
R74 source.n15 source.t5 1.3205
R75 source.n15 source.t11 1.3205
R76 source.n12 source.t18 1.3205
R77 source.n12 source.t4 1.3205
R78 source.n10 source.t3 1.3205
R79 source.n10 source.t0 1.3205
R80 source.n1 source.t1 1.3205
R81 source.n1 source.t16 1.3205
R82 source.n3 source.t15 1.3205
R83 source.n3 source.t2 1.3205
R84 source.n6 source.t9 1.3205
R85 source.n6 source.t7 1.3205
R86 source.n8 source.t13 1.3205
R87 source.n8 source.t10 1.3205
R88 source.n5 source.n4 0.87119
R89 source.n16 source.n14 0.87119
R90 source.n9 source.n7 0.802224
R91 source.n7 source.n5 0.802224
R92 source.n4 source.n2 0.802224
R93 source.n2 source.n0 0.802224
R94 source.n13 source.n11 0.802224
R95 source.n14 source.n13 0.802224
R96 source.n18 source.n16 0.802224
R97 source.n19 source.n18 0.802224
R98 source source.n20 0.188
R99 plus.n3 plus.t8 694.173
R100 plus.n13 plus.t0 694.173
R101 plus.n8 plus.t3 667.972
R102 plus.n6 plus.t5 667.972
R103 plus.n5 plus.t6 667.972
R104 plus.n4 plus.t7 667.972
R105 plus.n18 plus.t2 667.972
R106 plus.n16 plus.t1 667.972
R107 plus.n15 plus.t9 667.972
R108 plus.n14 plus.t4 667.972
R109 plus.n6 plus.n1 161.3
R110 plus.n7 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n16 plus.n11 161.3
R113 plus.n17 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n5 plus.n2 80.6037
R116 plus.n15 plus.n12 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n8 plus.n7 45.2793
R122 plus.n18 plus.n17 45.2793
R123 plus.n3 plus.n2 45.1669
R124 plus.n13 plus.n12 45.1669
R125 plus plus.n19 31.1789
R126 plus.n4 plus.n3 14.3992
R127 plus.n14 plus.n13 14.3992
R128 plus plus.n9 13.3812
R129 plus.n7 plus.n6 2.92171
R130 plus.n17 plus.n16 2.92171
R131 plus.n2 plus.n1 0.285035
R132 plus.n12 plus.n11 0.285035
R133 plus.n1 plus.n0 0.189894
R134 plus.n9 plus.n0 0.189894
R135 plus.n19 plus.n10 0.189894
R136 plus.n11 plus.n10 0.189894
R137 drain_left.n5 drain_left.t1 63.0015
R138 drain_left.n1 drain_left.t7 63.0013
R139 drain_left.n3 drain_left.n2 61.4255
R140 drain_left.n5 drain_left.n4 60.8798
R141 drain_left.n7 drain_left.n6 60.8796
R142 drain_left.n1 drain_left.n0 60.8796
R143 drain_left drain_left.n3 33.0471
R144 drain_left drain_left.n7 6.45494
R145 drain_left.n2 drain_left.t5 1.3205
R146 drain_left.n2 drain_left.t9 1.3205
R147 drain_left.n0 drain_left.t8 1.3205
R148 drain_left.n0 drain_left.t0 1.3205
R149 drain_left.n6 drain_left.t4 1.3205
R150 drain_left.n6 drain_left.t6 1.3205
R151 drain_left.n4 drain_left.t2 1.3205
R152 drain_left.n4 drain_left.t3 1.3205
R153 drain_left.n7 drain_left.n5 0.802224
R154 drain_left.n3 drain_left.n1 0.145585
C0 drain_right plus 0.335383f
C1 drain_left drain_right 0.910937f
C2 minus source 7.24892f
C3 plus minus 5.98535f
C4 plus source 7.26362f
C5 drain_left minus 0.172117f
C6 drain_right minus 7.59298f
C7 drain_left source 18.5994f
C8 drain_right source 18.589802f
C9 drain_left plus 7.76771f
C10 drain_right a_n1832_n3888# 7.72936f
C11 drain_left a_n1832_n3888# 8.01409f
C12 source a_n1832_n3888# 7.546754f
C13 minus a_n1832_n3888# 7.346212f
C14 plus a_n1832_n3888# 9.277519f
C15 drain_left.t7 a_n1832_n3888# 3.43778f
C16 drain_left.t8 a_n1832_n3888# 0.297578f
C17 drain_left.t0 a_n1832_n3888# 0.297578f
C18 drain_left.n0 a_n1832_n3888# 2.68975f
C19 drain_left.n1 a_n1832_n3888# 0.630368f
C20 drain_left.t5 a_n1832_n3888# 0.297578f
C21 drain_left.t9 a_n1832_n3888# 0.297578f
C22 drain_left.n2 a_n1832_n3888# 2.69265f
C23 drain_left.n3 a_n1832_n3888# 1.74369f
C24 drain_left.t1 a_n1832_n3888# 3.43778f
C25 drain_left.t2 a_n1832_n3888# 0.297578f
C26 drain_left.t3 a_n1832_n3888# 0.297578f
C27 drain_left.n4 a_n1832_n3888# 2.68976f
C28 drain_left.n5 a_n1832_n3888# 0.679469f
C29 drain_left.t4 a_n1832_n3888# 0.297578f
C30 drain_left.t6 a_n1832_n3888# 0.297578f
C31 drain_left.n6 a_n1832_n3888# 2.68975f
C32 drain_left.n7 a_n1832_n3888# 0.554249f
C33 plus.n0 a_n1832_n3888# 0.045695f
C34 plus.t3 a_n1832_n3888# 1.16868f
C35 plus.t5 a_n1832_n3888# 1.16868f
C36 plus.n1 a_n1832_n3888# 0.060975f
C37 plus.t6 a_n1832_n3888# 1.16868f
C38 plus.n2 a_n1832_n3888# 0.220867f
C39 plus.t7 a_n1832_n3888# 1.16868f
C40 plus.t8 a_n1832_n3888# 1.18578f
C41 plus.n3 a_n1832_n3888# 0.438214f
C42 plus.n4 a_n1832_n3888# 0.462804f
C43 plus.n5 a_n1832_n3888# 0.463571f
C44 plus.n6 a_n1832_n3888# 0.453765f
C45 plus.n7 a_n1832_n3888# 0.010369f
C46 plus.n8 a_n1832_n3888# 0.452638f
C47 plus.n9 a_n1832_n3888# 0.588281f
C48 plus.n10 a_n1832_n3888# 0.045695f
C49 plus.t2 a_n1832_n3888# 1.16868f
C50 plus.n11 a_n1832_n3888# 0.060975f
C51 plus.t1 a_n1832_n3888# 1.16868f
C52 plus.n12 a_n1832_n3888# 0.220867f
C53 plus.t9 a_n1832_n3888# 1.16868f
C54 plus.t0 a_n1832_n3888# 1.18578f
C55 plus.n13 a_n1832_n3888# 0.438214f
C56 plus.t4 a_n1832_n3888# 1.16868f
C57 plus.n14 a_n1832_n3888# 0.462804f
C58 plus.n15 a_n1832_n3888# 0.463571f
C59 plus.n16 a_n1832_n3888# 0.453765f
C60 plus.n17 a_n1832_n3888# 0.010369f
C61 plus.n18 a_n1832_n3888# 0.452638f
C62 plus.n19 a_n1832_n3888# 1.46207f
C63 source.t17 a_n1832_n3888# 3.43067f
C64 source.n0 a_n1832_n3888# 1.62371f
C65 source.t1 a_n1832_n3888# 0.306129f
C66 source.t16 a_n1832_n3888# 0.306129f
C67 source.n1 a_n1832_n3888# 2.68908f
C68 source.n2 a_n1832_n3888# 0.387825f
C69 source.t15 a_n1832_n3888# 0.306129f
C70 source.t2 a_n1832_n3888# 0.306129f
C71 source.n3 a_n1832_n3888# 2.68908f
C72 source.n4 a_n1832_n3888# 0.393564f
C73 source.t6 a_n1832_n3888# 3.43067f
C74 source.n5 a_n1832_n3888# 0.486875f
C75 source.t9 a_n1832_n3888# 0.306129f
C76 source.t7 a_n1832_n3888# 0.306129f
C77 source.n6 a_n1832_n3888# 2.68908f
C78 source.n7 a_n1832_n3888# 0.387825f
C79 source.t13 a_n1832_n3888# 0.306129f
C80 source.t10 a_n1832_n3888# 0.306129f
C81 source.n8 a_n1832_n3888# 2.68908f
C82 source.n9 a_n1832_n3888# 2.03485f
C83 source.t3 a_n1832_n3888# 0.306129f
C84 source.t0 a_n1832_n3888# 0.306129f
C85 source.n10 a_n1832_n3888# 2.68908f
C86 source.n11 a_n1832_n3888# 2.03485f
C87 source.t18 a_n1832_n3888# 0.306129f
C88 source.t4 a_n1832_n3888# 0.306129f
C89 source.n12 a_n1832_n3888# 2.68908f
C90 source.n13 a_n1832_n3888# 0.387829f
C91 source.t19 a_n1832_n3888# 3.43067f
C92 source.n14 a_n1832_n3888# 0.486879f
C93 source.t5 a_n1832_n3888# 0.306129f
C94 source.t11 a_n1832_n3888# 0.306129f
C95 source.n15 a_n1832_n3888# 2.68908f
C96 source.n16 a_n1832_n3888# 0.393568f
C97 source.t8 a_n1832_n3888# 0.306129f
C98 source.t14 a_n1832_n3888# 0.306129f
C99 source.n17 a_n1832_n3888# 2.68908f
C100 source.n18 a_n1832_n3888# 0.387829f
C101 source.t12 a_n1832_n3888# 3.43067f
C102 source.n19 a_n1832_n3888# 0.616364f
C103 source.n20 a_n1832_n3888# 1.90118f
C104 drain_right.t2 a_n1832_n3888# 3.42447f
C105 drain_right.t6 a_n1832_n3888# 0.296426f
C106 drain_right.t5 a_n1832_n3888# 0.296426f
C107 drain_right.n0 a_n1832_n3888# 2.67934f
C108 drain_right.n1 a_n1832_n3888# 0.627928f
C109 drain_right.t7 a_n1832_n3888# 0.296426f
C110 drain_right.t9 a_n1832_n3888# 0.296426f
C111 drain_right.n2 a_n1832_n3888# 2.68223f
C112 drain_right.n3 a_n1832_n3888# 1.68487f
C113 drain_right.t3 a_n1832_n3888# 0.296426f
C114 drain_right.t8 a_n1832_n3888# 0.296426f
C115 drain_right.n4 a_n1832_n3888# 2.68381f
C116 drain_right.t0 a_n1832_n3888# 0.296426f
C117 drain_right.t1 a_n1832_n3888# 0.296426f
C118 drain_right.n5 a_n1832_n3888# 2.67935f
C119 drain_right.n6 a_n1832_n3888# 0.673671f
C120 drain_right.t4 a_n1832_n3888# 3.42005f
C121 drain_right.n7 a_n1832_n3888# 0.571798f
C122 minus.n0 a_n1832_n3888# 0.044849f
C123 minus.t5 a_n1832_n3888# 1.14704f
C124 minus.n1 a_n1832_n3888# 0.454987f
C125 minus.t4 a_n1832_n3888# 1.14704f
C126 minus.t8 a_n1832_n3888# 1.16382f
C127 minus.t7 a_n1832_n3888# 1.14704f
C128 minus.n2 a_n1832_n3888# 0.454234f
C129 minus.n3 a_n1832_n3888# 0.430099f
C130 minus.n4 a_n1832_n3888# 0.216777f
C131 minus.n5 a_n1832_n3888# 0.059846f
C132 minus.n6 a_n1832_n3888# 0.445363f
C133 minus.n7 a_n1832_n3888# 0.010177f
C134 minus.t1 a_n1832_n3888# 1.14704f
C135 minus.n8 a_n1832_n3888# 0.444257f
C136 minus.n9 a_n1832_n3888# 1.74231f
C137 minus.n10 a_n1832_n3888# 0.044849f
C138 minus.t6 a_n1832_n3888# 1.14704f
C139 minus.n11 a_n1832_n3888# 0.454987f
C140 minus.t9 a_n1832_n3888# 1.16382f
C141 minus.t3 a_n1832_n3888# 1.14704f
C142 minus.n12 a_n1832_n3888# 0.454234f
C143 minus.n13 a_n1832_n3888# 0.430099f
C144 minus.n14 a_n1832_n3888# 0.216777f
C145 minus.n15 a_n1832_n3888# 0.059846f
C146 minus.t0 a_n1832_n3888# 1.14704f
C147 minus.n16 a_n1832_n3888# 0.445363f
C148 minus.n17 a_n1832_n3888# 0.010177f
C149 minus.t2 a_n1832_n3888# 1.14704f
C150 minus.n18 a_n1832_n3888# 0.444257f
C151 minus.n19 a_n1832_n3888# 0.303822f
C152 minus.n20 a_n1832_n3888# 2.09929f
.ends

