* NGSPICE file created from diffpair691.ext - technology: sky130A

.subckt diffpair691 minus drain_right drain_left source plus
X0 a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.6
X1 a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X2 drain_right minus source a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X3 a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X4 source plus drain_left a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X5 source minus drain_right a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X6 drain_right minus source a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X7 drain_left plus source a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X8 source plus drain_left a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X9 source minus drain_right a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X10 a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X11 drain_left plus source a_n1274_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
.ends

