* NGSPICE file created from diffpair501.ext - technology: sky130A

.subckt diffpair501 minus drain_right drain_left source plus
X0 drain_right minus source a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X1 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X2 source plus drain_left a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X3 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X4 drain_left plus source a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X5 drain_left plus source a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X6 source minus drain_right a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X7 source minus drain_right a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X9 source plus drain_left a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X10 drain_right minus source a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X11 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
.ends

