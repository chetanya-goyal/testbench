* NGSPICE file created from diffpair103.ext - technology: sky130A

.subckt diffpair103 minus drain_right drain_left source plus
X0 a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X1 drain_left.t7 plus.t0 source.t7 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X2 drain_left.t6 plus.t1 source.t12 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 drain_left.t5 plus.t2 source.t10 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 source.t14 minus.t0 drain_right.t7 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X5 source.t3 minus.t1 drain_right.t6 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 source.t11 plus.t3 drain_left.t4 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X7 source.t8 plus.t4 drain_left.t3 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X8 drain_right.t5 minus.t2 source.t0 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X9 a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X10 drain_right.t4 minus.t3 source.t15 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X11 a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X12 source.t1 minus.t4 drain_right.t3 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X13 source.t6 plus.t5 drain_left.t2 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X14 source.t2 minus.t5 drain_right.t2 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X15 drain_right.t1 minus.t6 source.t5 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X16 drain_right.t0 minus.t7 source.t4 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X17 source.t9 plus.t6 drain_left.t1 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X18 drain_left.t0 plus.t7 source.t13 a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X19 a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# a_n1296_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
R0 plus.n1 plus.t4 372.163
R1 plus.n5 plus.t0 372.163
R2 plus.n8 plus.t7 372.163
R3 plus.n12 plus.t3 372.163
R4 plus.n2 plus.t1 318.12
R5 plus.n4 plus.t5 318.12
R6 plus.n9 plus.t6 318.12
R7 plus.n11 plus.t2 318.12
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 24.124
R23 plus plus.n6 8.35656
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n66 source.n64 289.615
R27 source.n56 source.n54 289.615
R28 source.n48 source.n46 289.615
R29 source.n38 source.n36 289.615
R30 source.n2 source.n0 289.615
R31 source.n12 source.n10 289.615
R32 source.n20 source.n18 289.615
R33 source.n30 source.n28 289.615
R34 source.n67 source.n66 185
R35 source.n57 source.n56 185
R36 source.n49 source.n48 185
R37 source.n39 source.n38 185
R38 source.n3 source.n2 185
R39 source.n13 source.n12 185
R40 source.n21 source.n20 185
R41 source.n31 source.n30 185
R42 source.t15 source.n65 167.117
R43 source.t2 source.n55 167.117
R44 source.t13 source.n47 167.117
R45 source.t11 source.n37 167.117
R46 source.t7 source.n1 167.117
R47 source.t8 source.n11 167.117
R48 source.t4 source.n19 167.117
R49 source.t14 source.n29 167.117
R50 source.n9 source.n8 84.1169
R51 source.n27 source.n26 84.1169
R52 source.n63 source.n62 84.1168
R53 source.n45 source.n44 84.1168
R54 source.n66 source.t15 52.3082
R55 source.n56 source.t2 52.3082
R56 source.n48 source.t13 52.3082
R57 source.n38 source.t11 52.3082
R58 source.n2 source.t7 52.3082
R59 source.n12 source.t8 52.3082
R60 source.n20 source.t4 52.3082
R61 source.n30 source.t14 52.3082
R62 source.n71 source.n70 31.4096
R63 source.n61 source.n60 31.4096
R64 source.n53 source.n52 31.4096
R65 source.n43 source.n42 31.4096
R66 source.n7 source.n6 31.4096
R67 source.n17 source.n16 31.4096
R68 source.n25 source.n24 31.4096
R69 source.n35 source.n34 31.4096
R70 source.n43 source.n35 14.212
R71 source.n62 source.t0 9.9005
R72 source.n62 source.t1 9.9005
R73 source.n44 source.t10 9.9005
R74 source.n44 source.t9 9.9005
R75 source.n8 source.t12 9.9005
R76 source.n8 source.t6 9.9005
R77 source.n26 source.t5 9.9005
R78 source.n26 source.t3 9.9005
R79 source.n67 source.n65 9.71174
R80 source.n57 source.n55 9.71174
R81 source.n49 source.n47 9.71174
R82 source.n39 source.n37 9.71174
R83 source.n3 source.n1 9.71174
R84 source.n13 source.n11 9.71174
R85 source.n21 source.n19 9.71174
R86 source.n31 source.n29 9.71174
R87 source.n70 source.n69 9.45567
R88 source.n60 source.n59 9.45567
R89 source.n52 source.n51 9.45567
R90 source.n42 source.n41 9.45567
R91 source.n6 source.n5 9.45567
R92 source.n16 source.n15 9.45567
R93 source.n24 source.n23 9.45567
R94 source.n34 source.n33 9.45567
R95 source.n69 source.n68 9.3005
R96 source.n59 source.n58 9.3005
R97 source.n51 source.n50 9.3005
R98 source.n41 source.n40 9.3005
R99 source.n5 source.n4 9.3005
R100 source.n15 source.n14 9.3005
R101 source.n23 source.n22 9.3005
R102 source.n33 source.n32 9.3005
R103 source.n72 source.n7 8.69904
R104 source.n70 source.n64 8.14595
R105 source.n60 source.n54 8.14595
R106 source.n52 source.n46 8.14595
R107 source.n42 source.n36 8.14595
R108 source.n6 source.n0 8.14595
R109 source.n16 source.n10 8.14595
R110 source.n24 source.n18 8.14595
R111 source.n34 source.n28 8.14595
R112 source.n68 source.n67 7.3702
R113 source.n58 source.n57 7.3702
R114 source.n50 source.n49 7.3702
R115 source.n40 source.n39 7.3702
R116 source.n4 source.n3 7.3702
R117 source.n14 source.n13 7.3702
R118 source.n22 source.n21 7.3702
R119 source.n32 source.n31 7.3702
R120 source.n68 source.n64 5.81868
R121 source.n58 source.n54 5.81868
R122 source.n50 source.n46 5.81868
R123 source.n40 source.n36 5.81868
R124 source.n4 source.n0 5.81868
R125 source.n14 source.n10 5.81868
R126 source.n22 source.n18 5.81868
R127 source.n32 source.n28 5.81868
R128 source.n72 source.n71 5.51343
R129 source.n69 source.n65 3.44771
R130 source.n59 source.n55 3.44771
R131 source.n51 source.n47 3.44771
R132 source.n41 source.n37 3.44771
R133 source.n5 source.n1 3.44771
R134 source.n15 source.n11 3.44771
R135 source.n23 source.n19 3.44771
R136 source.n33 source.n29 3.44771
R137 source.n35 source.n27 0.5005
R138 source.n27 source.n25 0.5005
R139 source.n17 source.n9 0.5005
R140 source.n9 source.n7 0.5005
R141 source.n45 source.n43 0.5005
R142 source.n53 source.n45 0.5005
R143 source.n63 source.n61 0.5005
R144 source.n71 source.n63 0.5005
R145 source.n25 source.n17 0.470328
R146 source.n61 source.n53 0.470328
R147 source source.n72 0.188
R148 drain_left.n5 drain_left.n3 101.296
R149 drain_left.n2 drain_left.n1 100.99
R150 drain_left.n2 drain_left.n0 100.99
R151 drain_left.n5 drain_left.n4 100.796
R152 drain_left drain_left.n2 21.5413
R153 drain_left.n1 drain_left.t1 9.9005
R154 drain_left.n1 drain_left.t0 9.9005
R155 drain_left.n0 drain_left.t4 9.9005
R156 drain_left.n0 drain_left.t5 9.9005
R157 drain_left.n4 drain_left.t2 9.9005
R158 drain_left.n4 drain_left.t7 9.9005
R159 drain_left.n3 drain_left.t3 9.9005
R160 drain_left.n3 drain_left.t6 9.9005
R161 drain_left drain_left.n5 6.15322
R162 minus.n5 minus.t0 372.163
R163 minus.n1 minus.t7 372.163
R164 minus.n12 minus.t3 372.163
R165 minus.n8 minus.t5 372.163
R166 minus.n4 minus.t6 318.12
R167 minus.n2 minus.t1 318.12
R168 minus.n11 minus.t4 318.12
R169 minus.n9 minus.t2 318.12
R170 minus.n1 minus.n0 161.489
R171 minus.n8 minus.n7 161.489
R172 minus.n6 minus.n5 161.3
R173 minus.n3 minus.n0 161.3
R174 minus.n13 minus.n12 161.3
R175 minus.n10 minus.n7 161.3
R176 minus.n4 minus.n3 42.3581
R177 minus.n3 minus.n2 42.3581
R178 minus.n10 minus.n9 42.3581
R179 minus.n11 minus.n10 42.3581
R180 minus.n5 minus.n4 30.6732
R181 minus.n2 minus.n1 30.6732
R182 minus.n9 minus.n8 30.6732
R183 minus.n12 minus.n11 30.6732
R184 minus.n14 minus.n6 26.455
R185 minus.n14 minus.n13 6.5005
R186 minus.n6 minus.n0 0.189894
R187 minus.n13 minus.n7 0.189894
R188 minus minus.n14 0.188
R189 drain_right.n5 drain_right.n3 101.296
R190 drain_right.n2 drain_right.n1 100.99
R191 drain_right.n2 drain_right.n0 100.99
R192 drain_right.n5 drain_right.n4 100.796
R193 drain_right drain_right.n2 20.9881
R194 drain_right.n1 drain_right.t3 9.9005
R195 drain_right.n1 drain_right.t4 9.9005
R196 drain_right.n0 drain_right.t2 9.9005
R197 drain_right.n0 drain_right.t5 9.9005
R198 drain_right.n3 drain_right.t6 9.9005
R199 drain_right.n3 drain_right.t0 9.9005
R200 drain_right.n4 drain_right.t7 9.9005
R201 drain_right.n4 drain_right.t1 9.9005
R202 drain_right drain_right.n5 6.15322
C0 minus source 0.847864f
C1 minus drain_left 0.176215f
C2 plus minus 2.92188f
C3 source drain_left 4.48059f
C4 minus drain_right 0.793141f
C5 plus source 0.861827f
C6 plus drain_left 0.91516f
C7 drain_right source 4.47947f
C8 drain_right drain_left 0.605638f
C9 plus drain_right 0.281667f
C10 drain_right a_n1296_n1288# 3.12749f
C11 drain_left a_n1296_n1288# 3.28618f
C12 source a_n1296_n1288# 2.85049f
C13 minus a_n1296_n1288# 4.18613f
C14 plus a_n1296_n1288# 4.903523f
C15 drain_right.t2 a_n1296_n1288# 0.041253f
C16 drain_right.t5 a_n1296_n1288# 0.041253f
C17 drain_right.n0 a_n1296_n1288# 0.259687f
C18 drain_right.t3 a_n1296_n1288# 0.041253f
C19 drain_right.t4 a_n1296_n1288# 0.041253f
C20 drain_right.n1 a_n1296_n1288# 0.259687f
C21 drain_right.n2 a_n1296_n1288# 1.09209f
C22 drain_right.t6 a_n1296_n1288# 0.041253f
C23 drain_right.t0 a_n1296_n1288# 0.041253f
C24 drain_right.n3 a_n1296_n1288# 0.260617f
C25 drain_right.t7 a_n1296_n1288# 0.041253f
C26 drain_right.t1 a_n1296_n1288# 0.041253f
C27 drain_right.n4 a_n1296_n1288# 0.259164f
C28 drain_right.n5 a_n1296_n1288# 0.792282f
C29 minus.n0 a_n1296_n1288# 0.08201f
C30 minus.t0 a_n1296_n1288# 0.058416f
C31 minus.t6 a_n1296_n1288# 0.052448f
C32 minus.t1 a_n1296_n1288# 0.052448f
C33 minus.t7 a_n1296_n1288# 0.058416f
C34 minus.n1 a_n1296_n1288# 0.048769f
C35 minus.n2 a_n1296_n1288# 0.038462f
C36 minus.n3 a_n1296_n1288# 0.013584f
C37 minus.n4 a_n1296_n1288# 0.038462f
C38 minus.n5 a_n1296_n1288# 0.048715f
C39 minus.n6 a_n1296_n1288# 0.742738f
C40 minus.n7 a_n1296_n1288# 0.08201f
C41 minus.t4 a_n1296_n1288# 0.052448f
C42 minus.t2 a_n1296_n1288# 0.052448f
C43 minus.t5 a_n1296_n1288# 0.058416f
C44 minus.n8 a_n1296_n1288# 0.048769f
C45 minus.n9 a_n1296_n1288# 0.038462f
C46 minus.n10 a_n1296_n1288# 0.013584f
C47 minus.n11 a_n1296_n1288# 0.038462f
C48 minus.t3 a_n1296_n1288# 0.058416f
C49 minus.n12 a_n1296_n1288# 0.048715f
C50 minus.n13 a_n1296_n1288# 0.233097f
C51 minus.n14 a_n1296_n1288# 0.917293f
C52 drain_left.t4 a_n1296_n1288# 0.040338f
C53 drain_left.t5 a_n1296_n1288# 0.040338f
C54 drain_left.n0 a_n1296_n1288# 0.253925f
C55 drain_left.t1 a_n1296_n1288# 0.040338f
C56 drain_left.t0 a_n1296_n1288# 0.040338f
C57 drain_left.n1 a_n1296_n1288# 0.253925f
C58 drain_left.n2 a_n1296_n1288# 1.11814f
C59 drain_left.t3 a_n1296_n1288# 0.040338f
C60 drain_left.t6 a_n1296_n1288# 0.040338f
C61 drain_left.n3 a_n1296_n1288# 0.254835f
C62 drain_left.t2 a_n1296_n1288# 0.040338f
C63 drain_left.t7 a_n1296_n1288# 0.040338f
C64 drain_left.n4 a_n1296_n1288# 0.253414f
C65 drain_left.n5 a_n1296_n1288# 0.774704f
C66 source.n0 a_n1296_n1288# 0.0362f
C67 source.n1 a_n1296_n1288# 0.080097f
C68 source.t7 a_n1296_n1288# 0.060109f
C69 source.n2 a_n1296_n1288# 0.062687f
C70 source.n3 a_n1296_n1288# 0.020208f
C71 source.n4 a_n1296_n1288# 0.013327f
C72 source.n5 a_n1296_n1288# 0.176553f
C73 source.n6 a_n1296_n1288# 0.039683f
C74 source.n7 a_n1296_n1288# 0.368345f
C75 source.t12 a_n1296_n1288# 0.039198f
C76 source.t6 a_n1296_n1288# 0.039198f
C77 source.n8 a_n1296_n1288# 0.209554f
C78 source.n9 a_n1296_n1288# 0.272741f
C79 source.n10 a_n1296_n1288# 0.0362f
C80 source.n11 a_n1296_n1288# 0.080097f
C81 source.t8 a_n1296_n1288# 0.060109f
C82 source.n12 a_n1296_n1288# 0.062687f
C83 source.n13 a_n1296_n1288# 0.020208f
C84 source.n14 a_n1296_n1288# 0.013327f
C85 source.n15 a_n1296_n1288# 0.176553f
C86 source.n16 a_n1296_n1288# 0.039683f
C87 source.n17 a_n1296_n1288# 0.097924f
C88 source.n18 a_n1296_n1288# 0.0362f
C89 source.n19 a_n1296_n1288# 0.080097f
C90 source.t4 a_n1296_n1288# 0.060109f
C91 source.n20 a_n1296_n1288# 0.062687f
C92 source.n21 a_n1296_n1288# 0.020208f
C93 source.n22 a_n1296_n1288# 0.013327f
C94 source.n23 a_n1296_n1288# 0.176553f
C95 source.n24 a_n1296_n1288# 0.039683f
C96 source.n25 a_n1296_n1288# 0.097924f
C97 source.t5 a_n1296_n1288# 0.039198f
C98 source.t3 a_n1296_n1288# 0.039198f
C99 source.n26 a_n1296_n1288# 0.209554f
C100 source.n27 a_n1296_n1288# 0.272741f
C101 source.n28 a_n1296_n1288# 0.0362f
C102 source.n29 a_n1296_n1288# 0.080097f
C103 source.t14 a_n1296_n1288# 0.060109f
C104 source.n30 a_n1296_n1288# 0.062687f
C105 source.n31 a_n1296_n1288# 0.020208f
C106 source.n32 a_n1296_n1288# 0.013327f
C107 source.n33 a_n1296_n1288# 0.176553f
C108 source.n34 a_n1296_n1288# 0.039683f
C109 source.n35 a_n1296_n1288# 0.598808f
C110 source.n36 a_n1296_n1288# 0.0362f
C111 source.n37 a_n1296_n1288# 0.080097f
C112 source.t11 a_n1296_n1288# 0.060109f
C113 source.n38 a_n1296_n1288# 0.062687f
C114 source.n39 a_n1296_n1288# 0.020208f
C115 source.n40 a_n1296_n1288# 0.013327f
C116 source.n41 a_n1296_n1288# 0.176553f
C117 source.n42 a_n1296_n1288# 0.039683f
C118 source.n43 a_n1296_n1288# 0.598808f
C119 source.t10 a_n1296_n1288# 0.039198f
C120 source.t9 a_n1296_n1288# 0.039198f
C121 source.n44 a_n1296_n1288# 0.209553f
C122 source.n45 a_n1296_n1288# 0.272742f
C123 source.n46 a_n1296_n1288# 0.0362f
C124 source.n47 a_n1296_n1288# 0.080097f
C125 source.t13 a_n1296_n1288# 0.060109f
C126 source.n48 a_n1296_n1288# 0.062687f
C127 source.n49 a_n1296_n1288# 0.020208f
C128 source.n50 a_n1296_n1288# 0.013327f
C129 source.n51 a_n1296_n1288# 0.176553f
C130 source.n52 a_n1296_n1288# 0.039683f
C131 source.n53 a_n1296_n1288# 0.097924f
C132 source.n54 a_n1296_n1288# 0.0362f
C133 source.n55 a_n1296_n1288# 0.080097f
C134 source.t2 a_n1296_n1288# 0.060109f
C135 source.n56 a_n1296_n1288# 0.062687f
C136 source.n57 a_n1296_n1288# 0.020208f
C137 source.n58 a_n1296_n1288# 0.013327f
C138 source.n59 a_n1296_n1288# 0.176553f
C139 source.n60 a_n1296_n1288# 0.039683f
C140 source.n61 a_n1296_n1288# 0.097924f
C141 source.t0 a_n1296_n1288# 0.039198f
C142 source.t1 a_n1296_n1288# 0.039198f
C143 source.n62 a_n1296_n1288# 0.209553f
C144 source.n63 a_n1296_n1288# 0.272742f
C145 source.n64 a_n1296_n1288# 0.0362f
C146 source.n65 a_n1296_n1288# 0.080097f
C147 source.t15 a_n1296_n1288# 0.060109f
C148 source.n66 a_n1296_n1288# 0.062687f
C149 source.n67 a_n1296_n1288# 0.020208f
C150 source.n68 a_n1296_n1288# 0.013327f
C151 source.n69 a_n1296_n1288# 0.176553f
C152 source.n70 a_n1296_n1288# 0.039683f
C153 source.n71 a_n1296_n1288# 0.235173f
C154 source.n72 a_n1296_n1288# 0.61174f
C155 plus.n0 a_n1296_n1288# 0.084101f
C156 plus.t5 a_n1296_n1288# 0.053785f
C157 plus.t1 a_n1296_n1288# 0.053785f
C158 plus.t4 a_n1296_n1288# 0.059905f
C159 plus.n1 a_n1296_n1288# 0.050013f
C160 plus.n2 a_n1296_n1288# 0.039442f
C161 plus.n3 a_n1296_n1288# 0.01393f
C162 plus.n4 a_n1296_n1288# 0.039442f
C163 plus.t0 a_n1296_n1288# 0.059905f
C164 plus.n5 a_n1296_n1288# 0.049957f
C165 plus.n6 a_n1296_n1288# 0.261383f
C166 plus.n7 a_n1296_n1288# 0.084101f
C167 plus.t3 a_n1296_n1288# 0.059905f
C168 plus.t2 a_n1296_n1288# 0.053785f
C169 plus.t6 a_n1296_n1288# 0.053785f
C170 plus.t7 a_n1296_n1288# 0.059905f
C171 plus.n8 a_n1296_n1288# 0.050013f
C172 plus.n9 a_n1296_n1288# 0.039442f
C173 plus.n10 a_n1296_n1288# 0.01393f
C174 plus.n11 a_n1296_n1288# 0.039442f
C175 plus.n12 a_n1296_n1288# 0.049957f
C176 plus.n13 a_n1296_n1288# 0.732042f
.ends

