* NGSPICE file created from diffpair304.ext - technology: sky130A

.subckt diffpair304 minus drain_right drain_left source plus
X0 source.t17 plus.t0 drain_left.t6 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X1 drain_left.t8 plus.t1 source.t16 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X2 source.t18 minus.t0 drain_right.t9 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 drain_left.t1 plus.t2 source.t15 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X4 a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X5 drain_left.t9 plus.t3 source.t14 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X6 drain_left.t5 plus.t4 source.t13 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X7 drain_left.t2 plus.t5 source.t12 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X8 drain_right.t8 minus.t1 source.t5 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X9 a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X10 drain_left.t0 plus.t6 source.t11 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X11 drain_right.t7 minus.t2 source.t0 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 drain_right.t6 minus.t3 source.t19 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 source.t10 plus.t7 drain_left.t7 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X14 source.t9 plus.t8 drain_left.t3 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 source.t1 minus.t4 drain_right.t5 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X16 a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X17 a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X18 drain_right.t4 minus.t5 source.t2 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X19 drain_right.t3 minus.t6 source.t7 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X20 source.t8 plus.t9 drain_left.t4 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X21 drain_right.t2 minus.t7 source.t3 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X22 source.t6 minus.t8 drain_right.t1 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X23 source.t4 minus.t9 drain_right.t0 a_n1952_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n3 plus.t4 285.438
R1 plus.n17 plus.t6 285.438
R2 plus.n12 plus.t3 262.69
R3 plus.n10 plus.t8 262.69
R4 plus.n2 plus.t1 262.69
R5 plus.n4 plus.t9 262.69
R6 plus.n26 plus.t2 262.69
R7 plus.n24 plus.t0 262.69
R8 plus.n16 plus.t5 262.69
R9 plus.n18 plus.t7 262.69
R10 plus.n6 plus.n5 161.3
R11 plus.n7 plus.n2 161.3
R12 plus.n9 plus.n8 161.3
R13 plus.n10 plus.n1 161.3
R14 plus.n11 plus.n0 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n20 plus.n19 161.3
R17 plus.n21 plus.n16 161.3
R18 plus.n23 plus.n22 161.3
R19 plus.n24 plus.n15 161.3
R20 plus.n25 plus.n14 161.3
R21 plus.n27 plus.n26 161.3
R22 plus.n6 plus.n3 44.8741
R23 plus.n20 plus.n17 44.8741
R24 plus.n12 plus.n11 30.6732
R25 plus.n26 plus.n25 30.6732
R26 plus plus.n27 28.2623
R27 plus.n10 plus.n9 26.2914
R28 plus.n5 plus.n4 26.2914
R29 plus.n24 plus.n23 26.2914
R30 plus.n19 plus.n18 26.2914
R31 plus.n9 plus.n2 21.9096
R32 plus.n5 plus.n2 21.9096
R33 plus.n23 plus.n16 21.9096
R34 plus.n19 plus.n16 21.9096
R35 plus.n4 plus.n3 19.0667
R36 plus.n18 plus.n17 19.0667
R37 plus.n11 plus.n10 17.5278
R38 plus.n25 plus.n24 17.5278
R39 plus plus.n13 10.01
R40 plus.n7 plus.n6 0.189894
R41 plus.n8 plus.n7 0.189894
R42 plus.n8 plus.n1 0.189894
R43 plus.n1 plus.n0 0.189894
R44 plus.n13 plus.n0 0.189894
R45 plus.n27 plus.n14 0.189894
R46 plus.n15 plus.n14 0.189894
R47 plus.n22 plus.n15 0.189894
R48 plus.n22 plus.n21 0.189894
R49 plus.n21 plus.n20 0.189894
R50 drain_left.n26 drain_left.n0 289.615
R51 drain_left.n61 drain_left.n35 289.615
R52 drain_left.n11 drain_left.n10 185
R53 drain_left.n8 drain_left.n7 185
R54 drain_left.n17 drain_left.n16 185
R55 drain_left.n19 drain_left.n18 185
R56 drain_left.n4 drain_left.n3 185
R57 drain_left.n25 drain_left.n24 185
R58 drain_left.n27 drain_left.n26 185
R59 drain_left.n62 drain_left.n61 185
R60 drain_left.n60 drain_left.n59 185
R61 drain_left.n39 drain_left.n38 185
R62 drain_left.n54 drain_left.n53 185
R63 drain_left.n52 drain_left.n51 185
R64 drain_left.n43 drain_left.n42 185
R65 drain_left.n46 drain_left.n45 185
R66 drain_left.t1 drain_left.n9 147.661
R67 drain_left.t5 drain_left.n44 147.661
R68 drain_left.n10 drain_left.n7 104.615
R69 drain_left.n17 drain_left.n7 104.615
R70 drain_left.n18 drain_left.n17 104.615
R71 drain_left.n18 drain_left.n3 104.615
R72 drain_left.n25 drain_left.n3 104.615
R73 drain_left.n26 drain_left.n25 104.615
R74 drain_left.n61 drain_left.n60 104.615
R75 drain_left.n60 drain_left.n38 104.615
R76 drain_left.n53 drain_left.n38 104.615
R77 drain_left.n53 drain_left.n52 104.615
R78 drain_left.n52 drain_left.n42 104.615
R79 drain_left.n45 drain_left.n42 104.615
R80 drain_left.n34 drain_left.n33 67.8013
R81 drain_left.n67 drain_left.n66 67.1908
R82 drain_left.n69 drain_left.n68 67.1907
R83 drain_left.n32 drain_left.n31 67.1907
R84 drain_left.n10 drain_left.t1 52.3082
R85 drain_left.n45 drain_left.t5 52.3082
R86 drain_left.n32 drain_left.n30 49.7521
R87 drain_left.n67 drain_left.n65 49.7521
R88 drain_left drain_left.n34 26.5953
R89 drain_left.n11 drain_left.n9 15.6674
R90 drain_left.n46 drain_left.n44 15.6674
R91 drain_left.n12 drain_left.n8 12.8005
R92 drain_left.n47 drain_left.n43 12.8005
R93 drain_left.n16 drain_left.n15 12.0247
R94 drain_left.n51 drain_left.n50 12.0247
R95 drain_left.n19 drain_left.n6 11.249
R96 drain_left.n54 drain_left.n41 11.249
R97 drain_left.n20 drain_left.n4 10.4732
R98 drain_left.n55 drain_left.n39 10.4732
R99 drain_left.n24 drain_left.n23 9.69747
R100 drain_left.n59 drain_left.n58 9.69747
R101 drain_left.n30 drain_left.n29 9.45567
R102 drain_left.n65 drain_left.n64 9.45567
R103 drain_left.n29 drain_left.n28 9.3005
R104 drain_left.n2 drain_left.n1 9.3005
R105 drain_left.n23 drain_left.n22 9.3005
R106 drain_left.n21 drain_left.n20 9.3005
R107 drain_left.n6 drain_left.n5 9.3005
R108 drain_left.n15 drain_left.n14 9.3005
R109 drain_left.n13 drain_left.n12 9.3005
R110 drain_left.n64 drain_left.n63 9.3005
R111 drain_left.n37 drain_left.n36 9.3005
R112 drain_left.n58 drain_left.n57 9.3005
R113 drain_left.n56 drain_left.n55 9.3005
R114 drain_left.n41 drain_left.n40 9.3005
R115 drain_left.n50 drain_left.n49 9.3005
R116 drain_left.n48 drain_left.n47 9.3005
R117 drain_left.n27 drain_left.n2 8.92171
R118 drain_left.n62 drain_left.n37 8.92171
R119 drain_left.n28 drain_left.n0 8.14595
R120 drain_left.n63 drain_left.n35 8.14595
R121 drain_left drain_left.n69 6.54115
R122 drain_left.n30 drain_left.n0 5.81868
R123 drain_left.n65 drain_left.n35 5.81868
R124 drain_left.n28 drain_left.n27 5.04292
R125 drain_left.n63 drain_left.n62 5.04292
R126 drain_left.n13 drain_left.n9 4.38594
R127 drain_left.n48 drain_left.n44 4.38594
R128 drain_left.n24 drain_left.n2 4.26717
R129 drain_left.n59 drain_left.n37 4.26717
R130 drain_left.n23 drain_left.n4 3.49141
R131 drain_left.n58 drain_left.n39 3.49141
R132 drain_left.n33 drain_left.t7 3.3005
R133 drain_left.n33 drain_left.t0 3.3005
R134 drain_left.n31 drain_left.t6 3.3005
R135 drain_left.n31 drain_left.t2 3.3005
R136 drain_left.n68 drain_left.t3 3.3005
R137 drain_left.n68 drain_left.t9 3.3005
R138 drain_left.n66 drain_left.t4 3.3005
R139 drain_left.n66 drain_left.t8 3.3005
R140 drain_left.n20 drain_left.n19 2.71565
R141 drain_left.n55 drain_left.n54 2.71565
R142 drain_left.n16 drain_left.n6 1.93989
R143 drain_left.n51 drain_left.n41 1.93989
R144 drain_left.n15 drain_left.n8 1.16414
R145 drain_left.n50 drain_left.n43 1.16414
R146 drain_left.n69 drain_left.n67 0.888431
R147 drain_left.n12 drain_left.n11 0.388379
R148 drain_left.n47 drain_left.n46 0.388379
R149 drain_left.n34 drain_left.n32 0.167137
R150 drain_left.n14 drain_left.n13 0.155672
R151 drain_left.n14 drain_left.n5 0.155672
R152 drain_left.n21 drain_left.n5 0.155672
R153 drain_left.n22 drain_left.n21 0.155672
R154 drain_left.n22 drain_left.n1 0.155672
R155 drain_left.n29 drain_left.n1 0.155672
R156 drain_left.n64 drain_left.n36 0.155672
R157 drain_left.n57 drain_left.n36 0.155672
R158 drain_left.n57 drain_left.n56 0.155672
R159 drain_left.n56 drain_left.n40 0.155672
R160 drain_left.n49 drain_left.n40 0.155672
R161 drain_left.n49 drain_left.n48 0.155672
R162 source.n138 source.n112 289.615
R163 source.n102 source.n76 289.615
R164 source.n26 source.n0 289.615
R165 source.n62 source.n36 289.615
R166 source.n123 source.n122 185
R167 source.n120 source.n119 185
R168 source.n129 source.n128 185
R169 source.n131 source.n130 185
R170 source.n116 source.n115 185
R171 source.n137 source.n136 185
R172 source.n139 source.n138 185
R173 source.n87 source.n86 185
R174 source.n84 source.n83 185
R175 source.n93 source.n92 185
R176 source.n95 source.n94 185
R177 source.n80 source.n79 185
R178 source.n101 source.n100 185
R179 source.n103 source.n102 185
R180 source.n27 source.n26 185
R181 source.n25 source.n24 185
R182 source.n4 source.n3 185
R183 source.n19 source.n18 185
R184 source.n17 source.n16 185
R185 source.n8 source.n7 185
R186 source.n11 source.n10 185
R187 source.n63 source.n62 185
R188 source.n61 source.n60 185
R189 source.n40 source.n39 185
R190 source.n55 source.n54 185
R191 source.n53 source.n52 185
R192 source.n44 source.n43 185
R193 source.n47 source.n46 185
R194 source.t7 source.n121 147.661
R195 source.t11 source.n85 147.661
R196 source.t14 source.n9 147.661
R197 source.t2 source.n45 147.661
R198 source.n122 source.n119 104.615
R199 source.n129 source.n119 104.615
R200 source.n130 source.n129 104.615
R201 source.n130 source.n115 104.615
R202 source.n137 source.n115 104.615
R203 source.n138 source.n137 104.615
R204 source.n86 source.n83 104.615
R205 source.n93 source.n83 104.615
R206 source.n94 source.n93 104.615
R207 source.n94 source.n79 104.615
R208 source.n101 source.n79 104.615
R209 source.n102 source.n101 104.615
R210 source.n26 source.n25 104.615
R211 source.n25 source.n3 104.615
R212 source.n18 source.n3 104.615
R213 source.n18 source.n17 104.615
R214 source.n17 source.n7 104.615
R215 source.n10 source.n7 104.615
R216 source.n62 source.n61 104.615
R217 source.n61 source.n39 104.615
R218 source.n54 source.n39 104.615
R219 source.n54 source.n53 104.615
R220 source.n53 source.n43 104.615
R221 source.n46 source.n43 104.615
R222 source.n122 source.t7 52.3082
R223 source.n86 source.t11 52.3082
R224 source.n10 source.t14 52.3082
R225 source.n46 source.t2 52.3082
R226 source.n33 source.n32 50.512
R227 source.n35 source.n34 50.512
R228 source.n69 source.n68 50.512
R229 source.n71 source.n70 50.512
R230 source.n111 source.n110 50.5119
R231 source.n109 source.n108 50.5119
R232 source.n75 source.n74 50.5119
R233 source.n73 source.n72 50.5119
R234 source.n143 source.n142 32.1853
R235 source.n107 source.n106 32.1853
R236 source.n31 source.n30 32.1853
R237 source.n67 source.n66 32.1853
R238 source.n73 source.n71 18.5181
R239 source.n123 source.n121 15.6674
R240 source.n87 source.n85 15.6674
R241 source.n11 source.n9 15.6674
R242 source.n47 source.n45 15.6674
R243 source.n124 source.n120 12.8005
R244 source.n88 source.n84 12.8005
R245 source.n12 source.n8 12.8005
R246 source.n48 source.n44 12.8005
R247 source.n128 source.n127 12.0247
R248 source.n92 source.n91 12.0247
R249 source.n16 source.n15 12.0247
R250 source.n52 source.n51 12.0247
R251 source.n144 source.n31 11.9233
R252 source.n131 source.n118 11.249
R253 source.n95 source.n82 11.249
R254 source.n19 source.n6 11.249
R255 source.n55 source.n42 11.249
R256 source.n132 source.n116 10.4732
R257 source.n96 source.n80 10.4732
R258 source.n20 source.n4 10.4732
R259 source.n56 source.n40 10.4732
R260 source.n136 source.n135 9.69747
R261 source.n100 source.n99 9.69747
R262 source.n24 source.n23 9.69747
R263 source.n60 source.n59 9.69747
R264 source.n142 source.n141 9.45567
R265 source.n106 source.n105 9.45567
R266 source.n30 source.n29 9.45567
R267 source.n66 source.n65 9.45567
R268 source.n141 source.n140 9.3005
R269 source.n114 source.n113 9.3005
R270 source.n135 source.n134 9.3005
R271 source.n133 source.n132 9.3005
R272 source.n118 source.n117 9.3005
R273 source.n127 source.n126 9.3005
R274 source.n125 source.n124 9.3005
R275 source.n105 source.n104 9.3005
R276 source.n78 source.n77 9.3005
R277 source.n99 source.n98 9.3005
R278 source.n97 source.n96 9.3005
R279 source.n82 source.n81 9.3005
R280 source.n91 source.n90 9.3005
R281 source.n89 source.n88 9.3005
R282 source.n29 source.n28 9.3005
R283 source.n2 source.n1 9.3005
R284 source.n23 source.n22 9.3005
R285 source.n21 source.n20 9.3005
R286 source.n6 source.n5 9.3005
R287 source.n15 source.n14 9.3005
R288 source.n13 source.n12 9.3005
R289 source.n65 source.n64 9.3005
R290 source.n38 source.n37 9.3005
R291 source.n59 source.n58 9.3005
R292 source.n57 source.n56 9.3005
R293 source.n42 source.n41 9.3005
R294 source.n51 source.n50 9.3005
R295 source.n49 source.n48 9.3005
R296 source.n139 source.n114 8.92171
R297 source.n103 source.n78 8.92171
R298 source.n27 source.n2 8.92171
R299 source.n63 source.n38 8.92171
R300 source.n140 source.n112 8.14595
R301 source.n104 source.n76 8.14595
R302 source.n28 source.n0 8.14595
R303 source.n64 source.n36 8.14595
R304 source.n142 source.n112 5.81868
R305 source.n106 source.n76 5.81868
R306 source.n30 source.n0 5.81868
R307 source.n66 source.n36 5.81868
R308 source.n144 source.n143 5.7074
R309 source.n140 source.n139 5.04292
R310 source.n104 source.n103 5.04292
R311 source.n28 source.n27 5.04292
R312 source.n64 source.n63 5.04292
R313 source.n125 source.n121 4.38594
R314 source.n89 source.n85 4.38594
R315 source.n13 source.n9 4.38594
R316 source.n49 source.n45 4.38594
R317 source.n136 source.n114 4.26717
R318 source.n100 source.n78 4.26717
R319 source.n24 source.n2 4.26717
R320 source.n60 source.n38 4.26717
R321 source.n135 source.n116 3.49141
R322 source.n99 source.n80 3.49141
R323 source.n23 source.n4 3.49141
R324 source.n59 source.n40 3.49141
R325 source.n110 source.t19 3.3005
R326 source.n110 source.t1 3.3005
R327 source.n108 source.t3 3.3005
R328 source.n108 source.t6 3.3005
R329 source.n74 source.t12 3.3005
R330 source.n74 source.t10 3.3005
R331 source.n72 source.t15 3.3005
R332 source.n72 source.t17 3.3005
R333 source.n32 source.t16 3.3005
R334 source.n32 source.t9 3.3005
R335 source.n34 source.t13 3.3005
R336 source.n34 source.t8 3.3005
R337 source.n68 source.t0 3.3005
R338 source.n68 source.t18 3.3005
R339 source.n70 source.t5 3.3005
R340 source.n70 source.t4 3.3005
R341 source.n132 source.n131 2.71565
R342 source.n96 source.n95 2.71565
R343 source.n20 source.n19 2.71565
R344 source.n56 source.n55 2.71565
R345 source.n128 source.n118 1.93989
R346 source.n92 source.n82 1.93989
R347 source.n16 source.n6 1.93989
R348 source.n52 source.n42 1.93989
R349 source.n127 source.n120 1.16414
R350 source.n91 source.n84 1.16414
R351 source.n15 source.n8 1.16414
R352 source.n51 source.n44 1.16414
R353 source.n67 source.n35 0.914293
R354 source.n109 source.n107 0.914293
R355 source.n71 source.n69 0.888431
R356 source.n69 source.n67 0.888431
R357 source.n35 source.n33 0.888431
R358 source.n33 source.n31 0.888431
R359 source.n75 source.n73 0.888431
R360 source.n107 source.n75 0.888431
R361 source.n111 source.n109 0.888431
R362 source.n143 source.n111 0.888431
R363 source.n124 source.n123 0.388379
R364 source.n88 source.n87 0.388379
R365 source.n12 source.n11 0.388379
R366 source.n48 source.n47 0.388379
R367 source source.n144 0.188
R368 source.n126 source.n125 0.155672
R369 source.n126 source.n117 0.155672
R370 source.n133 source.n117 0.155672
R371 source.n134 source.n133 0.155672
R372 source.n134 source.n113 0.155672
R373 source.n141 source.n113 0.155672
R374 source.n90 source.n89 0.155672
R375 source.n90 source.n81 0.155672
R376 source.n97 source.n81 0.155672
R377 source.n98 source.n97 0.155672
R378 source.n98 source.n77 0.155672
R379 source.n105 source.n77 0.155672
R380 source.n29 source.n1 0.155672
R381 source.n22 source.n1 0.155672
R382 source.n22 source.n21 0.155672
R383 source.n21 source.n5 0.155672
R384 source.n14 source.n5 0.155672
R385 source.n14 source.n13 0.155672
R386 source.n65 source.n37 0.155672
R387 source.n58 source.n37 0.155672
R388 source.n58 source.n57 0.155672
R389 source.n57 source.n41 0.155672
R390 source.n50 source.n41 0.155672
R391 source.n50 source.n49 0.155672
R392 minus.n3 minus.t5 285.438
R393 minus.n17 minus.t7 285.438
R394 minus.n4 minus.t0 262.69
R395 minus.n6 minus.t2 262.69
R396 minus.n10 minus.t9 262.69
R397 minus.n12 minus.t1 262.69
R398 minus.n18 minus.t8 262.69
R399 minus.n20 minus.t3 262.69
R400 minus.n24 minus.t4 262.69
R401 minus.n26 minus.t6 262.69
R402 minus.n13 minus.n12 161.3
R403 minus.n11 minus.n0 161.3
R404 minus.n10 minus.n9 161.3
R405 minus.n8 minus.n1 161.3
R406 minus.n7 minus.n6 161.3
R407 minus.n5 minus.n2 161.3
R408 minus.n27 minus.n26 161.3
R409 minus.n25 minus.n14 161.3
R410 minus.n24 minus.n23 161.3
R411 minus.n22 minus.n15 161.3
R412 minus.n21 minus.n20 161.3
R413 minus.n19 minus.n16 161.3
R414 minus.n3 minus.n2 44.8741
R415 minus.n17 minus.n16 44.8741
R416 minus.n28 minus.n13 32.1085
R417 minus.n12 minus.n11 30.6732
R418 minus.n26 minus.n25 30.6732
R419 minus.n5 minus.n4 26.2914
R420 minus.n10 minus.n1 26.2914
R421 minus.n19 minus.n18 26.2914
R422 minus.n24 minus.n15 26.2914
R423 minus.n6 minus.n5 21.9096
R424 minus.n6 minus.n1 21.9096
R425 minus.n20 minus.n19 21.9096
R426 minus.n20 minus.n15 21.9096
R427 minus.n4 minus.n3 19.0667
R428 minus.n18 minus.n17 19.0667
R429 minus.n11 minus.n10 17.5278
R430 minus.n25 minus.n24 17.5278
R431 minus.n28 minus.n27 6.63876
R432 minus.n13 minus.n0 0.189894
R433 minus.n9 minus.n0 0.189894
R434 minus.n9 minus.n8 0.189894
R435 minus.n8 minus.n7 0.189894
R436 minus.n7 minus.n2 0.189894
R437 minus.n21 minus.n16 0.189894
R438 minus.n22 minus.n21 0.189894
R439 minus.n23 minus.n22 0.189894
R440 minus.n23 minus.n14 0.189894
R441 minus.n27 minus.n14 0.189894
R442 minus minus.n28 0.188
R443 drain_right.n26 drain_right.n0 289.615
R444 drain_right.n64 drain_right.n38 289.615
R445 drain_right.n11 drain_right.n10 185
R446 drain_right.n8 drain_right.n7 185
R447 drain_right.n17 drain_right.n16 185
R448 drain_right.n19 drain_right.n18 185
R449 drain_right.n4 drain_right.n3 185
R450 drain_right.n25 drain_right.n24 185
R451 drain_right.n27 drain_right.n26 185
R452 drain_right.n65 drain_right.n64 185
R453 drain_right.n63 drain_right.n62 185
R454 drain_right.n42 drain_right.n41 185
R455 drain_right.n57 drain_right.n56 185
R456 drain_right.n55 drain_right.n54 185
R457 drain_right.n46 drain_right.n45 185
R458 drain_right.n49 drain_right.n48 185
R459 drain_right.t2 drain_right.n9 147.661
R460 drain_right.t8 drain_right.n47 147.661
R461 drain_right.n10 drain_right.n7 104.615
R462 drain_right.n17 drain_right.n7 104.615
R463 drain_right.n18 drain_right.n17 104.615
R464 drain_right.n18 drain_right.n3 104.615
R465 drain_right.n25 drain_right.n3 104.615
R466 drain_right.n26 drain_right.n25 104.615
R467 drain_right.n64 drain_right.n63 104.615
R468 drain_right.n63 drain_right.n41 104.615
R469 drain_right.n56 drain_right.n41 104.615
R470 drain_right.n56 drain_right.n55 104.615
R471 drain_right.n55 drain_right.n45 104.615
R472 drain_right.n48 drain_right.n45 104.615
R473 drain_right.n37 drain_right.n35 68.0786
R474 drain_right.n34 drain_right.n33 67.8013
R475 drain_right.n37 drain_right.n36 67.1908
R476 drain_right.n32 drain_right.n31 67.1907
R477 drain_right.n10 drain_right.t2 52.3082
R478 drain_right.n48 drain_right.t8 52.3082
R479 drain_right.n32 drain_right.n30 49.7521
R480 drain_right.n69 drain_right.n68 48.8641
R481 drain_right drain_right.n34 26.0421
R482 drain_right.n11 drain_right.n9 15.6674
R483 drain_right.n49 drain_right.n47 15.6674
R484 drain_right.n12 drain_right.n8 12.8005
R485 drain_right.n50 drain_right.n46 12.8005
R486 drain_right.n16 drain_right.n15 12.0247
R487 drain_right.n54 drain_right.n53 12.0247
R488 drain_right.n19 drain_right.n6 11.249
R489 drain_right.n57 drain_right.n44 11.249
R490 drain_right.n20 drain_right.n4 10.4732
R491 drain_right.n58 drain_right.n42 10.4732
R492 drain_right.n24 drain_right.n23 9.69747
R493 drain_right.n62 drain_right.n61 9.69747
R494 drain_right.n30 drain_right.n29 9.45567
R495 drain_right.n68 drain_right.n67 9.45567
R496 drain_right.n29 drain_right.n28 9.3005
R497 drain_right.n2 drain_right.n1 9.3005
R498 drain_right.n23 drain_right.n22 9.3005
R499 drain_right.n21 drain_right.n20 9.3005
R500 drain_right.n6 drain_right.n5 9.3005
R501 drain_right.n15 drain_right.n14 9.3005
R502 drain_right.n13 drain_right.n12 9.3005
R503 drain_right.n67 drain_right.n66 9.3005
R504 drain_right.n40 drain_right.n39 9.3005
R505 drain_right.n61 drain_right.n60 9.3005
R506 drain_right.n59 drain_right.n58 9.3005
R507 drain_right.n44 drain_right.n43 9.3005
R508 drain_right.n53 drain_right.n52 9.3005
R509 drain_right.n51 drain_right.n50 9.3005
R510 drain_right.n27 drain_right.n2 8.92171
R511 drain_right.n65 drain_right.n40 8.92171
R512 drain_right.n28 drain_right.n0 8.14595
R513 drain_right.n66 drain_right.n38 8.14595
R514 drain_right drain_right.n69 6.09718
R515 drain_right.n30 drain_right.n0 5.81868
R516 drain_right.n68 drain_right.n38 5.81868
R517 drain_right.n28 drain_right.n27 5.04292
R518 drain_right.n66 drain_right.n65 5.04292
R519 drain_right.n13 drain_right.n9 4.38594
R520 drain_right.n51 drain_right.n47 4.38594
R521 drain_right.n24 drain_right.n2 4.26717
R522 drain_right.n62 drain_right.n40 4.26717
R523 drain_right.n23 drain_right.n4 3.49141
R524 drain_right.n61 drain_right.n42 3.49141
R525 drain_right.n33 drain_right.t5 3.3005
R526 drain_right.n33 drain_right.t3 3.3005
R527 drain_right.n31 drain_right.t1 3.3005
R528 drain_right.n31 drain_right.t6 3.3005
R529 drain_right.n35 drain_right.t9 3.3005
R530 drain_right.n35 drain_right.t4 3.3005
R531 drain_right.n36 drain_right.t0 3.3005
R532 drain_right.n36 drain_right.t7 3.3005
R533 drain_right.n20 drain_right.n19 2.71565
R534 drain_right.n58 drain_right.n57 2.71565
R535 drain_right.n16 drain_right.n6 1.93989
R536 drain_right.n54 drain_right.n44 1.93989
R537 drain_right.n15 drain_right.n8 1.16414
R538 drain_right.n53 drain_right.n46 1.16414
R539 drain_right.n69 drain_right.n37 0.888431
R540 drain_right.n12 drain_right.n11 0.388379
R541 drain_right.n50 drain_right.n49 0.388379
R542 drain_right.n34 drain_right.n32 0.167137
R543 drain_right.n14 drain_right.n13 0.155672
R544 drain_right.n14 drain_right.n5 0.155672
R545 drain_right.n21 drain_right.n5 0.155672
R546 drain_right.n22 drain_right.n21 0.155672
R547 drain_right.n22 drain_right.n1 0.155672
R548 drain_right.n29 drain_right.n1 0.155672
R549 drain_right.n67 drain_right.n39 0.155672
R550 drain_right.n60 drain_right.n39 0.155672
R551 drain_right.n60 drain_right.n59 0.155672
R552 drain_right.n59 drain_right.n43 0.155672
R553 drain_right.n52 drain_right.n43 0.155672
R554 drain_right.n52 drain_right.n51 0.155672
C0 drain_right source 8.46553f
C1 minus plus 4.46599f
C2 drain_right drain_left 0.967241f
C3 source plus 3.73563f
C4 source minus 3.72136f
C5 drain_left plus 3.76899f
C6 drain_right plus 0.346254f
C7 drain_left minus 0.171897f
C8 drain_right minus 3.57989f
C9 drain_left source 8.46826f
C10 drain_right a_n1952_n2088# 5.28012f
C11 drain_left a_n1952_n2088# 5.58467f
C12 source a_n1952_n2088# 4.155874f
C13 minus a_n1952_n2088# 7.144406f
C14 plus a_n1952_n2088# 8.5459f
C15 drain_right.n0 a_n1952_n2088# 0.034395f
C16 drain_right.n1 a_n1952_n2088# 0.02447f
C17 drain_right.n2 a_n1952_n2088# 0.013149f
C18 drain_right.n3 a_n1952_n2088# 0.03108f
C19 drain_right.n4 a_n1952_n2088# 0.013923f
C20 drain_right.n5 a_n1952_n2088# 0.02447f
C21 drain_right.n6 a_n1952_n2088# 0.013149f
C22 drain_right.n7 a_n1952_n2088# 0.03108f
C23 drain_right.n8 a_n1952_n2088# 0.013923f
C24 drain_right.n9 a_n1952_n2088# 0.104715f
C25 drain_right.t2 a_n1952_n2088# 0.050656f
C26 drain_right.n10 a_n1952_n2088# 0.02331f
C27 drain_right.n11 a_n1952_n2088# 0.018359f
C28 drain_right.n12 a_n1952_n2088# 0.013149f
C29 drain_right.n13 a_n1952_n2088# 0.582245f
C30 drain_right.n14 a_n1952_n2088# 0.02447f
C31 drain_right.n15 a_n1952_n2088# 0.013149f
C32 drain_right.n16 a_n1952_n2088# 0.013923f
C33 drain_right.n17 a_n1952_n2088# 0.03108f
C34 drain_right.n18 a_n1952_n2088# 0.03108f
C35 drain_right.n19 a_n1952_n2088# 0.013923f
C36 drain_right.n20 a_n1952_n2088# 0.013149f
C37 drain_right.n21 a_n1952_n2088# 0.02447f
C38 drain_right.n22 a_n1952_n2088# 0.02447f
C39 drain_right.n23 a_n1952_n2088# 0.013149f
C40 drain_right.n24 a_n1952_n2088# 0.013923f
C41 drain_right.n25 a_n1952_n2088# 0.03108f
C42 drain_right.n26 a_n1952_n2088# 0.067283f
C43 drain_right.n27 a_n1952_n2088# 0.013923f
C44 drain_right.n28 a_n1952_n2088# 0.013149f
C45 drain_right.n29 a_n1952_n2088# 0.056562f
C46 drain_right.n30 a_n1952_n2088# 0.056634f
C47 drain_right.t1 a_n1952_n2088# 0.116023f
C48 drain_right.t6 a_n1952_n2088# 0.116023f
C49 drain_right.n31 a_n1952_n2088# 0.967629f
C50 drain_right.n32 a_n1952_n2088# 0.400205f
C51 drain_right.t5 a_n1952_n2088# 0.116023f
C52 drain_right.t3 a_n1952_n2088# 0.116023f
C53 drain_right.n33 a_n1952_n2088# 0.970579f
C54 drain_right.n34 a_n1952_n2088# 1.20229f
C55 drain_right.t9 a_n1952_n2088# 0.116023f
C56 drain_right.t4 a_n1952_n2088# 0.116023f
C57 drain_right.n35 a_n1952_n2088# 0.972175f
C58 drain_right.t0 a_n1952_n2088# 0.116023f
C59 drain_right.t7 a_n1952_n2088# 0.116023f
C60 drain_right.n36 a_n1952_n2088# 0.967634f
C61 drain_right.n37 a_n1952_n2088# 0.682572f
C62 drain_right.n38 a_n1952_n2088# 0.034395f
C63 drain_right.n39 a_n1952_n2088# 0.02447f
C64 drain_right.n40 a_n1952_n2088# 0.013149f
C65 drain_right.n41 a_n1952_n2088# 0.03108f
C66 drain_right.n42 a_n1952_n2088# 0.013923f
C67 drain_right.n43 a_n1952_n2088# 0.02447f
C68 drain_right.n44 a_n1952_n2088# 0.013149f
C69 drain_right.n45 a_n1952_n2088# 0.03108f
C70 drain_right.n46 a_n1952_n2088# 0.013923f
C71 drain_right.n47 a_n1952_n2088# 0.104715f
C72 drain_right.t8 a_n1952_n2088# 0.050656f
C73 drain_right.n48 a_n1952_n2088# 0.02331f
C74 drain_right.n49 a_n1952_n2088# 0.018359f
C75 drain_right.n50 a_n1952_n2088# 0.013149f
C76 drain_right.n51 a_n1952_n2088# 0.582245f
C77 drain_right.n52 a_n1952_n2088# 0.02447f
C78 drain_right.n53 a_n1952_n2088# 0.013149f
C79 drain_right.n54 a_n1952_n2088# 0.013923f
C80 drain_right.n55 a_n1952_n2088# 0.03108f
C81 drain_right.n56 a_n1952_n2088# 0.03108f
C82 drain_right.n57 a_n1952_n2088# 0.013923f
C83 drain_right.n58 a_n1952_n2088# 0.013149f
C84 drain_right.n59 a_n1952_n2088# 0.02447f
C85 drain_right.n60 a_n1952_n2088# 0.02447f
C86 drain_right.n61 a_n1952_n2088# 0.013149f
C87 drain_right.n62 a_n1952_n2088# 0.013923f
C88 drain_right.n63 a_n1952_n2088# 0.03108f
C89 drain_right.n64 a_n1952_n2088# 0.067283f
C90 drain_right.n65 a_n1952_n2088# 0.013923f
C91 drain_right.n66 a_n1952_n2088# 0.013149f
C92 drain_right.n67 a_n1952_n2088# 0.056562f
C93 drain_right.n68 a_n1952_n2088# 0.054543f
C94 drain_right.n69 a_n1952_n2088# 0.342026f
C95 minus.n0 a_n1952_n2088# 0.043912f
C96 minus.n1 a_n1952_n2088# 0.009964f
C97 minus.t9 a_n1952_n2088# 0.534945f
C98 minus.n2 a_n1952_n2088# 0.18341f
C99 minus.t5 a_n1952_n2088# 0.554633f
C100 minus.n3 a_n1952_n2088# 0.231509f
C101 minus.t0 a_n1952_n2088# 0.534945f
C102 minus.n4 a_n1952_n2088# 0.251617f
C103 minus.n5 a_n1952_n2088# 0.009964f
C104 minus.t2 a_n1952_n2088# 0.534945f
C105 minus.n6 a_n1952_n2088# 0.247193f
C106 minus.n7 a_n1952_n2088# 0.043912f
C107 minus.n8 a_n1952_n2088# 0.043912f
C108 minus.n9 a_n1952_n2088# 0.043912f
C109 minus.n10 a_n1952_n2088# 0.247193f
C110 minus.n11 a_n1952_n2088# 0.009964f
C111 minus.t1 a_n1952_n2088# 0.534945f
C112 minus.n12 a_n1952_n2088# 0.244756f
C113 minus.n13 a_n1952_n2088# 1.28561f
C114 minus.n14 a_n1952_n2088# 0.043912f
C115 minus.n15 a_n1952_n2088# 0.009964f
C116 minus.n16 a_n1952_n2088# 0.18341f
C117 minus.t7 a_n1952_n2088# 0.554633f
C118 minus.n17 a_n1952_n2088# 0.231509f
C119 minus.t8 a_n1952_n2088# 0.534945f
C120 minus.n18 a_n1952_n2088# 0.251617f
C121 minus.n19 a_n1952_n2088# 0.009964f
C122 minus.t3 a_n1952_n2088# 0.534945f
C123 minus.n20 a_n1952_n2088# 0.247193f
C124 minus.n21 a_n1952_n2088# 0.043912f
C125 minus.n22 a_n1952_n2088# 0.043912f
C126 minus.n23 a_n1952_n2088# 0.043912f
C127 minus.t4 a_n1952_n2088# 0.534945f
C128 minus.n24 a_n1952_n2088# 0.247193f
C129 minus.n25 a_n1952_n2088# 0.009964f
C130 minus.t6 a_n1952_n2088# 0.534945f
C131 minus.n26 a_n1952_n2088# 0.244756f
C132 minus.n27 a_n1952_n2088# 0.301344f
C133 minus.n28 a_n1952_n2088# 1.57295f
C134 source.n0 a_n1952_n2088# 0.03848f
C135 source.n1 a_n1952_n2088# 0.027376f
C136 source.n2 a_n1952_n2088# 0.014711f
C137 source.n3 a_n1952_n2088# 0.034771f
C138 source.n4 a_n1952_n2088# 0.015576f
C139 source.n5 a_n1952_n2088# 0.027376f
C140 source.n6 a_n1952_n2088# 0.014711f
C141 source.n7 a_n1952_n2088# 0.034771f
C142 source.n8 a_n1952_n2088# 0.015576f
C143 source.n9 a_n1952_n2088# 0.117152f
C144 source.t14 a_n1952_n2088# 0.056673f
C145 source.n10 a_n1952_n2088# 0.026078f
C146 source.n11 a_n1952_n2088# 0.020539f
C147 source.n12 a_n1952_n2088# 0.014711f
C148 source.n13 a_n1952_n2088# 0.651398f
C149 source.n14 a_n1952_n2088# 0.027376f
C150 source.n15 a_n1952_n2088# 0.014711f
C151 source.n16 a_n1952_n2088# 0.015576f
C152 source.n17 a_n1952_n2088# 0.034771f
C153 source.n18 a_n1952_n2088# 0.034771f
C154 source.n19 a_n1952_n2088# 0.015576f
C155 source.n20 a_n1952_n2088# 0.014711f
C156 source.n21 a_n1952_n2088# 0.027376f
C157 source.n22 a_n1952_n2088# 0.027376f
C158 source.n23 a_n1952_n2088# 0.014711f
C159 source.n24 a_n1952_n2088# 0.015576f
C160 source.n25 a_n1952_n2088# 0.034771f
C161 source.n26 a_n1952_n2088# 0.075274f
C162 source.n27 a_n1952_n2088# 0.015576f
C163 source.n28 a_n1952_n2088# 0.014711f
C164 source.n29 a_n1952_n2088# 0.06328f
C165 source.n30 a_n1952_n2088# 0.042119f
C166 source.n31 a_n1952_n2088# 0.715173f
C167 source.t16 a_n1952_n2088# 0.129803f
C168 source.t9 a_n1952_n2088# 0.129803f
C169 source.n32 a_n1952_n2088# 1.01091f
C170 source.n33 a_n1952_n2088# 0.413283f
C171 source.t13 a_n1952_n2088# 0.129803f
C172 source.t8 a_n1952_n2088# 0.129803f
C173 source.n34 a_n1952_n2088# 1.01091f
C174 source.n35 a_n1952_n2088# 0.415565f
C175 source.n36 a_n1952_n2088# 0.03848f
C176 source.n37 a_n1952_n2088# 0.027376f
C177 source.n38 a_n1952_n2088# 0.014711f
C178 source.n39 a_n1952_n2088# 0.034771f
C179 source.n40 a_n1952_n2088# 0.015576f
C180 source.n41 a_n1952_n2088# 0.027376f
C181 source.n42 a_n1952_n2088# 0.014711f
C182 source.n43 a_n1952_n2088# 0.034771f
C183 source.n44 a_n1952_n2088# 0.015576f
C184 source.n45 a_n1952_n2088# 0.117152f
C185 source.t2 a_n1952_n2088# 0.056673f
C186 source.n46 a_n1952_n2088# 0.026078f
C187 source.n47 a_n1952_n2088# 0.020539f
C188 source.n48 a_n1952_n2088# 0.014711f
C189 source.n49 a_n1952_n2088# 0.651398f
C190 source.n50 a_n1952_n2088# 0.027376f
C191 source.n51 a_n1952_n2088# 0.014711f
C192 source.n52 a_n1952_n2088# 0.015576f
C193 source.n53 a_n1952_n2088# 0.034771f
C194 source.n54 a_n1952_n2088# 0.034771f
C195 source.n55 a_n1952_n2088# 0.015576f
C196 source.n56 a_n1952_n2088# 0.014711f
C197 source.n57 a_n1952_n2088# 0.027376f
C198 source.n58 a_n1952_n2088# 0.027376f
C199 source.n59 a_n1952_n2088# 0.014711f
C200 source.n60 a_n1952_n2088# 0.015576f
C201 source.n61 a_n1952_n2088# 0.034771f
C202 source.n62 a_n1952_n2088# 0.075274f
C203 source.n63 a_n1952_n2088# 0.015576f
C204 source.n64 a_n1952_n2088# 0.014711f
C205 source.n65 a_n1952_n2088# 0.06328f
C206 source.n66 a_n1952_n2088# 0.042119f
C207 source.n67 a_n1952_n2088# 0.182318f
C208 source.t0 a_n1952_n2088# 0.129803f
C209 source.t18 a_n1952_n2088# 0.129803f
C210 source.n68 a_n1952_n2088# 1.01091f
C211 source.n69 a_n1952_n2088# 0.413283f
C212 source.t5 a_n1952_n2088# 0.129803f
C213 source.t4 a_n1952_n2088# 0.129803f
C214 source.n70 a_n1952_n2088# 1.01091f
C215 source.n71 a_n1952_n2088# 1.38797f
C216 source.t15 a_n1952_n2088# 0.129803f
C217 source.t17 a_n1952_n2088# 0.129803f
C218 source.n72 a_n1952_n2088# 1.01091f
C219 source.n73 a_n1952_n2088# 1.38798f
C220 source.t12 a_n1952_n2088# 0.129803f
C221 source.t10 a_n1952_n2088# 0.129803f
C222 source.n74 a_n1952_n2088# 1.01091f
C223 source.n75 a_n1952_n2088# 0.41329f
C224 source.n76 a_n1952_n2088# 0.03848f
C225 source.n77 a_n1952_n2088# 0.027376f
C226 source.n78 a_n1952_n2088# 0.014711f
C227 source.n79 a_n1952_n2088# 0.034771f
C228 source.n80 a_n1952_n2088# 0.015576f
C229 source.n81 a_n1952_n2088# 0.027376f
C230 source.n82 a_n1952_n2088# 0.014711f
C231 source.n83 a_n1952_n2088# 0.034771f
C232 source.n84 a_n1952_n2088# 0.015576f
C233 source.n85 a_n1952_n2088# 0.117152f
C234 source.t11 a_n1952_n2088# 0.056673f
C235 source.n86 a_n1952_n2088# 0.026078f
C236 source.n87 a_n1952_n2088# 0.020539f
C237 source.n88 a_n1952_n2088# 0.014711f
C238 source.n89 a_n1952_n2088# 0.651398f
C239 source.n90 a_n1952_n2088# 0.027376f
C240 source.n91 a_n1952_n2088# 0.014711f
C241 source.n92 a_n1952_n2088# 0.015576f
C242 source.n93 a_n1952_n2088# 0.034771f
C243 source.n94 a_n1952_n2088# 0.034771f
C244 source.n95 a_n1952_n2088# 0.015576f
C245 source.n96 a_n1952_n2088# 0.014711f
C246 source.n97 a_n1952_n2088# 0.027376f
C247 source.n98 a_n1952_n2088# 0.027376f
C248 source.n99 a_n1952_n2088# 0.014711f
C249 source.n100 a_n1952_n2088# 0.015576f
C250 source.n101 a_n1952_n2088# 0.034771f
C251 source.n102 a_n1952_n2088# 0.075274f
C252 source.n103 a_n1952_n2088# 0.015576f
C253 source.n104 a_n1952_n2088# 0.014711f
C254 source.n105 a_n1952_n2088# 0.06328f
C255 source.n106 a_n1952_n2088# 0.042119f
C256 source.n107 a_n1952_n2088# 0.182318f
C257 source.t3 a_n1952_n2088# 0.129803f
C258 source.t6 a_n1952_n2088# 0.129803f
C259 source.n108 a_n1952_n2088# 1.01091f
C260 source.n109 a_n1952_n2088# 0.415572f
C261 source.t19 a_n1952_n2088# 0.129803f
C262 source.t1 a_n1952_n2088# 0.129803f
C263 source.n110 a_n1952_n2088# 1.01091f
C264 source.n111 a_n1952_n2088# 0.41329f
C265 source.n112 a_n1952_n2088# 0.03848f
C266 source.n113 a_n1952_n2088# 0.027376f
C267 source.n114 a_n1952_n2088# 0.014711f
C268 source.n115 a_n1952_n2088# 0.034771f
C269 source.n116 a_n1952_n2088# 0.015576f
C270 source.n117 a_n1952_n2088# 0.027376f
C271 source.n118 a_n1952_n2088# 0.014711f
C272 source.n119 a_n1952_n2088# 0.034771f
C273 source.n120 a_n1952_n2088# 0.015576f
C274 source.n121 a_n1952_n2088# 0.117152f
C275 source.t7 a_n1952_n2088# 0.056673f
C276 source.n122 a_n1952_n2088# 0.026078f
C277 source.n123 a_n1952_n2088# 0.020539f
C278 source.n124 a_n1952_n2088# 0.014711f
C279 source.n125 a_n1952_n2088# 0.651398f
C280 source.n126 a_n1952_n2088# 0.027376f
C281 source.n127 a_n1952_n2088# 0.014711f
C282 source.n128 a_n1952_n2088# 0.015576f
C283 source.n129 a_n1952_n2088# 0.034771f
C284 source.n130 a_n1952_n2088# 0.034771f
C285 source.n131 a_n1952_n2088# 0.015576f
C286 source.n132 a_n1952_n2088# 0.014711f
C287 source.n133 a_n1952_n2088# 0.027376f
C288 source.n134 a_n1952_n2088# 0.027376f
C289 source.n135 a_n1952_n2088# 0.014711f
C290 source.n136 a_n1952_n2088# 0.015576f
C291 source.n137 a_n1952_n2088# 0.034771f
C292 source.n138 a_n1952_n2088# 0.075274f
C293 source.n139 a_n1952_n2088# 0.015576f
C294 source.n140 a_n1952_n2088# 0.014711f
C295 source.n141 a_n1952_n2088# 0.06328f
C296 source.n142 a_n1952_n2088# 0.042119f
C297 source.n143 a_n1952_n2088# 0.321732f
C298 source.n144 a_n1952_n2088# 1.13536f
C299 drain_left.n0 a_n1952_n2088# 0.034689f
C300 drain_left.n1 a_n1952_n2088# 0.024679f
C301 drain_left.n2 a_n1952_n2088# 0.013262f
C302 drain_left.n3 a_n1952_n2088# 0.031346f
C303 drain_left.n4 a_n1952_n2088# 0.014042f
C304 drain_left.n5 a_n1952_n2088# 0.024679f
C305 drain_left.n6 a_n1952_n2088# 0.013262f
C306 drain_left.n7 a_n1952_n2088# 0.031346f
C307 drain_left.n8 a_n1952_n2088# 0.014042f
C308 drain_left.n9 a_n1952_n2088# 0.105611f
C309 drain_left.t1 a_n1952_n2088# 0.051089f
C310 drain_left.n10 a_n1952_n2088# 0.023509f
C311 drain_left.n11 a_n1952_n2088# 0.018516f
C312 drain_left.n12 a_n1952_n2088# 0.013262f
C313 drain_left.n13 a_n1952_n2088# 0.587223f
C314 drain_left.n14 a_n1952_n2088# 0.024679f
C315 drain_left.n15 a_n1952_n2088# 0.013262f
C316 drain_left.n16 a_n1952_n2088# 0.014042f
C317 drain_left.n17 a_n1952_n2088# 0.031346f
C318 drain_left.n18 a_n1952_n2088# 0.031346f
C319 drain_left.n19 a_n1952_n2088# 0.014042f
C320 drain_left.n20 a_n1952_n2088# 0.013262f
C321 drain_left.n21 a_n1952_n2088# 0.024679f
C322 drain_left.n22 a_n1952_n2088# 0.024679f
C323 drain_left.n23 a_n1952_n2088# 0.013262f
C324 drain_left.n24 a_n1952_n2088# 0.014042f
C325 drain_left.n25 a_n1952_n2088# 0.031346f
C326 drain_left.n26 a_n1952_n2088# 0.067858f
C327 drain_left.n27 a_n1952_n2088# 0.014042f
C328 drain_left.n28 a_n1952_n2088# 0.013262f
C329 drain_left.n29 a_n1952_n2088# 0.057045f
C330 drain_left.n30 a_n1952_n2088# 0.057118f
C331 drain_left.t6 a_n1952_n2088# 0.117015f
C332 drain_left.t2 a_n1952_n2088# 0.117015f
C333 drain_left.n31 a_n1952_n2088# 0.975903f
C334 drain_left.n32 a_n1952_n2088# 0.403627f
C335 drain_left.t7 a_n1952_n2088# 0.117015f
C336 drain_left.t0 a_n1952_n2088# 0.117015f
C337 drain_left.n33 a_n1952_n2088# 0.978878f
C338 drain_left.n34 a_n1952_n2088# 1.2626f
C339 drain_left.n35 a_n1952_n2088# 0.034689f
C340 drain_left.n36 a_n1952_n2088# 0.024679f
C341 drain_left.n37 a_n1952_n2088# 0.013262f
C342 drain_left.n38 a_n1952_n2088# 0.031346f
C343 drain_left.n39 a_n1952_n2088# 0.014042f
C344 drain_left.n40 a_n1952_n2088# 0.024679f
C345 drain_left.n41 a_n1952_n2088# 0.013262f
C346 drain_left.n42 a_n1952_n2088# 0.031346f
C347 drain_left.n43 a_n1952_n2088# 0.014042f
C348 drain_left.n44 a_n1952_n2088# 0.105611f
C349 drain_left.t5 a_n1952_n2088# 0.051089f
C350 drain_left.n45 a_n1952_n2088# 0.023509f
C351 drain_left.n46 a_n1952_n2088# 0.018516f
C352 drain_left.n47 a_n1952_n2088# 0.013262f
C353 drain_left.n48 a_n1952_n2088# 0.587223f
C354 drain_left.n49 a_n1952_n2088# 0.024679f
C355 drain_left.n50 a_n1952_n2088# 0.013262f
C356 drain_left.n51 a_n1952_n2088# 0.014042f
C357 drain_left.n52 a_n1952_n2088# 0.031346f
C358 drain_left.n53 a_n1952_n2088# 0.031346f
C359 drain_left.n54 a_n1952_n2088# 0.014042f
C360 drain_left.n55 a_n1952_n2088# 0.013262f
C361 drain_left.n56 a_n1952_n2088# 0.024679f
C362 drain_left.n57 a_n1952_n2088# 0.024679f
C363 drain_left.n58 a_n1952_n2088# 0.013262f
C364 drain_left.n59 a_n1952_n2088# 0.014042f
C365 drain_left.n60 a_n1952_n2088# 0.031346f
C366 drain_left.n61 a_n1952_n2088# 0.067858f
C367 drain_left.n62 a_n1952_n2088# 0.014042f
C368 drain_left.n63 a_n1952_n2088# 0.013262f
C369 drain_left.n64 a_n1952_n2088# 0.057045f
C370 drain_left.n65 a_n1952_n2088# 0.057118f
C371 drain_left.t4 a_n1952_n2088# 0.117015f
C372 drain_left.t8 a_n1952_n2088# 0.117015f
C373 drain_left.n66 a_n1952_n2088# 0.975907f
C374 drain_left.n67 a_n1952_n2088# 0.457548f
C375 drain_left.t3 a_n1952_n2088# 0.117015f
C376 drain_left.t9 a_n1952_n2088# 0.117015f
C377 drain_left.n68 a_n1952_n2088# 0.975903f
C378 drain_left.n69 a_n1952_n2088# 0.559819f
C379 plus.n0 a_n1952_n2088# 0.044994f
C380 plus.t3 a_n1952_n2088# 0.548137f
C381 plus.t8 a_n1952_n2088# 0.548137f
C382 plus.n1 a_n1952_n2088# 0.044994f
C383 plus.t1 a_n1952_n2088# 0.548137f
C384 plus.n2 a_n1952_n2088# 0.253289f
C385 plus.t4 a_n1952_n2088# 0.56831f
C386 plus.n3 a_n1952_n2088# 0.237218f
C387 plus.t9 a_n1952_n2088# 0.548137f
C388 plus.n4 a_n1952_n2088# 0.257822f
C389 plus.n5 a_n1952_n2088# 0.01021f
C390 plus.n6 a_n1952_n2088# 0.187933f
C391 plus.n7 a_n1952_n2088# 0.044994f
C392 plus.n8 a_n1952_n2088# 0.044994f
C393 plus.n9 a_n1952_n2088# 0.01021f
C394 plus.n10 a_n1952_n2088# 0.253289f
C395 plus.n11 a_n1952_n2088# 0.01021f
C396 plus.n12 a_n1952_n2088# 0.250792f
C397 plus.n13 a_n1952_n2088# 0.400825f
C398 plus.n14 a_n1952_n2088# 0.044994f
C399 plus.t2 a_n1952_n2088# 0.548137f
C400 plus.n15 a_n1952_n2088# 0.044994f
C401 plus.t0 a_n1952_n2088# 0.548137f
C402 plus.t5 a_n1952_n2088# 0.548137f
C403 plus.n16 a_n1952_n2088# 0.253289f
C404 plus.t6 a_n1952_n2088# 0.56831f
C405 plus.n17 a_n1952_n2088# 0.237218f
C406 plus.t7 a_n1952_n2088# 0.548137f
C407 plus.n18 a_n1952_n2088# 0.257822f
C408 plus.n19 a_n1952_n2088# 0.01021f
C409 plus.n20 a_n1952_n2088# 0.187933f
C410 plus.n21 a_n1952_n2088# 0.044994f
C411 plus.n22 a_n1952_n2088# 0.044994f
C412 plus.n23 a_n1952_n2088# 0.01021f
C413 plus.n24 a_n1952_n2088# 0.253289f
C414 plus.n25 a_n1952_n2088# 0.01021f
C415 plus.n26 a_n1952_n2088# 0.250792f
C416 plus.n27 a_n1952_n2088# 1.1913f
.ends

