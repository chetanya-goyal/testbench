* NGSPICE file created from diffpair264.ext - technology: sky130A

.subckt diffpair264 minus drain_right drain_left source plus
X0 source.t19 plus.t0 drain_left.t4 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 source.t18 plus.t1 drain_left.t8 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t6 plus.t2 source.t17 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 source.t4 minus.t0 drain_right.t9 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X4 source.t1 minus.t1 drain_right.t8 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X5 drain_left.t9 plus.t3 source.t16 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X6 source.t7 minus.t2 drain_right.t7 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X7 source.t15 plus.t4 drain_left.t7 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X8 a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X9 drain_right.t6 minus.t3 source.t9 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 drain_left.t2 plus.t5 source.t14 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X11 drain_left.t5 plus.t6 source.t13 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X12 a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X13 drain_left.t0 plus.t7 source.t12 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X14 drain_right.t5 minus.t4 source.t8 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 drain_right.t4 minus.t5 source.t2 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X16 drain_right.t3 minus.t6 source.t5 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X17 source.t11 plus.t8 drain_left.t3 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X18 a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X19 source.t6 minus.t7 drain_right.t2 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X20 drain_left.t1 plus.t9 source.t10 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X21 drain_right.t1 minus.t8 source.t0 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X22 a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X23 drain_right.t0 minus.t9 source.t3 a_n1412_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
R0 plus.n2 plus.t3 763.606
R1 plus.n8 plus.t5 763.606
R2 plus.n12 plus.t7 763.606
R3 plus.n18 plus.t9 763.606
R4 plus.n1 plus.t1 703.721
R5 plus.n5 plus.t6 703.721
R6 plus.n7 plus.t0 703.721
R7 plus.n11 plus.t4 703.721
R8 plus.n15 plus.t2 703.721
R9 plus.n17 plus.t8 703.721
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 26.0937
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 9.88686
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n26 drain_left.n0 289.615
R37 drain_left.n61 drain_left.n35 289.615
R38 drain_left.n11 drain_left.n10 185
R39 drain_left.n8 drain_left.n7 185
R40 drain_left.n17 drain_left.n16 185
R41 drain_left.n19 drain_left.n18 185
R42 drain_left.n4 drain_left.n3 185
R43 drain_left.n25 drain_left.n24 185
R44 drain_left.n27 drain_left.n26 185
R45 drain_left.n62 drain_left.n61 185
R46 drain_left.n60 drain_left.n59 185
R47 drain_left.n39 drain_left.n38 185
R48 drain_left.n54 drain_left.n53 185
R49 drain_left.n52 drain_left.n51 185
R50 drain_left.n43 drain_left.n42 185
R51 drain_left.n46 drain_left.n45 185
R52 drain_left.t1 drain_left.n9 147.661
R53 drain_left.t9 drain_left.n44 147.661
R54 drain_left.n10 drain_left.n7 104.615
R55 drain_left.n17 drain_left.n7 104.615
R56 drain_left.n18 drain_left.n17 104.615
R57 drain_left.n18 drain_left.n3 104.615
R58 drain_left.n25 drain_left.n3 104.615
R59 drain_left.n26 drain_left.n25 104.615
R60 drain_left.n61 drain_left.n60 104.615
R61 drain_left.n60 drain_left.n38 104.615
R62 drain_left.n53 drain_left.n38 104.615
R63 drain_left.n53 drain_left.n52 104.615
R64 drain_left.n52 drain_left.n42 104.615
R65 drain_left.n45 drain_left.n42 104.615
R66 drain_left.n34 drain_left.n33 67.5103
R67 drain_left.n67 drain_left.n66 67.1908
R68 drain_left.n69 drain_left.n68 67.1907
R69 drain_left.n32 drain_left.n31 67.1907
R70 drain_left.n10 drain_left.t1 52.3082
R71 drain_left.n45 drain_left.t9 52.3082
R72 drain_left.n32 drain_left.n30 49.3641
R73 drain_left.n67 drain_left.n65 49.3641
R74 drain_left drain_left.n34 24.9466
R75 drain_left.n11 drain_left.n9 15.6674
R76 drain_left.n46 drain_left.n44 15.6674
R77 drain_left.n12 drain_left.n8 12.8005
R78 drain_left.n47 drain_left.n43 12.8005
R79 drain_left.n16 drain_left.n15 12.0247
R80 drain_left.n51 drain_left.n50 12.0247
R81 drain_left.n19 drain_left.n6 11.249
R82 drain_left.n54 drain_left.n41 11.249
R83 drain_left.n20 drain_left.n4 10.4732
R84 drain_left.n55 drain_left.n39 10.4732
R85 drain_left.n24 drain_left.n23 9.69747
R86 drain_left.n59 drain_left.n58 9.69747
R87 drain_left.n30 drain_left.n29 9.45567
R88 drain_left.n65 drain_left.n64 9.45567
R89 drain_left.n29 drain_left.n28 9.3005
R90 drain_left.n2 drain_left.n1 9.3005
R91 drain_left.n23 drain_left.n22 9.3005
R92 drain_left.n21 drain_left.n20 9.3005
R93 drain_left.n6 drain_left.n5 9.3005
R94 drain_left.n15 drain_left.n14 9.3005
R95 drain_left.n13 drain_left.n12 9.3005
R96 drain_left.n64 drain_left.n63 9.3005
R97 drain_left.n37 drain_left.n36 9.3005
R98 drain_left.n58 drain_left.n57 9.3005
R99 drain_left.n56 drain_left.n55 9.3005
R100 drain_left.n41 drain_left.n40 9.3005
R101 drain_left.n50 drain_left.n49 9.3005
R102 drain_left.n48 drain_left.n47 9.3005
R103 drain_left.n27 drain_left.n2 8.92171
R104 drain_left.n62 drain_left.n37 8.92171
R105 drain_left.n28 drain_left.n0 8.14595
R106 drain_left.n63 drain_left.n35 8.14595
R107 drain_left drain_left.n69 6.15322
R108 drain_left.n30 drain_left.n0 5.81868
R109 drain_left.n65 drain_left.n35 5.81868
R110 drain_left.n28 drain_left.n27 5.04292
R111 drain_left.n63 drain_left.n62 5.04292
R112 drain_left.n13 drain_left.n9 4.38594
R113 drain_left.n48 drain_left.n44 4.38594
R114 drain_left.n24 drain_left.n2 4.26717
R115 drain_left.n59 drain_left.n37 4.26717
R116 drain_left.n23 drain_left.n4 3.49141
R117 drain_left.n58 drain_left.n39 3.49141
R118 drain_left.n33 drain_left.t7 3.3005
R119 drain_left.n33 drain_left.t0 3.3005
R120 drain_left.n31 drain_left.t3 3.3005
R121 drain_left.n31 drain_left.t6 3.3005
R122 drain_left.n68 drain_left.t4 3.3005
R123 drain_left.n68 drain_left.t2 3.3005
R124 drain_left.n66 drain_left.t8 3.3005
R125 drain_left.n66 drain_left.t5 3.3005
R126 drain_left.n20 drain_left.n19 2.71565
R127 drain_left.n55 drain_left.n54 2.71565
R128 drain_left.n16 drain_left.n6 1.93989
R129 drain_left.n51 drain_left.n41 1.93989
R130 drain_left.n15 drain_left.n8 1.16414
R131 drain_left.n50 drain_left.n43 1.16414
R132 drain_left.n69 drain_left.n67 0.5005
R133 drain_left.n12 drain_left.n11 0.388379
R134 drain_left.n47 drain_left.n46 0.388379
R135 drain_left.n14 drain_left.n13 0.155672
R136 drain_left.n14 drain_left.n5 0.155672
R137 drain_left.n21 drain_left.n5 0.155672
R138 drain_left.n22 drain_left.n21 0.155672
R139 drain_left.n22 drain_left.n1 0.155672
R140 drain_left.n29 drain_left.n1 0.155672
R141 drain_left.n64 drain_left.n36 0.155672
R142 drain_left.n57 drain_left.n36 0.155672
R143 drain_left.n57 drain_left.n56 0.155672
R144 drain_left.n56 drain_left.n40 0.155672
R145 drain_left.n49 drain_left.n40 0.155672
R146 drain_left.n49 drain_left.n48 0.155672
R147 drain_left.n34 drain_left.n32 0.070154
R148 source.n138 source.n112 289.615
R149 source.n102 source.n76 289.615
R150 source.n26 source.n0 289.615
R151 source.n62 source.n36 289.615
R152 source.n123 source.n122 185
R153 source.n120 source.n119 185
R154 source.n129 source.n128 185
R155 source.n131 source.n130 185
R156 source.n116 source.n115 185
R157 source.n137 source.n136 185
R158 source.n139 source.n138 185
R159 source.n87 source.n86 185
R160 source.n84 source.n83 185
R161 source.n93 source.n92 185
R162 source.n95 source.n94 185
R163 source.n80 source.n79 185
R164 source.n101 source.n100 185
R165 source.n103 source.n102 185
R166 source.n27 source.n26 185
R167 source.n25 source.n24 185
R168 source.n4 source.n3 185
R169 source.n19 source.n18 185
R170 source.n17 source.n16 185
R171 source.n8 source.n7 185
R172 source.n11 source.n10 185
R173 source.n63 source.n62 185
R174 source.n61 source.n60 185
R175 source.n40 source.n39 185
R176 source.n55 source.n54 185
R177 source.n53 source.n52 185
R178 source.n44 source.n43 185
R179 source.n47 source.n46 185
R180 source.t3 source.n121 147.661
R181 source.t12 source.n85 147.661
R182 source.t14 source.n9 147.661
R183 source.t5 source.n45 147.661
R184 source.n122 source.n119 104.615
R185 source.n129 source.n119 104.615
R186 source.n130 source.n129 104.615
R187 source.n130 source.n115 104.615
R188 source.n137 source.n115 104.615
R189 source.n138 source.n137 104.615
R190 source.n86 source.n83 104.615
R191 source.n93 source.n83 104.615
R192 source.n94 source.n93 104.615
R193 source.n94 source.n79 104.615
R194 source.n101 source.n79 104.615
R195 source.n102 source.n101 104.615
R196 source.n26 source.n25 104.615
R197 source.n25 source.n3 104.615
R198 source.n18 source.n3 104.615
R199 source.n18 source.n17 104.615
R200 source.n17 source.n7 104.615
R201 source.n10 source.n7 104.615
R202 source.n62 source.n61 104.615
R203 source.n61 source.n39 104.615
R204 source.n54 source.n39 104.615
R205 source.n54 source.n53 104.615
R206 source.n53 source.n43 104.615
R207 source.n46 source.n43 104.615
R208 source.n122 source.t3 52.3082
R209 source.n86 source.t12 52.3082
R210 source.n10 source.t14 52.3082
R211 source.n46 source.t5 52.3082
R212 source.n33 source.n32 50.512
R213 source.n35 source.n34 50.512
R214 source.n69 source.n68 50.512
R215 source.n71 source.n70 50.512
R216 source.n111 source.n110 50.5119
R217 source.n109 source.n108 50.5119
R218 source.n75 source.n74 50.5119
R219 source.n73 source.n72 50.5119
R220 source.n143 source.n142 32.1853
R221 source.n107 source.n106 32.1853
R222 source.n31 source.n30 32.1853
R223 source.n67 source.n66 32.1853
R224 source.n73 source.n71 17.7423
R225 source.n123 source.n121 15.6674
R226 source.n87 source.n85 15.6674
R227 source.n11 source.n9 15.6674
R228 source.n47 source.n45 15.6674
R229 source.n124 source.n120 12.8005
R230 source.n88 source.n84 12.8005
R231 source.n12 source.n8 12.8005
R232 source.n48 source.n44 12.8005
R233 source.n128 source.n127 12.0247
R234 source.n92 source.n91 12.0247
R235 source.n16 source.n15 12.0247
R236 source.n52 source.n51 12.0247
R237 source.n144 source.n31 11.7293
R238 source.n131 source.n118 11.249
R239 source.n95 source.n82 11.249
R240 source.n19 source.n6 11.249
R241 source.n55 source.n42 11.249
R242 source.n132 source.n116 10.4732
R243 source.n96 source.n80 10.4732
R244 source.n20 source.n4 10.4732
R245 source.n56 source.n40 10.4732
R246 source.n136 source.n135 9.69747
R247 source.n100 source.n99 9.69747
R248 source.n24 source.n23 9.69747
R249 source.n60 source.n59 9.69747
R250 source.n142 source.n141 9.45567
R251 source.n106 source.n105 9.45567
R252 source.n30 source.n29 9.45567
R253 source.n66 source.n65 9.45567
R254 source.n141 source.n140 9.3005
R255 source.n114 source.n113 9.3005
R256 source.n135 source.n134 9.3005
R257 source.n133 source.n132 9.3005
R258 source.n118 source.n117 9.3005
R259 source.n127 source.n126 9.3005
R260 source.n125 source.n124 9.3005
R261 source.n105 source.n104 9.3005
R262 source.n78 source.n77 9.3005
R263 source.n99 source.n98 9.3005
R264 source.n97 source.n96 9.3005
R265 source.n82 source.n81 9.3005
R266 source.n91 source.n90 9.3005
R267 source.n89 source.n88 9.3005
R268 source.n29 source.n28 9.3005
R269 source.n2 source.n1 9.3005
R270 source.n23 source.n22 9.3005
R271 source.n21 source.n20 9.3005
R272 source.n6 source.n5 9.3005
R273 source.n15 source.n14 9.3005
R274 source.n13 source.n12 9.3005
R275 source.n65 source.n64 9.3005
R276 source.n38 source.n37 9.3005
R277 source.n59 source.n58 9.3005
R278 source.n57 source.n56 9.3005
R279 source.n42 source.n41 9.3005
R280 source.n51 source.n50 9.3005
R281 source.n49 source.n48 9.3005
R282 source.n139 source.n114 8.92171
R283 source.n103 source.n78 8.92171
R284 source.n27 source.n2 8.92171
R285 source.n63 source.n38 8.92171
R286 source.n140 source.n112 8.14595
R287 source.n104 source.n76 8.14595
R288 source.n28 source.n0 8.14595
R289 source.n64 source.n36 8.14595
R290 source.n142 source.n112 5.81868
R291 source.n106 source.n76 5.81868
R292 source.n30 source.n0 5.81868
R293 source.n66 source.n36 5.81868
R294 source.n144 source.n143 5.51343
R295 source.n140 source.n139 5.04292
R296 source.n104 source.n103 5.04292
R297 source.n28 source.n27 5.04292
R298 source.n64 source.n63 5.04292
R299 source.n125 source.n121 4.38594
R300 source.n89 source.n85 4.38594
R301 source.n13 source.n9 4.38594
R302 source.n49 source.n45 4.38594
R303 source.n136 source.n114 4.26717
R304 source.n100 source.n78 4.26717
R305 source.n24 source.n2 4.26717
R306 source.n60 source.n38 4.26717
R307 source.n135 source.n116 3.49141
R308 source.n99 source.n80 3.49141
R309 source.n23 source.n4 3.49141
R310 source.n59 source.n40 3.49141
R311 source.n110 source.t9 3.3005
R312 source.n110 source.t7 3.3005
R313 source.n108 source.t2 3.3005
R314 source.n108 source.t6 3.3005
R315 source.n74 source.t17 3.3005
R316 source.n74 source.t15 3.3005
R317 source.n72 source.t10 3.3005
R318 source.n72 source.t11 3.3005
R319 source.n32 source.t13 3.3005
R320 source.n32 source.t19 3.3005
R321 source.n34 source.t16 3.3005
R322 source.n34 source.t18 3.3005
R323 source.n68 source.t8 3.3005
R324 source.n68 source.t1 3.3005
R325 source.n70 source.t0 3.3005
R326 source.n70 source.t4 3.3005
R327 source.n132 source.n131 2.71565
R328 source.n96 source.n95 2.71565
R329 source.n20 source.n19 2.71565
R330 source.n56 source.n55 2.71565
R331 source.n128 source.n118 1.93989
R332 source.n92 source.n82 1.93989
R333 source.n16 source.n6 1.93989
R334 source.n52 source.n42 1.93989
R335 source.n127 source.n120 1.16414
R336 source.n91 source.n84 1.16414
R337 source.n15 source.n8 1.16414
R338 source.n51 source.n44 1.16414
R339 source.n67 source.n35 0.720328
R340 source.n109 source.n107 0.720328
R341 source.n71 source.n69 0.5005
R342 source.n69 source.n67 0.5005
R343 source.n35 source.n33 0.5005
R344 source.n33 source.n31 0.5005
R345 source.n75 source.n73 0.5005
R346 source.n107 source.n75 0.5005
R347 source.n111 source.n109 0.5005
R348 source.n143 source.n111 0.5005
R349 source.n124 source.n123 0.388379
R350 source.n88 source.n87 0.388379
R351 source.n12 source.n11 0.388379
R352 source.n48 source.n47 0.388379
R353 source source.n144 0.188
R354 source.n126 source.n125 0.155672
R355 source.n126 source.n117 0.155672
R356 source.n133 source.n117 0.155672
R357 source.n134 source.n133 0.155672
R358 source.n134 source.n113 0.155672
R359 source.n141 source.n113 0.155672
R360 source.n90 source.n89 0.155672
R361 source.n90 source.n81 0.155672
R362 source.n97 source.n81 0.155672
R363 source.n98 source.n97 0.155672
R364 source.n98 source.n77 0.155672
R365 source.n105 source.n77 0.155672
R366 source.n29 source.n1 0.155672
R367 source.n22 source.n1 0.155672
R368 source.n22 source.n21 0.155672
R369 source.n21 source.n5 0.155672
R370 source.n14 source.n5 0.155672
R371 source.n14 source.n13 0.155672
R372 source.n65 source.n37 0.155672
R373 source.n58 source.n37 0.155672
R374 source.n58 source.n57 0.155672
R375 source.n57 source.n41 0.155672
R376 source.n50 source.n41 0.155672
R377 source.n50 source.n49 0.155672
R378 minus.n8 minus.t8 763.606
R379 minus.n2 minus.t6 763.606
R380 minus.n18 minus.t9 763.606
R381 minus.n12 minus.t5 763.606
R382 minus.n7 minus.t0 703.721
R383 minus.n5 minus.t4 703.721
R384 minus.n1 minus.t1 703.721
R385 minus.n17 minus.t2 703.721
R386 minus.n15 minus.t3 703.721
R387 minus.n11 minus.t7 703.721
R388 minus.n3 minus.n2 161.489
R389 minus.n13 minus.n12 161.489
R390 minus.n9 minus.n8 161.3
R391 minus.n6 minus.n0 161.3
R392 minus.n4 minus.n3 161.3
R393 minus.n19 minus.n18 161.3
R394 minus.n16 minus.n10 161.3
R395 minus.n14 minus.n13 161.3
R396 minus.n7 minus.n6 48.2005
R397 minus.n4 minus.n1 48.2005
R398 minus.n14 minus.n11 48.2005
R399 minus.n17 minus.n16 48.2005
R400 minus.n6 minus.n5 36.5157
R401 minus.n5 minus.n4 36.5157
R402 minus.n15 minus.n14 36.5157
R403 minus.n16 minus.n15 36.5157
R404 minus.n20 minus.n9 29.9399
R405 minus.n8 minus.n7 24.8308
R406 minus.n2 minus.n1 24.8308
R407 minus.n12 minus.n11 24.8308
R408 minus.n18 minus.n17 24.8308
R409 minus.n20 minus.n19 6.51565
R410 minus.n9 minus.n0 0.189894
R411 minus.n3 minus.n0 0.189894
R412 minus.n13 minus.n10 0.189894
R413 minus.n19 minus.n10 0.189894
R414 minus minus.n20 0.188
R415 drain_right.n26 drain_right.n0 289.615
R416 drain_right.n64 drain_right.n38 289.615
R417 drain_right.n11 drain_right.n10 185
R418 drain_right.n8 drain_right.n7 185
R419 drain_right.n17 drain_right.n16 185
R420 drain_right.n19 drain_right.n18 185
R421 drain_right.n4 drain_right.n3 185
R422 drain_right.n25 drain_right.n24 185
R423 drain_right.n27 drain_right.n26 185
R424 drain_right.n65 drain_right.n64 185
R425 drain_right.n63 drain_right.n62 185
R426 drain_right.n42 drain_right.n41 185
R427 drain_right.n57 drain_right.n56 185
R428 drain_right.n55 drain_right.n54 185
R429 drain_right.n46 drain_right.n45 185
R430 drain_right.n49 drain_right.n48 185
R431 drain_right.t4 drain_right.n9 147.661
R432 drain_right.t1 drain_right.n47 147.661
R433 drain_right.n10 drain_right.n7 104.615
R434 drain_right.n17 drain_right.n7 104.615
R435 drain_right.n18 drain_right.n17 104.615
R436 drain_right.n18 drain_right.n3 104.615
R437 drain_right.n25 drain_right.n3 104.615
R438 drain_right.n26 drain_right.n25 104.615
R439 drain_right.n64 drain_right.n63 104.615
R440 drain_right.n63 drain_right.n41 104.615
R441 drain_right.n56 drain_right.n41 104.615
R442 drain_right.n56 drain_right.n55 104.615
R443 drain_right.n55 drain_right.n45 104.615
R444 drain_right.n48 drain_right.n45 104.615
R445 drain_right.n37 drain_right.n35 67.6907
R446 drain_right.n34 drain_right.n33 67.5103
R447 drain_right.n37 drain_right.n36 67.1908
R448 drain_right.n32 drain_right.n31 67.1907
R449 drain_right.n10 drain_right.t4 52.3082
R450 drain_right.n48 drain_right.t1 52.3082
R451 drain_right.n32 drain_right.n30 49.3641
R452 drain_right.n69 drain_right.n68 48.8641
R453 drain_right drain_right.n34 24.3934
R454 drain_right.n11 drain_right.n9 15.6674
R455 drain_right.n49 drain_right.n47 15.6674
R456 drain_right.n12 drain_right.n8 12.8005
R457 drain_right.n50 drain_right.n46 12.8005
R458 drain_right.n16 drain_right.n15 12.0247
R459 drain_right.n54 drain_right.n53 12.0247
R460 drain_right.n19 drain_right.n6 11.249
R461 drain_right.n57 drain_right.n44 11.249
R462 drain_right.n20 drain_right.n4 10.4732
R463 drain_right.n58 drain_right.n42 10.4732
R464 drain_right.n24 drain_right.n23 9.69747
R465 drain_right.n62 drain_right.n61 9.69747
R466 drain_right.n30 drain_right.n29 9.45567
R467 drain_right.n68 drain_right.n67 9.45567
R468 drain_right.n29 drain_right.n28 9.3005
R469 drain_right.n2 drain_right.n1 9.3005
R470 drain_right.n23 drain_right.n22 9.3005
R471 drain_right.n21 drain_right.n20 9.3005
R472 drain_right.n6 drain_right.n5 9.3005
R473 drain_right.n15 drain_right.n14 9.3005
R474 drain_right.n13 drain_right.n12 9.3005
R475 drain_right.n67 drain_right.n66 9.3005
R476 drain_right.n40 drain_right.n39 9.3005
R477 drain_right.n61 drain_right.n60 9.3005
R478 drain_right.n59 drain_right.n58 9.3005
R479 drain_right.n44 drain_right.n43 9.3005
R480 drain_right.n53 drain_right.n52 9.3005
R481 drain_right.n51 drain_right.n50 9.3005
R482 drain_right.n27 drain_right.n2 8.92171
R483 drain_right.n65 drain_right.n40 8.92171
R484 drain_right.n28 drain_right.n0 8.14595
R485 drain_right.n66 drain_right.n38 8.14595
R486 drain_right drain_right.n69 5.90322
R487 drain_right.n30 drain_right.n0 5.81868
R488 drain_right.n68 drain_right.n38 5.81868
R489 drain_right.n28 drain_right.n27 5.04292
R490 drain_right.n66 drain_right.n65 5.04292
R491 drain_right.n13 drain_right.n9 4.38594
R492 drain_right.n51 drain_right.n47 4.38594
R493 drain_right.n24 drain_right.n2 4.26717
R494 drain_right.n62 drain_right.n40 4.26717
R495 drain_right.n23 drain_right.n4 3.49141
R496 drain_right.n61 drain_right.n42 3.49141
R497 drain_right.n33 drain_right.t7 3.3005
R498 drain_right.n33 drain_right.t0 3.3005
R499 drain_right.n31 drain_right.t2 3.3005
R500 drain_right.n31 drain_right.t6 3.3005
R501 drain_right.n35 drain_right.t8 3.3005
R502 drain_right.n35 drain_right.t3 3.3005
R503 drain_right.n36 drain_right.t9 3.3005
R504 drain_right.n36 drain_right.t5 3.3005
R505 drain_right.n20 drain_right.n19 2.71565
R506 drain_right.n58 drain_right.n57 2.71565
R507 drain_right.n16 drain_right.n6 1.93989
R508 drain_right.n54 drain_right.n44 1.93989
R509 drain_right.n15 drain_right.n8 1.16414
R510 drain_right.n53 drain_right.n46 1.16414
R511 drain_right.n69 drain_right.n37 0.5005
R512 drain_right.n12 drain_right.n11 0.388379
R513 drain_right.n50 drain_right.n49 0.388379
R514 drain_right.n14 drain_right.n13 0.155672
R515 drain_right.n14 drain_right.n5 0.155672
R516 drain_right.n21 drain_right.n5 0.155672
R517 drain_right.n22 drain_right.n21 0.155672
R518 drain_right.n22 drain_right.n1 0.155672
R519 drain_right.n29 drain_right.n1 0.155672
R520 drain_right.n67 drain_right.n39 0.155672
R521 drain_right.n60 drain_right.n39 0.155672
R522 drain_right.n60 drain_right.n59 0.155672
R523 drain_right.n59 drain_right.n43 0.155672
R524 drain_right.n52 drain_right.n43 0.155672
R525 drain_right.n52 drain_right.n51 0.155672
R526 drain_right.n34 drain_right.n32 0.070154
C0 drain_left minus 0.171039f
C1 source drain_right 12.4314f
C2 drain_left drain_right 0.691431f
C3 minus drain_right 1.96878f
C4 source plus 1.85702f
C5 drain_left plus 2.10149f
C6 minus plus 3.79895f
C7 source drain_left 12.4381f
C8 source minus 1.84266f
C9 plus drain_right 0.289092f
C10 drain_right a_n1412_n2088# 4.78087f
C11 drain_left a_n1412_n2088# 5.29846f
C12 source a_n1412_n2088# 3.849231f
C13 minus a_n1412_n2088# 4.96121f
C14 plus a_n1412_n2088# 6.15288f
C15 drain_right.n0 a_n1412_n2088# 0.037075f
C16 drain_right.n1 a_n1412_n2088# 0.026377f
C17 drain_right.n2 a_n1412_n2088# 0.014174f
C18 drain_right.n3 a_n1412_n2088# 0.033502f
C19 drain_right.n4 a_n1412_n2088# 0.015008f
C20 drain_right.n5 a_n1412_n2088# 0.026377f
C21 drain_right.n6 a_n1412_n2088# 0.014174f
C22 drain_right.n7 a_n1412_n2088# 0.033502f
C23 drain_right.n8 a_n1412_n2088# 0.015008f
C24 drain_right.n9 a_n1412_n2088# 0.112876f
C25 drain_right.t4 a_n1412_n2088# 0.054604f
C26 drain_right.n10 a_n1412_n2088# 0.025127f
C27 drain_right.n11 a_n1412_n2088# 0.019789f
C28 drain_right.n12 a_n1412_n2088# 0.014174f
C29 drain_right.n13 a_n1412_n2088# 0.627619f
C30 drain_right.n14 a_n1412_n2088# 0.026377f
C31 drain_right.n15 a_n1412_n2088# 0.014174f
C32 drain_right.n16 a_n1412_n2088# 0.015008f
C33 drain_right.n17 a_n1412_n2088# 0.033502f
C34 drain_right.n18 a_n1412_n2088# 0.033502f
C35 drain_right.n19 a_n1412_n2088# 0.015008f
C36 drain_right.n20 a_n1412_n2088# 0.014174f
C37 drain_right.n21 a_n1412_n2088# 0.026377f
C38 drain_right.n22 a_n1412_n2088# 0.026377f
C39 drain_right.n23 a_n1412_n2088# 0.014174f
C40 drain_right.n24 a_n1412_n2088# 0.015008f
C41 drain_right.n25 a_n1412_n2088# 0.033502f
C42 drain_right.n26 a_n1412_n2088# 0.072526f
C43 drain_right.n27 a_n1412_n2088# 0.015008f
C44 drain_right.n28 a_n1412_n2088# 0.014174f
C45 drain_right.n29 a_n1412_n2088# 0.06097f
C46 drain_right.n30 a_n1412_n2088# 0.059739f
C47 drain_right.t2 a_n1412_n2088# 0.125064f
C48 drain_right.t6 a_n1412_n2088# 0.125064f
C49 drain_right.n31 a_n1412_n2088# 1.04304f
C50 drain_right.n32 a_n1412_n2088# 0.363625f
C51 drain_right.t7 a_n1412_n2088# 0.125064f
C52 drain_right.t0 a_n1412_n2088# 0.125064f
C53 drain_right.n33 a_n1412_n2088# 1.04444f
C54 drain_right.n34 a_n1412_n2088# 1.06461f
C55 drain_right.t8 a_n1412_n2088# 0.125064f
C56 drain_right.t3 a_n1412_n2088# 0.125064f
C57 drain_right.n35 a_n1412_n2088# 1.04532f
C58 drain_right.t9 a_n1412_n2088# 0.125064f
C59 drain_right.t5 a_n1412_n2088# 0.125064f
C60 drain_right.n36 a_n1412_n2088# 1.04304f
C61 drain_right.n37 a_n1412_n2088# 0.60649f
C62 drain_right.n38 a_n1412_n2088# 0.037075f
C63 drain_right.n39 a_n1412_n2088# 0.026377f
C64 drain_right.n40 a_n1412_n2088# 0.014174f
C65 drain_right.n41 a_n1412_n2088# 0.033502f
C66 drain_right.n42 a_n1412_n2088# 0.015008f
C67 drain_right.n43 a_n1412_n2088# 0.026377f
C68 drain_right.n44 a_n1412_n2088# 0.014174f
C69 drain_right.n45 a_n1412_n2088# 0.033502f
C70 drain_right.n46 a_n1412_n2088# 0.015008f
C71 drain_right.n47 a_n1412_n2088# 0.112876f
C72 drain_right.t1 a_n1412_n2088# 0.054604f
C73 drain_right.n48 a_n1412_n2088# 0.025127f
C74 drain_right.n49 a_n1412_n2088# 0.019789f
C75 drain_right.n50 a_n1412_n2088# 0.014174f
C76 drain_right.n51 a_n1412_n2088# 0.627619f
C77 drain_right.n52 a_n1412_n2088# 0.026377f
C78 drain_right.n53 a_n1412_n2088# 0.014174f
C79 drain_right.n54 a_n1412_n2088# 0.015008f
C80 drain_right.n55 a_n1412_n2088# 0.033502f
C81 drain_right.n56 a_n1412_n2088# 0.033502f
C82 drain_right.n57 a_n1412_n2088# 0.015008f
C83 drain_right.n58 a_n1412_n2088# 0.014174f
C84 drain_right.n59 a_n1412_n2088# 0.026377f
C85 drain_right.n60 a_n1412_n2088# 0.026377f
C86 drain_right.n61 a_n1412_n2088# 0.014174f
C87 drain_right.n62 a_n1412_n2088# 0.015008f
C88 drain_right.n63 a_n1412_n2088# 0.033502f
C89 drain_right.n64 a_n1412_n2088# 0.072526f
C90 drain_right.n65 a_n1412_n2088# 0.015008f
C91 drain_right.n66 a_n1412_n2088# 0.014174f
C92 drain_right.n67 a_n1412_n2088# 0.06097f
C93 drain_right.n68 a_n1412_n2088# 0.058794f
C94 drain_right.n69 a_n1412_n2088# 0.31051f
C95 minus.n0 a_n1412_n2088# 0.027502f
C96 minus.t8 a_n1412_n2088# 0.122092f
C97 minus.t0 a_n1412_n2088# 0.117537f
C98 minus.t4 a_n1412_n2088# 0.117537f
C99 minus.t1 a_n1412_n2088# 0.117537f
C100 minus.n1 a_n1412_n2088# 0.055364f
C101 minus.t6 a_n1412_n2088# 0.122092f
C102 minus.n2 a_n1412_n2088# 0.064046f
C103 minus.n3 a_n1412_n2088# 0.064625f
C104 minus.n4 a_n1412_n2088# 0.01048f
C105 minus.n5 a_n1412_n2088# 0.055364f
C106 minus.n6 a_n1412_n2088# 0.01048f
C107 minus.n7 a_n1412_n2088# 0.055364f
C108 minus.n8 a_n1412_n2088# 0.064003f
C109 minus.n9 a_n1412_n2088# 0.713397f
C110 minus.n10 a_n1412_n2088# 0.027502f
C111 minus.t2 a_n1412_n2088# 0.117537f
C112 minus.t3 a_n1412_n2088# 0.117537f
C113 minus.t7 a_n1412_n2088# 0.117537f
C114 minus.n11 a_n1412_n2088# 0.055364f
C115 minus.t5 a_n1412_n2088# 0.122092f
C116 minus.n12 a_n1412_n2088# 0.064046f
C117 minus.n13 a_n1412_n2088# 0.064625f
C118 minus.n14 a_n1412_n2088# 0.01048f
C119 minus.n15 a_n1412_n2088# 0.055364f
C120 minus.n16 a_n1412_n2088# 0.01048f
C121 minus.n17 a_n1412_n2088# 0.055364f
C122 minus.t9 a_n1412_n2088# 0.122092f
C123 minus.n18 a_n1412_n2088# 0.064003f
C124 minus.n19 a_n1412_n2088# 0.180814f
C125 minus.n20 a_n1412_n2088# 0.879681f
C126 source.n0 a_n1412_n2088# 0.040473f
C127 source.n1 a_n1412_n2088# 0.028795f
C128 source.n2 a_n1412_n2088# 0.015473f
C129 source.n3 a_n1412_n2088# 0.036572f
C130 source.n4 a_n1412_n2088# 0.016383f
C131 source.n5 a_n1412_n2088# 0.028795f
C132 source.n6 a_n1412_n2088# 0.015473f
C133 source.n7 a_n1412_n2088# 0.036572f
C134 source.n8 a_n1412_n2088# 0.016383f
C135 source.n9 a_n1412_n2088# 0.12322f
C136 source.t14 a_n1412_n2088# 0.059608f
C137 source.n10 a_n1412_n2088# 0.027429f
C138 source.n11 a_n1412_n2088# 0.021603f
C139 source.n12 a_n1412_n2088# 0.015473f
C140 source.n13 a_n1412_n2088# 0.685138f
C141 source.n14 a_n1412_n2088# 0.028795f
C142 source.n15 a_n1412_n2088# 0.015473f
C143 source.n16 a_n1412_n2088# 0.016383f
C144 source.n17 a_n1412_n2088# 0.036572f
C145 source.n18 a_n1412_n2088# 0.036572f
C146 source.n19 a_n1412_n2088# 0.016383f
C147 source.n20 a_n1412_n2088# 0.015473f
C148 source.n21 a_n1412_n2088# 0.028795f
C149 source.n22 a_n1412_n2088# 0.028795f
C150 source.n23 a_n1412_n2088# 0.015473f
C151 source.n24 a_n1412_n2088# 0.016383f
C152 source.n25 a_n1412_n2088# 0.036572f
C153 source.n26 a_n1412_n2088# 0.079173f
C154 source.n27 a_n1412_n2088# 0.016383f
C155 source.n28 a_n1412_n2088# 0.015473f
C156 source.n29 a_n1412_n2088# 0.066557f
C157 source.n30 a_n1412_n2088# 0.0443f
C158 source.n31 a_n1412_n2088# 0.690603f
C159 source.t13 a_n1412_n2088# 0.136526f
C160 source.t19 a_n1412_n2088# 0.136526f
C161 source.n32 a_n1412_n2088# 1.06328f
C162 source.n33 a_n1412_n2088# 0.362704f
C163 source.t16 a_n1412_n2088# 0.136526f
C164 source.t18 a_n1412_n2088# 0.136526f
C165 source.n34 a_n1412_n2088# 1.06328f
C166 source.n35 a_n1412_n2088# 0.3831f
C167 source.n36 a_n1412_n2088# 0.040473f
C168 source.n37 a_n1412_n2088# 0.028795f
C169 source.n38 a_n1412_n2088# 0.015473f
C170 source.n39 a_n1412_n2088# 0.036572f
C171 source.n40 a_n1412_n2088# 0.016383f
C172 source.n41 a_n1412_n2088# 0.028795f
C173 source.n42 a_n1412_n2088# 0.015473f
C174 source.n43 a_n1412_n2088# 0.036572f
C175 source.n44 a_n1412_n2088# 0.016383f
C176 source.n45 a_n1412_n2088# 0.12322f
C177 source.t5 a_n1412_n2088# 0.059608f
C178 source.n46 a_n1412_n2088# 0.027429f
C179 source.n47 a_n1412_n2088# 0.021603f
C180 source.n48 a_n1412_n2088# 0.015473f
C181 source.n49 a_n1412_n2088# 0.685138f
C182 source.n50 a_n1412_n2088# 0.028795f
C183 source.n51 a_n1412_n2088# 0.015473f
C184 source.n52 a_n1412_n2088# 0.016383f
C185 source.n53 a_n1412_n2088# 0.036572f
C186 source.n54 a_n1412_n2088# 0.036572f
C187 source.n55 a_n1412_n2088# 0.016383f
C188 source.n56 a_n1412_n2088# 0.015473f
C189 source.n57 a_n1412_n2088# 0.028795f
C190 source.n58 a_n1412_n2088# 0.028795f
C191 source.n59 a_n1412_n2088# 0.015473f
C192 source.n60 a_n1412_n2088# 0.016383f
C193 source.n61 a_n1412_n2088# 0.036572f
C194 source.n62 a_n1412_n2088# 0.079173f
C195 source.n63 a_n1412_n2088# 0.016383f
C196 source.n64 a_n1412_n2088# 0.015473f
C197 source.n65 a_n1412_n2088# 0.066557f
C198 source.n66 a_n1412_n2088# 0.0443f
C199 source.n67 a_n1412_n2088# 0.137771f
C200 source.t8 a_n1412_n2088# 0.136526f
C201 source.t1 a_n1412_n2088# 0.136526f
C202 source.n68 a_n1412_n2088# 1.06328f
C203 source.n69 a_n1412_n2088# 0.362704f
C204 source.t0 a_n1412_n2088# 0.136526f
C205 source.t4 a_n1412_n2088# 0.136526f
C206 source.n70 a_n1412_n2088# 1.06328f
C207 source.n71 a_n1412_n2088# 1.35188f
C208 source.t10 a_n1412_n2088# 0.136526f
C209 source.t11 a_n1412_n2088# 0.136526f
C210 source.n72 a_n1412_n2088# 1.06327f
C211 source.n73 a_n1412_n2088# 1.35189f
C212 source.t17 a_n1412_n2088# 0.136526f
C213 source.t15 a_n1412_n2088# 0.136526f
C214 source.n74 a_n1412_n2088# 1.06327f
C215 source.n75 a_n1412_n2088# 0.362711f
C216 source.n76 a_n1412_n2088# 0.040473f
C217 source.n77 a_n1412_n2088# 0.028795f
C218 source.n78 a_n1412_n2088# 0.015473f
C219 source.n79 a_n1412_n2088# 0.036572f
C220 source.n80 a_n1412_n2088# 0.016383f
C221 source.n81 a_n1412_n2088# 0.028795f
C222 source.n82 a_n1412_n2088# 0.015473f
C223 source.n83 a_n1412_n2088# 0.036572f
C224 source.n84 a_n1412_n2088# 0.016383f
C225 source.n85 a_n1412_n2088# 0.12322f
C226 source.t12 a_n1412_n2088# 0.059608f
C227 source.n86 a_n1412_n2088# 0.027429f
C228 source.n87 a_n1412_n2088# 0.021603f
C229 source.n88 a_n1412_n2088# 0.015473f
C230 source.n89 a_n1412_n2088# 0.685138f
C231 source.n90 a_n1412_n2088# 0.028795f
C232 source.n91 a_n1412_n2088# 0.015473f
C233 source.n92 a_n1412_n2088# 0.016383f
C234 source.n93 a_n1412_n2088# 0.036572f
C235 source.n94 a_n1412_n2088# 0.036572f
C236 source.n95 a_n1412_n2088# 0.016383f
C237 source.n96 a_n1412_n2088# 0.015473f
C238 source.n97 a_n1412_n2088# 0.028795f
C239 source.n98 a_n1412_n2088# 0.028795f
C240 source.n99 a_n1412_n2088# 0.015473f
C241 source.n100 a_n1412_n2088# 0.016383f
C242 source.n101 a_n1412_n2088# 0.036572f
C243 source.n102 a_n1412_n2088# 0.079173f
C244 source.n103 a_n1412_n2088# 0.016383f
C245 source.n104 a_n1412_n2088# 0.015473f
C246 source.n105 a_n1412_n2088# 0.066557f
C247 source.n106 a_n1412_n2088# 0.0443f
C248 source.n107 a_n1412_n2088# 0.137771f
C249 source.t2 a_n1412_n2088# 0.136526f
C250 source.t6 a_n1412_n2088# 0.136526f
C251 source.n108 a_n1412_n2088# 1.06327f
C252 source.n109 a_n1412_n2088# 0.383107f
C253 source.t9 a_n1412_n2088# 0.136526f
C254 source.t7 a_n1412_n2088# 0.136526f
C255 source.n110 a_n1412_n2088# 1.06327f
C256 source.n111 a_n1412_n2088# 0.362711f
C257 source.n112 a_n1412_n2088# 0.040473f
C258 source.n113 a_n1412_n2088# 0.028795f
C259 source.n114 a_n1412_n2088# 0.015473f
C260 source.n115 a_n1412_n2088# 0.036572f
C261 source.n116 a_n1412_n2088# 0.016383f
C262 source.n117 a_n1412_n2088# 0.028795f
C263 source.n118 a_n1412_n2088# 0.015473f
C264 source.n119 a_n1412_n2088# 0.036572f
C265 source.n120 a_n1412_n2088# 0.016383f
C266 source.n121 a_n1412_n2088# 0.12322f
C267 source.t3 a_n1412_n2088# 0.059608f
C268 source.n122 a_n1412_n2088# 0.027429f
C269 source.n123 a_n1412_n2088# 0.021603f
C270 source.n124 a_n1412_n2088# 0.015473f
C271 source.n125 a_n1412_n2088# 0.685138f
C272 source.n126 a_n1412_n2088# 0.028795f
C273 source.n127 a_n1412_n2088# 0.015473f
C274 source.n128 a_n1412_n2088# 0.016383f
C275 source.n129 a_n1412_n2088# 0.036572f
C276 source.n130 a_n1412_n2088# 0.036572f
C277 source.n131 a_n1412_n2088# 0.016383f
C278 source.n132 a_n1412_n2088# 0.015473f
C279 source.n133 a_n1412_n2088# 0.028795f
C280 source.n134 a_n1412_n2088# 0.028795f
C281 source.n135 a_n1412_n2088# 0.015473f
C282 source.n136 a_n1412_n2088# 0.016383f
C283 source.n137 a_n1412_n2088# 0.036572f
C284 source.n138 a_n1412_n2088# 0.079173f
C285 source.n139 a_n1412_n2088# 0.016383f
C286 source.n140 a_n1412_n2088# 0.015473f
C287 source.n141 a_n1412_n2088# 0.066557f
C288 source.n142 a_n1412_n2088# 0.0443f
C289 source.n143 a_n1412_n2088# 0.273919f
C290 source.n144 a_n1412_n2088# 1.17628f
C291 drain_left.n0 a_n1412_n2088# 0.042997f
C292 drain_left.n1 a_n1412_n2088# 0.03059f
C293 drain_left.n2 a_n1412_n2088# 0.016438f
C294 drain_left.n3 a_n1412_n2088# 0.038853f
C295 drain_left.n4 a_n1412_n2088# 0.017404f
C296 drain_left.n5 a_n1412_n2088# 0.03059f
C297 drain_left.n6 a_n1412_n2088# 0.016438f
C298 drain_left.n7 a_n1412_n2088# 0.038853f
C299 drain_left.n8 a_n1412_n2088# 0.017404f
C300 drain_left.n9 a_n1412_n2088# 0.130902f
C301 drain_left.t1 a_n1412_n2088# 0.063325f
C302 drain_left.n10 a_n1412_n2088# 0.029139f
C303 drain_left.n11 a_n1412_n2088# 0.02295f
C304 drain_left.n12 a_n1412_n2088# 0.016438f
C305 drain_left.n13 a_n1412_n2088# 0.727853f
C306 drain_left.n14 a_n1412_n2088# 0.03059f
C307 drain_left.n15 a_n1412_n2088# 0.016438f
C308 drain_left.n16 a_n1412_n2088# 0.017404f
C309 drain_left.n17 a_n1412_n2088# 0.038853f
C310 drain_left.n18 a_n1412_n2088# 0.038853f
C311 drain_left.n19 a_n1412_n2088# 0.017404f
C312 drain_left.n20 a_n1412_n2088# 0.016438f
C313 drain_left.n21 a_n1412_n2088# 0.03059f
C314 drain_left.n22 a_n1412_n2088# 0.03059f
C315 drain_left.n23 a_n1412_n2088# 0.016438f
C316 drain_left.n24 a_n1412_n2088# 0.017404f
C317 drain_left.n25 a_n1412_n2088# 0.038853f
C318 drain_left.n26 a_n1412_n2088# 0.084109f
C319 drain_left.n27 a_n1412_n2088# 0.017404f
C320 drain_left.n28 a_n1412_n2088# 0.016438f
C321 drain_left.n29 a_n1412_n2088# 0.070707f
C322 drain_left.n30 a_n1412_n2088# 0.069279f
C323 drain_left.t3 a_n1412_n2088# 0.145038f
C324 drain_left.t6 a_n1412_n2088# 0.145038f
C325 drain_left.n31 a_n1412_n2088# 1.20961f
C326 drain_left.n32 a_n1412_n2088# 0.421698f
C327 drain_left.t7 a_n1412_n2088# 0.145038f
C328 drain_left.t0 a_n1412_n2088# 0.145038f
C329 drain_left.n33 a_n1412_n2088# 1.21124f
C330 drain_left.n34 a_n1412_n2088# 1.29719f
C331 drain_left.n35 a_n1412_n2088# 0.042997f
C332 drain_left.n36 a_n1412_n2088# 0.03059f
C333 drain_left.n37 a_n1412_n2088# 0.016438f
C334 drain_left.n38 a_n1412_n2088# 0.038853f
C335 drain_left.n39 a_n1412_n2088# 0.017404f
C336 drain_left.n40 a_n1412_n2088# 0.03059f
C337 drain_left.n41 a_n1412_n2088# 0.016438f
C338 drain_left.n42 a_n1412_n2088# 0.038853f
C339 drain_left.n43 a_n1412_n2088# 0.017404f
C340 drain_left.n44 a_n1412_n2088# 0.130902f
C341 drain_left.t9 a_n1412_n2088# 0.063325f
C342 drain_left.n45 a_n1412_n2088# 0.029139f
C343 drain_left.n46 a_n1412_n2088# 0.02295f
C344 drain_left.n47 a_n1412_n2088# 0.016438f
C345 drain_left.n48 a_n1412_n2088# 0.727853f
C346 drain_left.n49 a_n1412_n2088# 0.03059f
C347 drain_left.n50 a_n1412_n2088# 0.016438f
C348 drain_left.n51 a_n1412_n2088# 0.017404f
C349 drain_left.n52 a_n1412_n2088# 0.038853f
C350 drain_left.n53 a_n1412_n2088# 0.038853f
C351 drain_left.n54 a_n1412_n2088# 0.017404f
C352 drain_left.n55 a_n1412_n2088# 0.016438f
C353 drain_left.n56 a_n1412_n2088# 0.03059f
C354 drain_left.n57 a_n1412_n2088# 0.03059f
C355 drain_left.n58 a_n1412_n2088# 0.016438f
C356 drain_left.n59 a_n1412_n2088# 0.017404f
C357 drain_left.n60 a_n1412_n2088# 0.038853f
C358 drain_left.n61 a_n1412_n2088# 0.084109f
C359 drain_left.n62 a_n1412_n2088# 0.017404f
C360 drain_left.n63 a_n1412_n2088# 0.016438f
C361 drain_left.n64 a_n1412_n2088# 0.070707f
C362 drain_left.n65 a_n1412_n2088# 0.069279f
C363 drain_left.t8 a_n1412_n2088# 0.145038f
C364 drain_left.t5 a_n1412_n2088# 0.145038f
C365 drain_left.n66 a_n1412_n2088# 1.20962f
C366 drain_left.n67 a_n1412_n2088# 0.453928f
C367 drain_left.t4 a_n1412_n2088# 0.145038f
C368 drain_left.t2 a_n1412_n2088# 0.145038f
C369 drain_left.n68 a_n1412_n2088# 1.20961f
C370 drain_left.n69 a_n1412_n2088# 0.599341f
C371 plus.n0 a_n1412_n2088# 0.043335f
C372 plus.t0 a_n1412_n2088# 0.185202f
C373 plus.t6 a_n1412_n2088# 0.185202f
C374 plus.t1 a_n1412_n2088# 0.185202f
C375 plus.n1 a_n1412_n2088# 0.087237f
C376 plus.t3 a_n1412_n2088# 0.192379f
C377 plus.n2 a_n1412_n2088# 0.100917f
C378 plus.n3 a_n1412_n2088# 0.10183f
C379 plus.n4 a_n1412_n2088# 0.016513f
C380 plus.n5 a_n1412_n2088# 0.087237f
C381 plus.n6 a_n1412_n2088# 0.016513f
C382 plus.n7 a_n1412_n2088# 0.087237f
C383 plus.t5 a_n1412_n2088# 0.192379f
C384 plus.n8 a_n1412_n2088# 0.100848f
C385 plus.n9 a_n1412_n2088# 0.372998f
C386 plus.n10 a_n1412_n2088# 0.043335f
C387 plus.t9 a_n1412_n2088# 0.192379f
C388 plus.t8 a_n1412_n2088# 0.185202f
C389 plus.t2 a_n1412_n2088# 0.185202f
C390 plus.t4 a_n1412_n2088# 0.185202f
C391 plus.n11 a_n1412_n2088# 0.087237f
C392 plus.t7 a_n1412_n2088# 0.192379f
C393 plus.n12 a_n1412_n2088# 0.100917f
C394 plus.n13 a_n1412_n2088# 0.10183f
C395 plus.n14 a_n1412_n2088# 0.016513f
C396 plus.n15 a_n1412_n2088# 0.087237f
C397 plus.n16 a_n1412_n2088# 0.016513f
C398 plus.n17 a_n1412_n2088# 0.087237f
C399 plus.n18 a_n1412_n2088# 0.100848f
C400 plus.n19 a_n1412_n2088# 1.01642f
.ends

