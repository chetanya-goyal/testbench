* NGSPICE file created from diffpair393.ext - technology: sky130A

.subckt diffpair393 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t8 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X1 source.t7 plus.t0 drain_left.t7 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X2 a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X3 source.t5 plus.t1 drain_left.t6 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 drain_right.t6 minus.t1 source.t9 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X5 a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X6 a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X7 drain_right.t5 minus.t2 source.t10 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 drain_left.t5 plus.t2 source.t0 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X9 source.t11 minus.t3 drain_right.t4 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 source.t12 minus.t4 drain_right.t3 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 drain_right.t2 minus.t5 source.t13 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X12 source.t14 minus.t6 drain_right.t1 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X13 a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X14 drain_left.t4 plus.t3 source.t6 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X15 drain_left.t3 plus.t4 source.t4 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X16 source.t15 minus.t7 drain_right.t0 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X17 source.t2 plus.t5 drain_left.t2 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X18 drain_left.t1 plus.t6 source.t1 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 source.t3 plus.t7 drain_left.t0 a_n1846_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n2 minus.t5 340.832
R1 minus.n10 minus.t7 340.832
R2 minus.n1 minus.t3 320.229
R3 minus.n4 minus.t2 320.229
R4 minus.n6 minus.t6 320.229
R5 minus.n9 minus.t1 320.229
R6 minus.n12 minus.t4 320.229
R7 minus.n14 minus.t0 320.229
R8 minus.n7 minus.n6 161.3
R9 minus.n5 minus.n0 161.3
R10 minus.n15 minus.n14 161.3
R11 minus.n13 minus.n8 161.3
R12 minus.n4 minus.n3 80.6037
R13 minus.n12 minus.n11 80.6037
R14 minus.n4 minus.n1 48.2005
R15 minus.n12 minus.n9 48.2005
R16 minus.n5 minus.n4 41.6278
R17 minus.n13 minus.n12 41.6278
R18 minus.n16 minus.n7 33.9929
R19 minus.n3 minus.n2 31.6158
R20 minus.n11 minus.n10 31.6158
R21 minus.n2 minus.n1 17.6494
R22 minus.n10 minus.n9 17.6494
R23 minus.n16 minus.n15 6.65202
R24 minus.n6 minus.n5 6.57323
R25 minus.n14 minus.n13 6.57323
R26 minus.n3 minus.n0 0.285035
R27 minus.n11 minus.n8 0.285035
R28 minus.n7 minus.n0 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 source.n3 source.t3 51.0588
R32 source.n4 source.t13 51.0588
R33 source.n7 source.t14 51.0588
R34 source.n15 source.t8 51.0586
R35 source.n12 source.t15 51.0586
R36 source.n11 source.t6 51.0586
R37 source.n8 source.t7 51.0586
R38 source.n0 source.t4 51.0586
R39 source.n2 source.n1 48.8588
R40 source.n6 source.n5 48.8588
R41 source.n14 source.n13 48.8586
R42 source.n10 source.n9 48.8586
R43 source.n8 source.n7 19.9891
R44 source.n16 source.n0 14.2391
R45 source.n16 source.n15 5.7505
R46 source.n13 source.t9 2.2005
R47 source.n13 source.t12 2.2005
R48 source.n9 source.t0 2.2005
R49 source.n9 source.t5 2.2005
R50 source.n1 source.t1 2.2005
R51 source.n1 source.t2 2.2005
R52 source.n5 source.t10 2.2005
R53 source.n5 source.t11 2.2005
R54 source.n7 source.n6 0.974638
R55 source.n6 source.n4 0.974638
R56 source.n3 source.n2 0.974638
R57 source.n2 source.n0 0.974638
R58 source.n10 source.n8 0.974638
R59 source.n11 source.n10 0.974638
R60 source.n14 source.n12 0.974638
R61 source.n15 source.n14 0.974638
R62 source.n4 source.n3 0.470328
R63 source.n12 source.n11 0.470328
R64 source source.n16 0.188
R65 drain_right.n5 drain_right.n3 66.5116
R66 drain_right.n2 drain_right.n1 65.9691
R67 drain_right.n2 drain_right.n0 65.9691
R68 drain_right.n5 drain_right.n4 65.5376
R69 drain_right drain_right.n2 27.9506
R70 drain_right drain_right.n5 6.62735
R71 drain_right.n1 drain_right.t3 2.2005
R72 drain_right.n1 drain_right.t7 2.2005
R73 drain_right.n0 drain_right.t0 2.2005
R74 drain_right.n0 drain_right.t6 2.2005
R75 drain_right.n3 drain_right.t4 2.2005
R76 drain_right.n3 drain_right.t2 2.2005
R77 drain_right.n4 drain_right.t1 2.2005
R78 drain_right.n4 drain_right.t5 2.2005
R79 plus.n2 plus.t7 340.832
R80 plus.n10 plus.t3 340.832
R81 plus.n6 plus.t4 320.229
R82 plus.n4 plus.t5 320.229
R83 plus.n3 plus.t6 320.229
R84 plus.n14 plus.t0 320.229
R85 plus.n12 plus.t2 320.229
R86 plus.n11 plus.t1 320.229
R87 plus.n5 plus.n0 161.3
R88 plus.n7 plus.n6 161.3
R89 plus.n13 plus.n8 161.3
R90 plus.n15 plus.n14 161.3
R91 plus.n4 plus.n1 80.6037
R92 plus.n12 plus.n9 80.6037
R93 plus.n4 plus.n3 48.2005
R94 plus.n12 plus.n11 48.2005
R95 plus.n5 plus.n4 41.6278
R96 plus.n13 plus.n12 41.6278
R97 plus.n2 plus.n1 31.6158
R98 plus.n10 plus.n9 31.6158
R99 plus plus.n15 29.0104
R100 plus.n3 plus.n2 17.6494
R101 plus.n11 plus.n10 17.6494
R102 plus plus.n7 11.1596
R103 plus.n6 plus.n5 6.57323
R104 plus.n14 plus.n13 6.57323
R105 plus.n1 plus.n0 0.285035
R106 plus.n9 plus.n8 0.285035
R107 plus.n7 plus.n0 0.189894
R108 plus.n15 plus.n8 0.189894
R109 drain_left.n5 drain_left.n3 66.5117
R110 drain_left.n2 drain_left.n1 65.9691
R111 drain_left.n2 drain_left.n0 65.9691
R112 drain_left.n5 drain_left.n4 65.5374
R113 drain_left drain_left.n2 28.5038
R114 drain_left drain_left.n5 6.62735
R115 drain_left.n1 drain_left.t6 2.2005
R116 drain_left.n1 drain_left.t4 2.2005
R117 drain_left.n0 drain_left.t7 2.2005
R118 drain_left.n0 drain_left.t5 2.2005
R119 drain_left.n4 drain_left.t2 2.2005
R120 drain_left.n4 drain_left.t3 2.2005
R121 drain_left.n3 drain_left.t0 2.2005
R122 drain_left.n3 drain_left.t1 2.2005
C0 drain_right drain_left 0.873724f
C1 drain_left plus 4.70367f
C2 source drain_left 8.52236f
C3 minus drain_right 4.52442f
C4 minus plus 4.8877f
C5 source minus 4.43434f
C6 drain_right plus 0.333957f
C7 source drain_right 8.52475f
C8 source plus 4.44838f
C9 minus drain_left 0.17159f
C10 drain_right a_n1846_n2688# 5.15781f
C11 drain_left a_n1846_n2688# 5.43163f
C12 source a_n1846_n2688# 7.35702f
C13 minus a_n1846_n2688# 6.954864f
C14 plus a_n1846_n2688# 8.42878f
C15 drain_left.t7 a_n1846_n2688# 0.187833f
C16 drain_left.t5 a_n1846_n2688# 0.187833f
C17 drain_left.n0 a_n1846_n2688# 1.64516f
C18 drain_left.t6 a_n1846_n2688# 0.187833f
C19 drain_left.t4 a_n1846_n2688# 0.187833f
C20 drain_left.n1 a_n1846_n2688# 1.64516f
C21 drain_left.n2 a_n1846_n2688# 1.82749f
C22 drain_left.t0 a_n1846_n2688# 0.187833f
C23 drain_left.t1 a_n1846_n2688# 0.187833f
C24 drain_left.n3 a_n1846_n2688# 1.6486f
C25 drain_left.t2 a_n1846_n2688# 0.187833f
C26 drain_left.t3 a_n1846_n2688# 0.187833f
C27 drain_left.n4 a_n1846_n2688# 1.64291f
C28 drain_left.n5 a_n1846_n2688# 0.996478f
C29 plus.n0 a_n1846_n2688# 0.057215f
C30 plus.t4 a_n1846_n2688# 0.885361f
C31 plus.t5 a_n1846_n2688# 0.885361f
C32 plus.n1 a_n1846_n2688# 0.245403f
C33 plus.t6 a_n1846_n2688# 0.885361f
C34 plus.t7 a_n1846_n2688# 0.907845f
C35 plus.n2 a_n1846_n2688# 0.353061f
C36 plus.n3 a_n1846_n2688# 0.380739f
C37 plus.n4 a_n1846_n2688# 0.380041f
C38 plus.n5 a_n1846_n2688# 0.00973f
C39 plus.n6 a_n1846_n2688# 0.363966f
C40 plus.n7 a_n1846_n2688# 0.436926f
C41 plus.n8 a_n1846_n2688# 0.057215f
C42 plus.t0 a_n1846_n2688# 0.885361f
C43 plus.n9 a_n1846_n2688# 0.245403f
C44 plus.t2 a_n1846_n2688# 0.885361f
C45 plus.t3 a_n1846_n2688# 0.907845f
C46 plus.n10 a_n1846_n2688# 0.353061f
C47 plus.t1 a_n1846_n2688# 0.885361f
C48 plus.n11 a_n1846_n2688# 0.380739f
C49 plus.n12 a_n1846_n2688# 0.380041f
C50 plus.n13 a_n1846_n2688# 0.00973f
C51 plus.n14 a_n1846_n2688# 0.363966f
C52 plus.n15 a_n1846_n2688# 1.20294f
C53 drain_right.t0 a_n1846_n2688# 0.186447f
C54 drain_right.t6 a_n1846_n2688# 0.186447f
C55 drain_right.n0 a_n1846_n2688# 1.63302f
C56 drain_right.t3 a_n1846_n2688# 0.186447f
C57 drain_right.t7 a_n1846_n2688# 0.186447f
C58 drain_right.n1 a_n1846_n2688# 1.63302f
C59 drain_right.n2 a_n1846_n2688# 1.76001f
C60 drain_right.t4 a_n1846_n2688# 0.186447f
C61 drain_right.t2 a_n1846_n2688# 0.186447f
C62 drain_right.n3 a_n1846_n2688# 1.63642f
C63 drain_right.t1 a_n1846_n2688# 0.186447f
C64 drain_right.t5 a_n1846_n2688# 0.186447f
C65 drain_right.n4 a_n1846_n2688# 1.63079f
C66 drain_right.n5 a_n1846_n2688# 0.989121f
C67 source.t4 a_n1846_n2688# 1.53044f
C68 source.n0 a_n1846_n2688# 0.926896f
C69 source.t1 a_n1846_n2688# 0.143522f
C70 source.t2 a_n1846_n2688# 0.143522f
C71 source.n1 a_n1846_n2688# 1.20147f
C72 source.n2 a_n1846_n2688# 0.314768f
C73 source.t3 a_n1846_n2688# 1.53045f
C74 source.n3 a_n1846_n2688# 0.344426f
C75 source.t13 a_n1846_n2688# 1.53045f
C76 source.n4 a_n1846_n2688# 0.344426f
C77 source.t10 a_n1846_n2688# 0.143522f
C78 source.t11 a_n1846_n2688# 0.143522f
C79 source.n5 a_n1846_n2688# 1.20147f
C80 source.n6 a_n1846_n2688# 0.314768f
C81 source.t14 a_n1846_n2688# 1.53045f
C82 source.n7 a_n1846_n2688# 1.22931f
C83 source.t7 a_n1846_n2688# 1.53044f
C84 source.n8 a_n1846_n2688# 1.22932f
C85 source.t0 a_n1846_n2688# 0.143522f
C86 source.t5 a_n1846_n2688# 0.143522f
C87 source.n9 a_n1846_n2688# 1.20147f
C88 source.n10 a_n1846_n2688# 0.314771f
C89 source.t6 a_n1846_n2688# 1.53044f
C90 source.n11 a_n1846_n2688# 0.344429f
C91 source.t15 a_n1846_n2688# 1.53044f
C92 source.n12 a_n1846_n2688# 0.344429f
C93 source.t9 a_n1846_n2688# 0.143522f
C94 source.t12 a_n1846_n2688# 0.143522f
C95 source.n13 a_n1846_n2688# 1.20147f
C96 source.n14 a_n1846_n2688# 0.314771f
C97 source.t8 a_n1846_n2688# 1.53044f
C98 source.n15 a_n1846_n2688# 0.480434f
C99 source.n16 a_n1846_n2688# 1.06566f
C100 minus.n0 a_n1846_n2688# 0.05605f
C101 minus.t3 a_n1846_n2688# 0.867341f
C102 minus.n1 a_n1846_n2688# 0.37299f
C103 minus.t2 a_n1846_n2688# 0.867341f
C104 minus.t5 a_n1846_n2688# 0.889368f
C105 minus.n2 a_n1846_n2688# 0.345875f
C106 minus.n3 a_n1846_n2688# 0.240409f
C107 minus.n4 a_n1846_n2688# 0.372306f
C108 minus.n5 a_n1846_n2688# 0.009532f
C109 minus.t6 a_n1846_n2688# 0.867341f
C110 minus.n6 a_n1846_n2688# 0.356558f
C111 minus.n7 a_n1846_n2688# 1.34921f
C112 minus.n8 a_n1846_n2688# 0.05605f
C113 minus.t1 a_n1846_n2688# 0.867341f
C114 minus.n9 a_n1846_n2688# 0.37299f
C115 minus.t7 a_n1846_n2688# 0.889368f
C116 minus.n10 a_n1846_n2688# 0.345875f
C117 minus.n11 a_n1846_n2688# 0.240409f
C118 minus.t4 a_n1846_n2688# 0.867341f
C119 minus.n12 a_n1846_n2688# 0.372306f
C120 minus.n13 a_n1846_n2688# 0.009532f
C121 minus.t0 a_n1846_n2688# 0.867341f
C122 minus.n14 a_n1846_n2688# 0.356558f
C123 minus.n15 a_n1846_n2688# 0.289554f
C124 minus.n16 a_n1846_n2688# 1.64343f
.ends

