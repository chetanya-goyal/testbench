* NGSPICE file created from diffpair205.ext - technology: sky130A

.subckt diffpair205 minus drain_right drain_left source plus
X0 a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X1 a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X2 a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X3 source.t20 minus.t0 drain_right.t1 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X4 source.t19 minus.t1 drain_right.t6 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X5 drain_left.t11 plus.t0 source.t3 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X6 source.t2 plus.t1 drain_left.t10 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 source.t18 minus.t2 drain_right.t2 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X8 drain_right.t5 minus.t3 source.t17 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X9 drain_right.t9 minus.t4 source.t16 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X10 drain_left.t9 plus.t2 source.t7 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X11 drain_right.t7 minus.t5 source.t15 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X12 drain_left.t8 plus.t3 source.t1 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X13 drain_right.t8 minus.t6 source.t14 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X14 drain_right.t3 minus.t7 source.t13 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X15 source.t6 plus.t4 drain_left.t7 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X16 source.t12 minus.t8 drain_right.t0 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X17 source.t22 plus.t5 drain_left.t6 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X18 a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X19 source.t21 plus.t6 drain_left.t5 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X20 drain_right.t4 minus.t9 source.t11 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X21 drain_left.t4 plus.t7 source.t8 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X22 source.t10 minus.t10 drain_right.t11 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X23 source.t9 minus.t11 drain_right.t10 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X24 drain_left.t3 plus.t8 source.t0 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X25 source.t23 plus.t9 drain_left.t2 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X26 source.t5 plus.t10 drain_left.t1 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X27 drain_left.t0 plus.t11 source.t4 a_n1878_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
R0 minus.n3 minus.t9 249.835
R1 minus.n17 minus.t2 249.835
R2 minus.n4 minus.t1 223.167
R3 minus.n5 minus.t5 223.167
R4 minus.n1 minus.t11 223.167
R5 minus.n10 minus.t3 223.167
R6 minus.n12 minus.t8 223.167
R7 minus.n18 minus.t6 223.167
R8 minus.n19 minus.t0 223.167
R9 minus.n15 minus.t4 223.167
R10 minus.n24 minus.t10 223.167
R11 minus.n26 minus.t7 223.167
R12 minus.n13 minus.n12 161.3
R13 minus.n11 minus.n0 161.3
R14 minus.n10 minus.n9 161.3
R15 minus.n8 minus.n1 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n2 161.3
R18 minus.n27 minus.n26 161.3
R19 minus.n25 minus.n14 161.3
R20 minus.n24 minus.n23 161.3
R21 minus.n22 minus.n15 161.3
R22 minus.n21 minus.n20 161.3
R23 minus.n19 minus.n16 161.3
R24 minus.n5 minus.n4 48.2005
R25 minus.n10 minus.n1 48.2005
R26 minus.n19 minus.n18 48.2005
R27 minus.n24 minus.n15 48.2005
R28 minus.n12 minus.n11 47.4702
R29 minus.n26 minus.n25 47.4702
R30 minus.n3 minus.n2 45.1192
R31 minus.n17 minus.n16 45.1192
R32 minus.n28 minus.n13 29.4475
R33 minus.n6 minus.n1 24.1005
R34 minus.n6 minus.n5 24.1005
R35 minus.n20 minus.n19 24.1005
R36 minus.n20 minus.n15 24.1005
R37 minus.n4 minus.n3 13.6377
R38 minus.n18 minus.n17 13.6377
R39 minus.n28 minus.n27 6.5308
R40 minus.n11 minus.n10 0.730803
R41 minus.n25 minus.n24 0.730803
R42 minus.n13 minus.n0 0.189894
R43 minus.n9 minus.n0 0.189894
R44 minus.n9 minus.n8 0.189894
R45 minus.n8 minus.n7 0.189894
R46 minus.n7 minus.n2 0.189894
R47 minus.n21 minus.n16 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n14 0.189894
R51 minus.n27 minus.n14 0.189894
R52 minus minus.n28 0.188
R53 drain_right.n6 drain_right.n4 80.4886
R54 drain_right.n3 drain_right.n2 80.4332
R55 drain_right.n3 drain_right.n0 80.4332
R56 drain_right.n6 drain_right.n5 79.7731
R57 drain_right.n8 drain_right.n7 79.7731
R58 drain_right.n3 drain_right.n1 79.773
R59 drain_right drain_right.n3 23.5733
R60 drain_right.n1 drain_right.t1 6.6005
R61 drain_right.n1 drain_right.t9 6.6005
R62 drain_right.n2 drain_right.t11 6.6005
R63 drain_right.n2 drain_right.t3 6.6005
R64 drain_right.n0 drain_right.t2 6.6005
R65 drain_right.n0 drain_right.t8 6.6005
R66 drain_right.n4 drain_right.t6 6.6005
R67 drain_right.n4 drain_right.t4 6.6005
R68 drain_right.n5 drain_right.t10 6.6005
R69 drain_right.n5 drain_right.t7 6.6005
R70 drain_right.n7 drain_right.t0 6.6005
R71 drain_right.n7 drain_right.t5 6.6005
R72 drain_right drain_right.n8 6.36873
R73 drain_right.n8 drain_right.n6 0.716017
R74 source.n0 source.t4 69.6943
R75 source.n5 source.t2 69.6943
R76 source.n6 source.t11 69.6943
R77 source.n11 source.t12 69.6943
R78 source.n23 source.t13 69.6942
R79 source.n18 source.t18 69.6942
R80 source.n17 source.t7 69.6942
R81 source.n12 source.t6 69.6942
R82 source.n2 source.n1 63.0943
R83 source.n4 source.n3 63.0943
R84 source.n8 source.n7 63.0943
R85 source.n10 source.n9 63.0943
R86 source.n22 source.n21 63.0942
R87 source.n20 source.n19 63.0942
R88 source.n16 source.n15 63.0942
R89 source.n14 source.n13 63.0942
R90 source.n12 source.n11 15.1851
R91 source.n24 source.n0 9.56437
R92 source.n21 source.t16 6.6005
R93 source.n21 source.t10 6.6005
R94 source.n19 source.t14 6.6005
R95 source.n19 source.t20 6.6005
R96 source.n15 source.t3 6.6005
R97 source.n15 source.t22 6.6005
R98 source.n13 source.t0 6.6005
R99 source.n13 source.t21 6.6005
R100 source.n1 source.t1 6.6005
R101 source.n1 source.t23 6.6005
R102 source.n3 source.t8 6.6005
R103 source.n3 source.t5 6.6005
R104 source.n7 source.t15 6.6005
R105 source.n7 source.t19 6.6005
R106 source.n9 source.t17 6.6005
R107 source.n9 source.t9 6.6005
R108 source.n24 source.n23 5.62119
R109 source.n11 source.n10 0.716017
R110 source.n10 source.n8 0.716017
R111 source.n8 source.n6 0.716017
R112 source.n5 source.n4 0.716017
R113 source.n4 source.n2 0.716017
R114 source.n2 source.n0 0.716017
R115 source.n14 source.n12 0.716017
R116 source.n16 source.n14 0.716017
R117 source.n17 source.n16 0.716017
R118 source.n20 source.n18 0.716017
R119 source.n22 source.n20 0.716017
R120 source.n23 source.n22 0.716017
R121 source.n6 source.n5 0.470328
R122 source.n18 source.n17 0.470328
R123 source source.n24 0.188
R124 plus.n5 plus.t1 249.835
R125 plus.n19 plus.t2 249.835
R126 plus.n12 plus.t11 223.167
R127 plus.n10 plus.t9 223.167
R128 plus.n9 plus.t3 223.167
R129 plus.n3 plus.t10 223.167
R130 plus.n4 plus.t7 223.167
R131 plus.n26 plus.t4 223.167
R132 plus.n24 plus.t8 223.167
R133 plus.n23 plus.t6 223.167
R134 plus.n17 plus.t0 223.167
R135 plus.n18 plus.t5 223.167
R136 plus.n6 plus.n3 161.3
R137 plus.n8 plus.n7 161.3
R138 plus.n9 plus.n2 161.3
R139 plus.n10 plus.n1 161.3
R140 plus.n11 plus.n0 161.3
R141 plus.n13 plus.n12 161.3
R142 plus.n20 plus.n17 161.3
R143 plus.n22 plus.n21 161.3
R144 plus.n23 plus.n16 161.3
R145 plus.n24 plus.n15 161.3
R146 plus.n25 plus.n14 161.3
R147 plus.n27 plus.n26 161.3
R148 plus.n10 plus.n9 48.2005
R149 plus.n4 plus.n3 48.2005
R150 plus.n24 plus.n23 48.2005
R151 plus.n18 plus.n17 48.2005
R152 plus.n12 plus.n11 47.4702
R153 plus.n26 plus.n25 47.4702
R154 plus.n6 plus.n5 45.1192
R155 plus.n20 plus.n19 45.1192
R156 plus plus.n27 26.7377
R157 plus.n8 plus.n3 24.1005
R158 plus.n9 plus.n8 24.1005
R159 plus.n23 plus.n22 24.1005
R160 plus.n22 plus.n17 24.1005
R161 plus.n5 plus.n4 13.6377
R162 plus.n19 plus.n18 13.6377
R163 plus plus.n13 8.76565
R164 plus.n11 plus.n10 0.730803
R165 plus.n25 plus.n24 0.730803
R166 plus.n7 plus.n6 0.189894
R167 plus.n7 plus.n2 0.189894
R168 plus.n2 plus.n1 0.189894
R169 plus.n1 plus.n0 0.189894
R170 plus.n13 plus.n0 0.189894
R171 plus.n27 plus.n14 0.189894
R172 plus.n15 plus.n14 0.189894
R173 plus.n16 plus.n15 0.189894
R174 plus.n21 plus.n16 0.189894
R175 plus.n21 plus.n20 0.189894
R176 drain_left.n6 drain_left.n4 80.4886
R177 drain_left.n3 drain_left.n2 80.4332
R178 drain_left.n3 drain_left.n0 80.4332
R179 drain_left.n8 drain_left.n7 79.7731
R180 drain_left.n6 drain_left.n5 79.7731
R181 drain_left.n3 drain_left.n1 79.773
R182 drain_left drain_left.n3 24.1265
R183 drain_left.n1 drain_left.t5 6.6005
R184 drain_left.n1 drain_left.t11 6.6005
R185 drain_left.n2 drain_left.t6 6.6005
R186 drain_left.n2 drain_left.t9 6.6005
R187 drain_left.n0 drain_left.t7 6.6005
R188 drain_left.n0 drain_left.t3 6.6005
R189 drain_left.n7 drain_left.t2 6.6005
R190 drain_left.n7 drain_left.t0 6.6005
R191 drain_left.n5 drain_left.t1 6.6005
R192 drain_left.n5 drain_left.t8 6.6005
R193 drain_left.n4 drain_left.t10 6.6005
R194 drain_left.n4 drain_left.t4 6.6005
R195 drain_left drain_left.n8 6.36873
R196 drain_left.n8 drain_left.n6 0.716017
C0 drain_right drain_left 0.936369f
C1 drain_right source 6.48676f
C2 minus drain_left 0.176612f
C3 minus source 2.18962f
C4 drain_right plus 0.342826f
C5 minus plus 3.83316f
C6 source drain_left 6.48579f
C7 drain_left plus 2.15152f
C8 source plus 2.20362f
C9 drain_right minus 1.96896f
C10 drain_right a_n1878_n1488# 3.81272f
C11 drain_left a_n1878_n1488# 4.49471f
C12 source a_n1878_n1488# 3.702974f
C13 minus a_n1878_n1488# 6.635406f
C14 plus a_n1878_n1488# 7.94384f
C15 drain_left.t7 a_n1878_n1488# 0.067408f
C16 drain_left.t3 a_n1878_n1488# 0.067408f
C17 drain_left.n0 a_n1878_n1488# 0.489147f
C18 drain_left.t5 a_n1878_n1488# 0.067408f
C19 drain_left.t11 a_n1878_n1488# 0.067408f
C20 drain_left.n1 a_n1878_n1488# 0.486142f
C21 drain_left.t6 a_n1878_n1488# 0.067408f
C22 drain_left.t9 a_n1878_n1488# 0.067408f
C23 drain_left.n2 a_n1878_n1488# 0.489147f
C24 drain_left.n3 a_n1878_n1488# 1.90494f
C25 drain_left.t10 a_n1878_n1488# 0.067408f
C26 drain_left.t4 a_n1878_n1488# 0.067408f
C27 drain_left.n4 a_n1878_n1488# 0.489435f
C28 drain_left.t1 a_n1878_n1488# 0.067408f
C29 drain_left.t8 a_n1878_n1488# 0.067408f
C30 drain_left.n5 a_n1878_n1488# 0.486144f
C31 drain_left.n6 a_n1878_n1488# 0.725602f
C32 drain_left.t2 a_n1878_n1488# 0.067408f
C33 drain_left.t0 a_n1878_n1488# 0.067408f
C34 drain_left.n7 a_n1878_n1488# 0.486144f
C35 drain_left.n8 a_n1878_n1488# 0.603008f
C36 plus.n0 a_n1878_n1488# 0.049432f
C37 plus.t11 a_n1878_n1488# 0.222345f
C38 plus.t9 a_n1878_n1488# 0.222345f
C39 plus.n1 a_n1878_n1488# 0.049432f
C40 plus.t3 a_n1878_n1488# 0.222345f
C41 plus.n2 a_n1878_n1488# 0.049432f
C42 plus.t10 a_n1878_n1488# 0.222345f
C43 plus.n3 a_n1878_n1488# 0.138385f
C44 plus.t7 a_n1878_n1488# 0.222345f
C45 plus.n4 a_n1878_n1488# 0.144344f
C46 plus.t1 a_n1878_n1488# 0.236586f
C47 plus.n5 a_n1878_n1488# 0.120327f
C48 plus.n6 a_n1878_n1488# 0.20132f
C49 plus.n7 a_n1878_n1488# 0.049432f
C50 plus.n8 a_n1878_n1488# 0.011217f
C51 plus.n9 a_n1878_n1488# 0.138385f
C52 plus.n10 a_n1878_n1488# 0.133509f
C53 plus.n11 a_n1878_n1488# 0.011217f
C54 plus.n12 a_n1878_n1488# 0.133204f
C55 plus.n13 a_n1878_n1488# 0.373025f
C56 plus.n14 a_n1878_n1488# 0.049432f
C57 plus.t4 a_n1878_n1488# 0.222345f
C58 plus.n15 a_n1878_n1488# 0.049432f
C59 plus.t8 a_n1878_n1488# 0.222345f
C60 plus.n16 a_n1878_n1488# 0.049432f
C61 plus.t6 a_n1878_n1488# 0.222345f
C62 plus.t0 a_n1878_n1488# 0.222345f
C63 plus.n17 a_n1878_n1488# 0.138385f
C64 plus.t2 a_n1878_n1488# 0.236586f
C65 plus.t5 a_n1878_n1488# 0.222345f
C66 plus.n18 a_n1878_n1488# 0.144344f
C67 plus.n19 a_n1878_n1488# 0.120327f
C68 plus.n20 a_n1878_n1488# 0.20132f
C69 plus.n21 a_n1878_n1488# 0.049432f
C70 plus.n22 a_n1878_n1488# 0.011217f
C71 plus.n23 a_n1878_n1488# 0.138385f
C72 plus.n24 a_n1878_n1488# 0.133509f
C73 plus.n25 a_n1878_n1488# 0.011217f
C74 plus.n26 a_n1878_n1488# 0.133204f
C75 plus.n27 a_n1878_n1488# 1.17293f
C76 source.t4 a_n1878_n1488# 0.538927f
C77 source.n0 a_n1878_n1488# 0.762028f
C78 source.t1 a_n1878_n1488# 0.064901f
C79 source.t23 a_n1878_n1488# 0.064901f
C80 source.n1 a_n1878_n1488# 0.41151f
C81 source.n2 a_n1878_n1488# 0.36472f
C82 source.t8 a_n1878_n1488# 0.064901f
C83 source.t5 a_n1878_n1488# 0.064901f
C84 source.n3 a_n1878_n1488# 0.41151f
C85 source.n4 a_n1878_n1488# 0.36472f
C86 source.t2 a_n1878_n1488# 0.538927f
C87 source.n5 a_n1878_n1488# 0.392633f
C88 source.t11 a_n1878_n1488# 0.538927f
C89 source.n6 a_n1878_n1488# 0.392633f
C90 source.t15 a_n1878_n1488# 0.064901f
C91 source.t19 a_n1878_n1488# 0.064901f
C92 source.n7 a_n1878_n1488# 0.41151f
C93 source.n8 a_n1878_n1488# 0.36472f
C94 source.t17 a_n1878_n1488# 0.064901f
C95 source.t9 a_n1878_n1488# 0.064901f
C96 source.n9 a_n1878_n1488# 0.41151f
C97 source.n10 a_n1878_n1488# 0.36472f
C98 source.t12 a_n1878_n1488# 0.538927f
C99 source.n11 a_n1878_n1488# 1.05106f
C100 source.t6 a_n1878_n1488# 0.538925f
C101 source.n12 a_n1878_n1488# 1.05106f
C102 source.t0 a_n1878_n1488# 0.064901f
C103 source.t21 a_n1878_n1488# 0.064901f
C104 source.n13 a_n1878_n1488# 0.411507f
C105 source.n14 a_n1878_n1488# 0.364723f
C106 source.t3 a_n1878_n1488# 0.064901f
C107 source.t22 a_n1878_n1488# 0.064901f
C108 source.n15 a_n1878_n1488# 0.411507f
C109 source.n16 a_n1878_n1488# 0.364723f
C110 source.t7 a_n1878_n1488# 0.538925f
C111 source.n17 a_n1878_n1488# 0.392636f
C112 source.t18 a_n1878_n1488# 0.538925f
C113 source.n18 a_n1878_n1488# 0.392636f
C114 source.t14 a_n1878_n1488# 0.064901f
C115 source.t20 a_n1878_n1488# 0.064901f
C116 source.n19 a_n1878_n1488# 0.411507f
C117 source.n20 a_n1878_n1488# 0.364723f
C118 source.t16 a_n1878_n1488# 0.064901f
C119 source.t10 a_n1878_n1488# 0.064901f
C120 source.n21 a_n1878_n1488# 0.411507f
C121 source.n22 a_n1878_n1488# 0.364723f
C122 source.t13 a_n1878_n1488# 0.538925f
C123 source.n23 a_n1878_n1488# 0.559262f
C124 source.n24 a_n1878_n1488# 0.800301f
C125 drain_right.t2 a_n1878_n1488# 0.051015f
C126 drain_right.t8 a_n1878_n1488# 0.051015f
C127 drain_right.n0 a_n1878_n1488# 0.370187f
C128 drain_right.t1 a_n1878_n1488# 0.051015f
C129 drain_right.t9 a_n1878_n1488# 0.051015f
C130 drain_right.n1 a_n1878_n1488# 0.367913f
C131 drain_right.t11 a_n1878_n1488# 0.051015f
C132 drain_right.t3 a_n1878_n1488# 0.051015f
C133 drain_right.n2 a_n1878_n1488# 0.370187f
C134 drain_right.n3 a_n1878_n1488# 1.39904f
C135 drain_right.t6 a_n1878_n1488# 0.051015f
C136 drain_right.t4 a_n1878_n1488# 0.051015f
C137 drain_right.n4 a_n1878_n1488# 0.370405f
C138 drain_right.t10 a_n1878_n1488# 0.051015f
C139 drain_right.t7 a_n1878_n1488# 0.051015f
C140 drain_right.n5 a_n1878_n1488# 0.367915f
C141 drain_right.n6 a_n1878_n1488# 0.549137f
C142 drain_right.t0 a_n1878_n1488# 0.051015f
C143 drain_right.t5 a_n1878_n1488# 0.051015f
C144 drain_right.n7 a_n1878_n1488# 0.367915f
C145 drain_right.n8 a_n1878_n1488# 0.456358f
C146 minus.n0 a_n1878_n1488# 0.035734f
C147 minus.t11 a_n1878_n1488# 0.160732f
C148 minus.n1 a_n1878_n1488# 0.100038f
C149 minus.t3 a_n1878_n1488# 0.160732f
C150 minus.n2 a_n1878_n1488# 0.145533f
C151 minus.t9 a_n1878_n1488# 0.171027f
C152 minus.n3 a_n1878_n1488# 0.086984f
C153 minus.t1 a_n1878_n1488# 0.160732f
C154 minus.n4 a_n1878_n1488# 0.104345f
C155 minus.t5 a_n1878_n1488# 0.160732f
C156 minus.n5 a_n1878_n1488# 0.100038f
C157 minus.n6 a_n1878_n1488# 0.008109f
C158 minus.n7 a_n1878_n1488# 0.035734f
C159 minus.n8 a_n1878_n1488# 0.035734f
C160 minus.n9 a_n1878_n1488# 0.035734f
C161 minus.n10 a_n1878_n1488# 0.096513f
C162 minus.n11 a_n1878_n1488# 0.008109f
C163 minus.t8 a_n1878_n1488# 0.160732f
C164 minus.n12 a_n1878_n1488# 0.096293f
C165 minus.n13 a_n1878_n1488# 0.901464f
C166 minus.n14 a_n1878_n1488# 0.035734f
C167 minus.t4 a_n1878_n1488# 0.160732f
C168 minus.n15 a_n1878_n1488# 0.100038f
C169 minus.n16 a_n1878_n1488# 0.145533f
C170 minus.t2 a_n1878_n1488# 0.171027f
C171 minus.n17 a_n1878_n1488# 0.086984f
C172 minus.t6 a_n1878_n1488# 0.160732f
C173 minus.n18 a_n1878_n1488# 0.104345f
C174 minus.t0 a_n1878_n1488# 0.160732f
C175 minus.n19 a_n1878_n1488# 0.100038f
C176 minus.n20 a_n1878_n1488# 0.008109f
C177 minus.n21 a_n1878_n1488# 0.035734f
C178 minus.n22 a_n1878_n1488# 0.035734f
C179 minus.n23 a_n1878_n1488# 0.035734f
C180 minus.t10 a_n1878_n1488# 0.160732f
C181 minus.n24 a_n1878_n1488# 0.096513f
C182 minus.n25 a_n1878_n1488# 0.008109f
C183 minus.t7 a_n1878_n1488# 0.160732f
C184 minus.n26 a_n1878_n1488# 0.096293f
C185 minus.n27 a_n1878_n1488# 0.236212f
C186 minus.n28 a_n1878_n1488# 1.11169f
.ends

