* NGSPICE file created from diffpair436.ext - technology: sky130A

.subckt diffpair436 minus drain_right drain_left source plus
X0 a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.3
X1 drain_right.t13 minus.t0 source.t15 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X2 drain_right.t12 minus.t1 source.t21 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X3 source.t22 minus.t2 drain_right.t11 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X4 drain_right.t10 minus.t3 source.t17 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X5 drain_left.t13 plus.t0 source.t2 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X6 drain_left.t12 plus.t1 source.t6 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X7 drain_left.t11 plus.t2 source.t8 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X8 drain_right.t9 minus.t4 source.t26 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X9 drain_right.t8 minus.t5 source.t25 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X10 drain_right.t7 minus.t6 source.t23 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X11 a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X12 drain_left.t10 plus.t3 source.t1 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X13 source.t0 plus.t4 drain_left.t9 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X14 source.t11 plus.t5 drain_left.t8 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X15 source.t20 minus.t7 drain_right.t6 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X16 source.t7 plus.t6 drain_left.t7 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X17 source.t10 plus.t7 drain_left.t6 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X18 drain_right.t5 minus.t8 source.t19 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X19 source.t4 plus.t8 drain_left.t5 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X20 source.t18 minus.t9 drain_right.t4 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X21 source.t27 minus.t10 drain_right.t3 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X22 a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X23 drain_left.t4 plus.t9 source.t12 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X24 source.t24 minus.t11 drain_right.t2 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X25 drain_right.t1 minus.t12 source.t16 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X26 drain_left.t3 plus.t10 source.t13 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X27 drain_left.t2 plus.t11 source.t3 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X28 a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X29 source.t14 minus.t13 drain_right.t0 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X30 drain_left.t1 plus.t12 source.t9 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X31 source.t5 plus.t13 drain_left.t0 a_n1724_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
R0 minus.n15 minus.t4 1125.4
R1 minus.n3 minus.t8 1125.4
R2 minus.n32 minus.t5 1125.4
R3 minus.n20 minus.t1 1125.4
R4 minus.n1 minus.t7 1068.43
R5 minus.n14 minus.t2 1068.43
R6 minus.n12 minus.t12 1068.43
R7 minus.n6 minus.t3 1068.43
R8 minus.n4 minus.t13 1068.43
R9 minus.n18 minus.t9 1068.43
R10 minus.n31 minus.t11 1068.43
R11 minus.n29 minus.t6 1068.43
R12 minus.n23 minus.t0 1068.43
R13 minus.n21 minus.t10 1068.43
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n34 minus.n16 35.688
R41 minus.n15 minus.n14 35.055
R42 minus.n4 minus.n3 35.055
R43 minus.n21 minus.n20 35.055
R44 minus.n32 minus.n31 35.055
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 source.n282 source.n222 289.615
R62 source.n210 source.n150 289.615
R63 source.n60 source.n0 289.615
R64 source.n132 source.n72 289.615
R65 source.n242 source.n241 185
R66 source.n247 source.n246 185
R67 source.n249 source.n248 185
R68 source.n238 source.n237 185
R69 source.n255 source.n254 185
R70 source.n257 source.n256 185
R71 source.n234 source.n233 185
R72 source.n264 source.n263 185
R73 source.n265 source.n232 185
R74 source.n267 source.n266 185
R75 source.n230 source.n229 185
R76 source.n273 source.n272 185
R77 source.n275 source.n274 185
R78 source.n226 source.n225 185
R79 source.n281 source.n280 185
R80 source.n283 source.n282 185
R81 source.n170 source.n169 185
R82 source.n175 source.n174 185
R83 source.n177 source.n176 185
R84 source.n166 source.n165 185
R85 source.n183 source.n182 185
R86 source.n185 source.n184 185
R87 source.n162 source.n161 185
R88 source.n192 source.n191 185
R89 source.n193 source.n160 185
R90 source.n195 source.n194 185
R91 source.n158 source.n157 185
R92 source.n201 source.n200 185
R93 source.n203 source.n202 185
R94 source.n154 source.n153 185
R95 source.n209 source.n208 185
R96 source.n211 source.n210 185
R97 source.n61 source.n60 185
R98 source.n59 source.n58 185
R99 source.n4 source.n3 185
R100 source.n53 source.n52 185
R101 source.n51 source.n50 185
R102 source.n8 source.n7 185
R103 source.n45 source.n44 185
R104 source.n43 source.n10 185
R105 source.n42 source.n41 185
R106 source.n13 source.n11 185
R107 source.n36 source.n35 185
R108 source.n34 source.n33 185
R109 source.n17 source.n16 185
R110 source.n28 source.n27 185
R111 source.n26 source.n25 185
R112 source.n21 source.n20 185
R113 source.n133 source.n132 185
R114 source.n131 source.n130 185
R115 source.n76 source.n75 185
R116 source.n125 source.n124 185
R117 source.n123 source.n122 185
R118 source.n80 source.n79 185
R119 source.n117 source.n116 185
R120 source.n115 source.n82 185
R121 source.n114 source.n113 185
R122 source.n85 source.n83 185
R123 source.n108 source.n107 185
R124 source.n106 source.n105 185
R125 source.n89 source.n88 185
R126 source.n100 source.n99 185
R127 source.n98 source.n97 185
R128 source.n93 source.n92 185
R129 source.n243 source.t25 149.524
R130 source.n171 source.t13 149.524
R131 source.n22 source.t9 149.524
R132 source.n94 source.t19 149.524
R133 source.n247 source.n241 104.615
R134 source.n248 source.n247 104.615
R135 source.n248 source.n237 104.615
R136 source.n255 source.n237 104.615
R137 source.n256 source.n255 104.615
R138 source.n256 source.n233 104.615
R139 source.n264 source.n233 104.615
R140 source.n265 source.n264 104.615
R141 source.n266 source.n265 104.615
R142 source.n266 source.n229 104.615
R143 source.n273 source.n229 104.615
R144 source.n274 source.n273 104.615
R145 source.n274 source.n225 104.615
R146 source.n281 source.n225 104.615
R147 source.n282 source.n281 104.615
R148 source.n175 source.n169 104.615
R149 source.n176 source.n175 104.615
R150 source.n176 source.n165 104.615
R151 source.n183 source.n165 104.615
R152 source.n184 source.n183 104.615
R153 source.n184 source.n161 104.615
R154 source.n192 source.n161 104.615
R155 source.n193 source.n192 104.615
R156 source.n194 source.n193 104.615
R157 source.n194 source.n157 104.615
R158 source.n201 source.n157 104.615
R159 source.n202 source.n201 104.615
R160 source.n202 source.n153 104.615
R161 source.n209 source.n153 104.615
R162 source.n210 source.n209 104.615
R163 source.n60 source.n59 104.615
R164 source.n59 source.n3 104.615
R165 source.n52 source.n3 104.615
R166 source.n52 source.n51 104.615
R167 source.n51 source.n7 104.615
R168 source.n44 source.n7 104.615
R169 source.n44 source.n43 104.615
R170 source.n43 source.n42 104.615
R171 source.n42 source.n11 104.615
R172 source.n35 source.n11 104.615
R173 source.n35 source.n34 104.615
R174 source.n34 source.n16 104.615
R175 source.n27 source.n16 104.615
R176 source.n27 source.n26 104.615
R177 source.n26 source.n20 104.615
R178 source.n132 source.n131 104.615
R179 source.n131 source.n75 104.615
R180 source.n124 source.n75 104.615
R181 source.n124 source.n123 104.615
R182 source.n123 source.n79 104.615
R183 source.n116 source.n79 104.615
R184 source.n116 source.n115 104.615
R185 source.n115 source.n114 104.615
R186 source.n114 source.n83 104.615
R187 source.n107 source.n83 104.615
R188 source.n107 source.n106 104.615
R189 source.n106 source.n88 104.615
R190 source.n99 source.n88 104.615
R191 source.n99 source.n98 104.615
R192 source.n98 source.n92 104.615
R193 source.t25 source.n241 52.3082
R194 source.t13 source.n169 52.3082
R195 source.t9 source.n20 52.3082
R196 source.t19 source.n92 52.3082
R197 source.n67 source.n66 42.8739
R198 source.n69 source.n68 42.8739
R199 source.n71 source.n70 42.8739
R200 source.n139 source.n138 42.8739
R201 source.n141 source.n140 42.8739
R202 source.n143 source.n142 42.8739
R203 source.n221 source.n220 42.8737
R204 source.n219 source.n218 42.8737
R205 source.n217 source.n216 42.8737
R206 source.n149 source.n148 42.8737
R207 source.n147 source.n146 42.8737
R208 source.n145 source.n144 42.8737
R209 source.n287 source.n286 29.8581
R210 source.n215 source.n214 29.8581
R211 source.n65 source.n64 29.8581
R212 source.n137 source.n136 29.8581
R213 source.n145 source.n143 22.3739
R214 source.n288 source.n65 16.2963
R215 source.n267 source.n232 13.1884
R216 source.n195 source.n160 13.1884
R217 source.n45 source.n10 13.1884
R218 source.n117 source.n82 13.1884
R219 source.n263 source.n262 12.8005
R220 source.n268 source.n230 12.8005
R221 source.n191 source.n190 12.8005
R222 source.n196 source.n158 12.8005
R223 source.n46 source.n8 12.8005
R224 source.n41 source.n12 12.8005
R225 source.n118 source.n80 12.8005
R226 source.n113 source.n84 12.8005
R227 source.n261 source.n234 12.0247
R228 source.n272 source.n271 12.0247
R229 source.n189 source.n162 12.0247
R230 source.n200 source.n199 12.0247
R231 source.n50 source.n49 12.0247
R232 source.n40 source.n13 12.0247
R233 source.n122 source.n121 12.0247
R234 source.n112 source.n85 12.0247
R235 source.n258 source.n257 11.249
R236 source.n275 source.n228 11.249
R237 source.n186 source.n185 11.249
R238 source.n203 source.n156 11.249
R239 source.n53 source.n6 11.249
R240 source.n37 source.n36 11.249
R241 source.n125 source.n78 11.249
R242 source.n109 source.n108 11.249
R243 source.n254 source.n236 10.4732
R244 source.n276 source.n226 10.4732
R245 source.n182 source.n164 10.4732
R246 source.n204 source.n154 10.4732
R247 source.n54 source.n4 10.4732
R248 source.n33 source.n15 10.4732
R249 source.n126 source.n76 10.4732
R250 source.n105 source.n87 10.4732
R251 source.n243 source.n242 10.2747
R252 source.n171 source.n170 10.2747
R253 source.n22 source.n21 10.2747
R254 source.n94 source.n93 10.2747
R255 source.n253 source.n238 9.69747
R256 source.n280 source.n279 9.69747
R257 source.n181 source.n166 9.69747
R258 source.n208 source.n207 9.69747
R259 source.n58 source.n57 9.69747
R260 source.n32 source.n17 9.69747
R261 source.n130 source.n129 9.69747
R262 source.n104 source.n89 9.69747
R263 source.n286 source.n285 9.45567
R264 source.n214 source.n213 9.45567
R265 source.n64 source.n63 9.45567
R266 source.n136 source.n135 9.45567
R267 source.n285 source.n284 9.3005
R268 source.n224 source.n223 9.3005
R269 source.n279 source.n278 9.3005
R270 source.n277 source.n276 9.3005
R271 source.n228 source.n227 9.3005
R272 source.n271 source.n270 9.3005
R273 source.n269 source.n268 9.3005
R274 source.n245 source.n244 9.3005
R275 source.n240 source.n239 9.3005
R276 source.n251 source.n250 9.3005
R277 source.n253 source.n252 9.3005
R278 source.n236 source.n235 9.3005
R279 source.n259 source.n258 9.3005
R280 source.n261 source.n260 9.3005
R281 source.n262 source.n231 9.3005
R282 source.n213 source.n212 9.3005
R283 source.n152 source.n151 9.3005
R284 source.n207 source.n206 9.3005
R285 source.n205 source.n204 9.3005
R286 source.n156 source.n155 9.3005
R287 source.n199 source.n198 9.3005
R288 source.n197 source.n196 9.3005
R289 source.n173 source.n172 9.3005
R290 source.n168 source.n167 9.3005
R291 source.n179 source.n178 9.3005
R292 source.n181 source.n180 9.3005
R293 source.n164 source.n163 9.3005
R294 source.n187 source.n186 9.3005
R295 source.n189 source.n188 9.3005
R296 source.n190 source.n159 9.3005
R297 source.n24 source.n23 9.3005
R298 source.n19 source.n18 9.3005
R299 source.n30 source.n29 9.3005
R300 source.n32 source.n31 9.3005
R301 source.n15 source.n14 9.3005
R302 source.n38 source.n37 9.3005
R303 source.n40 source.n39 9.3005
R304 source.n12 source.n9 9.3005
R305 source.n63 source.n62 9.3005
R306 source.n2 source.n1 9.3005
R307 source.n57 source.n56 9.3005
R308 source.n55 source.n54 9.3005
R309 source.n6 source.n5 9.3005
R310 source.n49 source.n48 9.3005
R311 source.n47 source.n46 9.3005
R312 source.n96 source.n95 9.3005
R313 source.n91 source.n90 9.3005
R314 source.n102 source.n101 9.3005
R315 source.n104 source.n103 9.3005
R316 source.n87 source.n86 9.3005
R317 source.n110 source.n109 9.3005
R318 source.n112 source.n111 9.3005
R319 source.n84 source.n81 9.3005
R320 source.n135 source.n134 9.3005
R321 source.n74 source.n73 9.3005
R322 source.n129 source.n128 9.3005
R323 source.n127 source.n126 9.3005
R324 source.n78 source.n77 9.3005
R325 source.n121 source.n120 9.3005
R326 source.n119 source.n118 9.3005
R327 source.n250 source.n249 8.92171
R328 source.n283 source.n224 8.92171
R329 source.n178 source.n177 8.92171
R330 source.n211 source.n152 8.92171
R331 source.n61 source.n2 8.92171
R332 source.n29 source.n28 8.92171
R333 source.n133 source.n74 8.92171
R334 source.n101 source.n100 8.92171
R335 source.n246 source.n240 8.14595
R336 source.n284 source.n222 8.14595
R337 source.n174 source.n168 8.14595
R338 source.n212 source.n150 8.14595
R339 source.n62 source.n0 8.14595
R340 source.n25 source.n19 8.14595
R341 source.n134 source.n72 8.14595
R342 source.n97 source.n91 8.14595
R343 source.n245 source.n242 7.3702
R344 source.n173 source.n170 7.3702
R345 source.n24 source.n21 7.3702
R346 source.n96 source.n93 7.3702
R347 source.n246 source.n245 5.81868
R348 source.n286 source.n222 5.81868
R349 source.n174 source.n173 5.81868
R350 source.n214 source.n150 5.81868
R351 source.n64 source.n0 5.81868
R352 source.n25 source.n24 5.81868
R353 source.n136 source.n72 5.81868
R354 source.n97 source.n96 5.81868
R355 source.n288 source.n287 5.53498
R356 source.n249 source.n240 5.04292
R357 source.n284 source.n283 5.04292
R358 source.n177 source.n168 5.04292
R359 source.n212 source.n211 5.04292
R360 source.n62 source.n61 5.04292
R361 source.n28 source.n19 5.04292
R362 source.n134 source.n133 5.04292
R363 source.n100 source.n91 5.04292
R364 source.n250 source.n238 4.26717
R365 source.n280 source.n224 4.26717
R366 source.n178 source.n166 4.26717
R367 source.n208 source.n152 4.26717
R368 source.n58 source.n2 4.26717
R369 source.n29 source.n17 4.26717
R370 source.n130 source.n74 4.26717
R371 source.n101 source.n89 4.26717
R372 source.n254 source.n253 3.49141
R373 source.n279 source.n226 3.49141
R374 source.n182 source.n181 3.49141
R375 source.n207 source.n154 3.49141
R376 source.n57 source.n4 3.49141
R377 source.n33 source.n32 3.49141
R378 source.n129 source.n76 3.49141
R379 source.n105 source.n104 3.49141
R380 source.n244 source.n243 2.84303
R381 source.n172 source.n171 2.84303
R382 source.n23 source.n22 2.84303
R383 source.n95 source.n94 2.84303
R384 source.n257 source.n236 2.71565
R385 source.n276 source.n275 2.71565
R386 source.n185 source.n164 2.71565
R387 source.n204 source.n203 2.71565
R388 source.n54 source.n53 2.71565
R389 source.n36 source.n15 2.71565
R390 source.n126 source.n125 2.71565
R391 source.n108 source.n87 2.71565
R392 source.n258 source.n234 1.93989
R393 source.n272 source.n228 1.93989
R394 source.n186 source.n162 1.93989
R395 source.n200 source.n156 1.93989
R396 source.n50 source.n6 1.93989
R397 source.n37 source.n13 1.93989
R398 source.n122 source.n78 1.93989
R399 source.n109 source.n85 1.93989
R400 source.n220 source.t23 1.6505
R401 source.n220 source.t24 1.6505
R402 source.n218 source.t15 1.6505
R403 source.n218 source.t18 1.6505
R404 source.n216 source.t21 1.6505
R405 source.n216 source.t27 1.6505
R406 source.n148 source.t3 1.6505
R407 source.n148 source.t0 1.6505
R408 source.n146 source.t2 1.6505
R409 source.n146 source.t7 1.6505
R410 source.n144 source.t8 1.6505
R411 source.n144 source.t10 1.6505
R412 source.n66 source.t1 1.6505
R413 source.n66 source.t4 1.6505
R414 source.n68 source.t12 1.6505
R415 source.n68 source.t5 1.6505
R416 source.n70 source.t6 1.6505
R417 source.n70 source.t11 1.6505
R418 source.n138 source.t17 1.6505
R419 source.n138 source.t14 1.6505
R420 source.n140 source.t16 1.6505
R421 source.n140 source.t20 1.6505
R422 source.n142 source.t26 1.6505
R423 source.n142 source.t22 1.6505
R424 source.n263 source.n261 1.16414
R425 source.n271 source.n230 1.16414
R426 source.n191 source.n189 1.16414
R427 source.n199 source.n158 1.16414
R428 source.n49 source.n8 1.16414
R429 source.n41 source.n40 1.16414
R430 source.n121 source.n80 1.16414
R431 source.n113 source.n112 1.16414
R432 source.n137 source.n71 0.741879
R433 source.n217 source.n215 0.741879
R434 source.n143 source.n141 0.543603
R435 source.n141 source.n139 0.543603
R436 source.n139 source.n137 0.543603
R437 source.n71 source.n69 0.543603
R438 source.n69 source.n67 0.543603
R439 source.n67 source.n65 0.543603
R440 source.n147 source.n145 0.543603
R441 source.n149 source.n147 0.543603
R442 source.n215 source.n149 0.543603
R443 source.n219 source.n217 0.543603
R444 source.n221 source.n219 0.543603
R445 source.n287 source.n221 0.543603
R446 source.n262 source.n232 0.388379
R447 source.n268 source.n267 0.388379
R448 source.n190 source.n160 0.388379
R449 source.n196 source.n195 0.388379
R450 source.n46 source.n45 0.388379
R451 source.n12 source.n10 0.388379
R452 source.n118 source.n117 0.388379
R453 source.n84 source.n82 0.388379
R454 source source.n288 0.188
R455 source.n244 source.n239 0.155672
R456 source.n251 source.n239 0.155672
R457 source.n252 source.n251 0.155672
R458 source.n252 source.n235 0.155672
R459 source.n259 source.n235 0.155672
R460 source.n260 source.n259 0.155672
R461 source.n260 source.n231 0.155672
R462 source.n269 source.n231 0.155672
R463 source.n270 source.n269 0.155672
R464 source.n270 source.n227 0.155672
R465 source.n277 source.n227 0.155672
R466 source.n278 source.n277 0.155672
R467 source.n278 source.n223 0.155672
R468 source.n285 source.n223 0.155672
R469 source.n172 source.n167 0.155672
R470 source.n179 source.n167 0.155672
R471 source.n180 source.n179 0.155672
R472 source.n180 source.n163 0.155672
R473 source.n187 source.n163 0.155672
R474 source.n188 source.n187 0.155672
R475 source.n188 source.n159 0.155672
R476 source.n197 source.n159 0.155672
R477 source.n198 source.n197 0.155672
R478 source.n198 source.n155 0.155672
R479 source.n205 source.n155 0.155672
R480 source.n206 source.n205 0.155672
R481 source.n206 source.n151 0.155672
R482 source.n213 source.n151 0.155672
R483 source.n63 source.n1 0.155672
R484 source.n56 source.n1 0.155672
R485 source.n56 source.n55 0.155672
R486 source.n55 source.n5 0.155672
R487 source.n48 source.n5 0.155672
R488 source.n48 source.n47 0.155672
R489 source.n47 source.n9 0.155672
R490 source.n39 source.n9 0.155672
R491 source.n39 source.n38 0.155672
R492 source.n38 source.n14 0.155672
R493 source.n31 source.n14 0.155672
R494 source.n31 source.n30 0.155672
R495 source.n30 source.n18 0.155672
R496 source.n23 source.n18 0.155672
R497 source.n135 source.n73 0.155672
R498 source.n128 source.n73 0.155672
R499 source.n128 source.n127 0.155672
R500 source.n127 source.n77 0.155672
R501 source.n120 source.n77 0.155672
R502 source.n120 source.n119 0.155672
R503 source.n119 source.n81 0.155672
R504 source.n111 source.n81 0.155672
R505 source.n111 source.n110 0.155672
R506 source.n110 source.n86 0.155672
R507 source.n103 source.n86 0.155672
R508 source.n103 source.n102 0.155672
R509 source.n102 source.n90 0.155672
R510 source.n95 source.n90 0.155672
R511 drain_right.n60 drain_right.n0 289.615
R512 drain_right.n136 drain_right.n76 289.615
R513 drain_right.n20 drain_right.n19 185
R514 drain_right.n25 drain_right.n24 185
R515 drain_right.n27 drain_right.n26 185
R516 drain_right.n16 drain_right.n15 185
R517 drain_right.n33 drain_right.n32 185
R518 drain_right.n35 drain_right.n34 185
R519 drain_right.n12 drain_right.n11 185
R520 drain_right.n42 drain_right.n41 185
R521 drain_right.n43 drain_right.n10 185
R522 drain_right.n45 drain_right.n44 185
R523 drain_right.n8 drain_right.n7 185
R524 drain_right.n51 drain_right.n50 185
R525 drain_right.n53 drain_right.n52 185
R526 drain_right.n4 drain_right.n3 185
R527 drain_right.n59 drain_right.n58 185
R528 drain_right.n61 drain_right.n60 185
R529 drain_right.n137 drain_right.n136 185
R530 drain_right.n135 drain_right.n134 185
R531 drain_right.n80 drain_right.n79 185
R532 drain_right.n129 drain_right.n128 185
R533 drain_right.n127 drain_right.n126 185
R534 drain_right.n84 drain_right.n83 185
R535 drain_right.n121 drain_right.n120 185
R536 drain_right.n119 drain_right.n86 185
R537 drain_right.n118 drain_right.n117 185
R538 drain_right.n89 drain_right.n87 185
R539 drain_right.n112 drain_right.n111 185
R540 drain_right.n110 drain_right.n109 185
R541 drain_right.n93 drain_right.n92 185
R542 drain_right.n104 drain_right.n103 185
R543 drain_right.n102 drain_right.n101 185
R544 drain_right.n97 drain_right.n96 185
R545 drain_right.n21 drain_right.t12 149.524
R546 drain_right.n98 drain_right.t9 149.524
R547 drain_right.n25 drain_right.n19 104.615
R548 drain_right.n26 drain_right.n25 104.615
R549 drain_right.n26 drain_right.n15 104.615
R550 drain_right.n33 drain_right.n15 104.615
R551 drain_right.n34 drain_right.n33 104.615
R552 drain_right.n34 drain_right.n11 104.615
R553 drain_right.n42 drain_right.n11 104.615
R554 drain_right.n43 drain_right.n42 104.615
R555 drain_right.n44 drain_right.n43 104.615
R556 drain_right.n44 drain_right.n7 104.615
R557 drain_right.n51 drain_right.n7 104.615
R558 drain_right.n52 drain_right.n51 104.615
R559 drain_right.n52 drain_right.n3 104.615
R560 drain_right.n59 drain_right.n3 104.615
R561 drain_right.n60 drain_right.n59 104.615
R562 drain_right.n136 drain_right.n135 104.615
R563 drain_right.n135 drain_right.n79 104.615
R564 drain_right.n128 drain_right.n79 104.615
R565 drain_right.n128 drain_right.n127 104.615
R566 drain_right.n127 drain_right.n83 104.615
R567 drain_right.n120 drain_right.n83 104.615
R568 drain_right.n120 drain_right.n119 104.615
R569 drain_right.n119 drain_right.n118 104.615
R570 drain_right.n118 drain_right.n87 104.615
R571 drain_right.n111 drain_right.n87 104.615
R572 drain_right.n111 drain_right.n110 104.615
R573 drain_right.n110 drain_right.n92 104.615
R574 drain_right.n103 drain_right.n92 104.615
R575 drain_right.n103 drain_right.n102 104.615
R576 drain_right.n102 drain_right.n96 104.615
R577 drain_right.n69 drain_right.n67 60.0956
R578 drain_right.n73 drain_right.n71 60.0956
R579 drain_right.n73 drain_right.n72 59.5527
R580 drain_right.n75 drain_right.n74 59.5527
R581 drain_right.n69 drain_right.n68 59.5525
R582 drain_right.n66 drain_right.n65 59.5525
R583 drain_right.t12 drain_right.n19 52.3082
R584 drain_right.t9 drain_right.n96 52.3082
R585 drain_right.n66 drain_right.n64 47.08
R586 drain_right.n141 drain_right.n140 46.5369
R587 drain_right drain_right.n70 29.9367
R588 drain_right.n45 drain_right.n10 13.1884
R589 drain_right.n121 drain_right.n86 13.1884
R590 drain_right.n41 drain_right.n40 12.8005
R591 drain_right.n46 drain_right.n8 12.8005
R592 drain_right.n122 drain_right.n84 12.8005
R593 drain_right.n117 drain_right.n88 12.8005
R594 drain_right.n39 drain_right.n12 12.0247
R595 drain_right.n50 drain_right.n49 12.0247
R596 drain_right.n126 drain_right.n125 12.0247
R597 drain_right.n116 drain_right.n89 12.0247
R598 drain_right.n36 drain_right.n35 11.249
R599 drain_right.n53 drain_right.n6 11.249
R600 drain_right.n129 drain_right.n82 11.249
R601 drain_right.n113 drain_right.n112 11.249
R602 drain_right.n32 drain_right.n14 10.4732
R603 drain_right.n54 drain_right.n4 10.4732
R604 drain_right.n130 drain_right.n80 10.4732
R605 drain_right.n109 drain_right.n91 10.4732
R606 drain_right.n21 drain_right.n20 10.2747
R607 drain_right.n98 drain_right.n97 10.2747
R608 drain_right.n31 drain_right.n16 9.69747
R609 drain_right.n58 drain_right.n57 9.69747
R610 drain_right.n134 drain_right.n133 9.69747
R611 drain_right.n108 drain_right.n93 9.69747
R612 drain_right.n64 drain_right.n63 9.45567
R613 drain_right.n140 drain_right.n139 9.45567
R614 drain_right.n63 drain_right.n62 9.3005
R615 drain_right.n2 drain_right.n1 9.3005
R616 drain_right.n57 drain_right.n56 9.3005
R617 drain_right.n55 drain_right.n54 9.3005
R618 drain_right.n6 drain_right.n5 9.3005
R619 drain_right.n49 drain_right.n48 9.3005
R620 drain_right.n47 drain_right.n46 9.3005
R621 drain_right.n23 drain_right.n22 9.3005
R622 drain_right.n18 drain_right.n17 9.3005
R623 drain_right.n29 drain_right.n28 9.3005
R624 drain_right.n31 drain_right.n30 9.3005
R625 drain_right.n14 drain_right.n13 9.3005
R626 drain_right.n37 drain_right.n36 9.3005
R627 drain_right.n39 drain_right.n38 9.3005
R628 drain_right.n40 drain_right.n9 9.3005
R629 drain_right.n100 drain_right.n99 9.3005
R630 drain_right.n95 drain_right.n94 9.3005
R631 drain_right.n106 drain_right.n105 9.3005
R632 drain_right.n108 drain_right.n107 9.3005
R633 drain_right.n91 drain_right.n90 9.3005
R634 drain_right.n114 drain_right.n113 9.3005
R635 drain_right.n116 drain_right.n115 9.3005
R636 drain_right.n88 drain_right.n85 9.3005
R637 drain_right.n139 drain_right.n138 9.3005
R638 drain_right.n78 drain_right.n77 9.3005
R639 drain_right.n133 drain_right.n132 9.3005
R640 drain_right.n131 drain_right.n130 9.3005
R641 drain_right.n82 drain_right.n81 9.3005
R642 drain_right.n125 drain_right.n124 9.3005
R643 drain_right.n123 drain_right.n122 9.3005
R644 drain_right.n28 drain_right.n27 8.92171
R645 drain_right.n61 drain_right.n2 8.92171
R646 drain_right.n137 drain_right.n78 8.92171
R647 drain_right.n105 drain_right.n104 8.92171
R648 drain_right.n24 drain_right.n18 8.14595
R649 drain_right.n62 drain_right.n0 8.14595
R650 drain_right.n138 drain_right.n76 8.14595
R651 drain_right.n101 drain_right.n95 8.14595
R652 drain_right.n23 drain_right.n20 7.3702
R653 drain_right.n100 drain_right.n97 7.3702
R654 drain_right drain_right.n141 5.92477
R655 drain_right.n24 drain_right.n23 5.81868
R656 drain_right.n64 drain_right.n0 5.81868
R657 drain_right.n140 drain_right.n76 5.81868
R658 drain_right.n101 drain_right.n100 5.81868
R659 drain_right.n27 drain_right.n18 5.04292
R660 drain_right.n62 drain_right.n61 5.04292
R661 drain_right.n138 drain_right.n137 5.04292
R662 drain_right.n104 drain_right.n95 5.04292
R663 drain_right.n28 drain_right.n16 4.26717
R664 drain_right.n58 drain_right.n2 4.26717
R665 drain_right.n134 drain_right.n78 4.26717
R666 drain_right.n105 drain_right.n93 4.26717
R667 drain_right.n32 drain_right.n31 3.49141
R668 drain_right.n57 drain_right.n4 3.49141
R669 drain_right.n133 drain_right.n80 3.49141
R670 drain_right.n109 drain_right.n108 3.49141
R671 drain_right.n22 drain_right.n21 2.84303
R672 drain_right.n99 drain_right.n98 2.84303
R673 drain_right.n35 drain_right.n14 2.71565
R674 drain_right.n54 drain_right.n53 2.71565
R675 drain_right.n130 drain_right.n129 2.71565
R676 drain_right.n112 drain_right.n91 2.71565
R677 drain_right.n36 drain_right.n12 1.93989
R678 drain_right.n50 drain_right.n6 1.93989
R679 drain_right.n126 drain_right.n82 1.93989
R680 drain_right.n113 drain_right.n89 1.93989
R681 drain_right.n67 drain_right.t2 1.6505
R682 drain_right.n67 drain_right.t8 1.6505
R683 drain_right.n68 drain_right.t4 1.6505
R684 drain_right.n68 drain_right.t7 1.6505
R685 drain_right.n65 drain_right.t3 1.6505
R686 drain_right.n65 drain_right.t13 1.6505
R687 drain_right.n71 drain_right.t0 1.6505
R688 drain_right.n71 drain_right.t5 1.6505
R689 drain_right.n72 drain_right.t6 1.6505
R690 drain_right.n72 drain_right.t10 1.6505
R691 drain_right.n74 drain_right.t11 1.6505
R692 drain_right.n74 drain_right.t1 1.6505
R693 drain_right.n41 drain_right.n39 1.16414
R694 drain_right.n49 drain_right.n8 1.16414
R695 drain_right.n125 drain_right.n84 1.16414
R696 drain_right.n117 drain_right.n116 1.16414
R697 drain_right.n141 drain_right.n75 0.543603
R698 drain_right.n75 drain_right.n73 0.543603
R699 drain_right.n40 drain_right.n10 0.388379
R700 drain_right.n46 drain_right.n45 0.388379
R701 drain_right.n122 drain_right.n121 0.388379
R702 drain_right.n88 drain_right.n86 0.388379
R703 drain_right.n70 drain_right.n66 0.352482
R704 drain_right.n22 drain_right.n17 0.155672
R705 drain_right.n29 drain_right.n17 0.155672
R706 drain_right.n30 drain_right.n29 0.155672
R707 drain_right.n30 drain_right.n13 0.155672
R708 drain_right.n37 drain_right.n13 0.155672
R709 drain_right.n38 drain_right.n37 0.155672
R710 drain_right.n38 drain_right.n9 0.155672
R711 drain_right.n47 drain_right.n9 0.155672
R712 drain_right.n48 drain_right.n47 0.155672
R713 drain_right.n48 drain_right.n5 0.155672
R714 drain_right.n55 drain_right.n5 0.155672
R715 drain_right.n56 drain_right.n55 0.155672
R716 drain_right.n56 drain_right.n1 0.155672
R717 drain_right.n63 drain_right.n1 0.155672
R718 drain_right.n139 drain_right.n77 0.155672
R719 drain_right.n132 drain_right.n77 0.155672
R720 drain_right.n132 drain_right.n131 0.155672
R721 drain_right.n131 drain_right.n81 0.155672
R722 drain_right.n124 drain_right.n81 0.155672
R723 drain_right.n124 drain_right.n123 0.155672
R724 drain_right.n123 drain_right.n85 0.155672
R725 drain_right.n115 drain_right.n85 0.155672
R726 drain_right.n115 drain_right.n114 0.155672
R727 drain_right.n114 drain_right.n90 0.155672
R728 drain_right.n107 drain_right.n90 0.155672
R729 drain_right.n107 drain_right.n106 0.155672
R730 drain_right.n106 drain_right.n94 0.155672
R731 drain_right.n99 drain_right.n94 0.155672
R732 drain_right.n70 drain_right.n69 0.0809298
R733 plus.n3 plus.t1 1125.4
R734 plus.n15 plus.t12 1125.4
R735 plus.n20 plus.t10 1125.4
R736 plus.n32 plus.t2 1125.4
R737 plus.n1 plus.t13 1068.43
R738 plus.n4 plus.t5 1068.43
R739 plus.n6 plus.t9 1068.43
R740 plus.n12 plus.t3 1068.43
R741 plus.n14 plus.t8 1068.43
R742 plus.n18 plus.t6 1068.43
R743 plus.n21 plus.t4 1068.43
R744 plus.n23 plus.t11 1068.43
R745 plus.n29 plus.t0 1068.43
R746 plus.n31 plus.t7 1068.43
R747 plus.n3 plus.n2 161.489
R748 plus.n20 plus.n19 161.489
R749 plus.n5 plus.n2 161.3
R750 plus.n8 plus.n7 161.3
R751 plus.n9 plus.n1 161.3
R752 plus.n11 plus.n10 161.3
R753 plus.n13 plus.n0 161.3
R754 plus.n16 plus.n15 161.3
R755 plus.n22 plus.n19 161.3
R756 plus.n25 plus.n24 161.3
R757 plus.n26 plus.n18 161.3
R758 plus.n28 plus.n27 161.3
R759 plus.n30 plus.n17 161.3
R760 plus.n33 plus.n32 161.3
R761 plus.n7 plus.n1 73.0308
R762 plus.n11 plus.n1 73.0308
R763 plus.n28 plus.n18 73.0308
R764 plus.n24 plus.n18 73.0308
R765 plus.n6 plus.n5 54.0429
R766 plus.n13 plus.n12 54.0429
R767 plus.n30 plus.n29 54.0429
R768 plus.n23 plus.n22 54.0429
R769 plus.n5 plus.n4 37.9763
R770 plus.n14 plus.n13 37.9763
R771 plus.n31 plus.n30 37.9763
R772 plus.n22 plus.n21 37.9763
R773 plus.n4 plus.n3 35.055
R774 plus.n15 plus.n14 35.055
R775 plus.n32 plus.n31 35.055
R776 plus.n21 plus.n20 35.055
R777 plus plus.n33 29.5691
R778 plus.n7 plus.n6 18.9884
R779 plus.n12 plus.n11 18.9884
R780 plus.n29 plus.n28 18.9884
R781 plus.n24 plus.n23 18.9884
R782 plus plus.n16 12.1804
R783 plus.n8 plus.n2 0.189894
R784 plus.n9 plus.n8 0.189894
R785 plus.n10 plus.n9 0.189894
R786 plus.n10 plus.n0 0.189894
R787 plus.n16 plus.n0 0.189894
R788 plus.n33 plus.n17 0.189894
R789 plus.n27 plus.n17 0.189894
R790 plus.n27 plus.n26 0.189894
R791 plus.n26 plus.n25 0.189894
R792 plus.n25 plus.n19 0.189894
R793 drain_left.n60 drain_left.n0 289.615
R794 drain_left.n131 drain_left.n71 289.615
R795 drain_left.n20 drain_left.n19 185
R796 drain_left.n25 drain_left.n24 185
R797 drain_left.n27 drain_left.n26 185
R798 drain_left.n16 drain_left.n15 185
R799 drain_left.n33 drain_left.n32 185
R800 drain_left.n35 drain_left.n34 185
R801 drain_left.n12 drain_left.n11 185
R802 drain_left.n42 drain_left.n41 185
R803 drain_left.n43 drain_left.n10 185
R804 drain_left.n45 drain_left.n44 185
R805 drain_left.n8 drain_left.n7 185
R806 drain_left.n51 drain_left.n50 185
R807 drain_left.n53 drain_left.n52 185
R808 drain_left.n4 drain_left.n3 185
R809 drain_left.n59 drain_left.n58 185
R810 drain_left.n61 drain_left.n60 185
R811 drain_left.n132 drain_left.n131 185
R812 drain_left.n130 drain_left.n129 185
R813 drain_left.n75 drain_left.n74 185
R814 drain_left.n124 drain_left.n123 185
R815 drain_left.n122 drain_left.n121 185
R816 drain_left.n79 drain_left.n78 185
R817 drain_left.n116 drain_left.n115 185
R818 drain_left.n114 drain_left.n81 185
R819 drain_left.n113 drain_left.n112 185
R820 drain_left.n84 drain_left.n82 185
R821 drain_left.n107 drain_left.n106 185
R822 drain_left.n105 drain_left.n104 185
R823 drain_left.n88 drain_left.n87 185
R824 drain_left.n99 drain_left.n98 185
R825 drain_left.n97 drain_left.n96 185
R826 drain_left.n92 drain_left.n91 185
R827 drain_left.n21 drain_left.t11 149.524
R828 drain_left.n93 drain_left.t12 149.524
R829 drain_left.n25 drain_left.n19 104.615
R830 drain_left.n26 drain_left.n25 104.615
R831 drain_left.n26 drain_left.n15 104.615
R832 drain_left.n33 drain_left.n15 104.615
R833 drain_left.n34 drain_left.n33 104.615
R834 drain_left.n34 drain_left.n11 104.615
R835 drain_left.n42 drain_left.n11 104.615
R836 drain_left.n43 drain_left.n42 104.615
R837 drain_left.n44 drain_left.n43 104.615
R838 drain_left.n44 drain_left.n7 104.615
R839 drain_left.n51 drain_left.n7 104.615
R840 drain_left.n52 drain_left.n51 104.615
R841 drain_left.n52 drain_left.n3 104.615
R842 drain_left.n59 drain_left.n3 104.615
R843 drain_left.n60 drain_left.n59 104.615
R844 drain_left.n131 drain_left.n130 104.615
R845 drain_left.n130 drain_left.n74 104.615
R846 drain_left.n123 drain_left.n74 104.615
R847 drain_left.n123 drain_left.n122 104.615
R848 drain_left.n122 drain_left.n78 104.615
R849 drain_left.n115 drain_left.n78 104.615
R850 drain_left.n115 drain_left.n114 104.615
R851 drain_left.n114 drain_left.n113 104.615
R852 drain_left.n113 drain_left.n82 104.615
R853 drain_left.n106 drain_left.n82 104.615
R854 drain_left.n106 drain_left.n105 104.615
R855 drain_left.n105 drain_left.n87 104.615
R856 drain_left.n98 drain_left.n87 104.615
R857 drain_left.n98 drain_left.n97 104.615
R858 drain_left.n97 drain_left.n91 104.615
R859 drain_left.n69 drain_left.n67 60.0956
R860 drain_left.n139 drain_left.n138 59.5527
R861 drain_left.n137 drain_left.n136 59.5527
R862 drain_left.n69 drain_left.n68 59.5525
R863 drain_left.n66 drain_left.n65 59.5525
R864 drain_left.n141 drain_left.n140 59.5525
R865 drain_left.t11 drain_left.n19 52.3082
R866 drain_left.t12 drain_left.n91 52.3082
R867 drain_left.n66 drain_left.n64 47.08
R868 drain_left.n137 drain_left.n135 47.08
R869 drain_left drain_left.n70 30.4899
R870 drain_left.n45 drain_left.n10 13.1884
R871 drain_left.n116 drain_left.n81 13.1884
R872 drain_left.n41 drain_left.n40 12.8005
R873 drain_left.n46 drain_left.n8 12.8005
R874 drain_left.n117 drain_left.n79 12.8005
R875 drain_left.n112 drain_left.n83 12.8005
R876 drain_left.n39 drain_left.n12 12.0247
R877 drain_left.n50 drain_left.n49 12.0247
R878 drain_left.n121 drain_left.n120 12.0247
R879 drain_left.n111 drain_left.n84 12.0247
R880 drain_left.n36 drain_left.n35 11.249
R881 drain_left.n53 drain_left.n6 11.249
R882 drain_left.n124 drain_left.n77 11.249
R883 drain_left.n108 drain_left.n107 11.249
R884 drain_left.n32 drain_left.n14 10.4732
R885 drain_left.n54 drain_left.n4 10.4732
R886 drain_left.n125 drain_left.n75 10.4732
R887 drain_left.n104 drain_left.n86 10.4732
R888 drain_left.n21 drain_left.n20 10.2747
R889 drain_left.n93 drain_left.n92 10.2747
R890 drain_left.n31 drain_left.n16 9.69747
R891 drain_left.n58 drain_left.n57 9.69747
R892 drain_left.n129 drain_left.n128 9.69747
R893 drain_left.n103 drain_left.n88 9.69747
R894 drain_left.n64 drain_left.n63 9.45567
R895 drain_left.n135 drain_left.n134 9.45567
R896 drain_left.n63 drain_left.n62 9.3005
R897 drain_left.n2 drain_left.n1 9.3005
R898 drain_left.n57 drain_left.n56 9.3005
R899 drain_left.n55 drain_left.n54 9.3005
R900 drain_left.n6 drain_left.n5 9.3005
R901 drain_left.n49 drain_left.n48 9.3005
R902 drain_left.n47 drain_left.n46 9.3005
R903 drain_left.n23 drain_left.n22 9.3005
R904 drain_left.n18 drain_left.n17 9.3005
R905 drain_left.n29 drain_left.n28 9.3005
R906 drain_left.n31 drain_left.n30 9.3005
R907 drain_left.n14 drain_left.n13 9.3005
R908 drain_left.n37 drain_left.n36 9.3005
R909 drain_left.n39 drain_left.n38 9.3005
R910 drain_left.n40 drain_left.n9 9.3005
R911 drain_left.n95 drain_left.n94 9.3005
R912 drain_left.n90 drain_left.n89 9.3005
R913 drain_left.n101 drain_left.n100 9.3005
R914 drain_left.n103 drain_left.n102 9.3005
R915 drain_left.n86 drain_left.n85 9.3005
R916 drain_left.n109 drain_left.n108 9.3005
R917 drain_left.n111 drain_left.n110 9.3005
R918 drain_left.n83 drain_left.n80 9.3005
R919 drain_left.n134 drain_left.n133 9.3005
R920 drain_left.n73 drain_left.n72 9.3005
R921 drain_left.n128 drain_left.n127 9.3005
R922 drain_left.n126 drain_left.n125 9.3005
R923 drain_left.n77 drain_left.n76 9.3005
R924 drain_left.n120 drain_left.n119 9.3005
R925 drain_left.n118 drain_left.n117 9.3005
R926 drain_left.n28 drain_left.n27 8.92171
R927 drain_left.n61 drain_left.n2 8.92171
R928 drain_left.n132 drain_left.n73 8.92171
R929 drain_left.n100 drain_left.n99 8.92171
R930 drain_left.n24 drain_left.n18 8.14595
R931 drain_left.n62 drain_left.n0 8.14595
R932 drain_left.n133 drain_left.n71 8.14595
R933 drain_left.n96 drain_left.n90 8.14595
R934 drain_left.n23 drain_left.n20 7.3702
R935 drain_left.n95 drain_left.n92 7.3702
R936 drain_left drain_left.n141 6.19632
R937 drain_left.n24 drain_left.n23 5.81868
R938 drain_left.n64 drain_left.n0 5.81868
R939 drain_left.n135 drain_left.n71 5.81868
R940 drain_left.n96 drain_left.n95 5.81868
R941 drain_left.n27 drain_left.n18 5.04292
R942 drain_left.n62 drain_left.n61 5.04292
R943 drain_left.n133 drain_left.n132 5.04292
R944 drain_left.n99 drain_left.n90 5.04292
R945 drain_left.n28 drain_left.n16 4.26717
R946 drain_left.n58 drain_left.n2 4.26717
R947 drain_left.n129 drain_left.n73 4.26717
R948 drain_left.n100 drain_left.n88 4.26717
R949 drain_left.n32 drain_left.n31 3.49141
R950 drain_left.n57 drain_left.n4 3.49141
R951 drain_left.n128 drain_left.n75 3.49141
R952 drain_left.n104 drain_left.n103 3.49141
R953 drain_left.n22 drain_left.n21 2.84303
R954 drain_left.n94 drain_left.n93 2.84303
R955 drain_left.n35 drain_left.n14 2.71565
R956 drain_left.n54 drain_left.n53 2.71565
R957 drain_left.n125 drain_left.n124 2.71565
R958 drain_left.n107 drain_left.n86 2.71565
R959 drain_left.n36 drain_left.n12 1.93989
R960 drain_left.n50 drain_left.n6 1.93989
R961 drain_left.n121 drain_left.n77 1.93989
R962 drain_left.n108 drain_left.n84 1.93989
R963 drain_left.n67 drain_left.t9 1.6505
R964 drain_left.n67 drain_left.t3 1.6505
R965 drain_left.n68 drain_left.t7 1.6505
R966 drain_left.n68 drain_left.t2 1.6505
R967 drain_left.n65 drain_left.t6 1.6505
R968 drain_left.n65 drain_left.t13 1.6505
R969 drain_left.n140 drain_left.t5 1.6505
R970 drain_left.n140 drain_left.t1 1.6505
R971 drain_left.n138 drain_left.t0 1.6505
R972 drain_left.n138 drain_left.t10 1.6505
R973 drain_left.n136 drain_left.t8 1.6505
R974 drain_left.n136 drain_left.t4 1.6505
R975 drain_left.n41 drain_left.n39 1.16414
R976 drain_left.n49 drain_left.n8 1.16414
R977 drain_left.n120 drain_left.n79 1.16414
R978 drain_left.n112 drain_left.n111 1.16414
R979 drain_left.n139 drain_left.n137 0.543603
R980 drain_left.n141 drain_left.n139 0.543603
R981 drain_left.n40 drain_left.n10 0.388379
R982 drain_left.n46 drain_left.n45 0.388379
R983 drain_left.n117 drain_left.n116 0.388379
R984 drain_left.n83 drain_left.n81 0.388379
R985 drain_left.n70 drain_left.n66 0.352482
R986 drain_left.n22 drain_left.n17 0.155672
R987 drain_left.n29 drain_left.n17 0.155672
R988 drain_left.n30 drain_left.n29 0.155672
R989 drain_left.n30 drain_left.n13 0.155672
R990 drain_left.n37 drain_left.n13 0.155672
R991 drain_left.n38 drain_left.n37 0.155672
R992 drain_left.n38 drain_left.n9 0.155672
R993 drain_left.n47 drain_left.n9 0.155672
R994 drain_left.n48 drain_left.n47 0.155672
R995 drain_left.n48 drain_left.n5 0.155672
R996 drain_left.n55 drain_left.n5 0.155672
R997 drain_left.n56 drain_left.n55 0.155672
R998 drain_left.n56 drain_left.n1 0.155672
R999 drain_left.n63 drain_left.n1 0.155672
R1000 drain_left.n134 drain_left.n72 0.155672
R1001 drain_left.n127 drain_left.n72 0.155672
R1002 drain_left.n127 drain_left.n126 0.155672
R1003 drain_left.n126 drain_left.n76 0.155672
R1004 drain_left.n119 drain_left.n76 0.155672
R1005 drain_left.n119 drain_left.n118 0.155672
R1006 drain_left.n118 drain_left.n80 0.155672
R1007 drain_left.n110 drain_left.n80 0.155672
R1008 drain_left.n110 drain_left.n109 0.155672
R1009 drain_left.n109 drain_left.n85 0.155672
R1010 drain_left.n102 drain_left.n85 0.155672
R1011 drain_left.n102 drain_left.n101 0.155672
R1012 drain_left.n101 drain_left.n89 0.155672
R1013 drain_left.n94 drain_left.n89 0.155672
R1014 drain_left.n70 drain_left.n69 0.0809298
C0 minus plus 5.29917f
C1 source plus 4.9462f
C2 minus drain_right 5.26913f
C3 source drain_right 28.0045f
C4 drain_left minus 0.171678f
C5 drain_left source 28.015f
C6 source minus 4.931509f
C7 drain_right plus 0.323388f
C8 drain_left plus 5.43295f
C9 drain_left drain_right 0.883729f
C10 drain_right a_n1724_n3288# 7.36899f
C11 drain_left a_n1724_n3288# 7.641521f
C12 source a_n1724_n3288# 6.19225f
C13 minus a_n1724_n3288# 6.704053f
C14 plus a_n1724_n3288# 8.679029f
C15 drain_left.n0 a_n1724_n3288# 0.040782f
C16 drain_left.n1 a_n1724_n3288# 0.030787f
C17 drain_left.n2 a_n1724_n3288# 0.016544f
C18 drain_left.n3 a_n1724_n3288# 0.039103f
C19 drain_left.n4 a_n1724_n3288# 0.017517f
C20 drain_left.n5 a_n1724_n3288# 0.030787f
C21 drain_left.n6 a_n1724_n3288# 0.016544f
C22 drain_left.n7 a_n1724_n3288# 0.039103f
C23 drain_left.n8 a_n1724_n3288# 0.017517f
C24 drain_left.n9 a_n1724_n3288# 0.030787f
C25 drain_left.n10 a_n1724_n3288# 0.01703f
C26 drain_left.n11 a_n1724_n3288# 0.039103f
C27 drain_left.n12 a_n1724_n3288# 0.017517f
C28 drain_left.n13 a_n1724_n3288# 0.030787f
C29 drain_left.n14 a_n1724_n3288# 0.016544f
C30 drain_left.n15 a_n1724_n3288# 0.039103f
C31 drain_left.n16 a_n1724_n3288# 0.017517f
C32 drain_left.n17 a_n1724_n3288# 0.030787f
C33 drain_left.n18 a_n1724_n3288# 0.016544f
C34 drain_left.n19 a_n1724_n3288# 0.029327f
C35 drain_left.n20 a_n1724_n3288# 0.027643f
C36 drain_left.t11 a_n1724_n3288# 0.066043f
C37 drain_left.n21 a_n1724_n3288# 0.221972f
C38 drain_left.n22 a_n1724_n3288# 1.55316f
C39 drain_left.n23 a_n1724_n3288# 0.016544f
C40 drain_left.n24 a_n1724_n3288# 0.017517f
C41 drain_left.n25 a_n1724_n3288# 0.039103f
C42 drain_left.n26 a_n1724_n3288# 0.039103f
C43 drain_left.n27 a_n1724_n3288# 0.017517f
C44 drain_left.n28 a_n1724_n3288# 0.016544f
C45 drain_left.n29 a_n1724_n3288# 0.030787f
C46 drain_left.n30 a_n1724_n3288# 0.030787f
C47 drain_left.n31 a_n1724_n3288# 0.016544f
C48 drain_left.n32 a_n1724_n3288# 0.017517f
C49 drain_left.n33 a_n1724_n3288# 0.039103f
C50 drain_left.n34 a_n1724_n3288# 0.039103f
C51 drain_left.n35 a_n1724_n3288# 0.017517f
C52 drain_left.n36 a_n1724_n3288# 0.016544f
C53 drain_left.n37 a_n1724_n3288# 0.030787f
C54 drain_left.n38 a_n1724_n3288# 0.030787f
C55 drain_left.n39 a_n1724_n3288# 0.016544f
C56 drain_left.n40 a_n1724_n3288# 0.016544f
C57 drain_left.n41 a_n1724_n3288# 0.017517f
C58 drain_left.n42 a_n1724_n3288# 0.039103f
C59 drain_left.n43 a_n1724_n3288# 0.039103f
C60 drain_left.n44 a_n1724_n3288# 0.039103f
C61 drain_left.n45 a_n1724_n3288# 0.01703f
C62 drain_left.n46 a_n1724_n3288# 0.016544f
C63 drain_left.n47 a_n1724_n3288# 0.030787f
C64 drain_left.n48 a_n1724_n3288# 0.030787f
C65 drain_left.n49 a_n1724_n3288# 0.016544f
C66 drain_left.n50 a_n1724_n3288# 0.017517f
C67 drain_left.n51 a_n1724_n3288# 0.039103f
C68 drain_left.n52 a_n1724_n3288# 0.039103f
C69 drain_left.n53 a_n1724_n3288# 0.017517f
C70 drain_left.n54 a_n1724_n3288# 0.016544f
C71 drain_left.n55 a_n1724_n3288# 0.030787f
C72 drain_left.n56 a_n1724_n3288# 0.030787f
C73 drain_left.n57 a_n1724_n3288# 0.016544f
C74 drain_left.n58 a_n1724_n3288# 0.017517f
C75 drain_left.n59 a_n1724_n3288# 0.039103f
C76 drain_left.n60 a_n1724_n3288# 0.080244f
C77 drain_left.n61 a_n1724_n3288# 0.017517f
C78 drain_left.n62 a_n1724_n3288# 0.016544f
C79 drain_left.n63 a_n1724_n3288# 0.066116f
C80 drain_left.n64 a_n1724_n3288# 0.06686f
C81 drain_left.t6 a_n1724_n3288# 0.291947f
C82 drain_left.t13 a_n1724_n3288# 0.291947f
C83 drain_left.n65 a_n1724_n3288# 2.59788f
C84 drain_left.n66 a_n1724_n3288# 0.458207f
C85 drain_left.t9 a_n1724_n3288# 0.291947f
C86 drain_left.t3 a_n1724_n3288# 0.291947f
C87 drain_left.n67 a_n1724_n3288# 2.6013f
C88 drain_left.t7 a_n1724_n3288# 0.291947f
C89 drain_left.t2 a_n1724_n3288# 0.291947f
C90 drain_left.n68 a_n1724_n3288# 2.59788f
C91 drain_left.n69 a_n1724_n3288# 0.704231f
C92 drain_left.n70 a_n1724_n3288# 1.46446f
C93 drain_left.n71 a_n1724_n3288# 0.040782f
C94 drain_left.n72 a_n1724_n3288# 0.030787f
C95 drain_left.n73 a_n1724_n3288# 0.016544f
C96 drain_left.n74 a_n1724_n3288# 0.039103f
C97 drain_left.n75 a_n1724_n3288# 0.017517f
C98 drain_left.n76 a_n1724_n3288# 0.030787f
C99 drain_left.n77 a_n1724_n3288# 0.016544f
C100 drain_left.n78 a_n1724_n3288# 0.039103f
C101 drain_left.n79 a_n1724_n3288# 0.017517f
C102 drain_left.n80 a_n1724_n3288# 0.030787f
C103 drain_left.n81 a_n1724_n3288# 0.01703f
C104 drain_left.n82 a_n1724_n3288# 0.039103f
C105 drain_left.n83 a_n1724_n3288# 0.016544f
C106 drain_left.n84 a_n1724_n3288# 0.017517f
C107 drain_left.n85 a_n1724_n3288# 0.030787f
C108 drain_left.n86 a_n1724_n3288# 0.016544f
C109 drain_left.n87 a_n1724_n3288# 0.039103f
C110 drain_left.n88 a_n1724_n3288# 0.017517f
C111 drain_left.n89 a_n1724_n3288# 0.030787f
C112 drain_left.n90 a_n1724_n3288# 0.016544f
C113 drain_left.n91 a_n1724_n3288# 0.029327f
C114 drain_left.n92 a_n1724_n3288# 0.027643f
C115 drain_left.t12 a_n1724_n3288# 0.066043f
C116 drain_left.n93 a_n1724_n3288# 0.221972f
C117 drain_left.n94 a_n1724_n3288# 1.55316f
C118 drain_left.n95 a_n1724_n3288# 0.016544f
C119 drain_left.n96 a_n1724_n3288# 0.017517f
C120 drain_left.n97 a_n1724_n3288# 0.039103f
C121 drain_left.n98 a_n1724_n3288# 0.039103f
C122 drain_left.n99 a_n1724_n3288# 0.017517f
C123 drain_left.n100 a_n1724_n3288# 0.016544f
C124 drain_left.n101 a_n1724_n3288# 0.030787f
C125 drain_left.n102 a_n1724_n3288# 0.030787f
C126 drain_left.n103 a_n1724_n3288# 0.016544f
C127 drain_left.n104 a_n1724_n3288# 0.017517f
C128 drain_left.n105 a_n1724_n3288# 0.039103f
C129 drain_left.n106 a_n1724_n3288# 0.039103f
C130 drain_left.n107 a_n1724_n3288# 0.017517f
C131 drain_left.n108 a_n1724_n3288# 0.016544f
C132 drain_left.n109 a_n1724_n3288# 0.030787f
C133 drain_left.n110 a_n1724_n3288# 0.030787f
C134 drain_left.n111 a_n1724_n3288# 0.016544f
C135 drain_left.n112 a_n1724_n3288# 0.017517f
C136 drain_left.n113 a_n1724_n3288# 0.039103f
C137 drain_left.n114 a_n1724_n3288# 0.039103f
C138 drain_left.n115 a_n1724_n3288# 0.039103f
C139 drain_left.n116 a_n1724_n3288# 0.01703f
C140 drain_left.n117 a_n1724_n3288# 0.016544f
C141 drain_left.n118 a_n1724_n3288# 0.030787f
C142 drain_left.n119 a_n1724_n3288# 0.030787f
C143 drain_left.n120 a_n1724_n3288# 0.016544f
C144 drain_left.n121 a_n1724_n3288# 0.017517f
C145 drain_left.n122 a_n1724_n3288# 0.039103f
C146 drain_left.n123 a_n1724_n3288# 0.039103f
C147 drain_left.n124 a_n1724_n3288# 0.017517f
C148 drain_left.n125 a_n1724_n3288# 0.016544f
C149 drain_left.n126 a_n1724_n3288# 0.030787f
C150 drain_left.n127 a_n1724_n3288# 0.030787f
C151 drain_left.n128 a_n1724_n3288# 0.016544f
C152 drain_left.n129 a_n1724_n3288# 0.017517f
C153 drain_left.n130 a_n1724_n3288# 0.039103f
C154 drain_left.n131 a_n1724_n3288# 0.080244f
C155 drain_left.n132 a_n1724_n3288# 0.017517f
C156 drain_left.n133 a_n1724_n3288# 0.016544f
C157 drain_left.n134 a_n1724_n3288# 0.066116f
C158 drain_left.n135 a_n1724_n3288# 0.06686f
C159 drain_left.t8 a_n1724_n3288# 0.291947f
C160 drain_left.t4 a_n1724_n3288# 0.291947f
C161 drain_left.n136 a_n1724_n3288# 2.59789f
C162 drain_left.n137 a_n1724_n3288# 0.475128f
C163 drain_left.t0 a_n1724_n3288# 0.291947f
C164 drain_left.t10 a_n1724_n3288# 0.291947f
C165 drain_left.n138 a_n1724_n3288# 2.59789f
C166 drain_left.n139 a_n1724_n3288# 0.366127f
C167 drain_left.t5 a_n1724_n3288# 0.291947f
C168 drain_left.t1 a_n1724_n3288# 0.291947f
C169 drain_left.n140 a_n1724_n3288# 2.59788f
C170 drain_left.n141 a_n1724_n3288# 0.622398f
C171 plus.n0 a_n1724_n3288# 0.052065f
C172 plus.t8 a_n1724_n3288# 0.529658f
C173 plus.t3 a_n1724_n3288# 0.529658f
C174 plus.t13 a_n1724_n3288# 0.529658f
C175 plus.n1 a_n1724_n3288# 0.227384f
C176 plus.n2 a_n1724_n3288# 0.122666f
C177 plus.t9 a_n1724_n3288# 0.529658f
C178 plus.t5 a_n1724_n3288# 0.529658f
C179 plus.t1 a_n1724_n3288# 0.540602f
C180 plus.n3 a_n1724_n3288# 0.226795f
C181 plus.n4 a_n1724_n3288# 0.210112f
C182 plus.n5 a_n1724_n3288# 0.021445f
C183 plus.n6 a_n1724_n3288# 0.210112f
C184 plus.n7 a_n1724_n3288# 0.021445f
C185 plus.n8 a_n1724_n3288# 0.052065f
C186 plus.n9 a_n1724_n3288# 0.052065f
C187 plus.n10 a_n1724_n3288# 0.052065f
C188 plus.n11 a_n1724_n3288# 0.021445f
C189 plus.n12 a_n1724_n3288# 0.210112f
C190 plus.n13 a_n1724_n3288# 0.021445f
C191 plus.n14 a_n1724_n3288# 0.210112f
C192 plus.t12 a_n1724_n3288# 0.540602f
C193 plus.n15 a_n1724_n3288# 0.226712f
C194 plus.n16 a_n1724_n3288# 0.587069f
C195 plus.n17 a_n1724_n3288# 0.052065f
C196 plus.t2 a_n1724_n3288# 0.540602f
C197 plus.t7 a_n1724_n3288# 0.529658f
C198 plus.t0 a_n1724_n3288# 0.529658f
C199 plus.t6 a_n1724_n3288# 0.529658f
C200 plus.n18 a_n1724_n3288# 0.227384f
C201 plus.n19 a_n1724_n3288# 0.122666f
C202 plus.t11 a_n1724_n3288# 0.529658f
C203 plus.t4 a_n1724_n3288# 0.529658f
C204 plus.t10 a_n1724_n3288# 0.540602f
C205 plus.n20 a_n1724_n3288# 0.226795f
C206 plus.n21 a_n1724_n3288# 0.210112f
C207 plus.n22 a_n1724_n3288# 0.021445f
C208 plus.n23 a_n1724_n3288# 0.210112f
C209 plus.n24 a_n1724_n3288# 0.021445f
C210 plus.n25 a_n1724_n3288# 0.052065f
C211 plus.n26 a_n1724_n3288# 0.052065f
C212 plus.n27 a_n1724_n3288# 0.052065f
C213 plus.n28 a_n1724_n3288# 0.021445f
C214 plus.n29 a_n1724_n3288# 0.210112f
C215 plus.n30 a_n1724_n3288# 0.021445f
C216 plus.n31 a_n1724_n3288# 0.210112f
C217 plus.n32 a_n1724_n3288# 0.226712f
C218 plus.n33 a_n1724_n3288# 1.52237f
C219 drain_right.n0 a_n1724_n3288# 0.040807f
C220 drain_right.n1 a_n1724_n3288# 0.030806f
C221 drain_right.n2 a_n1724_n3288# 0.016554f
C222 drain_right.n3 a_n1724_n3288# 0.039127f
C223 drain_right.n4 a_n1724_n3288# 0.017528f
C224 drain_right.n5 a_n1724_n3288# 0.030806f
C225 drain_right.n6 a_n1724_n3288# 0.016554f
C226 drain_right.n7 a_n1724_n3288# 0.039127f
C227 drain_right.n8 a_n1724_n3288# 0.017528f
C228 drain_right.n9 a_n1724_n3288# 0.030806f
C229 drain_right.n10 a_n1724_n3288# 0.017041f
C230 drain_right.n11 a_n1724_n3288# 0.039127f
C231 drain_right.n12 a_n1724_n3288# 0.017528f
C232 drain_right.n13 a_n1724_n3288# 0.030806f
C233 drain_right.n14 a_n1724_n3288# 0.016554f
C234 drain_right.n15 a_n1724_n3288# 0.039127f
C235 drain_right.n16 a_n1724_n3288# 0.017528f
C236 drain_right.n17 a_n1724_n3288# 0.030806f
C237 drain_right.n18 a_n1724_n3288# 0.016554f
C238 drain_right.n19 a_n1724_n3288# 0.029345f
C239 drain_right.n20 a_n1724_n3288# 0.02766f
C240 drain_right.t12 a_n1724_n3288# 0.066083f
C241 drain_right.n21 a_n1724_n3288# 0.222108f
C242 drain_right.n22 a_n1724_n3288# 1.55411f
C243 drain_right.n23 a_n1724_n3288# 0.016554f
C244 drain_right.n24 a_n1724_n3288# 0.017528f
C245 drain_right.n25 a_n1724_n3288# 0.039127f
C246 drain_right.n26 a_n1724_n3288# 0.039127f
C247 drain_right.n27 a_n1724_n3288# 0.017528f
C248 drain_right.n28 a_n1724_n3288# 0.016554f
C249 drain_right.n29 a_n1724_n3288# 0.030806f
C250 drain_right.n30 a_n1724_n3288# 0.030806f
C251 drain_right.n31 a_n1724_n3288# 0.016554f
C252 drain_right.n32 a_n1724_n3288# 0.017528f
C253 drain_right.n33 a_n1724_n3288# 0.039127f
C254 drain_right.n34 a_n1724_n3288# 0.039127f
C255 drain_right.n35 a_n1724_n3288# 0.017528f
C256 drain_right.n36 a_n1724_n3288# 0.016554f
C257 drain_right.n37 a_n1724_n3288# 0.030806f
C258 drain_right.n38 a_n1724_n3288# 0.030806f
C259 drain_right.n39 a_n1724_n3288# 0.016554f
C260 drain_right.n40 a_n1724_n3288# 0.016554f
C261 drain_right.n41 a_n1724_n3288# 0.017528f
C262 drain_right.n42 a_n1724_n3288# 0.039127f
C263 drain_right.n43 a_n1724_n3288# 0.039127f
C264 drain_right.n44 a_n1724_n3288# 0.039127f
C265 drain_right.n45 a_n1724_n3288# 0.017041f
C266 drain_right.n46 a_n1724_n3288# 0.016554f
C267 drain_right.n47 a_n1724_n3288# 0.030806f
C268 drain_right.n48 a_n1724_n3288# 0.030806f
C269 drain_right.n49 a_n1724_n3288# 0.016554f
C270 drain_right.n50 a_n1724_n3288# 0.017528f
C271 drain_right.n51 a_n1724_n3288# 0.039127f
C272 drain_right.n52 a_n1724_n3288# 0.039127f
C273 drain_right.n53 a_n1724_n3288# 0.017528f
C274 drain_right.n54 a_n1724_n3288# 0.016554f
C275 drain_right.n55 a_n1724_n3288# 0.030806f
C276 drain_right.n56 a_n1724_n3288# 0.030806f
C277 drain_right.n57 a_n1724_n3288# 0.016554f
C278 drain_right.n58 a_n1724_n3288# 0.017528f
C279 drain_right.n59 a_n1724_n3288# 0.039127f
C280 drain_right.n60 a_n1724_n3288# 0.080293f
C281 drain_right.n61 a_n1724_n3288# 0.017528f
C282 drain_right.n62 a_n1724_n3288# 0.016554f
C283 drain_right.n63 a_n1724_n3288# 0.066157f
C284 drain_right.n64 a_n1724_n3288# 0.066901f
C285 drain_right.t3 a_n1724_n3288# 0.292127f
C286 drain_right.t13 a_n1724_n3288# 0.292127f
C287 drain_right.n65 a_n1724_n3288# 2.59948f
C288 drain_right.n66 a_n1724_n3288# 0.458489f
C289 drain_right.t2 a_n1724_n3288# 0.292127f
C290 drain_right.t8 a_n1724_n3288# 0.292127f
C291 drain_right.n67 a_n1724_n3288# 2.6029f
C292 drain_right.t4 a_n1724_n3288# 0.292127f
C293 drain_right.t7 a_n1724_n3288# 0.292127f
C294 drain_right.n68 a_n1724_n3288# 2.59948f
C295 drain_right.n69 a_n1724_n3288# 0.704664f
C296 drain_right.n70 a_n1724_n3288# 1.40133f
C297 drain_right.t0 a_n1724_n3288# 0.292127f
C298 drain_right.t5 a_n1724_n3288# 0.292127f
C299 drain_right.n71 a_n1724_n3288# 2.6029f
C300 drain_right.t6 a_n1724_n3288# 0.292127f
C301 drain_right.t10 a_n1724_n3288# 0.292127f
C302 drain_right.n72 a_n1724_n3288# 2.59949f
C303 drain_right.n73 a_n1724_n3288# 0.7417f
C304 drain_right.t11 a_n1724_n3288# 0.292127f
C305 drain_right.t1 a_n1724_n3288# 0.292127f
C306 drain_right.n74 a_n1724_n3288# 2.59949f
C307 drain_right.n75 a_n1724_n3288# 0.366352f
C308 drain_right.n76 a_n1724_n3288# 0.040807f
C309 drain_right.n77 a_n1724_n3288# 0.030806f
C310 drain_right.n78 a_n1724_n3288# 0.016554f
C311 drain_right.n79 a_n1724_n3288# 0.039127f
C312 drain_right.n80 a_n1724_n3288# 0.017528f
C313 drain_right.n81 a_n1724_n3288# 0.030806f
C314 drain_right.n82 a_n1724_n3288# 0.016554f
C315 drain_right.n83 a_n1724_n3288# 0.039127f
C316 drain_right.n84 a_n1724_n3288# 0.017528f
C317 drain_right.n85 a_n1724_n3288# 0.030806f
C318 drain_right.n86 a_n1724_n3288# 0.017041f
C319 drain_right.n87 a_n1724_n3288# 0.039127f
C320 drain_right.n88 a_n1724_n3288# 0.016554f
C321 drain_right.n89 a_n1724_n3288# 0.017528f
C322 drain_right.n90 a_n1724_n3288# 0.030806f
C323 drain_right.n91 a_n1724_n3288# 0.016554f
C324 drain_right.n92 a_n1724_n3288# 0.039127f
C325 drain_right.n93 a_n1724_n3288# 0.017528f
C326 drain_right.n94 a_n1724_n3288# 0.030806f
C327 drain_right.n95 a_n1724_n3288# 0.016554f
C328 drain_right.n96 a_n1724_n3288# 0.029345f
C329 drain_right.n97 a_n1724_n3288# 0.02766f
C330 drain_right.t9 a_n1724_n3288# 0.066083f
C331 drain_right.n98 a_n1724_n3288# 0.222108f
C332 drain_right.n99 a_n1724_n3288# 1.55411f
C333 drain_right.n100 a_n1724_n3288# 0.016554f
C334 drain_right.n101 a_n1724_n3288# 0.017528f
C335 drain_right.n102 a_n1724_n3288# 0.039127f
C336 drain_right.n103 a_n1724_n3288# 0.039127f
C337 drain_right.n104 a_n1724_n3288# 0.017528f
C338 drain_right.n105 a_n1724_n3288# 0.016554f
C339 drain_right.n106 a_n1724_n3288# 0.030806f
C340 drain_right.n107 a_n1724_n3288# 0.030806f
C341 drain_right.n108 a_n1724_n3288# 0.016554f
C342 drain_right.n109 a_n1724_n3288# 0.017528f
C343 drain_right.n110 a_n1724_n3288# 0.039127f
C344 drain_right.n111 a_n1724_n3288# 0.039127f
C345 drain_right.n112 a_n1724_n3288# 0.017528f
C346 drain_right.n113 a_n1724_n3288# 0.016554f
C347 drain_right.n114 a_n1724_n3288# 0.030806f
C348 drain_right.n115 a_n1724_n3288# 0.030806f
C349 drain_right.n116 a_n1724_n3288# 0.016554f
C350 drain_right.n117 a_n1724_n3288# 0.017528f
C351 drain_right.n118 a_n1724_n3288# 0.039127f
C352 drain_right.n119 a_n1724_n3288# 0.039127f
C353 drain_right.n120 a_n1724_n3288# 0.039127f
C354 drain_right.n121 a_n1724_n3288# 0.017041f
C355 drain_right.n122 a_n1724_n3288# 0.016554f
C356 drain_right.n123 a_n1724_n3288# 0.030806f
C357 drain_right.n124 a_n1724_n3288# 0.030806f
C358 drain_right.n125 a_n1724_n3288# 0.016554f
C359 drain_right.n126 a_n1724_n3288# 0.017528f
C360 drain_right.n127 a_n1724_n3288# 0.039127f
C361 drain_right.n128 a_n1724_n3288# 0.039127f
C362 drain_right.n129 a_n1724_n3288# 0.017528f
C363 drain_right.n130 a_n1724_n3288# 0.016554f
C364 drain_right.n131 a_n1724_n3288# 0.030806f
C365 drain_right.n132 a_n1724_n3288# 0.030806f
C366 drain_right.n133 a_n1724_n3288# 0.016554f
C367 drain_right.n134 a_n1724_n3288# 0.017528f
C368 drain_right.n135 a_n1724_n3288# 0.039127f
C369 drain_right.n136 a_n1724_n3288# 0.080293f
C370 drain_right.n137 a_n1724_n3288# 0.017528f
C371 drain_right.n138 a_n1724_n3288# 0.016554f
C372 drain_right.n139 a_n1724_n3288# 0.066157f
C373 drain_right.n140 a_n1724_n3288# 0.065628f
C374 drain_right.n141 a_n1724_n3288# 0.36734f
C375 source.n0 a_n1724_n3288# 0.042209f
C376 source.n1 a_n1724_n3288# 0.031865f
C377 source.n2 a_n1724_n3288# 0.017123f
C378 source.n3 a_n1724_n3288# 0.040472f
C379 source.n4 a_n1724_n3288# 0.01813f
C380 source.n5 a_n1724_n3288# 0.031865f
C381 source.n6 a_n1724_n3288# 0.017123f
C382 source.n7 a_n1724_n3288# 0.040472f
C383 source.n8 a_n1724_n3288# 0.01813f
C384 source.n9 a_n1724_n3288# 0.031865f
C385 source.n10 a_n1724_n3288# 0.017626f
C386 source.n11 a_n1724_n3288# 0.040472f
C387 source.n12 a_n1724_n3288# 0.017123f
C388 source.n13 a_n1724_n3288# 0.01813f
C389 source.n14 a_n1724_n3288# 0.031865f
C390 source.n15 a_n1724_n3288# 0.017123f
C391 source.n16 a_n1724_n3288# 0.040472f
C392 source.n17 a_n1724_n3288# 0.01813f
C393 source.n18 a_n1724_n3288# 0.031865f
C394 source.n19 a_n1724_n3288# 0.017123f
C395 source.n20 a_n1724_n3288# 0.030354f
C396 source.n21 a_n1724_n3288# 0.028611f
C397 source.t9 a_n1724_n3288# 0.068355f
C398 source.n22 a_n1724_n3288# 0.229743f
C399 source.n23 a_n1724_n3288# 1.60754f
C400 source.n24 a_n1724_n3288# 0.017123f
C401 source.n25 a_n1724_n3288# 0.01813f
C402 source.n26 a_n1724_n3288# 0.040472f
C403 source.n27 a_n1724_n3288# 0.040472f
C404 source.n28 a_n1724_n3288# 0.01813f
C405 source.n29 a_n1724_n3288# 0.017123f
C406 source.n30 a_n1724_n3288# 0.031865f
C407 source.n31 a_n1724_n3288# 0.031865f
C408 source.n32 a_n1724_n3288# 0.017123f
C409 source.n33 a_n1724_n3288# 0.01813f
C410 source.n34 a_n1724_n3288# 0.040472f
C411 source.n35 a_n1724_n3288# 0.040472f
C412 source.n36 a_n1724_n3288# 0.01813f
C413 source.n37 a_n1724_n3288# 0.017123f
C414 source.n38 a_n1724_n3288# 0.031865f
C415 source.n39 a_n1724_n3288# 0.031865f
C416 source.n40 a_n1724_n3288# 0.017123f
C417 source.n41 a_n1724_n3288# 0.01813f
C418 source.n42 a_n1724_n3288# 0.040472f
C419 source.n43 a_n1724_n3288# 0.040472f
C420 source.n44 a_n1724_n3288# 0.040472f
C421 source.n45 a_n1724_n3288# 0.017626f
C422 source.n46 a_n1724_n3288# 0.017123f
C423 source.n47 a_n1724_n3288# 0.031865f
C424 source.n48 a_n1724_n3288# 0.031865f
C425 source.n49 a_n1724_n3288# 0.017123f
C426 source.n50 a_n1724_n3288# 0.01813f
C427 source.n51 a_n1724_n3288# 0.040472f
C428 source.n52 a_n1724_n3288# 0.040472f
C429 source.n53 a_n1724_n3288# 0.01813f
C430 source.n54 a_n1724_n3288# 0.017123f
C431 source.n55 a_n1724_n3288# 0.031865f
C432 source.n56 a_n1724_n3288# 0.031865f
C433 source.n57 a_n1724_n3288# 0.017123f
C434 source.n58 a_n1724_n3288# 0.01813f
C435 source.n59 a_n1724_n3288# 0.040472f
C436 source.n60 a_n1724_n3288# 0.083053f
C437 source.n61 a_n1724_n3288# 0.01813f
C438 source.n62 a_n1724_n3288# 0.017123f
C439 source.n63 a_n1724_n3288# 0.068431f
C440 source.n64 a_n1724_n3288# 0.045836f
C441 source.n65 a_n1724_n3288# 1.28241f
C442 source.t1 a_n1724_n3288# 0.302169f
C443 source.t4 a_n1724_n3288# 0.302169f
C444 source.n66 a_n1724_n3288# 2.58717f
C445 source.n67 a_n1724_n3288# 0.437307f
C446 source.t12 a_n1724_n3288# 0.302169f
C447 source.t5 a_n1724_n3288# 0.302169f
C448 source.n68 a_n1724_n3288# 2.58717f
C449 source.n69 a_n1724_n3288# 0.437307f
C450 source.t6 a_n1724_n3288# 0.302169f
C451 source.t11 a_n1724_n3288# 0.302169f
C452 source.n70 a_n1724_n3288# 2.58717f
C453 source.n71 a_n1724_n3288# 0.457665f
C454 source.n72 a_n1724_n3288# 0.042209f
C455 source.n73 a_n1724_n3288# 0.031865f
C456 source.n74 a_n1724_n3288# 0.017123f
C457 source.n75 a_n1724_n3288# 0.040472f
C458 source.n76 a_n1724_n3288# 0.01813f
C459 source.n77 a_n1724_n3288# 0.031865f
C460 source.n78 a_n1724_n3288# 0.017123f
C461 source.n79 a_n1724_n3288# 0.040472f
C462 source.n80 a_n1724_n3288# 0.01813f
C463 source.n81 a_n1724_n3288# 0.031865f
C464 source.n82 a_n1724_n3288# 0.017626f
C465 source.n83 a_n1724_n3288# 0.040472f
C466 source.n84 a_n1724_n3288# 0.017123f
C467 source.n85 a_n1724_n3288# 0.01813f
C468 source.n86 a_n1724_n3288# 0.031865f
C469 source.n87 a_n1724_n3288# 0.017123f
C470 source.n88 a_n1724_n3288# 0.040472f
C471 source.n89 a_n1724_n3288# 0.01813f
C472 source.n90 a_n1724_n3288# 0.031865f
C473 source.n91 a_n1724_n3288# 0.017123f
C474 source.n92 a_n1724_n3288# 0.030354f
C475 source.n93 a_n1724_n3288# 0.028611f
C476 source.t19 a_n1724_n3288# 0.068355f
C477 source.n94 a_n1724_n3288# 0.229743f
C478 source.n95 a_n1724_n3288# 1.60754f
C479 source.n96 a_n1724_n3288# 0.017123f
C480 source.n97 a_n1724_n3288# 0.01813f
C481 source.n98 a_n1724_n3288# 0.040472f
C482 source.n99 a_n1724_n3288# 0.040472f
C483 source.n100 a_n1724_n3288# 0.01813f
C484 source.n101 a_n1724_n3288# 0.017123f
C485 source.n102 a_n1724_n3288# 0.031865f
C486 source.n103 a_n1724_n3288# 0.031865f
C487 source.n104 a_n1724_n3288# 0.017123f
C488 source.n105 a_n1724_n3288# 0.01813f
C489 source.n106 a_n1724_n3288# 0.040472f
C490 source.n107 a_n1724_n3288# 0.040472f
C491 source.n108 a_n1724_n3288# 0.01813f
C492 source.n109 a_n1724_n3288# 0.017123f
C493 source.n110 a_n1724_n3288# 0.031865f
C494 source.n111 a_n1724_n3288# 0.031865f
C495 source.n112 a_n1724_n3288# 0.017123f
C496 source.n113 a_n1724_n3288# 0.01813f
C497 source.n114 a_n1724_n3288# 0.040472f
C498 source.n115 a_n1724_n3288# 0.040472f
C499 source.n116 a_n1724_n3288# 0.040472f
C500 source.n117 a_n1724_n3288# 0.017626f
C501 source.n118 a_n1724_n3288# 0.017123f
C502 source.n119 a_n1724_n3288# 0.031865f
C503 source.n120 a_n1724_n3288# 0.031865f
C504 source.n121 a_n1724_n3288# 0.017123f
C505 source.n122 a_n1724_n3288# 0.01813f
C506 source.n123 a_n1724_n3288# 0.040472f
C507 source.n124 a_n1724_n3288# 0.040472f
C508 source.n125 a_n1724_n3288# 0.01813f
C509 source.n126 a_n1724_n3288# 0.017123f
C510 source.n127 a_n1724_n3288# 0.031865f
C511 source.n128 a_n1724_n3288# 0.031865f
C512 source.n129 a_n1724_n3288# 0.017123f
C513 source.n130 a_n1724_n3288# 0.01813f
C514 source.n131 a_n1724_n3288# 0.040472f
C515 source.n132 a_n1724_n3288# 0.083053f
C516 source.n133 a_n1724_n3288# 0.01813f
C517 source.n134 a_n1724_n3288# 0.017123f
C518 source.n135 a_n1724_n3288# 0.068431f
C519 source.n136 a_n1724_n3288# 0.045836f
C520 source.n137 a_n1724_n3288# 0.156158f
C521 source.t17 a_n1724_n3288# 0.302169f
C522 source.t14 a_n1724_n3288# 0.302169f
C523 source.n138 a_n1724_n3288# 2.58717f
C524 source.n139 a_n1724_n3288# 0.437307f
C525 source.t16 a_n1724_n3288# 0.302169f
C526 source.t20 a_n1724_n3288# 0.302169f
C527 source.n140 a_n1724_n3288# 2.58717f
C528 source.n141 a_n1724_n3288# 0.437307f
C529 source.t26 a_n1724_n3288# 0.302169f
C530 source.t22 a_n1724_n3288# 0.302169f
C531 source.n142 a_n1724_n3288# 2.58717f
C532 source.n143 a_n1724_n3288# 2.14073f
C533 source.t8 a_n1724_n3288# 0.302169f
C534 source.t10 a_n1724_n3288# 0.302169f
C535 source.n144 a_n1724_n3288# 2.58716f
C536 source.n145 a_n1724_n3288# 2.14075f
C537 source.t2 a_n1724_n3288# 0.302169f
C538 source.t7 a_n1724_n3288# 0.302169f
C539 source.n146 a_n1724_n3288# 2.58716f
C540 source.n147 a_n1724_n3288# 0.437323f
C541 source.t3 a_n1724_n3288# 0.302169f
C542 source.t0 a_n1724_n3288# 0.302169f
C543 source.n148 a_n1724_n3288# 2.58716f
C544 source.n149 a_n1724_n3288# 0.437323f
C545 source.n150 a_n1724_n3288# 0.042209f
C546 source.n151 a_n1724_n3288# 0.031865f
C547 source.n152 a_n1724_n3288# 0.017123f
C548 source.n153 a_n1724_n3288# 0.040472f
C549 source.n154 a_n1724_n3288# 0.01813f
C550 source.n155 a_n1724_n3288# 0.031865f
C551 source.n156 a_n1724_n3288# 0.017123f
C552 source.n157 a_n1724_n3288# 0.040472f
C553 source.n158 a_n1724_n3288# 0.01813f
C554 source.n159 a_n1724_n3288# 0.031865f
C555 source.n160 a_n1724_n3288# 0.017626f
C556 source.n161 a_n1724_n3288# 0.040472f
C557 source.n162 a_n1724_n3288# 0.01813f
C558 source.n163 a_n1724_n3288# 0.031865f
C559 source.n164 a_n1724_n3288# 0.017123f
C560 source.n165 a_n1724_n3288# 0.040472f
C561 source.n166 a_n1724_n3288# 0.01813f
C562 source.n167 a_n1724_n3288# 0.031865f
C563 source.n168 a_n1724_n3288# 0.017123f
C564 source.n169 a_n1724_n3288# 0.030354f
C565 source.n170 a_n1724_n3288# 0.028611f
C566 source.t13 a_n1724_n3288# 0.068355f
C567 source.n171 a_n1724_n3288# 0.229743f
C568 source.n172 a_n1724_n3288# 1.60754f
C569 source.n173 a_n1724_n3288# 0.017123f
C570 source.n174 a_n1724_n3288# 0.01813f
C571 source.n175 a_n1724_n3288# 0.040472f
C572 source.n176 a_n1724_n3288# 0.040472f
C573 source.n177 a_n1724_n3288# 0.01813f
C574 source.n178 a_n1724_n3288# 0.017123f
C575 source.n179 a_n1724_n3288# 0.031865f
C576 source.n180 a_n1724_n3288# 0.031865f
C577 source.n181 a_n1724_n3288# 0.017123f
C578 source.n182 a_n1724_n3288# 0.01813f
C579 source.n183 a_n1724_n3288# 0.040472f
C580 source.n184 a_n1724_n3288# 0.040472f
C581 source.n185 a_n1724_n3288# 0.01813f
C582 source.n186 a_n1724_n3288# 0.017123f
C583 source.n187 a_n1724_n3288# 0.031865f
C584 source.n188 a_n1724_n3288# 0.031865f
C585 source.n189 a_n1724_n3288# 0.017123f
C586 source.n190 a_n1724_n3288# 0.017123f
C587 source.n191 a_n1724_n3288# 0.01813f
C588 source.n192 a_n1724_n3288# 0.040472f
C589 source.n193 a_n1724_n3288# 0.040472f
C590 source.n194 a_n1724_n3288# 0.040472f
C591 source.n195 a_n1724_n3288# 0.017626f
C592 source.n196 a_n1724_n3288# 0.017123f
C593 source.n197 a_n1724_n3288# 0.031865f
C594 source.n198 a_n1724_n3288# 0.031865f
C595 source.n199 a_n1724_n3288# 0.017123f
C596 source.n200 a_n1724_n3288# 0.01813f
C597 source.n201 a_n1724_n3288# 0.040472f
C598 source.n202 a_n1724_n3288# 0.040472f
C599 source.n203 a_n1724_n3288# 0.01813f
C600 source.n204 a_n1724_n3288# 0.017123f
C601 source.n205 a_n1724_n3288# 0.031865f
C602 source.n206 a_n1724_n3288# 0.031865f
C603 source.n207 a_n1724_n3288# 0.017123f
C604 source.n208 a_n1724_n3288# 0.01813f
C605 source.n209 a_n1724_n3288# 0.040472f
C606 source.n210 a_n1724_n3288# 0.083053f
C607 source.n211 a_n1724_n3288# 0.01813f
C608 source.n212 a_n1724_n3288# 0.017123f
C609 source.n213 a_n1724_n3288# 0.068431f
C610 source.n214 a_n1724_n3288# 0.045836f
C611 source.n215 a_n1724_n3288# 0.156158f
C612 source.t21 a_n1724_n3288# 0.302169f
C613 source.t27 a_n1724_n3288# 0.302169f
C614 source.n216 a_n1724_n3288# 2.58716f
C615 source.n217 a_n1724_n3288# 0.457681f
C616 source.t15 a_n1724_n3288# 0.302169f
C617 source.t18 a_n1724_n3288# 0.302169f
C618 source.n218 a_n1724_n3288# 2.58716f
C619 source.n219 a_n1724_n3288# 0.437323f
C620 source.t23 a_n1724_n3288# 0.302169f
C621 source.t24 a_n1724_n3288# 0.302169f
C622 source.n220 a_n1724_n3288# 2.58716f
C623 source.n221 a_n1724_n3288# 0.437323f
C624 source.n222 a_n1724_n3288# 0.042209f
C625 source.n223 a_n1724_n3288# 0.031865f
C626 source.n224 a_n1724_n3288# 0.017123f
C627 source.n225 a_n1724_n3288# 0.040472f
C628 source.n226 a_n1724_n3288# 0.01813f
C629 source.n227 a_n1724_n3288# 0.031865f
C630 source.n228 a_n1724_n3288# 0.017123f
C631 source.n229 a_n1724_n3288# 0.040472f
C632 source.n230 a_n1724_n3288# 0.01813f
C633 source.n231 a_n1724_n3288# 0.031865f
C634 source.n232 a_n1724_n3288# 0.017626f
C635 source.n233 a_n1724_n3288# 0.040472f
C636 source.n234 a_n1724_n3288# 0.01813f
C637 source.n235 a_n1724_n3288# 0.031865f
C638 source.n236 a_n1724_n3288# 0.017123f
C639 source.n237 a_n1724_n3288# 0.040472f
C640 source.n238 a_n1724_n3288# 0.01813f
C641 source.n239 a_n1724_n3288# 0.031865f
C642 source.n240 a_n1724_n3288# 0.017123f
C643 source.n241 a_n1724_n3288# 0.030354f
C644 source.n242 a_n1724_n3288# 0.028611f
C645 source.t25 a_n1724_n3288# 0.068355f
C646 source.n243 a_n1724_n3288# 0.229743f
C647 source.n244 a_n1724_n3288# 1.60754f
C648 source.n245 a_n1724_n3288# 0.017123f
C649 source.n246 a_n1724_n3288# 0.01813f
C650 source.n247 a_n1724_n3288# 0.040472f
C651 source.n248 a_n1724_n3288# 0.040472f
C652 source.n249 a_n1724_n3288# 0.01813f
C653 source.n250 a_n1724_n3288# 0.017123f
C654 source.n251 a_n1724_n3288# 0.031865f
C655 source.n252 a_n1724_n3288# 0.031865f
C656 source.n253 a_n1724_n3288# 0.017123f
C657 source.n254 a_n1724_n3288# 0.01813f
C658 source.n255 a_n1724_n3288# 0.040472f
C659 source.n256 a_n1724_n3288# 0.040472f
C660 source.n257 a_n1724_n3288# 0.01813f
C661 source.n258 a_n1724_n3288# 0.017123f
C662 source.n259 a_n1724_n3288# 0.031865f
C663 source.n260 a_n1724_n3288# 0.031865f
C664 source.n261 a_n1724_n3288# 0.017123f
C665 source.n262 a_n1724_n3288# 0.017123f
C666 source.n263 a_n1724_n3288# 0.01813f
C667 source.n264 a_n1724_n3288# 0.040472f
C668 source.n265 a_n1724_n3288# 0.040472f
C669 source.n266 a_n1724_n3288# 0.040472f
C670 source.n267 a_n1724_n3288# 0.017626f
C671 source.n268 a_n1724_n3288# 0.017123f
C672 source.n269 a_n1724_n3288# 0.031865f
C673 source.n270 a_n1724_n3288# 0.031865f
C674 source.n271 a_n1724_n3288# 0.017123f
C675 source.n272 a_n1724_n3288# 0.01813f
C676 source.n273 a_n1724_n3288# 0.040472f
C677 source.n274 a_n1724_n3288# 0.040472f
C678 source.n275 a_n1724_n3288# 0.01813f
C679 source.n276 a_n1724_n3288# 0.017123f
C680 source.n277 a_n1724_n3288# 0.031865f
C681 source.n278 a_n1724_n3288# 0.031865f
C682 source.n279 a_n1724_n3288# 0.017123f
C683 source.n280 a_n1724_n3288# 0.01813f
C684 source.n281 a_n1724_n3288# 0.040472f
C685 source.n282 a_n1724_n3288# 0.083053f
C686 source.n283 a_n1724_n3288# 0.01813f
C687 source.n284 a_n1724_n3288# 0.017123f
C688 source.n285 a_n1724_n3288# 0.068431f
C689 source.n286 a_n1724_n3288# 0.045836f
C690 source.n287 a_n1724_n3288# 0.308154f
C691 source.n288 a_n1724_n3288# 1.99902f
C692 minus.n0 a_n1724_n3288# 0.051385f
C693 minus.t4 a_n1724_n3288# 0.533536f
C694 minus.t2 a_n1724_n3288# 0.522735f
C695 minus.t12 a_n1724_n3288# 0.522735f
C696 minus.t7 a_n1724_n3288# 0.522735f
C697 minus.n1 a_n1724_n3288# 0.224412f
C698 minus.n2 a_n1724_n3288# 0.121063f
C699 minus.t3 a_n1724_n3288# 0.522735f
C700 minus.t13 a_n1724_n3288# 0.522735f
C701 minus.t8 a_n1724_n3288# 0.533536f
C702 minus.n3 a_n1724_n3288# 0.223831f
C703 minus.n4 a_n1724_n3288# 0.207366f
C704 minus.n5 a_n1724_n3288# 0.021164f
C705 minus.n6 a_n1724_n3288# 0.207366f
C706 minus.n7 a_n1724_n3288# 0.021164f
C707 minus.n8 a_n1724_n3288# 0.051385f
C708 minus.n9 a_n1724_n3288# 0.051385f
C709 minus.n10 a_n1724_n3288# 0.051385f
C710 minus.n11 a_n1724_n3288# 0.021164f
C711 minus.n12 a_n1724_n3288# 0.207366f
C712 minus.n13 a_n1724_n3288# 0.021164f
C713 minus.n14 a_n1724_n3288# 0.207366f
C714 minus.n15 a_n1724_n3288# 0.223749f
C715 minus.n16 a_n1724_n3288# 1.77782f
C716 minus.n17 a_n1724_n3288# 0.051385f
C717 minus.t11 a_n1724_n3288# 0.522735f
C718 minus.t6 a_n1724_n3288# 0.522735f
C719 minus.t9 a_n1724_n3288# 0.522735f
C720 minus.n18 a_n1724_n3288# 0.224412f
C721 minus.n19 a_n1724_n3288# 0.121063f
C722 minus.t0 a_n1724_n3288# 0.522735f
C723 minus.t10 a_n1724_n3288# 0.522735f
C724 minus.t1 a_n1724_n3288# 0.533536f
C725 minus.n20 a_n1724_n3288# 0.223831f
C726 minus.n21 a_n1724_n3288# 0.207366f
C727 minus.n22 a_n1724_n3288# 0.021164f
C728 minus.n23 a_n1724_n3288# 0.207366f
C729 minus.n24 a_n1724_n3288# 0.021164f
C730 minus.n25 a_n1724_n3288# 0.051385f
C731 minus.n26 a_n1724_n3288# 0.051385f
C732 minus.n27 a_n1724_n3288# 0.051385f
C733 minus.n28 a_n1724_n3288# 0.021164f
C734 minus.n29 a_n1724_n3288# 0.207366f
C735 minus.n30 a_n1724_n3288# 0.021164f
C736 minus.n31 a_n1724_n3288# 0.207366f
C737 minus.t5 a_n1724_n3288# 0.533536f
C738 minus.n32 a_n1724_n3288# 0.223749f
C739 minus.n33 a_n1724_n3288# 0.340349f
C740 minus.n34 a_n1724_n3288# 2.16117f
.ends

