* NGSPICE file created from diffpair404.ext - technology: sky130A

.subckt diffpair404 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t9 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X1 drain_left.t9 plus.t0 source.t2 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X2 a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X3 a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X4 source.t4 plus.t1 drain_left.t8 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X5 drain_right.t8 minus.t1 source.t16 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X6 drain_left.t7 plus.t2 source.t5 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X7 source.t8 minus.t2 drain_right.t7 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X8 a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X9 drain_left.t6 plus.t3 source.t0 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X10 drain_right.t6 minus.t3 source.t10 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X11 drain_right.t5 minus.t4 source.t13 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X12 source.t14 minus.t5 drain_right.t4 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 source.t12 minus.t6 drain_right.t3 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X14 source.t1 plus.t4 drain_left.t5 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X15 drain_left.t4 plus.t5 source.t6 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X16 drain_right.t2 minus.t7 source.t11 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 source.t17 plus.t6 drain_left.t3 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X18 drain_right.t1 minus.t8 source.t15 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 drain_left.t2 plus.t7 source.t18 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X20 a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X21 source.t19 plus.t8 drain_left.t1 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X22 drain_left.t0 plus.t9 source.t3 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X23 source.t7 minus.t9 drain_right.t0 a_n1496_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
R0 minus.n9 minus.t4 2180.68
R1 minus.n3 minus.t3 2180.68
R2 minus.n20 minus.t1 2180.68
R3 minus.n14 minus.t0 2180.68
R4 minus.n6 minus.t7 2136.87
R5 minus.n8 minus.t6 2136.87
R6 minus.n2 minus.t2 2136.87
R7 minus.n17 minus.t8 2136.87
R8 minus.n19 minus.t9 2136.87
R9 minus.n13 minus.t5 2136.87
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 34.8016
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 source.n5 source.t10 45.3739
R42 source.n19 source.t16 45.3737
R43 source.n14 source.t5 45.3737
R44 source.n0 source.t3 45.3737
R45 source.n2 source.n1 42.8739
R46 source.n4 source.n3 42.8739
R47 source.n7 source.n6 42.8739
R48 source.n9 source.n8 42.8739
R49 source.n18 source.n17 42.8737
R50 source.n16 source.n15 42.8737
R51 source.n13 source.n12 42.8737
R52 source.n11 source.n10 42.8737
R53 source.n11 source.n9 22.4084
R54 source.n20 source.n0 16.305
R55 source.n20 source.n19 5.5436
R56 source.n17 source.t15 2.5005
R57 source.n17 source.t7 2.5005
R58 source.n15 source.t9 2.5005
R59 source.n15 source.t14 2.5005
R60 source.n12 source.t2 2.5005
R61 source.n12 source.t1 2.5005
R62 source.n10 source.t0 2.5005
R63 source.n10 source.t4 2.5005
R64 source.n1 source.t18 2.5005
R65 source.n1 source.t17 2.5005
R66 source.n3 source.t6 2.5005
R67 source.n3 source.t19 2.5005
R68 source.n6 source.t11 2.5005
R69 source.n6 source.t8 2.5005
R70 source.n8 source.t13 2.5005
R71 source.n8 source.t12 2.5005
R72 source.n5 source.n4 0.7505
R73 source.n16 source.n14 0.7505
R74 source.n9 source.n7 0.560845
R75 source.n7 source.n5 0.560845
R76 source.n4 source.n2 0.560845
R77 source.n2 source.n0 0.560845
R78 source.n13 source.n11 0.560845
R79 source.n14 source.n13 0.560845
R80 source.n18 source.n16 0.560845
R81 source.n19 source.n18 0.560845
R82 source source.n20 0.188
R83 drain_right.n1 drain_right.t9 62.6128
R84 drain_right.n7 drain_right.t5 62.0527
R85 drain_right.n6 drain_right.n4 60.1128
R86 drain_right.n3 drain_right.n2 59.9174
R87 drain_right.n6 drain_right.n5 59.5527
R88 drain_right.n1 drain_right.n0 59.5525
R89 drain_right drain_right.n3 29.1953
R90 drain_right drain_right.n7 5.93339
R91 drain_right.n2 drain_right.t0 2.5005
R92 drain_right.n2 drain_right.t8 2.5005
R93 drain_right.n0 drain_right.t4 2.5005
R94 drain_right.n0 drain_right.t1 2.5005
R95 drain_right.n4 drain_right.t7 2.5005
R96 drain_right.n4 drain_right.t6 2.5005
R97 drain_right.n5 drain_right.t3 2.5005
R98 drain_right.n5 drain_right.t2 2.5005
R99 drain_right.n7 drain_right.n6 0.560845
R100 drain_right.n3 drain_right.n1 0.0852402
R101 plus.n3 plus.t5 2180.68
R102 plus.n9 plus.t9 2180.68
R103 plus.n14 plus.t2 2180.68
R104 plus.n20 plus.t3 2180.68
R105 plus.n6 plus.t7 2136.87
R106 plus.n2 plus.t8 2136.87
R107 plus.n8 plus.t6 2136.87
R108 plus.n17 plus.t0 2136.87
R109 plus.n13 plus.t4 2136.87
R110 plus.n19 plus.t1 2136.87
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 28.6827
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 12.1577
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t4 62.613
R142 drain_left.n1 drain_left.t6 62.6128
R143 drain_left.n3 drain_left.n2 59.9174
R144 drain_left.n5 drain_left.n4 59.5527
R145 drain_left.n1 drain_left.n0 59.5525
R146 drain_left.n7 drain_left.n6 59.5525
R147 drain_left drain_left.n3 29.7485
R148 drain_left drain_left.n7 6.21356
R149 drain_left.n2 drain_left.t5 2.5005
R150 drain_left.n2 drain_left.t7 2.5005
R151 drain_left.n0 drain_left.t8 2.5005
R152 drain_left.n0 drain_left.t9 2.5005
R153 drain_left.n6 drain_left.t3 2.5005
R154 drain_left.n6 drain_left.t0 2.5005
R155 drain_left.n4 drain_left.t1 2.5005
R156 drain_left.n4 drain_left.t2 2.5005
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 minus drain_left 0.170828f
C1 drain_right drain_left 0.736455f
C2 source minus 1.98579f
C3 drain_right source 21.4566f
C4 plus drain_left 2.65644f
C5 drain_right minus 2.51628f
C6 source plus 2.00047f
C7 plus minus 5.00348f
C8 drain_right plus 0.298633f
C9 source drain_left 21.467402f
C10 drain_right a_n1496_n3288# 6.5503f
C11 drain_left a_n1496_n3288# 6.79411f
C12 source a_n1496_n3288# 6.15247f
C13 minus a_n1496_n3288# 5.492365f
C14 plus a_n1496_n3288# 7.6745f
C15 drain_left.t6 a_n1496_n3288# 2.95863f
C16 drain_left.t8 a_n1496_n3288# 0.366804f
C17 drain_left.t9 a_n1496_n3288# 0.366804f
C18 drain_left.n0 a_n1496_n3288# 2.40366f
C19 drain_left.n1 a_n1496_n3288# 0.650212f
C20 drain_left.t5 a_n1496_n3288# 0.366804f
C21 drain_left.t7 a_n1496_n3288# 0.366804f
C22 drain_left.n2 a_n1496_n3288# 2.4055f
C23 drain_left.n3 a_n1496_n3288# 1.45584f
C24 drain_left.t4 a_n1496_n3288# 2.95864f
C25 drain_left.t1 a_n1496_n3288# 0.366804f
C26 drain_left.t2 a_n1496_n3288# 0.366804f
C27 drain_left.n4 a_n1496_n3288# 2.40367f
C28 drain_left.n5 a_n1496_n3288# 0.682334f
C29 drain_left.t3 a_n1496_n3288# 0.366804f
C30 drain_left.t0 a_n1496_n3288# 0.366804f
C31 drain_left.n6 a_n1496_n3288# 2.40366f
C32 drain_left.n7 a_n1496_n3288# 0.519646f
C33 plus.n0 a_n1496_n3288# 0.059225f
C34 plus.t6 a_n1496_n3288# 0.301248f
C35 plus.t7 a_n1496_n3288# 0.301248f
C36 plus.n1 a_n1496_n3288# 0.025124f
C37 plus.t5 a_n1496_n3288# 0.303796f
C38 plus.t8 a_n1496_n3288# 0.301248f
C39 plus.n2 a_n1496_n3288# 0.128632f
C40 plus.n3 a_n1496_n3288# 0.149463f
C41 plus.n4 a_n1496_n3288# 0.127499f
C42 plus.n5 a_n1496_n3288# 0.059225f
C43 plus.n6 a_n1496_n3288# 0.148279f
C44 plus.n7 a_n1496_n3288# 0.025124f
C45 plus.n8 a_n1496_n3288# 0.128632f
C46 plus.t9 a_n1496_n3288# 0.303796f
C47 plus.n9 a_n1496_n3288# 0.149383f
C48 plus.n10 a_n1496_n3288# 0.664588f
C49 plus.n11 a_n1496_n3288# 0.059225f
C50 plus.t3 a_n1496_n3288# 0.303796f
C51 plus.t1 a_n1496_n3288# 0.301248f
C52 plus.t0 a_n1496_n3288# 0.301248f
C53 plus.n12 a_n1496_n3288# 0.025124f
C54 plus.t4 a_n1496_n3288# 0.301248f
C55 plus.n13 a_n1496_n3288# 0.128632f
C56 plus.t2 a_n1496_n3288# 0.303796f
C57 plus.n14 a_n1496_n3288# 0.149463f
C58 plus.n15 a_n1496_n3288# 0.127499f
C59 plus.n16 a_n1496_n3288# 0.059225f
C60 plus.n17 a_n1496_n3288# 0.148279f
C61 plus.n18 a_n1496_n3288# 0.025124f
C62 plus.n19 a_n1496_n3288# 0.128632f
C63 plus.n20 a_n1496_n3288# 0.149383f
C64 plus.n21 a_n1496_n3288# 1.66022f
C65 drain_right.t9 a_n1496_n3288# 2.94634f
C66 drain_right.t4 a_n1496_n3288# 0.36528f
C67 drain_right.t1 a_n1496_n3288# 0.36528f
C68 drain_right.n0 a_n1496_n3288# 2.39367f
C69 drain_right.n1 a_n1496_n3288# 0.647511f
C70 drain_right.t0 a_n1496_n3288# 0.36528f
C71 drain_right.t8 a_n1496_n3288# 0.36528f
C72 drain_right.n2 a_n1496_n3288# 2.3955f
C73 drain_right.n3 a_n1496_n3288# 1.39672f
C74 drain_right.t7 a_n1496_n3288# 0.36528f
C75 drain_right.t6 a_n1496_n3288# 0.36528f
C76 drain_right.n4 a_n1496_n3288# 2.39661f
C77 drain_right.t3 a_n1496_n3288# 0.36528f
C78 drain_right.t2 a_n1496_n3288# 0.36528f
C79 drain_right.n5 a_n1496_n3288# 2.39368f
C80 drain_right.n6 a_n1496_n3288# 0.61764f
C81 drain_right.t5 a_n1496_n3288# 2.94297f
C82 drain_right.n7 a_n1496_n3288# 0.590896f
C83 source.t3 a_n1496_n3288# 2.76996f
C84 source.n0 a_n1496_n3288# 1.38136f
C85 source.t18 a_n1496_n3288# 0.357968f
C86 source.t17 a_n1496_n3288# 0.357968f
C87 source.n1 a_n1496_n3288# 2.26627f
C88 source.n2 a_n1496_n3288# 0.344689f
C89 source.t6 a_n1496_n3288# 0.357968f
C90 source.t19 a_n1496_n3288# 0.357968f
C91 source.n3 a_n1496_n3288# 2.26627f
C92 source.n4 a_n1496_n3288# 0.359915f
C93 source.t10 a_n1496_n3288# 2.76997f
C94 source.n5 a_n1496_n3288# 0.500561f
C95 source.t11 a_n1496_n3288# 0.357968f
C96 source.t8 a_n1496_n3288# 0.357968f
C97 source.n6 a_n1496_n3288# 2.26627f
C98 source.n7 a_n1496_n3288# 0.344689f
C99 source.t13 a_n1496_n3288# 0.357968f
C100 source.t12 a_n1496_n3288# 0.357968f
C101 source.n8 a_n1496_n3288# 2.26627f
C102 source.n9 a_n1496_n3288# 1.67794f
C103 source.t0 a_n1496_n3288# 0.357968f
C104 source.t4 a_n1496_n3288# 0.357968f
C105 source.n10 a_n1496_n3288# 2.26626f
C106 source.n11 a_n1496_n3288# 1.67795f
C107 source.t2 a_n1496_n3288# 0.357968f
C108 source.t1 a_n1496_n3288# 0.357968f
C109 source.n12 a_n1496_n3288# 2.26626f
C110 source.n13 a_n1496_n3288# 0.344701f
C111 source.t5 a_n1496_n3288# 2.76996f
C112 source.n14 a_n1496_n3288# 0.500573f
C113 source.t9 a_n1496_n3288# 0.357968f
C114 source.t14 a_n1496_n3288# 0.357968f
C115 source.n15 a_n1496_n3288# 2.26626f
C116 source.n16 a_n1496_n3288# 0.359927f
C117 source.t15 a_n1496_n3288# 0.357968f
C118 source.t7 a_n1496_n3288# 0.357968f
C119 source.n17 a_n1496_n3288# 2.26626f
C120 source.n18 a_n1496_n3288# 0.344701f
C121 source.t16 a_n1496_n3288# 2.76996f
C122 source.n19 a_n1496_n3288# 0.619829f
C123 source.n20 a_n1496_n3288# 1.56377f
C124 minus.n0 a_n1496_n3288# 0.045234f
C125 minus.t4 a_n1496_n3288# 0.232029f
C126 minus.t6 a_n1496_n3288# 0.230083f
C127 minus.t7 a_n1496_n3288# 0.230083f
C128 minus.n1 a_n1496_n3288# 0.019189f
C129 minus.t2 a_n1496_n3288# 0.230083f
C130 minus.n2 a_n1496_n3288# 0.098245f
C131 minus.t3 a_n1496_n3288# 0.232029f
C132 minus.n3 a_n1496_n3288# 0.114154f
C133 minus.n4 a_n1496_n3288# 0.097379f
C134 minus.n5 a_n1496_n3288# 0.045234f
C135 minus.n6 a_n1496_n3288# 0.11325f
C136 minus.n7 a_n1496_n3288# 0.019189f
C137 minus.n8 a_n1496_n3288# 0.098245f
C138 minus.n9 a_n1496_n3288# 0.114093f
C139 minus.n10 a_n1496_n3288# 1.50324f
C140 minus.n11 a_n1496_n3288# 0.045234f
C141 minus.t9 a_n1496_n3288# 0.230083f
C142 minus.t8 a_n1496_n3288# 0.230083f
C143 minus.n12 a_n1496_n3288# 0.019189f
C144 minus.t0 a_n1496_n3288# 0.232029f
C145 minus.t5 a_n1496_n3288# 0.230083f
C146 minus.n13 a_n1496_n3288# 0.098245f
C147 minus.n14 a_n1496_n3288# 0.114154f
C148 minus.n15 a_n1496_n3288# 0.097379f
C149 minus.n16 a_n1496_n3288# 0.045234f
C150 minus.n17 a_n1496_n3288# 0.11325f
C151 minus.n18 a_n1496_n3288# 0.019189f
C152 minus.n19 a_n1496_n3288# 0.098245f
C153 minus.t1 a_n1496_n3288# 0.232029f
C154 minus.n20 a_n1496_n3288# 0.114093f
C155 minus.n21 a_n1496_n3288# 0.297195f
C156 minus.n22 a_n1496_n3288# 1.83282f
.ends

