* NGSPICE file created from diffpair628.ext - technology: sky130A

.subckt diffpair628 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t22 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 source.t15 minus.t0 drain_right.t19 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X2 source.t26 plus.t1 drain_left.t18 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t33 plus.t2 drain_left.t17 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 drain_right.t18 minus.t1 source.t3 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X5 source.t31 plus.t3 drain_left.t16 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 source.t7 minus.t2 drain_right.t17 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X8 drain_left.t15 plus.t4 source.t21 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X9 source.t8 minus.t3 drain_right.t16 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X10 source.t28 plus.t5 drain_left.t14 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X11 source.t36 plus.t6 drain_left.t13 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X12 source.t38 plus.t7 drain_left.t12 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X13 drain_left.t11 plus.t8 source.t24 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X14 drain_right.t15 minus.t4 source.t1 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X15 source.t9 minus.t5 drain_right.t14 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X16 drain_right.t13 minus.t6 source.t10 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X17 a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X18 drain_right.t12 minus.t7 source.t18 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 drain_right.t11 minus.t8 source.t19 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X20 drain_right.t10 minus.t9 source.t4 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X21 drain_left.t10 plus.t9 source.t32 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X22 drain_right.t9 minus.t10 source.t12 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 drain_left.t9 plus.t10 source.t39 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X24 drain_left.t8 plus.t11 source.t35 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X25 source.t23 plus.t12 drain_left.t7 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X26 drain_left.t6 plus.t13 source.t27 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X27 drain_right.t8 minus.t11 source.t5 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X28 drain_left.t5 plus.t14 source.t34 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X29 a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X30 drain_right.t7 minus.t12 source.t2 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X31 a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X32 source.t6 minus.t13 drain_right.t6 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X33 source.t16 minus.t14 drain_right.t5 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X34 drain_left.t4 plus.t15 source.t37 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X35 source.t25 plus.t16 drain_left.t3 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X36 drain_left.t2 plus.t17 source.t30 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X37 source.t0 minus.t15 drain_right.t4 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X38 drain_right.t3 minus.t16 source.t14 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X39 source.t11 minus.t17 drain_right.t2 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X40 source.t17 minus.t18 drain_right.t1 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X41 source.t13 minus.t19 drain_right.t0 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X42 source.t29 plus.t18 drain_left.t1 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X43 source.t20 plus.t19 drain_left.t0 a_n2982_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n9 plus.t6 770.083
R1 plus.n43 plus.t0 770.083
R2 plus.n32 plus.t4 744.691
R3 plus.n30 plus.t18 744.691
R4 plus.n2 plus.t9 744.691
R5 plus.n24 plus.t2 744.691
R6 plus.n4 plus.t11 744.691
R7 plus.n18 plus.t5 744.691
R8 plus.n6 plus.t10 744.691
R9 plus.n12 plus.t3 744.691
R10 plus.n8 plus.t14 744.691
R11 plus.n66 plus.t16 744.691
R12 plus.n64 plus.t15 744.691
R13 plus.n36 plus.t19 744.691
R14 plus.n58 plus.t8 744.691
R15 plus.n38 plus.t7 744.691
R16 plus.n52 plus.t13 744.691
R17 plus.n40 plus.t12 744.691
R18 plus.n46 plus.t17 744.691
R19 plus.n42 plus.t1 744.691
R20 plus.n11 plus.n10 161.3
R21 plus.n12 plus.n7 161.3
R22 plus.n14 plus.n13 161.3
R23 plus.n15 plus.n6 161.3
R24 plus.n17 plus.n16 161.3
R25 plus.n18 plus.n5 161.3
R26 plus.n20 plus.n19 161.3
R27 plus.n21 plus.n4 161.3
R28 plus.n23 plus.n22 161.3
R29 plus.n24 plus.n3 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n27 plus.n2 161.3
R32 plus.n29 plus.n28 161.3
R33 plus.n30 plus.n1 161.3
R34 plus.n31 plus.n0 161.3
R35 plus.n33 plus.n32 161.3
R36 plus.n45 plus.n44 161.3
R37 plus.n46 plus.n41 161.3
R38 plus.n48 plus.n47 161.3
R39 plus.n49 plus.n40 161.3
R40 plus.n51 plus.n50 161.3
R41 plus.n52 plus.n39 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n55 plus.n38 161.3
R44 plus.n57 plus.n56 161.3
R45 plus.n58 plus.n37 161.3
R46 plus.n60 plus.n59 161.3
R47 plus.n61 plus.n36 161.3
R48 plus.n63 plus.n62 161.3
R49 plus.n64 plus.n35 161.3
R50 plus.n65 plus.n34 161.3
R51 plus.n67 plus.n66 161.3
R52 plus.n10 plus.n9 45.0031
R53 plus.n44 plus.n43 45.0031
R54 plus.n32 plus.n31 41.6278
R55 plus.n66 plus.n65 41.6278
R56 plus plus.n67 37.4952
R57 plus.n30 plus.n29 37.246
R58 plus.n11 plus.n8 37.246
R59 plus.n64 plus.n63 37.246
R60 plus.n45 plus.n42 37.246
R61 plus.n25 plus.n2 32.8641
R62 plus.n13 plus.n12 32.8641
R63 plus.n59 plus.n36 32.8641
R64 plus.n47 plus.n46 32.8641
R65 plus.n24 plus.n23 28.4823
R66 plus.n17 plus.n6 28.4823
R67 plus.n58 plus.n57 28.4823
R68 plus.n51 plus.n40 28.4823
R69 plus.n19 plus.n18 24.1005
R70 plus.n19 plus.n4 24.1005
R71 plus.n53 plus.n38 24.1005
R72 plus.n53 plus.n52 24.1005
R73 plus.n23 plus.n4 19.7187
R74 plus.n18 plus.n17 19.7187
R75 plus.n57 plus.n38 19.7187
R76 plus.n52 plus.n51 19.7187
R77 plus.n9 plus.n8 15.6319
R78 plus.n43 plus.n42 15.6319
R79 plus plus.n33 15.3414
R80 plus.n25 plus.n24 15.3369
R81 plus.n13 plus.n6 15.3369
R82 plus.n59 plus.n58 15.3369
R83 plus.n47 plus.n40 15.3369
R84 plus.n29 plus.n2 10.955
R85 plus.n12 plus.n11 10.955
R86 plus.n63 plus.n36 10.955
R87 plus.n46 plus.n45 10.955
R88 plus.n31 plus.n30 6.57323
R89 plus.n65 plus.n64 6.57323
R90 plus.n10 plus.n7 0.189894
R91 plus.n14 plus.n7 0.189894
R92 plus.n15 plus.n14 0.189894
R93 plus.n16 plus.n15 0.189894
R94 plus.n16 plus.n5 0.189894
R95 plus.n20 plus.n5 0.189894
R96 plus.n21 plus.n20 0.189894
R97 plus.n22 plus.n21 0.189894
R98 plus.n22 plus.n3 0.189894
R99 plus.n26 plus.n3 0.189894
R100 plus.n27 plus.n26 0.189894
R101 plus.n28 plus.n27 0.189894
R102 plus.n28 plus.n1 0.189894
R103 plus.n1 plus.n0 0.189894
R104 plus.n33 plus.n0 0.189894
R105 plus.n67 plus.n34 0.189894
R106 plus.n35 plus.n34 0.189894
R107 plus.n62 plus.n35 0.189894
R108 plus.n62 plus.n61 0.189894
R109 plus.n61 plus.n60 0.189894
R110 plus.n60 plus.n37 0.189894
R111 plus.n56 plus.n37 0.189894
R112 plus.n56 plus.n55 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n39 0.189894
R115 plus.n50 plus.n39 0.189894
R116 plus.n50 plus.n49 0.189894
R117 plus.n49 plus.n48 0.189894
R118 plus.n48 plus.n41 0.189894
R119 plus.n44 plus.n41 0.189894
R120 source.n0 source.t21 44.1297
R121 source.n9 source.t36 44.1296
R122 source.n10 source.t5 44.1296
R123 source.n19 source.t6 44.1296
R124 source.n39 source.t19 44.1295
R125 source.n30 source.t9 44.1295
R126 source.n29 source.t22 44.1295
R127 source.n20 source.t25 44.1295
R128 source.n2 source.n1 43.1397
R129 source.n4 source.n3 43.1397
R130 source.n6 source.n5 43.1397
R131 source.n8 source.n7 43.1397
R132 source.n12 source.n11 43.1397
R133 source.n14 source.n13 43.1397
R134 source.n16 source.n15 43.1397
R135 source.n18 source.n17 43.1397
R136 source.n38 source.n37 43.1396
R137 source.n36 source.n35 43.1396
R138 source.n34 source.n33 43.1396
R139 source.n32 source.n31 43.1396
R140 source.n28 source.n27 43.1396
R141 source.n26 source.n25 43.1396
R142 source.n24 source.n23 43.1396
R143 source.n22 source.n21 43.1396
R144 source.n20 source.n19 28.2363
R145 source.n40 source.n0 22.5294
R146 source.n40 source.n39 5.7074
R147 source.n37 source.t2 0.9905
R148 source.n37 source.t16 0.9905
R149 source.n35 source.t14 0.9905
R150 source.n35 source.t13 0.9905
R151 source.n33 source.t3 0.9905
R152 source.n33 source.t8 0.9905
R153 source.n31 source.t1 0.9905
R154 source.n31 source.t15 0.9905
R155 source.n27 source.t30 0.9905
R156 source.n27 source.t26 0.9905
R157 source.n25 source.t27 0.9905
R158 source.n25 source.t23 0.9905
R159 source.n23 source.t24 0.9905
R160 source.n23 source.t38 0.9905
R161 source.n21 source.t37 0.9905
R162 source.n21 source.t20 0.9905
R163 source.n1 source.t32 0.9905
R164 source.n1 source.t29 0.9905
R165 source.n3 source.t35 0.9905
R166 source.n3 source.t33 0.9905
R167 source.n5 source.t39 0.9905
R168 source.n5 source.t28 0.9905
R169 source.n7 source.t34 0.9905
R170 source.n7 source.t31 0.9905
R171 source.n11 source.t12 0.9905
R172 source.n11 source.t7 0.9905
R173 source.n13 source.t4 0.9905
R174 source.n13 source.t11 0.9905
R175 source.n15 source.t18 0.9905
R176 source.n15 source.t17 0.9905
R177 source.n17 source.t10 0.9905
R178 source.n17 source.t0 0.9905
R179 source.n19 source.n18 0.888431
R180 source.n18 source.n16 0.888431
R181 source.n16 source.n14 0.888431
R182 source.n14 source.n12 0.888431
R183 source.n12 source.n10 0.888431
R184 source.n9 source.n8 0.888431
R185 source.n8 source.n6 0.888431
R186 source.n6 source.n4 0.888431
R187 source.n4 source.n2 0.888431
R188 source.n2 source.n0 0.888431
R189 source.n22 source.n20 0.888431
R190 source.n24 source.n22 0.888431
R191 source.n26 source.n24 0.888431
R192 source.n28 source.n26 0.888431
R193 source.n29 source.n28 0.888431
R194 source.n32 source.n30 0.888431
R195 source.n34 source.n32 0.888431
R196 source.n36 source.n34 0.888431
R197 source.n38 source.n36 0.888431
R198 source.n39 source.n38 0.888431
R199 source.n10 source.n9 0.470328
R200 source.n30 source.n29 0.470328
R201 source source.n40 0.188
R202 drain_left.n10 drain_left.n8 60.7064
R203 drain_left.n6 drain_left.n4 60.7063
R204 drain_left.n2 drain_left.n0 60.7063
R205 drain_left.n16 drain_left.n15 59.8185
R206 drain_left.n14 drain_left.n13 59.8185
R207 drain_left.n12 drain_left.n11 59.8185
R208 drain_left.n10 drain_left.n9 59.8185
R209 drain_left.n7 drain_left.n3 59.8184
R210 drain_left.n6 drain_left.n5 59.8184
R211 drain_left.n2 drain_left.n1 59.8184
R212 drain_left drain_left.n7 40.5311
R213 drain_left drain_left.n16 6.54115
R214 drain_left.n3 drain_left.t12 0.9905
R215 drain_left.n3 drain_left.t6 0.9905
R216 drain_left.n4 drain_left.t18 0.9905
R217 drain_left.n4 drain_left.t19 0.9905
R218 drain_left.n5 drain_left.t7 0.9905
R219 drain_left.n5 drain_left.t2 0.9905
R220 drain_left.n1 drain_left.t0 0.9905
R221 drain_left.n1 drain_left.t11 0.9905
R222 drain_left.n0 drain_left.t3 0.9905
R223 drain_left.n0 drain_left.t4 0.9905
R224 drain_left.n15 drain_left.t1 0.9905
R225 drain_left.n15 drain_left.t15 0.9905
R226 drain_left.n13 drain_left.t17 0.9905
R227 drain_left.n13 drain_left.t10 0.9905
R228 drain_left.n11 drain_left.t14 0.9905
R229 drain_left.n11 drain_left.t8 0.9905
R230 drain_left.n9 drain_left.t16 0.9905
R231 drain_left.n9 drain_left.t9 0.9905
R232 drain_left.n8 drain_left.t13 0.9905
R233 drain_left.n8 drain_left.t5 0.9905
R234 drain_left.n12 drain_left.n10 0.888431
R235 drain_left.n14 drain_left.n12 0.888431
R236 drain_left.n16 drain_left.n14 0.888431
R237 drain_left.n7 drain_left.n6 0.833085
R238 drain_left.n7 drain_left.n2 0.833085
R239 minus.n9 minus.t11 770.083
R240 minus.n43 minus.t5 770.083
R241 minus.n8 minus.t2 744.691
R242 minus.n12 minus.t10 744.691
R243 minus.n14 minus.t17 744.691
R244 minus.n18 minus.t9 744.691
R245 minus.n20 minus.t18 744.691
R246 minus.n24 minus.t7 744.691
R247 minus.n26 minus.t15 744.691
R248 minus.n30 minus.t6 744.691
R249 minus.n32 minus.t13 744.691
R250 minus.n42 minus.t4 744.691
R251 minus.n46 minus.t0 744.691
R252 minus.n48 minus.t1 744.691
R253 minus.n52 minus.t3 744.691
R254 minus.n54 minus.t16 744.691
R255 minus.n58 minus.t19 744.691
R256 minus.n60 minus.t12 744.691
R257 minus.n64 minus.t14 744.691
R258 minus.n66 minus.t8 744.691
R259 minus.n33 minus.n32 161.3
R260 minus.n31 minus.n0 161.3
R261 minus.n30 minus.n29 161.3
R262 minus.n28 minus.n1 161.3
R263 minus.n27 minus.n26 161.3
R264 minus.n25 minus.n2 161.3
R265 minus.n24 minus.n23 161.3
R266 minus.n22 minus.n3 161.3
R267 minus.n21 minus.n20 161.3
R268 minus.n19 minus.n4 161.3
R269 minus.n18 minus.n17 161.3
R270 minus.n16 minus.n5 161.3
R271 minus.n15 minus.n14 161.3
R272 minus.n13 minus.n6 161.3
R273 minus.n12 minus.n11 161.3
R274 minus.n10 minus.n7 161.3
R275 minus.n67 minus.n66 161.3
R276 minus.n65 minus.n34 161.3
R277 minus.n64 minus.n63 161.3
R278 minus.n62 minus.n35 161.3
R279 minus.n61 minus.n60 161.3
R280 minus.n59 minus.n36 161.3
R281 minus.n58 minus.n57 161.3
R282 minus.n56 minus.n37 161.3
R283 minus.n55 minus.n54 161.3
R284 minus.n53 minus.n38 161.3
R285 minus.n52 minus.n51 161.3
R286 minus.n50 minus.n39 161.3
R287 minus.n49 minus.n48 161.3
R288 minus.n47 minus.n40 161.3
R289 minus.n46 minus.n45 161.3
R290 minus.n44 minus.n41 161.3
R291 minus.n68 minus.n33 46.6444
R292 minus.n10 minus.n9 45.0031
R293 minus.n44 minus.n43 45.0031
R294 minus.n32 minus.n31 41.6278
R295 minus.n66 minus.n65 41.6278
R296 minus.n8 minus.n7 37.246
R297 minus.n30 minus.n1 37.246
R298 minus.n42 minus.n41 37.246
R299 minus.n64 minus.n35 37.246
R300 minus.n13 minus.n12 32.8641
R301 minus.n26 minus.n25 32.8641
R302 minus.n47 minus.n46 32.8641
R303 minus.n60 minus.n59 32.8641
R304 minus.n14 minus.n5 28.4823
R305 minus.n24 minus.n3 28.4823
R306 minus.n48 minus.n39 28.4823
R307 minus.n58 minus.n37 28.4823
R308 minus.n20 minus.n19 24.1005
R309 minus.n19 minus.n18 24.1005
R310 minus.n53 minus.n52 24.1005
R311 minus.n54 minus.n53 24.1005
R312 minus.n18 minus.n5 19.7187
R313 minus.n20 minus.n3 19.7187
R314 minus.n52 minus.n39 19.7187
R315 minus.n54 minus.n37 19.7187
R316 minus.n9 minus.n8 15.6319
R317 minus.n43 minus.n42 15.6319
R318 minus.n14 minus.n13 15.3369
R319 minus.n25 minus.n24 15.3369
R320 minus.n48 minus.n47 15.3369
R321 minus.n59 minus.n58 15.3369
R322 minus.n12 minus.n7 10.955
R323 minus.n26 minus.n1 10.955
R324 minus.n46 minus.n41 10.955
R325 minus.n60 minus.n35 10.955
R326 minus.n68 minus.n67 6.66717
R327 minus.n31 minus.n30 6.57323
R328 minus.n65 minus.n64 6.57323
R329 minus.n33 minus.n0 0.189894
R330 minus.n29 minus.n0 0.189894
R331 minus.n29 minus.n28 0.189894
R332 minus.n28 minus.n27 0.189894
R333 minus.n27 minus.n2 0.189894
R334 minus.n23 minus.n2 0.189894
R335 minus.n23 minus.n22 0.189894
R336 minus.n22 minus.n21 0.189894
R337 minus.n21 minus.n4 0.189894
R338 minus.n17 minus.n4 0.189894
R339 minus.n17 minus.n16 0.189894
R340 minus.n16 minus.n15 0.189894
R341 minus.n15 minus.n6 0.189894
R342 minus.n11 minus.n6 0.189894
R343 minus.n11 minus.n10 0.189894
R344 minus.n45 minus.n44 0.189894
R345 minus.n45 minus.n40 0.189894
R346 minus.n49 minus.n40 0.189894
R347 minus.n50 minus.n49 0.189894
R348 minus.n51 minus.n50 0.189894
R349 minus.n51 minus.n38 0.189894
R350 minus.n55 minus.n38 0.189894
R351 minus.n56 minus.n55 0.189894
R352 minus.n57 minus.n56 0.189894
R353 minus.n57 minus.n36 0.189894
R354 minus.n61 minus.n36 0.189894
R355 minus.n62 minus.n61 0.189894
R356 minus.n63 minus.n62 0.189894
R357 minus.n63 minus.n34 0.189894
R358 minus.n67 minus.n34 0.189894
R359 minus minus.n68 0.188
R360 drain_right.n10 drain_right.n8 60.7064
R361 drain_right.n6 drain_right.n4 60.7063
R362 drain_right.n2 drain_right.n0 60.7063
R363 drain_right.n10 drain_right.n9 59.8185
R364 drain_right.n12 drain_right.n11 59.8185
R365 drain_right.n14 drain_right.n13 59.8185
R366 drain_right.n16 drain_right.n15 59.8185
R367 drain_right.n7 drain_right.n3 59.8184
R368 drain_right.n6 drain_right.n5 59.8184
R369 drain_right.n2 drain_right.n1 59.8184
R370 drain_right drain_right.n7 39.9779
R371 drain_right drain_right.n16 6.54115
R372 drain_right.n3 drain_right.t16 0.9905
R373 drain_right.n3 drain_right.t3 0.9905
R374 drain_right.n4 drain_right.t5 0.9905
R375 drain_right.n4 drain_right.t11 0.9905
R376 drain_right.n5 drain_right.t0 0.9905
R377 drain_right.n5 drain_right.t7 0.9905
R378 drain_right.n1 drain_right.t19 0.9905
R379 drain_right.n1 drain_right.t18 0.9905
R380 drain_right.n0 drain_right.t14 0.9905
R381 drain_right.n0 drain_right.t15 0.9905
R382 drain_right.n8 drain_right.t17 0.9905
R383 drain_right.n8 drain_right.t8 0.9905
R384 drain_right.n9 drain_right.t2 0.9905
R385 drain_right.n9 drain_right.t9 0.9905
R386 drain_right.n11 drain_right.t1 0.9905
R387 drain_right.n11 drain_right.t10 0.9905
R388 drain_right.n13 drain_right.t4 0.9905
R389 drain_right.n13 drain_right.t12 0.9905
R390 drain_right.n15 drain_right.t6 0.9905
R391 drain_right.n15 drain_right.t13 0.9905
R392 drain_right.n16 drain_right.n14 0.888431
R393 drain_right.n14 drain_right.n12 0.888431
R394 drain_right.n12 drain_right.n10 0.888431
R395 drain_right.n7 drain_right.n6 0.833085
R396 drain_right.n7 drain_right.n2 0.833085
C0 drain_left drain_right 1.59885f
C1 plus drain_right 0.454687f
C2 plus drain_left 20.8236f
C3 source minus 20.3715f
C4 minus drain_right 20.5261f
C5 drain_left minus 0.173554f
C6 plus minus 8.34701f
C7 source drain_right 37.3771f
C8 source drain_left 37.3748f
C9 plus source 20.3856f
C10 drain_right a_n2982_n4888# 8.78104f
C11 drain_left a_n2982_n4888# 9.1962f
C12 source a_n2982_n4888# 13.895368f
C13 minus a_n2982_n4888# 12.540262f
C14 plus a_n2982_n4888# 14.74201f
C15 drain_right.t14 a_n2982_n4888# 0.429886f
C16 drain_right.t15 a_n2982_n4888# 0.429886f
C17 drain_right.n0 a_n2982_n4888# 3.93591f
C18 drain_right.t19 a_n2982_n4888# 0.429886f
C19 drain_right.t18 a_n2982_n4888# 0.429886f
C20 drain_right.n1 a_n2982_n4888# 3.93011f
C21 drain_right.n2 a_n2982_n4888# 0.771416f
C22 drain_right.t16 a_n2982_n4888# 0.429886f
C23 drain_right.t3 a_n2982_n4888# 0.429886f
C24 drain_right.n3 a_n2982_n4888# 3.93011f
C25 drain_right.t5 a_n2982_n4888# 0.429886f
C26 drain_right.t11 a_n2982_n4888# 0.429886f
C27 drain_right.n4 a_n2982_n4888# 3.93591f
C28 drain_right.t0 a_n2982_n4888# 0.429886f
C29 drain_right.t7 a_n2982_n4888# 0.429886f
C30 drain_right.n5 a_n2982_n4888# 3.93011f
C31 drain_right.n6 a_n2982_n4888# 0.771416f
C32 drain_right.n7 a_n2982_n4888# 2.46616f
C33 drain_right.t17 a_n2982_n4888# 0.429886f
C34 drain_right.t8 a_n2982_n4888# 0.429886f
C35 drain_right.n8 a_n2982_n4888# 3.9359f
C36 drain_right.t2 a_n2982_n4888# 0.429886f
C37 drain_right.t9 a_n2982_n4888# 0.429886f
C38 drain_right.n9 a_n2982_n4888# 3.93011f
C39 drain_right.n10 a_n2982_n4888# 0.775521f
C40 drain_right.t1 a_n2982_n4888# 0.429886f
C41 drain_right.t10 a_n2982_n4888# 0.429886f
C42 drain_right.n11 a_n2982_n4888# 3.93011f
C43 drain_right.n12 a_n2982_n4888# 0.38518f
C44 drain_right.t4 a_n2982_n4888# 0.429886f
C45 drain_right.t12 a_n2982_n4888# 0.429886f
C46 drain_right.n13 a_n2982_n4888# 3.93011f
C47 drain_right.n14 a_n2982_n4888# 0.38518f
C48 drain_right.t6 a_n2982_n4888# 0.429886f
C49 drain_right.t13 a_n2982_n4888# 0.429886f
C50 drain_right.n15 a_n2982_n4888# 3.93011f
C51 drain_right.n16 a_n2982_n4888# 0.625766f
C52 minus.n0 a_n2982_n4888# 0.039383f
C53 minus.n1 a_n2982_n4888# 0.008937f
C54 minus.t6 a_n2982_n4888# 1.5614f
C55 minus.n2 a_n2982_n4888# 0.039383f
C56 minus.n3 a_n2982_n4888# 0.008937f
C57 minus.t7 a_n2982_n4888# 1.5614f
C58 minus.n4 a_n2982_n4888# 0.039383f
C59 minus.n5 a_n2982_n4888# 0.008937f
C60 minus.t9 a_n2982_n4888# 1.5614f
C61 minus.n6 a_n2982_n4888# 0.039383f
C62 minus.n7 a_n2982_n4888# 0.008937f
C63 minus.t10 a_n2982_n4888# 1.5614f
C64 minus.t11 a_n2982_n4888# 1.58061f
C65 minus.t2 a_n2982_n4888# 1.5614f
C66 minus.n8 a_n2982_n4888# 0.588829f
C67 minus.n9 a_n2982_n4888# 0.565856f
C68 minus.n10 a_n2982_n4888# 0.168103f
C69 minus.n11 a_n2982_n4888# 0.039383f
C70 minus.n12 a_n2982_n4888# 0.582242f
C71 minus.n13 a_n2982_n4888# 0.008937f
C72 minus.t17 a_n2982_n4888# 1.5614f
C73 minus.n14 a_n2982_n4888# 0.582242f
C74 minus.n15 a_n2982_n4888# 0.039383f
C75 minus.n16 a_n2982_n4888# 0.039383f
C76 minus.n17 a_n2982_n4888# 0.039383f
C77 minus.n18 a_n2982_n4888# 0.582242f
C78 minus.n19 a_n2982_n4888# 0.008937f
C79 minus.t18 a_n2982_n4888# 1.5614f
C80 minus.n20 a_n2982_n4888# 0.582242f
C81 minus.n21 a_n2982_n4888# 0.039383f
C82 minus.n22 a_n2982_n4888# 0.039383f
C83 minus.n23 a_n2982_n4888# 0.039383f
C84 minus.n24 a_n2982_n4888# 0.582242f
C85 minus.n25 a_n2982_n4888# 0.008937f
C86 minus.t15 a_n2982_n4888# 1.5614f
C87 minus.n26 a_n2982_n4888# 0.582242f
C88 minus.n27 a_n2982_n4888# 0.039383f
C89 minus.n28 a_n2982_n4888# 0.039383f
C90 minus.n29 a_n2982_n4888# 0.039383f
C91 minus.n30 a_n2982_n4888# 0.582242f
C92 minus.n31 a_n2982_n4888# 0.008937f
C93 minus.t13 a_n2982_n4888# 1.5614f
C94 minus.n32 a_n2982_n4888# 0.581877f
C95 minus.n33 a_n2982_n4888# 2.03345f
C96 minus.n34 a_n2982_n4888# 0.039383f
C97 minus.n35 a_n2982_n4888# 0.008937f
C98 minus.n36 a_n2982_n4888# 0.039383f
C99 minus.n37 a_n2982_n4888# 0.008937f
C100 minus.n38 a_n2982_n4888# 0.039383f
C101 minus.n39 a_n2982_n4888# 0.008937f
C102 minus.n40 a_n2982_n4888# 0.039383f
C103 minus.n41 a_n2982_n4888# 0.008937f
C104 minus.t5 a_n2982_n4888# 1.58061f
C105 minus.t4 a_n2982_n4888# 1.5614f
C106 minus.n42 a_n2982_n4888# 0.588829f
C107 minus.n43 a_n2982_n4888# 0.565856f
C108 minus.n44 a_n2982_n4888# 0.168103f
C109 minus.n45 a_n2982_n4888# 0.039383f
C110 minus.t0 a_n2982_n4888# 1.5614f
C111 minus.n46 a_n2982_n4888# 0.582242f
C112 minus.n47 a_n2982_n4888# 0.008937f
C113 minus.t1 a_n2982_n4888# 1.5614f
C114 minus.n48 a_n2982_n4888# 0.582242f
C115 minus.n49 a_n2982_n4888# 0.039383f
C116 minus.n50 a_n2982_n4888# 0.039383f
C117 minus.n51 a_n2982_n4888# 0.039383f
C118 minus.t3 a_n2982_n4888# 1.5614f
C119 minus.n52 a_n2982_n4888# 0.582242f
C120 minus.n53 a_n2982_n4888# 0.008937f
C121 minus.t16 a_n2982_n4888# 1.5614f
C122 minus.n54 a_n2982_n4888# 0.582242f
C123 minus.n55 a_n2982_n4888# 0.039383f
C124 minus.n56 a_n2982_n4888# 0.039383f
C125 minus.n57 a_n2982_n4888# 0.039383f
C126 minus.t19 a_n2982_n4888# 1.5614f
C127 minus.n58 a_n2982_n4888# 0.582242f
C128 minus.n59 a_n2982_n4888# 0.008937f
C129 minus.t12 a_n2982_n4888# 1.5614f
C130 minus.n60 a_n2982_n4888# 0.582242f
C131 minus.n61 a_n2982_n4888# 0.039383f
C132 minus.n62 a_n2982_n4888# 0.039383f
C133 minus.n63 a_n2982_n4888# 0.039383f
C134 minus.t14 a_n2982_n4888# 1.5614f
C135 minus.n64 a_n2982_n4888# 0.582242f
C136 minus.n65 a_n2982_n4888# 0.008937f
C137 minus.t8 a_n2982_n4888# 1.5614f
C138 minus.n66 a_n2982_n4888# 0.581877f
C139 minus.n67 a_n2982_n4888# 0.272866f
C140 minus.n68 a_n2982_n4888# 2.39495f
C141 drain_left.t3 a_n2982_n4888# 0.431321f
C142 drain_left.t4 a_n2982_n4888# 0.431321f
C143 drain_left.n0 a_n2982_n4888# 3.94904f
C144 drain_left.t0 a_n2982_n4888# 0.431321f
C145 drain_left.t11 a_n2982_n4888# 0.431321f
C146 drain_left.n1 a_n2982_n4888# 3.94323f
C147 drain_left.n2 a_n2982_n4888# 0.773991f
C148 drain_left.t12 a_n2982_n4888# 0.431321f
C149 drain_left.t6 a_n2982_n4888# 0.431321f
C150 drain_left.n3 a_n2982_n4888# 3.94323f
C151 drain_left.t18 a_n2982_n4888# 0.431321f
C152 drain_left.t19 a_n2982_n4888# 0.431321f
C153 drain_left.n4 a_n2982_n4888# 3.94904f
C154 drain_left.t7 a_n2982_n4888# 0.431321f
C155 drain_left.t2 a_n2982_n4888# 0.431321f
C156 drain_left.n5 a_n2982_n4888# 3.94323f
C157 drain_left.n6 a_n2982_n4888# 0.773991f
C158 drain_left.n7 a_n2982_n4888# 2.53032f
C159 drain_left.t13 a_n2982_n4888# 0.431321f
C160 drain_left.t5 a_n2982_n4888# 0.431321f
C161 drain_left.n8 a_n2982_n4888# 3.94904f
C162 drain_left.t16 a_n2982_n4888# 0.431321f
C163 drain_left.t9 a_n2982_n4888# 0.431321f
C164 drain_left.n9 a_n2982_n4888# 3.94322f
C165 drain_left.n10 a_n2982_n4888# 0.778109f
C166 drain_left.t14 a_n2982_n4888# 0.431321f
C167 drain_left.t8 a_n2982_n4888# 0.431321f
C168 drain_left.n11 a_n2982_n4888# 3.94322f
C169 drain_left.n12 a_n2982_n4888# 0.386465f
C170 drain_left.t17 a_n2982_n4888# 0.431321f
C171 drain_left.t10 a_n2982_n4888# 0.431321f
C172 drain_left.n13 a_n2982_n4888# 3.94322f
C173 drain_left.n14 a_n2982_n4888# 0.386465f
C174 drain_left.t1 a_n2982_n4888# 0.431321f
C175 drain_left.t15 a_n2982_n4888# 0.431321f
C176 drain_left.n15 a_n2982_n4888# 3.94322f
C177 drain_left.n16 a_n2982_n4888# 0.627854f
C178 source.t21 a_n2982_n4888# 4.23479f
C179 source.n0 a_n2982_n4888# 1.84225f
C180 source.t32 a_n2982_n4888# 0.37055f
C181 source.t29 a_n2982_n4888# 0.37055f
C182 source.n1 a_n2982_n4888# 3.31288f
C183 source.n2 a_n2982_n4888# 0.374917f
C184 source.t35 a_n2982_n4888# 0.37055f
C185 source.t33 a_n2982_n4888# 0.37055f
C186 source.n3 a_n2982_n4888# 3.31288f
C187 source.n4 a_n2982_n4888# 0.374917f
C188 source.t39 a_n2982_n4888# 0.37055f
C189 source.t28 a_n2982_n4888# 0.37055f
C190 source.n5 a_n2982_n4888# 3.31288f
C191 source.n6 a_n2982_n4888# 0.374917f
C192 source.t34 a_n2982_n4888# 0.37055f
C193 source.t31 a_n2982_n4888# 0.37055f
C194 source.n7 a_n2982_n4888# 3.31288f
C195 source.n8 a_n2982_n4888# 0.374917f
C196 source.t36 a_n2982_n4888# 4.2348f
C197 source.n9 a_n2982_n4888# 0.432001f
C198 source.t5 a_n2982_n4888# 4.2348f
C199 source.n10 a_n2982_n4888# 0.432001f
C200 source.t12 a_n2982_n4888# 0.37055f
C201 source.t7 a_n2982_n4888# 0.37055f
C202 source.n11 a_n2982_n4888# 3.31288f
C203 source.n12 a_n2982_n4888# 0.374917f
C204 source.t4 a_n2982_n4888# 0.37055f
C205 source.t11 a_n2982_n4888# 0.37055f
C206 source.n13 a_n2982_n4888# 3.31288f
C207 source.n14 a_n2982_n4888# 0.374917f
C208 source.t18 a_n2982_n4888# 0.37055f
C209 source.t17 a_n2982_n4888# 0.37055f
C210 source.n15 a_n2982_n4888# 3.31288f
C211 source.n16 a_n2982_n4888# 0.374917f
C212 source.t10 a_n2982_n4888# 0.37055f
C213 source.t0 a_n2982_n4888# 0.37055f
C214 source.n17 a_n2982_n4888# 3.31288f
C215 source.n18 a_n2982_n4888# 0.374917f
C216 source.t6 a_n2982_n4888# 4.2348f
C217 source.n19 a_n2982_n4888# 2.26879f
C218 source.t25 a_n2982_n4888# 4.23477f
C219 source.n20 a_n2982_n4888# 2.26881f
C220 source.t37 a_n2982_n4888# 0.37055f
C221 source.t20 a_n2982_n4888# 0.37055f
C222 source.n21 a_n2982_n4888# 3.31288f
C223 source.n22 a_n2982_n4888# 0.37491f
C224 source.t24 a_n2982_n4888# 0.37055f
C225 source.t38 a_n2982_n4888# 0.37055f
C226 source.n23 a_n2982_n4888# 3.31288f
C227 source.n24 a_n2982_n4888# 0.37491f
C228 source.t27 a_n2982_n4888# 0.37055f
C229 source.t23 a_n2982_n4888# 0.37055f
C230 source.n25 a_n2982_n4888# 3.31288f
C231 source.n26 a_n2982_n4888# 0.37491f
C232 source.t30 a_n2982_n4888# 0.37055f
C233 source.t26 a_n2982_n4888# 0.37055f
C234 source.n27 a_n2982_n4888# 3.31288f
C235 source.n28 a_n2982_n4888# 0.37491f
C236 source.t22 a_n2982_n4888# 4.23477f
C237 source.n29 a_n2982_n4888# 0.432025f
C238 source.t9 a_n2982_n4888# 4.23477f
C239 source.n30 a_n2982_n4888# 0.432025f
C240 source.t1 a_n2982_n4888# 0.37055f
C241 source.t15 a_n2982_n4888# 0.37055f
C242 source.n31 a_n2982_n4888# 3.31288f
C243 source.n32 a_n2982_n4888# 0.37491f
C244 source.t3 a_n2982_n4888# 0.37055f
C245 source.t8 a_n2982_n4888# 0.37055f
C246 source.n33 a_n2982_n4888# 3.31288f
C247 source.n34 a_n2982_n4888# 0.37491f
C248 source.t14 a_n2982_n4888# 0.37055f
C249 source.t13 a_n2982_n4888# 0.37055f
C250 source.n35 a_n2982_n4888# 3.31288f
C251 source.n36 a_n2982_n4888# 0.37491f
C252 source.t2 a_n2982_n4888# 0.37055f
C253 source.t16 a_n2982_n4888# 0.37055f
C254 source.n37 a_n2982_n4888# 3.31288f
C255 source.n38 a_n2982_n4888# 0.37491f
C256 source.t19 a_n2982_n4888# 4.23477f
C257 source.n39 a_n2982_n4888# 0.584962f
C258 source.n40 a_n2982_n4888# 2.12707f
C259 plus.n0 a_n2982_n4888# 0.039687f
C260 plus.t4 a_n2982_n4888# 1.57347f
C261 plus.t18 a_n2982_n4888# 1.57347f
C262 plus.n1 a_n2982_n4888# 0.039687f
C263 plus.t9 a_n2982_n4888# 1.57347f
C264 plus.n2 a_n2982_n4888# 0.586742f
C265 plus.n3 a_n2982_n4888# 0.039687f
C266 plus.t2 a_n2982_n4888# 1.57347f
C267 plus.t11 a_n2982_n4888# 1.57347f
C268 plus.n4 a_n2982_n4888# 0.586742f
C269 plus.n5 a_n2982_n4888# 0.039687f
C270 plus.t5 a_n2982_n4888# 1.57347f
C271 plus.t10 a_n2982_n4888# 1.57347f
C272 plus.n6 a_n2982_n4888# 0.586742f
C273 plus.n7 a_n2982_n4888# 0.039687f
C274 plus.t3 a_n2982_n4888# 1.57347f
C275 plus.t14 a_n2982_n4888# 1.57347f
C276 plus.n8 a_n2982_n4888# 0.59338f
C277 plus.t6 a_n2982_n4888# 1.59283f
C278 plus.n9 a_n2982_n4888# 0.57023f
C279 plus.n10 a_n2982_n4888# 0.169402f
C280 plus.n11 a_n2982_n4888# 0.009006f
C281 plus.n12 a_n2982_n4888# 0.586742f
C282 plus.n13 a_n2982_n4888# 0.009006f
C283 plus.n14 a_n2982_n4888# 0.039687f
C284 plus.n15 a_n2982_n4888# 0.039687f
C285 plus.n16 a_n2982_n4888# 0.039687f
C286 plus.n17 a_n2982_n4888# 0.009006f
C287 plus.n18 a_n2982_n4888# 0.586742f
C288 plus.n19 a_n2982_n4888# 0.009006f
C289 plus.n20 a_n2982_n4888# 0.039687f
C290 plus.n21 a_n2982_n4888# 0.039687f
C291 plus.n22 a_n2982_n4888# 0.039687f
C292 plus.n23 a_n2982_n4888# 0.009006f
C293 plus.n24 a_n2982_n4888# 0.586742f
C294 plus.n25 a_n2982_n4888# 0.009006f
C295 plus.n26 a_n2982_n4888# 0.039687f
C296 plus.n27 a_n2982_n4888# 0.039687f
C297 plus.n28 a_n2982_n4888# 0.039687f
C298 plus.n29 a_n2982_n4888# 0.009006f
C299 plus.n30 a_n2982_n4888# 0.586742f
C300 plus.n31 a_n2982_n4888# 0.009006f
C301 plus.n32 a_n2982_n4888# 0.586375f
C302 plus.n33 a_n2982_n4888# 0.617839f
C303 plus.n34 a_n2982_n4888# 0.039687f
C304 plus.t16 a_n2982_n4888# 1.57347f
C305 plus.n35 a_n2982_n4888# 0.039687f
C306 plus.t15 a_n2982_n4888# 1.57347f
C307 plus.t19 a_n2982_n4888# 1.57347f
C308 plus.n36 a_n2982_n4888# 0.586742f
C309 plus.n37 a_n2982_n4888# 0.039687f
C310 plus.t8 a_n2982_n4888# 1.57347f
C311 plus.t7 a_n2982_n4888# 1.57347f
C312 plus.n38 a_n2982_n4888# 0.586742f
C313 plus.n39 a_n2982_n4888# 0.039687f
C314 plus.t13 a_n2982_n4888# 1.57347f
C315 plus.t12 a_n2982_n4888# 1.57347f
C316 plus.n40 a_n2982_n4888# 0.586742f
C317 plus.n41 a_n2982_n4888# 0.039687f
C318 plus.t17 a_n2982_n4888# 1.57347f
C319 plus.t1 a_n2982_n4888# 1.57347f
C320 plus.n42 a_n2982_n4888# 0.59338f
C321 plus.t0 a_n2982_n4888# 1.59283f
C322 plus.n43 a_n2982_n4888# 0.57023f
C323 plus.n44 a_n2982_n4888# 0.169402f
C324 plus.n45 a_n2982_n4888# 0.009006f
C325 plus.n46 a_n2982_n4888# 0.586742f
C326 plus.n47 a_n2982_n4888# 0.009006f
C327 plus.n48 a_n2982_n4888# 0.039687f
C328 plus.n49 a_n2982_n4888# 0.039687f
C329 plus.n50 a_n2982_n4888# 0.039687f
C330 plus.n51 a_n2982_n4888# 0.009006f
C331 plus.n52 a_n2982_n4888# 0.586742f
C332 plus.n53 a_n2982_n4888# 0.009006f
C333 plus.n54 a_n2982_n4888# 0.039687f
C334 plus.n55 a_n2982_n4888# 0.039687f
C335 plus.n56 a_n2982_n4888# 0.039687f
C336 plus.n57 a_n2982_n4888# 0.009006f
C337 plus.n58 a_n2982_n4888# 0.586742f
C338 plus.n59 a_n2982_n4888# 0.009006f
C339 plus.n60 a_n2982_n4888# 0.039687f
C340 plus.n61 a_n2982_n4888# 0.039687f
C341 plus.n62 a_n2982_n4888# 0.039687f
C342 plus.n63 a_n2982_n4888# 0.009006f
C343 plus.n64 a_n2982_n4888# 0.586742f
C344 plus.n65 a_n2982_n4888# 0.009006f
C345 plus.n66 a_n2982_n4888# 0.586375f
C346 plus.n67 a_n2982_n4888# 1.65115f
.ends

