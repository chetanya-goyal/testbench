* NGSPICE file created from diffpair543.ext - technology: sky130A

.subckt diffpair543 minus drain_right drain_left source plus
X0 a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X1 source.t15 minus.t0 drain_right.t2 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X2 drain_left.t7 plus.t0 source.t7 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X3 source.t6 plus.t1 drain_left.t6 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X4 source.t3 plus.t2 drain_left.t5 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 source.t14 minus.t1 drain_right.t5 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X6 drain_right.t0 minus.t2 source.t13 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X7 a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X8 source.t5 plus.t3 drain_left.t4 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X9 source.t12 minus.t3 drain_right.t1 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X10 drain_right.t6 minus.t4 source.t11 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X11 a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X12 drain_right.t4 minus.t5 source.t10 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X13 drain_left.t3 plus.t4 source.t4 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X14 drain_right.t3 minus.t6 source.t9 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X15 source.t0 plus.t5 drain_left.t2 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X16 drain_left.t1 plus.t6 source.t1 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X17 a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X18 drain_left.t0 plus.t7 source.t2 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X19 source.t8 minus.t7 drain_right.t7 a_n1746_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
R0 minus.n3 minus.t6 594.726
R1 minus.n13 minus.t3 594.726
R2 minus.n2 minus.t1 572.548
R3 minus.n6 minus.t5 572.548
R4 minus.n8 minus.t7 572.548
R5 minus.n12 minus.t4 572.548
R6 minus.n16 minus.t0 572.548
R7 minus.n18 minus.t2 572.548
R8 minus.n9 minus.n8 161.3
R9 minus.n7 minus.n0 161.3
R10 minus.n6 minus.n5 161.3
R11 minus.n4 minus.n1 161.3
R12 minus.n19 minus.n18 161.3
R13 minus.n17 minus.n10 161.3
R14 minus.n16 minus.n15 161.3
R15 minus.n14 minus.n11 161.3
R16 minus.n4 minus.n3 44.862
R17 minus.n14 minus.n13 44.862
R18 minus.n20 minus.n9 38.1406
R19 minus.n8 minus.n7 28.4823
R20 minus.n18 minus.n17 28.4823
R21 minus.n6 minus.n1 24.1005
R22 minus.n2 minus.n1 24.1005
R23 minus.n12 minus.n11 24.1005
R24 minus.n16 minus.n11 24.1005
R25 minus.n7 minus.n6 19.7187
R26 minus.n17 minus.n16 19.7187
R27 minus.n3 minus.n2 19.7081
R28 minus.n13 minus.n12 19.7081
R29 minus.n20 minus.n19 6.63308
R30 minus.n9 minus.n0 0.189894
R31 minus.n5 minus.n0 0.189894
R32 minus.n5 minus.n4 0.189894
R33 minus.n15 minus.n14 0.189894
R34 minus.n15 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 drain_right.n5 drain_right.n3 61.7676
R38 drain_right.n2 drain_right.n1 61.2682
R39 drain_right.n2 drain_right.n0 61.2682
R40 drain_right.n5 drain_right.n4 60.8798
R41 drain_right drain_right.n2 32.1943
R42 drain_right drain_right.n5 6.54115
R43 drain_right.n1 drain_right.t2 1.3205
R44 drain_right.n1 drain_right.t0 1.3205
R45 drain_right.n0 drain_right.t1 1.3205
R46 drain_right.n0 drain_right.t6 1.3205
R47 drain_right.n3 drain_right.t5 1.3205
R48 drain_right.n3 drain_right.t3 1.3205
R49 drain_right.n4 drain_right.t7 1.3205
R50 drain_right.n4 drain_right.t4 1.3205
R51 source.n3 source.t5 45.521
R52 source.n4 source.t9 45.521
R53 source.n7 source.t8 45.521
R54 source.n15 source.t13 45.5208
R55 source.n12 source.t12 45.5208
R56 source.n11 source.t7 45.5208
R57 source.n8 source.t0 45.5208
R58 source.n0 source.t4 45.5208
R59 source.n2 source.n1 44.201
R60 source.n6 source.n5 44.201
R61 source.n14 source.n13 44.2008
R62 source.n10 source.n9 44.2008
R63 source.n8 source.n7 24.4484
R64 source.n16 source.n0 18.7415
R65 source.n16 source.n15 5.7074
R66 source.n13 source.t11 1.3205
R67 source.n13 source.t15 1.3205
R68 source.n9 source.t2 1.3205
R69 source.n9 source.t6 1.3205
R70 source.n1 source.t1 1.3205
R71 source.n1 source.t3 1.3205
R72 source.n5 source.t10 1.3205
R73 source.n5 source.t14 1.3205
R74 source.n7 source.n6 0.888431
R75 source.n6 source.n4 0.888431
R76 source.n3 source.n2 0.888431
R77 source.n2 source.n0 0.888431
R78 source.n10 source.n8 0.888431
R79 source.n11 source.n10 0.888431
R80 source.n14 source.n12 0.888431
R81 source.n15 source.n14 0.888431
R82 source.n4 source.n3 0.470328
R83 source.n12 source.n11 0.470328
R84 source source.n16 0.188
R85 plus.n3 plus.t3 594.726
R86 plus.n13 plus.t0 594.726
R87 plus.n8 plus.t4 572.548
R88 plus.n6 plus.t2 572.548
R89 plus.n2 plus.t6 572.548
R90 plus.n18 plus.t5 572.548
R91 plus.n16 plus.t7 572.548
R92 plus.n12 plus.t1 572.548
R93 plus.n5 plus.n4 161.3
R94 plus.n6 plus.n1 161.3
R95 plus.n7 plus.n0 161.3
R96 plus.n9 plus.n8 161.3
R97 plus.n15 plus.n14 161.3
R98 plus.n16 plus.n11 161.3
R99 plus.n17 plus.n10 161.3
R100 plus.n19 plus.n18 161.3
R101 plus.n4 plus.n3 44.862
R102 plus.n14 plus.n13 44.862
R103 plus plus.n19 30.8854
R104 plus.n8 plus.n7 28.4823
R105 plus.n18 plus.n17 28.4823
R106 plus.n5 plus.n2 24.1005
R107 plus.n6 plus.n5 24.1005
R108 plus.n16 plus.n15 24.1005
R109 plus.n15 plus.n12 24.1005
R110 plus.n7 plus.n6 19.7187
R111 plus.n17 plus.n16 19.7187
R112 plus.n3 plus.n2 19.7081
R113 plus.n13 plus.n12 19.7081
R114 plus plus.n9 13.4134
R115 plus.n4 plus.n1 0.189894
R116 plus.n1 plus.n0 0.189894
R117 plus.n9 plus.n0 0.189894
R118 plus.n19 plus.n10 0.189894
R119 plus.n11 plus.n10 0.189894
R120 plus.n14 plus.n11 0.189894
R121 drain_left.n5 drain_left.n3 61.7677
R122 drain_left.n2 drain_left.n1 61.2682
R123 drain_left.n2 drain_left.n0 61.2682
R124 drain_left.n5 drain_left.n4 60.8796
R125 drain_left drain_left.n2 32.7476
R126 drain_left drain_left.n5 6.54115
R127 drain_left.n1 drain_left.t6 1.3205
R128 drain_left.n1 drain_left.t7 1.3205
R129 drain_left.n0 drain_left.t2 1.3205
R130 drain_left.n0 drain_left.t0 1.3205
R131 drain_left.n4 drain_left.t5 1.3205
R132 drain_left.n4 drain_left.t3 1.3205
R133 drain_left.n3 drain_left.t4 1.3205
R134 drain_left.n3 drain_left.t1 1.3205
C0 source minus 6.44367f
C1 drain_left source 13.4932f
C2 drain_right source 13.495f
C3 drain_left minus 0.171089f
C4 source plus 6.45771f
C5 drain_right minus 6.81873f
C6 drain_left drain_right 0.821811f
C7 plus minus 5.87497f
C8 drain_left plus 6.98757f
C9 drain_right plus 0.322995f
C10 drain_right a_n1746_n3888# 6.24063f
C11 drain_left a_n1746_n3888# 6.50199f
C12 source a_n1746_n3888# 10.655262f
C13 minus a_n1746_n3888# 6.965223f
C14 plus a_n1746_n3888# 8.826839f
C15 drain_left.t2 a_n1746_n3888# 0.323271f
C16 drain_left.t0 a_n1746_n3888# 0.323271f
C17 drain_left.n0 a_n1746_n3888# 2.9242f
C18 drain_left.t6 a_n1746_n3888# 0.323271f
C19 drain_left.t7 a_n1746_n3888# 0.323271f
C20 drain_left.n1 a_n1746_n3888# 2.9242f
C21 drain_left.n2 a_n1746_n3888# 2.21889f
C22 drain_left.t4 a_n1746_n3888# 0.323271f
C23 drain_left.t1 a_n1746_n3888# 0.323271f
C24 drain_left.n3 a_n1746_n3888# 2.92761f
C25 drain_left.t5 a_n1746_n3888# 0.323271f
C26 drain_left.t3 a_n1746_n3888# 0.323271f
C27 drain_left.n4 a_n1746_n3888# 2.92198f
C28 drain_left.n5 a_n1746_n3888# 1.00547f
C29 plus.n0 a_n1746_n3888# 0.04465f
C30 plus.t4 a_n1746_n3888# 1.33225f
C31 plus.t2 a_n1746_n3888# 1.33225f
C32 plus.n1 a_n1746_n3888# 0.04465f
C33 plus.t6 a_n1746_n3888# 1.33225f
C34 plus.n2 a_n1746_n3888# 0.518161f
C35 plus.t3 a_n1746_n3888# 1.35142f
C36 plus.n3 a_n1746_n3888# 0.499065f
C37 plus.n4 a_n1746_n3888# 0.185675f
C38 plus.n5 a_n1746_n3888# 0.010132f
C39 plus.n6 a_n1746_n3888# 0.51412f
C40 plus.n7 a_n1746_n3888# 0.010132f
C41 plus.n8 a_n1746_n3888# 0.51123f
C42 plus.n9 a_n1746_n3888# 0.578187f
C43 plus.n10 a_n1746_n3888# 0.04465f
C44 plus.t5 a_n1746_n3888# 1.33225f
C45 plus.n11 a_n1746_n3888# 0.04465f
C46 plus.t7 a_n1746_n3888# 1.33225f
C47 plus.t1 a_n1746_n3888# 1.33225f
C48 plus.n12 a_n1746_n3888# 0.518161f
C49 plus.t0 a_n1746_n3888# 1.35142f
C50 plus.n13 a_n1746_n3888# 0.499065f
C51 plus.n14 a_n1746_n3888# 0.185675f
C52 plus.n15 a_n1746_n3888# 0.010132f
C53 plus.n16 a_n1746_n3888# 0.51412f
C54 plus.n17 a_n1746_n3888# 0.010132f
C55 plus.n18 a_n1746_n3888# 0.51123f
C56 plus.n19 a_n1746_n3888# 1.41217f
C57 source.t4 a_n1746_n3888# 2.60894f
C58 source.n0 a_n1746_n3888# 1.24358f
C59 source.t1 a_n1746_n3888# 0.232803f
C60 source.t3 a_n1746_n3888# 0.232803f
C61 source.n1 a_n1746_n3888# 2.04498f
C62 source.n2 a_n1746_n3888# 0.305843f
C63 source.t5 a_n1746_n3888# 2.60894f
C64 source.n3 a_n1746_n3888# 0.350344f
C65 source.t9 a_n1746_n3888# 2.60894f
C66 source.n4 a_n1746_n3888# 0.350344f
C67 source.t10 a_n1746_n3888# 0.232803f
C68 source.t14 a_n1746_n3888# 0.232803f
C69 source.n5 a_n1746_n3888# 2.04498f
C70 source.n6 a_n1746_n3888# 0.305843f
C71 source.t8 a_n1746_n3888# 2.60894f
C72 source.n7 a_n1746_n3888# 1.57859f
C73 source.t0 a_n1746_n3888# 2.60894f
C74 source.n8 a_n1746_n3888# 1.57859f
C75 source.t2 a_n1746_n3888# 0.232803f
C76 source.t6 a_n1746_n3888# 0.232803f
C77 source.n9 a_n1746_n3888# 2.04498f
C78 source.n10 a_n1746_n3888# 0.305846f
C79 source.t7 a_n1746_n3888# 2.60894f
C80 source.n11 a_n1746_n3888# 0.350347f
C81 source.t12 a_n1746_n3888# 2.60894f
C82 source.n12 a_n1746_n3888# 0.350347f
C83 source.t11 a_n1746_n3888# 0.232803f
C84 source.t15 a_n1746_n3888# 0.232803f
C85 source.n13 a_n1746_n3888# 2.04498f
C86 source.n14 a_n1746_n3888# 0.305846f
C87 source.t13 a_n1746_n3888# 2.60894f
C88 source.n15 a_n1746_n3888# 0.47846f
C89 source.n16 a_n1746_n3888# 1.4491f
C90 drain_right.t1 a_n1746_n3888# 0.321792f
C91 drain_right.t6 a_n1746_n3888# 0.321792f
C92 drain_right.n0 a_n1746_n3888# 2.91082f
C93 drain_right.t2 a_n1746_n3888# 0.321792f
C94 drain_right.t0 a_n1746_n3888# 0.321792f
C95 drain_right.n1 a_n1746_n3888# 2.91082f
C96 drain_right.n2 a_n1746_n3888# 2.15212f
C97 drain_right.t5 a_n1746_n3888# 0.321792f
C98 drain_right.t3 a_n1746_n3888# 0.321792f
C99 drain_right.n3 a_n1746_n3888# 2.9142f
C100 drain_right.t7 a_n1746_n3888# 0.321792f
C101 drain_right.t4 a_n1746_n3888# 0.321792f
C102 drain_right.n4 a_n1746_n3888# 2.90862f
C103 drain_right.n5 a_n1746_n3888# 1.00087f
C104 minus.n0 a_n1746_n3888# 0.043756f
C105 minus.n1 a_n1746_n3888# 0.009929f
C106 minus.t5 a_n1746_n3888# 1.30558f
C107 minus.t6 a_n1746_n3888# 1.32436f
C108 minus.t1 a_n1746_n3888# 1.30558f
C109 minus.n2 a_n1746_n3888# 0.507785f
C110 minus.n3 a_n1746_n3888# 0.489071f
C111 minus.n4 a_n1746_n3888# 0.181957f
C112 minus.n5 a_n1746_n3888# 0.043756f
C113 minus.n6 a_n1746_n3888# 0.503825f
C114 minus.n7 a_n1746_n3888# 0.009929f
C115 minus.t7 a_n1746_n3888# 1.30558f
C116 minus.n8 a_n1746_n3888# 0.500993f
C117 minus.n9 a_n1746_n3888# 1.68113f
C118 minus.n10 a_n1746_n3888# 0.043756f
C119 minus.n11 a_n1746_n3888# 0.009929f
C120 minus.t3 a_n1746_n3888# 1.32436f
C121 minus.t4 a_n1746_n3888# 1.30558f
C122 minus.n12 a_n1746_n3888# 0.507785f
C123 minus.n13 a_n1746_n3888# 0.489071f
C124 minus.n14 a_n1746_n3888# 0.181957f
C125 minus.n15 a_n1746_n3888# 0.043756f
C126 minus.t0 a_n1746_n3888# 1.30558f
C127 minus.n16 a_n1746_n3888# 0.503825f
C128 minus.n17 a_n1746_n3888# 0.009929f
C129 minus.t2 a_n1746_n3888# 1.30558f
C130 minus.n18 a_n1746_n3888# 0.500993f
C131 minus.n19 a_n1746_n3888# 0.299696f
C132 minus.n20 a_n1746_n3888# 2.02628f
.ends

