* NGSPICE file created from diffpair364.ext - technology: sky130A

.subckt diffpair364 minus drain_right drain_left source plus
X0 a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X1 drain_right.t9 minus.t0 source.t6 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X2 a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X3 drain_left.t9 plus.t0 source.t17 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 source.t8 minus.t1 drain_right.t8 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 drain_left.t8 plus.t1 source.t18 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X6 drain_right.t7 minus.t2 source.t7 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X7 source.t10 minus.t3 drain_right.t6 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X8 drain_right.t5 minus.t4 source.t11 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 drain_right.t4 minus.t5 source.t14 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 source.t19 plus.t2 drain_left.t7 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X12 a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X13 drain_right.t3 minus.t6 source.t9 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X14 source.t1 plus.t3 drain_left.t6 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 drain_left.t5 plus.t4 source.t0 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X16 source.t2 plus.t5 drain_left.t4 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 source.t15 minus.t7 drain_right.t2 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 drain_left.t3 plus.t6 source.t4 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X19 source.t5 plus.t7 drain_left.t2 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 drain_left.t1 plus.t8 source.t3 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X21 drain_left.t0 plus.t9 source.t16 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X22 source.t12 minus.t8 drain_right.t1 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 drain_right.t0 minus.t9 source.t13 a_n1712_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n2 minus.t6 533.348
R1 minus.n14 minus.t9 533.348
R2 minus.n3 minus.t1 512.366
R3 minus.n1 minus.t4 512.366
R4 minus.n9 minus.t7 512.366
R5 minus.n10 minus.t2 512.366
R6 minus.n15 minus.t8 512.366
R7 minus.n13 minus.t5 512.366
R8 minus.n21 minus.t3 512.366
R9 minus.n22 minus.t0 512.366
R10 minus.n11 minus.n10 161.3
R11 minus.n9 minus.n0 161.3
R12 minus.n8 minus.n7 161.3
R13 minus.n6 minus.n1 161.3
R14 minus.n5 minus.n4 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n18 minus.n13 161.3
R19 minus.n17 minus.n16 161.3
R20 minus.n5 minus.n2 70.4033
R21 minus.n17 minus.n14 70.4033
R22 minus.n10 minus.n9 48.2005
R23 minus.n22 minus.n21 48.2005
R24 minus.n4 minus.n1 36.5157
R25 minus.n8 minus.n1 36.5157
R26 minus.n16 minus.n13 36.5157
R27 minus.n20 minus.n13 36.5157
R28 minus.n24 minus.n11 33.3963
R29 minus.n3 minus.n2 20.9576
R30 minus.n15 minus.n14 20.9576
R31 minus.n4 minus.n3 11.6853
R32 minus.n9 minus.n8 11.6853
R33 minus.n16 minus.n15 11.6853
R34 minus.n21 minus.n20 11.6853
R35 minus.n24 minus.n23 6.563
R36 minus.n11 minus.n0 0.189894
R37 minus.n7 minus.n0 0.189894
R38 minus.n7 minus.n6 0.189894
R39 minus.n6 minus.n5 0.189894
R40 minus.n18 minus.n17 0.189894
R41 minus.n19 minus.n18 0.189894
R42 minus.n19 minus.n12 0.189894
R43 minus.n23 minus.n12 0.189894
R44 minus minus.n24 0.188
R45 source.n5 source.t9 51.0588
R46 source.n19 source.t6 51.0586
R47 source.n14 source.t0 51.0586
R48 source.n0 source.t4 51.0586
R49 source.n2 source.n1 48.8588
R50 source.n4 source.n3 48.8588
R51 source.n7 source.n6 48.8588
R52 source.n9 source.n8 48.8588
R53 source.n18 source.n17 48.8586
R54 source.n16 source.n15 48.8586
R55 source.n13 source.n12 48.8586
R56 source.n11 source.n10 48.8586
R57 source.n11 source.n9 20.446
R58 source.n20 source.n0 14.1098
R59 source.n20 source.n19 5.62119
R60 source.n17 source.t14 2.2005
R61 source.n17 source.t10 2.2005
R62 source.n15 source.t13 2.2005
R63 source.n15 source.t12 2.2005
R64 source.n12 source.t17 2.2005
R65 source.n12 source.t2 2.2005
R66 source.n10 source.t3 2.2005
R67 source.n10 source.t5 2.2005
R68 source.n1 source.t16 2.2005
R69 source.n1 source.t19 2.2005
R70 source.n3 source.t18 2.2005
R71 source.n3 source.t1 2.2005
R72 source.n6 source.t11 2.2005
R73 source.n6 source.t8 2.2005
R74 source.n8 source.t7 2.2005
R75 source.n8 source.t15 2.2005
R76 source.n5 source.n4 0.828086
R77 source.n16 source.n14 0.828086
R78 source.n9 source.n7 0.716017
R79 source.n7 source.n5 0.716017
R80 source.n4 source.n2 0.716017
R81 source.n2 source.n0 0.716017
R82 source.n13 source.n11 0.716017
R83 source.n14 source.n13 0.716017
R84 source.n18 source.n16 0.716017
R85 source.n19 source.n18 0.716017
R86 source source.n20 0.188
R87 drain_right.n1 drain_right.t0 68.4529
R88 drain_right.n7 drain_right.t7 67.7376
R89 drain_right.n6 drain_right.n4 66.2529
R90 drain_right.n3 drain_right.n2 66.0186
R91 drain_right.n6 drain_right.n5 65.5376
R92 drain_right.n1 drain_right.n0 65.5373
R93 drain_right drain_right.n3 27.5821
R94 drain_right drain_right.n7 6.01097
R95 drain_right.n2 drain_right.t6 2.2005
R96 drain_right.n2 drain_right.t9 2.2005
R97 drain_right.n0 drain_right.t1 2.2005
R98 drain_right.n0 drain_right.t4 2.2005
R99 drain_right.n4 drain_right.t8 2.2005
R100 drain_right.n4 drain_right.t3 2.2005
R101 drain_right.n5 drain_right.t2 2.2005
R102 drain_right.n5 drain_right.t5 2.2005
R103 drain_right.n7 drain_right.n6 0.716017
R104 drain_right.n3 drain_right.n1 0.124033
R105 plus.n2 plus.t1 533.348
R106 plus.n14 plus.t4 533.348
R107 plus.n10 plus.t6 512.366
R108 plus.n9 plus.t2 512.366
R109 plus.n1 plus.t9 512.366
R110 plus.n3 plus.t3 512.366
R111 plus.n22 plus.t8 512.366
R112 plus.n21 plus.t7 512.366
R113 plus.n13 plus.t0 512.366
R114 plus.n15 plus.t5 512.366
R115 plus.n5 plus.n4 161.3
R116 plus.n6 plus.n1 161.3
R117 plus.n8 plus.n7 161.3
R118 plus.n9 plus.n0 161.3
R119 plus.n11 plus.n10 161.3
R120 plus.n17 plus.n16 161.3
R121 plus.n18 plus.n13 161.3
R122 plus.n20 plus.n19 161.3
R123 plus.n21 plus.n12 161.3
R124 plus.n23 plus.n22 161.3
R125 plus.n5 plus.n2 70.4033
R126 plus.n17 plus.n14 70.4033
R127 plus.n10 plus.n9 48.2005
R128 plus.n22 plus.n21 48.2005
R129 plus.n8 plus.n1 36.5157
R130 plus.n4 plus.n1 36.5157
R131 plus.n20 plus.n13 36.5157
R132 plus.n16 plus.n13 36.5157
R133 plus plus.n23 28.4138
R134 plus.n3 plus.n2 20.9576
R135 plus.n15 plus.n14 20.9576
R136 plus.n9 plus.n8 11.6853
R137 plus.n4 plus.n3 11.6853
R138 plus.n21 plus.n20 11.6853
R139 plus.n16 plus.n15 11.6853
R140 plus plus.n11 11.0706
R141 plus.n6 plus.n5 0.189894
R142 plus.n7 plus.n6 0.189894
R143 plus.n7 plus.n0 0.189894
R144 plus.n11 plus.n0 0.189894
R145 plus.n23 plus.n12 0.189894
R146 plus.n19 plus.n12 0.189894
R147 plus.n19 plus.n18 0.189894
R148 plus.n18 plus.n17 0.189894
R149 drain_left.n5 drain_left.t8 68.4531
R150 drain_left.n1 drain_left.t1 68.4529
R151 drain_left.n3 drain_left.n2 66.0186
R152 drain_left.n5 drain_left.n4 65.5376
R153 drain_left.n7 drain_left.n6 65.5374
R154 drain_left.n1 drain_left.n0 65.5373
R155 drain_left drain_left.n3 28.1353
R156 drain_left drain_left.n7 6.36873
R157 drain_left.n2 drain_left.t4 2.2005
R158 drain_left.n2 drain_left.t5 2.2005
R159 drain_left.n0 drain_left.t2 2.2005
R160 drain_left.n0 drain_left.t9 2.2005
R161 drain_left.n6 drain_left.t7 2.2005
R162 drain_left.n6 drain_left.t3 2.2005
R163 drain_left.n4 drain_left.t6 2.2005
R164 drain_left.n4 drain_left.t0 2.2005
R165 drain_left.n7 drain_left.n5 0.716017
R166 drain_left.n3 drain_left.n1 0.124033
C0 plus source 4.11124f
C1 drain_left source 13.109599f
C2 drain_right minus 4.25568f
C3 plus drain_right 0.321603f
C4 drain_right drain_left 0.846116f
C5 drain_right source 13.103f
C6 plus minus 4.72692f
C7 minus drain_left 0.171781f
C8 plus drain_left 4.41905f
C9 minus source 4.09677f
C10 drain_right a_n1712_n2688# 5.99024f
C11 drain_left a_n1712_n2688# 6.25199f
C12 source a_n1712_n2688# 5.266892f
C13 minus a_n1712_n2688# 6.458999f
C14 plus a_n1712_n2688# 8.094259f
C15 drain_left.t1 a_n1712_n2688# 2.06025f
C16 drain_left.t2 a_n1712_n2688# 0.184725f
C17 drain_left.t9 a_n1712_n2688# 0.184725f
C18 drain_left.n0 a_n1712_n2688# 1.61573f
C19 drain_left.n1 a_n1712_n2688# 0.620815f
C20 drain_left.t4 a_n1712_n2688# 0.184725f
C21 drain_left.t5 a_n1712_n2688# 0.184725f
C22 drain_left.n2 a_n1712_n2688# 1.61806f
C23 drain_left.n3 a_n1712_n2688# 1.38859f
C24 drain_left.t8 a_n1712_n2688# 2.06026f
C25 drain_left.t6 a_n1712_n2688# 0.184725f
C26 drain_left.t0 a_n1712_n2688# 0.184725f
C27 drain_left.n4 a_n1712_n2688# 1.61573f
C28 drain_left.n5 a_n1712_n2688# 0.665479f
C29 drain_left.t7 a_n1712_n2688# 0.184725f
C30 drain_left.t3 a_n1712_n2688# 0.184725f
C31 drain_left.n6 a_n1712_n2688# 1.61573f
C32 drain_left.n7 a_n1712_n2688# 0.550969f
C33 plus.n0 a_n1712_n2688# 0.048475f
C34 plus.t6 a_n1712_n2688# 0.625586f
C35 plus.t2 a_n1712_n2688# 0.625586f
C36 plus.t9 a_n1712_n2688# 0.625586f
C37 plus.n1 a_n1712_n2688# 0.271704f
C38 plus.t1 a_n1712_n2688# 0.636077f
C39 plus.n2 a_n1712_n2688# 0.256486f
C40 plus.t3 a_n1712_n2688# 0.625586f
C41 plus.n3 a_n1712_n2688# 0.269014f
C42 plus.n4 a_n1712_n2688# 0.011f
C43 plus.n5 a_n1712_n2688# 0.154634f
C44 plus.n6 a_n1712_n2688# 0.048475f
C45 plus.n7 a_n1712_n2688# 0.048475f
C46 plus.n8 a_n1712_n2688# 0.011f
C47 plus.n9 a_n1712_n2688# 0.269014f
C48 plus.n10 a_n1712_n2688# 0.266623f
C49 plus.n11 a_n1712_n2688# 0.483562f
C50 plus.n12 a_n1712_n2688# 0.048475f
C51 plus.t8 a_n1712_n2688# 0.625586f
C52 plus.t7 a_n1712_n2688# 0.625586f
C53 plus.t0 a_n1712_n2688# 0.625586f
C54 plus.n13 a_n1712_n2688# 0.271704f
C55 plus.t4 a_n1712_n2688# 0.636077f
C56 plus.n14 a_n1712_n2688# 0.256486f
C57 plus.t5 a_n1712_n2688# 0.625586f
C58 plus.n15 a_n1712_n2688# 0.269014f
C59 plus.n16 a_n1712_n2688# 0.011f
C60 plus.n17 a_n1712_n2688# 0.154634f
C61 plus.n18 a_n1712_n2688# 0.048475f
C62 plus.n19 a_n1712_n2688# 0.048475f
C63 plus.n20 a_n1712_n2688# 0.011f
C64 plus.n21 a_n1712_n2688# 0.269014f
C65 plus.n22 a_n1712_n2688# 0.266623f
C66 plus.n23 a_n1712_n2688# 1.31686f
C67 drain_right.t0 a_n1712_n2688# 2.06044f
C68 drain_right.t1 a_n1712_n2688# 0.184742f
C69 drain_right.t4 a_n1712_n2688# 0.184742f
C70 drain_right.n0 a_n1712_n2688# 1.61588f
C71 drain_right.n1 a_n1712_n2688# 0.620872f
C72 drain_right.t6 a_n1712_n2688# 0.184742f
C73 drain_right.t9 a_n1712_n2688# 0.184742f
C74 drain_right.n2 a_n1712_n2688# 1.61821f
C75 drain_right.n3 a_n1712_n2688# 1.33511f
C76 drain_right.t8 a_n1712_n2688# 0.184742f
C77 drain_right.t3 a_n1712_n2688# 0.184742f
C78 drain_right.n4 a_n1712_n2688# 1.61953f
C79 drain_right.t2 a_n1712_n2688# 0.184742f
C80 drain_right.t5 a_n1712_n2688# 0.184742f
C81 drain_right.n5 a_n1712_n2688# 1.61588f
C82 drain_right.n6 a_n1712_n2688# 0.662504f
C83 drain_right.t7 a_n1712_n2688# 2.05688f
C84 drain_right.n7 a_n1712_n2688# 0.569036f
C85 source.t4 a_n1712_n2688# 2.08651f
C86 source.n0 a_n1712_n2688# 1.22537f
C87 source.t16 a_n1712_n2688# 0.195669f
C88 source.t19 a_n1712_n2688# 0.195669f
C89 source.n1 a_n1712_n2688# 1.63801f
C90 source.n2 a_n1712_n2688# 0.38328f
C91 source.t18 a_n1712_n2688# 0.195669f
C92 source.t1 a_n1712_n2688# 0.195669f
C93 source.n3 a_n1712_n2688# 1.63801f
C94 source.n4 a_n1712_n2688# 0.393215f
C95 source.t9 a_n1712_n2688# 2.08651f
C96 source.n5 a_n1712_n2688# 0.478356f
C97 source.t11 a_n1712_n2688# 0.195669f
C98 source.t8 a_n1712_n2688# 0.195669f
C99 source.n6 a_n1712_n2688# 1.63801f
C100 source.n7 a_n1712_n2688# 0.38328f
C101 source.t7 a_n1712_n2688# 0.195669f
C102 source.t15 a_n1712_n2688# 0.195669f
C103 source.n8 a_n1712_n2688# 1.63801f
C104 source.n9 a_n1712_n2688# 1.6084f
C105 source.t3 a_n1712_n2688# 0.195669f
C106 source.t5 a_n1712_n2688# 0.195669f
C107 source.n10 a_n1712_n2688# 1.63801f
C108 source.n11 a_n1712_n2688# 1.60841f
C109 source.t17 a_n1712_n2688# 0.195669f
C110 source.t2 a_n1712_n2688# 0.195669f
C111 source.n12 a_n1712_n2688# 1.63801f
C112 source.n13 a_n1712_n2688# 0.383285f
C113 source.t0 a_n1712_n2688# 2.08651f
C114 source.n14 a_n1712_n2688# 0.478361f
C115 source.t13 a_n1712_n2688# 0.195669f
C116 source.t12 a_n1712_n2688# 0.195669f
C117 source.n15 a_n1712_n2688# 1.63801f
C118 source.n16 a_n1712_n2688# 0.39322f
C119 source.t14 a_n1712_n2688# 0.195669f
C120 source.t10 a_n1712_n2688# 0.195669f
C121 source.n17 a_n1712_n2688# 1.63801f
C122 source.n18 a_n1712_n2688# 0.383285f
C123 source.t6 a_n1712_n2688# 2.08651f
C124 source.n19 a_n1712_n2688# 0.614098f
C125 source.n20 a_n1712_n2688# 1.44034f
C126 minus.n0 a_n1712_n2688# 0.047753f
C127 minus.t4 a_n1712_n2688# 0.61627f
C128 minus.n1 a_n1712_n2688# 0.267658f
C129 minus.t6 a_n1712_n2688# 0.626605f
C130 minus.n2 a_n1712_n2688# 0.252666f
C131 minus.t1 a_n1712_n2688# 0.61627f
C132 minus.n3 a_n1712_n2688# 0.265008f
C133 minus.n4 a_n1712_n2688# 0.010836f
C134 minus.n5 a_n1712_n2688# 0.152331f
C135 minus.n6 a_n1712_n2688# 0.047753f
C136 minus.n7 a_n1712_n2688# 0.047753f
C137 minus.n8 a_n1712_n2688# 0.010836f
C138 minus.t7 a_n1712_n2688# 0.61627f
C139 minus.n9 a_n1712_n2688# 0.265008f
C140 minus.t2 a_n1712_n2688# 0.61627f
C141 minus.n10 a_n1712_n2688# 0.262652f
C142 minus.n11 a_n1712_n2688# 1.48734f
C143 minus.n12 a_n1712_n2688# 0.047753f
C144 minus.t5 a_n1712_n2688# 0.61627f
C145 minus.n13 a_n1712_n2688# 0.267658f
C146 minus.t9 a_n1712_n2688# 0.626605f
C147 minus.n14 a_n1712_n2688# 0.252666f
C148 minus.t8 a_n1712_n2688# 0.61627f
C149 minus.n15 a_n1712_n2688# 0.265008f
C150 minus.n16 a_n1712_n2688# 0.010836f
C151 minus.n17 a_n1712_n2688# 0.152331f
C152 minus.n18 a_n1712_n2688# 0.047753f
C153 minus.n19 a_n1712_n2688# 0.047753f
C154 minus.n20 a_n1712_n2688# 0.010836f
C155 minus.t3 a_n1712_n2688# 0.61627f
C156 minus.n21 a_n1712_n2688# 0.265008f
C157 minus.t0 a_n1712_n2688# 0.61627f
C158 minus.n22 a_n1712_n2688# 0.262652f
C159 minus.n23 a_n1712_n2688# 0.319263f
C160 minus.n24 a_n1712_n2688# 1.81816f
.ends

