* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X2 drain_right.t5 minus.t0 source.t7 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X3 drain_left.t5 plus.t0 source.t4 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X4 a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X5 source.t5 plus.t1 drain_left.t4 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right.t4 minus.t1 source.t6 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X7 source.t8 minus.t2 drain_right.t3 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X8 drain_left.t3 plus.t2 source.t0 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X9 drain_right.t2 minus.t3 source.t11 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X10 drain_right.t1 minus.t4 source.t10 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X11 source.t1 plus.t3 drain_left.t2 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X12 drain_left.t1 plus.t4 source.t3 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X13 a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X14 source.t9 minus.t5 drain_right.t0 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 drain_left.t0 plus.t5 source.t2 a_n1460_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
R0 minus.n0 minus.t3 172.626
R1 minus.n4 minus.t0 172.626
R2 minus.n3 minus.n2 161.3
R3 minus.n7 minus.n6 161.3
R4 minus.n1 minus.t2 145.805
R5 minus.n2 minus.t1 145.805
R6 minus.n5 minus.t5 145.805
R7 minus.n6 minus.t4 145.805
R8 minus.n2 minus.n1 48.2005
R9 minus.n6 minus.n5 48.2005
R10 minus.n3 minus.n0 45.1367
R11 minus.n7 minus.n4 45.1367
R12 minus.n8 minus.n3 27.2032
R13 minus.n1 minus.n0 13.3799
R14 minus.n5 minus.n4 13.3799
R15 minus.n8 minus.n7 6.62739
R16 minus minus.n8 0.188
R17 source.n34 source.n32 289.615
R18 source.n24 source.n22 289.615
R19 source.n2 source.n0 289.615
R20 source.n12 source.n10 289.615
R21 source.n35 source.n34 185
R22 source.n25 source.n24 185
R23 source.n3 source.n2 185
R24 source.n13 source.n12 185
R25 source.t10 source.n33 167.117
R26 source.t2 source.n23 167.117
R27 source.t0 source.n1 167.117
R28 source.t11 source.n11 167.117
R29 source.n9 source.n8 84.1169
R30 source.n19 source.n18 84.1169
R31 source.n31 source.n30 84.1168
R32 source.n21 source.n20 84.1168
R33 source.n34 source.t10 52.3082
R34 source.n24 source.t2 52.3082
R35 source.n2 source.t0 52.3082
R36 source.n12 source.t11 52.3082
R37 source.n39 source.n38 31.4096
R38 source.n29 source.n28 31.4096
R39 source.n7 source.n6 31.4096
R40 source.n17 source.n16 31.4096
R41 source.n21 source.n19 15.3154
R42 source.n30 source.t7 9.9005
R43 source.n30 source.t9 9.9005
R44 source.n20 source.t4 9.9005
R45 source.n20 source.t5 9.9005
R46 source.n8 source.t3 9.9005
R47 source.n8 source.t1 9.9005
R48 source.n18 source.t6 9.9005
R49 source.n18 source.t8 9.9005
R50 source.n35 source.n33 9.71174
R51 source.n25 source.n23 9.71174
R52 source.n3 source.n1 9.71174
R53 source.n13 source.n11 9.71174
R54 source.n38 source.n37 9.45567
R55 source.n28 source.n27 9.45567
R56 source.n6 source.n5 9.45567
R57 source.n16 source.n15 9.45567
R58 source.n37 source.n36 9.3005
R59 source.n27 source.n26 9.3005
R60 source.n5 source.n4 9.3005
R61 source.n15 source.n14 9.3005
R62 source.n40 source.n7 8.8499
R63 source.n38 source.n32 8.14595
R64 source.n28 source.n22 8.14595
R65 source.n6 source.n0 8.14595
R66 source.n16 source.n10 8.14595
R67 source.n36 source.n35 7.3702
R68 source.n26 source.n25 7.3702
R69 source.n4 source.n3 7.3702
R70 source.n14 source.n13 7.3702
R71 source.n36 source.n32 5.81868
R72 source.n26 source.n22 5.81868
R73 source.n4 source.n0 5.81868
R74 source.n14 source.n10 5.81868
R75 source.n40 source.n39 5.66429
R76 source.n37 source.n33 3.44771
R77 source.n27 source.n23 3.44771
R78 source.n5 source.n1 3.44771
R79 source.n15 source.n11 3.44771
R80 source.n17 source.n9 0.87119
R81 source.n31 source.n29 0.87119
R82 source.n19 source.n17 0.802224
R83 source.n9 source.n7 0.802224
R84 source.n29 source.n21 0.802224
R85 source.n39 source.n31 0.802224
R86 source source.n40 0.188
R87 drain_right.n2 drain_right.n0 289.615
R88 drain_right.n12 drain_right.n10 289.615
R89 drain_right.n3 drain_right.n2 185
R90 drain_right.n13 drain_right.n12 185
R91 drain_right.t5 drain_right.n1 167.117
R92 drain_right.t4 drain_right.n11 167.117
R93 drain_right.n17 drain_right.n9 101.597
R94 drain_right.n8 drain_right.n7 100.941
R95 drain_right.n2 drain_right.t5 52.3082
R96 drain_right.n12 drain_right.t4 52.3082
R97 drain_right.n8 drain_right.n6 48.6343
R98 drain_right.n17 drain_right.n16 48.0884
R99 drain_right drain_right.n8 21.4428
R100 drain_right.n7 drain_right.t0 9.9005
R101 drain_right.n7 drain_right.t1 9.9005
R102 drain_right.n9 drain_right.t3 9.9005
R103 drain_right.n9 drain_right.t2 9.9005
R104 drain_right.n3 drain_right.n1 9.71174
R105 drain_right.n13 drain_right.n11 9.71174
R106 drain_right.n6 drain_right.n5 9.45567
R107 drain_right.n16 drain_right.n15 9.45567
R108 drain_right.n5 drain_right.n4 9.3005
R109 drain_right.n15 drain_right.n14 9.3005
R110 drain_right.n6 drain_right.n0 8.14595
R111 drain_right.n16 drain_right.n10 8.14595
R112 drain_right.n4 drain_right.n3 7.3702
R113 drain_right.n14 drain_right.n13 7.3702
R114 drain_right drain_right.n17 6.05408
R115 drain_right.n4 drain_right.n0 5.81868
R116 drain_right.n14 drain_right.n10 5.81868
R117 drain_right.n5 drain_right.n1 3.44771
R118 drain_right.n15 drain_right.n11 3.44771
R119 plus.n0 plus.t4 172.626
R120 plus.n4 plus.t5 172.626
R121 plus.n3 plus.n2 161.3
R122 plus.n7 plus.n6 161.3
R123 plus.n2 plus.t2 145.805
R124 plus.n1 plus.t3 145.805
R125 plus.n6 plus.t0 145.805
R126 plus.n5 plus.t1 145.805
R127 plus.n2 plus.n1 48.2005
R128 plus.n6 plus.n5 48.2005
R129 plus.n3 plus.n0 45.1367
R130 plus.n7 plus.n4 45.1367
R131 plus plus.n7 24.8721
R132 plus.n1 plus.n0 13.3799
R133 plus.n5 plus.n4 13.3799
R134 plus plus.n3 8.48345
R135 drain_left.n2 drain_left.n0 289.615
R136 drain_left.n11 drain_left.n9 289.615
R137 drain_left.n3 drain_left.n2 185
R138 drain_left.n12 drain_left.n11 185
R139 drain_left.t5 drain_left.n1 167.117
R140 drain_left.t1 drain_left.n10 167.117
R141 drain_left.n8 drain_left.n7 100.941
R142 drain_left.n17 drain_left.n16 100.796
R143 drain_left.n2 drain_left.t5 52.3082
R144 drain_left.n11 drain_left.t1 52.3082
R145 drain_left.n17 drain_left.n15 48.8901
R146 drain_left.n8 drain_left.n6 48.6343
R147 drain_left drain_left.n8 21.9961
R148 drain_left.n7 drain_left.t4 9.9005
R149 drain_left.n7 drain_left.t0 9.9005
R150 drain_left.n16 drain_left.t2 9.9005
R151 drain_left.n16 drain_left.t3 9.9005
R152 drain_left.n3 drain_left.n1 9.71174
R153 drain_left.n12 drain_left.n10 9.71174
R154 drain_left.n6 drain_left.n5 9.45567
R155 drain_left.n15 drain_left.n14 9.45567
R156 drain_left.n5 drain_left.n4 9.3005
R157 drain_left.n14 drain_left.n13 9.3005
R158 drain_left.n6 drain_left.n0 8.14595
R159 drain_left.n15 drain_left.n9 8.14595
R160 drain_left.n4 drain_left.n3 7.3702
R161 drain_left.n13 drain_left.n12 7.3702
R162 drain_left drain_left.n17 6.45494
R163 drain_left.n4 drain_left.n0 5.81868
R164 drain_left.n13 drain_left.n9 5.81868
R165 drain_left.n5 drain_left.n1 3.44771
R166 drain_left.n14 drain_left.n10 3.44771
C0 drain_right minus 0.946846f
C1 drain_right source 3.32086f
C2 drain_left drain_right 0.671331f
C3 minus source 1.11179f
C4 drain_left minus 0.177626f
C5 drain_left source 3.32226f
C6 plus drain_right 0.300636f
C7 plus minus 3.11697f
C8 plus source 1.12584f
C9 plus drain_left 1.08543f
C10 drain_right a_n1460_n1288# 3.16395f
C11 drain_left a_n1460_n1288# 3.35767f
C12 source a_n1460_n1288# 2.448311f
C13 minus a_n1460_n1288# 4.768833f
C14 plus a_n1460_n1288# 5.394262f
C15 drain_left.n0 a_n1460_n1288# 0.026018f
C16 drain_left.n1 a_n1460_n1288# 0.057567f
C17 drain_left.t5 a_n1460_n1288# 0.043201f
C18 drain_left.n2 a_n1460_n1288# 0.045054f
C19 drain_left.n3 a_n1460_n1288# 0.014524f
C20 drain_left.n4 a_n1460_n1288# 0.009579f
C21 drain_left.n5 a_n1460_n1288# 0.126892f
C22 drain_left.n6 a_n1460_n1288# 0.041577f
C23 drain_left.t4 a_n1460_n1288# 0.028173f
C24 drain_left.t0 a_n1460_n1288# 0.028173f
C25 drain_left.n7 a_n1460_n1288# 0.177278f
C26 drain_left.n8 a_n1460_n1288# 0.718479f
C27 drain_left.n9 a_n1460_n1288# 0.026018f
C28 drain_left.n10 a_n1460_n1288# 0.057567f
C29 drain_left.t1 a_n1460_n1288# 0.043201f
C30 drain_left.n11 a_n1460_n1288# 0.045054f
C31 drain_left.n12 a_n1460_n1288# 0.014524f
C32 drain_left.n13 a_n1460_n1288# 0.009579f
C33 drain_left.n14 a_n1460_n1288# 0.126892f
C34 drain_left.n15 a_n1460_n1288# 0.042146f
C35 drain_left.t2 a_n1460_n1288# 0.028173f
C36 drain_left.t3 a_n1460_n1288# 0.028173f
C37 drain_left.n16 a_n1460_n1288# 0.17699f
C38 drain_left.n17 a_n1460_n1288# 0.462479f
C39 plus.t4 a_n1460_n1288# 0.128277f
C40 plus.n0 a_n1460_n1288# 0.069763f
C41 plus.t2 a_n1460_n1288# 0.11555f
C42 plus.t3 a_n1460_n1288# 0.11555f
C43 plus.n1 a_n1460_n1288# 0.08888f
C44 plus.n2 a_n1460_n1288# 0.081824f
C45 plus.n3 a_n1460_n1288# 0.333512f
C46 plus.t5 a_n1460_n1288# 0.128277f
C47 plus.n4 a_n1460_n1288# 0.069763f
C48 plus.t0 a_n1460_n1288# 0.11555f
C49 plus.t1 a_n1460_n1288# 0.11555f
C50 plus.n5 a_n1460_n1288# 0.08888f
C51 plus.n6 a_n1460_n1288# 0.081824f
C52 plus.n7 a_n1460_n1288# 0.758931f
C53 drain_right.n0 a_n1460_n1288# 0.026579f
C54 drain_right.n1 a_n1460_n1288# 0.05881f
C55 drain_right.t5 a_n1460_n1288# 0.044134f
C56 drain_right.n2 a_n1460_n1288# 0.046027f
C57 drain_right.n3 a_n1460_n1288# 0.014837f
C58 drain_right.n4 a_n1460_n1288# 0.009785f
C59 drain_right.n5 a_n1460_n1288# 0.129631f
C60 drain_right.n6 a_n1460_n1288# 0.042475f
C61 drain_right.t0 a_n1460_n1288# 0.028781f
C62 drain_right.t1 a_n1460_n1288# 0.028781f
C63 drain_right.n7 a_n1460_n1288# 0.181105f
C64 drain_right.n8 a_n1460_n1288# 0.698166f
C65 drain_right.t3 a_n1460_n1288# 0.028781f
C66 drain_right.t2 a_n1460_n1288# 0.028781f
C67 drain_right.n9 a_n1460_n1288# 0.182711f
C68 drain_right.n10 a_n1460_n1288# 0.026579f
C69 drain_right.n11 a_n1460_n1288# 0.05881f
C70 drain_right.t4 a_n1460_n1288# 0.044134f
C71 drain_right.n12 a_n1460_n1288# 0.046027f
C72 drain_right.n13 a_n1460_n1288# 0.014837f
C73 drain_right.n14 a_n1460_n1288# 0.009785f
C74 drain_right.n15 a_n1460_n1288# 0.129631f
C75 drain_right.n16 a_n1460_n1288# 0.041719f
C76 drain_right.n17 a_n1460_n1288# 0.483973f
C77 source.n0 a_n1460_n1288# 0.033235f
C78 source.n1 a_n1460_n1288# 0.073536f
C79 source.t0 a_n1460_n1288# 0.055185f
C80 source.n2 a_n1460_n1288# 0.057552f
C81 source.n3 a_n1460_n1288# 0.018553f
C82 source.n4 a_n1460_n1288# 0.012236f
C83 source.n5 a_n1460_n1288# 0.162091f
C84 source.n6 a_n1460_n1288# 0.036433f
C85 source.n7 a_n1460_n1288# 0.37744f
C86 source.t3 a_n1460_n1288# 0.035988f
C87 source.t1 a_n1460_n1288# 0.035988f
C88 source.n8 a_n1460_n1288# 0.192389f
C89 source.n9 a_n1460_n1288# 0.299736f
C90 source.n10 a_n1460_n1288# 0.033235f
C91 source.n11 a_n1460_n1288# 0.073536f
C92 source.t11 a_n1460_n1288# 0.055185f
C93 source.n12 a_n1460_n1288# 0.057552f
C94 source.n13 a_n1460_n1288# 0.018553f
C95 source.n14 a_n1460_n1288# 0.012236f
C96 source.n15 a_n1460_n1288# 0.162091f
C97 source.n16 a_n1460_n1288# 0.036433f
C98 source.n17 a_n1460_n1288# 0.141453f
C99 source.t6 a_n1460_n1288# 0.035988f
C100 source.t8 a_n1460_n1288# 0.035988f
C101 source.n18 a_n1460_n1288# 0.192389f
C102 source.n19 a_n1460_n1288# 0.811142f
C103 source.t4 a_n1460_n1288# 0.035988f
C104 source.t5 a_n1460_n1288# 0.035988f
C105 source.n20 a_n1460_n1288# 0.192388f
C106 source.n21 a_n1460_n1288# 0.811143f
C107 source.n22 a_n1460_n1288# 0.033235f
C108 source.n23 a_n1460_n1288# 0.073536f
C109 source.t2 a_n1460_n1288# 0.055185f
C110 source.n24 a_n1460_n1288# 0.057552f
C111 source.n25 a_n1460_n1288# 0.018553f
C112 source.n26 a_n1460_n1288# 0.012236f
C113 source.n27 a_n1460_n1288# 0.162091f
C114 source.n28 a_n1460_n1288# 0.036433f
C115 source.n29 a_n1460_n1288# 0.141453f
C116 source.t7 a_n1460_n1288# 0.035988f
C117 source.t9 a_n1460_n1288# 0.035988f
C118 source.n30 a_n1460_n1288# 0.192388f
C119 source.n31 a_n1460_n1288# 0.299737f
C120 source.n32 a_n1460_n1288# 0.033235f
C121 source.n33 a_n1460_n1288# 0.073536f
C122 source.t10 a_n1460_n1288# 0.055185f
C123 source.n34 a_n1460_n1288# 0.057552f
C124 source.n35 a_n1460_n1288# 0.018553f
C125 source.n36 a_n1460_n1288# 0.012236f
C126 source.n37 a_n1460_n1288# 0.162091f
C127 source.n38 a_n1460_n1288# 0.036433f
C128 source.n39 a_n1460_n1288# 0.255616f
C129 source.n40 a_n1460_n1288# 0.57121f
C130 minus.t3 a_n1460_n1288# 0.125726f
C131 minus.n0 a_n1460_n1288# 0.068376f
C132 minus.t2 a_n1460_n1288# 0.113253f
C133 minus.n1 a_n1460_n1288# 0.087113f
C134 minus.t1 a_n1460_n1288# 0.113253f
C135 minus.n2 a_n1460_n1288# 0.080197f
C136 minus.n3 a_n1460_n1288# 0.771301f
C137 minus.t0 a_n1460_n1288# 0.125726f
C138 minus.n4 a_n1460_n1288# 0.068376f
C139 minus.t5 a_n1460_n1288# 0.113253f
C140 minus.n5 a_n1460_n1288# 0.087113f
C141 minus.t4 a_n1460_n1288# 0.113253f
C142 minus.n6 a_n1460_n1288# 0.080197f
C143 minus.n7 a_n1460_n1288# 0.307759f
C144 minus.n8 a_n1460_n1288# 0.825093f
.ends

