* NGSPICE file created from diffpair49.ext - technology: sky130A

.subckt diffpair49 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t38 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X1 source.t34 plus.t1 drain_left.t22 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 drain_right.t23 minus.t0 source.t13 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_left.t21 plus.t2 source.t45 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X5 source.t40 plus.t3 drain_left.t20 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X6 source.t19 minus.t1 drain_right.t22 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 drain_right.t21 minus.t2 source.t2 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 source.t35 plus.t4 drain_left.t19 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 source.t27 plus.t5 drain_left.t18 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 source.t33 plus.t6 drain_left.t17 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X11 source.t23 minus.t3 drain_right.t20 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X13 a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X14 drain_right.t19 minus.t4 source.t18 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X15 source.t25 plus.t7 drain_left.t16 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 drain_right.t18 minus.t5 source.t9 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 drain_right.t17 minus.t6 source.t17 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 source.t22 minus.t7 drain_right.t16 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 drain_right.t15 minus.t8 source.t6 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X20 drain_left.t15 plus.t8 source.t28 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X21 drain_left.t14 plus.t9 source.t30 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 source.t21 minus.t9 drain_right.t14 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X23 source.t31 plus.t10 drain_left.t13 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X24 source.t8 minus.t10 drain_right.t13 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 drain_right.t12 minus.t11 source.t12 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 source.t16 minus.t12 drain_right.t11 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 drain_left.t12 plus.t11 source.t26 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X28 source.t5 minus.t13 drain_right.t10 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 drain_left.t11 plus.t12 source.t32 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 drain_left.t10 plus.t13 source.t43 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 drain_right.t9 minus.t14 source.t1 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X32 drain_right.t8 minus.t15 source.t4 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X33 a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X34 drain_right.t7 minus.t16 source.t7 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X35 drain_right.t6 minus.t17 source.t11 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X36 drain_left.t9 plus.t14 source.t42 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X37 drain_right.t5 minus.t18 source.t15 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X38 source.t0 minus.t19 drain_right.t4 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X39 source.t44 plus.t15 drain_left.t8 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X40 source.t47 plus.t16 drain_left.t7 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X41 source.t20 minus.t20 drain_right.t3 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X42 source.t29 plus.t17 drain_left.t6 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X43 source.t24 plus.t18 drain_left.t5 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X44 source.t3 minus.t21 drain_right.t2 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X45 drain_left.t4 plus.t19 source.t36 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X46 source.t10 minus.t22 drain_right.t1 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X47 drain_left.t3 plus.t20 source.t46 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X48 source.t37 plus.t21 drain_left.t2 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X49 source.t14 minus.t23 drain_right.t0 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X50 drain_left.t1 plus.t22 source.t39 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X51 drain_left.t0 plus.t23 source.t41 a_n2874_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
R0 plus.n12 plus.n9 161.3
R1 plus.n14 plus.n13 161.3
R2 plus.n15 plus.n8 161.3
R3 plus.n16 plus.n7 161.3
R4 plus.n18 plus.n17 161.3
R5 plus.n19 plus.n6 161.3
R6 plus.n21 plus.n20 161.3
R7 plus.n22 plus.n5 161.3
R8 plus.n23 plus.n4 161.3
R9 plus.n25 plus.n24 161.3
R10 plus.n26 plus.n3 161.3
R11 plus.n28 plus.n27 161.3
R12 plus.n29 plus.n2 161.3
R13 plus.n30 plus.n1 161.3
R14 plus.n31 plus.n0 161.3
R15 plus.n33 plus.n32 161.3
R16 plus.n46 plus.n43 161.3
R17 plus.n48 plus.n47 161.3
R18 plus.n49 plus.n42 161.3
R19 plus.n50 plus.n41 161.3
R20 plus.n52 plus.n51 161.3
R21 plus.n53 plus.n40 161.3
R22 plus.n55 plus.n54 161.3
R23 plus.n56 plus.n39 161.3
R24 plus.n57 plus.n38 161.3
R25 plus.n59 plus.n58 161.3
R26 plus.n60 plus.n37 161.3
R27 plus.n62 plus.n61 161.3
R28 plus.n63 plus.n36 161.3
R29 plus.n64 plus.n35 161.3
R30 plus.n65 plus.n34 161.3
R31 plus.n67 plus.n66 161.3
R32 plus.n11 plus.t6 153.125
R33 plus.n45 plus.t11 153.125
R34 plus.n32 plus.t2 126.766
R35 plus.n30 plus.t3 126.766
R36 plus.n29 plus.t13 126.766
R37 plus.n3 plus.t5 126.766
R38 plus.n23 plus.t20 126.766
R39 plus.n22 plus.t10 126.766
R40 plus.n6 plus.t23 126.766
R41 plus.n17 plus.t18 126.766
R42 plus.n15 plus.t8 126.766
R43 plus.n9 plus.t21 126.766
R44 plus.n10 plus.t14 126.766
R45 plus.n66 plus.t1 126.766
R46 plus.n64 plus.t12 126.766
R47 plus.n63 plus.t4 126.766
R48 plus.n37 plus.t22 126.766
R49 plus.n57 plus.t7 126.766
R50 plus.n56 plus.t19 126.766
R51 plus.n40 plus.t16 126.766
R52 plus.n51 plus.t0 126.766
R53 plus.n49 plus.t17 126.766
R54 plus.n43 plus.t9 126.766
R55 plus.n44 plus.t15 126.766
R56 plus.n30 plus.n29 48.2005
R57 plus.n23 plus.n22 48.2005
R58 plus.n17 plus.n6 48.2005
R59 plus.n10 plus.n9 48.2005
R60 plus.n64 plus.n63 48.2005
R61 plus.n57 plus.n56 48.2005
R62 plus.n51 plus.n40 48.2005
R63 plus.n44 plus.n43 48.2005
R64 plus.n24 plus.n3 47.4702
R65 plus.n16 plus.n15 47.4702
R66 plus.n58 plus.n37 47.4702
R67 plus.n50 plus.n49 47.4702
R68 plus.n32 plus.n31 46.0096
R69 plus.n66 plus.n65 46.0096
R70 plus.n12 plus.n11 45.0871
R71 plus.n46 plus.n45 45.0871
R72 plus plus.n67 29.749
R73 plus.n28 plus.n3 25.5611
R74 plus.n15 plus.n14 25.5611
R75 plus.n62 plus.n37 25.5611
R76 plus.n49 plus.n48 25.5611
R77 plus.n21 plus.n6 24.1005
R78 plus.n22 plus.n21 24.1005
R79 plus.n56 plus.n55 24.1005
R80 plus.n55 plus.n40 24.1005
R81 plus.n29 plus.n28 22.6399
R82 plus.n14 plus.n9 22.6399
R83 plus.n63 plus.n62 22.6399
R84 plus.n48 plus.n43 22.6399
R85 plus.n11 plus.n10 14.1472
R86 plus.n45 plus.n44 14.1472
R87 plus plus.n33 8.00429
R88 plus.n31 plus.n30 2.19141
R89 plus.n65 plus.n64 2.19141
R90 plus.n24 plus.n23 0.730803
R91 plus.n17 plus.n16 0.730803
R92 plus.n58 plus.n57 0.730803
R93 plus.n51 plus.n50 0.730803
R94 plus.n13 plus.n12 0.189894
R95 plus.n13 plus.n8 0.189894
R96 plus.n8 plus.n7 0.189894
R97 plus.n18 plus.n7 0.189894
R98 plus.n19 plus.n18 0.189894
R99 plus.n20 plus.n19 0.189894
R100 plus.n20 plus.n5 0.189894
R101 plus.n5 plus.n4 0.189894
R102 plus.n25 plus.n4 0.189894
R103 plus.n26 plus.n25 0.189894
R104 plus.n27 plus.n26 0.189894
R105 plus.n27 plus.n2 0.189894
R106 plus.n2 plus.n1 0.189894
R107 plus.n1 plus.n0 0.189894
R108 plus.n33 plus.n0 0.189894
R109 plus.n67 plus.n34 0.189894
R110 plus.n35 plus.n34 0.189894
R111 plus.n36 plus.n35 0.189894
R112 plus.n61 plus.n36 0.189894
R113 plus.n61 plus.n60 0.189894
R114 plus.n60 plus.n59 0.189894
R115 plus.n59 plus.n38 0.189894
R116 plus.n39 plus.n38 0.189894
R117 plus.n54 plus.n39 0.189894
R118 plus.n54 plus.n53 0.189894
R119 plus.n53 plus.n52 0.189894
R120 plus.n52 plus.n41 0.189894
R121 plus.n42 plus.n41 0.189894
R122 plus.n47 plus.n42 0.189894
R123 plus.n47 plus.n46 0.189894
R124 source.n0 source.t45 243.255
R125 source.n11 source.t33 243.255
R126 source.n12 source.t1 243.255
R127 source.n23 source.t10 243.255
R128 source.n47 source.t6 243.254
R129 source.n36 source.t21 243.254
R130 source.n35 source.t26 243.254
R131 source.n24 source.t34 243.254
R132 source.n2 source.n1 223.454
R133 source.n4 source.n3 223.454
R134 source.n6 source.n5 223.454
R135 source.n8 source.n7 223.454
R136 source.n10 source.n9 223.454
R137 source.n14 source.n13 223.454
R138 source.n16 source.n15 223.454
R139 source.n18 source.n17 223.454
R140 source.n20 source.n19 223.454
R141 source.n22 source.n21 223.454
R142 source.n46 source.n45 223.453
R143 source.n44 source.n43 223.453
R144 source.n42 source.n41 223.453
R145 source.n40 source.n39 223.453
R146 source.n38 source.n37 223.453
R147 source.n34 source.n33 223.453
R148 source.n32 source.n31 223.453
R149 source.n30 source.n29 223.453
R150 source.n28 source.n27 223.453
R151 source.n26 source.n25 223.453
R152 source.n45 source.t2 19.8005
R153 source.n45 source.t5 19.8005
R154 source.n43 source.t9 19.8005
R155 source.n43 source.t0 19.8005
R156 source.n41 source.t11 19.8005
R157 source.n41 source.t3 19.8005
R158 source.n39 source.t12 19.8005
R159 source.n39 source.t14 19.8005
R160 source.n37 source.t7 19.8005
R161 source.n37 source.t22 19.8005
R162 source.n33 source.t30 19.8005
R163 source.n33 source.t44 19.8005
R164 source.n31 source.t38 19.8005
R165 source.n31 source.t29 19.8005
R166 source.n29 source.t36 19.8005
R167 source.n29 source.t47 19.8005
R168 source.n27 source.t39 19.8005
R169 source.n27 source.t25 19.8005
R170 source.n25 source.t32 19.8005
R171 source.n25 source.t35 19.8005
R172 source.n1 source.t43 19.8005
R173 source.n1 source.t40 19.8005
R174 source.n3 source.t46 19.8005
R175 source.n3 source.t27 19.8005
R176 source.n5 source.t41 19.8005
R177 source.n5 source.t31 19.8005
R178 source.n7 source.t28 19.8005
R179 source.n7 source.t24 19.8005
R180 source.n9 source.t42 19.8005
R181 source.n9 source.t37 19.8005
R182 source.n13 source.t17 19.8005
R183 source.n13 source.t19 19.8005
R184 source.n15 source.t18 19.8005
R185 source.n15 source.t20 19.8005
R186 source.n17 source.t13 19.8005
R187 source.n17 source.t8 19.8005
R188 source.n19 source.t15 19.8005
R189 source.n19 source.t16 19.8005
R190 source.n21 source.t4 19.8005
R191 source.n21 source.t23 19.8005
R192 source.n24 source.n23 13.6699
R193 source.n48 source.n0 8.04922
R194 source.n48 source.n47 5.62119
R195 source.n23 source.n22 0.716017
R196 source.n22 source.n20 0.716017
R197 source.n20 source.n18 0.716017
R198 source.n18 source.n16 0.716017
R199 source.n16 source.n14 0.716017
R200 source.n14 source.n12 0.716017
R201 source.n11 source.n10 0.716017
R202 source.n10 source.n8 0.716017
R203 source.n8 source.n6 0.716017
R204 source.n6 source.n4 0.716017
R205 source.n4 source.n2 0.716017
R206 source.n2 source.n0 0.716017
R207 source.n26 source.n24 0.716017
R208 source.n28 source.n26 0.716017
R209 source.n30 source.n28 0.716017
R210 source.n32 source.n30 0.716017
R211 source.n34 source.n32 0.716017
R212 source.n35 source.n34 0.716017
R213 source.n38 source.n36 0.716017
R214 source.n40 source.n38 0.716017
R215 source.n42 source.n40 0.716017
R216 source.n44 source.n42 0.716017
R217 source.n46 source.n44 0.716017
R218 source.n47 source.n46 0.716017
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 240.849
R223 drain_left.n7 drain_left.n5 240.847
R224 drain_left.n2 drain_left.n0 240.847
R225 drain_left.n21 drain_left.n20 240.132
R226 drain_left.n19 drain_left.n18 240.132
R227 drain_left.n17 drain_left.n16 240.132
R228 drain_left.n15 drain_left.n14 240.132
R229 drain_left.n13 drain_left.n12 240.132
R230 drain_left.n7 drain_left.n6 240.131
R231 drain_left.n9 drain_left.n8 240.131
R232 drain_left.n4 drain_left.n3 240.131
R233 drain_left.n2 drain_left.n1 240.131
R234 drain_left drain_left.n10 25.8312
R235 drain_left.n5 drain_left.t8 19.8005
R236 drain_left.n5 drain_left.t12 19.8005
R237 drain_left.n6 drain_left.t6 19.8005
R238 drain_left.n6 drain_left.t14 19.8005
R239 drain_left.n8 drain_left.t7 19.8005
R240 drain_left.n8 drain_left.t23 19.8005
R241 drain_left.n3 drain_left.t16 19.8005
R242 drain_left.n3 drain_left.t4 19.8005
R243 drain_left.n1 drain_left.t19 19.8005
R244 drain_left.n1 drain_left.t1 19.8005
R245 drain_left.n0 drain_left.t22 19.8005
R246 drain_left.n0 drain_left.t11 19.8005
R247 drain_left.n20 drain_left.t20 19.8005
R248 drain_left.n20 drain_left.t21 19.8005
R249 drain_left.n18 drain_left.t18 19.8005
R250 drain_left.n18 drain_left.t10 19.8005
R251 drain_left.n16 drain_left.t13 19.8005
R252 drain_left.n16 drain_left.t3 19.8005
R253 drain_left.n14 drain_left.t5 19.8005
R254 drain_left.n14 drain_left.t0 19.8005
R255 drain_left.n12 drain_left.t2 19.8005
R256 drain_left.n12 drain_left.t15 19.8005
R257 drain_left.n11 drain_left.t17 19.8005
R258 drain_left.n11 drain_left.t9 19.8005
R259 drain_left drain_left.n21 6.36873
R260 drain_left.n9 drain_left.n7 0.716017
R261 drain_left.n4 drain_left.n2 0.716017
R262 drain_left.n15 drain_left.n13 0.716017
R263 drain_left.n17 drain_left.n15 0.716017
R264 drain_left.n19 drain_left.n17 0.716017
R265 drain_left.n21 drain_left.n19 0.716017
R266 drain_left.n10 drain_left.n9 0.302913
R267 drain_left.n10 drain_left.n4 0.302913
R268 minus.n33 minus.n32 161.3
R269 minus.n31 minus.n0 161.3
R270 minus.n30 minus.n29 161.3
R271 minus.n28 minus.n1 161.3
R272 minus.n27 minus.n26 161.3
R273 minus.n25 minus.n2 161.3
R274 minus.n24 minus.n23 161.3
R275 minus.n22 minus.n3 161.3
R276 minus.n21 minus.n20 161.3
R277 minus.n19 minus.n4 161.3
R278 minus.n18 minus.n17 161.3
R279 minus.n16 minus.n5 161.3
R280 minus.n15 minus.n14 161.3
R281 minus.n13 minus.n6 161.3
R282 minus.n12 minus.n11 161.3
R283 minus.n10 minus.n7 161.3
R284 minus.n67 minus.n66 161.3
R285 minus.n65 minus.n34 161.3
R286 minus.n64 minus.n63 161.3
R287 minus.n62 minus.n35 161.3
R288 minus.n61 minus.n60 161.3
R289 minus.n59 minus.n36 161.3
R290 minus.n58 minus.n57 161.3
R291 minus.n56 minus.n37 161.3
R292 minus.n55 minus.n54 161.3
R293 minus.n53 minus.n38 161.3
R294 minus.n52 minus.n51 161.3
R295 minus.n50 minus.n39 161.3
R296 minus.n49 minus.n48 161.3
R297 minus.n47 minus.n40 161.3
R298 minus.n46 minus.n45 161.3
R299 minus.n44 minus.n41 161.3
R300 minus.n9 minus.t14 153.125
R301 minus.n43 minus.t9 153.125
R302 minus.n8 minus.t1 126.766
R303 minus.n7 minus.t6 126.766
R304 minus.n13 minus.t20 126.766
R305 minus.n5 minus.t4 126.766
R306 minus.n18 minus.t10 126.766
R307 minus.n20 minus.t0 126.766
R308 minus.n3 minus.t12 126.766
R309 minus.n25 minus.t18 126.766
R310 minus.n1 minus.t3 126.766
R311 minus.n30 minus.t15 126.766
R312 minus.n32 minus.t22 126.766
R313 minus.n42 minus.t16 126.766
R314 minus.n41 minus.t7 126.766
R315 minus.n47 minus.t11 126.766
R316 minus.n39 minus.t23 126.766
R317 minus.n52 minus.t17 126.766
R318 minus.n54 minus.t21 126.766
R319 minus.n37 minus.t5 126.766
R320 minus.n59 minus.t19 126.766
R321 minus.n35 minus.t2 126.766
R322 minus.n64 minus.t13 126.766
R323 minus.n66 minus.t8 126.766
R324 minus.n8 minus.n7 48.2005
R325 minus.n18 minus.n5 48.2005
R326 minus.n20 minus.n3 48.2005
R327 minus.n30 minus.n1 48.2005
R328 minus.n42 minus.n41 48.2005
R329 minus.n52 minus.n39 48.2005
R330 minus.n54 minus.n37 48.2005
R331 minus.n64 minus.n35 48.2005
R332 minus.n14 minus.n13 47.4702
R333 minus.n25 minus.n24 47.4702
R334 minus.n48 minus.n47 47.4702
R335 minus.n59 minus.n58 47.4702
R336 minus.n32 minus.n31 46.0096
R337 minus.n66 minus.n65 46.0096
R338 minus.n10 minus.n9 45.0871
R339 minus.n44 minus.n43 45.0871
R340 minus.n68 minus.n33 31.7013
R341 minus.n13 minus.n12 25.5611
R342 minus.n26 minus.n25 25.5611
R343 minus.n47 minus.n46 25.5611
R344 minus.n60 minus.n59 25.5611
R345 minus.n20 minus.n19 24.1005
R346 minus.n19 minus.n18 24.1005
R347 minus.n53 minus.n52 24.1005
R348 minus.n54 minus.n53 24.1005
R349 minus.n12 minus.n7 22.6399
R350 minus.n26 minus.n1 22.6399
R351 minus.n46 minus.n41 22.6399
R352 minus.n60 minus.n35 22.6399
R353 minus.n9 minus.n8 14.1472
R354 minus.n43 minus.n42 14.1472
R355 minus.n68 minus.n67 6.52702
R356 minus.n31 minus.n30 2.19141
R357 minus.n65 minus.n64 2.19141
R358 minus.n14 minus.n5 0.730803
R359 minus.n24 minus.n3 0.730803
R360 minus.n48 minus.n39 0.730803
R361 minus.n58 minus.n37 0.730803
R362 minus.n33 minus.n0 0.189894
R363 minus.n29 minus.n0 0.189894
R364 minus.n29 minus.n28 0.189894
R365 minus.n28 minus.n27 0.189894
R366 minus.n27 minus.n2 0.189894
R367 minus.n23 minus.n2 0.189894
R368 minus.n23 minus.n22 0.189894
R369 minus.n22 minus.n21 0.189894
R370 minus.n21 minus.n4 0.189894
R371 minus.n17 minus.n4 0.189894
R372 minus.n17 minus.n16 0.189894
R373 minus.n16 minus.n15 0.189894
R374 minus.n15 minus.n6 0.189894
R375 minus.n11 minus.n6 0.189894
R376 minus.n11 minus.n10 0.189894
R377 minus.n45 minus.n44 0.189894
R378 minus.n45 minus.n40 0.189894
R379 minus.n49 minus.n40 0.189894
R380 minus.n50 minus.n49 0.189894
R381 minus.n51 minus.n50 0.189894
R382 minus.n51 minus.n38 0.189894
R383 minus.n55 minus.n38 0.189894
R384 minus.n56 minus.n55 0.189894
R385 minus.n57 minus.n56 0.189894
R386 minus.n57 minus.n36 0.189894
R387 minus.n61 minus.n36 0.189894
R388 minus.n62 minus.n61 0.189894
R389 minus.n63 minus.n62 0.189894
R390 minus.n63 minus.n34 0.189894
R391 minus.n67 minus.n34 0.189894
R392 minus minus.n68 0.188
R393 drain_right.n13 drain_right.n11 240.849
R394 drain_right.n7 drain_right.n5 240.847
R395 drain_right.n2 drain_right.n0 240.847
R396 drain_right.n13 drain_right.n12 240.132
R397 drain_right.n15 drain_right.n14 240.132
R398 drain_right.n17 drain_right.n16 240.132
R399 drain_right.n19 drain_right.n18 240.132
R400 drain_right.n21 drain_right.n20 240.132
R401 drain_right.n7 drain_right.n6 240.131
R402 drain_right.n9 drain_right.n8 240.131
R403 drain_right.n4 drain_right.n3 240.131
R404 drain_right.n2 drain_right.n1 240.131
R405 drain_right drain_right.n10 25.2779
R406 drain_right.n5 drain_right.t10 19.8005
R407 drain_right.n5 drain_right.t15 19.8005
R408 drain_right.n6 drain_right.t4 19.8005
R409 drain_right.n6 drain_right.t21 19.8005
R410 drain_right.n8 drain_right.t2 19.8005
R411 drain_right.n8 drain_right.t18 19.8005
R412 drain_right.n3 drain_right.t0 19.8005
R413 drain_right.n3 drain_right.t6 19.8005
R414 drain_right.n1 drain_right.t16 19.8005
R415 drain_right.n1 drain_right.t12 19.8005
R416 drain_right.n0 drain_right.t14 19.8005
R417 drain_right.n0 drain_right.t7 19.8005
R418 drain_right.n11 drain_right.t22 19.8005
R419 drain_right.n11 drain_right.t9 19.8005
R420 drain_right.n12 drain_right.t3 19.8005
R421 drain_right.n12 drain_right.t17 19.8005
R422 drain_right.n14 drain_right.t13 19.8005
R423 drain_right.n14 drain_right.t19 19.8005
R424 drain_right.n16 drain_right.t11 19.8005
R425 drain_right.n16 drain_right.t23 19.8005
R426 drain_right.n18 drain_right.t20 19.8005
R427 drain_right.n18 drain_right.t5 19.8005
R428 drain_right.n20 drain_right.t1 19.8005
R429 drain_right.n20 drain_right.t8 19.8005
R430 drain_right drain_right.n21 6.36873
R431 drain_right.n9 drain_right.n7 0.716017
R432 drain_right.n4 drain_right.n2 0.716017
R433 drain_right.n21 drain_right.n19 0.716017
R434 drain_right.n19 drain_right.n17 0.716017
R435 drain_right.n17 drain_right.n15 0.716017
R436 drain_right.n15 drain_right.n13 0.716017
R437 drain_right.n10 drain_right.n9 0.302913
R438 drain_right.n10 drain_right.n4 0.302913
C0 minus plus 4.71453f
C1 plus source 2.41973f
C2 minus drain_left 0.181087f
C3 source drain_left 6.72479f
C4 minus source 2.40586f
C5 plus drain_right 0.452367f
C6 drain_left drain_right 1.55985f
C7 minus drain_right 1.68928f
C8 source drain_right 6.72631f
C9 plus drain_left 1.97535f
C10 drain_right a_n2874_n1088# 4.88226f
C11 drain_left a_n2874_n1088# 5.25235f
C12 source a_n2874_n1088# 2.931975f
C13 minus a_n2874_n1088# 10.60857f
C14 plus a_n2874_n1088# 11.651681f
C15 drain_right.t14 a_n2874_n1088# 0.017737f
C16 drain_right.t7 a_n2874_n1088# 0.017737f
C17 drain_right.n0 a_n2874_n1088# 0.069721f
C18 drain_right.t16 a_n2874_n1088# 0.017737f
C19 drain_right.t12 a_n2874_n1088# 0.017737f
C20 drain_right.n1 a_n2874_n1088# 0.068921f
C21 drain_right.n2 a_n2874_n1088# 0.529162f
C22 drain_right.t0 a_n2874_n1088# 0.017737f
C23 drain_right.t6 a_n2874_n1088# 0.017737f
C24 drain_right.n3 a_n2874_n1088# 0.068921f
C25 drain_right.n4 a_n2874_n1088# 0.232305f
C26 drain_right.t10 a_n2874_n1088# 0.017737f
C27 drain_right.t15 a_n2874_n1088# 0.017737f
C28 drain_right.n5 a_n2874_n1088# 0.069721f
C29 drain_right.t4 a_n2874_n1088# 0.017737f
C30 drain_right.t21 a_n2874_n1088# 0.017737f
C31 drain_right.n6 a_n2874_n1088# 0.068921f
C32 drain_right.n7 a_n2874_n1088# 0.529162f
C33 drain_right.t2 a_n2874_n1088# 0.017737f
C34 drain_right.t18 a_n2874_n1088# 0.017737f
C35 drain_right.n8 a_n2874_n1088# 0.068921f
C36 drain_right.n9 a_n2874_n1088# 0.232305f
C37 drain_right.n10 a_n2874_n1088# 0.797423f
C38 drain_right.t22 a_n2874_n1088# 0.017737f
C39 drain_right.t9 a_n2874_n1088# 0.017737f
C40 drain_right.n11 a_n2874_n1088# 0.069722f
C41 drain_right.t3 a_n2874_n1088# 0.017737f
C42 drain_right.t17 a_n2874_n1088# 0.017737f
C43 drain_right.n12 a_n2874_n1088# 0.068921f
C44 drain_right.n13 a_n2874_n1088# 0.529162f
C45 drain_right.t13 a_n2874_n1088# 0.017737f
C46 drain_right.t19 a_n2874_n1088# 0.017737f
C47 drain_right.n14 a_n2874_n1088# 0.068921f
C48 drain_right.n15 a_n2874_n1088# 0.260461f
C49 drain_right.t11 a_n2874_n1088# 0.017737f
C50 drain_right.t23 a_n2874_n1088# 0.017737f
C51 drain_right.n16 a_n2874_n1088# 0.068921f
C52 drain_right.n17 a_n2874_n1088# 0.260461f
C53 drain_right.t20 a_n2874_n1088# 0.017737f
C54 drain_right.t5 a_n2874_n1088# 0.017737f
C55 drain_right.n18 a_n2874_n1088# 0.068921f
C56 drain_right.n19 a_n2874_n1088# 0.260461f
C57 drain_right.t1 a_n2874_n1088# 0.017737f
C58 drain_right.t8 a_n2874_n1088# 0.017737f
C59 drain_right.n20 a_n2874_n1088# 0.068921f
C60 drain_right.n21 a_n2874_n1088# 0.453299f
C61 minus.n0 a_n2874_n1088# 0.036503f
C62 minus.t3 a_n2874_n1088# 0.061891f
C63 minus.n1 a_n2874_n1088# 0.067865f
C64 minus.t15 a_n2874_n1088# 0.061891f
C65 minus.n2 a_n2874_n1088# 0.036503f
C66 minus.t12 a_n2874_n1088# 0.061891f
C67 minus.n3 a_n2874_n1088# 0.06449f
C68 minus.n4 a_n2874_n1088# 0.036503f
C69 minus.t4 a_n2874_n1088# 0.061891f
C70 minus.n5 a_n2874_n1088# 0.06449f
C71 minus.t10 a_n2874_n1088# 0.061891f
C72 minus.n6 a_n2874_n1088# 0.036503f
C73 minus.t6 a_n2874_n1088# 0.061891f
C74 minus.n7 a_n2874_n1088# 0.067865f
C75 minus.t14 a_n2874_n1088# 0.072963f
C76 minus.t1 a_n2874_n1088# 0.061891f
C77 minus.n8 a_n2874_n1088# 0.072185f
C78 minus.n9 a_n2874_n1088# 0.0545f
C79 minus.n10 a_n2874_n1088# 0.148217f
C80 minus.n11 a_n2874_n1088# 0.036503f
C81 minus.n12 a_n2874_n1088# 0.008283f
C82 minus.t20 a_n2874_n1088# 0.061891f
C83 minus.n13 a_n2874_n1088# 0.068203f
C84 minus.n14 a_n2874_n1088# 0.008283f
C85 minus.n15 a_n2874_n1088# 0.036503f
C86 minus.n16 a_n2874_n1088# 0.036503f
C87 minus.n17 a_n2874_n1088# 0.036503f
C88 minus.n18 a_n2874_n1088# 0.06809f
C89 minus.n19 a_n2874_n1088# 0.008283f
C90 minus.t0 a_n2874_n1088# 0.061891f
C91 minus.n20 a_n2874_n1088# 0.06809f
C92 minus.n21 a_n2874_n1088# 0.036503f
C93 minus.n22 a_n2874_n1088# 0.036503f
C94 minus.n23 a_n2874_n1088# 0.036503f
C95 minus.n24 a_n2874_n1088# 0.008283f
C96 minus.t18 a_n2874_n1088# 0.061891f
C97 minus.n25 a_n2874_n1088# 0.068203f
C98 minus.n26 a_n2874_n1088# 0.008283f
C99 minus.n27 a_n2874_n1088# 0.036503f
C100 minus.n28 a_n2874_n1088# 0.036503f
C101 minus.n29 a_n2874_n1088# 0.036503f
C102 minus.n30 a_n2874_n1088# 0.064715f
C103 minus.n31 a_n2874_n1088# 0.008283f
C104 minus.t22 a_n2874_n1088# 0.061891f
C105 minus.n32 a_n2874_n1088# 0.064039f
C106 minus.n33 a_n2874_n1088# 1.04291f
C107 minus.n34 a_n2874_n1088# 0.036503f
C108 minus.t2 a_n2874_n1088# 0.061891f
C109 minus.n35 a_n2874_n1088# 0.067865f
C110 minus.n36 a_n2874_n1088# 0.036503f
C111 minus.t5 a_n2874_n1088# 0.061891f
C112 minus.n37 a_n2874_n1088# 0.06449f
C113 minus.n38 a_n2874_n1088# 0.036503f
C114 minus.t23 a_n2874_n1088# 0.061891f
C115 minus.n39 a_n2874_n1088# 0.06449f
C116 minus.n40 a_n2874_n1088# 0.036503f
C117 minus.t7 a_n2874_n1088# 0.061891f
C118 minus.n41 a_n2874_n1088# 0.067865f
C119 minus.t9 a_n2874_n1088# 0.072963f
C120 minus.t16 a_n2874_n1088# 0.061891f
C121 minus.n42 a_n2874_n1088# 0.072185f
C122 minus.n43 a_n2874_n1088# 0.0545f
C123 minus.n44 a_n2874_n1088# 0.148217f
C124 minus.n45 a_n2874_n1088# 0.036503f
C125 minus.n46 a_n2874_n1088# 0.008283f
C126 minus.t11 a_n2874_n1088# 0.061891f
C127 minus.n47 a_n2874_n1088# 0.068203f
C128 minus.n48 a_n2874_n1088# 0.008283f
C129 minus.n49 a_n2874_n1088# 0.036503f
C130 minus.n50 a_n2874_n1088# 0.036503f
C131 minus.n51 a_n2874_n1088# 0.036503f
C132 minus.t17 a_n2874_n1088# 0.061891f
C133 minus.n52 a_n2874_n1088# 0.06809f
C134 minus.n53 a_n2874_n1088# 0.008283f
C135 minus.t21 a_n2874_n1088# 0.061891f
C136 minus.n54 a_n2874_n1088# 0.06809f
C137 minus.n55 a_n2874_n1088# 0.036503f
C138 minus.n56 a_n2874_n1088# 0.036503f
C139 minus.n57 a_n2874_n1088# 0.036503f
C140 minus.n58 a_n2874_n1088# 0.008283f
C141 minus.t19 a_n2874_n1088# 0.061891f
C142 minus.n59 a_n2874_n1088# 0.068203f
C143 minus.n60 a_n2874_n1088# 0.008283f
C144 minus.n61 a_n2874_n1088# 0.036503f
C145 minus.n62 a_n2874_n1088# 0.036503f
C146 minus.n63 a_n2874_n1088# 0.036503f
C147 minus.t13 a_n2874_n1088# 0.061891f
C148 minus.n64 a_n2874_n1088# 0.064715f
C149 minus.n65 a_n2874_n1088# 0.008283f
C150 minus.t8 a_n2874_n1088# 0.061891f
C151 minus.n66 a_n2874_n1088# 0.064039f
C152 minus.n67 a_n2874_n1088# 0.240968f
C153 minus.n68 a_n2874_n1088# 1.28124f
C154 drain_left.t22 a_n2874_n1088# 0.017508f
C155 drain_left.t11 a_n2874_n1088# 0.017508f
C156 drain_left.n0 a_n2874_n1088# 0.06882f
C157 drain_left.t19 a_n2874_n1088# 0.017508f
C158 drain_left.t1 a_n2874_n1088# 0.017508f
C159 drain_left.n1 a_n2874_n1088# 0.068029f
C160 drain_left.n2 a_n2874_n1088# 0.522317f
C161 drain_left.t16 a_n2874_n1088# 0.017508f
C162 drain_left.t4 a_n2874_n1088# 0.017508f
C163 drain_left.n3 a_n2874_n1088# 0.068029f
C164 drain_left.n4 a_n2874_n1088# 0.2293f
C165 drain_left.t8 a_n2874_n1088# 0.017508f
C166 drain_left.t12 a_n2874_n1088# 0.017508f
C167 drain_left.n5 a_n2874_n1088# 0.06882f
C168 drain_left.t6 a_n2874_n1088# 0.017508f
C169 drain_left.t14 a_n2874_n1088# 0.017508f
C170 drain_left.n6 a_n2874_n1088# 0.068029f
C171 drain_left.n7 a_n2874_n1088# 0.522318f
C172 drain_left.t7 a_n2874_n1088# 0.017508f
C173 drain_left.t23 a_n2874_n1088# 0.017508f
C174 drain_left.n8 a_n2874_n1088# 0.068029f
C175 drain_left.n9 a_n2874_n1088# 0.2293f
C176 drain_left.n10 a_n2874_n1088# 0.829623f
C177 drain_left.t17 a_n2874_n1088# 0.017508f
C178 drain_left.t9 a_n2874_n1088# 0.017508f
C179 drain_left.n11 a_n2874_n1088# 0.06882f
C180 drain_left.t2 a_n2874_n1088# 0.017508f
C181 drain_left.t15 a_n2874_n1088# 0.017508f
C182 drain_left.n12 a_n2874_n1088# 0.068029f
C183 drain_left.n13 a_n2874_n1088# 0.522317f
C184 drain_left.t5 a_n2874_n1088# 0.017508f
C185 drain_left.t0 a_n2874_n1088# 0.017508f
C186 drain_left.n14 a_n2874_n1088# 0.068029f
C187 drain_left.n15 a_n2874_n1088# 0.257092f
C188 drain_left.t13 a_n2874_n1088# 0.017508f
C189 drain_left.t3 a_n2874_n1088# 0.017508f
C190 drain_left.n16 a_n2874_n1088# 0.068029f
C191 drain_left.n17 a_n2874_n1088# 0.257092f
C192 drain_left.t18 a_n2874_n1088# 0.017508f
C193 drain_left.t10 a_n2874_n1088# 0.017508f
C194 drain_left.n18 a_n2874_n1088# 0.068029f
C195 drain_left.n19 a_n2874_n1088# 0.257092f
C196 drain_left.t20 a_n2874_n1088# 0.017508f
C197 drain_left.t21 a_n2874_n1088# 0.017508f
C198 drain_left.n20 a_n2874_n1088# 0.068029f
C199 drain_left.n21 a_n2874_n1088# 0.447435f
C200 source.t45 a_n2874_n1088# 0.163812f
C201 source.n0 a_n2874_n1088# 0.740397f
C202 source.t43 a_n2874_n1088# 0.029432f
C203 source.t40 a_n2874_n1088# 0.029432f
C204 source.n1 a_n2874_n1088# 0.095451f
C205 source.n2 a_n2874_n1088# 0.40048f
C206 source.t46 a_n2874_n1088# 0.029432f
C207 source.t27 a_n2874_n1088# 0.029432f
C208 source.n3 a_n2874_n1088# 0.095451f
C209 source.n4 a_n2874_n1088# 0.40048f
C210 source.t41 a_n2874_n1088# 0.029432f
C211 source.t31 a_n2874_n1088# 0.029432f
C212 source.n5 a_n2874_n1088# 0.095451f
C213 source.n6 a_n2874_n1088# 0.40048f
C214 source.t28 a_n2874_n1088# 0.029432f
C215 source.t24 a_n2874_n1088# 0.029432f
C216 source.n7 a_n2874_n1088# 0.095451f
C217 source.n8 a_n2874_n1088# 0.40048f
C218 source.t42 a_n2874_n1088# 0.029432f
C219 source.t37 a_n2874_n1088# 0.029432f
C220 source.n9 a_n2874_n1088# 0.095451f
C221 source.n10 a_n2874_n1088# 0.40048f
C222 source.t33 a_n2874_n1088# 0.163812f
C223 source.n11 a_n2874_n1088# 0.382902f
C224 source.t1 a_n2874_n1088# 0.163812f
C225 source.n12 a_n2874_n1088# 0.382902f
C226 source.t17 a_n2874_n1088# 0.029432f
C227 source.t19 a_n2874_n1088# 0.029432f
C228 source.n13 a_n2874_n1088# 0.095451f
C229 source.n14 a_n2874_n1088# 0.40048f
C230 source.t18 a_n2874_n1088# 0.029432f
C231 source.t20 a_n2874_n1088# 0.029432f
C232 source.n15 a_n2874_n1088# 0.095451f
C233 source.n16 a_n2874_n1088# 0.40048f
C234 source.t13 a_n2874_n1088# 0.029432f
C235 source.t8 a_n2874_n1088# 0.029432f
C236 source.n17 a_n2874_n1088# 0.095451f
C237 source.n18 a_n2874_n1088# 0.40048f
C238 source.t15 a_n2874_n1088# 0.029432f
C239 source.t16 a_n2874_n1088# 0.029432f
C240 source.n19 a_n2874_n1088# 0.095451f
C241 source.n20 a_n2874_n1088# 0.40048f
C242 source.t4 a_n2874_n1088# 0.029432f
C243 source.t23 a_n2874_n1088# 0.029432f
C244 source.n21 a_n2874_n1088# 0.095451f
C245 source.n22 a_n2874_n1088# 0.40048f
C246 source.t10 a_n2874_n1088# 0.163812f
C247 source.n23 a_n2874_n1088# 1.0432f
C248 source.t34 a_n2874_n1088# 0.163812f
C249 source.n24 a_n2874_n1088# 1.0432f
C250 source.t32 a_n2874_n1088# 0.029432f
C251 source.t35 a_n2874_n1088# 0.029432f
C252 source.n25 a_n2874_n1088# 0.095451f
C253 source.n26 a_n2874_n1088# 0.40048f
C254 source.t39 a_n2874_n1088# 0.029432f
C255 source.t25 a_n2874_n1088# 0.029432f
C256 source.n27 a_n2874_n1088# 0.095451f
C257 source.n28 a_n2874_n1088# 0.40048f
C258 source.t36 a_n2874_n1088# 0.029432f
C259 source.t47 a_n2874_n1088# 0.029432f
C260 source.n29 a_n2874_n1088# 0.095451f
C261 source.n30 a_n2874_n1088# 0.40048f
C262 source.t38 a_n2874_n1088# 0.029432f
C263 source.t29 a_n2874_n1088# 0.029432f
C264 source.n31 a_n2874_n1088# 0.095451f
C265 source.n32 a_n2874_n1088# 0.40048f
C266 source.t30 a_n2874_n1088# 0.029432f
C267 source.t44 a_n2874_n1088# 0.029432f
C268 source.n33 a_n2874_n1088# 0.095451f
C269 source.n34 a_n2874_n1088# 0.40048f
C270 source.t26 a_n2874_n1088# 0.163812f
C271 source.n35 a_n2874_n1088# 0.382902f
C272 source.t21 a_n2874_n1088# 0.163812f
C273 source.n36 a_n2874_n1088# 0.382902f
C274 source.t7 a_n2874_n1088# 0.029432f
C275 source.t22 a_n2874_n1088# 0.029432f
C276 source.n37 a_n2874_n1088# 0.095451f
C277 source.n38 a_n2874_n1088# 0.40048f
C278 source.t12 a_n2874_n1088# 0.029432f
C279 source.t14 a_n2874_n1088# 0.029432f
C280 source.n39 a_n2874_n1088# 0.095451f
C281 source.n40 a_n2874_n1088# 0.40048f
C282 source.t11 a_n2874_n1088# 0.029432f
C283 source.t3 a_n2874_n1088# 0.029432f
C284 source.n41 a_n2874_n1088# 0.095451f
C285 source.n42 a_n2874_n1088# 0.40048f
C286 source.t9 a_n2874_n1088# 0.029432f
C287 source.t0 a_n2874_n1088# 0.029432f
C288 source.n43 a_n2874_n1088# 0.095451f
C289 source.n44 a_n2874_n1088# 0.40048f
C290 source.t2 a_n2874_n1088# 0.029432f
C291 source.t5 a_n2874_n1088# 0.029432f
C292 source.n45 a_n2874_n1088# 0.095451f
C293 source.n46 a_n2874_n1088# 0.40048f
C294 source.t6 a_n2874_n1088# 0.163812f
C295 source.n47 a_n2874_n1088# 0.609589f
C296 source.n48 a_n2874_n1088# 0.762914f
C297 plus.n0 a_n2874_n1088# 0.036887f
C298 plus.t2 a_n2874_n1088# 0.062541f
C299 plus.t3 a_n2874_n1088# 0.062541f
C300 plus.n1 a_n2874_n1088# 0.036887f
C301 plus.t13 a_n2874_n1088# 0.062541f
C302 plus.n2 a_n2874_n1088# 0.036887f
C303 plus.t5 a_n2874_n1088# 0.062541f
C304 plus.n3 a_n2874_n1088# 0.06892f
C305 plus.n4 a_n2874_n1088# 0.036887f
C306 plus.t20 a_n2874_n1088# 0.062541f
C307 plus.t10 a_n2874_n1088# 0.062541f
C308 plus.n5 a_n2874_n1088# 0.036887f
C309 plus.t23 a_n2874_n1088# 0.062541f
C310 plus.n6 a_n2874_n1088# 0.068806f
C311 plus.n7 a_n2874_n1088# 0.036887f
C312 plus.t18 a_n2874_n1088# 0.062541f
C313 plus.t8 a_n2874_n1088# 0.062541f
C314 plus.n8 a_n2874_n1088# 0.036887f
C315 plus.t21 a_n2874_n1088# 0.062541f
C316 plus.n9 a_n2874_n1088# 0.068578f
C317 plus.t14 a_n2874_n1088# 0.062541f
C318 plus.n10 a_n2874_n1088# 0.072943f
C319 plus.t6 a_n2874_n1088# 0.07373f
C320 plus.n11 a_n2874_n1088# 0.055073f
C321 plus.n12 a_n2874_n1088# 0.149775f
C322 plus.n13 a_n2874_n1088# 0.036887f
C323 plus.n14 a_n2874_n1088# 0.00837f
C324 plus.n15 a_n2874_n1088# 0.06892f
C325 plus.n16 a_n2874_n1088# 0.00837f
C326 plus.n17 a_n2874_n1088# 0.065167f
C327 plus.n18 a_n2874_n1088# 0.036887f
C328 plus.n19 a_n2874_n1088# 0.036887f
C329 plus.n20 a_n2874_n1088# 0.036887f
C330 plus.n21 a_n2874_n1088# 0.00837f
C331 plus.n22 a_n2874_n1088# 0.068806f
C332 plus.n23 a_n2874_n1088# 0.065167f
C333 plus.n24 a_n2874_n1088# 0.00837f
C334 plus.n25 a_n2874_n1088# 0.036887f
C335 plus.n26 a_n2874_n1088# 0.036887f
C336 plus.n27 a_n2874_n1088# 0.036887f
C337 plus.n28 a_n2874_n1088# 0.00837f
C338 plus.n29 a_n2874_n1088# 0.068578f
C339 plus.n30 a_n2874_n1088# 0.065395f
C340 plus.n31 a_n2874_n1088# 0.00837f
C341 plus.n32 a_n2874_n1088# 0.064712f
C342 plus.n33 a_n2874_n1088# 0.255365f
C343 plus.n34 a_n2874_n1088# 0.036887f
C344 plus.t1 a_n2874_n1088# 0.062541f
C345 plus.n35 a_n2874_n1088# 0.036887f
C346 plus.t12 a_n2874_n1088# 0.062541f
C347 plus.n36 a_n2874_n1088# 0.036887f
C348 plus.t4 a_n2874_n1088# 0.062541f
C349 plus.t22 a_n2874_n1088# 0.062541f
C350 plus.n37 a_n2874_n1088# 0.06892f
C351 plus.n38 a_n2874_n1088# 0.036887f
C352 plus.t7 a_n2874_n1088# 0.062541f
C353 plus.n39 a_n2874_n1088# 0.036887f
C354 plus.t19 a_n2874_n1088# 0.062541f
C355 plus.t16 a_n2874_n1088# 0.062541f
C356 plus.n40 a_n2874_n1088# 0.068806f
C357 plus.n41 a_n2874_n1088# 0.036887f
C358 plus.t0 a_n2874_n1088# 0.062541f
C359 plus.n42 a_n2874_n1088# 0.036887f
C360 plus.t17 a_n2874_n1088# 0.062541f
C361 plus.t9 a_n2874_n1088# 0.062541f
C362 plus.n43 a_n2874_n1088# 0.068578f
C363 plus.t11 a_n2874_n1088# 0.07373f
C364 plus.t15 a_n2874_n1088# 0.062541f
C365 plus.n44 a_n2874_n1088# 0.072943f
C366 plus.n45 a_n2874_n1088# 0.055073f
C367 plus.n46 a_n2874_n1088# 0.149775f
C368 plus.n47 a_n2874_n1088# 0.036887f
C369 plus.n48 a_n2874_n1088# 0.00837f
C370 plus.n49 a_n2874_n1088# 0.06892f
C371 plus.n50 a_n2874_n1088# 0.00837f
C372 plus.n51 a_n2874_n1088# 0.065167f
C373 plus.n52 a_n2874_n1088# 0.036887f
C374 plus.n53 a_n2874_n1088# 0.036887f
C375 plus.n54 a_n2874_n1088# 0.036887f
C376 plus.n55 a_n2874_n1088# 0.00837f
C377 plus.n56 a_n2874_n1088# 0.068806f
C378 plus.n57 a_n2874_n1088# 0.065167f
C379 plus.n58 a_n2874_n1088# 0.00837f
C380 plus.n59 a_n2874_n1088# 0.036887f
C381 plus.n60 a_n2874_n1088# 0.036887f
C382 plus.n61 a_n2874_n1088# 0.036887f
C383 plus.n62 a_n2874_n1088# 0.00837f
C384 plus.n63 a_n2874_n1088# 0.068578f
C385 plus.n64 a_n2874_n1088# 0.065395f
C386 plus.n65 a_n2874_n1088# 0.00837f
C387 plus.n66 a_n2874_n1088# 0.064712f
C388 plus.n67 a_n2874_n1088# 1.01505f
.ends

