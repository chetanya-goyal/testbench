* NGSPICE file created from diffpair270.ext - technology: sky130A

.subckt diffpair270 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=0.3
X1 drain_right.t0 minus.t1 source.t3 a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=0.3
X2 a_n968_n2092# a_n968_n2092# a_n968_n2092# a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X3 a_n968_n2092# a_n968_n2092# a_n968_n2092# a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X4 drain_left.t1 plus.t0 source.t1 a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=0.3
X5 a_n968_n2092# a_n968_n2092# a_n968_n2092# a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X6 a_n968_n2092# a_n968_n2092# a_n968_n2092# a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X7 drain_left.t0 plus.t1 source.t0 a_n968_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=0.3
R0 minus.n0 minus.t0 799.98
R1 minus.n0 minus.t1 778.222
R2 minus minus.n0 0.188
R3 source.n122 source.n96 289.615
R4 source.n90 source.n64 289.615
R5 source.n26 source.n0 289.615
R6 source.n58 source.n32 289.615
R7 source.n107 source.n106 185
R8 source.n104 source.n103 185
R9 source.n113 source.n112 185
R10 source.n115 source.n114 185
R11 source.n100 source.n99 185
R12 source.n121 source.n120 185
R13 source.n123 source.n122 185
R14 source.n75 source.n74 185
R15 source.n72 source.n71 185
R16 source.n81 source.n80 185
R17 source.n83 source.n82 185
R18 source.n68 source.n67 185
R19 source.n89 source.n88 185
R20 source.n91 source.n90 185
R21 source.n27 source.n26 185
R22 source.n25 source.n24 185
R23 source.n4 source.n3 185
R24 source.n19 source.n18 185
R25 source.n17 source.n16 185
R26 source.n8 source.n7 185
R27 source.n11 source.n10 185
R28 source.n59 source.n58 185
R29 source.n57 source.n56 185
R30 source.n36 source.n35 185
R31 source.n51 source.n50 185
R32 source.n49 source.n48 185
R33 source.n40 source.n39 185
R34 source.n43 source.n42 185
R35 source.t3 source.n105 147.661
R36 source.t0 source.n73 147.661
R37 source.t1 source.n9 147.661
R38 source.t2 source.n41 147.661
R39 source.n106 source.n103 104.615
R40 source.n113 source.n103 104.615
R41 source.n114 source.n113 104.615
R42 source.n114 source.n99 104.615
R43 source.n121 source.n99 104.615
R44 source.n122 source.n121 104.615
R45 source.n74 source.n71 104.615
R46 source.n81 source.n71 104.615
R47 source.n82 source.n81 104.615
R48 source.n82 source.n67 104.615
R49 source.n89 source.n67 104.615
R50 source.n90 source.n89 104.615
R51 source.n26 source.n25 104.615
R52 source.n25 source.n3 104.615
R53 source.n18 source.n3 104.615
R54 source.n18 source.n17 104.615
R55 source.n17 source.n7 104.615
R56 source.n10 source.n7 104.615
R57 source.n58 source.n57 104.615
R58 source.n57 source.n35 104.615
R59 source.n50 source.n35 104.615
R60 source.n50 source.n49 104.615
R61 source.n49 source.n39 104.615
R62 source.n42 source.n39 104.615
R63 source.n106 source.t3 52.3082
R64 source.n74 source.t0 52.3082
R65 source.n10 source.t1 52.3082
R66 source.n42 source.t2 52.3082
R67 source.n127 source.n126 32.1853
R68 source.n95 source.n94 32.1853
R69 source.n31 source.n30 32.1853
R70 source.n63 source.n62 32.1853
R71 source.n95 source.n63 17.8436
R72 source.n107 source.n105 15.6674
R73 source.n75 source.n73 15.6674
R74 source.n11 source.n9 15.6674
R75 source.n43 source.n41 15.6674
R76 source.n108 source.n104 12.8005
R77 source.n76 source.n72 12.8005
R78 source.n12 source.n8 12.8005
R79 source.n44 source.n40 12.8005
R80 source.n112 source.n111 12.0247
R81 source.n80 source.n79 12.0247
R82 source.n16 source.n15 12.0247
R83 source.n48 source.n47 12.0247
R84 source.n128 source.n31 11.766
R85 source.n115 source.n102 11.249
R86 source.n83 source.n70 11.249
R87 source.n19 source.n6 11.249
R88 source.n51 source.n38 11.249
R89 source.n116 source.n100 10.4732
R90 source.n84 source.n68 10.4732
R91 source.n20 source.n4 10.4732
R92 source.n52 source.n36 10.4732
R93 source.n120 source.n119 9.69747
R94 source.n88 source.n87 9.69747
R95 source.n24 source.n23 9.69747
R96 source.n56 source.n55 9.69747
R97 source.n126 source.n125 9.45567
R98 source.n94 source.n93 9.45567
R99 source.n30 source.n29 9.45567
R100 source.n62 source.n61 9.45567
R101 source.n125 source.n124 9.3005
R102 source.n98 source.n97 9.3005
R103 source.n119 source.n118 9.3005
R104 source.n117 source.n116 9.3005
R105 source.n102 source.n101 9.3005
R106 source.n111 source.n110 9.3005
R107 source.n109 source.n108 9.3005
R108 source.n93 source.n92 9.3005
R109 source.n66 source.n65 9.3005
R110 source.n87 source.n86 9.3005
R111 source.n85 source.n84 9.3005
R112 source.n70 source.n69 9.3005
R113 source.n79 source.n78 9.3005
R114 source.n77 source.n76 9.3005
R115 source.n29 source.n28 9.3005
R116 source.n2 source.n1 9.3005
R117 source.n23 source.n22 9.3005
R118 source.n21 source.n20 9.3005
R119 source.n6 source.n5 9.3005
R120 source.n15 source.n14 9.3005
R121 source.n13 source.n12 9.3005
R122 source.n61 source.n60 9.3005
R123 source.n34 source.n33 9.3005
R124 source.n55 source.n54 9.3005
R125 source.n53 source.n52 9.3005
R126 source.n38 source.n37 9.3005
R127 source.n47 source.n46 9.3005
R128 source.n45 source.n44 9.3005
R129 source.n123 source.n98 8.92171
R130 source.n91 source.n66 8.92171
R131 source.n27 source.n2 8.92171
R132 source.n59 source.n34 8.92171
R133 source.n124 source.n96 8.14595
R134 source.n92 source.n64 8.14595
R135 source.n28 source.n0 8.14595
R136 source.n60 source.n32 8.14595
R137 source.n126 source.n96 5.81868
R138 source.n94 source.n64 5.81868
R139 source.n30 source.n0 5.81868
R140 source.n62 source.n32 5.81868
R141 source.n128 source.n127 5.53498
R142 source.n124 source.n123 5.04292
R143 source.n92 source.n91 5.04292
R144 source.n28 source.n27 5.04292
R145 source.n60 source.n59 5.04292
R146 source.n109 source.n105 4.38594
R147 source.n77 source.n73 4.38594
R148 source.n13 source.n9 4.38594
R149 source.n45 source.n41 4.38594
R150 source.n120 source.n98 4.26717
R151 source.n88 source.n66 4.26717
R152 source.n24 source.n2 4.26717
R153 source.n56 source.n34 4.26717
R154 source.n119 source.n100 3.49141
R155 source.n87 source.n68 3.49141
R156 source.n23 source.n4 3.49141
R157 source.n55 source.n36 3.49141
R158 source.n116 source.n115 2.71565
R159 source.n84 source.n83 2.71565
R160 source.n20 source.n19 2.71565
R161 source.n52 source.n51 2.71565
R162 source.n112 source.n102 1.93989
R163 source.n80 source.n70 1.93989
R164 source.n16 source.n6 1.93989
R165 source.n48 source.n38 1.93989
R166 source.n111 source.n104 1.16414
R167 source.n79 source.n72 1.16414
R168 source.n15 source.n8 1.16414
R169 source.n47 source.n40 1.16414
R170 source.n63 source.n31 0.741879
R171 source.n127 source.n95 0.741879
R172 source.n108 source.n107 0.388379
R173 source.n76 source.n75 0.388379
R174 source.n12 source.n11 0.388379
R175 source.n44 source.n43 0.388379
R176 source source.n128 0.188
R177 source.n110 source.n109 0.155672
R178 source.n110 source.n101 0.155672
R179 source.n117 source.n101 0.155672
R180 source.n118 source.n117 0.155672
R181 source.n118 source.n97 0.155672
R182 source.n125 source.n97 0.155672
R183 source.n78 source.n77 0.155672
R184 source.n78 source.n69 0.155672
R185 source.n85 source.n69 0.155672
R186 source.n86 source.n85 0.155672
R187 source.n86 source.n65 0.155672
R188 source.n93 source.n65 0.155672
R189 source.n29 source.n1 0.155672
R190 source.n22 source.n1 0.155672
R191 source.n22 source.n21 0.155672
R192 source.n21 source.n5 0.155672
R193 source.n14 source.n5 0.155672
R194 source.n14 source.n13 0.155672
R195 source.n61 source.n33 0.155672
R196 source.n54 source.n33 0.155672
R197 source.n54 source.n53 0.155672
R198 source.n53 source.n37 0.155672
R199 source.n46 source.n37 0.155672
R200 source.n46 source.n45 0.155672
R201 drain_right.n26 drain_right.n0 289.615
R202 drain_right.n57 drain_right.n31 289.615
R203 drain_right.n11 drain_right.n10 185
R204 drain_right.n8 drain_right.n7 185
R205 drain_right.n17 drain_right.n16 185
R206 drain_right.n19 drain_right.n18 185
R207 drain_right.n4 drain_right.n3 185
R208 drain_right.n25 drain_right.n24 185
R209 drain_right.n27 drain_right.n26 185
R210 drain_right.n58 drain_right.n57 185
R211 drain_right.n56 drain_right.n55 185
R212 drain_right.n35 drain_right.n34 185
R213 drain_right.n50 drain_right.n49 185
R214 drain_right.n48 drain_right.n47 185
R215 drain_right.n39 drain_right.n38 185
R216 drain_right.n42 drain_right.n41 185
R217 drain_right.t0 drain_right.n9 147.661
R218 drain_right.t1 drain_right.n40 147.661
R219 drain_right.n10 drain_right.n7 104.615
R220 drain_right.n17 drain_right.n7 104.615
R221 drain_right.n18 drain_right.n17 104.615
R222 drain_right.n18 drain_right.n3 104.615
R223 drain_right.n25 drain_right.n3 104.615
R224 drain_right.n26 drain_right.n25 104.615
R225 drain_right.n57 drain_right.n56 104.615
R226 drain_right.n56 drain_right.n34 104.615
R227 drain_right.n49 drain_right.n34 104.615
R228 drain_right.n49 drain_right.n48 104.615
R229 drain_right.n48 drain_right.n38 104.615
R230 drain_right.n41 drain_right.n38 104.615
R231 drain_right drain_right.n30 71.9065
R232 drain_right drain_right.n61 54.7884
R233 drain_right.n10 drain_right.t0 52.3082
R234 drain_right.n41 drain_right.t1 52.3082
R235 drain_right.n11 drain_right.n9 15.6674
R236 drain_right.n42 drain_right.n40 15.6674
R237 drain_right.n12 drain_right.n8 12.8005
R238 drain_right.n43 drain_right.n39 12.8005
R239 drain_right.n16 drain_right.n15 12.0247
R240 drain_right.n47 drain_right.n46 12.0247
R241 drain_right.n19 drain_right.n6 11.249
R242 drain_right.n50 drain_right.n37 11.249
R243 drain_right.n20 drain_right.n4 10.4732
R244 drain_right.n51 drain_right.n35 10.4732
R245 drain_right.n24 drain_right.n23 9.69747
R246 drain_right.n55 drain_right.n54 9.69747
R247 drain_right.n30 drain_right.n29 9.45567
R248 drain_right.n61 drain_right.n60 9.45567
R249 drain_right.n29 drain_right.n28 9.3005
R250 drain_right.n2 drain_right.n1 9.3005
R251 drain_right.n23 drain_right.n22 9.3005
R252 drain_right.n21 drain_right.n20 9.3005
R253 drain_right.n6 drain_right.n5 9.3005
R254 drain_right.n15 drain_right.n14 9.3005
R255 drain_right.n13 drain_right.n12 9.3005
R256 drain_right.n60 drain_right.n59 9.3005
R257 drain_right.n33 drain_right.n32 9.3005
R258 drain_right.n54 drain_right.n53 9.3005
R259 drain_right.n52 drain_right.n51 9.3005
R260 drain_right.n37 drain_right.n36 9.3005
R261 drain_right.n46 drain_right.n45 9.3005
R262 drain_right.n44 drain_right.n43 9.3005
R263 drain_right.n27 drain_right.n2 8.92171
R264 drain_right.n58 drain_right.n33 8.92171
R265 drain_right.n28 drain_right.n0 8.14595
R266 drain_right.n59 drain_right.n31 8.14595
R267 drain_right.n30 drain_right.n0 5.81868
R268 drain_right.n61 drain_right.n31 5.81868
R269 drain_right.n28 drain_right.n27 5.04292
R270 drain_right.n59 drain_right.n58 5.04292
R271 drain_right.n13 drain_right.n9 4.38594
R272 drain_right.n44 drain_right.n40 4.38594
R273 drain_right.n24 drain_right.n2 4.26717
R274 drain_right.n55 drain_right.n33 4.26717
R275 drain_right.n23 drain_right.n4 3.49141
R276 drain_right.n54 drain_right.n35 3.49141
R277 drain_right.n20 drain_right.n19 2.71565
R278 drain_right.n51 drain_right.n50 2.71565
R279 drain_right.n16 drain_right.n6 1.93989
R280 drain_right.n47 drain_right.n37 1.93989
R281 drain_right.n15 drain_right.n8 1.16414
R282 drain_right.n46 drain_right.n39 1.16414
R283 drain_right.n12 drain_right.n11 0.388379
R284 drain_right.n43 drain_right.n42 0.388379
R285 drain_right.n14 drain_right.n13 0.155672
R286 drain_right.n14 drain_right.n5 0.155672
R287 drain_right.n21 drain_right.n5 0.155672
R288 drain_right.n22 drain_right.n21 0.155672
R289 drain_right.n22 drain_right.n1 0.155672
R290 drain_right.n29 drain_right.n1 0.155672
R291 drain_right.n60 drain_right.n32 0.155672
R292 drain_right.n53 drain_right.n32 0.155672
R293 drain_right.n53 drain_right.n52 0.155672
R294 drain_right.n52 drain_right.n36 0.155672
R295 drain_right.n45 drain_right.n36 0.155672
R296 drain_right.n45 drain_right.n44 0.155672
R297 plus plus.t1 796.134
R298 plus plus.t0 781.593
R299 drain_left.n26 drain_left.n0 289.615
R300 drain_left.n57 drain_left.n31 289.615
R301 drain_left.n11 drain_left.n10 185
R302 drain_left.n8 drain_left.n7 185
R303 drain_left.n17 drain_left.n16 185
R304 drain_left.n19 drain_left.n18 185
R305 drain_left.n4 drain_left.n3 185
R306 drain_left.n25 drain_left.n24 185
R307 drain_left.n27 drain_left.n26 185
R308 drain_left.n58 drain_left.n57 185
R309 drain_left.n56 drain_left.n55 185
R310 drain_left.n35 drain_left.n34 185
R311 drain_left.n50 drain_left.n49 185
R312 drain_left.n48 drain_left.n47 185
R313 drain_left.n39 drain_left.n38 185
R314 drain_left.n42 drain_left.n41 185
R315 drain_left.t0 drain_left.n9 147.661
R316 drain_left.t1 drain_left.n40 147.661
R317 drain_left.n10 drain_left.n7 104.615
R318 drain_left.n17 drain_left.n7 104.615
R319 drain_left.n18 drain_left.n17 104.615
R320 drain_left.n18 drain_left.n3 104.615
R321 drain_left.n25 drain_left.n3 104.615
R322 drain_left.n26 drain_left.n25 104.615
R323 drain_left.n57 drain_left.n56 104.615
R324 drain_left.n56 drain_left.n34 104.615
R325 drain_left.n49 drain_left.n34 104.615
R326 drain_left.n49 drain_left.n48 104.615
R327 drain_left.n48 drain_left.n38 104.615
R328 drain_left.n41 drain_left.n38 104.615
R329 drain_left drain_left.n30 72.4597
R330 drain_left drain_left.n61 55.06
R331 drain_left.n10 drain_left.t0 52.3082
R332 drain_left.n41 drain_left.t1 52.3082
R333 drain_left.n11 drain_left.n9 15.6674
R334 drain_left.n42 drain_left.n40 15.6674
R335 drain_left.n12 drain_left.n8 12.8005
R336 drain_left.n43 drain_left.n39 12.8005
R337 drain_left.n16 drain_left.n15 12.0247
R338 drain_left.n47 drain_left.n46 12.0247
R339 drain_left.n19 drain_left.n6 11.249
R340 drain_left.n50 drain_left.n37 11.249
R341 drain_left.n20 drain_left.n4 10.4732
R342 drain_left.n51 drain_left.n35 10.4732
R343 drain_left.n24 drain_left.n23 9.69747
R344 drain_left.n55 drain_left.n54 9.69747
R345 drain_left.n30 drain_left.n29 9.45567
R346 drain_left.n61 drain_left.n60 9.45567
R347 drain_left.n29 drain_left.n28 9.3005
R348 drain_left.n2 drain_left.n1 9.3005
R349 drain_left.n23 drain_left.n22 9.3005
R350 drain_left.n21 drain_left.n20 9.3005
R351 drain_left.n6 drain_left.n5 9.3005
R352 drain_left.n15 drain_left.n14 9.3005
R353 drain_left.n13 drain_left.n12 9.3005
R354 drain_left.n60 drain_left.n59 9.3005
R355 drain_left.n33 drain_left.n32 9.3005
R356 drain_left.n54 drain_left.n53 9.3005
R357 drain_left.n52 drain_left.n51 9.3005
R358 drain_left.n37 drain_left.n36 9.3005
R359 drain_left.n46 drain_left.n45 9.3005
R360 drain_left.n44 drain_left.n43 9.3005
R361 drain_left.n27 drain_left.n2 8.92171
R362 drain_left.n58 drain_left.n33 8.92171
R363 drain_left.n28 drain_left.n0 8.14595
R364 drain_left.n59 drain_left.n31 8.14595
R365 drain_left.n30 drain_left.n0 5.81868
R366 drain_left.n61 drain_left.n31 5.81868
R367 drain_left.n28 drain_left.n27 5.04292
R368 drain_left.n59 drain_left.n58 5.04292
R369 drain_left.n13 drain_left.n9 4.38594
R370 drain_left.n44 drain_left.n40 4.38594
R371 drain_left.n24 drain_left.n2 4.26717
R372 drain_left.n55 drain_left.n33 4.26717
R373 drain_left.n23 drain_left.n4 3.49141
R374 drain_left.n54 drain_left.n35 3.49141
R375 drain_left.n20 drain_left.n19 2.71565
R376 drain_left.n51 drain_left.n50 2.71565
R377 drain_left.n16 drain_left.n6 1.93989
R378 drain_left.n47 drain_left.n37 1.93989
R379 drain_left.n15 drain_left.n8 1.16414
R380 drain_left.n46 drain_left.n39 1.16414
R381 drain_left.n12 drain_left.n11 0.388379
R382 drain_left.n43 drain_left.n42 0.388379
R383 drain_left.n14 drain_left.n13 0.155672
R384 drain_left.n14 drain_left.n5 0.155672
R385 drain_left.n21 drain_left.n5 0.155672
R386 drain_left.n22 drain_left.n21 0.155672
R387 drain_left.n22 drain_left.n1 0.155672
R388 drain_left.n29 drain_left.n1 0.155672
R389 drain_left.n60 drain_left.n32 0.155672
R390 drain_left.n53 drain_left.n32 0.155672
R391 drain_left.n53 drain_left.n52 0.155672
R392 drain_left.n52 drain_left.n36 0.155672
R393 drain_left.n45 drain_left.n36 0.155672
R394 drain_left.n45 drain_left.n44 0.155672
C0 source minus 0.581732f
C1 drain_left minus 0.171671f
C2 plus minus 3.25187f
C3 source drain_right 4.13061f
C4 drain_left drain_right 0.423956f
C5 plus drain_right 0.243327f
C6 source drain_left 4.1349f
C7 source plus 0.596076f
C8 plus drain_left 0.933311f
C9 drain_right minus 0.846828f
C10 drain_right a_n968_n2092# 4.19111f
C11 drain_left a_n968_n2092# 4.31376f
C12 source a_n968_n2092# 3.557659f
C13 minus a_n968_n2092# 3.225472f
C14 plus a_n968_n2092# 5.81133f
C15 drain_left.n0 a_n968_n2092# 0.02591f
C16 drain_left.n1 a_n968_n2092# 0.018434f
C17 drain_left.n2 a_n968_n2092# 0.009905f
C18 drain_left.n3 a_n968_n2092# 0.023413f
C19 drain_left.n4 a_n968_n2092# 0.010488f
C20 drain_left.n5 a_n968_n2092# 0.018434f
C21 drain_left.n6 a_n968_n2092# 0.009905f
C22 drain_left.n7 a_n968_n2092# 0.023413f
C23 drain_left.n8 a_n968_n2092# 0.010488f
C24 drain_left.n9 a_n968_n2092# 0.078883f
C25 drain_left.t0 a_n968_n2092# 0.03816f
C26 drain_left.n10 a_n968_n2092# 0.01756f
C27 drain_left.n11 a_n968_n2092# 0.01383f
C28 drain_left.n12 a_n968_n2092# 0.009905f
C29 drain_left.n13 a_n968_n2092# 0.438609f
C30 drain_left.n14 a_n968_n2092# 0.018434f
C31 drain_left.n15 a_n968_n2092# 0.009905f
C32 drain_left.n16 a_n968_n2092# 0.010488f
C33 drain_left.n17 a_n968_n2092# 0.023413f
C34 drain_left.n18 a_n968_n2092# 0.023413f
C35 drain_left.n19 a_n968_n2092# 0.010488f
C36 drain_left.n20 a_n968_n2092# 0.009905f
C37 drain_left.n21 a_n968_n2092# 0.018434f
C38 drain_left.n22 a_n968_n2092# 0.018434f
C39 drain_left.n23 a_n968_n2092# 0.009905f
C40 drain_left.n24 a_n968_n2092# 0.010488f
C41 drain_left.n25 a_n968_n2092# 0.023413f
C42 drain_left.n26 a_n968_n2092# 0.050685f
C43 drain_left.n27 a_n968_n2092# 0.010488f
C44 drain_left.n28 a_n968_n2092# 0.009905f
C45 drain_left.n29 a_n968_n2092# 0.042608f
C46 drain_left.n30 a_n968_n2092# 0.207935f
C47 drain_left.n31 a_n968_n2092# 0.02591f
C48 drain_left.n32 a_n968_n2092# 0.018434f
C49 drain_left.n33 a_n968_n2092# 0.009905f
C50 drain_left.n34 a_n968_n2092# 0.023413f
C51 drain_left.n35 a_n968_n2092# 0.010488f
C52 drain_left.n36 a_n968_n2092# 0.018434f
C53 drain_left.n37 a_n968_n2092# 0.009905f
C54 drain_left.n38 a_n968_n2092# 0.023413f
C55 drain_left.n39 a_n968_n2092# 0.010488f
C56 drain_left.n40 a_n968_n2092# 0.078883f
C57 drain_left.t1 a_n968_n2092# 0.03816f
C58 drain_left.n41 a_n968_n2092# 0.01756f
C59 drain_left.n42 a_n968_n2092# 0.01383f
C60 drain_left.n43 a_n968_n2092# 0.009905f
C61 drain_left.n44 a_n968_n2092# 0.438609f
C62 drain_left.n45 a_n968_n2092# 0.018434f
C63 drain_left.n46 a_n968_n2092# 0.009905f
C64 drain_left.n47 a_n968_n2092# 0.010488f
C65 drain_left.n48 a_n968_n2092# 0.023413f
C66 drain_left.n49 a_n968_n2092# 0.023413f
C67 drain_left.n50 a_n968_n2092# 0.010488f
C68 drain_left.n51 a_n968_n2092# 0.009905f
C69 drain_left.n52 a_n968_n2092# 0.018434f
C70 drain_left.n53 a_n968_n2092# 0.018434f
C71 drain_left.n54 a_n968_n2092# 0.009905f
C72 drain_left.n55 a_n968_n2092# 0.010488f
C73 drain_left.n56 a_n968_n2092# 0.023413f
C74 drain_left.n57 a_n968_n2092# 0.050685f
C75 drain_left.n58 a_n968_n2092# 0.010488f
C76 drain_left.n59 a_n968_n2092# 0.009905f
C77 drain_left.n60 a_n968_n2092# 0.042608f
C78 drain_left.n61 a_n968_n2092# 0.065978f
C79 plus.t0 a_n968_n2092# 0.268054f
C80 plus.t1 a_n968_n2092# 0.29421f
C81 drain_right.n0 a_n968_n2092# 0.026374f
C82 drain_right.n1 a_n968_n2092# 0.018764f
C83 drain_right.n2 a_n968_n2092# 0.010083f
C84 drain_right.n3 a_n968_n2092# 0.023832f
C85 drain_right.n4 a_n968_n2092# 0.010676f
C86 drain_right.n5 a_n968_n2092# 0.018764f
C87 drain_right.n6 a_n968_n2092# 0.010083f
C88 drain_right.n7 a_n968_n2092# 0.023832f
C89 drain_right.n8 a_n968_n2092# 0.010676f
C90 drain_right.n9 a_n968_n2092# 0.080295f
C91 drain_right.t0 a_n968_n2092# 0.038843f
C92 drain_right.n10 a_n968_n2092# 0.017874f
C93 drain_right.n11 a_n968_n2092# 0.014077f
C94 drain_right.n12 a_n968_n2092# 0.010083f
C95 drain_right.n13 a_n968_n2092# 0.446462f
C96 drain_right.n14 a_n968_n2092# 0.018764f
C97 drain_right.n15 a_n968_n2092# 0.010083f
C98 drain_right.n16 a_n968_n2092# 0.010676f
C99 drain_right.n17 a_n968_n2092# 0.023832f
C100 drain_right.n18 a_n968_n2092# 0.023832f
C101 drain_right.n19 a_n968_n2092# 0.010676f
C102 drain_right.n20 a_n968_n2092# 0.010083f
C103 drain_right.n21 a_n968_n2092# 0.018764f
C104 drain_right.n22 a_n968_n2092# 0.018764f
C105 drain_right.n23 a_n968_n2092# 0.010083f
C106 drain_right.n24 a_n968_n2092# 0.010676f
C107 drain_right.n25 a_n968_n2092# 0.023832f
C108 drain_right.n26 a_n968_n2092# 0.051592f
C109 drain_right.n27 a_n968_n2092# 0.010676f
C110 drain_right.n28 a_n968_n2092# 0.010083f
C111 drain_right.n29 a_n968_n2092# 0.043371f
C112 drain_right.n30 a_n968_n2092# 0.19658f
C113 drain_right.n31 a_n968_n2092# 0.026374f
C114 drain_right.n32 a_n968_n2092# 0.018764f
C115 drain_right.n33 a_n968_n2092# 0.010083f
C116 drain_right.n34 a_n968_n2092# 0.023832f
C117 drain_right.n35 a_n968_n2092# 0.010676f
C118 drain_right.n36 a_n968_n2092# 0.018764f
C119 drain_right.n37 a_n968_n2092# 0.010083f
C120 drain_right.n38 a_n968_n2092# 0.023832f
C121 drain_right.n39 a_n968_n2092# 0.010676f
C122 drain_right.n40 a_n968_n2092# 0.080295f
C123 drain_right.t1 a_n968_n2092# 0.038843f
C124 drain_right.n41 a_n968_n2092# 0.017874f
C125 drain_right.n42 a_n968_n2092# 0.014077f
C126 drain_right.n43 a_n968_n2092# 0.010083f
C127 drain_right.n44 a_n968_n2092# 0.446462f
C128 drain_right.n45 a_n968_n2092# 0.018764f
C129 drain_right.n46 a_n968_n2092# 0.010083f
C130 drain_right.n47 a_n968_n2092# 0.010676f
C131 drain_right.n48 a_n968_n2092# 0.023832f
C132 drain_right.n49 a_n968_n2092# 0.023832f
C133 drain_right.n50 a_n968_n2092# 0.010676f
C134 drain_right.n51 a_n968_n2092# 0.010083f
C135 drain_right.n52 a_n968_n2092# 0.018764f
C136 drain_right.n53 a_n968_n2092# 0.018764f
C137 drain_right.n54 a_n968_n2092# 0.010083f
C138 drain_right.n55 a_n968_n2092# 0.010676f
C139 drain_right.n56 a_n968_n2092# 0.023832f
C140 drain_right.n57 a_n968_n2092# 0.051592f
C141 drain_right.n58 a_n968_n2092# 0.010676f
C142 drain_right.n59 a_n968_n2092# 0.010083f
C143 drain_right.n60 a_n968_n2092# 0.043371f
C144 drain_right.n61 a_n968_n2092# 0.067024f
C145 source.n0 a_n968_n2092# 0.029508f
C146 source.n1 a_n968_n2092# 0.020994f
C147 source.n2 a_n968_n2092# 0.011281f
C148 source.n3 a_n968_n2092# 0.026664f
C149 source.n4 a_n968_n2092# 0.011945f
C150 source.n5 a_n968_n2092# 0.020994f
C151 source.n6 a_n968_n2092# 0.011281f
C152 source.n7 a_n968_n2092# 0.026664f
C153 source.n8 a_n968_n2092# 0.011945f
C154 source.n9 a_n968_n2092# 0.089838f
C155 source.t1 a_n968_n2092# 0.043459f
C156 source.n10 a_n968_n2092# 0.019998f
C157 source.n11 a_n968_n2092# 0.01575f
C158 source.n12 a_n968_n2092# 0.011281f
C159 source.n13 a_n968_n2092# 0.499521f
C160 source.n14 a_n968_n2092# 0.020994f
C161 source.n15 a_n968_n2092# 0.011281f
C162 source.n16 a_n968_n2092# 0.011945f
C163 source.n17 a_n968_n2092# 0.026664f
C164 source.n18 a_n968_n2092# 0.026664f
C165 source.n19 a_n968_n2092# 0.011945f
C166 source.n20 a_n968_n2092# 0.011281f
C167 source.n21 a_n968_n2092# 0.020994f
C168 source.n22 a_n968_n2092# 0.020994f
C169 source.n23 a_n968_n2092# 0.011281f
C170 source.n24 a_n968_n2092# 0.011945f
C171 source.n25 a_n968_n2092# 0.026664f
C172 source.n26 a_n968_n2092# 0.057724f
C173 source.n27 a_n968_n2092# 0.011945f
C174 source.n28 a_n968_n2092# 0.011281f
C175 source.n29 a_n968_n2092# 0.048526f
C176 source.n30 a_n968_n2092# 0.032299f
C177 source.n31 a_n968_n2092# 0.522969f
C178 source.n32 a_n968_n2092# 0.029508f
C179 source.n33 a_n968_n2092# 0.020994f
C180 source.n34 a_n968_n2092# 0.011281f
C181 source.n35 a_n968_n2092# 0.026664f
C182 source.n36 a_n968_n2092# 0.011945f
C183 source.n37 a_n968_n2092# 0.020994f
C184 source.n38 a_n968_n2092# 0.011281f
C185 source.n39 a_n968_n2092# 0.026664f
C186 source.n40 a_n968_n2092# 0.011945f
C187 source.n41 a_n968_n2092# 0.089838f
C188 source.t2 a_n968_n2092# 0.043459f
C189 source.n42 a_n968_n2092# 0.019998f
C190 source.n43 a_n968_n2092# 0.01575f
C191 source.n44 a_n968_n2092# 0.011281f
C192 source.n45 a_n968_n2092# 0.499521f
C193 source.n46 a_n968_n2092# 0.020994f
C194 source.n47 a_n968_n2092# 0.011281f
C195 source.n48 a_n968_n2092# 0.011945f
C196 source.n49 a_n968_n2092# 0.026664f
C197 source.n50 a_n968_n2092# 0.026664f
C198 source.n51 a_n968_n2092# 0.011945f
C199 source.n52 a_n968_n2092# 0.011281f
C200 source.n53 a_n968_n2092# 0.020994f
C201 source.n54 a_n968_n2092# 0.020994f
C202 source.n55 a_n968_n2092# 0.011281f
C203 source.n56 a_n968_n2092# 0.011945f
C204 source.n57 a_n968_n2092# 0.026664f
C205 source.n58 a_n968_n2092# 0.057724f
C206 source.n59 a_n968_n2092# 0.011945f
C207 source.n60 a_n968_n2092# 0.011281f
C208 source.n61 a_n968_n2092# 0.048526f
C209 source.n62 a_n968_n2092# 0.032299f
C210 source.n63 a_n968_n2092# 0.830255f
C211 source.n64 a_n968_n2092# 0.029508f
C212 source.n65 a_n968_n2092# 0.020994f
C213 source.n66 a_n968_n2092# 0.011281f
C214 source.n67 a_n968_n2092# 0.026664f
C215 source.n68 a_n968_n2092# 0.011945f
C216 source.n69 a_n968_n2092# 0.020994f
C217 source.n70 a_n968_n2092# 0.011281f
C218 source.n71 a_n968_n2092# 0.026664f
C219 source.n72 a_n968_n2092# 0.011945f
C220 source.n73 a_n968_n2092# 0.089838f
C221 source.t0 a_n968_n2092# 0.043459f
C222 source.n74 a_n968_n2092# 0.019998f
C223 source.n75 a_n968_n2092# 0.01575f
C224 source.n76 a_n968_n2092# 0.011281f
C225 source.n77 a_n968_n2092# 0.499521f
C226 source.n78 a_n968_n2092# 0.020994f
C227 source.n79 a_n968_n2092# 0.011281f
C228 source.n80 a_n968_n2092# 0.011945f
C229 source.n81 a_n968_n2092# 0.026664f
C230 source.n82 a_n968_n2092# 0.026664f
C231 source.n83 a_n968_n2092# 0.011945f
C232 source.n84 a_n968_n2092# 0.011281f
C233 source.n85 a_n968_n2092# 0.020994f
C234 source.n86 a_n968_n2092# 0.020994f
C235 source.n87 a_n968_n2092# 0.011281f
C236 source.n88 a_n968_n2092# 0.011945f
C237 source.n89 a_n968_n2092# 0.026664f
C238 source.n90 a_n968_n2092# 0.057724f
C239 source.n91 a_n968_n2092# 0.011945f
C240 source.n92 a_n968_n2092# 0.011281f
C241 source.n93 a_n968_n2092# 0.048526f
C242 source.n94 a_n968_n2092# 0.032299f
C243 source.n95 a_n968_n2092# 0.830254f
C244 source.n96 a_n968_n2092# 0.029508f
C245 source.n97 a_n968_n2092# 0.020994f
C246 source.n98 a_n968_n2092# 0.011281f
C247 source.n99 a_n968_n2092# 0.026664f
C248 source.n100 a_n968_n2092# 0.011945f
C249 source.n101 a_n968_n2092# 0.020994f
C250 source.n102 a_n968_n2092# 0.011281f
C251 source.n103 a_n968_n2092# 0.026664f
C252 source.n104 a_n968_n2092# 0.011945f
C253 source.n105 a_n968_n2092# 0.089838f
C254 source.t3 a_n968_n2092# 0.043459f
C255 source.n106 a_n968_n2092# 0.019998f
C256 source.n107 a_n968_n2092# 0.01575f
C257 source.n108 a_n968_n2092# 0.011281f
C258 source.n109 a_n968_n2092# 0.499521f
C259 source.n110 a_n968_n2092# 0.020994f
C260 source.n111 a_n968_n2092# 0.011281f
C261 source.n112 a_n968_n2092# 0.011945f
C262 source.n113 a_n968_n2092# 0.026664f
C263 source.n114 a_n968_n2092# 0.026664f
C264 source.n115 a_n968_n2092# 0.011945f
C265 source.n116 a_n968_n2092# 0.011281f
C266 source.n117 a_n968_n2092# 0.020994f
C267 source.n118 a_n968_n2092# 0.020994f
C268 source.n119 a_n968_n2092# 0.011281f
C269 source.n120 a_n968_n2092# 0.011945f
C270 source.n121 a_n968_n2092# 0.026664f
C271 source.n122 a_n968_n2092# 0.057724f
C272 source.n123 a_n968_n2092# 0.011945f
C273 source.n124 a_n968_n2092# 0.011281f
C274 source.n125 a_n968_n2092# 0.048526f
C275 source.n126 a_n968_n2092# 0.032299f
C276 source.n127 a_n968_n2092# 0.218372f
C277 source.n128 a_n968_n2092# 0.860623f
C278 minus.t0 a_n968_n2092# 0.294304f
C279 minus.t1 a_n968_n2092# 0.258053f
C280 minus.n0 a_n968_n2092# 2.71832f
.ends

