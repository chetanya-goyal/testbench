* NGSPICE file created from diffpair431.ext - technology: sky130A

.subckt diffpair431 minus drain_right drain_left source plus
X0 drain_right minus source a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X1 drain_right minus source a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X2 source minus drain_right a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X3 drain_left plus source a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X4 a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.3
X5 a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X6 source minus drain_right a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X7 a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X8 a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X9 source plus drain_left a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X10 drain_left plus source a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X11 source plus drain_left a_n1094_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
.ends

