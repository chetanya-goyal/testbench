* NGSPICE file created from diffpair622.ext - technology: sky130A

.subckt diffpair622 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t11 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 drain_right.t5 minus.t0 source.t5 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X2 source.t6 plus.t1 drain_left.t4 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 drain_left.t3 plus.t2 source.t9 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X4 source.t0 minus.t1 drain_right.t4 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X5 drain_left.t2 plus.t3 source.t10 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X6 source.t1 minus.t2 drain_right.t3 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 drain_right.t2 minus.t3 source.t4 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X8 a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X9 a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X10 drain_right.t1 minus.t4 source.t3 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X11 a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X12 drain_right.t0 minus.t5 source.t2 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X13 source.t8 plus.t4 drain_left.t1 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X14 a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X15 drain_left.t0 plus.t5 source.t7 a_n1540_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n1 plus.t3 766.284
R1 plus.n7 plus.t0 766.284
R2 plus.n4 plus.t2 744.691
R3 plus.n2 plus.t4 744.691
R4 plus.n10 plus.t5 744.691
R5 plus.n8 plus.t1 744.691
R6 plus.n3 plus.n0 161.3
R7 plus.n5 plus.n4 161.3
R8 plus.n9 plus.n6 161.3
R9 plus.n11 plus.n10 161.3
R10 plus.n1 plus.n0 44.8545
R11 plus.n7 plus.n6 44.8545
R12 plus plus.n11 31.9933
R13 plus.n4 plus.n3 26.2914
R14 plus.n10 plus.n9 26.2914
R15 plus.n3 plus.n2 21.9096
R16 plus.n9 plus.n8 21.9096
R17 plus.n2 plus.n1 20.3348
R18 plus.n8 plus.n7 20.3348
R19 plus plus.n5 15.3016
R20 plus.n5 plus.n0 0.189894
R21 plus.n11 plus.n6 0.189894
R22 source.n0 source.t9 44.1297
R23 source.n3 source.t2 44.1296
R24 source.n11 source.t5 44.1295
R25 source.n8 source.t11 44.1295
R26 source.n2 source.n1 43.1397
R27 source.n5 source.n4 43.1397
R28 source.n10 source.n9 43.1396
R29 source.n7 source.n6 43.1396
R30 source.n7 source.n5 29.1242
R31 source.n12 source.n0 22.5294
R32 source.n12 source.n11 5.7074
R33 source.n9 source.t4 0.9905
R34 source.n9 source.t1 0.9905
R35 source.n6 source.t7 0.9905
R36 source.n6 source.t6 0.9905
R37 source.n1 source.t10 0.9905
R38 source.n1 source.t8 0.9905
R39 source.n4 source.t3 0.9905
R40 source.n4 source.t0 0.9905
R41 source.n3 source.n2 0.914293
R42 source.n10 source.n8 0.914293
R43 source.n5 source.n3 0.888431
R44 source.n2 source.n0 0.888431
R45 source.n8 source.n7 0.888431
R46 source.n11 source.n10 0.888431
R47 source source.n12 0.188
R48 drain_left.n3 drain_left.t2 61.6963
R49 drain_left.n1 drain_left.t0 61.4189
R50 drain_left.n1 drain_left.n0 59.985
R51 drain_left.n3 drain_left.n2 59.8185
R52 drain_left drain_left.n1 35.8695
R53 drain_left drain_left.n3 6.54115
R54 drain_left.n0 drain_left.t4 0.9905
R55 drain_left.n0 drain_left.t5 0.9905
R56 drain_left.n2 drain_left.t1 0.9905
R57 drain_left.n2 drain_left.t3 0.9905
R58 minus.n1 minus.t5 766.284
R59 minus.n7 minus.t3 766.284
R60 minus.n2 minus.t1 744.691
R61 minus.n4 minus.t4 744.691
R62 minus.n8 minus.t2 744.691
R63 minus.n10 minus.t0 744.691
R64 minus.n5 minus.n4 161.3
R65 minus.n3 minus.n0 161.3
R66 minus.n11 minus.n10 161.3
R67 minus.n9 minus.n6 161.3
R68 minus.n1 minus.n0 44.8545
R69 minus.n7 minus.n6 44.8545
R70 minus.n12 minus.n5 41.1425
R71 minus.n4 minus.n3 26.2914
R72 minus.n10 minus.n9 26.2914
R73 minus.n3 minus.n2 21.9096
R74 minus.n9 minus.n8 21.9096
R75 minus.n2 minus.n1 20.3348
R76 minus.n8 minus.n7 20.3348
R77 minus.n12 minus.n11 6.62739
R78 minus.n5 minus.n0 0.189894
R79 minus.n11 minus.n6 0.189894
R80 minus minus.n12 0.188
R81 drain_right.n1 drain_right.t2 61.4189
R82 drain_right.n3 drain_right.t1 60.8084
R83 drain_right.n3 drain_right.n2 60.7064
R84 drain_right.n1 drain_right.n0 59.985
R85 drain_right drain_right.n1 35.3163
R86 drain_right drain_right.n3 6.09718
R87 drain_right.n0 drain_right.t3 0.9905
R88 drain_right.n0 drain_right.t5 0.9905
R89 drain_right.n2 drain_right.t4 0.9905
R90 drain_right.n2 drain_right.t0 0.9905
C0 drain_left source 15.524402f
C1 drain_right source 15.5123f
C2 plus source 6.40305f
C3 drain_left minus 0.171172f
C4 drain_right minus 7.03731f
C5 plus minus 6.5432f
C6 source minus 6.38818f
C7 drain_right drain_left 0.71116f
C8 drain_left plus 7.1808f
C9 drain_right plus 0.304583f
C10 drain_right a_n1540_n4888# 8.466479f
C11 drain_left a_n1540_n4888# 8.71325f
C12 source a_n1540_n4888# 9.377603f
C13 minus a_n1540_n4888# 6.428829f
C14 plus a_n1540_n4888# 8.5907f
C15 drain_right.t2 a_n1540_n4888# 4.27051f
C16 drain_right.t3 a_n1540_n4888# 0.364968f
C17 drain_right.t5 a_n1540_n4888# 0.364968f
C18 drain_right.n0 a_n1540_n4888# 3.33741f
C19 drain_right.n1 a_n1540_n4888# 2.0802f
C20 drain_right.t4 a_n1540_n4888# 0.364968f
C21 drain_right.t0 a_n1540_n4888# 0.364968f
C22 drain_right.n2 a_n1540_n4888# 3.34153f
C23 drain_right.t1 a_n1540_n4888# 4.2674f
C24 drain_right.n3 a_n1540_n4888# 0.87845f
C25 minus.n0 a_n1540_n4888# 0.188316f
C26 minus.t5 a_n1540_n4888# 1.82227f
C27 minus.n1 a_n1540_n4888# 0.657704f
C28 minus.t1 a_n1540_n4888# 1.80333f
C29 minus.n2 a_n1540_n4888# 0.676137f
C30 minus.n3 a_n1540_n4888# 0.010321f
C31 minus.t4 a_n1540_n4888# 1.80333f
C32 minus.n4 a_n1540_n4888# 0.66909f
C33 minus.n5 a_n1540_n4888# 1.95781f
C34 minus.n6 a_n1540_n4888# 0.188316f
C35 minus.t3 a_n1540_n4888# 1.82227f
C36 minus.n7 a_n1540_n4888# 0.657704f
C37 minus.t2 a_n1540_n4888# 1.80333f
C38 minus.n8 a_n1540_n4888# 0.676137f
C39 minus.n9 a_n1540_n4888# 0.010321f
C40 minus.t0 a_n1540_n4888# 1.80333f
C41 minus.n10 a_n1540_n4888# 0.66909f
C42 minus.n11 a_n1540_n4888# 0.31094f
C43 minus.n12 a_n1540_n4888# 2.34038f
C44 drain_left.t0 a_n1540_n4888# 4.29124f
C45 drain_left.t4 a_n1540_n4888# 0.366739f
C46 drain_left.t5 a_n1540_n4888# 0.366739f
C47 drain_left.n0 a_n1540_n4888# 3.35361f
C48 drain_left.n1 a_n1540_n4888# 2.13884f
C49 drain_left.t2 a_n1540_n4888# 4.29296f
C50 drain_left.t1 a_n1540_n4888# 0.366739f
C51 drain_left.t3 a_n1540_n4888# 0.366739f
C52 drain_left.n2 a_n1540_n4888# 3.35281f
C53 drain_left.n3 a_n1540_n4888# 0.865452f
C54 source.t9 a_n1540_n4888# 4.22245f
C55 source.n0 a_n1540_n4888# 1.83688f
C56 source.t10 a_n1540_n4888# 0.36947f
C57 source.t8 a_n1540_n4888# 0.36947f
C58 source.n1 a_n1540_n4888# 3.30322f
C59 source.n2 a_n1540_n4888# 0.375772f
C60 source.t2 a_n1540_n4888# 4.22246f
C61 source.n3 a_n1540_n4888# 0.464185f
C62 source.t3 a_n1540_n4888# 0.36947f
C63 source.t0 a_n1540_n4888# 0.36947f
C64 source.n4 a_n1540_n4888# 3.30322f
C65 source.n5 a_n1540_n4888# 2.24065f
C66 source.t7 a_n1540_n4888# 0.36947f
C67 source.t6 a_n1540_n4888# 0.36947f
C68 source.n6 a_n1540_n4888# 3.30323f
C69 source.n7 a_n1540_n4888# 2.24064f
C70 source.t11 a_n1540_n4888# 4.22243f
C71 source.n8 a_n1540_n4888# 0.464208f
C72 source.t4 a_n1540_n4888# 0.36947f
C73 source.t1 a_n1540_n4888# 0.36947f
C74 source.n9 a_n1540_n4888# 3.30323f
C75 source.n10 a_n1540_n4888# 0.375766f
C76 source.t5 a_n1540_n4888# 4.22243f
C77 source.n11 a_n1540_n4888# 0.583257f
C78 source.n12 a_n1540_n4888# 2.12087f
C79 plus.n0 a_n1540_n4888# 0.191092f
C80 plus.t2 a_n1540_n4888# 1.82991f
C81 plus.t4 a_n1540_n4888# 1.82991f
C82 plus.t3 a_n1540_n4888# 1.84913f
C83 plus.n1 a_n1540_n4888# 0.667399f
C84 plus.n2 a_n1540_n4888# 0.686104f
C85 plus.n3 a_n1540_n4888# 0.010474f
C86 plus.n4 a_n1540_n4888# 0.678953f
C87 plus.n5 a_n1540_n4888# 0.714335f
C88 plus.n6 a_n1540_n4888# 0.191092f
C89 plus.t5 a_n1540_n4888# 1.82991f
C90 plus.t0 a_n1540_n4888# 1.84913f
C91 plus.n7 a_n1540_n4888# 0.667399f
C92 plus.t1 a_n1540_n4888# 1.82991f
C93 plus.n8 a_n1540_n4888# 0.686104f
C94 plus.n9 a_n1540_n4888# 0.010474f
C95 plus.n10 a_n1540_n4888# 0.678953f
C96 plus.n11 a_n1540_n4888# 1.56722f
.ends

