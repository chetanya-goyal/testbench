* NGSPICE file created from diffpair254.ext - technology: sky130A

.subckt diffpair254 minus drain_right drain_left source plus
X0 a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X1 drain_right.t9 minus.t0 source.t14 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 drain_right.t8 minus.t1 source.t15 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X3 a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X4 source.t9 plus.t0 drain_left.t9 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X5 a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X6 source.t2 plus.t1 drain_left.t8 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 source.t10 minus.t2 drain_right.t7 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X8 drain_left.t7 plus.t2 source.t1 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X9 drain_left.t6 plus.t3 source.t3 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X10 drain_left.t5 plus.t4 source.t4 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X11 drain_left.t4 plus.t5 source.t5 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X12 drain_right.t6 minus.t3 source.t18 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X13 drain_right.t5 minus.t4 source.t11 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X14 source.t6 plus.t6 drain_left.t3 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X15 drain_left.t2 plus.t7 source.t0 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X16 source.t8 plus.t8 drain_left.t1 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X17 drain_right.t4 minus.t5 source.t17 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X18 drain_right.t3 minus.t6 source.t12 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X19 source.t13 minus.t7 drain_right.t2 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X20 a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X21 source.t16 minus.t8 drain_right.t1 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X22 source.t19 minus.t9 drain_right.t0 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X23 drain_left.t0 plus.t9 source.t7 a_n1352_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n8 minus.t4 924.929
R1 minus.n2 minus.t3 924.929
R2 minus.n18 minus.t1 924.929
R3 minus.n12 minus.t6 924.929
R4 minus.n7 minus.t7 879.65
R5 minus.n5 minus.t0 879.65
R6 minus.n1 minus.t2 879.65
R7 minus.n17 minus.t8 879.65
R8 minus.n15 minus.t5 879.65
R9 minus.n11 minus.t9 879.65
R10 minus.n3 minus.n2 161.489
R11 minus.n13 minus.n12 161.489
R12 minus.n9 minus.n8 161.3
R13 minus.n6 minus.n0 161.3
R14 minus.n4 minus.n3 161.3
R15 minus.n19 minus.n18 161.3
R16 minus.n16 minus.n10 161.3
R17 minus.n14 minus.n13 161.3
R18 minus.n7 minus.n6 40.8975
R19 minus.n4 minus.n1 40.8975
R20 minus.n14 minus.n11 40.8975
R21 minus.n17 minus.n16 40.8975
R22 minus.n6 minus.n5 36.5157
R23 minus.n5 minus.n4 36.5157
R24 minus.n15 minus.n14 36.5157
R25 minus.n16 minus.n15 36.5157
R26 minus.n8 minus.n7 32.1338
R27 minus.n2 minus.n1 32.1338
R28 minus.n12 minus.n11 32.1338
R29 minus.n18 minus.n17 32.1338
R30 minus.n20 minus.n9 29.6463
R31 minus.n20 minus.n19 6.44936
R32 minus.n9 minus.n0 0.189894
R33 minus.n3 minus.n0 0.189894
R34 minus.n13 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n138 source.n112 289.615
R38 source.n102 source.n76 289.615
R39 source.n26 source.n0 289.615
R40 source.n62 source.n36 289.615
R41 source.n123 source.n122 185
R42 source.n120 source.n119 185
R43 source.n129 source.n128 185
R44 source.n131 source.n130 185
R45 source.n116 source.n115 185
R46 source.n137 source.n136 185
R47 source.n139 source.n138 185
R48 source.n87 source.n86 185
R49 source.n84 source.n83 185
R50 source.n93 source.n92 185
R51 source.n95 source.n94 185
R52 source.n80 source.n79 185
R53 source.n101 source.n100 185
R54 source.n103 source.n102 185
R55 source.n27 source.n26 185
R56 source.n25 source.n24 185
R57 source.n4 source.n3 185
R58 source.n19 source.n18 185
R59 source.n17 source.n16 185
R60 source.n8 source.n7 185
R61 source.n11 source.n10 185
R62 source.n63 source.n62 185
R63 source.n61 source.n60 185
R64 source.n40 source.n39 185
R65 source.n55 source.n54 185
R66 source.n53 source.n52 185
R67 source.n44 source.n43 185
R68 source.n47 source.n46 185
R69 source.t15 source.n121 147.661
R70 source.t5 source.n85 147.661
R71 source.t0 source.n9 147.661
R72 source.t18 source.n45 147.661
R73 source.n122 source.n119 104.615
R74 source.n129 source.n119 104.615
R75 source.n130 source.n129 104.615
R76 source.n130 source.n115 104.615
R77 source.n137 source.n115 104.615
R78 source.n138 source.n137 104.615
R79 source.n86 source.n83 104.615
R80 source.n93 source.n83 104.615
R81 source.n94 source.n93 104.615
R82 source.n94 source.n79 104.615
R83 source.n101 source.n79 104.615
R84 source.n102 source.n101 104.615
R85 source.n26 source.n25 104.615
R86 source.n25 source.n3 104.615
R87 source.n18 source.n3 104.615
R88 source.n18 source.n17 104.615
R89 source.n17 source.n7 104.615
R90 source.n10 source.n7 104.615
R91 source.n62 source.n61 104.615
R92 source.n61 source.n39 104.615
R93 source.n54 source.n39 104.615
R94 source.n54 source.n53 104.615
R95 source.n53 source.n43 104.615
R96 source.n46 source.n43 104.615
R97 source.n122 source.t15 52.3082
R98 source.n86 source.t5 52.3082
R99 source.n10 source.t0 52.3082
R100 source.n46 source.t18 52.3082
R101 source.n33 source.n32 50.512
R102 source.n35 source.n34 50.512
R103 source.n69 source.n68 50.512
R104 source.n71 source.n70 50.512
R105 source.n111 source.n110 50.5119
R106 source.n109 source.n108 50.5119
R107 source.n75 source.n74 50.5119
R108 source.n73 source.n72 50.5119
R109 source.n143 source.n142 32.1853
R110 source.n107 source.n106 32.1853
R111 source.n31 source.n30 32.1853
R112 source.n67 source.n66 32.1853
R113 source.n73 source.n71 17.6561
R114 source.n123 source.n121 15.6674
R115 source.n87 source.n85 15.6674
R116 source.n11 source.n9 15.6674
R117 source.n47 source.n45 15.6674
R118 source.n124 source.n120 12.8005
R119 source.n88 source.n84 12.8005
R120 source.n12 source.n8 12.8005
R121 source.n48 source.n44 12.8005
R122 source.n128 source.n127 12.0247
R123 source.n92 source.n91 12.0247
R124 source.n16 source.n15 12.0247
R125 source.n52 source.n51 12.0247
R126 source.n144 source.n31 11.7078
R127 source.n131 source.n118 11.249
R128 source.n95 source.n82 11.249
R129 source.n19 source.n6 11.249
R130 source.n55 source.n42 11.249
R131 source.n132 source.n116 10.4732
R132 source.n96 source.n80 10.4732
R133 source.n20 source.n4 10.4732
R134 source.n56 source.n40 10.4732
R135 source.n136 source.n135 9.69747
R136 source.n100 source.n99 9.69747
R137 source.n24 source.n23 9.69747
R138 source.n60 source.n59 9.69747
R139 source.n142 source.n141 9.45567
R140 source.n106 source.n105 9.45567
R141 source.n30 source.n29 9.45567
R142 source.n66 source.n65 9.45567
R143 source.n141 source.n140 9.3005
R144 source.n114 source.n113 9.3005
R145 source.n135 source.n134 9.3005
R146 source.n133 source.n132 9.3005
R147 source.n118 source.n117 9.3005
R148 source.n127 source.n126 9.3005
R149 source.n125 source.n124 9.3005
R150 source.n105 source.n104 9.3005
R151 source.n78 source.n77 9.3005
R152 source.n99 source.n98 9.3005
R153 source.n97 source.n96 9.3005
R154 source.n82 source.n81 9.3005
R155 source.n91 source.n90 9.3005
R156 source.n89 source.n88 9.3005
R157 source.n29 source.n28 9.3005
R158 source.n2 source.n1 9.3005
R159 source.n23 source.n22 9.3005
R160 source.n21 source.n20 9.3005
R161 source.n6 source.n5 9.3005
R162 source.n15 source.n14 9.3005
R163 source.n13 source.n12 9.3005
R164 source.n65 source.n64 9.3005
R165 source.n38 source.n37 9.3005
R166 source.n59 source.n58 9.3005
R167 source.n57 source.n56 9.3005
R168 source.n42 source.n41 9.3005
R169 source.n51 source.n50 9.3005
R170 source.n49 source.n48 9.3005
R171 source.n139 source.n114 8.92171
R172 source.n103 source.n78 8.92171
R173 source.n27 source.n2 8.92171
R174 source.n63 source.n38 8.92171
R175 source.n140 source.n112 8.14595
R176 source.n104 source.n76 8.14595
R177 source.n28 source.n0 8.14595
R178 source.n64 source.n36 8.14595
R179 source.n142 source.n112 5.81868
R180 source.n106 source.n76 5.81868
R181 source.n30 source.n0 5.81868
R182 source.n66 source.n36 5.81868
R183 source.n144 source.n143 5.49188
R184 source.n140 source.n139 5.04292
R185 source.n104 source.n103 5.04292
R186 source.n28 source.n27 5.04292
R187 source.n64 source.n63 5.04292
R188 source.n125 source.n121 4.38594
R189 source.n89 source.n85 4.38594
R190 source.n13 source.n9 4.38594
R191 source.n49 source.n45 4.38594
R192 source.n136 source.n114 4.26717
R193 source.n100 source.n78 4.26717
R194 source.n24 source.n2 4.26717
R195 source.n60 source.n38 4.26717
R196 source.n135 source.n116 3.49141
R197 source.n99 source.n80 3.49141
R198 source.n23 source.n4 3.49141
R199 source.n59 source.n40 3.49141
R200 source.n110 source.t17 3.3005
R201 source.n110 source.t16 3.3005
R202 source.n108 source.t12 3.3005
R203 source.n108 source.t19 3.3005
R204 source.n74 source.t3 3.3005
R205 source.n74 source.t6 3.3005
R206 source.n72 source.t4 3.3005
R207 source.n72 source.t2 3.3005
R208 source.n32 source.t7 3.3005
R209 source.n32 source.t8 3.3005
R210 source.n34 source.t1 3.3005
R211 source.n34 source.t9 3.3005
R212 source.n68 source.t14 3.3005
R213 source.n68 source.t10 3.3005
R214 source.n70 source.t11 3.3005
R215 source.n70 source.t13 3.3005
R216 source.n132 source.n131 2.71565
R217 source.n96 source.n95 2.71565
R218 source.n20 source.n19 2.71565
R219 source.n56 source.n55 2.71565
R220 source.n128 source.n118 1.93989
R221 source.n92 source.n82 1.93989
R222 source.n16 source.n6 1.93989
R223 source.n52 source.n42 1.93989
R224 source.n127 source.n120 1.16414
R225 source.n91 source.n84 1.16414
R226 source.n15 source.n8 1.16414
R227 source.n51 source.n44 1.16414
R228 source.n67 source.n35 0.698776
R229 source.n109 source.n107 0.698776
R230 source.n71 source.n69 0.457397
R231 source.n69 source.n67 0.457397
R232 source.n35 source.n33 0.457397
R233 source.n33 source.n31 0.457397
R234 source.n75 source.n73 0.457397
R235 source.n107 source.n75 0.457397
R236 source.n111 source.n109 0.457397
R237 source.n143 source.n111 0.457397
R238 source.n124 source.n123 0.388379
R239 source.n88 source.n87 0.388379
R240 source.n12 source.n11 0.388379
R241 source.n48 source.n47 0.388379
R242 source source.n144 0.188
R243 source.n126 source.n125 0.155672
R244 source.n126 source.n117 0.155672
R245 source.n133 source.n117 0.155672
R246 source.n134 source.n133 0.155672
R247 source.n134 source.n113 0.155672
R248 source.n141 source.n113 0.155672
R249 source.n90 source.n89 0.155672
R250 source.n90 source.n81 0.155672
R251 source.n97 source.n81 0.155672
R252 source.n98 source.n97 0.155672
R253 source.n98 source.n77 0.155672
R254 source.n105 source.n77 0.155672
R255 source.n29 source.n1 0.155672
R256 source.n22 source.n1 0.155672
R257 source.n22 source.n21 0.155672
R258 source.n21 source.n5 0.155672
R259 source.n14 source.n5 0.155672
R260 source.n14 source.n13 0.155672
R261 source.n65 source.n37 0.155672
R262 source.n58 source.n37 0.155672
R263 source.n58 source.n57 0.155672
R264 source.n57 source.n41 0.155672
R265 source.n50 source.n41 0.155672
R266 source.n50 source.n49 0.155672
R267 drain_right.n26 drain_right.n0 289.615
R268 drain_right.n64 drain_right.n38 289.615
R269 drain_right.n11 drain_right.n10 185
R270 drain_right.n8 drain_right.n7 185
R271 drain_right.n17 drain_right.n16 185
R272 drain_right.n19 drain_right.n18 185
R273 drain_right.n4 drain_right.n3 185
R274 drain_right.n25 drain_right.n24 185
R275 drain_right.n27 drain_right.n26 185
R276 drain_right.n65 drain_right.n64 185
R277 drain_right.n63 drain_right.n62 185
R278 drain_right.n42 drain_right.n41 185
R279 drain_right.n57 drain_right.n56 185
R280 drain_right.n55 drain_right.n54 185
R281 drain_right.n46 drain_right.n45 185
R282 drain_right.n49 drain_right.n48 185
R283 drain_right.t3 drain_right.n9 147.661
R284 drain_right.t5 drain_right.n47 147.661
R285 drain_right.n10 drain_right.n7 104.615
R286 drain_right.n17 drain_right.n7 104.615
R287 drain_right.n18 drain_right.n17 104.615
R288 drain_right.n18 drain_right.n3 104.615
R289 drain_right.n25 drain_right.n3 104.615
R290 drain_right.n26 drain_right.n25 104.615
R291 drain_right.n64 drain_right.n63 104.615
R292 drain_right.n63 drain_right.n41 104.615
R293 drain_right.n56 drain_right.n41 104.615
R294 drain_right.n56 drain_right.n55 104.615
R295 drain_right.n55 drain_right.n45 104.615
R296 drain_right.n48 drain_right.n45 104.615
R297 drain_right.n37 drain_right.n35 67.6476
R298 drain_right.n34 drain_right.n33 67.478
R299 drain_right.n37 drain_right.n36 67.1908
R300 drain_right.n32 drain_right.n31 67.1907
R301 drain_right.n10 drain_right.t3 52.3082
R302 drain_right.n48 drain_right.t5 52.3082
R303 drain_right.n32 drain_right.n30 49.321
R304 drain_right.n69 drain_right.n68 48.8641
R305 drain_right drain_right.n34 24.2102
R306 drain_right.n11 drain_right.n9 15.6674
R307 drain_right.n49 drain_right.n47 15.6674
R308 drain_right.n12 drain_right.n8 12.8005
R309 drain_right.n50 drain_right.n46 12.8005
R310 drain_right.n16 drain_right.n15 12.0247
R311 drain_right.n54 drain_right.n53 12.0247
R312 drain_right.n19 drain_right.n6 11.249
R313 drain_right.n57 drain_right.n44 11.249
R314 drain_right.n20 drain_right.n4 10.4732
R315 drain_right.n58 drain_right.n42 10.4732
R316 drain_right.n24 drain_right.n23 9.69747
R317 drain_right.n62 drain_right.n61 9.69747
R318 drain_right.n30 drain_right.n29 9.45567
R319 drain_right.n68 drain_right.n67 9.45567
R320 drain_right.n29 drain_right.n28 9.3005
R321 drain_right.n2 drain_right.n1 9.3005
R322 drain_right.n23 drain_right.n22 9.3005
R323 drain_right.n21 drain_right.n20 9.3005
R324 drain_right.n6 drain_right.n5 9.3005
R325 drain_right.n15 drain_right.n14 9.3005
R326 drain_right.n13 drain_right.n12 9.3005
R327 drain_right.n67 drain_right.n66 9.3005
R328 drain_right.n40 drain_right.n39 9.3005
R329 drain_right.n61 drain_right.n60 9.3005
R330 drain_right.n59 drain_right.n58 9.3005
R331 drain_right.n44 drain_right.n43 9.3005
R332 drain_right.n53 drain_right.n52 9.3005
R333 drain_right.n51 drain_right.n50 9.3005
R334 drain_right.n27 drain_right.n2 8.92171
R335 drain_right.n65 drain_right.n40 8.92171
R336 drain_right.n28 drain_right.n0 8.14595
R337 drain_right.n66 drain_right.n38 8.14595
R338 drain_right drain_right.n69 5.88166
R339 drain_right.n30 drain_right.n0 5.81868
R340 drain_right.n68 drain_right.n38 5.81868
R341 drain_right.n28 drain_right.n27 5.04292
R342 drain_right.n66 drain_right.n65 5.04292
R343 drain_right.n13 drain_right.n9 4.38594
R344 drain_right.n51 drain_right.n47 4.38594
R345 drain_right.n24 drain_right.n2 4.26717
R346 drain_right.n62 drain_right.n40 4.26717
R347 drain_right.n23 drain_right.n4 3.49141
R348 drain_right.n61 drain_right.n42 3.49141
R349 drain_right.n33 drain_right.t1 3.3005
R350 drain_right.n33 drain_right.t8 3.3005
R351 drain_right.n31 drain_right.t0 3.3005
R352 drain_right.n31 drain_right.t4 3.3005
R353 drain_right.n35 drain_right.t7 3.3005
R354 drain_right.n35 drain_right.t6 3.3005
R355 drain_right.n36 drain_right.t2 3.3005
R356 drain_right.n36 drain_right.t9 3.3005
R357 drain_right.n20 drain_right.n19 2.71565
R358 drain_right.n58 drain_right.n57 2.71565
R359 drain_right.n16 drain_right.n6 1.93989
R360 drain_right.n54 drain_right.n44 1.93989
R361 drain_right.n15 drain_right.n8 1.16414
R362 drain_right.n53 drain_right.n46 1.16414
R363 drain_right.n69 drain_right.n37 0.457397
R364 drain_right.n12 drain_right.n11 0.388379
R365 drain_right.n50 drain_right.n49 0.388379
R366 drain_right.n14 drain_right.n13 0.155672
R367 drain_right.n14 drain_right.n5 0.155672
R368 drain_right.n21 drain_right.n5 0.155672
R369 drain_right.n22 drain_right.n21 0.155672
R370 drain_right.n22 drain_right.n1 0.155672
R371 drain_right.n29 drain_right.n1 0.155672
R372 drain_right.n67 drain_right.n39 0.155672
R373 drain_right.n60 drain_right.n39 0.155672
R374 drain_right.n60 drain_right.n59 0.155672
R375 drain_right.n59 drain_right.n43 0.155672
R376 drain_right.n52 drain_right.n43 0.155672
R377 drain_right.n52 drain_right.n51 0.155672
R378 drain_right.n34 drain_right.n32 0.0593781
R379 plus.n2 plus.t2 924.929
R380 plus.n8 plus.t7 924.929
R381 plus.n12 plus.t5 924.929
R382 plus.n18 plus.t4 924.929
R383 plus.n1 plus.t0 879.65
R384 plus.n5 plus.t9 879.65
R385 plus.n7 plus.t8 879.65
R386 plus.n11 plus.t6 879.65
R387 plus.n15 plus.t3 879.65
R388 plus.n17 plus.t1 879.65
R389 plus.n3 plus.n2 161.489
R390 plus.n13 plus.n12 161.489
R391 plus.n4 plus.n3 161.3
R392 plus.n6 plus.n0 161.3
R393 plus.n9 plus.n8 161.3
R394 plus.n14 plus.n13 161.3
R395 plus.n16 plus.n10 161.3
R396 plus.n19 plus.n18 161.3
R397 plus.n4 plus.n1 40.8975
R398 plus.n7 plus.n6 40.8975
R399 plus.n17 plus.n16 40.8975
R400 plus.n14 plus.n11 40.8975
R401 plus.n5 plus.n4 36.5157
R402 plus.n6 plus.n5 36.5157
R403 plus.n16 plus.n15 36.5157
R404 plus.n15 plus.n14 36.5157
R405 plus.n2 plus.n1 32.1338
R406 plus.n8 plus.n7 32.1338
R407 plus.n18 plus.n17 32.1338
R408 plus.n12 plus.n11 32.1338
R409 plus plus.n19 25.8002
R410 plus plus.n9 9.82058
R411 plus.n3 plus.n0 0.189894
R412 plus.n9 plus.n0 0.189894
R413 plus.n19 plus.n10 0.189894
R414 plus.n13 plus.n10 0.189894
R415 drain_left.n26 drain_left.n0 289.615
R416 drain_left.n61 drain_left.n35 289.615
R417 drain_left.n11 drain_left.n10 185
R418 drain_left.n8 drain_left.n7 185
R419 drain_left.n17 drain_left.n16 185
R420 drain_left.n19 drain_left.n18 185
R421 drain_left.n4 drain_left.n3 185
R422 drain_left.n25 drain_left.n24 185
R423 drain_left.n27 drain_left.n26 185
R424 drain_left.n62 drain_left.n61 185
R425 drain_left.n60 drain_left.n59 185
R426 drain_left.n39 drain_left.n38 185
R427 drain_left.n54 drain_left.n53 185
R428 drain_left.n52 drain_left.n51 185
R429 drain_left.n43 drain_left.n42 185
R430 drain_left.n46 drain_left.n45 185
R431 drain_left.t5 drain_left.n9 147.661
R432 drain_left.t7 drain_left.n44 147.661
R433 drain_left.n10 drain_left.n7 104.615
R434 drain_left.n17 drain_left.n7 104.615
R435 drain_left.n18 drain_left.n17 104.615
R436 drain_left.n18 drain_left.n3 104.615
R437 drain_left.n25 drain_left.n3 104.615
R438 drain_left.n26 drain_left.n25 104.615
R439 drain_left.n61 drain_left.n60 104.615
R440 drain_left.n60 drain_left.n38 104.615
R441 drain_left.n53 drain_left.n38 104.615
R442 drain_left.n53 drain_left.n52 104.615
R443 drain_left.n52 drain_left.n42 104.615
R444 drain_left.n45 drain_left.n42 104.615
R445 drain_left.n34 drain_left.n33 67.478
R446 drain_left.n67 drain_left.n66 67.1908
R447 drain_left.n69 drain_left.n68 67.1907
R448 drain_left.n32 drain_left.n31 67.1907
R449 drain_left.n10 drain_left.t5 52.3082
R450 drain_left.n45 drain_left.t7 52.3082
R451 drain_left.n32 drain_left.n30 49.321
R452 drain_left.n67 drain_left.n65 49.321
R453 drain_left drain_left.n34 24.7634
R454 drain_left.n11 drain_left.n9 15.6674
R455 drain_left.n46 drain_left.n44 15.6674
R456 drain_left.n12 drain_left.n8 12.8005
R457 drain_left.n47 drain_left.n43 12.8005
R458 drain_left.n16 drain_left.n15 12.0247
R459 drain_left.n51 drain_left.n50 12.0247
R460 drain_left.n19 drain_left.n6 11.249
R461 drain_left.n54 drain_left.n41 11.249
R462 drain_left.n20 drain_left.n4 10.4732
R463 drain_left.n55 drain_left.n39 10.4732
R464 drain_left.n24 drain_left.n23 9.69747
R465 drain_left.n59 drain_left.n58 9.69747
R466 drain_left.n30 drain_left.n29 9.45567
R467 drain_left.n65 drain_left.n64 9.45567
R468 drain_left.n29 drain_left.n28 9.3005
R469 drain_left.n2 drain_left.n1 9.3005
R470 drain_left.n23 drain_left.n22 9.3005
R471 drain_left.n21 drain_left.n20 9.3005
R472 drain_left.n6 drain_left.n5 9.3005
R473 drain_left.n15 drain_left.n14 9.3005
R474 drain_left.n13 drain_left.n12 9.3005
R475 drain_left.n64 drain_left.n63 9.3005
R476 drain_left.n37 drain_left.n36 9.3005
R477 drain_left.n58 drain_left.n57 9.3005
R478 drain_left.n56 drain_left.n55 9.3005
R479 drain_left.n41 drain_left.n40 9.3005
R480 drain_left.n50 drain_left.n49 9.3005
R481 drain_left.n48 drain_left.n47 9.3005
R482 drain_left.n27 drain_left.n2 8.92171
R483 drain_left.n62 drain_left.n37 8.92171
R484 drain_left.n28 drain_left.n0 8.14595
R485 drain_left.n63 drain_left.n35 8.14595
R486 drain_left drain_left.n69 6.11011
R487 drain_left.n30 drain_left.n0 5.81868
R488 drain_left.n65 drain_left.n35 5.81868
R489 drain_left.n28 drain_left.n27 5.04292
R490 drain_left.n63 drain_left.n62 5.04292
R491 drain_left.n13 drain_left.n9 4.38594
R492 drain_left.n48 drain_left.n44 4.38594
R493 drain_left.n24 drain_left.n2 4.26717
R494 drain_left.n59 drain_left.n37 4.26717
R495 drain_left.n23 drain_left.n4 3.49141
R496 drain_left.n58 drain_left.n39 3.49141
R497 drain_left.n33 drain_left.t3 3.3005
R498 drain_left.n33 drain_left.t4 3.3005
R499 drain_left.n31 drain_left.t8 3.3005
R500 drain_left.n31 drain_left.t6 3.3005
R501 drain_left.n68 drain_left.t1 3.3005
R502 drain_left.n68 drain_left.t2 3.3005
R503 drain_left.n66 drain_left.t9 3.3005
R504 drain_left.n66 drain_left.t0 3.3005
R505 drain_left.n20 drain_left.n19 2.71565
R506 drain_left.n55 drain_left.n54 2.71565
R507 drain_left.n16 drain_left.n6 1.93989
R508 drain_left.n51 drain_left.n41 1.93989
R509 drain_left.n15 drain_left.n8 1.16414
R510 drain_left.n50 drain_left.n43 1.16414
R511 drain_left.n69 drain_left.n67 0.457397
R512 drain_left.n12 drain_left.n11 0.388379
R513 drain_left.n47 drain_left.n46 0.388379
R514 drain_left.n14 drain_left.n13 0.155672
R515 drain_left.n14 drain_left.n5 0.155672
R516 drain_left.n21 drain_left.n5 0.155672
R517 drain_left.n22 drain_left.n21 0.155672
R518 drain_left.n22 drain_left.n1 0.155672
R519 drain_left.n29 drain_left.n1 0.155672
R520 drain_left.n64 drain_left.n36 0.155672
R521 drain_left.n57 drain_left.n36 0.155672
R522 drain_left.n57 drain_left.n56 0.155672
R523 drain_left.n56 drain_left.n40 0.155672
R524 drain_left.n49 drain_left.n40 0.155672
R525 drain_left.n49 drain_left.n48 0.155672
R526 drain_left.n34 drain_left.n32 0.0593781
C0 minus plus 3.72944f
C1 source drain_left 13.5005f
C2 source minus 1.57086f
C3 plus drain_right 0.282549f
C4 drain_left minus 0.170748f
C5 source drain_right 13.4933f
C6 drain_left drain_right 0.660358f
C7 minus drain_right 1.72961f
C8 source plus 1.58522f
C9 drain_left plus 1.85605f
C10 drain_right a_n1352_n2088# 4.869051f
C11 drain_left a_n1352_n2088# 5.06191f
C12 source a_n1352_n2088# 3.804386f
C13 minus a_n1352_n2088# 4.737616f
C14 plus a_n1352_n2088# 5.508046f
C15 drain_left.n0 a_n1352_n2088# 0.040261f
C16 drain_left.n1 a_n1352_n2088# 0.028644f
C17 drain_left.n2 a_n1352_n2088# 0.015392f
C18 drain_left.n3 a_n1352_n2088# 0.036381f
C19 drain_left.n4 a_n1352_n2088# 0.016297f
C20 drain_left.n5 a_n1352_n2088# 0.028644f
C21 drain_left.n6 a_n1352_n2088# 0.015392f
C22 drain_left.n7 a_n1352_n2088# 0.036381f
C23 drain_left.n8 a_n1352_n2088# 0.016297f
C24 drain_left.n9 a_n1352_n2088# 0.122575f
C25 drain_left.t5 a_n1352_n2088# 0.059296f
C26 drain_left.n10 a_n1352_n2088# 0.027286f
C27 drain_left.n11 a_n1352_n2088# 0.02149f
C28 drain_left.n12 a_n1352_n2088# 0.015392f
C29 drain_left.n13 a_n1352_n2088# 0.68155f
C30 drain_left.n14 a_n1352_n2088# 0.028644f
C31 drain_left.n15 a_n1352_n2088# 0.015392f
C32 drain_left.n16 a_n1352_n2088# 0.016297f
C33 drain_left.n17 a_n1352_n2088# 0.036381f
C34 drain_left.n18 a_n1352_n2088# 0.036381f
C35 drain_left.n19 a_n1352_n2088# 0.016297f
C36 drain_left.n20 a_n1352_n2088# 0.015392f
C37 drain_left.n21 a_n1352_n2088# 0.028644f
C38 drain_left.n22 a_n1352_n2088# 0.028644f
C39 drain_left.n23 a_n1352_n2088# 0.015392f
C40 drain_left.n24 a_n1352_n2088# 0.016297f
C41 drain_left.n25 a_n1352_n2088# 0.036381f
C42 drain_left.n26 a_n1352_n2088# 0.078758f
C43 drain_left.n27 a_n1352_n2088# 0.016297f
C44 drain_left.n28 a_n1352_n2088# 0.015392f
C45 drain_left.n29 a_n1352_n2088# 0.066209f
C46 drain_left.n30 a_n1352_n2088# 0.064748f
C47 drain_left.t8 a_n1352_n2088# 0.135811f
C48 drain_left.t6 a_n1352_n2088# 0.135811f
C49 drain_left.n31 a_n1352_n2088# 1.13266f
C50 drain_left.n32 a_n1352_n2088# 0.387789f
C51 drain_left.t3 a_n1352_n2088# 0.135811f
C52 drain_left.t4 a_n1352_n2088# 0.135811f
C53 drain_left.n33 a_n1352_n2088# 1.13401f
C54 drain_left.n34 a_n1352_n2088# 1.18567f
C55 drain_left.n35 a_n1352_n2088# 0.040261f
C56 drain_left.n36 a_n1352_n2088# 0.028644f
C57 drain_left.n37 a_n1352_n2088# 0.015392f
C58 drain_left.n38 a_n1352_n2088# 0.036381f
C59 drain_left.n39 a_n1352_n2088# 0.016297f
C60 drain_left.n40 a_n1352_n2088# 0.028644f
C61 drain_left.n41 a_n1352_n2088# 0.015392f
C62 drain_left.n42 a_n1352_n2088# 0.036381f
C63 drain_left.n43 a_n1352_n2088# 0.016297f
C64 drain_left.n44 a_n1352_n2088# 0.122575f
C65 drain_left.t7 a_n1352_n2088# 0.059296f
C66 drain_left.n45 a_n1352_n2088# 0.027286f
C67 drain_left.n46 a_n1352_n2088# 0.02149f
C68 drain_left.n47 a_n1352_n2088# 0.015392f
C69 drain_left.n48 a_n1352_n2088# 0.68155f
C70 drain_left.n49 a_n1352_n2088# 0.028644f
C71 drain_left.n50 a_n1352_n2088# 0.015392f
C72 drain_left.n51 a_n1352_n2088# 0.016297f
C73 drain_left.n52 a_n1352_n2088# 0.036381f
C74 drain_left.n53 a_n1352_n2088# 0.036381f
C75 drain_left.n54 a_n1352_n2088# 0.016297f
C76 drain_left.n55 a_n1352_n2088# 0.015392f
C77 drain_left.n56 a_n1352_n2088# 0.028644f
C78 drain_left.n57 a_n1352_n2088# 0.028644f
C79 drain_left.n58 a_n1352_n2088# 0.015392f
C80 drain_left.n59 a_n1352_n2088# 0.016297f
C81 drain_left.n60 a_n1352_n2088# 0.036381f
C82 drain_left.n61 a_n1352_n2088# 0.078758f
C83 drain_left.n62 a_n1352_n2088# 0.016297f
C84 drain_left.n63 a_n1352_n2088# 0.015392f
C85 drain_left.n64 a_n1352_n2088# 0.066209f
C86 drain_left.n65 a_n1352_n2088# 0.064748f
C87 drain_left.t9 a_n1352_n2088# 0.135811f
C88 drain_left.t0 a_n1352_n2088# 0.135811f
C89 drain_left.n66 a_n1352_n2088# 1.13267f
C90 drain_left.n67 a_n1352_n2088# 0.413241f
C91 drain_left.t1 a_n1352_n2088# 0.135811f
C92 drain_left.t2 a_n1352_n2088# 0.135811f
C93 drain_left.n68 a_n1352_n2088# 1.13266f
C94 drain_left.n69 a_n1352_n2088# 0.551244f
C95 plus.n0 a_n1352_n2088# 0.030304f
C96 plus.t8 a_n1352_n2088# 0.10361f
C97 plus.t9 a_n1352_n2088# 0.10361f
C98 plus.t0 a_n1352_n2088# 0.10361f
C99 plus.n1 a_n1352_n2088# 0.050673f
C100 plus.t2 a_n1352_n2088# 0.1061f
C101 plus.n2 a_n1352_n2088# 0.059026f
C102 plus.n3 a_n1352_n2088# 0.066544f
C103 plus.n4 a_n1352_n2088# 0.010613f
C104 plus.n5 a_n1352_n2088# 0.050673f
C105 plus.n6 a_n1352_n2088# 0.010613f
C106 plus.n7 a_n1352_n2088# 0.050673f
C107 plus.t7 a_n1352_n2088# 0.1061f
C108 plus.n8 a_n1352_n2088# 0.058983f
C109 plus.n9 a_n1352_n2088# 0.255896f
C110 plus.n10 a_n1352_n2088# 0.030304f
C111 plus.t4 a_n1352_n2088# 0.1061f
C112 plus.t1 a_n1352_n2088# 0.10361f
C113 plus.t3 a_n1352_n2088# 0.10361f
C114 plus.t6 a_n1352_n2088# 0.10361f
C115 plus.n11 a_n1352_n2088# 0.050673f
C116 plus.t5 a_n1352_n2088# 0.1061f
C117 plus.n12 a_n1352_n2088# 0.059026f
C118 plus.n13 a_n1352_n2088# 0.066544f
C119 plus.n14 a_n1352_n2088# 0.010613f
C120 plus.n15 a_n1352_n2088# 0.050673f
C121 plus.n16 a_n1352_n2088# 0.010613f
C122 plus.n17 a_n1352_n2088# 0.050673f
C123 plus.n18 a_n1352_n2088# 0.058983f
C124 plus.n19 a_n1352_n2088# 0.696959f
C125 drain_right.n0 a_n1352_n2088# 0.040598f
C126 drain_right.n1 a_n1352_n2088# 0.028884f
C127 drain_right.n2 a_n1352_n2088# 0.015521f
C128 drain_right.n3 a_n1352_n2088# 0.036685f
C129 drain_right.n4 a_n1352_n2088# 0.016434f
C130 drain_right.n5 a_n1352_n2088# 0.028884f
C131 drain_right.n6 a_n1352_n2088# 0.015521f
C132 drain_right.n7 a_n1352_n2088# 0.036685f
C133 drain_right.n8 a_n1352_n2088# 0.016434f
C134 drain_right.n9 a_n1352_n2088# 0.123601f
C135 drain_right.t3 a_n1352_n2088# 0.059792f
C136 drain_right.n10 a_n1352_n2088# 0.027514f
C137 drain_right.n11 a_n1352_n2088# 0.02167f
C138 drain_right.n12 a_n1352_n2088# 0.015521f
C139 drain_right.n13 a_n1352_n2088# 0.687254f
C140 drain_right.n14 a_n1352_n2088# 0.028884f
C141 drain_right.n15 a_n1352_n2088# 0.015521f
C142 drain_right.n16 a_n1352_n2088# 0.016434f
C143 drain_right.n17 a_n1352_n2088# 0.036685f
C144 drain_right.n18 a_n1352_n2088# 0.036685f
C145 drain_right.n19 a_n1352_n2088# 0.016434f
C146 drain_right.n20 a_n1352_n2088# 0.015521f
C147 drain_right.n21 a_n1352_n2088# 0.028884f
C148 drain_right.n22 a_n1352_n2088# 0.028884f
C149 drain_right.n23 a_n1352_n2088# 0.015521f
C150 drain_right.n24 a_n1352_n2088# 0.016434f
C151 drain_right.n25 a_n1352_n2088# 0.036685f
C152 drain_right.n26 a_n1352_n2088# 0.079418f
C153 drain_right.n27 a_n1352_n2088# 0.016434f
C154 drain_right.n28 a_n1352_n2088# 0.015521f
C155 drain_right.n29 a_n1352_n2088# 0.066763f
C156 drain_right.n30 a_n1352_n2088# 0.06529f
C157 drain_right.t0 a_n1352_n2088# 0.136948f
C158 drain_right.t4 a_n1352_n2088# 0.136948f
C159 drain_right.n31 a_n1352_n2088# 1.14214f
C160 drain_right.n32 a_n1352_n2088# 0.391035f
C161 drain_right.t1 a_n1352_n2088# 0.136948f
C162 drain_right.t8 a_n1352_n2088# 0.136948f
C163 drain_right.n33 a_n1352_n2088# 1.1435f
C164 drain_right.n34 a_n1352_n2088# 1.13647f
C165 drain_right.t7 a_n1352_n2088# 0.136948f
C166 drain_right.t6 a_n1352_n2088# 0.136948f
C167 drain_right.n35 a_n1352_n2088# 1.14438f
C168 drain_right.t2 a_n1352_n2088# 0.136948f
C169 drain_right.t9 a_n1352_n2088# 0.136948f
C170 drain_right.n36 a_n1352_n2088# 1.14215f
C171 drain_right.n37 a_n1352_n2088# 0.64834f
C172 drain_right.n38 a_n1352_n2088# 0.040598f
C173 drain_right.n39 a_n1352_n2088# 0.028884f
C174 drain_right.n40 a_n1352_n2088# 0.015521f
C175 drain_right.n41 a_n1352_n2088# 0.036685f
C176 drain_right.n42 a_n1352_n2088# 0.016434f
C177 drain_right.n43 a_n1352_n2088# 0.028884f
C178 drain_right.n44 a_n1352_n2088# 0.015521f
C179 drain_right.n45 a_n1352_n2088# 0.036685f
C180 drain_right.n46 a_n1352_n2088# 0.016434f
C181 drain_right.n47 a_n1352_n2088# 0.123601f
C182 drain_right.t5 a_n1352_n2088# 0.059792f
C183 drain_right.n48 a_n1352_n2088# 0.027514f
C184 drain_right.n49 a_n1352_n2088# 0.02167f
C185 drain_right.n50 a_n1352_n2088# 0.015521f
C186 drain_right.n51 a_n1352_n2088# 0.687254f
C187 drain_right.n52 a_n1352_n2088# 0.028884f
C188 drain_right.n53 a_n1352_n2088# 0.015521f
C189 drain_right.n54 a_n1352_n2088# 0.016434f
C190 drain_right.n55 a_n1352_n2088# 0.036685f
C191 drain_right.n56 a_n1352_n2088# 0.036685f
C192 drain_right.n57 a_n1352_n2088# 0.016434f
C193 drain_right.n58 a_n1352_n2088# 0.015521f
C194 drain_right.n59 a_n1352_n2088# 0.028884f
C195 drain_right.n60 a_n1352_n2088# 0.028884f
C196 drain_right.n61 a_n1352_n2088# 0.015521f
C197 drain_right.n62 a_n1352_n2088# 0.016434f
C198 drain_right.n63 a_n1352_n2088# 0.036685f
C199 drain_right.n64 a_n1352_n2088# 0.079418f
C200 drain_right.n65 a_n1352_n2088# 0.016434f
C201 drain_right.n66 a_n1352_n2088# 0.015521f
C202 drain_right.n67 a_n1352_n2088# 0.066763f
C203 drain_right.n68 a_n1352_n2088# 0.06438f
C204 drain_right.n69 a_n1352_n2088# 0.332898f
C205 source.n0 a_n1352_n2088# 0.044235f
C206 source.n1 a_n1352_n2088# 0.031471f
C207 source.n2 a_n1352_n2088# 0.016911f
C208 source.n3 a_n1352_n2088# 0.039971f
C209 source.n4 a_n1352_n2088# 0.017906f
C210 source.n5 a_n1352_n2088# 0.031471f
C211 source.n6 a_n1352_n2088# 0.016911f
C212 source.n7 a_n1352_n2088# 0.039971f
C213 source.n8 a_n1352_n2088# 0.017906f
C214 source.n9 a_n1352_n2088# 0.134672f
C215 source.t0 a_n1352_n2088# 0.065148f
C216 source.n10 a_n1352_n2088# 0.029979f
C217 source.n11 a_n1352_n2088# 0.023611f
C218 source.n12 a_n1352_n2088# 0.016911f
C219 source.n13 a_n1352_n2088# 0.748815f
C220 source.n14 a_n1352_n2088# 0.031471f
C221 source.n15 a_n1352_n2088# 0.016911f
C222 source.n16 a_n1352_n2088# 0.017906f
C223 source.n17 a_n1352_n2088# 0.039971f
C224 source.n18 a_n1352_n2088# 0.039971f
C225 source.n19 a_n1352_n2088# 0.017906f
C226 source.n20 a_n1352_n2088# 0.016911f
C227 source.n21 a_n1352_n2088# 0.031471f
C228 source.n22 a_n1352_n2088# 0.031471f
C229 source.n23 a_n1352_n2088# 0.016911f
C230 source.n24 a_n1352_n2088# 0.017906f
C231 source.n25 a_n1352_n2088# 0.039971f
C232 source.n26 a_n1352_n2088# 0.086531f
C233 source.n27 a_n1352_n2088# 0.017906f
C234 source.n28 a_n1352_n2088# 0.016911f
C235 source.n29 a_n1352_n2088# 0.072743f
C236 source.n30 a_n1352_n2088# 0.048418f
C237 source.n31 a_n1352_n2088# 0.747288f
C238 source.t7 a_n1352_n2088# 0.149215f
C239 source.t8 a_n1352_n2088# 0.149215f
C240 source.n32 a_n1352_n2088# 1.1621f
C241 source.n33 a_n1352_n2088# 0.387671f
C242 source.t1 a_n1352_n2088# 0.149215f
C243 source.t9 a_n1352_n2088# 0.149215f
C244 source.n34 a_n1352_n2088# 1.1621f
C245 source.n35 a_n1352_n2088# 0.412149f
C246 source.n36 a_n1352_n2088# 0.044235f
C247 source.n37 a_n1352_n2088# 0.031471f
C248 source.n38 a_n1352_n2088# 0.016911f
C249 source.n39 a_n1352_n2088# 0.039971f
C250 source.n40 a_n1352_n2088# 0.017906f
C251 source.n41 a_n1352_n2088# 0.031471f
C252 source.n42 a_n1352_n2088# 0.016911f
C253 source.n43 a_n1352_n2088# 0.039971f
C254 source.n44 a_n1352_n2088# 0.017906f
C255 source.n45 a_n1352_n2088# 0.134672f
C256 source.t18 a_n1352_n2088# 0.065148f
C257 source.n46 a_n1352_n2088# 0.029979f
C258 source.n47 a_n1352_n2088# 0.023611f
C259 source.n48 a_n1352_n2088# 0.016911f
C260 source.n49 a_n1352_n2088# 0.748815f
C261 source.n50 a_n1352_n2088# 0.031471f
C262 source.n51 a_n1352_n2088# 0.016911f
C263 source.n52 a_n1352_n2088# 0.017906f
C264 source.n53 a_n1352_n2088# 0.039971f
C265 source.n54 a_n1352_n2088# 0.039971f
C266 source.n55 a_n1352_n2088# 0.017906f
C267 source.n56 a_n1352_n2088# 0.016911f
C268 source.n57 a_n1352_n2088# 0.031471f
C269 source.n58 a_n1352_n2088# 0.031471f
C270 source.n59 a_n1352_n2088# 0.016911f
C271 source.n60 a_n1352_n2088# 0.017906f
C272 source.n61 a_n1352_n2088# 0.039971f
C273 source.n62 a_n1352_n2088# 0.086531f
C274 source.n63 a_n1352_n2088# 0.017906f
C275 source.n64 a_n1352_n2088# 0.016911f
C276 source.n65 a_n1352_n2088# 0.072743f
C277 source.n66 a_n1352_n2088# 0.048418f
C278 source.n67 a_n1352_n2088# 0.144019f
C279 source.t14 a_n1352_n2088# 0.149215f
C280 source.t10 a_n1352_n2088# 0.149215f
C281 source.n68 a_n1352_n2088# 1.1621f
C282 source.n69 a_n1352_n2088# 0.387671f
C283 source.t11 a_n1352_n2088# 0.149215f
C284 source.t13 a_n1352_n2088# 0.149215f
C285 source.n70 a_n1352_n2088# 1.1621f
C286 source.n71 a_n1352_n2088# 1.46441f
C287 source.t4 a_n1352_n2088# 0.149215f
C288 source.t2 a_n1352_n2088# 0.149215f
C289 source.n72 a_n1352_n2088# 1.16209f
C290 source.n73 a_n1352_n2088# 1.46442f
C291 source.t3 a_n1352_n2088# 0.149215f
C292 source.t6 a_n1352_n2088# 0.149215f
C293 source.n74 a_n1352_n2088# 1.16209f
C294 source.n75 a_n1352_n2088# 0.387679f
C295 source.n76 a_n1352_n2088# 0.044235f
C296 source.n77 a_n1352_n2088# 0.031471f
C297 source.n78 a_n1352_n2088# 0.016911f
C298 source.n79 a_n1352_n2088# 0.039971f
C299 source.n80 a_n1352_n2088# 0.017906f
C300 source.n81 a_n1352_n2088# 0.031471f
C301 source.n82 a_n1352_n2088# 0.016911f
C302 source.n83 a_n1352_n2088# 0.039971f
C303 source.n84 a_n1352_n2088# 0.017906f
C304 source.n85 a_n1352_n2088# 0.134672f
C305 source.t5 a_n1352_n2088# 0.065148f
C306 source.n86 a_n1352_n2088# 0.029979f
C307 source.n87 a_n1352_n2088# 0.023611f
C308 source.n88 a_n1352_n2088# 0.016911f
C309 source.n89 a_n1352_n2088# 0.748815f
C310 source.n90 a_n1352_n2088# 0.031471f
C311 source.n91 a_n1352_n2088# 0.016911f
C312 source.n92 a_n1352_n2088# 0.017906f
C313 source.n93 a_n1352_n2088# 0.039971f
C314 source.n94 a_n1352_n2088# 0.039971f
C315 source.n95 a_n1352_n2088# 0.017906f
C316 source.n96 a_n1352_n2088# 0.016911f
C317 source.n97 a_n1352_n2088# 0.031471f
C318 source.n98 a_n1352_n2088# 0.031471f
C319 source.n99 a_n1352_n2088# 0.016911f
C320 source.n100 a_n1352_n2088# 0.017906f
C321 source.n101 a_n1352_n2088# 0.039971f
C322 source.n102 a_n1352_n2088# 0.086531f
C323 source.n103 a_n1352_n2088# 0.017906f
C324 source.n104 a_n1352_n2088# 0.016911f
C325 source.n105 a_n1352_n2088# 0.072743f
C326 source.n106 a_n1352_n2088# 0.048418f
C327 source.n107 a_n1352_n2088# 0.144019f
C328 source.t12 a_n1352_n2088# 0.149215f
C329 source.t19 a_n1352_n2088# 0.149215f
C330 source.n108 a_n1352_n2088# 1.16209f
C331 source.n109 a_n1352_n2088# 0.412157f
C332 source.t17 a_n1352_n2088# 0.149215f
C333 source.t16 a_n1352_n2088# 0.149215f
C334 source.n110 a_n1352_n2088# 1.16209f
C335 source.n111 a_n1352_n2088# 0.387679f
C336 source.n112 a_n1352_n2088# 0.044235f
C337 source.n113 a_n1352_n2088# 0.031471f
C338 source.n114 a_n1352_n2088# 0.016911f
C339 source.n115 a_n1352_n2088# 0.039971f
C340 source.n116 a_n1352_n2088# 0.017906f
C341 source.n117 a_n1352_n2088# 0.031471f
C342 source.n118 a_n1352_n2088# 0.016911f
C343 source.n119 a_n1352_n2088# 0.039971f
C344 source.n120 a_n1352_n2088# 0.017906f
C345 source.n121 a_n1352_n2088# 0.134672f
C346 source.t15 a_n1352_n2088# 0.065148f
C347 source.n122 a_n1352_n2088# 0.029979f
C348 source.n123 a_n1352_n2088# 0.023611f
C349 source.n124 a_n1352_n2088# 0.016911f
C350 source.n125 a_n1352_n2088# 0.748815f
C351 source.n126 a_n1352_n2088# 0.031471f
C352 source.n127 a_n1352_n2088# 0.016911f
C353 source.n128 a_n1352_n2088# 0.017906f
C354 source.n129 a_n1352_n2088# 0.039971f
C355 source.n130 a_n1352_n2088# 0.039971f
C356 source.n131 a_n1352_n2088# 0.017906f
C357 source.n132 a_n1352_n2088# 0.016911f
C358 source.n133 a_n1352_n2088# 0.031471f
C359 source.n134 a_n1352_n2088# 0.031471f
C360 source.n135 a_n1352_n2088# 0.016911f
C361 source.n136 a_n1352_n2088# 0.017906f
C362 source.n137 a_n1352_n2088# 0.039971f
C363 source.n138 a_n1352_n2088# 0.086531f
C364 source.n139 a_n1352_n2088# 0.017906f
C365 source.n140 a_n1352_n2088# 0.016911f
C366 source.n141 a_n1352_n2088# 0.072743f
C367 source.n142 a_n1352_n2088# 0.048418f
C368 source.n143 a_n1352_n2088# 0.291497f
C369 source.n144 a_n1352_n2088# 1.2835f
C370 minus.n0 a_n1352_n2088# 0.02981f
C371 minus.t4 a_n1352_n2088# 0.104371f
C372 minus.t7 a_n1352_n2088# 0.101922f
C373 minus.t0 a_n1352_n2088# 0.101922f
C374 minus.t2 a_n1352_n2088# 0.101922f
C375 minus.n1 a_n1352_n2088# 0.049847f
C376 minus.t3 a_n1352_n2088# 0.104371f
C377 minus.n2 a_n1352_n2088# 0.058064f
C378 minus.n3 a_n1352_n2088# 0.06546f
C379 minus.n4 a_n1352_n2088# 0.01044f
C380 minus.n5 a_n1352_n2088# 0.049847f
C381 minus.n6 a_n1352_n2088# 0.01044f
C382 minus.n7 a_n1352_n2088# 0.049847f
C383 minus.n8 a_n1352_n2088# 0.058022f
C384 minus.n9 a_n1352_n2088# 0.758477f
C385 minus.n10 a_n1352_n2088# 0.02981f
C386 minus.t8 a_n1352_n2088# 0.101922f
C387 minus.t5 a_n1352_n2088# 0.101922f
C388 minus.t9 a_n1352_n2088# 0.101922f
C389 minus.n11 a_n1352_n2088# 0.049847f
C390 minus.t6 a_n1352_n2088# 0.104371f
C391 minus.n12 a_n1352_n2088# 0.058064f
C392 minus.n13 a_n1352_n2088# 0.06546f
C393 minus.n14 a_n1352_n2088# 0.01044f
C394 minus.n15 a_n1352_n2088# 0.049847f
C395 minus.n16 a_n1352_n2088# 0.01044f
C396 minus.n17 a_n1352_n2088# 0.049847f
C397 minus.t1 a_n1352_n2088# 0.104371f
C398 minus.n18 a_n1352_n2088# 0.058022f
C399 minus.n19 a_n1352_n2088# 0.191327f
C400 minus.n20 a_n1352_n2088# 0.938052f
.ends

