* NGSPICE file created from diffpair398.ext - technology: sky130A

.subckt diffpair398 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t31 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X1 a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X2 a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X3 drain_right.t18 minus.t1 source.t32 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 source.t15 plus.t0 drain_left.t19 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X5 drain_left.t18 plus.t1 source.t2 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X7 source.t9 plus.t2 drain_left.t17 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 drain_right.t17 minus.t2 source.t33 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X9 drain_left.t16 plus.t3 source.t11 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X11 source.t34 minus.t3 drain_right.t16 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X12 drain_right.t15 minus.t4 source.t35 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X13 drain_left.t15 plus.t4 source.t10 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X14 drain_left.t14 plus.t5 source.t8 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X15 drain_left.t13 plus.t6 source.t4 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X16 source.t36 minus.t5 drain_right.t14 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X17 source.t20 minus.t6 drain_right.t13 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X18 drain_right.t12 minus.t7 source.t25 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 source.t27 minus.t8 drain_right.t11 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X20 drain_right.t10 minus.t9 source.t21 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X21 source.t29 minus.t10 drain_right.t9 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X22 source.t3 plus.t7 drain_left.t12 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X23 source.t28 minus.t11 drain_right.t8 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X24 source.t39 plus.t8 drain_left.t11 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X25 drain_left.t10 plus.t9 source.t12 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X26 source.t37 minus.t12 drain_right.t7 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X27 drain_right.t6 minus.t13 source.t19 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X28 drain_left.t9 plus.t10 source.t5 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X29 drain_right.t5 minus.t14 source.t22 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X30 source.t17 plus.t11 drain_left.t8 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X31 source.t24 minus.t15 drain_right.t4 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X32 drain_left.t7 plus.t12 source.t18 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X33 drain_left.t6 plus.t13 source.t13 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X34 source.t30 minus.t16 drain_right.t3 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X35 source.t38 minus.t17 drain_right.t2 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X36 source.t16 plus.t14 drain_left.t5 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X37 source.t1 plus.t15 drain_left.t4 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X38 drain_right.t1 minus.t18 source.t26 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X39 source.t0 plus.t16 drain_left.t3 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X40 drain_left.t2 plus.t17 source.t14 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X41 drain_right.t0 minus.t19 source.t23 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X42 source.t7 plus.t18 drain_left.t1 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X43 source.t6 plus.t19 drain_left.t0 a_n3202_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n7 minus.t9 342.019
R1 minus.n37 minus.t17 342.019
R2 minus.n8 minus.t5 320.229
R3 minus.n10 minus.t4 320.229
R4 minus.n5 minus.t12 320.229
R5 minus.n15 minus.t14 320.229
R6 minus.n3 minus.t11 320.229
R7 minus.n21 minus.t7 320.229
R8 minus.n22 minus.t16 320.229
R9 minus.n26 minus.t13 320.229
R10 minus.n28 minus.t3 320.229
R11 minus.n38 minus.t2 320.229
R12 minus.n40 minus.t8 320.229
R13 minus.n35 minus.t1 320.229
R14 minus.n45 minus.t15 320.229
R15 minus.n33 minus.t0 320.229
R16 minus.n51 minus.t6 320.229
R17 minus.n52 minus.t18 320.229
R18 minus.n56 minus.t10 320.229
R19 minus.n58 minus.t19 320.229
R20 minus.n29 minus.n28 161.3
R21 minus.n27 minus.n0 161.3
R22 minus.n26 minus.n25 161.3
R23 minus.n24 minus.n1 161.3
R24 minus.n20 minus.n19 161.3
R25 minus.n18 minus.n3 161.3
R26 minus.n17 minus.n16 161.3
R27 minus.n15 minus.n4 161.3
R28 minus.n14 minus.n13 161.3
R29 minus.n9 minus.n6 161.3
R30 minus.n59 minus.n58 161.3
R31 minus.n57 minus.n30 161.3
R32 minus.n56 minus.n55 161.3
R33 minus.n54 minus.n31 161.3
R34 minus.n50 minus.n49 161.3
R35 minus.n48 minus.n33 161.3
R36 minus.n47 minus.n46 161.3
R37 minus.n45 minus.n34 161.3
R38 minus.n44 minus.n43 161.3
R39 minus.n39 minus.n36 161.3
R40 minus.n23 minus.n22 80.6037
R41 minus.n21 minus.n2 80.6037
R42 minus.n12 minus.n5 80.6037
R43 minus.n11 minus.n10 80.6037
R44 minus.n53 minus.n52 80.6037
R45 minus.n51 minus.n32 80.6037
R46 minus.n42 minus.n35 80.6037
R47 minus.n41 minus.n40 80.6037
R48 minus.n10 minus.n5 48.2005
R49 minus.n22 minus.n21 48.2005
R50 minus.n40 minus.n35 48.2005
R51 minus.n52 minus.n51 48.2005
R52 minus.n7 minus.n6 44.8565
R53 minus.n37 minus.n36 44.8565
R54 minus.n14 minus.n5 43.0884
R55 minus.n21 minus.n20 43.0884
R56 minus.n44 minus.n35 43.0884
R57 minus.n51 minus.n50 43.0884
R58 minus.n10 minus.n9 40.1672
R59 minus.n22 minus.n1 40.1672
R60 minus.n40 minus.n39 40.1672
R61 minus.n52 minus.n31 40.1672
R62 minus.n60 minus.n29 39.1823
R63 minus.n28 minus.n27 27.0217
R64 minus.n58 minus.n57 27.0217
R65 minus.n16 minus.n3 24.1005
R66 minus.n16 minus.n15 24.1005
R67 minus.n46 minus.n45 24.1005
R68 minus.n46 minus.n33 24.1005
R69 minus.n27 minus.n26 21.1793
R70 minus.n57 minus.n56 21.1793
R71 minus.n8 minus.n7 20.1275
R72 minus.n38 minus.n37 20.1275
R73 minus.n9 minus.n8 8.03383
R74 minus.n26 minus.n1 8.03383
R75 minus.n39 minus.n38 8.03383
R76 minus.n56 minus.n31 8.03383
R77 minus.n60 minus.n59 6.70505
R78 minus.n15 minus.n14 5.11262
R79 minus.n20 minus.n3 5.11262
R80 minus.n45 minus.n44 5.11262
R81 minus.n50 minus.n33 5.11262
R82 minus.n23 minus.n2 0.380177
R83 minus.n12 minus.n11 0.380177
R84 minus.n42 minus.n41 0.380177
R85 minus.n53 minus.n32 0.380177
R86 minus.n24 minus.n23 0.285035
R87 minus.n19 minus.n2 0.285035
R88 minus.n13 minus.n12 0.285035
R89 minus.n11 minus.n6 0.285035
R90 minus.n41 minus.n36 0.285035
R91 minus.n43 minus.n42 0.285035
R92 minus.n49 minus.n32 0.285035
R93 minus.n54 minus.n53 0.285035
R94 minus.n29 minus.n0 0.189894
R95 minus.n25 minus.n0 0.189894
R96 minus.n25 minus.n24 0.189894
R97 minus.n19 minus.n18 0.189894
R98 minus.n18 minus.n17 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n13 minus.n4 0.189894
R101 minus.n43 minus.n34 0.189894
R102 minus.n47 minus.n34 0.189894
R103 minus.n48 minus.n47 0.189894
R104 minus.n49 minus.n48 0.189894
R105 minus.n55 minus.n54 0.189894
R106 minus.n55 minus.n30 0.189894
R107 minus.n59 minus.n30 0.189894
R108 minus minus.n60 0.188
R109 source.n9 source.t7 51.0588
R110 source.n10 source.t21 51.0588
R111 source.n19 source.t34 51.0588
R112 source.n39 source.t23 51.0586
R113 source.n30 source.t38 51.0586
R114 source.n29 source.t5 51.0586
R115 source.n20 source.t39 51.0586
R116 source.n0 source.t4 51.0586
R117 source.n2 source.n1 48.8588
R118 source.n4 source.n3 48.8588
R119 source.n6 source.n5 48.8588
R120 source.n8 source.n7 48.8588
R121 source.n12 source.n11 48.8588
R122 source.n14 source.n13 48.8588
R123 source.n16 source.n15 48.8588
R124 source.n18 source.n17 48.8588
R125 source.n38 source.n37 48.8586
R126 source.n36 source.n35 48.8586
R127 source.n34 source.n33 48.8586
R128 source.n32 source.n31 48.8586
R129 source.n28 source.n27 48.8586
R130 source.n26 source.n25 48.8586
R131 source.n24 source.n23 48.8586
R132 source.n22 source.n21 48.8586
R133 source.n20 source.n19 19.9891
R134 source.n40 source.n0 14.2391
R135 source.n40 source.n39 5.7505
R136 source.n37 source.t26 2.2005
R137 source.n37 source.t29 2.2005
R138 source.n35 source.t31 2.2005
R139 source.n35 source.t20 2.2005
R140 source.n33 source.t32 2.2005
R141 source.n33 source.t24 2.2005
R142 source.n31 source.t33 2.2005
R143 source.n31 source.t27 2.2005
R144 source.n27 source.t8 2.2005
R145 source.n27 source.t9 2.2005
R146 source.n25 source.t10 2.2005
R147 source.n25 source.t15 2.2005
R148 source.n23 source.t11 2.2005
R149 source.n23 source.t16 2.2005
R150 source.n21 source.t2 2.2005
R151 source.n21 source.t6 2.2005
R152 source.n1 source.t12 2.2005
R153 source.n1 source.t3 2.2005
R154 source.n3 source.t18 2.2005
R155 source.n3 source.t17 2.2005
R156 source.n5 source.t13 2.2005
R157 source.n5 source.t0 2.2005
R158 source.n7 source.t14 2.2005
R159 source.n7 source.t1 2.2005
R160 source.n11 source.t35 2.2005
R161 source.n11 source.t36 2.2005
R162 source.n13 source.t22 2.2005
R163 source.n13 source.t37 2.2005
R164 source.n15 source.t25 2.2005
R165 source.n15 source.t28 2.2005
R166 source.n17 source.t19 2.2005
R167 source.n17 source.t30 2.2005
R168 source.n19 source.n18 0.974638
R169 source.n18 source.n16 0.974638
R170 source.n16 source.n14 0.974638
R171 source.n14 source.n12 0.974638
R172 source.n12 source.n10 0.974638
R173 source.n9 source.n8 0.974638
R174 source.n8 source.n6 0.974638
R175 source.n6 source.n4 0.974638
R176 source.n4 source.n2 0.974638
R177 source.n2 source.n0 0.974638
R178 source.n22 source.n20 0.974638
R179 source.n24 source.n22 0.974638
R180 source.n26 source.n24 0.974638
R181 source.n28 source.n26 0.974638
R182 source.n29 source.n28 0.974638
R183 source.n32 source.n30 0.974638
R184 source.n34 source.n32 0.974638
R185 source.n36 source.n34 0.974638
R186 source.n38 source.n36 0.974638
R187 source.n39 source.n38 0.974638
R188 source.n10 source.n9 0.470328
R189 source.n30 source.n29 0.470328
R190 source source.n40 0.188
R191 drain_right.n10 drain_right.n8 66.5116
R192 drain_right.n6 drain_right.n4 66.5115
R193 drain_right.n2 drain_right.n0 66.5115
R194 drain_right.n10 drain_right.n9 65.5376
R195 drain_right.n12 drain_right.n11 65.5376
R196 drain_right.n14 drain_right.n13 65.5376
R197 drain_right.n16 drain_right.n15 65.5376
R198 drain_right.n7 drain_right.n3 65.5373
R199 drain_right.n6 drain_right.n5 65.5373
R200 drain_right.n2 drain_right.n1 65.5373
R201 drain_right drain_right.n7 32.3342
R202 drain_right drain_right.n16 6.62735
R203 drain_right.n3 drain_right.t4 2.2005
R204 drain_right.n3 drain_right.t19 2.2005
R205 drain_right.n4 drain_right.t9 2.2005
R206 drain_right.n4 drain_right.t0 2.2005
R207 drain_right.n5 drain_right.t13 2.2005
R208 drain_right.n5 drain_right.t1 2.2005
R209 drain_right.n1 drain_right.t11 2.2005
R210 drain_right.n1 drain_right.t18 2.2005
R211 drain_right.n0 drain_right.t2 2.2005
R212 drain_right.n0 drain_right.t17 2.2005
R213 drain_right.n8 drain_right.t14 2.2005
R214 drain_right.n8 drain_right.t10 2.2005
R215 drain_right.n9 drain_right.t7 2.2005
R216 drain_right.n9 drain_right.t15 2.2005
R217 drain_right.n11 drain_right.t8 2.2005
R218 drain_right.n11 drain_right.t5 2.2005
R219 drain_right.n13 drain_right.t3 2.2005
R220 drain_right.n13 drain_right.t12 2.2005
R221 drain_right.n15 drain_right.t16 2.2005
R222 drain_right.n15 drain_right.t6 2.2005
R223 drain_right.n16 drain_right.n14 0.974638
R224 drain_right.n14 drain_right.n12 0.974638
R225 drain_right.n12 drain_right.n10 0.974638
R226 drain_right.n7 drain_right.n6 0.919292
R227 drain_right.n7 drain_right.n2 0.919292
R228 plus.n9 plus.t18 342.019
R229 plus.n39 plus.t10 342.019
R230 plus.n28 plus.t6 320.229
R231 plus.n26 plus.t7 320.229
R232 plus.n2 plus.t9 320.229
R233 plus.n21 plus.t11 320.229
R234 plus.n19 plus.t12 320.229
R235 plus.n5 plus.t16 320.229
R236 plus.n13 plus.t13 320.229
R237 plus.n12 plus.t15 320.229
R238 plus.n8 plus.t17 320.229
R239 plus.n58 plus.t8 320.229
R240 plus.n56 plus.t1 320.229
R241 plus.n32 plus.t19 320.229
R242 plus.n51 plus.t3 320.229
R243 plus.n49 plus.t14 320.229
R244 plus.n35 plus.t4 320.229
R245 plus.n43 plus.t0 320.229
R246 plus.n42 plus.t5 320.229
R247 plus.n38 plus.t2 320.229
R248 plus.n11 plus.n10 161.3
R249 plus.n15 plus.n14 161.3
R250 plus.n16 plus.n5 161.3
R251 plus.n18 plus.n17 161.3
R252 plus.n19 plus.n4 161.3
R253 plus.n20 plus.n3 161.3
R254 plus.n25 plus.n24 161.3
R255 plus.n26 plus.n1 161.3
R256 plus.n27 plus.n0 161.3
R257 plus.n29 plus.n28 161.3
R258 plus.n41 plus.n40 161.3
R259 plus.n45 plus.n44 161.3
R260 plus.n46 plus.n35 161.3
R261 plus.n48 plus.n47 161.3
R262 plus.n49 plus.n34 161.3
R263 plus.n50 plus.n33 161.3
R264 plus.n55 plus.n54 161.3
R265 plus.n56 plus.n31 161.3
R266 plus.n57 plus.n30 161.3
R267 plus.n59 plus.n58 161.3
R268 plus.n12 plus.n7 80.6037
R269 plus.n13 plus.n6 80.6037
R270 plus.n22 plus.n21 80.6037
R271 plus.n23 plus.n2 80.6037
R272 plus.n42 plus.n37 80.6037
R273 plus.n43 plus.n36 80.6037
R274 plus.n52 plus.n51 80.6037
R275 plus.n53 plus.n32 80.6037
R276 plus.n21 plus.n2 48.2005
R277 plus.n13 plus.n12 48.2005
R278 plus.n51 plus.n32 48.2005
R279 plus.n43 plus.n42 48.2005
R280 plus.n40 plus.n39 44.8565
R281 plus.n10 plus.n9 44.8565
R282 plus.n21 plus.n20 43.0884
R283 plus.n14 plus.n13 43.0884
R284 plus.n51 plus.n50 43.0884
R285 plus.n44 plus.n43 43.0884
R286 plus.n25 plus.n2 40.1672
R287 plus.n12 plus.n11 40.1672
R288 plus.n55 plus.n32 40.1672
R289 plus.n42 plus.n41 40.1672
R290 plus plus.n59 34.1998
R291 plus.n28 plus.n27 27.0217
R292 plus.n58 plus.n57 27.0217
R293 plus.n18 plus.n5 24.1005
R294 plus.n19 plus.n18 24.1005
R295 plus.n49 plus.n48 24.1005
R296 plus.n48 plus.n35 24.1005
R297 plus.n27 plus.n26 21.1793
R298 plus.n57 plus.n56 21.1793
R299 plus.n39 plus.n38 20.1275
R300 plus.n9 plus.n8 20.1275
R301 plus plus.n29 11.2126
R302 plus.n26 plus.n25 8.03383
R303 plus.n11 plus.n8 8.03383
R304 plus.n56 plus.n55 8.03383
R305 plus.n41 plus.n38 8.03383
R306 plus.n20 plus.n19 5.11262
R307 plus.n14 plus.n5 5.11262
R308 plus.n50 plus.n49 5.11262
R309 plus.n44 plus.n35 5.11262
R310 plus.n7 plus.n6 0.380177
R311 plus.n23 plus.n22 0.380177
R312 plus.n53 plus.n52 0.380177
R313 plus.n37 plus.n36 0.380177
R314 plus.n10 plus.n7 0.285035
R315 plus.n15 plus.n6 0.285035
R316 plus.n22 plus.n3 0.285035
R317 plus.n24 plus.n23 0.285035
R318 plus.n54 plus.n53 0.285035
R319 plus.n52 plus.n33 0.285035
R320 plus.n45 plus.n36 0.285035
R321 plus.n40 plus.n37 0.285035
R322 plus.n16 plus.n15 0.189894
R323 plus.n17 plus.n16 0.189894
R324 plus.n17 plus.n4 0.189894
R325 plus.n4 plus.n3 0.189894
R326 plus.n24 plus.n1 0.189894
R327 plus.n1 plus.n0 0.189894
R328 plus.n29 plus.n0 0.189894
R329 plus.n59 plus.n30 0.189894
R330 plus.n31 plus.n30 0.189894
R331 plus.n54 plus.n31 0.189894
R332 plus.n34 plus.n33 0.189894
R333 plus.n47 plus.n34 0.189894
R334 plus.n47 plus.n46 0.189894
R335 plus.n46 plus.n45 0.189894
R336 drain_left.n10 drain_left.n8 66.5117
R337 drain_left.n6 drain_left.n4 66.5115
R338 drain_left.n2 drain_left.n0 66.5115
R339 drain_left.n14 drain_left.n13 65.5376
R340 drain_left.n12 drain_left.n11 65.5376
R341 drain_left.n10 drain_left.n9 65.5376
R342 drain_left.n16 drain_left.n15 65.5374
R343 drain_left.n7 drain_left.n3 65.5373
R344 drain_left.n6 drain_left.n5 65.5373
R345 drain_left.n2 drain_left.n1 65.5373
R346 drain_left drain_left.n7 32.8875
R347 drain_left drain_left.n16 6.62735
R348 drain_left.n3 drain_left.t5 2.2005
R349 drain_left.n3 drain_left.t15 2.2005
R350 drain_left.n4 drain_left.t17 2.2005
R351 drain_left.n4 drain_left.t9 2.2005
R352 drain_left.n5 drain_left.t19 2.2005
R353 drain_left.n5 drain_left.t14 2.2005
R354 drain_left.n1 drain_left.t0 2.2005
R355 drain_left.n1 drain_left.t16 2.2005
R356 drain_left.n0 drain_left.t11 2.2005
R357 drain_left.n0 drain_left.t18 2.2005
R358 drain_left.n15 drain_left.t12 2.2005
R359 drain_left.n15 drain_left.t13 2.2005
R360 drain_left.n13 drain_left.t8 2.2005
R361 drain_left.n13 drain_left.t10 2.2005
R362 drain_left.n11 drain_left.t3 2.2005
R363 drain_left.n11 drain_left.t7 2.2005
R364 drain_left.n9 drain_left.t4 2.2005
R365 drain_left.n9 drain_left.t6 2.2005
R366 drain_left.n8 drain_left.t1 2.2005
R367 drain_left.n8 drain_left.t2 2.2005
R368 drain_left.n12 drain_left.n10 0.974638
R369 drain_left.n14 drain_left.n12 0.974638
R370 drain_left.n16 drain_left.n14 0.974638
R371 drain_left.n7 drain_left.n6 0.919292
R372 drain_left.n7 drain_left.n2 0.919292
C0 drain_right plus 0.478206f
C1 minus source 10.687f
C2 minus plus 6.58275f
C3 plus source 10.7011f
C4 drain_right drain_left 1.72917f
C5 minus drain_left 0.17405f
C6 drain_left source 17.9505f
C7 plus drain_left 10.648901f
C8 drain_right minus 10.328501f
C9 drain_right source 17.9534f
C10 drain_right a_n3202_n2688# 6.96503f
C11 drain_left a_n3202_n2688# 7.4105f
C12 source a_n3202_n2688# 7.881482f
C13 minus a_n3202_n2688# 12.733248f
C14 plus a_n3202_n2688# 14.37077f
C15 drain_left.t11 a_n3202_n2688# 0.189679f
C16 drain_left.t18 a_n3202_n2688# 0.189679f
C17 drain_left.n0 a_n3202_n2688# 1.6648f
C18 drain_left.t0 a_n3202_n2688# 0.189679f
C19 drain_left.t16 a_n3202_n2688# 0.189679f
C20 drain_left.n1 a_n3202_n2688# 1.65906f
C21 drain_left.n2 a_n3202_n2688# 0.763037f
C22 drain_left.t5 a_n3202_n2688# 0.189679f
C23 drain_left.t15 a_n3202_n2688# 0.189679f
C24 drain_left.n3 a_n3202_n2688# 1.65906f
C25 drain_left.t17 a_n3202_n2688# 0.189679f
C26 drain_left.t9 a_n3202_n2688# 0.189679f
C27 drain_left.n4 a_n3202_n2688# 1.6648f
C28 drain_left.t19 a_n3202_n2688# 0.189679f
C29 drain_left.t14 a_n3202_n2688# 0.189679f
C30 drain_left.n5 a_n3202_n2688# 1.65906f
C31 drain_left.n6 a_n3202_n2688# 0.763037f
C32 drain_left.n7 a_n3202_n2688# 1.82935f
C33 drain_left.t1 a_n3202_n2688# 0.189679f
C34 drain_left.t2 a_n3202_n2688# 0.189679f
C35 drain_left.n8 a_n3202_n2688# 1.6648f
C36 drain_left.t4 a_n3202_n2688# 0.189679f
C37 drain_left.t6 a_n3202_n2688# 0.189679f
C38 drain_left.n9 a_n3202_n2688# 1.65906f
C39 drain_left.n10 a_n3202_n2688# 0.767114f
C40 drain_left.t3 a_n3202_n2688# 0.189679f
C41 drain_left.t7 a_n3202_n2688# 0.189679f
C42 drain_left.n11 a_n3202_n2688# 1.65906f
C43 drain_left.n12 a_n3202_n2688# 0.381055f
C44 drain_left.t8 a_n3202_n2688# 0.189679f
C45 drain_left.t10 a_n3202_n2688# 0.189679f
C46 drain_left.n13 a_n3202_n2688# 1.65906f
C47 drain_left.n14 a_n3202_n2688# 0.381055f
C48 drain_left.t12 a_n3202_n2688# 0.189679f
C49 drain_left.t13 a_n3202_n2688# 0.189679f
C50 drain_left.n15 a_n3202_n2688# 1.65906f
C51 drain_left.n16 a_n3202_n2688# 0.620211f
C52 plus.n0 a_n3202_n2688# 0.038512f
C53 plus.t6 a_n3202_n2688# 0.795222f
C54 plus.t7 a_n3202_n2688# 0.795222f
C55 plus.n1 a_n3202_n2688# 0.038512f
C56 plus.t9 a_n3202_n2688# 0.795222f
C57 plus.n2 a_n3202_n2688# 0.341111f
C58 plus.n3 a_n3202_n2688# 0.05139f
C59 plus.t11 a_n3202_n2688# 0.795222f
C60 plus.t12 a_n3202_n2688# 0.795222f
C61 plus.n4 a_n3202_n2688# 0.038512f
C62 plus.t16 a_n3202_n2688# 0.795222f
C63 plus.n5 a_n3202_n2688# 0.330591f
C64 plus.n6 a_n3202_n2688# 0.064147f
C65 plus.t13 a_n3202_n2688# 0.795222f
C66 plus.t15 a_n3202_n2688# 0.795222f
C67 plus.n7 a_n3202_n2688# 0.064147f
C68 plus.t17 a_n3202_n2688# 0.795222f
C69 plus.n8 a_n3202_n2688# 0.333828f
C70 plus.t18 a_n3202_n2688# 0.816422f
C71 plus.n9 a_n3202_n2688# 0.315354f
C72 plus.n10 a_n3202_n2688# 0.177271f
C73 plus.n11 a_n3202_n2688# 0.008739f
C74 plus.n12 a_n3202_n2688# 0.341111f
C75 plus.n13 a_n3202_n2688# 0.341586f
C76 plus.n14 a_n3202_n2688# 0.008739f
C77 plus.n15 a_n3202_n2688# 0.05139f
C78 plus.n16 a_n3202_n2688# 0.038512f
C79 plus.n17 a_n3202_n2688# 0.038512f
C80 plus.n18 a_n3202_n2688# 0.008739f
C81 plus.n19 a_n3202_n2688# 0.330591f
C82 plus.n20 a_n3202_n2688# 0.008739f
C83 plus.n21 a_n3202_n2688# 0.341586f
C84 plus.n22 a_n3202_n2688# 0.064147f
C85 plus.n23 a_n3202_n2688# 0.064147f
C86 plus.n24 a_n3202_n2688# 0.05139f
C87 plus.n25 a_n3202_n2688# 0.008739f
C88 plus.n26 a_n3202_n2688# 0.330591f
C89 plus.n27 a_n3202_n2688# 0.008739f
C90 plus.n28 a_n3202_n2688# 0.330235f
C91 plus.n29 a_n3202_n2688# 0.397345f
C92 plus.n30 a_n3202_n2688# 0.038512f
C93 plus.t8 a_n3202_n2688# 0.795222f
C94 plus.n31 a_n3202_n2688# 0.038512f
C95 plus.t1 a_n3202_n2688# 0.795222f
C96 plus.t19 a_n3202_n2688# 0.795222f
C97 plus.n32 a_n3202_n2688# 0.341111f
C98 plus.n33 a_n3202_n2688# 0.05139f
C99 plus.t3 a_n3202_n2688# 0.795222f
C100 plus.n34 a_n3202_n2688# 0.038512f
C101 plus.t14 a_n3202_n2688# 0.795222f
C102 plus.t4 a_n3202_n2688# 0.795222f
C103 plus.n35 a_n3202_n2688# 0.330591f
C104 plus.n36 a_n3202_n2688# 0.064147f
C105 plus.t0 a_n3202_n2688# 0.795222f
C106 plus.n37 a_n3202_n2688# 0.064147f
C107 plus.t5 a_n3202_n2688# 0.795222f
C108 plus.t2 a_n3202_n2688# 0.795222f
C109 plus.n38 a_n3202_n2688# 0.333828f
C110 plus.t10 a_n3202_n2688# 0.816422f
C111 plus.n39 a_n3202_n2688# 0.315354f
C112 plus.n40 a_n3202_n2688# 0.177271f
C113 plus.n41 a_n3202_n2688# 0.008739f
C114 plus.n42 a_n3202_n2688# 0.341111f
C115 plus.n43 a_n3202_n2688# 0.341586f
C116 plus.n44 a_n3202_n2688# 0.008739f
C117 plus.n45 a_n3202_n2688# 0.05139f
C118 plus.n46 a_n3202_n2688# 0.038512f
C119 plus.n47 a_n3202_n2688# 0.038512f
C120 plus.n48 a_n3202_n2688# 0.008739f
C121 plus.n49 a_n3202_n2688# 0.330591f
C122 plus.n50 a_n3202_n2688# 0.008739f
C123 plus.n51 a_n3202_n2688# 0.341586f
C124 plus.n52 a_n3202_n2688# 0.064147f
C125 plus.n53 a_n3202_n2688# 0.064147f
C126 plus.n54 a_n3202_n2688# 0.05139f
C127 plus.n55 a_n3202_n2688# 0.008739f
C128 plus.n56 a_n3202_n2688# 0.330591f
C129 plus.n57 a_n3202_n2688# 0.008739f
C130 plus.n58 a_n3202_n2688# 0.330235f
C131 plus.n59 a_n3202_n2688# 1.36032f
C132 drain_right.t2 a_n3202_n2688# 0.188377f
C133 drain_right.t17 a_n3202_n2688# 0.188377f
C134 drain_right.n0 a_n3202_n2688# 1.65337f
C135 drain_right.t11 a_n3202_n2688# 0.188377f
C136 drain_right.t18 a_n3202_n2688# 0.188377f
C137 drain_right.n1 a_n3202_n2688# 1.64767f
C138 drain_right.n2 a_n3202_n2688# 0.757798f
C139 drain_right.t4 a_n3202_n2688# 0.188377f
C140 drain_right.t19 a_n3202_n2688# 0.188377f
C141 drain_right.n3 a_n3202_n2688# 1.64767f
C142 drain_right.t9 a_n3202_n2688# 0.188377f
C143 drain_right.t0 a_n3202_n2688# 0.188377f
C144 drain_right.n4 a_n3202_n2688# 1.65337f
C145 drain_right.t13 a_n3202_n2688# 0.188377f
C146 drain_right.t1 a_n3202_n2688# 0.188377f
C147 drain_right.n5 a_n3202_n2688# 1.64767f
C148 drain_right.n6 a_n3202_n2688# 0.757798f
C149 drain_right.n7 a_n3202_n2688# 1.76342f
C150 drain_right.t14 a_n3202_n2688# 0.188377f
C151 drain_right.t10 a_n3202_n2688# 0.188377f
C152 drain_right.n8 a_n3202_n2688# 1.65336f
C153 drain_right.t7 a_n3202_n2688# 0.188377f
C154 drain_right.t15 a_n3202_n2688# 0.188377f
C155 drain_right.n9 a_n3202_n2688# 1.64767f
C156 drain_right.n10 a_n3202_n2688# 0.761854f
C157 drain_right.t8 a_n3202_n2688# 0.188377f
C158 drain_right.t5 a_n3202_n2688# 0.188377f
C159 drain_right.n11 a_n3202_n2688# 1.64767f
C160 drain_right.n12 a_n3202_n2688# 0.378439f
C161 drain_right.t3 a_n3202_n2688# 0.188377f
C162 drain_right.t12 a_n3202_n2688# 0.188377f
C163 drain_right.n13 a_n3202_n2688# 1.64767f
C164 drain_right.n14 a_n3202_n2688# 0.378439f
C165 drain_right.t16 a_n3202_n2688# 0.188377f
C166 drain_right.t6 a_n3202_n2688# 0.188377f
C167 drain_right.n15 a_n3202_n2688# 1.64767f
C168 drain_right.n16 a_n3202_n2688# 0.615945f
C169 source.t4 a_n3202_n2688# 1.85178f
C170 source.n0 a_n3202_n2688# 1.12151f
C171 source.t12 a_n3202_n2688# 0.173657f
C172 source.t3 a_n3202_n2688# 0.173657f
C173 source.n1 a_n3202_n2688# 1.45374f
C174 source.n2 a_n3202_n2688# 0.380858f
C175 source.t18 a_n3202_n2688# 0.173657f
C176 source.t17 a_n3202_n2688# 0.173657f
C177 source.n3 a_n3202_n2688# 1.45374f
C178 source.n4 a_n3202_n2688# 0.380858f
C179 source.t13 a_n3202_n2688# 0.173657f
C180 source.t0 a_n3202_n2688# 0.173657f
C181 source.n5 a_n3202_n2688# 1.45374f
C182 source.n6 a_n3202_n2688# 0.380858f
C183 source.t14 a_n3202_n2688# 0.173657f
C184 source.t1 a_n3202_n2688# 0.173657f
C185 source.n7 a_n3202_n2688# 1.45374f
C186 source.n8 a_n3202_n2688# 0.380858f
C187 source.t7 a_n3202_n2688# 1.85179f
C188 source.n9 a_n3202_n2688# 0.416743f
C189 source.t21 a_n3202_n2688# 1.85179f
C190 source.n10 a_n3202_n2688# 0.416743f
C191 source.t35 a_n3202_n2688# 0.173657f
C192 source.t36 a_n3202_n2688# 0.173657f
C193 source.n11 a_n3202_n2688# 1.45374f
C194 source.n12 a_n3202_n2688# 0.380858f
C195 source.t22 a_n3202_n2688# 0.173657f
C196 source.t37 a_n3202_n2688# 0.173657f
C197 source.n13 a_n3202_n2688# 1.45374f
C198 source.n14 a_n3202_n2688# 0.380858f
C199 source.t25 a_n3202_n2688# 0.173657f
C200 source.t28 a_n3202_n2688# 0.173657f
C201 source.n15 a_n3202_n2688# 1.45374f
C202 source.n16 a_n3202_n2688# 0.380858f
C203 source.t19 a_n3202_n2688# 0.173657f
C204 source.t30 a_n3202_n2688# 0.173657f
C205 source.n17 a_n3202_n2688# 1.45374f
C206 source.n18 a_n3202_n2688# 0.380858f
C207 source.t34 a_n3202_n2688# 1.85179f
C208 source.n19 a_n3202_n2688# 1.48743f
C209 source.t39 a_n3202_n2688# 1.85178f
C210 source.n20 a_n3202_n2688# 1.48743f
C211 source.t2 a_n3202_n2688# 0.173657f
C212 source.t6 a_n3202_n2688# 0.173657f
C213 source.n21 a_n3202_n2688# 1.45374f
C214 source.n22 a_n3202_n2688# 0.380862f
C215 source.t11 a_n3202_n2688# 0.173657f
C216 source.t16 a_n3202_n2688# 0.173657f
C217 source.n23 a_n3202_n2688# 1.45374f
C218 source.n24 a_n3202_n2688# 0.380862f
C219 source.t10 a_n3202_n2688# 0.173657f
C220 source.t15 a_n3202_n2688# 0.173657f
C221 source.n25 a_n3202_n2688# 1.45374f
C222 source.n26 a_n3202_n2688# 0.380862f
C223 source.t8 a_n3202_n2688# 0.173657f
C224 source.t9 a_n3202_n2688# 0.173657f
C225 source.n27 a_n3202_n2688# 1.45374f
C226 source.n28 a_n3202_n2688# 0.380862f
C227 source.t5 a_n3202_n2688# 1.85178f
C228 source.n29 a_n3202_n2688# 0.416747f
C229 source.t38 a_n3202_n2688# 1.85178f
C230 source.n30 a_n3202_n2688# 0.416747f
C231 source.t33 a_n3202_n2688# 0.173657f
C232 source.t27 a_n3202_n2688# 0.173657f
C233 source.n31 a_n3202_n2688# 1.45374f
C234 source.n32 a_n3202_n2688# 0.380862f
C235 source.t32 a_n3202_n2688# 0.173657f
C236 source.t24 a_n3202_n2688# 0.173657f
C237 source.n33 a_n3202_n2688# 1.45374f
C238 source.n34 a_n3202_n2688# 0.380862f
C239 source.t31 a_n3202_n2688# 0.173657f
C240 source.t20 a_n3202_n2688# 0.173657f
C241 source.n35 a_n3202_n2688# 1.45374f
C242 source.n36 a_n3202_n2688# 0.380862f
C243 source.t26 a_n3202_n2688# 0.173657f
C244 source.t29 a_n3202_n2688# 0.173657f
C245 source.n37 a_n3202_n2688# 1.45374f
C246 source.n38 a_n3202_n2688# 0.380862f
C247 source.t23 a_n3202_n2688# 1.85178f
C248 source.n39 a_n3202_n2688# 0.581307f
C249 source.n40 a_n3202_n2688# 1.28941f
C250 minus.n0 a_n3202_n2688# 0.037992f
C251 minus.n1 a_n3202_n2688# 0.008621f
C252 minus.t13 a_n3202_n2688# 0.784482f
C253 minus.n2 a_n3202_n2688# 0.063281f
C254 minus.t11 a_n3202_n2688# 0.784482f
C255 minus.n3 a_n3202_n2688# 0.326126f
C256 minus.n4 a_n3202_n2688# 0.037992f
C257 minus.t12 a_n3202_n2688# 0.784482f
C258 minus.n5 a_n3202_n2688# 0.336973f
C259 minus.n6 a_n3202_n2688# 0.174876f
C260 minus.t9 a_n3202_n2688# 0.805394f
C261 minus.n7 a_n3202_n2688# 0.311094f
C262 minus.t5 a_n3202_n2688# 0.784482f
C263 minus.n8 a_n3202_n2688# 0.329319f
C264 minus.n9 a_n3202_n2688# 0.008621f
C265 minus.t4 a_n3202_n2688# 0.784482f
C266 minus.n10 a_n3202_n2688# 0.336504f
C267 minus.n11 a_n3202_n2688# 0.063281f
C268 minus.n12 a_n3202_n2688# 0.063281f
C269 minus.n13 a_n3202_n2688# 0.050696f
C270 minus.n14 a_n3202_n2688# 0.008621f
C271 minus.t14 a_n3202_n2688# 0.784482f
C272 minus.n15 a_n3202_n2688# 0.326126f
C273 minus.n16 a_n3202_n2688# 0.008621f
C274 minus.n17 a_n3202_n2688# 0.037992f
C275 minus.n18 a_n3202_n2688# 0.037992f
C276 minus.n19 a_n3202_n2688# 0.050696f
C277 minus.n20 a_n3202_n2688# 0.008621f
C278 minus.t7 a_n3202_n2688# 0.784482f
C279 minus.n21 a_n3202_n2688# 0.336973f
C280 minus.t16 a_n3202_n2688# 0.784482f
C281 minus.n22 a_n3202_n2688# 0.336504f
C282 minus.n23 a_n3202_n2688# 0.063281f
C283 minus.n24 a_n3202_n2688# 0.050696f
C284 minus.n25 a_n3202_n2688# 0.037992f
C285 minus.n26 a_n3202_n2688# 0.326126f
C286 minus.n27 a_n3202_n2688# 0.008621f
C287 minus.t3 a_n3202_n2688# 0.784482f
C288 minus.n28 a_n3202_n2688# 0.325775f
C289 minus.n29 a_n3202_n2688# 1.52245f
C290 minus.n30 a_n3202_n2688# 0.037992f
C291 minus.n31 a_n3202_n2688# 0.008621f
C292 minus.n32 a_n3202_n2688# 0.063281f
C293 minus.t0 a_n3202_n2688# 0.784482f
C294 minus.n33 a_n3202_n2688# 0.326126f
C295 minus.n34 a_n3202_n2688# 0.037992f
C296 minus.t1 a_n3202_n2688# 0.784482f
C297 minus.n35 a_n3202_n2688# 0.336973f
C298 minus.n36 a_n3202_n2688# 0.174876f
C299 minus.t17 a_n3202_n2688# 0.805394f
C300 minus.n37 a_n3202_n2688# 0.311094f
C301 minus.t2 a_n3202_n2688# 0.784482f
C302 minus.n38 a_n3202_n2688# 0.329319f
C303 minus.n39 a_n3202_n2688# 0.008621f
C304 minus.t8 a_n3202_n2688# 0.784482f
C305 minus.n40 a_n3202_n2688# 0.336504f
C306 minus.n41 a_n3202_n2688# 0.063281f
C307 minus.n42 a_n3202_n2688# 0.063281f
C308 minus.n43 a_n3202_n2688# 0.050696f
C309 minus.n44 a_n3202_n2688# 0.008621f
C310 minus.t15 a_n3202_n2688# 0.784482f
C311 minus.n45 a_n3202_n2688# 0.326126f
C312 minus.n46 a_n3202_n2688# 0.008621f
C313 minus.n47 a_n3202_n2688# 0.037992f
C314 minus.n48 a_n3202_n2688# 0.037992f
C315 minus.n49 a_n3202_n2688# 0.050696f
C316 minus.n50 a_n3202_n2688# 0.008621f
C317 minus.t6 a_n3202_n2688# 0.784482f
C318 minus.n51 a_n3202_n2688# 0.336973f
C319 minus.t18 a_n3202_n2688# 0.784482f
C320 minus.n52 a_n3202_n2688# 0.336504f
C321 minus.n53 a_n3202_n2688# 0.063281f
C322 minus.n54 a_n3202_n2688# 0.050696f
C323 minus.n55 a_n3202_n2688# 0.037992f
C324 minus.t10 a_n3202_n2688# 0.784482f
C325 minus.n56 a_n3202_n2688# 0.326126f
C326 minus.n57 a_n3202_n2688# 0.008621f
C327 minus.t19 a_n3202_n2688# 0.784482f
C328 minus.n58 a_n3202_n2688# 0.325775f
C329 minus.n59 a_n3202_n2688# 0.266561f
C330 minus.n60 a_n3202_n2688# 1.828f
.ends

