* NGSPICE file created from diffpair246.ext - technology: sky130A

.subckt diffpair246 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t6 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X1 drain_right.t13 minus.t0 source.t7 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X2 drain_left.t3 plus.t1 source.t26 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X3 drain_left.t11 plus.t2 source.t25 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X4 source.t2 minus.t1 drain_right.t12 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X5 a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X6 source.t0 minus.t2 drain_right.t11 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 source.t24 plus.t3 drain_left.t8 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 drain_right.t10 minus.t3 source.t1 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X9 a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X10 drain_right.t9 minus.t4 source.t4 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X11 source.t10 minus.t5 drain_right.t8 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X12 drain_right.t7 minus.t6 source.t6 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X13 drain_right.t6 minus.t7 source.t12 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X14 source.t13 minus.t8 drain_right.t5 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 source.t5 minus.t9 drain_right.t4 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X16 drain_left.t4 plus.t4 source.t23 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X17 drain_right.t3 minus.t10 source.t8 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_right.t2 minus.t11 source.t11 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X19 drain_right.t1 minus.t12 source.t3 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X20 source.t22 plus.t5 drain_left.t1 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X21 source.t21 plus.t6 drain_left.t9 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 source.t9 minus.t13 drain_right.t0 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X23 drain_left.t13 plus.t7 source.t20 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X24 drain_left.t7 plus.t8 source.t19 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X25 a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X26 drain_left.t2 plus.t9 source.t18 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X27 source.t17 plus.t10 drain_left.t12 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X28 source.t16 plus.t11 drain_left.t10 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X29 a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X30 drain_left.t5 plus.t12 source.t15 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X31 drain_left.t0 plus.t13 source.t14 a_n1756_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
R0 plus.n3 plus.t4 1238.59
R1 plus.n15 plus.t7 1238.59
R2 plus.n20 plus.t1 1238.59
R3 plus.n32 plus.t12 1238.59
R4 plus.n1 plus.t6 1172.87
R5 plus.n4 plus.t11 1172.87
R6 plus.n6 plus.t8 1172.87
R7 plus.n12 plus.t13 1172.87
R8 plus.n14 plus.t10 1172.87
R9 plus.n18 plus.t0 1172.87
R10 plus.n21 plus.t3 1172.87
R11 plus.n23 plus.t9 1172.87
R12 plus.n29 plus.t2 1172.87
R13 plus.n31 plus.t5 1172.87
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 51.1217
R33 plus.n13 plus.n12 51.1217
R34 plus.n30 plus.n29 51.1217
R35 plus.n23 plus.n22 51.1217
R36 plus.n5 plus.n4 43.8187
R37 plus.n14 plus.n13 43.8187
R38 plus.n31 plus.n30 43.8187
R39 plus.n22 plus.n21 43.8187
R40 plus.n4 plus.n3 29.2126
R41 plus.n15 plus.n14 29.2126
R42 plus.n32 plus.n31 29.2126
R43 plus.n21 plus.n20 29.2126
R44 plus plus.n33 27.4517
R45 plus.n7 plus.n6 21.9096
R46 plus.n12 plus.n11 21.9096
R47 plus.n29 plus.n28 21.9096
R48 plus.n24 plus.n23 21.9096
R49 plus plus.n16 9.94179
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t4 72.7512
R61 drain_left.n1 drain_left.t5 72.751
R62 drain_left.n4 drain_left.n2 67.751
R63 drain_left.n9 drain_left.n8 67.1908
R64 drain_left.n7 drain_left.n6 67.1908
R65 drain_left.n11 drain_left.n10 67.1907
R66 drain_left.n4 drain_left.n3 67.1907
R67 drain_left.n1 drain_left.n0 67.1907
R68 drain_left drain_left.n5 26.0436
R69 drain_left drain_left.n11 6.21356
R70 drain_left.n2 drain_left.t8 5.0005
R71 drain_left.n2 drain_left.t3 5.0005
R72 drain_left.n3 drain_left.t6 5.0005
R73 drain_left.n3 drain_left.t2 5.0005
R74 drain_left.n0 drain_left.t1 5.0005
R75 drain_left.n0 drain_left.t11 5.0005
R76 drain_left.n10 drain_left.t12 5.0005
R77 drain_left.n10 drain_left.t13 5.0005
R78 drain_left.n8 drain_left.t9 5.0005
R79 drain_left.n8 drain_left.t0 5.0005
R80 drain_left.n6 drain_left.t10 5.0005
R81 drain_left.n6 drain_left.t7 5.0005
R82 drain_left.n9 drain_left.n7 0.560845
R83 drain_left.n11 drain_left.n9 0.560845
R84 drain_left.n5 drain_left.n1 0.365413
R85 drain_left.n5 drain_left.n4 0.0852402
R86 source.n7 source.t6 55.512
R87 source.n0 source.t20 55.5119
R88 source.n27 source.t4 55.5119
R89 source.n20 source.t26 55.5119
R90 source.n2 source.n1 50.512
R91 source.n4 source.n3 50.512
R92 source.n6 source.n5 50.512
R93 source.n9 source.n8 50.512
R94 source.n11 source.n10 50.512
R95 source.n13 source.n12 50.512
R96 source.n26 source.n25 50.5119
R97 source.n24 source.n23 50.5119
R98 source.n22 source.n21 50.5119
R99 source.n19 source.n18 50.5119
R100 source.n17 source.n16 50.5119
R101 source.n15 source.n14 50.5119
R102 source.n15 source.n13 17.863
R103 source.n28 source.n0 11.7595
R104 source.n28 source.n27 5.5436
R105 source.n25 source.t7 5.0005
R106 source.n25 source.t0 5.0005
R107 source.n23 source.t1 5.0005
R108 source.n23 source.t13 5.0005
R109 source.n21 source.t3 5.0005
R110 source.n21 source.t2 5.0005
R111 source.n18 source.t18 5.0005
R112 source.n18 source.t24 5.0005
R113 source.n16 source.t25 5.0005
R114 source.n16 source.t27 5.0005
R115 source.n14 source.t15 5.0005
R116 source.n14 source.t22 5.0005
R117 source.n1 source.t14 5.0005
R118 source.n1 source.t17 5.0005
R119 source.n3 source.t19 5.0005
R120 source.n3 source.t21 5.0005
R121 source.n5 source.t23 5.0005
R122 source.n5 source.t16 5.0005
R123 source.n8 source.t8 5.0005
R124 source.n8 source.t10 5.0005
R125 source.n10 source.t12 5.0005
R126 source.n10 source.t5 5.0005
R127 source.n12 source.t11 5.0005
R128 source.n12 source.t9 5.0005
R129 source.n7 source.n6 0.7505
R130 source.n22 source.n20 0.7505
R131 source.n13 source.n11 0.560845
R132 source.n11 source.n9 0.560845
R133 source.n9 source.n7 0.560845
R134 source.n6 source.n4 0.560845
R135 source.n4 source.n2 0.560845
R136 source.n2 source.n0 0.560845
R137 source.n17 source.n15 0.560845
R138 source.n19 source.n17 0.560845
R139 source.n20 source.n19 0.560845
R140 source.n24 source.n22 0.560845
R141 source.n26 source.n24 0.560845
R142 source.n27 source.n26 0.560845
R143 source source.n28 0.188
R144 minus.n15 minus.t11 1238.59
R145 minus.n3 minus.t6 1238.59
R146 minus.n32 minus.t4 1238.59
R147 minus.n20 minus.t12 1238.59
R148 minus.n1 minus.t9 1172.87
R149 minus.n14 minus.t13 1172.87
R150 minus.n12 minus.t7 1172.87
R151 minus.n6 minus.t10 1172.87
R152 minus.n4 minus.t5 1172.87
R153 minus.n18 minus.t8 1172.87
R154 minus.n31 minus.t2 1172.87
R155 minus.n29 minus.t0 1172.87
R156 minus.n23 minus.t3 1172.87
R157 minus.n21 minus.t1 1172.87
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 51.1217
R177 minus.n6 minus.n5 51.1217
R178 minus.n23 minus.n22 51.1217
R179 minus.n30 minus.n29 51.1217
R180 minus.n14 minus.n13 43.8187
R181 minus.n5 minus.n4 43.8187
R182 minus.n22 minus.n21 43.8187
R183 minus.n31 minus.n30 43.8187
R184 minus.n34 minus.n16 31.2978
R185 minus.n15 minus.n14 29.2126
R186 minus.n4 minus.n3 29.2126
R187 minus.n21 minus.n20 29.2126
R188 minus.n32 minus.n31 29.2126
R189 minus.n12 minus.n11 21.9096
R190 minus.n7 minus.n6 21.9096
R191 minus.n24 minus.n23 21.9096
R192 minus.n29 minus.n28 21.9096
R193 minus.n34 minus.n33 6.57058
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t1 72.751
R206 drain_right.n11 drain_right.t2 72.1908
R207 drain_right.n8 drain_right.n6 67.751
R208 drain_right.n4 drain_right.n2 67.751
R209 drain_right.n8 drain_right.n7 67.1908
R210 drain_right.n10 drain_right.n9 67.1908
R211 drain_right.n4 drain_right.n3 67.1907
R212 drain_right.n1 drain_right.n0 67.1907
R213 drain_right drain_right.n5 25.4904
R214 drain_right drain_right.n11 5.93339
R215 drain_right.n2 drain_right.t11 5.0005
R216 drain_right.n2 drain_right.t9 5.0005
R217 drain_right.n3 drain_right.t5 5.0005
R218 drain_right.n3 drain_right.t13 5.0005
R219 drain_right.n0 drain_right.t12 5.0005
R220 drain_right.n0 drain_right.t10 5.0005
R221 drain_right.n6 drain_right.t8 5.0005
R222 drain_right.n6 drain_right.t7 5.0005
R223 drain_right.n7 drain_right.t4 5.0005
R224 drain_right.n7 drain_right.t3 5.0005
R225 drain_right.n9 drain_right.t0 5.0005
R226 drain_right.n9 drain_right.t6 5.0005
R227 drain_right.n11 drain_right.n10 0.560845
R228 drain_right.n10 drain_right.n8 0.560845
R229 drain_right.n5 drain_right.n1 0.365413
R230 drain_right.n5 drain_right.n4 0.0852402
C0 drain_right minus 1.83538f
C1 drain_right plus 0.325058f
C2 plus minus 4.21286f
C3 drain_right drain_left 0.898966f
C4 drain_right source 15.6431f
C5 minus drain_left 0.171187f
C6 plus drain_left 2.00403f
C7 minus source 1.68136f
C8 plus source 1.6957f
C9 source drain_left 15.6486f
C10 drain_right a_n1756_n2088# 5.0588f
C11 drain_left a_n1756_n2088# 5.52754f
C12 source a_n1756_n2088# 4.068465f
C13 minus a_n1756_n2088# 5.970701f
C14 plus a_n1756_n2088# 7.28496f
C15 drain_right.t1 a_n1756_n2088# 1.25857f
C16 drain_right.t12 a_n1756_n2088# 0.167465f
C17 drain_right.t10 a_n1756_n2088# 0.167465f
C18 drain_right.n0 a_n1756_n2088# 1.03567f
C19 drain_right.n1 a_n1756_n2088# 0.579394f
C20 drain_right.t11 a_n1756_n2088# 0.167465f
C21 drain_right.t9 a_n1756_n2088# 0.167465f
C22 drain_right.n2 a_n1756_n2088# 1.03801f
C23 drain_right.t5 a_n1756_n2088# 0.167465f
C24 drain_right.t13 a_n1756_n2088# 0.167465f
C25 drain_right.n3 a_n1756_n2088# 1.03567f
C26 drain_right.n4 a_n1756_n2088# 0.524463f
C27 drain_right.n5 a_n1756_n2088# 0.767118f
C28 drain_right.t8 a_n1756_n2088# 0.167465f
C29 drain_right.t7 a_n1756_n2088# 0.167465f
C30 drain_right.n6 a_n1756_n2088# 1.03801f
C31 drain_right.t4 a_n1756_n2088# 0.167465f
C32 drain_right.t3 a_n1756_n2088# 0.167465f
C33 drain_right.n7 a_n1756_n2088# 1.03567f
C34 drain_right.n8 a_n1756_n2088# 0.553806f
C35 drain_right.t0 a_n1756_n2088# 0.167465f
C36 drain_right.t6 a_n1756_n2088# 0.167465f
C37 drain_right.n9 a_n1756_n2088# 1.03567f
C38 drain_right.n10 a_n1756_n2088# 0.273376f
C39 drain_right.t2 a_n1756_n2088# 1.2561f
C40 drain_right.n11 a_n1756_n2088# 0.517156f
C41 minus.n0 a_n1756_n2088# 0.029376f
C42 minus.t11 a_n1756_n2088# 0.0775f
C43 minus.t13 a_n1756_n2088# 0.075329f
C44 minus.t7 a_n1756_n2088# 0.075329f
C45 minus.t9 a_n1756_n2088# 0.075329f
C46 minus.n1 a_n1756_n2088# 0.04885f
C47 minus.n2 a_n1756_n2088# 0.068668f
C48 minus.t10 a_n1756_n2088# 0.075329f
C49 minus.t5 a_n1756_n2088# 0.075329f
C50 minus.t6 a_n1756_n2088# 0.0775f
C51 minus.n3 a_n1756_n2088# 0.051253f
C52 minus.n4 a_n1756_n2088# 0.039105f
C53 minus.n5 a_n1756_n2088# 0.012462f
C54 minus.n6 a_n1756_n2088# 0.039105f
C55 minus.n7 a_n1756_n2088# 0.012462f
C56 minus.n8 a_n1756_n2088# 0.029376f
C57 minus.n9 a_n1756_n2088# 0.029376f
C58 minus.n10 a_n1756_n2088# 0.029376f
C59 minus.n11 a_n1756_n2088# 0.012462f
C60 minus.n12 a_n1756_n2088# 0.039105f
C61 minus.n13 a_n1756_n2088# 0.012462f
C62 minus.n14 a_n1756_n2088# 0.039105f
C63 minus.n15 a_n1756_n2088# 0.051207f
C64 minus.n16 a_n1756_n2088# 0.822741f
C65 minus.n17 a_n1756_n2088# 0.029376f
C66 minus.t2 a_n1756_n2088# 0.075329f
C67 minus.t0 a_n1756_n2088# 0.075329f
C68 minus.t8 a_n1756_n2088# 0.075329f
C69 minus.n18 a_n1756_n2088# 0.04885f
C70 minus.n19 a_n1756_n2088# 0.068668f
C71 minus.t3 a_n1756_n2088# 0.075329f
C72 minus.t1 a_n1756_n2088# 0.075329f
C73 minus.t12 a_n1756_n2088# 0.0775f
C74 minus.n20 a_n1756_n2088# 0.051253f
C75 minus.n21 a_n1756_n2088# 0.039105f
C76 minus.n22 a_n1756_n2088# 0.012462f
C77 minus.n23 a_n1756_n2088# 0.039105f
C78 minus.n24 a_n1756_n2088# 0.012462f
C79 minus.n25 a_n1756_n2088# 0.029376f
C80 minus.n26 a_n1756_n2088# 0.029376f
C81 minus.n27 a_n1756_n2088# 0.029376f
C82 minus.n28 a_n1756_n2088# 0.012462f
C83 minus.n29 a_n1756_n2088# 0.039105f
C84 minus.n30 a_n1756_n2088# 0.012462f
C85 minus.n31 a_n1756_n2088# 0.039105f
C86 minus.t4 a_n1756_n2088# 0.0775f
C87 minus.n32 a_n1756_n2088# 0.051207f
C88 minus.n33 a_n1756_n2088# 0.196924f
C89 minus.n34 a_n1756_n2088# 1.01025f
C90 source.t20 a_n1756_n2088# 1.26929f
C91 source.n0 a_n1756_n2088# 0.933789f
C92 source.t14 a_n1756_n2088# 0.180713f
C93 source.t17 a_n1756_n2088# 0.180713f
C94 source.n1 a_n1756_n2088# 1.05177f
C95 source.n2 a_n1756_n2088# 0.326644f
C96 source.t19 a_n1756_n2088# 0.180713f
C97 source.t21 a_n1756_n2088# 0.180713f
C98 source.n3 a_n1756_n2088# 1.05177f
C99 source.n4 a_n1756_n2088# 0.326644f
C100 source.t23 a_n1756_n2088# 0.180713f
C101 source.t16 a_n1756_n2088# 0.180713f
C102 source.n5 a_n1756_n2088# 1.05177f
C103 source.n6 a_n1756_n2088# 0.342017f
C104 source.t6 a_n1756_n2088# 1.2693f
C105 source.n7 a_n1756_n2088# 0.449773f
C106 source.t8 a_n1756_n2088# 0.180713f
C107 source.t10 a_n1756_n2088# 0.180713f
C108 source.n8 a_n1756_n2088# 1.05177f
C109 source.n9 a_n1756_n2088# 0.326644f
C110 source.t12 a_n1756_n2088# 0.180713f
C111 source.t5 a_n1756_n2088# 0.180713f
C112 source.n10 a_n1756_n2088# 1.05177f
C113 source.n11 a_n1756_n2088# 0.326644f
C114 source.t11 a_n1756_n2088# 0.180713f
C115 source.t9 a_n1756_n2088# 0.180713f
C116 source.n12 a_n1756_n2088# 1.05177f
C117 source.n13 a_n1756_n2088# 1.19569f
C118 source.t15 a_n1756_n2088# 0.180713f
C119 source.t22 a_n1756_n2088# 0.180713f
C120 source.n14 a_n1756_n2088# 1.05177f
C121 source.n15 a_n1756_n2088# 1.1957f
C122 source.t25 a_n1756_n2088# 0.180713f
C123 source.t27 a_n1756_n2088# 0.180713f
C124 source.n16 a_n1756_n2088# 1.05177f
C125 source.n17 a_n1756_n2088# 0.326651f
C126 source.t18 a_n1756_n2088# 0.180713f
C127 source.t24 a_n1756_n2088# 0.180713f
C128 source.n18 a_n1756_n2088# 1.05177f
C129 source.n19 a_n1756_n2088# 0.326651f
C130 source.t26 a_n1756_n2088# 1.26929f
C131 source.n20 a_n1756_n2088# 0.449779f
C132 source.t3 a_n1756_n2088# 0.180713f
C133 source.t2 a_n1756_n2088# 0.180713f
C134 source.n21 a_n1756_n2088# 1.05177f
C135 source.n22 a_n1756_n2088# 0.342023f
C136 source.t1 a_n1756_n2088# 0.180713f
C137 source.t13 a_n1756_n2088# 0.180713f
C138 source.n23 a_n1756_n2088# 1.05177f
C139 source.n24 a_n1756_n2088# 0.326651f
C140 source.t7 a_n1756_n2088# 0.180713f
C141 source.t0 a_n1756_n2088# 0.180713f
C142 source.n25 a_n1756_n2088# 1.05177f
C143 source.n26 a_n1756_n2088# 0.326651f
C144 source.t4 a_n1756_n2088# 1.26929f
C145 source.n27 a_n1756_n2088# 0.570187f
C146 source.n28 a_n1756_n2088# 1.02999f
C147 drain_left.t5 a_n1756_n2088# 1.41168f
C148 drain_left.t1 a_n1756_n2088# 0.187837f
C149 drain_left.t11 a_n1756_n2088# 0.187837f
C150 drain_left.n0 a_n1756_n2088# 1.16166f
C151 drain_left.n1 a_n1756_n2088# 0.649877f
C152 drain_left.t8 a_n1756_n2088# 0.187837f
C153 drain_left.t3 a_n1756_n2088# 0.187837f
C154 drain_left.n2 a_n1756_n2088# 1.16428f
C155 drain_left.t6 a_n1756_n2088# 0.187837f
C156 drain_left.t2 a_n1756_n2088# 0.187837f
C157 drain_left.n3 a_n1756_n2088# 1.16166f
C158 drain_left.n4 a_n1756_n2088# 0.588264f
C159 drain_left.n5 a_n1756_n2088# 0.913585f
C160 drain_left.t4 a_n1756_n2088# 1.41168f
C161 drain_left.t10 a_n1756_n2088# 0.187837f
C162 drain_left.t7 a_n1756_n2088# 0.187837f
C163 drain_left.n6 a_n1756_n2088# 1.16166f
C164 drain_left.n7 a_n1756_n2088# 0.664671f
C165 drain_left.t9 a_n1756_n2088# 0.187837f
C166 drain_left.t0 a_n1756_n2088# 0.187837f
C167 drain_left.n8 a_n1756_n2088# 1.16166f
C168 drain_left.n9 a_n1756_n2088# 0.306631f
C169 drain_left.t12 a_n1756_n2088# 0.187837f
C170 drain_left.t13 a_n1756_n2088# 0.187837f
C171 drain_left.n10 a_n1756_n2088# 1.16166f
C172 drain_left.n11 a_n1756_n2088# 0.52499f
C173 plus.n0 a_n1756_n2088# 0.043988f
C174 plus.t10 a_n1756_n2088# 0.112795f
C175 plus.t13 a_n1756_n2088# 0.112795f
C176 plus.t6 a_n1756_n2088# 0.112795f
C177 plus.n1 a_n1756_n2088# 0.073147f
C178 plus.n2 a_n1756_n2088# 0.102822f
C179 plus.t8 a_n1756_n2088# 0.112795f
C180 plus.t11 a_n1756_n2088# 0.112795f
C181 plus.t4 a_n1756_n2088# 0.116046f
C182 plus.n3 a_n1756_n2088# 0.076745f
C183 plus.n4 a_n1756_n2088# 0.058555f
C184 plus.n5 a_n1756_n2088# 0.01866f
C185 plus.n6 a_n1756_n2088# 0.058555f
C186 plus.n7 a_n1756_n2088# 0.01866f
C187 plus.n8 a_n1756_n2088# 0.043988f
C188 plus.n9 a_n1756_n2088# 0.043988f
C189 plus.n10 a_n1756_n2088# 0.043988f
C190 plus.n11 a_n1756_n2088# 0.01866f
C191 plus.n12 a_n1756_n2088# 0.058555f
C192 plus.n13 a_n1756_n2088# 0.01866f
C193 plus.n14 a_n1756_n2088# 0.058555f
C194 plus.t7 a_n1756_n2088# 0.116046f
C195 plus.n15 a_n1756_n2088# 0.076676f
C196 plus.n16 a_n1756_n2088# 0.384536f
C197 plus.n17 a_n1756_n2088# 0.043988f
C198 plus.t12 a_n1756_n2088# 0.116046f
C199 plus.t5 a_n1756_n2088# 0.112795f
C200 plus.t2 a_n1756_n2088# 0.112795f
C201 plus.t0 a_n1756_n2088# 0.112795f
C202 plus.n18 a_n1756_n2088# 0.073147f
C203 plus.n19 a_n1756_n2088# 0.102822f
C204 plus.t9 a_n1756_n2088# 0.112795f
C205 plus.t3 a_n1756_n2088# 0.112795f
C206 plus.t1 a_n1756_n2088# 0.116046f
C207 plus.n20 a_n1756_n2088# 0.076745f
C208 plus.n21 a_n1756_n2088# 0.058555f
C209 plus.n22 a_n1756_n2088# 0.01866f
C210 plus.n23 a_n1756_n2088# 0.058555f
C211 plus.n24 a_n1756_n2088# 0.01866f
C212 plus.n25 a_n1756_n2088# 0.043988f
C213 plus.n26 a_n1756_n2088# 0.043988f
C214 plus.n27 a_n1756_n2088# 0.043988f
C215 plus.n28 a_n1756_n2088# 0.01866f
C216 plus.n29 a_n1756_n2088# 0.058555f
C217 plus.n30 a_n1756_n2088# 0.01866f
C218 plus.n31 a_n1756_n2088# 0.058555f
C219 plus.n32 a_n1756_n2088# 0.076676f
C220 plus.n33 a_n1756_n2088# 1.11355f
.ends

