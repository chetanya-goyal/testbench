* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X1 source.t36 plus.t0 drain_left.t0 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X2 a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X3 drain_right.t19 minus.t0 source.t10 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X4 a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X5 drain_right.t18 minus.t1 source.t16 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X6 drain_right.t17 minus.t2 source.t12 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X7 a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X8 drain_right.t16 minus.t3 source.t38 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X9 source.t35 plus.t1 drain_left.t12 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X10 source.t34 plus.t2 drain_left.t2 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X11 source.t33 plus.t3 drain_left.t3 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X12 source.t7 minus.t4 drain_right.t15 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X13 drain_right.t14 minus.t5 source.t39 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X14 source.t32 plus.t4 drain_left.t16 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X15 drain_right.t13 minus.t6 source.t8 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X16 drain_left.t13 plus.t5 source.t31 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X17 source.t15 minus.t7 drain_right.t12 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X18 drain_right.t11 minus.t8 source.t11 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X19 drain_right.t10 minus.t9 source.t37 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X20 source.t1 minus.t10 drain_right.t9 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X21 source.t30 plus.t6 drain_left.t4 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X22 source.t3 minus.t11 drain_right.t8 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X23 source.t4 minus.t12 drain_right.t7 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X24 drain_left.t8 plus.t7 source.t29 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X25 drain_left.t17 plus.t8 source.t28 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X26 source.t5 minus.t13 drain_right.t6 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X27 drain_right.t5 minus.t14 source.t13 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X28 drain_left.t5 plus.t9 source.t27 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X29 drain_right.t4 minus.t15 source.t0 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X30 drain_left.t14 plus.t10 source.t26 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X31 source.t25 plus.t11 drain_left.t1 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X32 source.t14 minus.t16 drain_right.t3 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X33 drain_left.t6 plus.t12 source.t24 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X34 drain_left.t18 plus.t13 source.t23 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X35 source.t9 minus.t17 drain_right.t2 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X36 source.t2 minus.t18 drain_right.t1 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X37 source.t22 plus.t14 drain_left.t15 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X38 source.t6 minus.t19 drain_right.t0 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X39 source.t21 plus.t15 drain_left.t19 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X40 drain_left.t9 plus.t16 source.t20 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X41 drain_left.t10 plus.t17 source.t19 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X42 source.t18 plus.t18 drain_left.t11 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X43 drain_left.t7 plus.t19 source.t17 a_n3202_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 plus.n11 plus.n10 161.3
R1 plus.n15 plus.n14 161.3
R2 plus.n16 plus.n5 161.3
R3 plus.n18 plus.n17 161.3
R4 plus.n19 plus.n4 161.3
R5 plus.n20 plus.n3 161.3
R6 plus.n25 plus.n24 161.3
R7 plus.n26 plus.n1 161.3
R8 plus.n27 plus.n0 161.3
R9 plus.n29 plus.n28 161.3
R10 plus.n41 plus.n40 161.3
R11 plus.n45 plus.n44 161.3
R12 plus.n46 plus.n35 161.3
R13 plus.n48 plus.n47 161.3
R14 plus.n49 plus.n34 161.3
R15 plus.n50 plus.n33 161.3
R16 plus.n55 plus.n54 161.3
R17 plus.n56 plus.n31 161.3
R18 plus.n57 plus.n30 161.3
R19 plus.n59 plus.n58 161.3
R20 plus.n9 plus.t18 131.144
R21 plus.n39 plus.t17 131.144
R22 plus.n28 plus.t5 109.355
R23 plus.n26 plus.t6 109.355
R24 plus.n2 plus.t8 109.355
R25 plus.n21 plus.t11 109.355
R26 plus.n19 plus.t12 109.355
R27 plus.n5 plus.t15 109.355
R28 plus.n13 plus.t13 109.355
R29 plus.n12 plus.t14 109.355
R30 plus.n8 plus.t16 109.355
R31 plus.n58 plus.t4 109.355
R32 plus.n56 plus.t10 109.355
R33 plus.n32 plus.t0 109.355
R34 plus.n51 plus.t9 109.355
R35 plus.n49 plus.t3 109.355
R36 plus.n35 plus.t7 109.355
R37 plus.n43 plus.t2 109.355
R38 plus.n42 plus.t19 109.355
R39 plus.n38 plus.t1 109.355
R40 plus.n12 plus.n7 80.6037
R41 plus.n13 plus.n6 80.6037
R42 plus.n22 plus.n21 80.6037
R43 plus.n23 plus.n2 80.6037
R44 plus.n42 plus.n37 80.6037
R45 plus.n43 plus.n36 80.6037
R46 plus.n52 plus.n51 80.6037
R47 plus.n53 plus.n32 80.6037
R48 plus.n21 plus.n2 48.2005
R49 plus.n13 plus.n12 48.2005
R50 plus.n51 plus.n32 48.2005
R51 plus.n43 plus.n42 48.2005
R52 plus.n40 plus.n39 44.8565
R53 plus.n10 plus.n9 44.8565
R54 plus.n21 plus.n20 43.0884
R55 plus.n14 plus.n13 43.0884
R56 plus.n51 plus.n50 43.0884
R57 plus.n44 plus.n43 43.0884
R58 plus.n25 plus.n2 40.1672
R59 plus.n12 plus.n11 40.1672
R60 plus.n55 plus.n32 40.1672
R61 plus.n42 plus.n41 40.1672
R62 plus plus.n59 31.5483
R63 plus.n28 plus.n27 27.0217
R64 plus.n58 plus.n57 27.0217
R65 plus.n18 plus.n5 24.1005
R66 plus.n19 plus.n18 24.1005
R67 plus.n49 plus.n48 24.1005
R68 plus.n48 plus.n35 24.1005
R69 plus.n27 plus.n26 21.1793
R70 plus.n57 plus.n56 21.1793
R71 plus.n39 plus.n38 20.1275
R72 plus.n9 plus.n8 20.1275
R73 plus plus.n29 8.56111
R74 plus.n26 plus.n25 8.03383
R75 plus.n11 plus.n8 8.03383
R76 plus.n56 plus.n55 8.03383
R77 plus.n41 plus.n38 8.03383
R78 plus.n20 plus.n19 5.11262
R79 plus.n14 plus.n5 5.11262
R80 plus.n50 plus.n49 5.11262
R81 plus.n44 plus.n35 5.11262
R82 plus.n7 plus.n6 0.380177
R83 plus.n23 plus.n22 0.380177
R84 plus.n53 plus.n52 0.380177
R85 plus.n37 plus.n36 0.380177
R86 plus.n10 plus.n7 0.285035
R87 plus.n15 plus.n6 0.285035
R88 plus.n22 plus.n3 0.285035
R89 plus.n24 plus.n23 0.285035
R90 plus.n54 plus.n53 0.285035
R91 plus.n52 plus.n33 0.285035
R92 plus.n45 plus.n36 0.285035
R93 plus.n40 plus.n37 0.285035
R94 plus.n16 plus.n15 0.189894
R95 plus.n17 plus.n16 0.189894
R96 plus.n17 plus.n4 0.189894
R97 plus.n4 plus.n3 0.189894
R98 plus.n24 plus.n1 0.189894
R99 plus.n1 plus.n0 0.189894
R100 plus.n29 plus.n0 0.189894
R101 plus.n59 plus.n30 0.189894
R102 plus.n31 plus.n30 0.189894
R103 plus.n54 plus.n31 0.189894
R104 plus.n34 plus.n33 0.189894
R105 plus.n47 plus.n34 0.189894
R106 plus.n47 plus.n46 0.189894
R107 plus.n46 plus.n45 0.189894
R108 drain_left.n10 drain_left.n8 101.769
R109 drain_left.n6 drain_left.n4 101.769
R110 drain_left.n2 drain_left.n0 101.769
R111 drain_left.n16 drain_left.n15 100.796
R112 drain_left.n14 drain_left.n13 100.796
R113 drain_left.n12 drain_left.n11 100.796
R114 drain_left.n10 drain_left.n9 100.796
R115 drain_left.n7 drain_left.n3 100.796
R116 drain_left.n6 drain_left.n5 100.796
R117 drain_left.n2 drain_left.n1 100.796
R118 drain_left drain_left.n7 27.5844
R119 drain_left.n3 drain_left.t3 9.9005
R120 drain_left.n3 drain_left.t8 9.9005
R121 drain_left.n4 drain_left.t12 9.9005
R122 drain_left.n4 drain_left.t10 9.9005
R123 drain_left.n5 drain_left.t2 9.9005
R124 drain_left.n5 drain_left.t7 9.9005
R125 drain_left.n1 drain_left.t0 9.9005
R126 drain_left.n1 drain_left.t5 9.9005
R127 drain_left.n0 drain_left.t16 9.9005
R128 drain_left.n0 drain_left.t14 9.9005
R129 drain_left.n15 drain_left.t4 9.9005
R130 drain_left.n15 drain_left.t13 9.9005
R131 drain_left.n13 drain_left.t1 9.9005
R132 drain_left.n13 drain_left.t17 9.9005
R133 drain_left.n11 drain_left.t19 9.9005
R134 drain_left.n11 drain_left.t6 9.9005
R135 drain_left.n9 drain_left.t15 9.9005
R136 drain_left.n9 drain_left.t18 9.9005
R137 drain_left.n8 drain_left.t11 9.9005
R138 drain_left.n8 drain_left.t9 9.9005
R139 drain_left drain_left.n16 6.62735
R140 drain_left.n12 drain_left.n10 0.974638
R141 drain_left.n14 drain_left.n12 0.974638
R142 drain_left.n16 drain_left.n14 0.974638
R143 drain_left.n7 drain_left.n6 0.919292
R144 drain_left.n7 drain_left.n2 0.919292
R145 source.n90 source.n88 289.615
R146 source.n74 source.n72 289.615
R147 source.n66 source.n64 289.615
R148 source.n50 source.n48 289.615
R149 source.n2 source.n0 289.615
R150 source.n18 source.n16 289.615
R151 source.n26 source.n24 289.615
R152 source.n42 source.n40 289.615
R153 source.n91 source.n90 185
R154 source.n75 source.n74 185
R155 source.n67 source.n66 185
R156 source.n51 source.n50 185
R157 source.n3 source.n2 185
R158 source.n19 source.n18 185
R159 source.n27 source.n26 185
R160 source.n43 source.n42 185
R161 source.t39 source.n89 167.117
R162 source.t2 source.n73 167.117
R163 source.t19 source.n65 167.117
R164 source.t32 source.n49 167.117
R165 source.t31 source.n1 167.117
R166 source.t18 source.n17 167.117
R167 source.t37 source.n25 167.117
R168 source.t7 source.n41 167.117
R169 source.n9 source.n8 84.1169
R170 source.n11 source.n10 84.1169
R171 source.n13 source.n12 84.1169
R172 source.n15 source.n14 84.1169
R173 source.n33 source.n32 84.1169
R174 source.n35 source.n34 84.1169
R175 source.n37 source.n36 84.1169
R176 source.n39 source.n38 84.1169
R177 source.n87 source.n86 84.1168
R178 source.n85 source.n84 84.1168
R179 source.n83 source.n82 84.1168
R180 source.n81 source.n80 84.1168
R181 source.n63 source.n62 84.1168
R182 source.n61 source.n60 84.1168
R183 source.n59 source.n58 84.1168
R184 source.n57 source.n56 84.1168
R185 source.n90 source.t39 52.3082
R186 source.n74 source.t2 52.3082
R187 source.n66 source.t19 52.3082
R188 source.n50 source.t32 52.3082
R189 source.n2 source.t31 52.3082
R190 source.n18 source.t18 52.3082
R191 source.n26 source.t37 52.3082
R192 source.n42 source.t7 52.3082
R193 source.n95 source.n94 31.4096
R194 source.n79 source.n78 31.4096
R195 source.n71 source.n70 31.4096
R196 source.n55 source.n54 31.4096
R197 source.n7 source.n6 31.4096
R198 source.n23 source.n22 31.4096
R199 source.n31 source.n30 31.4096
R200 source.n47 source.n46 31.4096
R201 source.n55 source.n47 14.6861
R202 source.n86 source.t38 9.9005
R203 source.n86 source.t14 9.9005
R204 source.n84 source.t12 9.9005
R205 source.n84 source.t4 9.9005
R206 source.n82 source.t16 9.9005
R207 source.n82 source.t1 9.9005
R208 source.n80 source.t10 9.9005
R209 source.n80 source.t6 9.9005
R210 source.n62 source.t17 9.9005
R211 source.n62 source.t35 9.9005
R212 source.n60 source.t29 9.9005
R213 source.n60 source.t34 9.9005
R214 source.n58 source.t27 9.9005
R215 source.n58 source.t33 9.9005
R216 source.n56 source.t26 9.9005
R217 source.n56 source.t36 9.9005
R218 source.n8 source.t28 9.9005
R219 source.n8 source.t30 9.9005
R220 source.n10 source.t24 9.9005
R221 source.n10 source.t25 9.9005
R222 source.n12 source.t23 9.9005
R223 source.n12 source.t21 9.9005
R224 source.n14 source.t20 9.9005
R225 source.n14 source.t22 9.9005
R226 source.n32 source.t8 9.9005
R227 source.n32 source.t15 9.9005
R228 source.n34 source.t0 9.9005
R229 source.n34 source.t5 9.9005
R230 source.n36 source.t11 9.9005
R231 source.n36 source.t3 9.9005
R232 source.n38 source.t13 9.9005
R233 source.n38 source.t9 9.9005
R234 source.n91 source.n89 9.71174
R235 source.n75 source.n73 9.71174
R236 source.n67 source.n65 9.71174
R237 source.n51 source.n49 9.71174
R238 source.n3 source.n1 9.71174
R239 source.n19 source.n17 9.71174
R240 source.n27 source.n25 9.71174
R241 source.n43 source.n41 9.71174
R242 source.n94 source.n93 9.45567
R243 source.n78 source.n77 9.45567
R244 source.n70 source.n69 9.45567
R245 source.n54 source.n53 9.45567
R246 source.n6 source.n5 9.45567
R247 source.n22 source.n21 9.45567
R248 source.n30 source.n29 9.45567
R249 source.n46 source.n45 9.45567
R250 source.n93 source.n92 9.3005
R251 source.n77 source.n76 9.3005
R252 source.n69 source.n68 9.3005
R253 source.n53 source.n52 9.3005
R254 source.n5 source.n4 9.3005
R255 source.n21 source.n20 9.3005
R256 source.n29 source.n28 9.3005
R257 source.n45 source.n44 9.3005
R258 source.n96 source.n7 8.93611
R259 source.n94 source.n88 8.14595
R260 source.n78 source.n72 8.14595
R261 source.n70 source.n64 8.14595
R262 source.n54 source.n48 8.14595
R263 source.n6 source.n0 8.14595
R264 source.n22 source.n16 8.14595
R265 source.n30 source.n24 8.14595
R266 source.n46 source.n40 8.14595
R267 source.n92 source.n91 7.3702
R268 source.n76 source.n75 7.3702
R269 source.n68 source.n67 7.3702
R270 source.n52 source.n51 7.3702
R271 source.n4 source.n3 7.3702
R272 source.n20 source.n19 7.3702
R273 source.n28 source.n27 7.3702
R274 source.n44 source.n43 7.3702
R275 source.n92 source.n88 5.81868
R276 source.n76 source.n72 5.81868
R277 source.n68 source.n64 5.81868
R278 source.n52 source.n48 5.81868
R279 source.n4 source.n0 5.81868
R280 source.n20 source.n16 5.81868
R281 source.n28 source.n24 5.81868
R282 source.n44 source.n40 5.81868
R283 source.n96 source.n95 5.7505
R284 source.n93 source.n89 3.44771
R285 source.n77 source.n73 3.44771
R286 source.n69 source.n65 3.44771
R287 source.n53 source.n49 3.44771
R288 source.n5 source.n1 3.44771
R289 source.n21 source.n17 3.44771
R290 source.n29 source.n25 3.44771
R291 source.n45 source.n41 3.44771
R292 source.n47 source.n39 0.974638
R293 source.n39 source.n37 0.974638
R294 source.n37 source.n35 0.974638
R295 source.n35 source.n33 0.974638
R296 source.n33 source.n31 0.974638
R297 source.n23 source.n15 0.974638
R298 source.n15 source.n13 0.974638
R299 source.n13 source.n11 0.974638
R300 source.n11 source.n9 0.974638
R301 source.n9 source.n7 0.974638
R302 source.n57 source.n55 0.974638
R303 source.n59 source.n57 0.974638
R304 source.n61 source.n59 0.974638
R305 source.n63 source.n61 0.974638
R306 source.n71 source.n63 0.974638
R307 source.n81 source.n79 0.974638
R308 source.n83 source.n81 0.974638
R309 source.n85 source.n83 0.974638
R310 source.n87 source.n85 0.974638
R311 source.n95 source.n87 0.974638
R312 source.n31 source.n23 0.470328
R313 source.n79 source.n71 0.470328
R314 source source.n96 0.188
R315 minus.n29 minus.n28 161.3
R316 minus.n27 minus.n0 161.3
R317 minus.n26 minus.n25 161.3
R318 minus.n24 minus.n1 161.3
R319 minus.n20 minus.n19 161.3
R320 minus.n18 minus.n3 161.3
R321 minus.n17 minus.n16 161.3
R322 minus.n15 minus.n4 161.3
R323 minus.n14 minus.n13 161.3
R324 minus.n9 minus.n6 161.3
R325 minus.n59 minus.n58 161.3
R326 minus.n57 minus.n30 161.3
R327 minus.n56 minus.n55 161.3
R328 minus.n54 minus.n31 161.3
R329 minus.n50 minus.n49 161.3
R330 minus.n48 minus.n33 161.3
R331 minus.n47 minus.n46 161.3
R332 minus.n45 minus.n34 161.3
R333 minus.n44 minus.n43 161.3
R334 minus.n39 minus.n36 161.3
R335 minus.n7 minus.t9 131.144
R336 minus.n37 minus.t18 131.144
R337 minus.n8 minus.t7 109.355
R338 minus.n10 minus.t6 109.355
R339 minus.n5 minus.t13 109.355
R340 minus.n15 minus.t15 109.355
R341 minus.n3 minus.t11 109.355
R342 minus.n21 minus.t8 109.355
R343 minus.n22 minus.t17 109.355
R344 minus.n26 minus.t14 109.355
R345 minus.n28 minus.t4 109.355
R346 minus.n38 minus.t0 109.355
R347 minus.n40 minus.t19 109.355
R348 minus.n35 minus.t1 109.355
R349 minus.n45 minus.t10 109.355
R350 minus.n33 minus.t2 109.355
R351 minus.n51 minus.t12 109.355
R352 minus.n52 minus.t3 109.355
R353 minus.n56 minus.t16 109.355
R354 minus.n58 minus.t5 109.355
R355 minus.n23 minus.n22 80.6037
R356 minus.n21 minus.n2 80.6037
R357 minus.n12 minus.n5 80.6037
R358 minus.n11 minus.n10 80.6037
R359 minus.n53 minus.n52 80.6037
R360 minus.n51 minus.n32 80.6037
R361 minus.n42 minus.n35 80.6037
R362 minus.n41 minus.n40 80.6037
R363 minus.n10 minus.n5 48.2005
R364 minus.n22 minus.n21 48.2005
R365 minus.n40 minus.n35 48.2005
R366 minus.n52 minus.n51 48.2005
R367 minus.n7 minus.n6 44.8565
R368 minus.n37 minus.n36 44.8565
R369 minus.n14 minus.n5 43.0884
R370 minus.n21 minus.n20 43.0884
R371 minus.n44 minus.n35 43.0884
R372 minus.n51 minus.n50 43.0884
R373 minus.n10 minus.n9 40.1672
R374 minus.n22 minus.n1 40.1672
R375 minus.n40 minus.n39 40.1672
R376 minus.n52 minus.n31 40.1672
R377 minus.n60 minus.n29 33.8793
R378 minus.n28 minus.n27 27.0217
R379 minus.n58 minus.n57 27.0217
R380 minus.n16 minus.n3 24.1005
R381 minus.n16 minus.n15 24.1005
R382 minus.n46 minus.n45 24.1005
R383 minus.n46 minus.n33 24.1005
R384 minus.n27 minus.n26 21.1793
R385 minus.n57 minus.n56 21.1793
R386 minus.n8 minus.n7 20.1275
R387 minus.n38 minus.n37 20.1275
R388 minus.n9 minus.n8 8.03383
R389 minus.n26 minus.n1 8.03383
R390 minus.n39 minus.n38 8.03383
R391 minus.n56 minus.n31 8.03383
R392 minus.n60 minus.n59 6.70505
R393 minus.n15 minus.n14 5.11262
R394 minus.n20 minus.n3 5.11262
R395 minus.n45 minus.n44 5.11262
R396 minus.n50 minus.n33 5.11262
R397 minus.n23 minus.n2 0.380177
R398 minus.n12 minus.n11 0.380177
R399 minus.n42 minus.n41 0.380177
R400 minus.n53 minus.n32 0.380177
R401 minus.n24 minus.n23 0.285035
R402 minus.n19 minus.n2 0.285035
R403 minus.n13 minus.n12 0.285035
R404 minus.n11 minus.n6 0.285035
R405 minus.n41 minus.n36 0.285035
R406 minus.n43 minus.n42 0.285035
R407 minus.n49 minus.n32 0.285035
R408 minus.n54 minus.n53 0.285035
R409 minus.n29 minus.n0 0.189894
R410 minus.n25 minus.n0 0.189894
R411 minus.n25 minus.n24 0.189894
R412 minus.n19 minus.n18 0.189894
R413 minus.n18 minus.n17 0.189894
R414 minus.n17 minus.n4 0.189894
R415 minus.n13 minus.n4 0.189894
R416 minus.n43 minus.n34 0.189894
R417 minus.n47 minus.n34 0.189894
R418 minus.n48 minus.n47 0.189894
R419 minus.n49 minus.n48 0.189894
R420 minus.n55 minus.n54 0.189894
R421 minus.n55 minus.n30 0.189894
R422 minus.n59 minus.n30 0.189894
R423 minus minus.n60 0.188
R424 drain_right.n10 drain_right.n8 101.769
R425 drain_right.n6 drain_right.n4 101.769
R426 drain_right.n2 drain_right.n0 101.769
R427 drain_right.n10 drain_right.n9 100.796
R428 drain_right.n12 drain_right.n11 100.796
R429 drain_right.n14 drain_right.n13 100.796
R430 drain_right.n16 drain_right.n15 100.796
R431 drain_right.n7 drain_right.n3 100.796
R432 drain_right.n6 drain_right.n5 100.796
R433 drain_right.n2 drain_right.n1 100.796
R434 drain_right drain_right.n7 27.0312
R435 drain_right.n3 drain_right.t9 9.9005
R436 drain_right.n3 drain_right.t17 9.9005
R437 drain_right.n4 drain_right.t3 9.9005
R438 drain_right.n4 drain_right.t14 9.9005
R439 drain_right.n5 drain_right.t7 9.9005
R440 drain_right.n5 drain_right.t16 9.9005
R441 drain_right.n1 drain_right.t0 9.9005
R442 drain_right.n1 drain_right.t18 9.9005
R443 drain_right.n0 drain_right.t1 9.9005
R444 drain_right.n0 drain_right.t19 9.9005
R445 drain_right.n8 drain_right.t12 9.9005
R446 drain_right.n8 drain_right.t10 9.9005
R447 drain_right.n9 drain_right.t6 9.9005
R448 drain_right.n9 drain_right.t13 9.9005
R449 drain_right.n11 drain_right.t8 9.9005
R450 drain_right.n11 drain_right.t4 9.9005
R451 drain_right.n13 drain_right.t2 9.9005
R452 drain_right.n13 drain_right.t11 9.9005
R453 drain_right.n15 drain_right.t15 9.9005
R454 drain_right.n15 drain_right.t5 9.9005
R455 drain_right drain_right.n16 6.62735
R456 drain_right.n16 drain_right.n14 0.974638
R457 drain_right.n14 drain_right.n12 0.974638
R458 drain_right.n12 drain_right.n10 0.974638
R459 drain_right.n7 drain_right.n6 0.919292
R460 drain_right.n7 drain_right.n2 0.919292
C0 source drain_left 7.35231f
C1 source plus 3.6953f
C2 plus drain_left 3.16757f
C3 drain_right source 7.35519f
C4 drain_right drain_left 1.72942f
C5 drain_right plus 0.4852f
C6 source minus 3.68134f
C7 minus drain_left 0.180041f
C8 minus plus 5.29449f
C9 drain_right minus 2.84731f
C10 drain_right a_n3202_n1288# 5.62049f
C11 drain_left a_n3202_n1288# 6.10373f
C12 source a_n3202_n1288# 3.596681f
C13 minus a_n3202_n1288# 12.083856f
C14 plus a_n3202_n1288# 13.466599f
C15 drain_right.t1 a_n3202_n1288# 0.041631f
C16 drain_right.t19 a_n3202_n1288# 0.041631f
C17 drain_right.n0 a_n3202_n1288# 0.265154f
C18 drain_right.t0 a_n3202_n1288# 0.041631f
C19 drain_right.t18 a_n3202_n1288# 0.041631f
C20 drain_right.n1 a_n3202_n1288# 0.26154f
C21 drain_right.n2 a_n3202_n1288# 0.736918f
C22 drain_right.t9 a_n3202_n1288# 0.041631f
C23 drain_right.t17 a_n3202_n1288# 0.041631f
C24 drain_right.n3 a_n3202_n1288# 0.26154f
C25 drain_right.t3 a_n3202_n1288# 0.041631f
C26 drain_right.t14 a_n3202_n1288# 0.041631f
C27 drain_right.n4 a_n3202_n1288# 0.265154f
C28 drain_right.t7 a_n3202_n1288# 0.041631f
C29 drain_right.t16 a_n3202_n1288# 0.041631f
C30 drain_right.n5 a_n3202_n1288# 0.26154f
C31 drain_right.n6 a_n3202_n1288# 0.736918f
C32 drain_right.n7 a_n3202_n1288# 1.37145f
C33 drain_right.t12 a_n3202_n1288# 0.041631f
C34 drain_right.t10 a_n3202_n1288# 0.041631f
C35 drain_right.n8 a_n3202_n1288# 0.265156f
C36 drain_right.t6 a_n3202_n1288# 0.041631f
C37 drain_right.t13 a_n3202_n1288# 0.041631f
C38 drain_right.n9 a_n3202_n1288# 0.261541f
C39 drain_right.n10 a_n3202_n1288# 0.740948f
C40 drain_right.t8 a_n3202_n1288# 0.041631f
C41 drain_right.t4 a_n3202_n1288# 0.041631f
C42 drain_right.n11 a_n3202_n1288# 0.261541f
C43 drain_right.n12 a_n3202_n1288# 0.366976f
C44 drain_right.t2 a_n3202_n1288# 0.041631f
C45 drain_right.t11 a_n3202_n1288# 0.041631f
C46 drain_right.n13 a_n3202_n1288# 0.261541f
C47 drain_right.n14 a_n3202_n1288# 0.366976f
C48 drain_right.t15 a_n3202_n1288# 0.041631f
C49 drain_right.t5 a_n3202_n1288# 0.041631f
C50 drain_right.n15 a_n3202_n1288# 0.261541f
C51 drain_right.n16 a_n3202_n1288# 0.603176f
C52 minus.n0 a_n3202_n1288# 0.040591f
C53 minus.n1 a_n3202_n1288# 0.009211f
C54 minus.t14 a_n3202_n1288# 0.20112f
C55 minus.n2 a_n3202_n1288# 0.06761f
C56 minus.t11 a_n3202_n1288# 0.20112f
C57 minus.n3 a_n3202_n1288# 0.136094f
C58 minus.n4 a_n3202_n1288# 0.040591f
C59 minus.t13 a_n3202_n1288# 0.20112f
C60 minus.n5 a_n3202_n1288# 0.147683f
C61 minus.n6 a_n3202_n1288# 0.18684f
C62 minus.t9 a_n3202_n1288# 0.224109f
C63 minus.n7 a_n3202_n1288# 0.119388f
C64 minus.t7 a_n3202_n1288# 0.20112f
C65 minus.n8 a_n3202_n1288# 0.139506f
C66 minus.n9 a_n3202_n1288# 0.009211f
C67 minus.t6 a_n3202_n1288# 0.20112f
C68 minus.n10 a_n3202_n1288# 0.147182f
C69 minus.n11 a_n3202_n1288# 0.06761f
C70 minus.n12 a_n3202_n1288# 0.06761f
C71 minus.n13 a_n3202_n1288# 0.054164f
C72 minus.n14 a_n3202_n1288# 0.009211f
C73 minus.t15 a_n3202_n1288# 0.20112f
C74 minus.n15 a_n3202_n1288# 0.136094f
C75 minus.n16 a_n3202_n1288# 0.009211f
C76 minus.n17 a_n3202_n1288# 0.040591f
C77 minus.n18 a_n3202_n1288# 0.040591f
C78 minus.n19 a_n3202_n1288# 0.054164f
C79 minus.n20 a_n3202_n1288# 0.009211f
C80 minus.t8 a_n3202_n1288# 0.20112f
C81 minus.n21 a_n3202_n1288# 0.147683f
C82 minus.t17 a_n3202_n1288# 0.20112f
C83 minus.n22 a_n3202_n1288# 0.147182f
C84 minus.n23 a_n3202_n1288# 0.06761f
C85 minus.n24 a_n3202_n1288# 0.054164f
C86 minus.n25 a_n3202_n1288# 0.040591f
C87 minus.n26 a_n3202_n1288# 0.136094f
C88 minus.n27 a_n3202_n1288# 0.009211f
C89 minus.t4 a_n3202_n1288# 0.20112f
C90 minus.n28 a_n3202_n1288# 0.135719f
C91 minus.n29 a_n3202_n1288# 1.29862f
C92 minus.n30 a_n3202_n1288# 0.040591f
C93 minus.n31 a_n3202_n1288# 0.009211f
C94 minus.n32 a_n3202_n1288# 0.06761f
C95 minus.t2 a_n3202_n1288# 0.20112f
C96 minus.n33 a_n3202_n1288# 0.136094f
C97 minus.n34 a_n3202_n1288# 0.040591f
C98 minus.t1 a_n3202_n1288# 0.20112f
C99 minus.n35 a_n3202_n1288# 0.147683f
C100 minus.n36 a_n3202_n1288# 0.18684f
C101 minus.t18 a_n3202_n1288# 0.224109f
C102 minus.n37 a_n3202_n1288# 0.119388f
C103 minus.t0 a_n3202_n1288# 0.20112f
C104 minus.n38 a_n3202_n1288# 0.139506f
C105 minus.n39 a_n3202_n1288# 0.009211f
C106 minus.t19 a_n3202_n1288# 0.20112f
C107 minus.n40 a_n3202_n1288# 0.147182f
C108 minus.n41 a_n3202_n1288# 0.06761f
C109 minus.n42 a_n3202_n1288# 0.06761f
C110 minus.n43 a_n3202_n1288# 0.054164f
C111 minus.n44 a_n3202_n1288# 0.009211f
C112 minus.t10 a_n3202_n1288# 0.20112f
C113 minus.n45 a_n3202_n1288# 0.136094f
C114 minus.n46 a_n3202_n1288# 0.009211f
C115 minus.n47 a_n3202_n1288# 0.040591f
C116 minus.n48 a_n3202_n1288# 0.040591f
C117 minus.n49 a_n3202_n1288# 0.054164f
C118 minus.n50 a_n3202_n1288# 0.009211f
C119 minus.t12 a_n3202_n1288# 0.20112f
C120 minus.n51 a_n3202_n1288# 0.147683f
C121 minus.t3 a_n3202_n1288# 0.20112f
C122 minus.n52 a_n3202_n1288# 0.147182f
C123 minus.n53 a_n3202_n1288# 0.06761f
C124 minus.n54 a_n3202_n1288# 0.054164f
C125 minus.n55 a_n3202_n1288# 0.040591f
C126 minus.t16 a_n3202_n1288# 0.20112f
C127 minus.n56 a_n3202_n1288# 0.136094f
C128 minus.n57 a_n3202_n1288# 0.009211f
C129 minus.t5 a_n3202_n1288# 0.20112f
C130 minus.n58 a_n3202_n1288# 0.135719f
C131 minus.n59 a_n3202_n1288# 0.284798f
C132 minus.n60 a_n3202_n1288# 1.58032f
C133 source.n0 a_n3202_n1288# 0.046198f
C134 source.n1 a_n3202_n1288# 0.102219f
C135 source.t31 a_n3202_n1288# 0.07671f
C136 source.n2 a_n3202_n1288# 0.08f
C137 source.n3 a_n3202_n1288# 0.025789f
C138 source.n4 a_n3202_n1288# 0.017008f
C139 source.n5 a_n3202_n1288# 0.225315f
C140 source.n6 a_n3202_n1288# 0.050644f
C141 source.n7 a_n3202_n1288# 0.555723f
C142 source.t28 a_n3202_n1288# 0.050025f
C143 source.t30 a_n3202_n1288# 0.050025f
C144 source.n8 a_n3202_n1288# 0.26743f
C145 source.n9 a_n3202_n1288# 0.444783f
C146 source.t24 a_n3202_n1288# 0.050025f
C147 source.t25 a_n3202_n1288# 0.050025f
C148 source.n10 a_n3202_n1288# 0.26743f
C149 source.n11 a_n3202_n1288# 0.444783f
C150 source.t23 a_n3202_n1288# 0.050025f
C151 source.t21 a_n3202_n1288# 0.050025f
C152 source.n12 a_n3202_n1288# 0.26743f
C153 source.n13 a_n3202_n1288# 0.444783f
C154 source.t20 a_n3202_n1288# 0.050025f
C155 source.t22 a_n3202_n1288# 0.050025f
C156 source.n14 a_n3202_n1288# 0.26743f
C157 source.n15 a_n3202_n1288# 0.444783f
C158 source.n16 a_n3202_n1288# 0.046198f
C159 source.n17 a_n3202_n1288# 0.102219f
C160 source.t18 a_n3202_n1288# 0.07671f
C161 source.n18 a_n3202_n1288# 0.08f
C162 source.n19 a_n3202_n1288# 0.025789f
C163 source.n20 a_n3202_n1288# 0.017008f
C164 source.n21 a_n3202_n1288# 0.225315f
C165 source.n22 a_n3202_n1288# 0.050644f
C166 source.n23 a_n3202_n1288# 0.173327f
C167 source.n24 a_n3202_n1288# 0.046198f
C168 source.n25 a_n3202_n1288# 0.102219f
C169 source.t37 a_n3202_n1288# 0.07671f
C170 source.n26 a_n3202_n1288# 0.08f
C171 source.n27 a_n3202_n1288# 0.025789f
C172 source.n28 a_n3202_n1288# 0.017008f
C173 source.n29 a_n3202_n1288# 0.225315f
C174 source.n30 a_n3202_n1288# 0.050644f
C175 source.n31 a_n3202_n1288# 0.173327f
C176 source.t8 a_n3202_n1288# 0.050025f
C177 source.t15 a_n3202_n1288# 0.050025f
C178 source.n32 a_n3202_n1288# 0.26743f
C179 source.n33 a_n3202_n1288# 0.444783f
C180 source.t0 a_n3202_n1288# 0.050025f
C181 source.t5 a_n3202_n1288# 0.050025f
C182 source.n34 a_n3202_n1288# 0.26743f
C183 source.n35 a_n3202_n1288# 0.444783f
C184 source.t11 a_n3202_n1288# 0.050025f
C185 source.t3 a_n3202_n1288# 0.050025f
C186 source.n36 a_n3202_n1288# 0.26743f
C187 source.n37 a_n3202_n1288# 0.444783f
C188 source.t13 a_n3202_n1288# 0.050025f
C189 source.t9 a_n3202_n1288# 0.050025f
C190 source.n38 a_n3202_n1288# 0.26743f
C191 source.n39 a_n3202_n1288# 0.444783f
C192 source.n40 a_n3202_n1288# 0.046198f
C193 source.n41 a_n3202_n1288# 0.102219f
C194 source.t7 a_n3202_n1288# 0.07671f
C195 source.n42 a_n3202_n1288# 0.08f
C196 source.n43 a_n3202_n1288# 0.025789f
C197 source.n44 a_n3202_n1288# 0.017008f
C198 source.n45 a_n3202_n1288# 0.225315f
C199 source.n46 a_n3202_n1288# 0.050644f
C200 source.n47 a_n3202_n1288# 0.860907f
C201 source.n48 a_n3202_n1288# 0.046198f
C202 source.n49 a_n3202_n1288# 0.102219f
C203 source.t32 a_n3202_n1288# 0.07671f
C204 source.n50 a_n3202_n1288# 0.08f
C205 source.n51 a_n3202_n1288# 0.025789f
C206 source.n52 a_n3202_n1288# 0.017008f
C207 source.n53 a_n3202_n1288# 0.225315f
C208 source.n54 a_n3202_n1288# 0.050644f
C209 source.n55 a_n3202_n1288# 0.860907f
C210 source.t26 a_n3202_n1288# 0.050025f
C211 source.t36 a_n3202_n1288# 0.050025f
C212 source.n56 a_n3202_n1288# 0.267429f
C213 source.n57 a_n3202_n1288# 0.444785f
C214 source.t27 a_n3202_n1288# 0.050025f
C215 source.t33 a_n3202_n1288# 0.050025f
C216 source.n58 a_n3202_n1288# 0.267429f
C217 source.n59 a_n3202_n1288# 0.444785f
C218 source.t29 a_n3202_n1288# 0.050025f
C219 source.t34 a_n3202_n1288# 0.050025f
C220 source.n60 a_n3202_n1288# 0.267429f
C221 source.n61 a_n3202_n1288# 0.444785f
C222 source.t17 a_n3202_n1288# 0.050025f
C223 source.t35 a_n3202_n1288# 0.050025f
C224 source.n62 a_n3202_n1288# 0.267429f
C225 source.n63 a_n3202_n1288# 0.444785f
C226 source.n64 a_n3202_n1288# 0.046198f
C227 source.n65 a_n3202_n1288# 0.102219f
C228 source.t19 a_n3202_n1288# 0.07671f
C229 source.n66 a_n3202_n1288# 0.08f
C230 source.n67 a_n3202_n1288# 0.025789f
C231 source.n68 a_n3202_n1288# 0.017008f
C232 source.n69 a_n3202_n1288# 0.225315f
C233 source.n70 a_n3202_n1288# 0.050644f
C234 source.n71 a_n3202_n1288# 0.173327f
C235 source.n72 a_n3202_n1288# 0.046198f
C236 source.n73 a_n3202_n1288# 0.102219f
C237 source.t2 a_n3202_n1288# 0.07671f
C238 source.n74 a_n3202_n1288# 0.08f
C239 source.n75 a_n3202_n1288# 0.025789f
C240 source.n76 a_n3202_n1288# 0.017008f
C241 source.n77 a_n3202_n1288# 0.225315f
C242 source.n78 a_n3202_n1288# 0.050644f
C243 source.n79 a_n3202_n1288# 0.173327f
C244 source.t10 a_n3202_n1288# 0.050025f
C245 source.t6 a_n3202_n1288# 0.050025f
C246 source.n80 a_n3202_n1288# 0.267429f
C247 source.n81 a_n3202_n1288# 0.444785f
C248 source.t16 a_n3202_n1288# 0.050025f
C249 source.t1 a_n3202_n1288# 0.050025f
C250 source.n82 a_n3202_n1288# 0.267429f
C251 source.n83 a_n3202_n1288# 0.444785f
C252 source.t12 a_n3202_n1288# 0.050025f
C253 source.t4 a_n3202_n1288# 0.050025f
C254 source.n84 a_n3202_n1288# 0.267429f
C255 source.n85 a_n3202_n1288# 0.444785f
C256 source.t38 a_n3202_n1288# 0.050025f
C257 source.t14 a_n3202_n1288# 0.050025f
C258 source.n86 a_n3202_n1288# 0.267429f
C259 source.n87 a_n3202_n1288# 0.444785f
C260 source.n88 a_n3202_n1288# 0.046198f
C261 source.n89 a_n3202_n1288# 0.102219f
C262 source.t39 a_n3202_n1288# 0.07671f
C263 source.n90 a_n3202_n1288# 0.08f
C264 source.n91 a_n3202_n1288# 0.025789f
C265 source.n92 a_n3202_n1288# 0.017008f
C266 source.n93 a_n3202_n1288# 0.225315f
C267 source.n94 a_n3202_n1288# 0.050644f
C268 source.n95 a_n3202_n1288# 0.386646f
C269 source.n96 a_n3202_n1288# 0.801959f
C270 drain_left.t16 a_n3202_n1288# 0.042831f
C271 drain_left.t14 a_n3202_n1288# 0.042831f
C272 drain_left.n0 a_n3202_n1288# 0.272797f
C273 drain_left.t0 a_n3202_n1288# 0.042831f
C274 drain_left.t5 a_n3202_n1288# 0.042831f
C275 drain_left.n1 a_n3202_n1288# 0.269078f
C276 drain_left.n2 a_n3202_n1288# 0.758157f
C277 drain_left.t3 a_n3202_n1288# 0.042831f
C278 drain_left.t8 a_n3202_n1288# 0.042831f
C279 drain_left.n3 a_n3202_n1288# 0.269078f
C280 drain_left.t12 a_n3202_n1288# 0.042831f
C281 drain_left.t10 a_n3202_n1288# 0.042831f
C282 drain_left.n4 a_n3202_n1288# 0.272797f
C283 drain_left.t2 a_n3202_n1288# 0.042831f
C284 drain_left.t7 a_n3202_n1288# 0.042831f
C285 drain_left.n5 a_n3202_n1288# 0.269078f
C286 drain_left.n6 a_n3202_n1288# 0.758157f
C287 drain_left.n7 a_n3202_n1288# 1.4634f
C288 drain_left.t11 a_n3202_n1288# 0.042831f
C289 drain_left.t9 a_n3202_n1288# 0.042831f
C290 drain_left.n8 a_n3202_n1288# 0.272798f
C291 drain_left.t15 a_n3202_n1288# 0.042831f
C292 drain_left.t18 a_n3202_n1288# 0.042831f
C293 drain_left.n9 a_n3202_n1288# 0.26908f
C294 drain_left.n10 a_n3202_n1288# 0.762304f
C295 drain_left.t19 a_n3202_n1288# 0.042831f
C296 drain_left.t6 a_n3202_n1288# 0.042831f
C297 drain_left.n11 a_n3202_n1288# 0.26908f
C298 drain_left.n12 a_n3202_n1288# 0.377554f
C299 drain_left.t1 a_n3202_n1288# 0.042831f
C300 drain_left.t17 a_n3202_n1288# 0.042831f
C301 drain_left.n13 a_n3202_n1288# 0.26908f
C302 drain_left.n14 a_n3202_n1288# 0.377554f
C303 drain_left.t4 a_n3202_n1288# 0.042831f
C304 drain_left.t13 a_n3202_n1288# 0.042831f
C305 drain_left.n15 a_n3202_n1288# 0.26908f
C306 drain_left.n16 a_n3202_n1288# 0.620561f
C307 plus.n0 a_n3202_n1288# 0.042261f
C308 plus.t5 a_n3202_n1288# 0.209394f
C309 plus.t6 a_n3202_n1288# 0.209394f
C310 plus.n1 a_n3202_n1288# 0.042261f
C311 plus.t8 a_n3202_n1288# 0.209394f
C312 plus.n2 a_n3202_n1288# 0.153237f
C313 plus.n3 a_n3202_n1288# 0.056392f
C314 plus.t11 a_n3202_n1288# 0.209394f
C315 plus.t12 a_n3202_n1288# 0.209394f
C316 plus.n4 a_n3202_n1288# 0.042261f
C317 plus.t15 a_n3202_n1288# 0.209394f
C318 plus.n5 a_n3202_n1288# 0.141693f
C319 plus.n6 a_n3202_n1288# 0.070391f
C320 plus.t13 a_n3202_n1288# 0.209394f
C321 plus.t14 a_n3202_n1288# 0.209394f
C322 plus.n7 a_n3202_n1288# 0.070391f
C323 plus.t16 a_n3202_n1288# 0.209394f
C324 plus.n8 a_n3202_n1288# 0.145245f
C325 plus.t18 a_n3202_n1288# 0.233329f
C326 plus.n9 a_n3202_n1288# 0.1243f
C327 plus.n10 a_n3202_n1288# 0.194527f
C328 plus.n11 a_n3202_n1288# 0.00959f
C329 plus.n12 a_n3202_n1288# 0.153237f
C330 plus.n13 a_n3202_n1288# 0.153758f
C331 plus.n14 a_n3202_n1288# 0.00959f
C332 plus.n15 a_n3202_n1288# 0.056392f
C333 plus.n16 a_n3202_n1288# 0.042261f
C334 plus.n17 a_n3202_n1288# 0.042261f
C335 plus.n18 a_n3202_n1288# 0.00959f
C336 plus.n19 a_n3202_n1288# 0.141693f
C337 plus.n20 a_n3202_n1288# 0.00959f
C338 plus.n21 a_n3202_n1288# 0.153758f
C339 plus.n22 a_n3202_n1288# 0.070391f
C340 plus.n23 a_n3202_n1288# 0.070391f
C341 plus.n24 a_n3202_n1288# 0.056392f
C342 plus.n25 a_n3202_n1288# 0.00959f
C343 plus.n26 a_n3202_n1288# 0.141693f
C344 plus.n27 a_n3202_n1288# 0.00959f
C345 plus.n28 a_n3202_n1288# 0.141302f
C346 plus.n29 a_n3202_n1288# 0.323456f
C347 plus.n30 a_n3202_n1288# 0.042261f
C348 plus.t4 a_n3202_n1288# 0.209394f
C349 plus.n31 a_n3202_n1288# 0.042261f
C350 plus.t10 a_n3202_n1288# 0.209394f
C351 plus.t0 a_n3202_n1288# 0.209394f
C352 plus.n32 a_n3202_n1288# 0.153237f
C353 plus.n33 a_n3202_n1288# 0.056392f
C354 plus.t9 a_n3202_n1288# 0.209394f
C355 plus.n34 a_n3202_n1288# 0.042261f
C356 plus.t3 a_n3202_n1288# 0.209394f
C357 plus.t7 a_n3202_n1288# 0.209394f
C358 plus.n35 a_n3202_n1288# 0.141693f
C359 plus.n36 a_n3202_n1288# 0.070391f
C360 plus.t2 a_n3202_n1288# 0.209394f
C361 plus.n37 a_n3202_n1288# 0.070391f
C362 plus.t19 a_n3202_n1288# 0.209394f
C363 plus.t1 a_n3202_n1288# 0.209394f
C364 plus.n38 a_n3202_n1288# 0.145245f
C365 plus.t17 a_n3202_n1288# 0.233329f
C366 plus.n39 a_n3202_n1288# 0.1243f
C367 plus.n40 a_n3202_n1288# 0.194527f
C368 plus.n41 a_n3202_n1288# 0.00959f
C369 plus.n42 a_n3202_n1288# 0.153237f
C370 plus.n43 a_n3202_n1288# 0.153758f
C371 plus.n44 a_n3202_n1288# 0.00959f
C372 plus.n45 a_n3202_n1288# 0.056392f
C373 plus.n46 a_n3202_n1288# 0.042261f
C374 plus.n47 a_n3202_n1288# 0.042261f
C375 plus.n48 a_n3202_n1288# 0.00959f
C376 plus.n49 a_n3202_n1288# 0.141693f
C377 plus.n50 a_n3202_n1288# 0.00959f
C378 plus.n51 a_n3202_n1288# 0.153758f
C379 plus.n52 a_n3202_n1288# 0.070391f
C380 plus.n53 a_n3202_n1288# 0.070391f
C381 plus.n54 a_n3202_n1288# 0.056392f
C382 plus.n55 a_n3202_n1288# 0.00959f
C383 plus.n56 a_n3202_n1288# 0.141693f
C384 plus.n57 a_n3202_n1288# 0.00959f
C385 plus.n58 a_n3202_n1288# 0.141302f
C386 plus.n59 a_n3202_n1288# 1.28522f
.ends

