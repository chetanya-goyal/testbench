* NGSPICE file created from diffpair355.ext - technology: sky130A

.subckt diffpair355 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t7 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X1 drain_left.t11 plus.t0 source.t11 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 drain_right.t4 minus.t1 source.t22 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X3 a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X4 a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X5 a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X6 source.t6 plus.t1 drain_left.t10 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X7 source.t21 minus.t2 drain_right.t1 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X8 source.t3 plus.t2 drain_left.t9 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X10 source.t4 plus.t3 drain_left.t8 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 source.t7 plus.t4 drain_left.t7 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X12 source.t8 plus.t5 drain_left.t6 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X13 drain_left.t5 plus.t6 source.t0 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X14 drain_right.t0 minus.t3 source.t20 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 drain_right.t2 minus.t4 source.t19 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X16 source.t18 minus.t5 drain_right.t8 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X17 drain_right.t6 minus.t6 source.t17 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X18 drain_right.t5 minus.t7 source.t16 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X19 drain_left.t4 plus.t7 source.t10 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X20 drain_left.t3 plus.t8 source.t2 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X21 source.t1 plus.t9 drain_left.t2 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X22 drain_left.t1 plus.t10 source.t5 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X23 drain_right.t11 minus.t8 source.t15 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X24 source.t14 minus.t9 drain_right.t10 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X25 source.t13 minus.t10 drain_right.t9 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X26 source.t12 minus.t11 drain_right.t3 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X27 drain_left.t0 plus.t11 source.t9 a_n1598_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 minus.n13 minus.t0 874.904
R1 minus.n2 minus.t7 874.904
R2 minus.n28 minus.t6 874.904
R3 minus.n17 minus.t11 874.904
R4 minus.n12 minus.t8 827.433
R5 minus.n10 minus.t5 827.433
R6 minus.n3 minus.t1 827.433
R7 minus.n4 minus.t9 827.433
R8 minus.n27 minus.t2 827.433
R9 minus.n25 minus.t3 827.433
R10 minus.n19 minus.t10 827.433
R11 minus.n18 minus.t4 827.433
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n13 minus.n12 44.549
R31 minus.n4 minus.n2 44.549
R32 minus.n18 minus.n17 44.549
R33 minus.n28 minus.n27 44.549
R34 minus.n30 minus.n14 32.9134
R35 minus.n12 minus.n11 28.4823
R36 minus.n5 minus.n4 28.4823
R37 minus.n20 minus.n18 28.4823
R38 minus.n27 minus.n26 28.4823
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 66.0805
R54 drain_right.n3 drain_right.n2 66.0251
R55 drain_right.n3 drain_right.n0 66.0251
R56 drain_right.n6 drain_right.n5 65.5376
R57 drain_right.n8 drain_right.n7 65.5376
R58 drain_right.n3 drain_right.n1 65.5373
R59 drain_right drain_right.n3 27.2566
R60 drain_right drain_right.n8 6.19632
R61 drain_right.n1 drain_right.t9 2.2005
R62 drain_right.n1 drain_right.t0 2.2005
R63 drain_right.n2 drain_right.t1 2.2005
R64 drain_right.n2 drain_right.t6 2.2005
R65 drain_right.n0 drain_right.t3 2.2005
R66 drain_right.n0 drain_right.t2 2.2005
R67 drain_right.n4 drain_right.t10 2.2005
R68 drain_right.n4 drain_right.t5 2.2005
R69 drain_right.n5 drain_right.t8 2.2005
R70 drain_right.n5 drain_right.t4 2.2005
R71 drain_right.n7 drain_right.t7 2.2005
R72 drain_right.n7 drain_right.t11 2.2005
R73 drain_right.n8 drain_right.n6 0.543603
R74 source.n5 source.t6 51.0588
R75 source.n6 source.t16 51.0588
R76 source.n11 source.t23 51.0588
R77 source.n23 source.t17 51.0586
R78 source.n18 source.t12 51.0586
R79 source.n17 source.t2 51.0586
R80 source.n12 source.t8 51.0586
R81 source.n0 source.t10 51.0586
R82 source.n2 source.n1 48.8588
R83 source.n4 source.n3 48.8588
R84 source.n8 source.n7 48.8588
R85 source.n10 source.n9 48.8588
R86 source.n22 source.n21 48.8586
R87 source.n20 source.n19 48.8586
R88 source.n16 source.n15 48.8586
R89 source.n14 source.n13 48.8586
R90 source.n12 source.n11 19.5581
R91 source.n24 source.n0 14.0236
R92 source.n24 source.n23 5.53498
R93 source.n21 source.t20 2.2005
R94 source.n21 source.t21 2.2005
R95 source.n19 source.t19 2.2005
R96 source.n19 source.t13 2.2005
R97 source.n15 source.t5 2.2005
R98 source.n15 source.t3 2.2005
R99 source.n13 source.t11 2.2005
R100 source.n13 source.t7 2.2005
R101 source.n1 source.t9 2.2005
R102 source.n1 source.t4 2.2005
R103 source.n3 source.t0 2.2005
R104 source.n3 source.t1 2.2005
R105 source.n7 source.t22 2.2005
R106 source.n7 source.t14 2.2005
R107 source.n9 source.t15 2.2005
R108 source.n9 source.t18 2.2005
R109 source.n11 source.n10 0.543603
R110 source.n10 source.n8 0.543603
R111 source.n8 source.n6 0.543603
R112 source.n5 source.n4 0.543603
R113 source.n4 source.n2 0.543603
R114 source.n2 source.n0 0.543603
R115 source.n14 source.n12 0.543603
R116 source.n16 source.n14 0.543603
R117 source.n17 source.n16 0.543603
R118 source.n20 source.n18 0.543603
R119 source.n22 source.n20 0.543603
R120 source.n23 source.n22 0.543603
R121 source.n6 source.n5 0.470328
R122 source.n18 source.n17 0.470328
R123 source source.n24 0.188
R124 plus.n2 plus.t1 874.904
R125 plus.n13 plus.t7 874.904
R126 plus.n17 plus.t8 874.904
R127 plus.n28 plus.t5 874.904
R128 plus.n3 plus.t6 827.433
R129 plus.n4 plus.t9 827.433
R130 plus.n10 plus.t11 827.433
R131 plus.n12 plus.t3 827.433
R132 plus.n19 plus.t2 827.433
R133 plus.n18 plus.t10 827.433
R134 plus.n25 plus.t4 827.433
R135 plus.n27 plus.t0 827.433
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 63.5369
R151 plus.n11 plus.n10 63.5369
R152 plus.n26 plus.n25 63.5369
R153 plus.n20 plus.n18 63.5369
R154 plus.n3 plus.n2 44.549
R155 plus.n13 plus.n12 44.549
R156 plus.n28 plus.n27 44.549
R157 plus.n19 plus.n17 44.549
R158 plus.n5 plus.n3 28.4823
R159 plus.n12 plus.n11 28.4823
R160 plus.n27 plus.n26 28.4823
R161 plus.n20 plus.n19 28.4823
R162 plus plus.n29 27.9308
R163 plus plus.n14 11.0194
R164 plus.n4 plus.n1 9.49444
R165 plus.n10 plus.n9 9.49444
R166 plus.n25 plus.n24 9.49444
R167 plus.n18 plus.n16 9.49444
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 66.0807
R177 drain_left.n3 drain_left.n2 66.0251
R178 drain_left.n3 drain_left.n0 66.0251
R179 drain_left.n6 drain_left.n5 65.5376
R180 drain_left.n8 drain_left.n7 65.5374
R181 drain_left.n3 drain_left.n1 65.5373
R182 drain_left drain_left.n3 27.8099
R183 drain_left drain_left.n8 6.19632
R184 drain_left.n1 drain_left.t7 2.2005
R185 drain_left.n1 drain_left.t1 2.2005
R186 drain_left.n2 drain_left.t9 2.2005
R187 drain_left.n2 drain_left.t3 2.2005
R188 drain_left.n0 drain_left.t6 2.2005
R189 drain_left.n0 drain_left.t11 2.2005
R190 drain_left.n7 drain_left.t8 2.2005
R191 drain_left.n7 drain_left.t4 2.2005
R192 drain_left.n5 drain_left.t2 2.2005
R193 drain_left.n5 drain_left.t0 2.2005
R194 drain_left.n4 drain_left.t10 2.2005
R195 drain_left.n4 drain_left.t5 2.2005
R196 drain_left.n8 drain_left.n6 0.543603
C0 source minus 3.33482f
C1 source plus 3.34886f
C2 drain_right drain_left 0.785787f
C3 minus drain_left 0.170859f
C4 plus drain_left 3.73938f
C5 minus drain_right 3.58592f
C6 plus drain_right 0.30725f
C7 source drain_left 18.2222f
C8 minus plus 4.58797f
C9 source drain_right 18.221899f
C10 drain_right a_n1598_n2688# 5.48901f
C11 drain_left a_n1598_n2688# 5.73511f
C12 source a_n1598_n2688# 6.994413f
C13 minus a_n1598_n2688# 5.997251f
C14 plus a_n1598_n2688# 7.756259f
C15 drain_left.t6 a_n1598_n2688# 0.236453f
C16 drain_left.t11 a_n1598_n2688# 0.236453f
C17 drain_left.n0 a_n1598_n2688# 2.07107f
C18 drain_left.t7 a_n1598_n2688# 0.236453f
C19 drain_left.t1 a_n1598_n2688# 0.236453f
C20 drain_left.n1 a_n1598_n2688# 2.06818f
C21 drain_left.t9 a_n1598_n2688# 0.236453f
C22 drain_left.t3 a_n1598_n2688# 0.236453f
C23 drain_left.n2 a_n1598_n2688# 2.07107f
C24 drain_left.n3 a_n1598_n2688# 2.42471f
C25 drain_left.t10 a_n1598_n2688# 0.236453f
C26 drain_left.t5 a_n1598_n2688# 0.236453f
C27 drain_left.n4 a_n1598_n2688# 2.07144f
C28 drain_left.t2 a_n1598_n2688# 0.236453f
C29 drain_left.t0 a_n1598_n2688# 0.236453f
C30 drain_left.n5 a_n1598_n2688# 2.06818f
C31 drain_left.n6 a_n1598_n2688# 0.775475f
C32 drain_left.t8 a_n1598_n2688# 0.236453f
C33 drain_left.t4 a_n1598_n2688# 0.236453f
C34 drain_left.n7 a_n1598_n2688# 2.06817f
C35 drain_left.n8 a_n1598_n2688# 0.659411f
C36 plus.n0 a_n1598_n2688# 0.053066f
C37 plus.t3 a_n1598_n2688# 0.405997f
C38 plus.t11 a_n1598_n2688# 0.405997f
C39 plus.n1 a_n1598_n2688# 0.01973f
C40 plus.t1 a_n1598_n2688# 0.415417f
C41 plus.n2 a_n1598_n2688# 0.186143f
C42 plus.t6 a_n1598_n2688# 0.405997f
C43 plus.n3 a_n1598_n2688# 0.169537f
C44 plus.t9 a_n1598_n2688# 0.405997f
C45 plus.n4 a_n1598_n2688# 0.169537f
C46 plus.n5 a_n1598_n2688# 0.021857f
C47 plus.n6 a_n1598_n2688# 0.120776f
C48 plus.n7 a_n1598_n2688# 0.053066f
C49 plus.n8 a_n1598_n2688# 0.053066f
C50 plus.n9 a_n1598_n2688# 0.01973f
C51 plus.n10 a_n1598_n2688# 0.169537f
C52 plus.n11 a_n1598_n2688# 0.021857f
C53 plus.n12 a_n1598_n2688# 0.169537f
C54 plus.t7 a_n1598_n2688# 0.415417f
C55 plus.n13 a_n1598_n2688# 0.186063f
C56 plus.n14 a_n1598_n2688# 0.522796f
C57 plus.n15 a_n1598_n2688# 0.053066f
C58 plus.t5 a_n1598_n2688# 0.415417f
C59 plus.t0 a_n1598_n2688# 0.405997f
C60 plus.t4 a_n1598_n2688# 0.405997f
C61 plus.n16 a_n1598_n2688# 0.01973f
C62 plus.t8 a_n1598_n2688# 0.415417f
C63 plus.n17 a_n1598_n2688# 0.186143f
C64 plus.t10 a_n1598_n2688# 0.405997f
C65 plus.n18 a_n1598_n2688# 0.169537f
C66 plus.t2 a_n1598_n2688# 0.405997f
C67 plus.n19 a_n1598_n2688# 0.169537f
C68 plus.n20 a_n1598_n2688# 0.021857f
C69 plus.n21 a_n1598_n2688# 0.120776f
C70 plus.n22 a_n1598_n2688# 0.053066f
C71 plus.n23 a_n1598_n2688# 0.053066f
C72 plus.n24 a_n1598_n2688# 0.01973f
C73 plus.n25 a_n1598_n2688# 0.169537f
C74 plus.n26 a_n1598_n2688# 0.021857f
C75 plus.n27 a_n1598_n2688# 0.169537f
C76 plus.n28 a_n1598_n2688# 0.186063f
C77 plus.n29 a_n1598_n2688# 1.40464f
C78 source.t10 a_n1598_n2688# 2.04196f
C79 source.n0 a_n1598_n2688# 1.17418f
C80 source.t9 a_n1598_n2688# 0.191491f
C81 source.t4 a_n1598_n2688# 0.191491f
C82 source.n1 a_n1598_n2688# 1.60304f
C83 source.n2 a_n1598_n2688# 0.345181f
C84 source.t0 a_n1598_n2688# 0.191491f
C85 source.t1 a_n1598_n2688# 0.191491f
C86 source.n3 a_n1598_n2688# 1.60304f
C87 source.n4 a_n1598_n2688# 0.345181f
C88 source.t6 a_n1598_n2688# 2.04197f
C89 source.n5 a_n1598_n2688# 0.422147f
C90 source.t16 a_n1598_n2688# 2.04197f
C91 source.n6 a_n1598_n2688# 0.422147f
C92 source.t22 a_n1598_n2688# 0.191491f
C93 source.t14 a_n1598_n2688# 0.191491f
C94 source.n7 a_n1598_n2688# 1.60304f
C95 source.n8 a_n1598_n2688# 0.345181f
C96 source.t15 a_n1598_n2688# 0.191491f
C97 source.t18 a_n1598_n2688# 0.191491f
C98 source.n9 a_n1598_n2688# 1.60304f
C99 source.n10 a_n1598_n2688# 0.345181f
C100 source.t23 a_n1598_n2688# 2.04197f
C101 source.n11 a_n1598_n2688# 1.5654f
C102 source.t8 a_n1598_n2688# 2.04196f
C103 source.n12 a_n1598_n2688# 1.5654f
C104 source.t11 a_n1598_n2688# 0.191491f
C105 source.t7 a_n1598_n2688# 0.191491f
C106 source.n13 a_n1598_n2688# 1.60304f
C107 source.n14 a_n1598_n2688# 0.345186f
C108 source.t5 a_n1598_n2688# 0.191491f
C109 source.t3 a_n1598_n2688# 0.191491f
C110 source.n15 a_n1598_n2688# 1.60304f
C111 source.n16 a_n1598_n2688# 0.345186f
C112 source.t2 a_n1598_n2688# 2.04196f
C113 source.n17 a_n1598_n2688# 0.422152f
C114 source.t12 a_n1598_n2688# 2.04196f
C115 source.n18 a_n1598_n2688# 0.422152f
C116 source.t19 a_n1598_n2688# 0.191491f
C117 source.t13 a_n1598_n2688# 0.191491f
C118 source.n19 a_n1598_n2688# 1.60304f
C119 source.n20 a_n1598_n2688# 0.345186f
C120 source.t20 a_n1598_n2688# 0.191491f
C121 source.t21 a_n1598_n2688# 0.191491f
C122 source.n21 a_n1598_n2688# 1.60304f
C123 source.n22 a_n1598_n2688# 0.345186f
C124 source.t17 a_n1598_n2688# 2.04196f
C125 source.n23 a_n1598_n2688# 0.574143f
C126 source.n24 a_n1598_n2688# 1.40163f
C127 drain_right.t3 a_n1598_n2688# 0.23678f
C128 drain_right.t2 a_n1598_n2688# 0.23678f
C129 drain_right.n0 a_n1598_n2688# 2.07393f
C130 drain_right.t9 a_n1598_n2688# 0.23678f
C131 drain_right.t0 a_n1598_n2688# 0.23678f
C132 drain_right.n1 a_n1598_n2688# 2.07103f
C133 drain_right.t1 a_n1598_n2688# 0.23678f
C134 drain_right.t6 a_n1598_n2688# 0.23678f
C135 drain_right.n2 a_n1598_n2688# 2.07393f
C136 drain_right.n3 a_n1598_n2688# 2.35922f
C137 drain_right.t10 a_n1598_n2688# 0.23678f
C138 drain_right.t5 a_n1598_n2688# 0.23678f
C139 drain_right.n4 a_n1598_n2688# 2.07429f
C140 drain_right.t8 a_n1598_n2688# 0.23678f
C141 drain_right.t4 a_n1598_n2688# 0.23678f
C142 drain_right.n5 a_n1598_n2688# 2.07104f
C143 drain_right.n6 a_n1598_n2688# 0.776555f
C144 drain_right.t7 a_n1598_n2688# 0.23678f
C145 drain_right.t11 a_n1598_n2688# 0.23678f
C146 drain_right.n7 a_n1598_n2688# 2.07104f
C147 drain_right.n8 a_n1598_n2688# 0.660313f
C148 minus.n0 a_n1598_n2688# 0.052127f
C149 minus.t0 a_n1598_n2688# 0.408061f
C150 minus.t8 a_n1598_n2688# 0.398807f
C151 minus.t5 a_n1598_n2688# 0.398807f
C152 minus.n1 a_n1598_n2688# 0.019381f
C153 minus.t7 a_n1598_n2688# 0.408061f
C154 minus.n2 a_n1598_n2688# 0.182847f
C155 minus.t1 a_n1598_n2688# 0.398807f
C156 minus.n3 a_n1598_n2688# 0.166535f
C157 minus.t9 a_n1598_n2688# 0.398807f
C158 minus.n4 a_n1598_n2688# 0.166535f
C159 minus.n5 a_n1598_n2688# 0.02147f
C160 minus.n6 a_n1598_n2688# 0.118637f
C161 minus.n7 a_n1598_n2688# 0.052127f
C162 minus.n8 a_n1598_n2688# 0.052127f
C163 minus.n9 a_n1598_n2688# 0.019381f
C164 minus.n10 a_n1598_n2688# 0.166535f
C165 minus.n11 a_n1598_n2688# 0.02147f
C166 minus.n12 a_n1598_n2688# 0.166535f
C167 minus.n13 a_n1598_n2688# 0.182769f
C168 minus.n14 a_n1598_n2688# 1.5834f
C169 minus.n15 a_n1598_n2688# 0.052127f
C170 minus.t2 a_n1598_n2688# 0.398807f
C171 minus.t3 a_n1598_n2688# 0.398807f
C172 minus.n16 a_n1598_n2688# 0.019381f
C173 minus.t11 a_n1598_n2688# 0.408061f
C174 minus.n17 a_n1598_n2688# 0.182847f
C175 minus.t4 a_n1598_n2688# 0.398807f
C176 minus.n18 a_n1598_n2688# 0.166535f
C177 minus.t10 a_n1598_n2688# 0.398807f
C178 minus.n19 a_n1598_n2688# 0.166535f
C179 minus.n20 a_n1598_n2688# 0.02147f
C180 minus.n21 a_n1598_n2688# 0.118637f
C181 minus.n22 a_n1598_n2688# 0.052127f
C182 minus.n23 a_n1598_n2688# 0.052127f
C183 minus.n24 a_n1598_n2688# 0.019381f
C184 minus.n25 a_n1598_n2688# 0.166535f
C185 minus.n26 a_n1598_n2688# 0.02147f
C186 minus.n27 a_n1598_n2688# 0.166535f
C187 minus.t6 a_n1598_n2688# 0.408061f
C188 minus.n28 a_n1598_n2688# 0.182769f
C189 minus.n29 a_n1598_n2688# 0.342247f
C190 minus.n30 a_n1598_n2688# 1.94048f
.ends

