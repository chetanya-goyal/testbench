* NGSPICE file created from diffpair546.ext - technology: sky130A

.subckt diffpair546 minus drain_right drain_left source plus
X0 a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X1 drain_left.t13 plus.t0 source.t15 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X2 drain_right.t13 minus.t0 source.t5 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X3 drain_left.t12 plus.t1 source.t21 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X4 source.t23 plus.t2 drain_left.t11 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 drain_left.t10 plus.t3 source.t22 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X6 source.t7 minus.t1 drain_right.t12 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X7 source.t0 minus.t2 drain_right.t11 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X8 drain_left.t9 plus.t4 source.t20 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X9 drain_left.t8 plus.t5 source.t18 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X10 drain_right.t10 minus.t3 source.t10 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X11 source.t16 plus.t6 drain_left.t7 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X12 drain_left.t6 plus.t7 source.t14 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X13 drain_right.t9 minus.t4 source.t2 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X14 a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X15 source.t1 minus.t5 drain_right.t8 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X16 drain_right.t7 minus.t6 source.t4 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X17 drain_right.t6 minus.t7 source.t9 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X18 drain_right.t5 minus.t8 source.t12 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X19 source.t17 plus.t8 drain_left.t5 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X20 source.t24 plus.t9 drain_left.t4 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X21 drain_right.t4 minus.t9 source.t11 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X22 a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X23 source.t19 plus.t10 drain_left.t3 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X24 drain_left.t2 plus.t11 source.t27 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X25 source.t26 plus.t12 drain_left.t1 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X26 a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X27 drain_left.t0 plus.t13 source.t25 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X28 source.t3 minus.t10 drain_right.t3 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X29 source.t6 minus.t11 drain_right.t2 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X30 drain_right.t1 minus.t12 source.t8 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X31 source.t13 minus.t13 drain_right.t0 a_n2364_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
R0 plus.n5 plus.t5 596.394
R1 plus.n27 plus.t1 596.394
R2 plus.n20 plus.t0 572.548
R3 plus.n18 plus.t9 572.548
R4 plus.n2 plus.t4 572.548
R5 plus.n12 plus.t8 572.548
R6 plus.n4 plus.t3 572.548
R7 plus.n6 plus.t12 572.548
R8 plus.n42 plus.t7 572.548
R9 plus.n40 plus.t6 572.548
R10 plus.n24 plus.t11 572.548
R11 plus.n34 plus.t10 572.548
R12 plus.n26 plus.t13 572.548
R13 plus.n28 plus.t2 572.548
R14 plus.n8 plus.n7 161.3
R15 plus.n9 plus.n4 161.3
R16 plus.n11 plus.n10 161.3
R17 plus.n12 plus.n3 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n15 plus.n2 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n18 plus.n1 161.3
R22 plus.n19 plus.n0 161.3
R23 plus.n21 plus.n20 161.3
R24 plus.n30 plus.n29 161.3
R25 plus.n31 plus.n26 161.3
R26 plus.n33 plus.n32 161.3
R27 plus.n34 plus.n25 161.3
R28 plus.n36 plus.n35 161.3
R29 plus.n37 plus.n24 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n40 plus.n23 161.3
R32 plus.n41 plus.n22 161.3
R33 plus.n43 plus.n42 161.3
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus plus.n43 33.2433
R39 plus.n18 plus.n17 30.6732
R40 plus.n7 plus.n6 30.6732
R41 plus.n40 plus.n39 30.6732
R42 plus.n29 plus.n28 30.6732
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus plus.n21 13.4304
R58 plus.n19 plus.n18 13.146
R59 plus.n41 plus.n40 13.146
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n7 source.t11 45.521
R79 source.n27 source.t8 45.5208
R80 source.n20 source.t21 45.5208
R81 source.n0 source.t15 45.5208
R82 source.n2 source.n1 44.201
R83 source.n4 source.n3 44.201
R84 source.n6 source.n5 44.201
R85 source.n9 source.n8 44.201
R86 source.n11 source.n10 44.201
R87 source.n13 source.n12 44.201
R88 source.n26 source.n25 44.2008
R89 source.n24 source.n23 44.2008
R90 source.n22 source.n21 44.2008
R91 source.n19 source.n18 44.2008
R92 source.n17 source.n16 44.2008
R93 source.n15 source.n14 44.2008
R94 source.n15 source.n13 25.3363
R95 source.n28 source.n0 18.7415
R96 source.n28 source.n27 5.7074
R97 source.n25 source.t10 1.3205
R98 source.n25 source.t13 1.3205
R99 source.n23 source.t5 1.3205
R100 source.n23 source.t0 1.3205
R101 source.n21 source.t2 1.3205
R102 source.n21 source.t1 1.3205
R103 source.n18 source.t25 1.3205
R104 source.n18 source.t23 1.3205
R105 source.n16 source.t27 1.3205
R106 source.n16 source.t19 1.3205
R107 source.n14 source.t14 1.3205
R108 source.n14 source.t16 1.3205
R109 source.n1 source.t20 1.3205
R110 source.n1 source.t24 1.3205
R111 source.n3 source.t22 1.3205
R112 source.n3 source.t17 1.3205
R113 source.n5 source.t18 1.3205
R114 source.n5 source.t26 1.3205
R115 source.n8 source.t12 1.3205
R116 source.n8 source.t7 1.3205
R117 source.n10 source.t9 1.3205
R118 source.n10 source.t3 1.3205
R119 source.n12 source.t4 1.3205
R120 source.n12 source.t6 1.3205
R121 source.n7 source.n6 0.914293
R122 source.n22 source.n20 0.914293
R123 source.n13 source.n11 0.888431
R124 source.n11 source.n9 0.888431
R125 source.n9 source.n7 0.888431
R126 source.n6 source.n4 0.888431
R127 source.n4 source.n2 0.888431
R128 source.n2 source.n0 0.888431
R129 source.n17 source.n15 0.888431
R130 source.n19 source.n17 0.888431
R131 source.n20 source.n19 0.888431
R132 source.n24 source.n22 0.888431
R133 source.n26 source.n24 0.888431
R134 source.n27 source.n26 0.888431
R135 source source.n28 0.188
R136 drain_left.n7 drain_left.t8 63.0877
R137 drain_left.n1 drain_left.t6 63.0875
R138 drain_left.n4 drain_left.n2 61.7675
R139 drain_left.n9 drain_left.n8 60.8798
R140 drain_left.n7 drain_left.n6 60.8798
R141 drain_left.n11 drain_left.n10 60.8796
R142 drain_left.n4 drain_left.n3 60.8796
R143 drain_left.n1 drain_left.n0 60.8796
R144 drain_left drain_left.n5 34.7454
R145 drain_left drain_left.n11 6.54115
R146 drain_left.n2 drain_left.t11 1.3205
R147 drain_left.n2 drain_left.t12 1.3205
R148 drain_left.n3 drain_left.t3 1.3205
R149 drain_left.n3 drain_left.t0 1.3205
R150 drain_left.n0 drain_left.t7 1.3205
R151 drain_left.n0 drain_left.t2 1.3205
R152 drain_left.n10 drain_left.t4 1.3205
R153 drain_left.n10 drain_left.t13 1.3205
R154 drain_left.n8 drain_left.t5 1.3205
R155 drain_left.n8 drain_left.t9 1.3205
R156 drain_left.n6 drain_left.t1 1.3205
R157 drain_left.n6 drain_left.t10 1.3205
R158 drain_left.n9 drain_left.n7 0.888431
R159 drain_left.n11 drain_left.n9 0.888431
R160 drain_left.n5 drain_left.n1 0.611102
R161 drain_left.n5 drain_left.n4 0.167137
R162 minus.n5 minus.t9 596.394
R163 minus.n27 minus.t4 596.394
R164 minus.n6 minus.t1 572.548
R165 minus.n8 minus.t8 572.548
R166 minus.n12 minus.t10 572.548
R167 minus.n14 minus.t7 572.548
R168 minus.n18 minus.t11 572.548
R169 minus.n20 minus.t6 572.548
R170 minus.n28 minus.t5 572.548
R171 minus.n30 minus.t0 572.548
R172 minus.n34 minus.t2 572.548
R173 minus.n36 minus.t3 572.548
R174 minus.n40 minus.t13 572.548
R175 minus.n42 minus.t12 572.548
R176 minus.n21 minus.n20 161.3
R177 minus.n19 minus.n0 161.3
R178 minus.n18 minus.n17 161.3
R179 minus.n16 minus.n1 161.3
R180 minus.n15 minus.n14 161.3
R181 minus.n13 minus.n2 161.3
R182 minus.n12 minus.n11 161.3
R183 minus.n10 minus.n3 161.3
R184 minus.n9 minus.n8 161.3
R185 minus.n7 minus.n4 161.3
R186 minus.n43 minus.n42 161.3
R187 minus.n41 minus.n22 161.3
R188 minus.n40 minus.n39 161.3
R189 minus.n38 minus.n23 161.3
R190 minus.n37 minus.n36 161.3
R191 minus.n35 minus.n24 161.3
R192 minus.n34 minus.n33 161.3
R193 minus.n32 minus.n25 161.3
R194 minus.n31 minus.n30 161.3
R195 minus.n29 minus.n26 161.3
R196 minus.n5 minus.n4 44.9119
R197 minus.n27 minus.n26 44.9119
R198 minus.n44 minus.n21 40.4986
R199 minus.n20 minus.n19 35.055
R200 minus.n42 minus.n41 35.055
R201 minus.n7 minus.n6 30.6732
R202 minus.n18 minus.n1 30.6732
R203 minus.n29 minus.n28 30.6732
R204 minus.n40 minus.n23 30.6732
R205 minus.n8 minus.n3 26.2914
R206 minus.n14 minus.n13 26.2914
R207 minus.n30 minus.n25 26.2914
R208 minus.n36 minus.n35 26.2914
R209 minus.n12 minus.n3 21.9096
R210 minus.n13 minus.n12 21.9096
R211 minus.n34 minus.n25 21.9096
R212 minus.n35 minus.n34 21.9096
R213 minus.n6 minus.n5 17.739
R214 minus.n28 minus.n27 17.739
R215 minus.n8 minus.n7 17.5278
R216 minus.n14 minus.n1 17.5278
R217 minus.n30 minus.n29 17.5278
R218 minus.n36 minus.n23 17.5278
R219 minus.n19 minus.n18 13.146
R220 minus.n41 minus.n40 13.146
R221 minus.n44 minus.n43 6.65012
R222 minus.n21 minus.n0 0.189894
R223 minus.n17 minus.n0 0.189894
R224 minus.n17 minus.n16 0.189894
R225 minus.n16 minus.n15 0.189894
R226 minus.n15 minus.n2 0.189894
R227 minus.n11 minus.n2 0.189894
R228 minus.n11 minus.n10 0.189894
R229 minus.n10 minus.n9 0.189894
R230 minus.n9 minus.n4 0.189894
R231 minus.n31 minus.n26 0.189894
R232 minus.n32 minus.n31 0.189894
R233 minus.n33 minus.n32 0.189894
R234 minus.n33 minus.n24 0.189894
R235 minus.n37 minus.n24 0.189894
R236 minus.n38 minus.n37 0.189894
R237 minus.n39 minus.n38 0.189894
R238 minus.n39 minus.n22 0.189894
R239 minus.n43 minus.n22 0.189894
R240 minus minus.n44 0.188
R241 drain_right.n1 drain_right.t9 63.0875
R242 drain_right.n11 drain_right.t7 62.1998
R243 drain_right.n8 drain_right.n6 61.7676
R244 drain_right.n4 drain_right.n2 61.7675
R245 drain_right.n8 drain_right.n7 60.8798
R246 drain_right.n10 drain_right.n9 60.8798
R247 drain_right.n4 drain_right.n3 60.8796
R248 drain_right.n1 drain_right.n0 60.8796
R249 drain_right drain_right.n5 34.1922
R250 drain_right drain_right.n11 6.09718
R251 drain_right.n2 drain_right.t0 1.3205
R252 drain_right.n2 drain_right.t1 1.3205
R253 drain_right.n3 drain_right.t11 1.3205
R254 drain_right.n3 drain_right.t10 1.3205
R255 drain_right.n0 drain_right.t8 1.3205
R256 drain_right.n0 drain_right.t13 1.3205
R257 drain_right.n6 drain_right.t12 1.3205
R258 drain_right.n6 drain_right.t4 1.3205
R259 drain_right.n7 drain_right.t3 1.3205
R260 drain_right.n7 drain_right.t5 1.3205
R261 drain_right.n9 drain_right.t2 1.3205
R262 drain_right.n9 drain_right.t6 1.3205
R263 drain_right.n11 drain_right.n10 0.888431
R264 drain_right.n10 drain_right.n8 0.888431
R265 drain_right.n5 drain_right.n1 0.611102
R266 drain_right.n5 drain_right.n4 0.167137
C0 minus drain_right 11.197599f
C1 minus source 11.0425f
C2 drain_left drain_right 1.23484f
C3 drain_left source 22.501999f
C4 plus minus 6.64803f
C5 drain_right source 22.493801f
C6 drain_left plus 11.4278f
C7 drain_left minus 0.172675f
C8 plus drain_right 0.391476f
C9 plus source 11.0572f
C10 drain_right a_n2364_n3888# 8.38399f
C11 drain_left a_n2364_n3888# 8.73299f
C12 source a_n2364_n3888# 7.762824f
C13 minus a_n2364_n3888# 9.584849f
C14 plus a_n2364_n3888# 11.46142f
C15 drain_right.t9 a_n2364_n3888# 3.41588f
C16 drain_right.t8 a_n2364_n3888# 0.295633f
C17 drain_right.t13 a_n2364_n3888# 0.295633f
C18 drain_right.n0 a_n2364_n3888# 2.67218f
C19 drain_right.n1 a_n2364_n3888# 0.673913f
C20 drain_right.t0 a_n2364_n3888# 0.295633f
C21 drain_right.t1 a_n2364_n3888# 0.295633f
C22 drain_right.n2 a_n2364_n3888# 2.67731f
C23 drain_right.t11 a_n2364_n3888# 0.295633f
C24 drain_right.t10 a_n2364_n3888# 0.295633f
C25 drain_right.n3 a_n2364_n3888# 2.67218f
C26 drain_right.n4 a_n2364_n3888# 0.644408f
C27 drain_right.n5 a_n2364_n3888# 1.50396f
C28 drain_right.t12 a_n2364_n3888# 0.295633f
C29 drain_right.t4 a_n2364_n3888# 0.295633f
C30 drain_right.n6 a_n2364_n3888# 2.67731f
C31 drain_right.t3 a_n2364_n3888# 0.295633f
C32 drain_right.t5 a_n2364_n3888# 0.295633f
C33 drain_right.n7 a_n2364_n3888# 2.67218f
C34 drain_right.n8 a_n2364_n3888# 0.698909f
C35 drain_right.t2 a_n2364_n3888# 0.295633f
C36 drain_right.t6 a_n2364_n3888# 0.295633f
C37 drain_right.n9 a_n2364_n3888# 2.67218f
C38 drain_right.n10 a_n2364_n3888# 0.346994f
C39 drain_right.t7 a_n2364_n3888# 3.41091f
C40 drain_right.n11 a_n2364_n3888# 0.582446f
C41 minus.n0 a_n2364_n3888# 0.040796f
C42 minus.n1 a_n2364_n3888# 0.009258f
C43 minus.t11 a_n2364_n3888# 1.21728f
C44 minus.n2 a_n2364_n3888# 0.040796f
C45 minus.n3 a_n2364_n3888# 0.009258f
C46 minus.t10 a_n2364_n3888# 1.21728f
C47 minus.n4 a_n2364_n3888# 0.171893f
C48 minus.t9 a_n2364_n3888# 1.23606f
C49 minus.n5 a_n2364_n3888# 0.454512f
C50 minus.t1 a_n2364_n3888# 1.21728f
C51 minus.n6 a_n2364_n3888# 0.474805f
C52 minus.n7 a_n2364_n3888# 0.009258f
C53 minus.t8 a_n2364_n3888# 1.21728f
C54 minus.n8 a_n2364_n3888# 0.469751f
C55 minus.n9 a_n2364_n3888# 0.040796f
C56 minus.n10 a_n2364_n3888# 0.040796f
C57 minus.n11 a_n2364_n3888# 0.040796f
C58 minus.n12 a_n2364_n3888# 0.469751f
C59 minus.n13 a_n2364_n3888# 0.009258f
C60 minus.t7 a_n2364_n3888# 1.21728f
C61 minus.n14 a_n2364_n3888# 0.469751f
C62 minus.n15 a_n2364_n3888# 0.040796f
C63 minus.n16 a_n2364_n3888# 0.040796f
C64 minus.n17 a_n2364_n3888# 0.040796f
C65 minus.n18 a_n2364_n3888# 0.469751f
C66 minus.n19 a_n2364_n3888# 0.009258f
C67 minus.t6 a_n2364_n3888# 1.21728f
C68 minus.n20 a_n2364_n3888# 0.468242f
C69 minus.n21 a_n2364_n3888# 1.71602f
C70 minus.n22 a_n2364_n3888# 0.040796f
C71 minus.n23 a_n2364_n3888# 0.009258f
C72 minus.n24 a_n2364_n3888# 0.040796f
C73 minus.n25 a_n2364_n3888# 0.009258f
C74 minus.n26 a_n2364_n3888# 0.171893f
C75 minus.t4 a_n2364_n3888# 1.23606f
C76 minus.n27 a_n2364_n3888# 0.454512f
C77 minus.t5 a_n2364_n3888# 1.21728f
C78 minus.n28 a_n2364_n3888# 0.474805f
C79 minus.n29 a_n2364_n3888# 0.009258f
C80 minus.t0 a_n2364_n3888# 1.21728f
C81 minus.n30 a_n2364_n3888# 0.469751f
C82 minus.n31 a_n2364_n3888# 0.040796f
C83 minus.n32 a_n2364_n3888# 0.040796f
C84 minus.n33 a_n2364_n3888# 0.040796f
C85 minus.t2 a_n2364_n3888# 1.21728f
C86 minus.n34 a_n2364_n3888# 0.469751f
C87 minus.n35 a_n2364_n3888# 0.009258f
C88 minus.t3 a_n2364_n3888# 1.21728f
C89 minus.n36 a_n2364_n3888# 0.469751f
C90 minus.n37 a_n2364_n3888# 0.040796f
C91 minus.n38 a_n2364_n3888# 0.040796f
C92 minus.n39 a_n2364_n3888# 0.040796f
C93 minus.t13 a_n2364_n3888# 1.21728f
C94 minus.n40 a_n2364_n3888# 0.469751f
C95 minus.n41 a_n2364_n3888# 0.009258f
C96 minus.t12 a_n2364_n3888# 1.21728f
C97 minus.n42 a_n2364_n3888# 0.468242f
C98 minus.n43 a_n2364_n3888# 0.281044f
C99 minus.n44 a_n2364_n3888# 2.05445f
C100 drain_left.t6 a_n2364_n3888# 3.42623f
C101 drain_left.t7 a_n2364_n3888# 0.296529f
C102 drain_left.t2 a_n2364_n3888# 0.296529f
C103 drain_left.n0 a_n2364_n3888# 2.68028f
C104 drain_left.n1 a_n2364_n3888# 0.675956f
C105 drain_left.t11 a_n2364_n3888# 0.296529f
C106 drain_left.t12 a_n2364_n3888# 0.296529f
C107 drain_left.n2 a_n2364_n3888# 2.68543f
C108 drain_left.t3 a_n2364_n3888# 0.296529f
C109 drain_left.t0 a_n2364_n3888# 0.296529f
C110 drain_left.n3 a_n2364_n3888# 2.68028f
C111 drain_left.n4 a_n2364_n3888# 0.646361f
C112 drain_left.n5 a_n2364_n3888# 1.56016f
C113 drain_left.t8 a_n2364_n3888# 3.42623f
C114 drain_left.t1 a_n2364_n3888# 0.296529f
C115 drain_left.t10 a_n2364_n3888# 0.296529f
C116 drain_left.n6 a_n2364_n3888# 2.68028f
C117 drain_left.n7 a_n2364_n3888# 0.697356f
C118 drain_left.t5 a_n2364_n3888# 0.296529f
C119 drain_left.t9 a_n2364_n3888# 0.296529f
C120 drain_left.n8 a_n2364_n3888# 2.68028f
C121 drain_left.n9 a_n2364_n3888# 0.348045f
C122 drain_left.t4 a_n2364_n3888# 0.296529f
C123 drain_left.t13 a_n2364_n3888# 0.296529f
C124 drain_left.n10 a_n2364_n3888# 2.68027f
C125 drain_left.n11 a_n2364_n3888# 0.569325f
C126 source.t15 a_n2364_n3888# 3.45195f
C127 source.n0 a_n2364_n3888# 1.64542f
C128 source.t20 a_n2364_n3888# 0.308028f
C129 source.t24 a_n2364_n3888# 0.308028f
C130 source.n1 a_n2364_n3888# 2.70577f
C131 source.n2 a_n2364_n3888# 0.404669f
C132 source.t22 a_n2364_n3888# 0.308028f
C133 source.t17 a_n2364_n3888# 0.308028f
C134 source.n3 a_n2364_n3888# 2.70577f
C135 source.n4 a_n2364_n3888# 0.404669f
C136 source.t18 a_n2364_n3888# 0.308028f
C137 source.t26 a_n2364_n3888# 0.308028f
C138 source.n5 a_n2364_n3888# 2.70577f
C139 source.n6 a_n2364_n3888# 0.406834f
C140 source.t11 a_n2364_n3888# 3.45195f
C141 source.n7 a_n2364_n3888# 0.500724f
C142 source.t12 a_n2364_n3888# 0.308028f
C143 source.t7 a_n2364_n3888# 0.308028f
C144 source.n8 a_n2364_n3888# 2.70577f
C145 source.n9 a_n2364_n3888# 0.404669f
C146 source.t9 a_n2364_n3888# 0.308028f
C147 source.t3 a_n2364_n3888# 0.308028f
C148 source.n10 a_n2364_n3888# 2.70577f
C149 source.n11 a_n2364_n3888# 0.404669f
C150 source.t4 a_n2364_n3888# 0.308028f
C151 source.t6 a_n2364_n3888# 0.308028f
C152 source.n12 a_n2364_n3888# 2.70577f
C153 source.n13 a_n2364_n3888# 2.06913f
C154 source.t14 a_n2364_n3888# 0.308028f
C155 source.t16 a_n2364_n3888# 0.308028f
C156 source.n14 a_n2364_n3888# 2.70576f
C157 source.n15 a_n2364_n3888# 2.06913f
C158 source.t27 a_n2364_n3888# 0.308028f
C159 source.t19 a_n2364_n3888# 0.308028f
C160 source.n16 a_n2364_n3888# 2.70576f
C161 source.n17 a_n2364_n3888# 0.404672f
C162 source.t25 a_n2364_n3888# 0.308028f
C163 source.t23 a_n2364_n3888# 0.308028f
C164 source.n18 a_n2364_n3888# 2.70576f
C165 source.n19 a_n2364_n3888# 0.404672f
C166 source.t21 a_n2364_n3888# 3.45195f
C167 source.n20 a_n2364_n3888# 0.500728f
C168 source.t2 a_n2364_n3888# 0.308028f
C169 source.t1 a_n2364_n3888# 0.308028f
C170 source.n21 a_n2364_n3888# 2.70576f
C171 source.n22 a_n2364_n3888# 0.406838f
C172 source.t5 a_n2364_n3888# 0.308028f
C173 source.t0 a_n2364_n3888# 0.308028f
C174 source.n23 a_n2364_n3888# 2.70576f
C175 source.n24 a_n2364_n3888# 0.404672f
C176 source.t10 a_n2364_n3888# 0.308028f
C177 source.t13 a_n2364_n3888# 0.308028f
C178 source.n25 a_n2364_n3888# 2.70576f
C179 source.n26 a_n2364_n3888# 0.404672f
C180 source.t8 a_n2364_n3888# 3.45195f
C181 source.n27 a_n2364_n3888# 0.633063f
C182 source.n28 a_n2364_n3888# 1.91735f
C183 plus.n0 a_n2364_n3888# 0.04134f
C184 plus.t0 a_n2364_n3888# 1.23349f
C185 plus.t9 a_n2364_n3888# 1.23349f
C186 plus.n1 a_n2364_n3888# 0.04134f
C187 plus.t4 a_n2364_n3888# 1.23349f
C188 plus.n2 a_n2364_n3888# 0.476008f
C189 plus.n3 a_n2364_n3888# 0.04134f
C190 plus.t8 a_n2364_n3888# 1.23349f
C191 plus.t3 a_n2364_n3888# 1.23349f
C192 plus.n4 a_n2364_n3888# 0.476008f
C193 plus.t5 a_n2364_n3888# 1.25253f
C194 plus.n5 a_n2364_n3888# 0.460566f
C195 plus.t12 a_n2364_n3888# 1.23349f
C196 plus.n6 a_n2364_n3888# 0.481129f
C197 plus.n7 a_n2364_n3888# 0.009381f
C198 plus.n8 a_n2364_n3888# 0.174183f
C199 plus.n9 a_n2364_n3888# 0.04134f
C200 plus.n10 a_n2364_n3888# 0.04134f
C201 plus.n11 a_n2364_n3888# 0.009381f
C202 plus.n12 a_n2364_n3888# 0.476008f
C203 plus.n13 a_n2364_n3888# 0.009381f
C204 plus.n14 a_n2364_n3888# 0.04134f
C205 plus.n15 a_n2364_n3888# 0.04134f
C206 plus.n16 a_n2364_n3888# 0.04134f
C207 plus.n17 a_n2364_n3888# 0.009381f
C208 plus.n18 a_n2364_n3888# 0.476008f
C209 plus.n19 a_n2364_n3888# 0.009381f
C210 plus.n20 a_n2364_n3888# 0.474479f
C211 plus.n21 a_n2364_n3888# 0.536974f
C212 plus.n22 a_n2364_n3888# 0.04134f
C213 plus.t7 a_n2364_n3888# 1.23349f
C214 plus.n23 a_n2364_n3888# 0.04134f
C215 plus.t6 a_n2364_n3888# 1.23349f
C216 plus.t11 a_n2364_n3888# 1.23349f
C217 plus.n24 a_n2364_n3888# 0.476008f
C218 plus.n25 a_n2364_n3888# 0.04134f
C219 plus.t10 a_n2364_n3888# 1.23349f
C220 plus.t13 a_n2364_n3888# 1.23349f
C221 plus.n26 a_n2364_n3888# 0.476008f
C222 plus.t1 a_n2364_n3888# 1.25253f
C223 plus.n27 a_n2364_n3888# 0.460566f
C224 plus.t2 a_n2364_n3888# 1.23349f
C225 plus.n28 a_n2364_n3888# 0.481129f
C226 plus.n29 a_n2364_n3888# 0.009381f
C227 plus.n30 a_n2364_n3888# 0.174183f
C228 plus.n31 a_n2364_n3888# 0.04134f
C229 plus.n32 a_n2364_n3888# 0.04134f
C230 plus.n33 a_n2364_n3888# 0.009381f
C231 plus.n34 a_n2364_n3888# 0.476008f
C232 plus.n35 a_n2364_n3888# 0.009381f
C233 plus.n36 a_n2364_n3888# 0.04134f
C234 plus.n37 a_n2364_n3888# 0.04134f
C235 plus.n38 a_n2364_n3888# 0.04134f
C236 plus.n39 a_n2364_n3888# 0.009381f
C237 plus.n40 a_n2364_n3888# 0.476008f
C238 plus.n41 a_n2364_n3888# 0.009381f
C239 plus.n42 a_n2364_n3888# 0.474479f
C240 plus.n43 a_n2364_n3888# 1.44157f
.ends

