* NGSPICE file created from diffpair105.ext - technology: sky130A

.subckt diffpair105 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t18 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_left.t10 plus.t1 source.t13 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t9 plus.t2 source.t11 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t12 plus.t3 drain_left.t8 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X4 source.t4 minus.t0 drain_right.t11 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X5 source.t5 minus.t1 drain_right.t10 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X7 source.t14 plus.t4 drain_left.t7 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X8 source.t10 plus.t5 drain_left.t6 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X9 drain_right.t9 minus.t2 source.t8 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X10 source.t3 minus.t3 drain_right.t8 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X11 drain_right.t7 minus.t4 source.t6 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X13 source.t7 minus.t5 drain_right.t6 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X14 source.t15 plus.t6 drain_left.t5 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X15 source.t19 plus.t7 drain_left.t4 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X16 a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X17 source.t0 minus.t6 drain_right.t5 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X18 source.t1 minus.t7 drain_right.t4 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X19 drain_right.t3 minus.t8 source.t2 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X20 drain_right.t2 minus.t9 source.t9 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X21 drain_right.t1 minus.t10 source.t22 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X22 source.t20 plus.t8 drain_left.t3 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X23 drain_right.t0 minus.t11 source.t23 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X24 a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X25 drain_left.t2 plus.t9 source.t21 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X26 drain_left.t1 plus.t10 source.t16 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X27 drain_left.t0 plus.t11 source.t17 a_n1528_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
R0 plus.n2 plus.t5 347.332
R1 plus.n13 plus.t11 347.332
R2 plus.n17 plus.t10 347.332
R3 plus.n28 plus.t3 347.332
R4 plus.n3 plus.t1 318.12
R5 plus.n4 plus.t7 318.12
R6 plus.n10 plus.t0 318.12
R7 plus.n12 plus.t6 318.12
R8 plus.n19 plus.t8 318.12
R9 plus.n18 plus.t2 318.12
R10 plus.n25 plus.t4 318.12
R11 plus.n27 plus.t9 318.12
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 24.9384
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 8.29217
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n74 source.n72 289.615
R53 source.n62 source.n60 289.615
R54 source.n54 source.n52 289.615
R55 source.n42 source.n40 289.615
R56 source.n2 source.n0 289.615
R57 source.n14 source.n12 289.615
R58 source.n22 source.n20 289.615
R59 source.n34 source.n32 289.615
R60 source.n75 source.n74 185
R61 source.n63 source.n62 185
R62 source.n55 source.n54 185
R63 source.n43 source.n42 185
R64 source.n3 source.n2 185
R65 source.n15 source.n14 185
R66 source.n23 source.n22 185
R67 source.n35 source.n34 185
R68 source.t22 source.n73 167.117
R69 source.t1 source.n61 167.117
R70 source.t16 source.n53 167.117
R71 source.t12 source.n41 167.117
R72 source.t17 source.n1 167.117
R73 source.t10 source.n13 167.117
R74 source.t9 source.n21 167.117
R75 source.t3 source.n33 167.117
R76 source.n9 source.n8 84.1169
R77 source.n11 source.n10 84.1169
R78 source.n29 source.n28 84.1169
R79 source.n31 source.n30 84.1169
R80 source.n71 source.n70 84.1168
R81 source.n69 source.n68 84.1168
R82 source.n51 source.n50 84.1168
R83 source.n49 source.n48 84.1168
R84 source.n74 source.t22 52.3082
R85 source.n62 source.t1 52.3082
R86 source.n54 source.t16 52.3082
R87 source.n42 source.t12 52.3082
R88 source.n2 source.t17 52.3082
R89 source.n14 source.t10 52.3082
R90 source.n22 source.t9 52.3082
R91 source.n34 source.t3 52.3082
R92 source.n79 source.n78 31.4096
R93 source.n67 source.n66 31.4096
R94 source.n59 source.n58 31.4096
R95 source.n47 source.n46 31.4096
R96 source.n7 source.n6 31.4096
R97 source.n19 source.n18 31.4096
R98 source.n27 source.n26 31.4096
R99 source.n39 source.n38 31.4096
R100 source.n47 source.n39 14.212
R101 source.n70 source.t6 9.9005
R102 source.n70 source.t0 9.9005
R103 source.n68 source.t8 9.9005
R104 source.n68 source.t7 9.9005
R105 source.n50 source.t11 9.9005
R106 source.n50 source.t20 9.9005
R107 source.n48 source.t21 9.9005
R108 source.n48 source.t14 9.9005
R109 source.n8 source.t18 9.9005
R110 source.n8 source.t15 9.9005
R111 source.n10 source.t13 9.9005
R112 source.n10 source.t19 9.9005
R113 source.n28 source.t2 9.9005
R114 source.n28 source.t5 9.9005
R115 source.n30 source.t23 9.9005
R116 source.n30 source.t4 9.9005
R117 source.n75 source.n73 9.71174
R118 source.n63 source.n61 9.71174
R119 source.n55 source.n53 9.71174
R120 source.n43 source.n41 9.71174
R121 source.n3 source.n1 9.71174
R122 source.n15 source.n13 9.71174
R123 source.n23 source.n21 9.71174
R124 source.n35 source.n33 9.71174
R125 source.n78 source.n77 9.45567
R126 source.n66 source.n65 9.45567
R127 source.n58 source.n57 9.45567
R128 source.n46 source.n45 9.45567
R129 source.n6 source.n5 9.45567
R130 source.n18 source.n17 9.45567
R131 source.n26 source.n25 9.45567
R132 source.n38 source.n37 9.45567
R133 source.n77 source.n76 9.3005
R134 source.n65 source.n64 9.3005
R135 source.n57 source.n56 9.3005
R136 source.n45 source.n44 9.3005
R137 source.n5 source.n4 9.3005
R138 source.n17 source.n16 9.3005
R139 source.n25 source.n24 9.3005
R140 source.n37 source.n36 9.3005
R141 source.n80 source.n7 8.69904
R142 source.n78 source.n72 8.14595
R143 source.n66 source.n60 8.14595
R144 source.n58 source.n52 8.14595
R145 source.n46 source.n40 8.14595
R146 source.n6 source.n0 8.14595
R147 source.n18 source.n12 8.14595
R148 source.n26 source.n20 8.14595
R149 source.n38 source.n32 8.14595
R150 source.n76 source.n75 7.3702
R151 source.n64 source.n63 7.3702
R152 source.n56 source.n55 7.3702
R153 source.n44 source.n43 7.3702
R154 source.n4 source.n3 7.3702
R155 source.n16 source.n15 7.3702
R156 source.n24 source.n23 7.3702
R157 source.n36 source.n35 7.3702
R158 source.n76 source.n72 5.81868
R159 source.n64 source.n60 5.81868
R160 source.n56 source.n52 5.81868
R161 source.n44 source.n40 5.81868
R162 source.n4 source.n0 5.81868
R163 source.n16 source.n12 5.81868
R164 source.n24 source.n20 5.81868
R165 source.n36 source.n32 5.81868
R166 source.n80 source.n79 5.51343
R167 source.n77 source.n73 3.44771
R168 source.n65 source.n61 3.44771
R169 source.n57 source.n53 3.44771
R170 source.n45 source.n41 3.44771
R171 source.n5 source.n1 3.44771
R172 source.n17 source.n13 3.44771
R173 source.n25 source.n21 3.44771
R174 source.n37 source.n33 3.44771
R175 source.n39 source.n31 0.5005
R176 source.n31 source.n29 0.5005
R177 source.n29 source.n27 0.5005
R178 source.n19 source.n11 0.5005
R179 source.n11 source.n9 0.5005
R180 source.n9 source.n7 0.5005
R181 source.n49 source.n47 0.5005
R182 source.n51 source.n49 0.5005
R183 source.n59 source.n51 0.5005
R184 source.n69 source.n67 0.5005
R185 source.n71 source.n69 0.5005
R186 source.n79 source.n71 0.5005
R187 source.n27 source.n19 0.470328
R188 source.n67 source.n59 0.470328
R189 source source.n80 0.188
R190 drain_left.n6 drain_left.n4 101.296
R191 drain_left.n3 drain_left.n2 101.24
R192 drain_left.n3 drain_left.n0 101.24
R193 drain_left.n8 drain_left.n7 100.796
R194 drain_left.n6 drain_left.n5 100.796
R195 drain_left.n3 drain_left.n1 100.796
R196 drain_left drain_left.n3 22.2913
R197 drain_left.n1 drain_left.t7 9.9005
R198 drain_left.n1 drain_left.t9 9.9005
R199 drain_left.n2 drain_left.t3 9.9005
R200 drain_left.n2 drain_left.t1 9.9005
R201 drain_left.n0 drain_left.t8 9.9005
R202 drain_left.n0 drain_left.t2 9.9005
R203 drain_left.n7 drain_left.t5 9.9005
R204 drain_left.n7 drain_left.t0 9.9005
R205 drain_left.n5 drain_left.t4 9.9005
R206 drain_left.n5 drain_left.t11 9.9005
R207 drain_left.n4 drain_left.t6 9.9005
R208 drain_left.n4 drain_left.t10 9.9005
R209 drain_left drain_left.n8 6.15322
R210 drain_left.n8 drain_left.n6 0.5005
R211 minus.n13 minus.t3 347.332
R212 minus.n2 minus.t9 347.332
R213 minus.n28 minus.t10 347.332
R214 minus.n17 minus.t7 347.332
R215 minus.n12 minus.t11 318.12
R216 minus.n10 minus.t0 318.12
R217 minus.n3 minus.t8 318.12
R218 minus.n4 minus.t1 318.12
R219 minus.n27 minus.t6 318.12
R220 minus.n25 minus.t4 318.12
R221 minus.n19 minus.t5 318.12
R222 minus.n18 minus.t2 318.12
R223 minus.n6 minus.n2 161.489
R224 minus.n21 minus.n17 161.489
R225 minus.n14 minus.n13 161.3
R226 minus.n11 minus.n0 161.3
R227 minus.n9 minus.n8 161.3
R228 minus.n7 minus.n1 161.3
R229 minus.n6 minus.n5 161.3
R230 minus.n29 minus.n28 161.3
R231 minus.n26 minus.n15 161.3
R232 minus.n24 minus.n23 161.3
R233 minus.n22 minus.n16 161.3
R234 minus.n21 minus.n20 161.3
R235 minus.n9 minus.n1 73.0308
R236 minus.n24 minus.n16 73.0308
R237 minus.n11 minus.n10 67.1884
R238 minus.n5 minus.n3 67.1884
R239 minus.n20 minus.n19 67.1884
R240 minus.n26 minus.n25 67.1884
R241 minus.n13 minus.n12 55.5035
R242 minus.n4 minus.n2 55.5035
R243 minus.n18 minus.n17 55.5035
R244 minus.n28 minus.n27 55.5035
R245 minus.n30 minus.n14 27.2694
R246 minus.n12 minus.n11 17.5278
R247 minus.n5 minus.n4 17.5278
R248 minus.n20 minus.n18 17.5278
R249 minus.n27 minus.n26 17.5278
R250 minus.n30 minus.n29 6.43611
R251 minus.n10 minus.n9 5.84292
R252 minus.n3 minus.n1 5.84292
R253 minus.n19 minus.n16 5.84292
R254 minus.n25 minus.n24 5.84292
R255 minus.n14 minus.n0 0.189894
R256 minus.n8 minus.n0 0.189894
R257 minus.n8 minus.n7 0.189894
R258 minus.n7 minus.n6 0.189894
R259 minus.n22 minus.n21 0.189894
R260 minus.n23 minus.n22 0.189894
R261 minus.n23 minus.n15 0.189894
R262 minus.n29 minus.n15 0.189894
R263 minus minus.n30 0.188
R264 drain_right.n6 drain_right.n4 101.296
R265 drain_right.n3 drain_right.n2 101.24
R266 drain_right.n3 drain_right.n0 101.24
R267 drain_right.n6 drain_right.n5 100.796
R268 drain_right.n8 drain_right.n7 100.796
R269 drain_right.n3 drain_right.n1 100.796
R270 drain_right drain_right.n3 21.7381
R271 drain_right.n1 drain_right.t6 9.9005
R272 drain_right.n1 drain_right.t7 9.9005
R273 drain_right.n2 drain_right.t5 9.9005
R274 drain_right.n2 drain_right.t1 9.9005
R275 drain_right.n0 drain_right.t4 9.9005
R276 drain_right.n0 drain_right.t9 9.9005
R277 drain_right.n4 drain_right.t10 9.9005
R278 drain_right.n4 drain_right.t2 9.9005
R279 drain_right.n5 drain_right.t11 9.9005
R280 drain_right.n5 drain_right.t3 9.9005
R281 drain_right.n7 drain_right.t8 9.9005
R282 drain_right.n7 drain_right.t0 9.9005
R283 drain_right drain_right.n8 6.15322
R284 drain_right.n8 drain_right.n6 0.5005
C0 drain_right plus 0.306604f
C1 source minus 1.14245f
C2 source drain_left 6.15348f
C3 minus drain_left 0.176852f
C4 source plus 1.15642f
C5 minus plus 3.21812f
C6 drain_left plus 1.1825f
C7 drain_right source 6.15293f
C8 drain_right minus 1.03636f
C9 drain_right drain_left 0.751334f
C10 drain_right a_n1528_n1288# 3.5352f
C11 drain_left a_n1528_n1288# 3.74583f
C12 source a_n1528_n1288# 2.977508f
C13 minus a_n1528_n1288# 5.128845f
C14 plus a_n1528_n1288# 5.786765f
C15 drain_right.t4 a_n1528_n1288# 0.043518f
C16 drain_right.t9 a_n1528_n1288# 0.043518f
C17 drain_right.n0 a_n1528_n1288# 0.274743f
C18 drain_right.t6 a_n1528_n1288# 0.043518f
C19 drain_right.t7 a_n1528_n1288# 0.043518f
C20 drain_right.n1 a_n1528_n1288# 0.273394f
C21 drain_right.t5 a_n1528_n1288# 0.043518f
C22 drain_right.t1 a_n1528_n1288# 0.043518f
C23 drain_right.n2 a_n1528_n1288# 0.274743f
C24 drain_right.n3 a_n1528_n1288# 1.51237f
C25 drain_right.t10 a_n1528_n1288# 0.043518f
C26 drain_right.t2 a_n1528_n1288# 0.043518f
C27 drain_right.n4 a_n1528_n1288# 0.274928f
C28 drain_right.t11 a_n1528_n1288# 0.043518f
C29 drain_right.t3 a_n1528_n1288# 0.043518f
C30 drain_right.n5 a_n1528_n1288# 0.273395f
C31 drain_right.n6 a_n1528_n1288# 0.608505f
C32 drain_right.t8 a_n1528_n1288# 0.043518f
C33 drain_right.t0 a_n1528_n1288# 0.043518f
C34 drain_right.n7 a_n1528_n1288# 0.273395f
C35 drain_right.n8 a_n1528_n1288# 0.526757f
C36 minus.n0 a_n1528_n1288# 0.031576f
C37 minus.t3 a_n1528_n1288# 0.049241f
C38 minus.t11 a_n1528_n1288# 0.046457f
C39 minus.t0 a_n1528_n1288# 0.046457f
C40 minus.n1 a_n1528_n1288# 0.011253f
C41 minus.t9 a_n1528_n1288# 0.049241f
C42 minus.n2 a_n1528_n1288# 0.042384f
C43 minus.t8 a_n1528_n1288# 0.046457f
C44 minus.n3 a_n1528_n1288# 0.034069f
C45 minus.t1 a_n1528_n1288# 0.046457f
C46 minus.n4 a_n1528_n1288# 0.034069f
C47 minus.n5 a_n1528_n1288# 0.012032f
C48 minus.n6 a_n1528_n1288# 0.066031f
C49 minus.n7 a_n1528_n1288# 0.031576f
C50 minus.n8 a_n1528_n1288# 0.031576f
C51 minus.n9 a_n1528_n1288# 0.011253f
C52 minus.n10 a_n1528_n1288# 0.034069f
C53 minus.n11 a_n1528_n1288# 0.012032f
C54 minus.n12 a_n1528_n1288# 0.034069f
C55 minus.n13 a_n1528_n1288# 0.042344f
C56 minus.n14 a_n1528_n1288# 0.692958f
C57 minus.n15 a_n1528_n1288# 0.031576f
C58 minus.t6 a_n1528_n1288# 0.046457f
C59 minus.t4 a_n1528_n1288# 0.046457f
C60 minus.n16 a_n1528_n1288# 0.011253f
C61 minus.t7 a_n1528_n1288# 0.049241f
C62 minus.n17 a_n1528_n1288# 0.042384f
C63 minus.t2 a_n1528_n1288# 0.046457f
C64 minus.n18 a_n1528_n1288# 0.034069f
C65 minus.t5 a_n1528_n1288# 0.046457f
C66 minus.n19 a_n1528_n1288# 0.034069f
C67 minus.n20 a_n1528_n1288# 0.012032f
C68 minus.n21 a_n1528_n1288# 0.066031f
C69 minus.n22 a_n1528_n1288# 0.031576f
C70 minus.n23 a_n1528_n1288# 0.031576f
C71 minus.n24 a_n1528_n1288# 0.011253f
C72 minus.n25 a_n1528_n1288# 0.034069f
C73 minus.n26 a_n1528_n1288# 0.012032f
C74 minus.n27 a_n1528_n1288# 0.034069f
C75 minus.t10 a_n1528_n1288# 0.049241f
C76 minus.n28 a_n1528_n1288# 0.042344f
C77 minus.n29 a_n1528_n1288# 0.201667f
C78 minus.n30 a_n1528_n1288# 0.859355f
C79 drain_left.t8 a_n1528_n1288# 0.042775f
C80 drain_left.t2 a_n1528_n1288# 0.042775f
C81 drain_left.n0 a_n1528_n1288# 0.270051f
C82 drain_left.t7 a_n1528_n1288# 0.042775f
C83 drain_left.t9 a_n1528_n1288# 0.042775f
C84 drain_left.n1 a_n1528_n1288# 0.268725f
C85 drain_left.t3 a_n1528_n1288# 0.042775f
C86 drain_left.t1 a_n1528_n1288# 0.042775f
C87 drain_left.n2 a_n1528_n1288# 0.270051f
C88 drain_left.n3 a_n1528_n1288# 1.53974f
C89 drain_left.t6 a_n1528_n1288# 0.042775f
C90 drain_left.t10 a_n1528_n1288# 0.042775f
C91 drain_left.n4 a_n1528_n1288# 0.270233f
C92 drain_left.t4 a_n1528_n1288# 0.042775f
C93 drain_left.t11 a_n1528_n1288# 0.042775f
C94 drain_left.n5 a_n1528_n1288# 0.268726f
C95 drain_left.n6 a_n1528_n1288# 0.598114f
C96 drain_left.t5 a_n1528_n1288# 0.042775f
C97 drain_left.t0 a_n1528_n1288# 0.042775f
C98 drain_left.n7 a_n1528_n1288# 0.268726f
C99 drain_left.n8 a_n1528_n1288# 0.517761f
C100 source.n0 a_n1528_n1288# 0.039926f
C101 source.n1 a_n1528_n1288# 0.088341f
C102 source.t17 a_n1528_n1288# 0.066296f
C103 source.n2 a_n1528_n1288# 0.069139f
C104 source.n3 a_n1528_n1288# 0.022288f
C105 source.n4 a_n1528_n1288# 0.014699f
C106 source.n5 a_n1528_n1288# 0.194726f
C107 source.n6 a_n1528_n1288# 0.043768f
C108 source.n7 a_n1528_n1288# 0.406259f
C109 source.t18 a_n1528_n1288# 0.043233f
C110 source.t15 a_n1528_n1288# 0.043233f
C111 source.n8 a_n1528_n1288# 0.231124f
C112 source.n9 a_n1528_n1288# 0.300814f
C113 source.t13 a_n1528_n1288# 0.043233f
C114 source.t19 a_n1528_n1288# 0.043233f
C115 source.n10 a_n1528_n1288# 0.231124f
C116 source.n11 a_n1528_n1288# 0.300814f
C117 source.n12 a_n1528_n1288# 0.039926f
C118 source.n13 a_n1528_n1288# 0.088341f
C119 source.t10 a_n1528_n1288# 0.066296f
C120 source.n14 a_n1528_n1288# 0.069139f
C121 source.n15 a_n1528_n1288# 0.022288f
C122 source.n16 a_n1528_n1288# 0.014699f
C123 source.n17 a_n1528_n1288# 0.194726f
C124 source.n18 a_n1528_n1288# 0.043768f
C125 source.n19 a_n1528_n1288# 0.108003f
C126 source.n20 a_n1528_n1288# 0.039926f
C127 source.n21 a_n1528_n1288# 0.088341f
C128 source.t9 a_n1528_n1288# 0.066296f
C129 source.n22 a_n1528_n1288# 0.069139f
C130 source.n23 a_n1528_n1288# 0.022288f
C131 source.n24 a_n1528_n1288# 0.014699f
C132 source.n25 a_n1528_n1288# 0.194726f
C133 source.n26 a_n1528_n1288# 0.043768f
C134 source.n27 a_n1528_n1288# 0.108003f
C135 source.t2 a_n1528_n1288# 0.043233f
C136 source.t5 a_n1528_n1288# 0.043233f
C137 source.n28 a_n1528_n1288# 0.231124f
C138 source.n29 a_n1528_n1288# 0.300814f
C139 source.t23 a_n1528_n1288# 0.043233f
C140 source.t4 a_n1528_n1288# 0.043233f
C141 source.n30 a_n1528_n1288# 0.231124f
C142 source.n31 a_n1528_n1288# 0.300814f
C143 source.n32 a_n1528_n1288# 0.039926f
C144 source.n33 a_n1528_n1288# 0.088341f
C145 source.t3 a_n1528_n1288# 0.066296f
C146 source.n34 a_n1528_n1288# 0.069139f
C147 source.n35 a_n1528_n1288# 0.022288f
C148 source.n36 a_n1528_n1288# 0.014699f
C149 source.n37 a_n1528_n1288# 0.194726f
C150 source.n38 a_n1528_n1288# 0.043768f
C151 source.n39 a_n1528_n1288# 0.660444f
C152 source.n40 a_n1528_n1288# 0.039926f
C153 source.n41 a_n1528_n1288# 0.088341f
C154 source.t12 a_n1528_n1288# 0.066296f
C155 source.n42 a_n1528_n1288# 0.069139f
C156 source.n43 a_n1528_n1288# 0.022288f
C157 source.n44 a_n1528_n1288# 0.014699f
C158 source.n45 a_n1528_n1288# 0.194726f
C159 source.n46 a_n1528_n1288# 0.043768f
C160 source.n47 a_n1528_n1288# 0.660445f
C161 source.t21 a_n1528_n1288# 0.043233f
C162 source.t14 a_n1528_n1288# 0.043233f
C163 source.n48 a_n1528_n1288# 0.231122f
C164 source.n49 a_n1528_n1288# 0.300816f
C165 source.t11 a_n1528_n1288# 0.043233f
C166 source.t20 a_n1528_n1288# 0.043233f
C167 source.n50 a_n1528_n1288# 0.231122f
C168 source.n51 a_n1528_n1288# 0.300816f
C169 source.n52 a_n1528_n1288# 0.039926f
C170 source.n53 a_n1528_n1288# 0.088341f
C171 source.t16 a_n1528_n1288# 0.066296f
C172 source.n54 a_n1528_n1288# 0.069139f
C173 source.n55 a_n1528_n1288# 0.022288f
C174 source.n56 a_n1528_n1288# 0.014699f
C175 source.n57 a_n1528_n1288# 0.194726f
C176 source.n58 a_n1528_n1288# 0.043768f
C177 source.n59 a_n1528_n1288# 0.108003f
C178 source.n60 a_n1528_n1288# 0.039926f
C179 source.n61 a_n1528_n1288# 0.088341f
C180 source.t1 a_n1528_n1288# 0.066296f
C181 source.n62 a_n1528_n1288# 0.069139f
C182 source.n63 a_n1528_n1288# 0.022288f
C183 source.n64 a_n1528_n1288# 0.014699f
C184 source.n65 a_n1528_n1288# 0.194726f
C185 source.n66 a_n1528_n1288# 0.043768f
C186 source.n67 a_n1528_n1288# 0.108003f
C187 source.t8 a_n1528_n1288# 0.043233f
C188 source.t7 a_n1528_n1288# 0.043233f
C189 source.n68 a_n1528_n1288# 0.231122f
C190 source.n69 a_n1528_n1288# 0.300816f
C191 source.t6 a_n1528_n1288# 0.043233f
C192 source.t0 a_n1528_n1288# 0.043233f
C193 source.n70 a_n1528_n1288# 0.231122f
C194 source.n71 a_n1528_n1288# 0.300816f
C195 source.n72 a_n1528_n1288# 0.039926f
C196 source.n73 a_n1528_n1288# 0.088341f
C197 source.t22 a_n1528_n1288# 0.066296f
C198 source.n74 a_n1528_n1288# 0.069139f
C199 source.n75 a_n1528_n1288# 0.022288f
C200 source.n76 a_n1528_n1288# 0.014699f
C201 source.n77 a_n1528_n1288# 0.194726f
C202 source.n78 a_n1528_n1288# 0.043768f
C203 source.n79 a_n1528_n1288# 0.25938f
C204 source.n80 a_n1528_n1288# 0.674707f
C205 plus.n0 a_n1528_n1288# 0.032219f
C206 plus.t6 a_n1528_n1288# 0.047403f
C207 plus.t0 a_n1528_n1288# 0.047403f
C208 plus.n1 a_n1528_n1288# 0.011483f
C209 plus.t5 a_n1528_n1288# 0.050243f
C210 plus.n2 a_n1528_n1288# 0.043247f
C211 plus.t1 a_n1528_n1288# 0.047403f
C212 plus.n3 a_n1528_n1288# 0.034762f
C213 plus.t7 a_n1528_n1288# 0.047403f
C214 plus.n4 a_n1528_n1288# 0.034762f
C215 plus.n5 a_n1528_n1288# 0.012277f
C216 plus.n6 a_n1528_n1288# 0.067376f
C217 plus.n7 a_n1528_n1288# 0.032219f
C218 plus.n8 a_n1528_n1288# 0.032219f
C219 plus.n9 a_n1528_n1288# 0.011483f
C220 plus.n10 a_n1528_n1288# 0.034762f
C221 plus.n11 a_n1528_n1288# 0.012277f
C222 plus.n12 a_n1528_n1288# 0.034762f
C223 plus.t11 a_n1528_n1288# 0.050243f
C224 plus.n13 a_n1528_n1288# 0.043206f
C225 plus.n14 a_n1528_n1288# 0.225204f
C226 plus.n15 a_n1528_n1288# 0.032219f
C227 plus.t3 a_n1528_n1288# 0.050243f
C228 plus.t9 a_n1528_n1288# 0.047403f
C229 plus.t4 a_n1528_n1288# 0.047403f
C230 plus.n16 a_n1528_n1288# 0.011483f
C231 plus.t10 a_n1528_n1288# 0.050243f
C232 plus.n17 a_n1528_n1288# 0.043247f
C233 plus.t2 a_n1528_n1288# 0.047403f
C234 plus.n18 a_n1528_n1288# 0.034762f
C235 plus.t8 a_n1528_n1288# 0.047403f
C236 plus.n19 a_n1528_n1288# 0.034762f
C237 plus.n20 a_n1528_n1288# 0.012277f
C238 plus.n21 a_n1528_n1288# 0.067376f
C239 plus.n22 a_n1528_n1288# 0.032219f
C240 plus.n23 a_n1528_n1288# 0.032219f
C241 plus.n24 a_n1528_n1288# 0.011483f
C242 plus.n25 a_n1528_n1288# 0.034762f
C243 plus.n26 a_n1528_n1288# 0.012277f
C244 plus.n27 a_n1528_n1288# 0.034762f
C245 plus.n28 a_n1528_n1288# 0.043206f
C246 plus.n29 a_n1528_n1288# 0.677165f
.ends

