* NGSPICE file created from diffpair67.ext - technology: sky130A

.subckt diffpair67 minus drain_right drain_left source plus
X0 source.t30 plus.t0 drain_left.t7 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X1 source.t29 plus.t1 drain_left.t10 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X2 source.t9 minus.t0 drain_right.t15 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X3 source.t28 plus.t2 drain_left.t13 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X4 drain_left.t3 plus.t3 source.t27 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X5 source.t26 plus.t4 drain_left.t1 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X6 source.t25 plus.t5 drain_left.t12 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X7 drain_right.t14 minus.t1 source.t6 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X8 a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X9 source.t8 minus.t2 drain_right.t13 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X10 source.t24 plus.t6 drain_left.t4 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X11 drain_right.t12 minus.t3 source.t7 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X12 drain_right.t11 minus.t4 source.t14 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X13 drain_right.t10 minus.t5 source.t5 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X14 source.t4 minus.t6 drain_right.t9 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X15 drain_left.t11 plus.t7 source.t23 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X16 source.t3 minus.t7 drain_right.t8 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X17 source.t22 plus.t8 drain_left.t9 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X18 drain_right.t7 minus.t8 source.t13 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X19 drain_left.t6 plus.t9 source.t21 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X20 drain_left.t14 plus.t10 source.t20 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X21 drain_left.t5 plus.t11 source.t19 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X22 drain_right.t6 minus.t9 source.t11 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X23 drain_left.t15 plus.t12 source.t18 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X24 a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X25 source.t10 minus.t10 drain_right.t5 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X26 drain_right.t4 minus.t11 source.t12 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X27 drain_left.t0 plus.t13 source.t17 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X28 source.t2 minus.t12 drain_right.t3 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X29 a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X30 a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X31 source.t1 minus.t13 drain_right.t2 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X32 source.t0 minus.t14 drain_right.t1 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X33 drain_right.t0 minus.t15 source.t31 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X34 source.t16 plus.t14 drain_left.t8 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X35 drain_left.t2 plus.t15 source.t15 a_n2570_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n9 plus.n8 161.3
R1 plus.n10 plus.n5 161.3
R2 plus.n12 plus.n11 161.3
R3 plus.n13 plus.n4 161.3
R4 plus.n15 plus.n14 161.3
R5 plus.n16 plus.n3 161.3
R6 plus.n18 plus.n17 161.3
R7 plus.n19 plus.n2 161.3
R8 plus.n21 plus.n20 161.3
R9 plus.n22 plus.n1 161.3
R10 plus.n23 plus.n0 161.3
R11 plus.n25 plus.n24 161.3
R12 plus.n35 plus.n34 161.3
R13 plus.n36 plus.n31 161.3
R14 plus.n38 plus.n37 161.3
R15 plus.n39 plus.n30 161.3
R16 plus.n41 plus.n40 161.3
R17 plus.n42 plus.n29 161.3
R18 plus.n44 plus.n43 161.3
R19 plus.n45 plus.n28 161.3
R20 plus.n47 plus.n46 161.3
R21 plus.n48 plus.n27 161.3
R22 plus.n49 plus.n26 161.3
R23 plus.n51 plus.n50 161.3
R24 plus.n7 plus.t5 114.922
R25 plus.n33 plus.t9 114.922
R26 plus.n24 plus.t7 90.5476
R27 plus.n22 plus.t0 90.5476
R28 plus.n2 plus.t11 90.5476
R29 plus.n16 plus.t4 90.5476
R30 plus.n4 plus.t10 90.5476
R31 plus.n10 plus.t1 90.5476
R32 plus.n6 plus.t12 90.5476
R33 plus.n50 plus.t6 90.5476
R34 plus.n48 plus.t3 90.5476
R35 plus.n28 plus.t2 90.5476
R36 plus.n42 plus.t15 90.5476
R37 plus.n30 plus.t14 90.5476
R38 plus.n36 plus.t13 90.5476
R39 plus.n32 plus.t8 90.5476
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus.n22 plus.n21 32.8641
R45 plus.n9 plus.n6 32.8641
R46 plus.n48 plus.n47 32.8641
R47 plus.n35 plus.n32 32.8641
R48 plus plus.n51 28.7263
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus.n23 plus.n22 10.955
R68 plus.n49 plus.n48 10.955
R69 plus plus.n25 8.13308
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 drain_left.n9 drain_left.n7 241.02
R93 drain_left.n5 drain_left.n3 241.019
R94 drain_left.n2 drain_left.n0 241.019
R95 drain_left.n13 drain_left.n12 240.132
R96 drain_left.n11 drain_left.n10 240.132
R97 drain_left.n9 drain_left.n8 240.132
R98 drain_left.n5 drain_left.n4 240.131
R99 drain_left.n2 drain_left.n1 240.131
R100 drain_left drain_left.n6 24.8053
R101 drain_left.n3 drain_left.t9 19.8005
R102 drain_left.n3 drain_left.t6 19.8005
R103 drain_left.n4 drain_left.t8 19.8005
R104 drain_left.n4 drain_left.t0 19.8005
R105 drain_left.n1 drain_left.t13 19.8005
R106 drain_left.n1 drain_left.t2 19.8005
R107 drain_left.n0 drain_left.t4 19.8005
R108 drain_left.n0 drain_left.t3 19.8005
R109 drain_left.n12 drain_left.t7 19.8005
R110 drain_left.n12 drain_left.t11 19.8005
R111 drain_left.n10 drain_left.t1 19.8005
R112 drain_left.n10 drain_left.t5 19.8005
R113 drain_left.n8 drain_left.t10 19.8005
R114 drain_left.n8 drain_left.t14 19.8005
R115 drain_left.n7 drain_left.t12 19.8005
R116 drain_left.n7 drain_left.t15 19.8005
R117 drain_left drain_left.n13 6.54115
R118 drain_left.n11 drain_left.n9 0.888431
R119 drain_left.n13 drain_left.n11 0.888431
R120 drain_left.n6 drain_left.n5 0.389119
R121 drain_left.n6 drain_left.n2 0.389119
R122 source.n0 source.t23 243.255
R123 source.n7 source.t25 243.255
R124 source.n8 source.t11 243.255
R125 source.n15 source.t2 243.255
R126 source.n31 source.t31 243.254
R127 source.n24 source.t8 243.254
R128 source.n23 source.t21 243.254
R129 source.n16 source.t24 243.254
R130 source.n2 source.n1 223.454
R131 source.n4 source.n3 223.454
R132 source.n6 source.n5 223.454
R133 source.n10 source.n9 223.454
R134 source.n12 source.n11 223.454
R135 source.n14 source.n13 223.454
R136 source.n30 source.n29 223.453
R137 source.n28 source.n27 223.453
R138 source.n26 source.n25 223.453
R139 source.n22 source.n21 223.453
R140 source.n20 source.n19 223.453
R141 source.n18 source.n17 223.453
R142 source.n29 source.t12 19.8005
R143 source.n29 source.t10 19.8005
R144 source.n27 source.t5 19.8005
R145 source.n27 source.t3 19.8005
R146 source.n25 source.t6 19.8005
R147 source.n25 source.t4 19.8005
R148 source.n21 source.t17 19.8005
R149 source.n21 source.t22 19.8005
R150 source.n19 source.t15 19.8005
R151 source.n19 source.t16 19.8005
R152 source.n17 source.t27 19.8005
R153 source.n17 source.t28 19.8005
R154 source.n1 source.t19 19.8005
R155 source.n1 source.t30 19.8005
R156 source.n3 source.t20 19.8005
R157 source.n3 source.t26 19.8005
R158 source.n5 source.t18 19.8005
R159 source.n5 source.t29 19.8005
R160 source.n9 source.t13 19.8005
R161 source.n9 source.t9 19.8005
R162 source.n11 source.t14 19.8005
R163 source.n11 source.t1 19.8005
R164 source.n13 source.t7 19.8005
R165 source.n13 source.t0 19.8005
R166 source.n16 source.n15 13.8423
R167 source.n32 source.n0 8.13543
R168 source.n32 source.n31 5.7074
R169 source.n15 source.n14 0.888431
R170 source.n14 source.n12 0.888431
R171 source.n12 source.n10 0.888431
R172 source.n10 source.n8 0.888431
R173 source.n7 source.n6 0.888431
R174 source.n6 source.n4 0.888431
R175 source.n4 source.n2 0.888431
R176 source.n2 source.n0 0.888431
R177 source.n18 source.n16 0.888431
R178 source.n20 source.n18 0.888431
R179 source.n22 source.n20 0.888431
R180 source.n23 source.n22 0.888431
R181 source.n26 source.n24 0.888431
R182 source.n28 source.n26 0.888431
R183 source.n30 source.n28 0.888431
R184 source.n31 source.n30 0.888431
R185 source.n8 source.n7 0.470328
R186 source.n24 source.n23 0.470328
R187 source source.n32 0.188
R188 minus.n25 minus.n24 161.3
R189 minus.n23 minus.n0 161.3
R190 minus.n22 minus.n21 161.3
R191 minus.n20 minus.n1 161.3
R192 minus.n19 minus.n18 161.3
R193 minus.n17 minus.n2 161.3
R194 minus.n16 minus.n15 161.3
R195 minus.n14 minus.n3 161.3
R196 minus.n13 minus.n12 161.3
R197 minus.n11 minus.n4 161.3
R198 minus.n10 minus.n9 161.3
R199 minus.n8 minus.n5 161.3
R200 minus.n51 minus.n50 161.3
R201 minus.n49 minus.n26 161.3
R202 minus.n48 minus.n47 161.3
R203 minus.n46 minus.n27 161.3
R204 minus.n45 minus.n44 161.3
R205 minus.n43 minus.n28 161.3
R206 minus.n42 minus.n41 161.3
R207 minus.n40 minus.n29 161.3
R208 minus.n39 minus.n38 161.3
R209 minus.n37 minus.n30 161.3
R210 minus.n36 minus.n35 161.3
R211 minus.n34 minus.n31 161.3
R212 minus.n7 minus.t9 114.922
R213 minus.n33 minus.t2 114.922
R214 minus.n6 minus.t0 90.5476
R215 minus.n10 minus.t8 90.5476
R216 minus.n12 minus.t13 90.5476
R217 minus.n16 minus.t4 90.5476
R218 minus.n18 minus.t14 90.5476
R219 minus.n22 minus.t3 90.5476
R220 minus.n24 minus.t12 90.5476
R221 minus.n32 minus.t1 90.5476
R222 minus.n36 minus.t6 90.5476
R223 minus.n38 minus.t5 90.5476
R224 minus.n42 minus.t7 90.5476
R225 minus.n44 minus.t11 90.5476
R226 minus.n48 minus.t10 90.5476
R227 minus.n50 minus.t15 90.5476
R228 minus.n8 minus.n7 44.9377
R229 minus.n34 minus.n33 44.9377
R230 minus.n24 minus.n23 37.246
R231 minus.n50 minus.n49 37.246
R232 minus.n6 minus.n5 32.8641
R233 minus.n22 minus.n1 32.8641
R234 minus.n32 minus.n31 32.8641
R235 minus.n48 minus.n27 32.8641
R236 minus.n52 minus.n25 30.6785
R237 minus.n11 minus.n10 28.4823
R238 minus.n18 minus.n17 28.4823
R239 minus.n37 minus.n36 28.4823
R240 minus.n44 minus.n43 28.4823
R241 minus.n16 minus.n3 24.1005
R242 minus.n12 minus.n3 24.1005
R243 minus.n38 minus.n29 24.1005
R244 minus.n42 minus.n29 24.1005
R245 minus.n12 minus.n11 19.7187
R246 minus.n17 minus.n16 19.7187
R247 minus.n38 minus.n37 19.7187
R248 minus.n43 minus.n42 19.7187
R249 minus.n7 minus.n6 17.0522
R250 minus.n33 minus.n32 17.0522
R251 minus.n10 minus.n5 15.3369
R252 minus.n18 minus.n1 15.3369
R253 minus.n36 minus.n31 15.3369
R254 minus.n44 minus.n27 15.3369
R255 minus.n23 minus.n22 10.955
R256 minus.n49 minus.n48 10.955
R257 minus.n52 minus.n51 6.6558
R258 minus.n25 minus.n0 0.189894
R259 minus.n21 minus.n0 0.189894
R260 minus.n21 minus.n20 0.189894
R261 minus.n20 minus.n19 0.189894
R262 minus.n19 minus.n2 0.189894
R263 minus.n15 minus.n2 0.189894
R264 minus.n15 minus.n14 0.189894
R265 minus.n14 minus.n13 0.189894
R266 minus.n13 minus.n4 0.189894
R267 minus.n9 minus.n4 0.189894
R268 minus.n9 minus.n8 0.189894
R269 minus.n35 minus.n34 0.189894
R270 minus.n35 minus.n30 0.189894
R271 minus.n39 minus.n30 0.189894
R272 minus.n40 minus.n39 0.189894
R273 minus.n41 minus.n40 0.189894
R274 minus.n41 minus.n28 0.189894
R275 minus.n45 minus.n28 0.189894
R276 minus.n46 minus.n45 0.189894
R277 minus.n47 minus.n46 0.189894
R278 minus.n47 minus.n26 0.189894
R279 minus.n51 minus.n26 0.189894
R280 minus minus.n52 0.188
R281 drain_right.n9 drain_right.n7 241.02
R282 drain_right.n5 drain_right.n3 241.019
R283 drain_right.n2 drain_right.n0 241.019
R284 drain_right.n9 drain_right.n8 240.132
R285 drain_right.n11 drain_right.n10 240.132
R286 drain_right.n13 drain_right.n12 240.132
R287 drain_right.n5 drain_right.n4 240.131
R288 drain_right.n2 drain_right.n1 240.131
R289 drain_right drain_right.n6 24.2521
R290 drain_right.n3 drain_right.t5 19.8005
R291 drain_right.n3 drain_right.t0 19.8005
R292 drain_right.n4 drain_right.t8 19.8005
R293 drain_right.n4 drain_right.t4 19.8005
R294 drain_right.n1 drain_right.t9 19.8005
R295 drain_right.n1 drain_right.t10 19.8005
R296 drain_right.n0 drain_right.t13 19.8005
R297 drain_right.n0 drain_right.t14 19.8005
R298 drain_right.n7 drain_right.t15 19.8005
R299 drain_right.n7 drain_right.t6 19.8005
R300 drain_right.n8 drain_right.t2 19.8005
R301 drain_right.n8 drain_right.t7 19.8005
R302 drain_right.n10 drain_right.t1 19.8005
R303 drain_right.n10 drain_right.t11 19.8005
R304 drain_right.n12 drain_right.t3 19.8005
R305 drain_right.n12 drain_right.t12 19.8005
R306 drain_right drain_right.n13 6.54115
R307 drain_right.n13 drain_right.n11 0.888431
R308 drain_right.n11 drain_right.n9 0.888431
R309 drain_right.n6 drain_right.n5 0.389119
R310 drain_right.n6 drain_right.n2 0.389119
C0 minus source 2.08087f
C1 plus drain_left 1.65558f
C2 plus drain_right 0.419367f
C3 source drain_left 4.82159f
C4 source drain_right 4.82382f
C5 minus drain_left 0.179948f
C6 minus drain_right 1.40112f
C7 drain_left drain_right 1.34357f
C8 source plus 2.09474f
C9 minus plus 4.32273f
C10 drain_right a_n2570_n1088# 4.25102f
C11 drain_left a_n2570_n1088# 4.57292f
C12 source a_n2570_n1088# 2.750302f
C13 minus a_n2570_n1088# 9.330372f
C14 plus a_n2570_n1088# 10.314101f
C15 drain_right.t13 a_n2570_n1088# 0.016051f
C16 drain_right.t14 a_n2570_n1088# 0.016051f
C17 drain_right.n0 a_n2570_n1088# 0.063351f
C18 drain_right.t9 a_n2570_n1088# 0.016051f
C19 drain_right.t10 a_n2570_n1088# 0.016051f
C20 drain_right.n1 a_n2570_n1088# 0.06237f
C21 drain_right.n2 a_n2570_n1088# 0.492277f
C22 drain_right.t5 a_n2570_n1088# 0.016051f
C23 drain_right.t0 a_n2570_n1088# 0.016051f
C24 drain_right.n3 a_n2570_n1088# 0.063351f
C25 drain_right.t8 a_n2570_n1088# 0.016051f
C26 drain_right.t4 a_n2570_n1088# 0.016051f
C27 drain_right.n4 a_n2570_n1088# 0.06237f
C28 drain_right.n5 a_n2570_n1088# 0.492277f
C29 drain_right.n6 a_n2570_n1088# 0.670068f
C30 drain_right.t15 a_n2570_n1088# 0.016051f
C31 drain_right.t6 a_n2570_n1088# 0.016051f
C32 drain_right.n7 a_n2570_n1088# 0.063351f
C33 drain_right.t2 a_n2570_n1088# 0.016051f
C34 drain_right.t7 a_n2570_n1088# 0.016051f
C35 drain_right.n8 a_n2570_n1088# 0.06237f
C36 drain_right.n9 a_n2570_n1088# 0.523745f
C37 drain_right.t1 a_n2570_n1088# 0.016051f
C38 drain_right.t11 a_n2570_n1088# 0.016051f
C39 drain_right.n10 a_n2570_n1088# 0.06237f
C40 drain_right.n11 a_n2570_n1088# 0.258273f
C41 drain_right.t3 a_n2570_n1088# 0.016051f
C42 drain_right.t12 a_n2570_n1088# 0.016051f
C43 drain_right.n12 a_n2570_n1088# 0.06237f
C44 drain_right.n13 a_n2570_n1088# 0.437933f
C45 minus.n0 a_n2570_n1088# 0.036504f
C46 minus.n1 a_n2570_n1088# 0.008283f
C47 minus.t3 a_n2570_n1088# 0.086648f
C48 minus.n2 a_n2570_n1088# 0.036504f
C49 minus.n3 a_n2570_n1088# 0.008283f
C50 minus.t4 a_n2570_n1088# 0.086648f
C51 minus.n4 a_n2570_n1088# 0.036504f
C52 minus.n5 a_n2570_n1088# 0.008283f
C53 minus.t8 a_n2570_n1088# 0.086648f
C54 minus.t9 a_n2570_n1088# 0.104949f
C55 minus.t0 a_n2570_n1088# 0.086648f
C56 minus.n6 a_n2570_n1088# 0.091141f
C57 minus.n7 a_n2570_n1088# 0.070878f
C58 minus.n8 a_n2570_n1088# 0.154474f
C59 minus.n9 a_n2570_n1088# 0.036504f
C60 minus.n10 a_n2570_n1088# 0.086141f
C61 minus.n11 a_n2570_n1088# 0.008283f
C62 minus.t13 a_n2570_n1088# 0.086648f
C63 minus.n12 a_n2570_n1088# 0.086141f
C64 minus.n13 a_n2570_n1088# 0.036504f
C65 minus.n14 a_n2570_n1088# 0.036504f
C66 minus.n15 a_n2570_n1088# 0.036504f
C67 minus.n16 a_n2570_n1088# 0.086141f
C68 minus.n17 a_n2570_n1088# 0.008283f
C69 minus.t14 a_n2570_n1088# 0.086648f
C70 minus.n18 a_n2570_n1088# 0.086141f
C71 minus.n19 a_n2570_n1088# 0.036504f
C72 minus.n20 a_n2570_n1088# 0.036504f
C73 minus.n21 a_n2570_n1088# 0.036504f
C74 minus.n22 a_n2570_n1088# 0.086141f
C75 minus.n23 a_n2570_n1088# 0.008283f
C76 minus.t12 a_n2570_n1088# 0.086648f
C77 minus.n24 a_n2570_n1088# 0.085128f
C78 minus.n25 a_n2570_n1088# 0.991544f
C79 minus.n26 a_n2570_n1088# 0.036504f
C80 minus.n27 a_n2570_n1088# 0.008283f
C81 minus.n28 a_n2570_n1088# 0.036504f
C82 minus.n29 a_n2570_n1088# 0.008283f
C83 minus.n30 a_n2570_n1088# 0.036504f
C84 minus.n31 a_n2570_n1088# 0.008283f
C85 minus.t2 a_n2570_n1088# 0.104949f
C86 minus.t1 a_n2570_n1088# 0.086648f
C87 minus.n32 a_n2570_n1088# 0.091141f
C88 minus.n33 a_n2570_n1088# 0.070878f
C89 minus.n34 a_n2570_n1088# 0.154474f
C90 minus.n35 a_n2570_n1088# 0.036504f
C91 minus.t6 a_n2570_n1088# 0.086648f
C92 minus.n36 a_n2570_n1088# 0.086141f
C93 minus.n37 a_n2570_n1088# 0.008283f
C94 minus.t5 a_n2570_n1088# 0.086648f
C95 minus.n38 a_n2570_n1088# 0.086141f
C96 minus.n39 a_n2570_n1088# 0.036504f
C97 minus.n40 a_n2570_n1088# 0.036504f
C98 minus.n41 a_n2570_n1088# 0.036504f
C99 minus.t7 a_n2570_n1088# 0.086648f
C100 minus.n42 a_n2570_n1088# 0.086141f
C101 minus.n43 a_n2570_n1088# 0.008283f
C102 minus.t11 a_n2570_n1088# 0.086648f
C103 minus.n44 a_n2570_n1088# 0.086141f
C104 minus.n45 a_n2570_n1088# 0.036504f
C105 minus.n46 a_n2570_n1088# 0.036504f
C106 minus.n47 a_n2570_n1088# 0.036504f
C107 minus.t10 a_n2570_n1088# 0.086648f
C108 minus.n48 a_n2570_n1088# 0.086141f
C109 minus.n49 a_n2570_n1088# 0.008283f
C110 minus.t15 a_n2570_n1088# 0.086648f
C111 minus.n50 a_n2570_n1088# 0.085128f
C112 minus.n51 a_n2570_n1088# 0.251953f
C113 minus.n52 a_n2570_n1088# 1.21543f
C114 source.t23 a_n2570_n1088# 0.155834f
C115 source.n0 a_n2570_n1088# 0.739427f
C116 source.t19 a_n2570_n1088# 0.027998f
C117 source.t30 a_n2570_n1088# 0.027998f
C118 source.n1 a_n2570_n1088# 0.090802f
C119 source.n2 a_n2570_n1088# 0.420342f
C120 source.t20 a_n2570_n1088# 0.027998f
C121 source.t26 a_n2570_n1088# 0.027998f
C122 source.n3 a_n2570_n1088# 0.090802f
C123 source.n4 a_n2570_n1088# 0.420342f
C124 source.t18 a_n2570_n1088# 0.027998f
C125 source.t29 a_n2570_n1088# 0.027998f
C126 source.n5 a_n2570_n1088# 0.090802f
C127 source.n6 a_n2570_n1088# 0.420342f
C128 source.t25 a_n2570_n1088# 0.155834f
C129 source.n7 a_n2570_n1088# 0.383937f
C130 source.t11 a_n2570_n1088# 0.155834f
C131 source.n8 a_n2570_n1088# 0.383937f
C132 source.t13 a_n2570_n1088# 0.027998f
C133 source.t9 a_n2570_n1088# 0.027998f
C134 source.n9 a_n2570_n1088# 0.090802f
C135 source.n10 a_n2570_n1088# 0.420342f
C136 source.t14 a_n2570_n1088# 0.027998f
C137 source.t1 a_n2570_n1088# 0.027998f
C138 source.n11 a_n2570_n1088# 0.090802f
C139 source.n12 a_n2570_n1088# 0.420342f
C140 source.t7 a_n2570_n1088# 0.027998f
C141 source.t0 a_n2570_n1088# 0.027998f
C142 source.n13 a_n2570_n1088# 0.090802f
C143 source.n14 a_n2570_n1088# 0.420342f
C144 source.t2 a_n2570_n1088# 0.155834f
C145 source.n15 a_n2570_n1088# 1.03176f
C146 source.t24 a_n2570_n1088# 0.155834f
C147 source.n16 a_n2570_n1088# 1.03176f
C148 source.t27 a_n2570_n1088# 0.027998f
C149 source.t28 a_n2570_n1088# 0.027998f
C150 source.n17 a_n2570_n1088# 0.090802f
C151 source.n18 a_n2570_n1088# 0.420342f
C152 source.t15 a_n2570_n1088# 0.027998f
C153 source.t16 a_n2570_n1088# 0.027998f
C154 source.n19 a_n2570_n1088# 0.090802f
C155 source.n20 a_n2570_n1088# 0.420342f
C156 source.t17 a_n2570_n1088# 0.027998f
C157 source.t22 a_n2570_n1088# 0.027998f
C158 source.n21 a_n2570_n1088# 0.090802f
C159 source.n22 a_n2570_n1088# 0.420342f
C160 source.t21 a_n2570_n1088# 0.155834f
C161 source.n23 a_n2570_n1088# 0.383937f
C162 source.t8 a_n2570_n1088# 0.155834f
C163 source.n24 a_n2570_n1088# 0.383937f
C164 source.t6 a_n2570_n1088# 0.027998f
C165 source.t4 a_n2570_n1088# 0.027998f
C166 source.n25 a_n2570_n1088# 0.090802f
C167 source.n26 a_n2570_n1088# 0.420342f
C168 source.t5 a_n2570_n1088# 0.027998f
C169 source.t3 a_n2570_n1088# 0.027998f
C170 source.n27 a_n2570_n1088# 0.090802f
C171 source.n28 a_n2570_n1088# 0.420342f
C172 source.t12 a_n2570_n1088# 0.027998f
C173 source.t10 a_n2570_n1088# 0.027998f
C174 source.n29 a_n2570_n1088# 0.090802f
C175 source.n30 a_n2570_n1088# 0.420342f
C176 source.t31 a_n2570_n1088# 0.155834f
C177 source.n31 a_n2570_n1088# 0.615051f
C178 source.n32 a_n2570_n1088# 0.73425f
C179 drain_left.t4 a_n2570_n1088# 0.01579f
C180 drain_left.t3 a_n2570_n1088# 0.01579f
C181 drain_left.n0 a_n2570_n1088# 0.06232f
C182 drain_left.t13 a_n2570_n1088# 0.01579f
C183 drain_left.t2 a_n2570_n1088# 0.01579f
C184 drain_left.n1 a_n2570_n1088# 0.061354f
C185 drain_left.n2 a_n2570_n1088# 0.484261f
C186 drain_left.t9 a_n2570_n1088# 0.01579f
C187 drain_left.t6 a_n2570_n1088# 0.01579f
C188 drain_left.n3 a_n2570_n1088# 0.06232f
C189 drain_left.t8 a_n2570_n1088# 0.01579f
C190 drain_left.t0 a_n2570_n1088# 0.01579f
C191 drain_left.n4 a_n2570_n1088# 0.061354f
C192 drain_left.n5 a_n2570_n1088# 0.484261f
C193 drain_left.n6 a_n2570_n1088# 0.697586f
C194 drain_left.t12 a_n2570_n1088# 0.01579f
C195 drain_left.t15 a_n2570_n1088# 0.01579f
C196 drain_left.n7 a_n2570_n1088# 0.06232f
C197 drain_left.t10 a_n2570_n1088# 0.01579f
C198 drain_left.t14 a_n2570_n1088# 0.01579f
C199 drain_left.n8 a_n2570_n1088# 0.061354f
C200 drain_left.n9 a_n2570_n1088# 0.515216f
C201 drain_left.t1 a_n2570_n1088# 0.01579f
C202 drain_left.t5 a_n2570_n1088# 0.01579f
C203 drain_left.n10 a_n2570_n1088# 0.061354f
C204 drain_left.n11 a_n2570_n1088# 0.254067f
C205 drain_left.t7 a_n2570_n1088# 0.01579f
C206 drain_left.t11 a_n2570_n1088# 0.01579f
C207 drain_left.n12 a_n2570_n1088# 0.061354f
C208 drain_left.n13 a_n2570_n1088# 0.430802f
C209 plus.n0 a_n2570_n1088# 0.03693f
C210 plus.t7 a_n2570_n1088# 0.087659f
C211 plus.t0 a_n2570_n1088# 0.087659f
C212 plus.n1 a_n2570_n1088# 0.03693f
C213 plus.t11 a_n2570_n1088# 0.087659f
C214 plus.n2 a_n2570_n1088# 0.087146f
C215 plus.n3 a_n2570_n1088# 0.03693f
C216 plus.t4 a_n2570_n1088# 0.087659f
C217 plus.t10 a_n2570_n1088# 0.087659f
C218 plus.n4 a_n2570_n1088# 0.087146f
C219 plus.n5 a_n2570_n1088# 0.03693f
C220 plus.t1 a_n2570_n1088# 0.087659f
C221 plus.t12 a_n2570_n1088# 0.087659f
C222 plus.n6 a_n2570_n1088# 0.092205f
C223 plus.t5 a_n2570_n1088# 0.106174f
C224 plus.n7 a_n2570_n1088# 0.071705f
C225 plus.n8 a_n2570_n1088# 0.156277f
C226 plus.n9 a_n2570_n1088# 0.00838f
C227 plus.n10 a_n2570_n1088# 0.087146f
C228 plus.n11 a_n2570_n1088# 0.00838f
C229 plus.n12 a_n2570_n1088# 0.03693f
C230 plus.n13 a_n2570_n1088# 0.03693f
C231 plus.n14 a_n2570_n1088# 0.03693f
C232 plus.n15 a_n2570_n1088# 0.00838f
C233 plus.n16 a_n2570_n1088# 0.087146f
C234 plus.n17 a_n2570_n1088# 0.00838f
C235 plus.n18 a_n2570_n1088# 0.03693f
C236 plus.n19 a_n2570_n1088# 0.03693f
C237 plus.n20 a_n2570_n1088# 0.03693f
C238 plus.n21 a_n2570_n1088# 0.00838f
C239 plus.n22 a_n2570_n1088# 0.087146f
C240 plus.n23 a_n2570_n1088# 0.00838f
C241 plus.n24 a_n2570_n1088# 0.086121f
C242 plus.n25 a_n2570_n1088# 0.267379f
C243 plus.n26 a_n2570_n1088# 0.03693f
C244 plus.t6 a_n2570_n1088# 0.087659f
C245 plus.n27 a_n2570_n1088# 0.03693f
C246 plus.t3 a_n2570_n1088# 0.087659f
C247 plus.t2 a_n2570_n1088# 0.087659f
C248 plus.n28 a_n2570_n1088# 0.087146f
C249 plus.n29 a_n2570_n1088# 0.03693f
C250 plus.t15 a_n2570_n1088# 0.087659f
C251 plus.t14 a_n2570_n1088# 0.087659f
C252 plus.n30 a_n2570_n1088# 0.087146f
C253 plus.n31 a_n2570_n1088# 0.03693f
C254 plus.t13 a_n2570_n1088# 0.087659f
C255 plus.t8 a_n2570_n1088# 0.087659f
C256 plus.n32 a_n2570_n1088# 0.092205f
C257 plus.t9 a_n2570_n1088# 0.106174f
C258 plus.n33 a_n2570_n1088# 0.071705f
C259 plus.n34 a_n2570_n1088# 0.156277f
C260 plus.n35 a_n2570_n1088# 0.00838f
C261 plus.n36 a_n2570_n1088# 0.087146f
C262 plus.n37 a_n2570_n1088# 0.00838f
C263 plus.n38 a_n2570_n1088# 0.03693f
C264 plus.n39 a_n2570_n1088# 0.03693f
C265 plus.n40 a_n2570_n1088# 0.03693f
C266 plus.n41 a_n2570_n1088# 0.00838f
C267 plus.n42 a_n2570_n1088# 0.087146f
C268 plus.n43 a_n2570_n1088# 0.00838f
C269 plus.n44 a_n2570_n1088# 0.03693f
C270 plus.n45 a_n2570_n1088# 0.03693f
C271 plus.n46 a_n2570_n1088# 0.03693f
C272 plus.n47 a_n2570_n1088# 0.00838f
C273 plus.n48 a_n2570_n1088# 0.087146f
C274 plus.n49 a_n2570_n1088# 0.00838f
C275 plus.n50 a_n2570_n1088# 0.086121f
C276 plus.n51 a_n2570_n1088# 0.967692f
.ends

