* NGSPICE file created from diffpair268.ext - technology: sky130A

.subckt diffpair268 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t21 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_left.t18 plus.t1 source.t24 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t17 plus.t2 source.t29 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 drain_left.t16 plus.t3 source.t30 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X4 source.t10 minus.t0 drain_right.t19 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X5 drain_left.t15 plus.t4 source.t25 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X6 source.t12 minus.t1 drain_right.t18 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X7 a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X8 a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X9 source.t13 minus.t2 drain_right.t17 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 source.t26 plus.t5 drain_left.t14 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X11 source.t35 plus.t6 drain_left.t13 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X12 drain_right.t16 minus.t3 source.t16 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X13 source.t2 minus.t4 drain_right.t15 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X14 drain_right.t14 minus.t5 source.t7 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 drain_left.t12 plus.t7 source.t19 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X16 source.t1 minus.t6 drain_right.t13 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X17 source.t5 minus.t7 drain_right.t12 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X18 source.t20 plus.t8 drain_left.t11 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 drain_left.t10 plus.t9 source.t32 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X20 source.t11 minus.t8 drain_right.t11 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X21 source.t15 minus.t9 drain_right.t10 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X22 source.t27 plus.t10 drain_left.t9 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X23 source.t31 plus.t11 drain_left.t8 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X24 source.t22 plus.t12 drain_left.t7 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X25 source.t37 plus.t13 drain_left.t6 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X26 drain_left.t5 plus.t14 source.t34 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X27 drain_right.t9 minus.t10 source.t9 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X28 drain_right.t8 minus.t11 source.t8 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X29 source.t38 minus.t12 drain_right.t7 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X30 source.t36 plus.t15 drain_left.t4 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X31 drain_right.t6 minus.t13 source.t39 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X32 a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X33 source.t28 plus.t16 drain_left.t3 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X34 a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X35 drain_right.t5 minus.t14 source.t4 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X36 drain_right.t4 minus.t15 source.t0 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X37 drain_left.t2 plus.t17 source.t18 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X38 drain_right.t3 minus.t16 source.t3 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X39 drain_right.t2 minus.t17 source.t17 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X40 drain_right.t1 minus.t18 source.t14 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X41 source.t6 minus.t19 drain_right.t0 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X42 drain_left.t1 plus.t18 source.t23 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X43 source.t33 plus.t19 drain_left.t0 a_n1992_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
R0 plus.n6 plus.t5 756.303
R1 plus.n25 plus.t3 756.303
R2 plus.n33 plus.t14 756.303
R3 plus.n52 plus.t6 756.303
R4 plus.n5 plus.t1 703.721
R5 plus.n9 plus.t13 703.721
R6 plus.n11 plus.t0 703.721
R7 plus.n3 plus.t12 703.721
R8 plus.n17 plus.t18 703.721
R9 plus.n1 plus.t11 703.721
R10 plus.n22 plus.t4 703.721
R11 plus.n24 plus.t15 703.721
R12 plus.n32 plus.t8 703.721
R13 plus.n36 plus.t2 703.721
R14 plus.n38 plus.t16 703.721
R15 plus.n30 plus.t17 703.721
R16 plus.n44 plus.t10 703.721
R17 plus.n28 plus.t7 703.721
R18 plus.n49 plus.t19 703.721
R19 plus.n51 plus.t9 703.721
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus.n10 plus.n9 29.2126
R63 plus.n22 plus.n21 29.2126
R64 plus.n49 plus.n48 29.2126
R65 plus.n37 plus.n36 29.2126
R66 plus plus.n53 28.2717
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 9.86792
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n282 source.n256 289.615
R93 source.n242 source.n216 289.615
R94 source.n210 source.n184 289.615
R95 source.n170 source.n144 289.615
R96 source.n26 source.n0 289.615
R97 source.n66 source.n40 289.615
R98 source.n98 source.n72 289.615
R99 source.n138 source.n112 289.615
R100 source.n267 source.n266 185
R101 source.n264 source.n263 185
R102 source.n273 source.n272 185
R103 source.n275 source.n274 185
R104 source.n260 source.n259 185
R105 source.n281 source.n280 185
R106 source.n283 source.n282 185
R107 source.n227 source.n226 185
R108 source.n224 source.n223 185
R109 source.n233 source.n232 185
R110 source.n235 source.n234 185
R111 source.n220 source.n219 185
R112 source.n241 source.n240 185
R113 source.n243 source.n242 185
R114 source.n195 source.n194 185
R115 source.n192 source.n191 185
R116 source.n201 source.n200 185
R117 source.n203 source.n202 185
R118 source.n188 source.n187 185
R119 source.n209 source.n208 185
R120 source.n211 source.n210 185
R121 source.n155 source.n154 185
R122 source.n152 source.n151 185
R123 source.n161 source.n160 185
R124 source.n163 source.n162 185
R125 source.n148 source.n147 185
R126 source.n169 source.n168 185
R127 source.n171 source.n170 185
R128 source.n27 source.n26 185
R129 source.n25 source.n24 185
R130 source.n4 source.n3 185
R131 source.n19 source.n18 185
R132 source.n17 source.n16 185
R133 source.n8 source.n7 185
R134 source.n11 source.n10 185
R135 source.n67 source.n66 185
R136 source.n65 source.n64 185
R137 source.n44 source.n43 185
R138 source.n59 source.n58 185
R139 source.n57 source.n56 185
R140 source.n48 source.n47 185
R141 source.n51 source.n50 185
R142 source.n99 source.n98 185
R143 source.n97 source.n96 185
R144 source.n76 source.n75 185
R145 source.n91 source.n90 185
R146 source.n89 source.n88 185
R147 source.n80 source.n79 185
R148 source.n83 source.n82 185
R149 source.n139 source.n138 185
R150 source.n137 source.n136 185
R151 source.n116 source.n115 185
R152 source.n131 source.n130 185
R153 source.n129 source.n128 185
R154 source.n120 source.n119 185
R155 source.n123 source.n122 185
R156 source.t0 source.n265 147.661
R157 source.t38 source.n225 147.661
R158 source.t34 source.n193 147.661
R159 source.t35 source.n153 147.661
R160 source.t30 source.n9 147.661
R161 source.t26 source.n49 147.661
R162 source.t39 source.n81 147.661
R163 source.t11 source.n121 147.661
R164 source.n266 source.n263 104.615
R165 source.n273 source.n263 104.615
R166 source.n274 source.n273 104.615
R167 source.n274 source.n259 104.615
R168 source.n281 source.n259 104.615
R169 source.n282 source.n281 104.615
R170 source.n226 source.n223 104.615
R171 source.n233 source.n223 104.615
R172 source.n234 source.n233 104.615
R173 source.n234 source.n219 104.615
R174 source.n241 source.n219 104.615
R175 source.n242 source.n241 104.615
R176 source.n194 source.n191 104.615
R177 source.n201 source.n191 104.615
R178 source.n202 source.n201 104.615
R179 source.n202 source.n187 104.615
R180 source.n209 source.n187 104.615
R181 source.n210 source.n209 104.615
R182 source.n154 source.n151 104.615
R183 source.n161 source.n151 104.615
R184 source.n162 source.n161 104.615
R185 source.n162 source.n147 104.615
R186 source.n169 source.n147 104.615
R187 source.n170 source.n169 104.615
R188 source.n26 source.n25 104.615
R189 source.n25 source.n3 104.615
R190 source.n18 source.n3 104.615
R191 source.n18 source.n17 104.615
R192 source.n17 source.n7 104.615
R193 source.n10 source.n7 104.615
R194 source.n66 source.n65 104.615
R195 source.n65 source.n43 104.615
R196 source.n58 source.n43 104.615
R197 source.n58 source.n57 104.615
R198 source.n57 source.n47 104.615
R199 source.n50 source.n47 104.615
R200 source.n98 source.n97 104.615
R201 source.n97 source.n75 104.615
R202 source.n90 source.n75 104.615
R203 source.n90 source.n89 104.615
R204 source.n89 source.n79 104.615
R205 source.n82 source.n79 104.615
R206 source.n138 source.n137 104.615
R207 source.n137 source.n115 104.615
R208 source.n130 source.n115 104.615
R209 source.n130 source.n129 104.615
R210 source.n129 source.n119 104.615
R211 source.n122 source.n119 104.615
R212 source.n266 source.t0 52.3082
R213 source.n226 source.t38 52.3082
R214 source.n194 source.t34 52.3082
R215 source.n154 source.t35 52.3082
R216 source.n10 source.t30 52.3082
R217 source.n50 source.t26 52.3082
R218 source.n82 source.t39 52.3082
R219 source.n122 source.t11 52.3082
R220 source.n33 source.n32 50.512
R221 source.n35 source.n34 50.512
R222 source.n37 source.n36 50.512
R223 source.n39 source.n38 50.512
R224 source.n105 source.n104 50.512
R225 source.n107 source.n106 50.512
R226 source.n109 source.n108 50.512
R227 source.n111 source.n110 50.512
R228 source.n255 source.n254 50.5119
R229 source.n253 source.n252 50.5119
R230 source.n251 source.n250 50.5119
R231 source.n249 source.n248 50.5119
R232 source.n183 source.n182 50.5119
R233 source.n181 source.n180 50.5119
R234 source.n179 source.n178 50.5119
R235 source.n177 source.n176 50.5119
R236 source.n287 source.n286 32.1853
R237 source.n247 source.n246 32.1853
R238 source.n215 source.n214 32.1853
R239 source.n175 source.n174 32.1853
R240 source.n31 source.n30 32.1853
R241 source.n71 source.n70 32.1853
R242 source.n103 source.n102 32.1853
R243 source.n143 source.n142 32.1853
R244 source.n175 source.n143 17.2423
R245 source.n267 source.n265 15.6674
R246 source.n227 source.n225 15.6674
R247 source.n195 source.n193 15.6674
R248 source.n155 source.n153 15.6674
R249 source.n11 source.n9 15.6674
R250 source.n51 source.n49 15.6674
R251 source.n83 source.n81 15.6674
R252 source.n123 source.n121 15.6674
R253 source.n268 source.n264 12.8005
R254 source.n228 source.n224 12.8005
R255 source.n196 source.n192 12.8005
R256 source.n156 source.n152 12.8005
R257 source.n12 source.n8 12.8005
R258 source.n52 source.n48 12.8005
R259 source.n84 source.n80 12.8005
R260 source.n124 source.n120 12.8005
R261 source.n272 source.n271 12.0247
R262 source.n232 source.n231 12.0247
R263 source.n200 source.n199 12.0247
R264 source.n160 source.n159 12.0247
R265 source.n16 source.n15 12.0247
R266 source.n56 source.n55 12.0247
R267 source.n88 source.n87 12.0247
R268 source.n128 source.n127 12.0247
R269 source.n288 source.n31 11.7293
R270 source.n275 source.n262 11.249
R271 source.n235 source.n222 11.249
R272 source.n203 source.n190 11.249
R273 source.n163 source.n150 11.249
R274 source.n19 source.n6 11.249
R275 source.n59 source.n46 11.249
R276 source.n91 source.n78 11.249
R277 source.n131 source.n118 11.249
R278 source.n276 source.n260 10.4732
R279 source.n236 source.n220 10.4732
R280 source.n204 source.n188 10.4732
R281 source.n164 source.n148 10.4732
R282 source.n20 source.n4 10.4732
R283 source.n60 source.n44 10.4732
R284 source.n92 source.n76 10.4732
R285 source.n132 source.n116 10.4732
R286 source.n280 source.n279 9.69747
R287 source.n240 source.n239 9.69747
R288 source.n208 source.n207 9.69747
R289 source.n168 source.n167 9.69747
R290 source.n24 source.n23 9.69747
R291 source.n64 source.n63 9.69747
R292 source.n96 source.n95 9.69747
R293 source.n136 source.n135 9.69747
R294 source.n286 source.n285 9.45567
R295 source.n246 source.n245 9.45567
R296 source.n214 source.n213 9.45567
R297 source.n174 source.n173 9.45567
R298 source.n30 source.n29 9.45567
R299 source.n70 source.n69 9.45567
R300 source.n102 source.n101 9.45567
R301 source.n142 source.n141 9.45567
R302 source.n285 source.n284 9.3005
R303 source.n258 source.n257 9.3005
R304 source.n279 source.n278 9.3005
R305 source.n277 source.n276 9.3005
R306 source.n262 source.n261 9.3005
R307 source.n271 source.n270 9.3005
R308 source.n269 source.n268 9.3005
R309 source.n245 source.n244 9.3005
R310 source.n218 source.n217 9.3005
R311 source.n239 source.n238 9.3005
R312 source.n237 source.n236 9.3005
R313 source.n222 source.n221 9.3005
R314 source.n231 source.n230 9.3005
R315 source.n229 source.n228 9.3005
R316 source.n213 source.n212 9.3005
R317 source.n186 source.n185 9.3005
R318 source.n207 source.n206 9.3005
R319 source.n205 source.n204 9.3005
R320 source.n190 source.n189 9.3005
R321 source.n199 source.n198 9.3005
R322 source.n197 source.n196 9.3005
R323 source.n173 source.n172 9.3005
R324 source.n146 source.n145 9.3005
R325 source.n167 source.n166 9.3005
R326 source.n165 source.n164 9.3005
R327 source.n150 source.n149 9.3005
R328 source.n159 source.n158 9.3005
R329 source.n157 source.n156 9.3005
R330 source.n29 source.n28 9.3005
R331 source.n2 source.n1 9.3005
R332 source.n23 source.n22 9.3005
R333 source.n21 source.n20 9.3005
R334 source.n6 source.n5 9.3005
R335 source.n15 source.n14 9.3005
R336 source.n13 source.n12 9.3005
R337 source.n69 source.n68 9.3005
R338 source.n42 source.n41 9.3005
R339 source.n63 source.n62 9.3005
R340 source.n61 source.n60 9.3005
R341 source.n46 source.n45 9.3005
R342 source.n55 source.n54 9.3005
R343 source.n53 source.n52 9.3005
R344 source.n101 source.n100 9.3005
R345 source.n74 source.n73 9.3005
R346 source.n95 source.n94 9.3005
R347 source.n93 source.n92 9.3005
R348 source.n78 source.n77 9.3005
R349 source.n87 source.n86 9.3005
R350 source.n85 source.n84 9.3005
R351 source.n141 source.n140 9.3005
R352 source.n114 source.n113 9.3005
R353 source.n135 source.n134 9.3005
R354 source.n133 source.n132 9.3005
R355 source.n118 source.n117 9.3005
R356 source.n127 source.n126 9.3005
R357 source.n125 source.n124 9.3005
R358 source.n283 source.n258 8.92171
R359 source.n243 source.n218 8.92171
R360 source.n211 source.n186 8.92171
R361 source.n171 source.n146 8.92171
R362 source.n27 source.n2 8.92171
R363 source.n67 source.n42 8.92171
R364 source.n99 source.n74 8.92171
R365 source.n139 source.n114 8.92171
R366 source.n284 source.n256 8.14595
R367 source.n244 source.n216 8.14595
R368 source.n212 source.n184 8.14595
R369 source.n172 source.n144 8.14595
R370 source.n28 source.n0 8.14595
R371 source.n68 source.n40 8.14595
R372 source.n100 source.n72 8.14595
R373 source.n140 source.n112 8.14595
R374 source.n286 source.n256 5.81868
R375 source.n246 source.n216 5.81868
R376 source.n214 source.n184 5.81868
R377 source.n174 source.n144 5.81868
R378 source.n30 source.n0 5.81868
R379 source.n70 source.n40 5.81868
R380 source.n102 source.n72 5.81868
R381 source.n142 source.n112 5.81868
R382 source.n288 source.n287 5.51343
R383 source.n284 source.n283 5.04292
R384 source.n244 source.n243 5.04292
R385 source.n212 source.n211 5.04292
R386 source.n172 source.n171 5.04292
R387 source.n28 source.n27 5.04292
R388 source.n68 source.n67 5.04292
R389 source.n100 source.n99 5.04292
R390 source.n140 source.n139 5.04292
R391 source.n269 source.n265 4.38594
R392 source.n229 source.n225 4.38594
R393 source.n197 source.n193 4.38594
R394 source.n157 source.n153 4.38594
R395 source.n13 source.n9 4.38594
R396 source.n53 source.n49 4.38594
R397 source.n85 source.n81 4.38594
R398 source.n125 source.n121 4.38594
R399 source.n280 source.n258 4.26717
R400 source.n240 source.n218 4.26717
R401 source.n208 source.n186 4.26717
R402 source.n168 source.n146 4.26717
R403 source.n24 source.n2 4.26717
R404 source.n64 source.n42 4.26717
R405 source.n96 source.n74 4.26717
R406 source.n136 source.n114 4.26717
R407 source.n279 source.n260 3.49141
R408 source.n239 source.n220 3.49141
R409 source.n207 source.n188 3.49141
R410 source.n167 source.n148 3.49141
R411 source.n23 source.n4 3.49141
R412 source.n63 source.n44 3.49141
R413 source.n95 source.n76 3.49141
R414 source.n135 source.n116 3.49141
R415 source.n254 source.t7 3.3005
R416 source.n254 source.t13 3.3005
R417 source.n252 source.t9 3.3005
R418 source.n252 source.t5 3.3005
R419 source.n250 source.t16 3.3005
R420 source.n250 source.t6 3.3005
R421 source.n248 source.t4 3.3005
R422 source.n248 source.t15 3.3005
R423 source.n182 source.t29 3.3005
R424 source.n182 source.t20 3.3005
R425 source.n180 source.t18 3.3005
R426 source.n180 source.t28 3.3005
R427 source.n178 source.t19 3.3005
R428 source.n178 source.t27 3.3005
R429 source.n176 source.t32 3.3005
R430 source.n176 source.t33 3.3005
R431 source.n32 source.t25 3.3005
R432 source.n32 source.t36 3.3005
R433 source.n34 source.t23 3.3005
R434 source.n34 source.t31 3.3005
R435 source.n36 source.t21 3.3005
R436 source.n36 source.t22 3.3005
R437 source.n38 source.t24 3.3005
R438 source.n38 source.t37 3.3005
R439 source.n104 source.t8 3.3005
R440 source.n104 source.t12 3.3005
R441 source.n106 source.t3 3.3005
R442 source.n106 source.t10 3.3005
R443 source.n108 source.t17 3.3005
R444 source.n108 source.t1 3.3005
R445 source.n110 source.t14 3.3005
R446 source.n110 source.t2 3.3005
R447 source.n276 source.n275 2.71565
R448 source.n236 source.n235 2.71565
R449 source.n204 source.n203 2.71565
R450 source.n164 source.n163 2.71565
R451 source.n20 source.n19 2.71565
R452 source.n60 source.n59 2.71565
R453 source.n92 source.n91 2.71565
R454 source.n132 source.n131 2.71565
R455 source.n272 source.n262 1.93989
R456 source.n232 source.n222 1.93989
R457 source.n200 source.n190 1.93989
R458 source.n160 source.n150 1.93989
R459 source.n16 source.n6 1.93989
R460 source.n56 source.n46 1.93989
R461 source.n88 source.n78 1.93989
R462 source.n128 source.n118 1.93989
R463 source.n271 source.n264 1.16414
R464 source.n231 source.n224 1.16414
R465 source.n199 source.n192 1.16414
R466 source.n159 source.n152 1.16414
R467 source.n15 source.n8 1.16414
R468 source.n55 source.n48 1.16414
R469 source.n87 source.n80 1.16414
R470 source.n127 source.n120 1.16414
R471 source.n143 source.n111 0.5005
R472 source.n111 source.n109 0.5005
R473 source.n109 source.n107 0.5005
R474 source.n107 source.n105 0.5005
R475 source.n105 source.n103 0.5005
R476 source.n71 source.n39 0.5005
R477 source.n39 source.n37 0.5005
R478 source.n37 source.n35 0.5005
R479 source.n35 source.n33 0.5005
R480 source.n33 source.n31 0.5005
R481 source.n177 source.n175 0.5005
R482 source.n179 source.n177 0.5005
R483 source.n181 source.n179 0.5005
R484 source.n183 source.n181 0.5005
R485 source.n215 source.n183 0.5005
R486 source.n249 source.n247 0.5005
R487 source.n251 source.n249 0.5005
R488 source.n253 source.n251 0.5005
R489 source.n255 source.n253 0.5005
R490 source.n287 source.n255 0.5005
R491 source.n103 source.n71 0.470328
R492 source.n247 source.n215 0.470328
R493 source.n268 source.n267 0.388379
R494 source.n228 source.n227 0.388379
R495 source.n196 source.n195 0.388379
R496 source.n156 source.n155 0.388379
R497 source.n12 source.n11 0.388379
R498 source.n52 source.n51 0.388379
R499 source.n84 source.n83 0.388379
R500 source.n124 source.n123 0.388379
R501 source source.n288 0.188
R502 source.n270 source.n269 0.155672
R503 source.n270 source.n261 0.155672
R504 source.n277 source.n261 0.155672
R505 source.n278 source.n277 0.155672
R506 source.n278 source.n257 0.155672
R507 source.n285 source.n257 0.155672
R508 source.n230 source.n229 0.155672
R509 source.n230 source.n221 0.155672
R510 source.n237 source.n221 0.155672
R511 source.n238 source.n237 0.155672
R512 source.n238 source.n217 0.155672
R513 source.n245 source.n217 0.155672
R514 source.n198 source.n197 0.155672
R515 source.n198 source.n189 0.155672
R516 source.n205 source.n189 0.155672
R517 source.n206 source.n205 0.155672
R518 source.n206 source.n185 0.155672
R519 source.n213 source.n185 0.155672
R520 source.n158 source.n157 0.155672
R521 source.n158 source.n149 0.155672
R522 source.n165 source.n149 0.155672
R523 source.n166 source.n165 0.155672
R524 source.n166 source.n145 0.155672
R525 source.n173 source.n145 0.155672
R526 source.n29 source.n1 0.155672
R527 source.n22 source.n1 0.155672
R528 source.n22 source.n21 0.155672
R529 source.n21 source.n5 0.155672
R530 source.n14 source.n5 0.155672
R531 source.n14 source.n13 0.155672
R532 source.n69 source.n41 0.155672
R533 source.n62 source.n41 0.155672
R534 source.n62 source.n61 0.155672
R535 source.n61 source.n45 0.155672
R536 source.n54 source.n45 0.155672
R537 source.n54 source.n53 0.155672
R538 source.n101 source.n73 0.155672
R539 source.n94 source.n73 0.155672
R540 source.n94 source.n93 0.155672
R541 source.n93 source.n77 0.155672
R542 source.n86 source.n77 0.155672
R543 source.n86 source.n85 0.155672
R544 source.n141 source.n113 0.155672
R545 source.n134 source.n113 0.155672
R546 source.n134 source.n133 0.155672
R547 source.n133 source.n117 0.155672
R548 source.n126 source.n117 0.155672
R549 source.n126 source.n125 0.155672
R550 drain_left.n10 drain_left.n8 67.6908
R551 drain_left.n6 drain_left.n4 67.6907
R552 drain_left.n2 drain_left.n0 67.6907
R553 drain_left.n14 drain_left.n13 67.1908
R554 drain_left.n12 drain_left.n11 67.1908
R555 drain_left.n10 drain_left.n9 67.1908
R556 drain_left.n16 drain_left.n15 67.1907
R557 drain_left.n7 drain_left.n3 67.1907
R558 drain_left.n6 drain_left.n5 67.1907
R559 drain_left.n2 drain_left.n1 67.1907
R560 drain_left drain_left.n7 26.8216
R561 drain_left drain_left.n16 6.15322
R562 drain_left.n3 drain_left.t9 3.3005
R563 drain_left.n3 drain_left.t2 3.3005
R564 drain_left.n4 drain_left.t11 3.3005
R565 drain_left.n4 drain_left.t5 3.3005
R566 drain_left.n5 drain_left.t3 3.3005
R567 drain_left.n5 drain_left.t17 3.3005
R568 drain_left.n1 drain_left.t0 3.3005
R569 drain_left.n1 drain_left.t12 3.3005
R570 drain_left.n0 drain_left.t13 3.3005
R571 drain_left.n0 drain_left.t10 3.3005
R572 drain_left.n15 drain_left.t4 3.3005
R573 drain_left.n15 drain_left.t16 3.3005
R574 drain_left.n13 drain_left.t8 3.3005
R575 drain_left.n13 drain_left.t15 3.3005
R576 drain_left.n11 drain_left.t7 3.3005
R577 drain_left.n11 drain_left.t1 3.3005
R578 drain_left.n9 drain_left.t6 3.3005
R579 drain_left.n9 drain_left.t19 3.3005
R580 drain_left.n8 drain_left.t14 3.3005
R581 drain_left.n8 drain_left.t18 3.3005
R582 drain_left.n12 drain_left.n10 0.5005
R583 drain_left.n14 drain_left.n12 0.5005
R584 drain_left.n16 drain_left.n14 0.5005
R585 drain_left.n7 drain_left.n6 0.445154
R586 drain_left.n7 drain_left.n2 0.445154
R587 minus.n25 minus.t8 756.303
R588 minus.n6 minus.t13 756.303
R589 minus.n52 minus.t15 756.303
R590 minus.n33 minus.t12 756.303
R591 minus.n24 minus.t18 703.721
R592 minus.n22 minus.t4 703.721
R593 minus.n1 minus.t17 703.721
R594 minus.n17 minus.t6 703.721
R595 minus.n3 minus.t16 703.721
R596 minus.n11 minus.t0 703.721
R597 minus.n9 minus.t11 703.721
R598 minus.n5 minus.t1 703.721
R599 minus.n51 minus.t2 703.721
R600 minus.n49 minus.t5 703.721
R601 minus.n28 minus.t7 703.721
R602 minus.n44 minus.t10 703.721
R603 minus.n30 minus.t19 703.721
R604 minus.n38 minus.t3 703.721
R605 minus.n36 minus.t9 703.721
R606 minus.n32 minus.t14 703.721
R607 minus.n7 minus.n6 161.489
R608 minus.n34 minus.n33 161.489
R609 minus.n26 minus.n25 161.3
R610 minus.n23 minus.n0 161.3
R611 minus.n21 minus.n20 161.3
R612 minus.n19 minus.n18 161.3
R613 minus.n16 minus.n2 161.3
R614 minus.n15 minus.n14 161.3
R615 minus.n13 minus.n12 161.3
R616 minus.n10 minus.n4 161.3
R617 minus.n8 minus.n7 161.3
R618 minus.n53 minus.n52 161.3
R619 minus.n50 minus.n27 161.3
R620 minus.n48 minus.n47 161.3
R621 minus.n46 minus.n45 161.3
R622 minus.n43 minus.n29 161.3
R623 minus.n42 minus.n41 161.3
R624 minus.n40 minus.n39 161.3
R625 minus.n37 minus.n31 161.3
R626 minus.n35 minus.n34 161.3
R627 minus.n16 minus.n15 73.0308
R628 minus.n43 minus.n42 73.0308
R629 minus.n18 minus.n17 67.1884
R630 minus.n12 minus.n3 67.1884
R631 minus.n39 minus.n30 67.1884
R632 minus.n45 minus.n44 67.1884
R633 minus.n21 minus.n1 55.5035
R634 minus.n11 minus.n10 55.5035
R635 minus.n38 minus.n37 55.5035
R636 minus.n48 minus.n28 55.5035
R637 minus.n23 minus.n22 43.8187
R638 minus.n9 minus.n8 43.8187
R639 minus.n36 minus.n35 43.8187
R640 minus.n50 minus.n49 43.8187
R641 minus.n24 minus.n23 40.8975
R642 minus.n8 minus.n5 40.8975
R643 minus.n35 minus.n32 40.8975
R644 minus.n51 minus.n50 40.8975
R645 minus.n25 minus.n24 32.1338
R646 minus.n6 minus.n5 32.1338
R647 minus.n33 minus.n32 32.1338
R648 minus.n52 minus.n51 32.1338
R649 minus.n54 minus.n26 32.1179
R650 minus.n22 minus.n21 29.2126
R651 minus.n10 minus.n9 29.2126
R652 minus.n37 minus.n36 29.2126
R653 minus.n49 minus.n48 29.2126
R654 minus.n18 minus.n1 17.5278
R655 minus.n12 minus.n11 17.5278
R656 minus.n39 minus.n38 17.5278
R657 minus.n45 minus.n28 17.5278
R658 minus.n54 minus.n53 6.49671
R659 minus.n17 minus.n16 5.84292
R660 minus.n15 minus.n3 5.84292
R661 minus.n42 minus.n30 5.84292
R662 minus.n44 minus.n43 5.84292
R663 minus.n26 minus.n0 0.189894
R664 minus.n20 minus.n0 0.189894
R665 minus.n20 minus.n19 0.189894
R666 minus.n19 minus.n2 0.189894
R667 minus.n14 minus.n2 0.189894
R668 minus.n14 minus.n13 0.189894
R669 minus.n13 minus.n4 0.189894
R670 minus.n7 minus.n4 0.189894
R671 minus.n34 minus.n31 0.189894
R672 minus.n40 minus.n31 0.189894
R673 minus.n41 minus.n40 0.189894
R674 minus.n41 minus.n29 0.189894
R675 minus.n46 minus.n29 0.189894
R676 minus.n47 minus.n46 0.189894
R677 minus.n47 minus.n27 0.189894
R678 minus.n53 minus.n27 0.189894
R679 minus minus.n54 0.188
R680 drain_right.n10 drain_right.n8 67.6907
R681 drain_right.n6 drain_right.n4 67.6907
R682 drain_right.n2 drain_right.n0 67.6907
R683 drain_right.n10 drain_right.n9 67.1908
R684 drain_right.n12 drain_right.n11 67.1908
R685 drain_right.n14 drain_right.n13 67.1908
R686 drain_right.n16 drain_right.n15 67.1908
R687 drain_right.n7 drain_right.n3 67.1907
R688 drain_right.n6 drain_right.n5 67.1907
R689 drain_right.n2 drain_right.n1 67.1907
R690 drain_right drain_right.n7 26.2684
R691 drain_right drain_right.n16 6.15322
R692 drain_right.n3 drain_right.t0 3.3005
R693 drain_right.n3 drain_right.t9 3.3005
R694 drain_right.n4 drain_right.t17 3.3005
R695 drain_right.n4 drain_right.t4 3.3005
R696 drain_right.n5 drain_right.t12 3.3005
R697 drain_right.n5 drain_right.t14 3.3005
R698 drain_right.n1 drain_right.t10 3.3005
R699 drain_right.n1 drain_right.t16 3.3005
R700 drain_right.n0 drain_right.t7 3.3005
R701 drain_right.n0 drain_right.t5 3.3005
R702 drain_right.n8 drain_right.t18 3.3005
R703 drain_right.n8 drain_right.t6 3.3005
R704 drain_right.n9 drain_right.t19 3.3005
R705 drain_right.n9 drain_right.t8 3.3005
R706 drain_right.n11 drain_right.t13 3.3005
R707 drain_right.n11 drain_right.t3 3.3005
R708 drain_right.n13 drain_right.t15 3.3005
R709 drain_right.n13 drain_right.t2 3.3005
R710 drain_right.n15 drain_right.t11 3.3005
R711 drain_right.n15 drain_right.t1 3.3005
R712 drain_right.n16 drain_right.n14 0.5005
R713 drain_right.n14 drain_right.n12 0.5005
R714 drain_right.n12 drain_right.n10 0.5005
R715 drain_right.n7 drain_right.n6 0.445154
R716 drain_right.n7 drain_right.n2 0.445154
C0 minus plus 4.52695f
C1 drain_left plus 3.62371f
C2 minus drain_right 3.42921f
C3 drain_left drain_right 1.04652f
C4 source plus 3.45425f
C5 drain_right source 22.0644f
C6 drain_right plus 0.349242f
C7 minus drain_left 0.171712f
C8 minus source 3.44023f
C9 drain_left source 22.0641f
C10 drain_right a_n1992_n2088# 5.59602f
C11 drain_left a_n1992_n2088# 5.90796f
C12 source a_n1992_n2088# 5.378997f
C13 minus a_n1992_n2088# 7.298873f
C14 plus a_n1992_n2088# 8.95028f
C15 drain_right.t7 a_n1992_n2088# 0.167931f
C16 drain_right.t5 a_n1992_n2088# 0.167931f
C17 drain_right.n0 a_n1992_n2088# 1.40362f
C18 drain_right.t10 a_n1992_n2088# 0.167931f
C19 drain_right.t16 a_n1992_n2088# 0.167931f
C20 drain_right.n1 a_n1992_n2088# 1.40054f
C21 drain_right.n2 a_n1992_n2088# 0.809906f
C22 drain_right.t0 a_n1992_n2088# 0.167931f
C23 drain_right.t9 a_n1992_n2088# 0.167931f
C24 drain_right.n3 a_n1992_n2088# 1.40054f
C25 drain_right.t17 a_n1992_n2088# 0.167931f
C26 drain_right.t4 a_n1992_n2088# 0.167931f
C27 drain_right.n4 a_n1992_n2088# 1.40362f
C28 drain_right.t12 a_n1992_n2088# 0.167931f
C29 drain_right.t14 a_n1992_n2088# 0.167931f
C30 drain_right.n5 a_n1992_n2088# 1.40054f
C31 drain_right.n6 a_n1992_n2088# 0.809906f
C32 drain_right.n7 a_n1992_n2088# 1.59856f
C33 drain_right.t18 a_n1992_n2088# 0.167931f
C34 drain_right.t6 a_n1992_n2088# 0.167931f
C35 drain_right.n8 a_n1992_n2088# 1.40362f
C36 drain_right.t19 a_n1992_n2088# 0.167931f
C37 drain_right.t8 a_n1992_n2088# 0.167931f
C38 drain_right.n9 a_n1992_n2088# 1.40055f
C39 drain_right.n10 a_n1992_n2088# 0.814369f
C40 drain_right.t13 a_n1992_n2088# 0.167931f
C41 drain_right.t3 a_n1992_n2088# 0.167931f
C42 drain_right.n11 a_n1992_n2088# 1.40055f
C43 drain_right.n12 a_n1992_n2088# 0.401584f
C44 drain_right.t15 a_n1992_n2088# 0.167931f
C45 drain_right.t2 a_n1992_n2088# 0.167931f
C46 drain_right.n13 a_n1992_n2088# 1.40055f
C47 drain_right.n14 a_n1992_n2088# 0.401584f
C48 drain_right.t11 a_n1992_n2088# 0.167931f
C49 drain_right.t1 a_n1992_n2088# 0.167931f
C50 drain_right.n15 a_n1992_n2088# 1.40055f
C51 drain_right.n16 a_n1992_n2088# 0.693937f
C52 minus.n0 a_n1992_n2088# 0.05038f
C53 minus.t8 a_n1992_n2088# 0.2226f
C54 minus.t18 a_n1992_n2088# 0.215311f
C55 minus.t4 a_n1992_n2088# 0.215311f
C56 minus.t17 a_n1992_n2088# 0.215311f
C57 minus.n1 a_n1992_n2088# 0.10142f
C58 minus.n2 a_n1992_n2088# 0.05038f
C59 minus.t6 a_n1992_n2088# 0.215311f
C60 minus.t16 a_n1992_n2088# 0.215311f
C61 minus.n3 a_n1992_n2088# 0.10142f
C62 minus.n4 a_n1992_n2088# 0.05038f
C63 minus.t0 a_n1992_n2088# 0.215311f
C64 minus.t11 a_n1992_n2088# 0.215311f
C65 minus.t1 a_n1992_n2088# 0.215311f
C66 minus.n5 a_n1992_n2088# 0.10142f
C67 minus.t13 a_n1992_n2088# 0.2226f
C68 minus.n6 a_n1992_n2088# 0.116822f
C69 minus.n7 a_n1992_n2088# 0.115282f
C70 minus.n8 a_n1992_n2088# 0.019198f
C71 minus.n9 a_n1992_n2088# 0.10142f
C72 minus.n10 a_n1992_n2088# 0.019198f
C73 minus.n11 a_n1992_n2088# 0.10142f
C74 minus.n12 a_n1992_n2088# 0.019198f
C75 minus.n13 a_n1992_n2088# 0.05038f
C76 minus.n14 a_n1992_n2088# 0.05038f
C77 minus.n15 a_n1992_n2088# 0.017955f
C78 minus.n16 a_n1992_n2088# 0.017955f
C79 minus.n17 a_n1992_n2088# 0.10142f
C80 minus.n18 a_n1992_n2088# 0.019198f
C81 minus.n19 a_n1992_n2088# 0.05038f
C82 minus.n20 a_n1992_n2088# 0.05038f
C83 minus.n21 a_n1992_n2088# 0.019198f
C84 minus.n22 a_n1992_n2088# 0.10142f
C85 minus.n23 a_n1992_n2088# 0.019198f
C86 minus.n24 a_n1992_n2088# 0.10142f
C87 minus.n25 a_n1992_n2088# 0.116745f
C88 minus.n26 a_n1992_n2088# 1.46947f
C89 minus.n27 a_n1992_n2088# 0.05038f
C90 minus.t2 a_n1992_n2088# 0.215311f
C91 minus.t5 a_n1992_n2088# 0.215311f
C92 minus.t7 a_n1992_n2088# 0.215311f
C93 minus.n28 a_n1992_n2088# 0.10142f
C94 minus.n29 a_n1992_n2088# 0.05038f
C95 minus.t10 a_n1992_n2088# 0.215311f
C96 minus.t19 a_n1992_n2088# 0.215311f
C97 minus.n30 a_n1992_n2088# 0.10142f
C98 minus.n31 a_n1992_n2088# 0.05038f
C99 minus.t3 a_n1992_n2088# 0.215311f
C100 minus.t9 a_n1992_n2088# 0.215311f
C101 minus.t14 a_n1992_n2088# 0.215311f
C102 minus.n32 a_n1992_n2088# 0.10142f
C103 minus.t12 a_n1992_n2088# 0.2226f
C104 minus.n33 a_n1992_n2088# 0.116822f
C105 minus.n34 a_n1992_n2088# 0.115282f
C106 minus.n35 a_n1992_n2088# 0.019198f
C107 minus.n36 a_n1992_n2088# 0.10142f
C108 minus.n37 a_n1992_n2088# 0.019198f
C109 minus.n38 a_n1992_n2088# 0.10142f
C110 minus.n39 a_n1992_n2088# 0.019198f
C111 minus.n40 a_n1992_n2088# 0.05038f
C112 minus.n41 a_n1992_n2088# 0.05038f
C113 minus.n42 a_n1992_n2088# 0.017955f
C114 minus.n43 a_n1992_n2088# 0.017955f
C115 minus.n44 a_n1992_n2088# 0.10142f
C116 minus.n45 a_n1992_n2088# 0.019198f
C117 minus.n46 a_n1992_n2088# 0.05038f
C118 minus.n47 a_n1992_n2088# 0.05038f
C119 minus.n48 a_n1992_n2088# 0.019198f
C120 minus.n49 a_n1992_n2088# 0.10142f
C121 minus.n50 a_n1992_n2088# 0.019198f
C122 minus.n51 a_n1992_n2088# 0.10142f
C123 minus.t15 a_n1992_n2088# 0.2226f
C124 minus.n52 a_n1992_n2088# 0.116745f
C125 minus.n53 a_n1992_n2088# 0.32898f
C126 minus.n54 a_n1992_n2088# 1.80517f
C127 drain_left.t13 a_n1992_n2088# 0.168333f
C128 drain_left.t10 a_n1992_n2088# 0.168333f
C129 drain_left.n0 a_n1992_n2088# 1.40698f
C130 drain_left.t0 a_n1992_n2088# 0.168333f
C131 drain_left.t12 a_n1992_n2088# 0.168333f
C132 drain_left.n1 a_n1992_n2088# 1.4039f
C133 drain_left.n2 a_n1992_n2088# 0.811847f
C134 drain_left.t9 a_n1992_n2088# 0.168333f
C135 drain_left.t2 a_n1992_n2088# 0.168333f
C136 drain_left.n3 a_n1992_n2088# 1.4039f
C137 drain_left.t11 a_n1992_n2088# 0.168333f
C138 drain_left.t5 a_n1992_n2088# 0.168333f
C139 drain_left.n4 a_n1992_n2088# 1.40698f
C140 drain_left.t3 a_n1992_n2088# 0.168333f
C141 drain_left.t17 a_n1992_n2088# 0.168333f
C142 drain_left.n5 a_n1992_n2088# 1.4039f
C143 drain_left.n6 a_n1992_n2088# 0.811847f
C144 drain_left.n7 a_n1992_n2088# 1.67427f
C145 drain_left.t14 a_n1992_n2088# 0.168333f
C146 drain_left.t18 a_n1992_n2088# 0.168333f
C147 drain_left.n8 a_n1992_n2088# 1.40699f
C148 drain_left.t6 a_n1992_n2088# 0.168333f
C149 drain_left.t19 a_n1992_n2088# 0.168333f
C150 drain_left.n9 a_n1992_n2088# 1.40391f
C151 drain_left.n10 a_n1992_n2088# 0.816314f
C152 drain_left.t7 a_n1992_n2088# 0.168333f
C153 drain_left.t1 a_n1992_n2088# 0.168333f
C154 drain_left.n11 a_n1992_n2088# 1.40391f
C155 drain_left.n12 a_n1992_n2088# 0.402547f
C156 drain_left.t8 a_n1992_n2088# 0.168333f
C157 drain_left.t15 a_n1992_n2088# 0.168333f
C158 drain_left.n13 a_n1992_n2088# 1.40391f
C159 drain_left.n14 a_n1992_n2088# 0.402547f
C160 drain_left.t4 a_n1992_n2088# 0.168333f
C161 drain_left.t16 a_n1992_n2088# 0.168333f
C162 drain_left.n15 a_n1992_n2088# 1.4039f
C163 drain_left.n16 a_n1992_n2088# 0.695607f
C164 source.n0 a_n1992_n2088# 0.045555f
C165 source.n1 a_n1992_n2088# 0.03241f
C166 source.n2 a_n1992_n2088# 0.017416f
C167 source.n3 a_n1992_n2088# 0.041164f
C168 source.n4 a_n1992_n2088# 0.01844f
C169 source.n5 a_n1992_n2088# 0.03241f
C170 source.n6 a_n1992_n2088# 0.017416f
C171 source.n7 a_n1992_n2088# 0.041164f
C172 source.n8 a_n1992_n2088# 0.01844f
C173 source.n9 a_n1992_n2088# 0.138691f
C174 source.t30 a_n1992_n2088# 0.067092f
C175 source.n10 a_n1992_n2088# 0.030873f
C176 source.n11 a_n1992_n2088# 0.024315f
C177 source.n12 a_n1992_n2088# 0.017416f
C178 source.n13 a_n1992_n2088# 0.771158f
C179 source.n14 a_n1992_n2088# 0.03241f
C180 source.n15 a_n1992_n2088# 0.017416f
C181 source.n16 a_n1992_n2088# 0.01844f
C182 source.n17 a_n1992_n2088# 0.041164f
C183 source.n18 a_n1992_n2088# 0.041164f
C184 source.n19 a_n1992_n2088# 0.01844f
C185 source.n20 a_n1992_n2088# 0.017416f
C186 source.n21 a_n1992_n2088# 0.03241f
C187 source.n22 a_n1992_n2088# 0.03241f
C188 source.n23 a_n1992_n2088# 0.017416f
C189 source.n24 a_n1992_n2088# 0.01844f
C190 source.n25 a_n1992_n2088# 0.041164f
C191 source.n26 a_n1992_n2088# 0.089113f
C192 source.n27 a_n1992_n2088# 0.01844f
C193 source.n28 a_n1992_n2088# 0.017416f
C194 source.n29 a_n1992_n2088# 0.074914f
C195 source.n30 a_n1992_n2088# 0.049862f
C196 source.n31 a_n1992_n2088# 0.777309f
C197 source.t25 a_n1992_n2088# 0.153667f
C198 source.t36 a_n1992_n2088# 0.153667f
C199 source.n32 a_n1992_n2088# 1.19677f
C200 source.n33 a_n1992_n2088# 0.408242f
C201 source.t23 a_n1992_n2088# 0.153667f
C202 source.t31 a_n1992_n2088# 0.153667f
C203 source.n34 a_n1992_n2088# 1.19677f
C204 source.n35 a_n1992_n2088# 0.408242f
C205 source.t21 a_n1992_n2088# 0.153667f
C206 source.t22 a_n1992_n2088# 0.153667f
C207 source.n36 a_n1992_n2088# 1.19677f
C208 source.n37 a_n1992_n2088# 0.408242f
C209 source.t24 a_n1992_n2088# 0.153667f
C210 source.t37 a_n1992_n2088# 0.153667f
C211 source.n38 a_n1992_n2088# 1.19677f
C212 source.n39 a_n1992_n2088# 0.408242f
C213 source.n40 a_n1992_n2088# 0.045555f
C214 source.n41 a_n1992_n2088# 0.03241f
C215 source.n42 a_n1992_n2088# 0.017416f
C216 source.n43 a_n1992_n2088# 0.041164f
C217 source.n44 a_n1992_n2088# 0.01844f
C218 source.n45 a_n1992_n2088# 0.03241f
C219 source.n46 a_n1992_n2088# 0.017416f
C220 source.n47 a_n1992_n2088# 0.041164f
C221 source.n48 a_n1992_n2088# 0.01844f
C222 source.n49 a_n1992_n2088# 0.138691f
C223 source.t26 a_n1992_n2088# 0.067092f
C224 source.n50 a_n1992_n2088# 0.030873f
C225 source.n51 a_n1992_n2088# 0.024315f
C226 source.n52 a_n1992_n2088# 0.017416f
C227 source.n53 a_n1992_n2088# 0.771158f
C228 source.n54 a_n1992_n2088# 0.03241f
C229 source.n55 a_n1992_n2088# 0.017416f
C230 source.n56 a_n1992_n2088# 0.01844f
C231 source.n57 a_n1992_n2088# 0.041164f
C232 source.n58 a_n1992_n2088# 0.041164f
C233 source.n59 a_n1992_n2088# 0.01844f
C234 source.n60 a_n1992_n2088# 0.017416f
C235 source.n61 a_n1992_n2088# 0.03241f
C236 source.n62 a_n1992_n2088# 0.03241f
C237 source.n63 a_n1992_n2088# 0.017416f
C238 source.n64 a_n1992_n2088# 0.01844f
C239 source.n65 a_n1992_n2088# 0.041164f
C240 source.n66 a_n1992_n2088# 0.089113f
C241 source.n67 a_n1992_n2088# 0.01844f
C242 source.n68 a_n1992_n2088# 0.017416f
C243 source.n69 a_n1992_n2088# 0.074914f
C244 source.n70 a_n1992_n2088# 0.049862f
C245 source.n71 a_n1992_n2088# 0.128961f
C246 source.n72 a_n1992_n2088# 0.045555f
C247 source.n73 a_n1992_n2088# 0.03241f
C248 source.n74 a_n1992_n2088# 0.017416f
C249 source.n75 a_n1992_n2088# 0.041164f
C250 source.n76 a_n1992_n2088# 0.01844f
C251 source.n77 a_n1992_n2088# 0.03241f
C252 source.n78 a_n1992_n2088# 0.017416f
C253 source.n79 a_n1992_n2088# 0.041164f
C254 source.n80 a_n1992_n2088# 0.01844f
C255 source.n81 a_n1992_n2088# 0.138691f
C256 source.t39 a_n1992_n2088# 0.067092f
C257 source.n82 a_n1992_n2088# 0.030873f
C258 source.n83 a_n1992_n2088# 0.024315f
C259 source.n84 a_n1992_n2088# 0.017416f
C260 source.n85 a_n1992_n2088# 0.771158f
C261 source.n86 a_n1992_n2088# 0.03241f
C262 source.n87 a_n1992_n2088# 0.017416f
C263 source.n88 a_n1992_n2088# 0.01844f
C264 source.n89 a_n1992_n2088# 0.041164f
C265 source.n90 a_n1992_n2088# 0.041164f
C266 source.n91 a_n1992_n2088# 0.01844f
C267 source.n92 a_n1992_n2088# 0.017416f
C268 source.n93 a_n1992_n2088# 0.03241f
C269 source.n94 a_n1992_n2088# 0.03241f
C270 source.n95 a_n1992_n2088# 0.017416f
C271 source.n96 a_n1992_n2088# 0.01844f
C272 source.n97 a_n1992_n2088# 0.041164f
C273 source.n98 a_n1992_n2088# 0.089113f
C274 source.n99 a_n1992_n2088# 0.01844f
C275 source.n100 a_n1992_n2088# 0.017416f
C276 source.n101 a_n1992_n2088# 0.074914f
C277 source.n102 a_n1992_n2088# 0.049862f
C278 source.n103 a_n1992_n2088# 0.128961f
C279 source.t8 a_n1992_n2088# 0.153667f
C280 source.t12 a_n1992_n2088# 0.153667f
C281 source.n104 a_n1992_n2088# 1.19677f
C282 source.n105 a_n1992_n2088# 0.408242f
C283 source.t3 a_n1992_n2088# 0.153667f
C284 source.t10 a_n1992_n2088# 0.153667f
C285 source.n106 a_n1992_n2088# 1.19677f
C286 source.n107 a_n1992_n2088# 0.408242f
C287 source.t17 a_n1992_n2088# 0.153667f
C288 source.t1 a_n1992_n2088# 0.153667f
C289 source.n108 a_n1992_n2088# 1.19677f
C290 source.n109 a_n1992_n2088# 0.408242f
C291 source.t14 a_n1992_n2088# 0.153667f
C292 source.t2 a_n1992_n2088# 0.153667f
C293 source.n110 a_n1992_n2088# 1.19677f
C294 source.n111 a_n1992_n2088# 0.408242f
C295 source.n112 a_n1992_n2088# 0.045555f
C296 source.n113 a_n1992_n2088# 0.03241f
C297 source.n114 a_n1992_n2088# 0.017416f
C298 source.n115 a_n1992_n2088# 0.041164f
C299 source.n116 a_n1992_n2088# 0.01844f
C300 source.n117 a_n1992_n2088# 0.03241f
C301 source.n118 a_n1992_n2088# 0.017416f
C302 source.n119 a_n1992_n2088# 0.041164f
C303 source.n120 a_n1992_n2088# 0.01844f
C304 source.n121 a_n1992_n2088# 0.138691f
C305 source.t11 a_n1992_n2088# 0.067092f
C306 source.n122 a_n1992_n2088# 0.030873f
C307 source.n123 a_n1992_n2088# 0.024315f
C308 source.n124 a_n1992_n2088# 0.017416f
C309 source.n125 a_n1992_n2088# 0.771158f
C310 source.n126 a_n1992_n2088# 0.03241f
C311 source.n127 a_n1992_n2088# 0.017416f
C312 source.n128 a_n1992_n2088# 0.01844f
C313 source.n129 a_n1992_n2088# 0.041164f
C314 source.n130 a_n1992_n2088# 0.041164f
C315 source.n131 a_n1992_n2088# 0.01844f
C316 source.n132 a_n1992_n2088# 0.017416f
C317 source.n133 a_n1992_n2088# 0.03241f
C318 source.n134 a_n1992_n2088# 0.03241f
C319 source.n135 a_n1992_n2088# 0.017416f
C320 source.n136 a_n1992_n2088# 0.01844f
C321 source.n137 a_n1992_n2088# 0.041164f
C322 source.n138 a_n1992_n2088# 0.089113f
C323 source.n139 a_n1992_n2088# 0.01844f
C324 source.n140 a_n1992_n2088# 0.017416f
C325 source.n141 a_n1992_n2088# 0.074914f
C326 source.n142 a_n1992_n2088# 0.049862f
C327 source.n143 a_n1992_n2088# 1.19327f
C328 source.n144 a_n1992_n2088# 0.045555f
C329 source.n145 a_n1992_n2088# 0.03241f
C330 source.n146 a_n1992_n2088# 0.017416f
C331 source.n147 a_n1992_n2088# 0.041164f
C332 source.n148 a_n1992_n2088# 0.01844f
C333 source.n149 a_n1992_n2088# 0.03241f
C334 source.n150 a_n1992_n2088# 0.017416f
C335 source.n151 a_n1992_n2088# 0.041164f
C336 source.n152 a_n1992_n2088# 0.01844f
C337 source.n153 a_n1992_n2088# 0.138691f
C338 source.t35 a_n1992_n2088# 0.067092f
C339 source.n154 a_n1992_n2088# 0.030873f
C340 source.n155 a_n1992_n2088# 0.024315f
C341 source.n156 a_n1992_n2088# 0.017416f
C342 source.n157 a_n1992_n2088# 0.771158f
C343 source.n158 a_n1992_n2088# 0.03241f
C344 source.n159 a_n1992_n2088# 0.017416f
C345 source.n160 a_n1992_n2088# 0.01844f
C346 source.n161 a_n1992_n2088# 0.041164f
C347 source.n162 a_n1992_n2088# 0.041164f
C348 source.n163 a_n1992_n2088# 0.01844f
C349 source.n164 a_n1992_n2088# 0.017416f
C350 source.n165 a_n1992_n2088# 0.03241f
C351 source.n166 a_n1992_n2088# 0.03241f
C352 source.n167 a_n1992_n2088# 0.017416f
C353 source.n168 a_n1992_n2088# 0.01844f
C354 source.n169 a_n1992_n2088# 0.041164f
C355 source.n170 a_n1992_n2088# 0.089113f
C356 source.n171 a_n1992_n2088# 0.01844f
C357 source.n172 a_n1992_n2088# 0.017416f
C358 source.n173 a_n1992_n2088# 0.074914f
C359 source.n174 a_n1992_n2088# 0.049862f
C360 source.n175 a_n1992_n2088# 1.19327f
C361 source.t32 a_n1992_n2088# 0.153667f
C362 source.t33 a_n1992_n2088# 0.153667f
C363 source.n176 a_n1992_n2088# 1.19676f
C364 source.n177 a_n1992_n2088# 0.40825f
C365 source.t19 a_n1992_n2088# 0.153667f
C366 source.t27 a_n1992_n2088# 0.153667f
C367 source.n178 a_n1992_n2088# 1.19676f
C368 source.n179 a_n1992_n2088# 0.40825f
C369 source.t18 a_n1992_n2088# 0.153667f
C370 source.t28 a_n1992_n2088# 0.153667f
C371 source.n180 a_n1992_n2088# 1.19676f
C372 source.n181 a_n1992_n2088# 0.40825f
C373 source.t29 a_n1992_n2088# 0.153667f
C374 source.t20 a_n1992_n2088# 0.153667f
C375 source.n182 a_n1992_n2088# 1.19676f
C376 source.n183 a_n1992_n2088# 0.40825f
C377 source.n184 a_n1992_n2088# 0.045555f
C378 source.n185 a_n1992_n2088# 0.03241f
C379 source.n186 a_n1992_n2088# 0.017416f
C380 source.n187 a_n1992_n2088# 0.041164f
C381 source.n188 a_n1992_n2088# 0.01844f
C382 source.n189 a_n1992_n2088# 0.03241f
C383 source.n190 a_n1992_n2088# 0.017416f
C384 source.n191 a_n1992_n2088# 0.041164f
C385 source.n192 a_n1992_n2088# 0.01844f
C386 source.n193 a_n1992_n2088# 0.138691f
C387 source.t34 a_n1992_n2088# 0.067092f
C388 source.n194 a_n1992_n2088# 0.030873f
C389 source.n195 a_n1992_n2088# 0.024315f
C390 source.n196 a_n1992_n2088# 0.017416f
C391 source.n197 a_n1992_n2088# 0.771158f
C392 source.n198 a_n1992_n2088# 0.03241f
C393 source.n199 a_n1992_n2088# 0.017416f
C394 source.n200 a_n1992_n2088# 0.01844f
C395 source.n201 a_n1992_n2088# 0.041164f
C396 source.n202 a_n1992_n2088# 0.041164f
C397 source.n203 a_n1992_n2088# 0.01844f
C398 source.n204 a_n1992_n2088# 0.017416f
C399 source.n205 a_n1992_n2088# 0.03241f
C400 source.n206 a_n1992_n2088# 0.03241f
C401 source.n207 a_n1992_n2088# 0.017416f
C402 source.n208 a_n1992_n2088# 0.01844f
C403 source.n209 a_n1992_n2088# 0.041164f
C404 source.n210 a_n1992_n2088# 0.089113f
C405 source.n211 a_n1992_n2088# 0.01844f
C406 source.n212 a_n1992_n2088# 0.017416f
C407 source.n213 a_n1992_n2088# 0.074914f
C408 source.n214 a_n1992_n2088# 0.049862f
C409 source.n215 a_n1992_n2088# 0.128961f
C410 source.n216 a_n1992_n2088# 0.045555f
C411 source.n217 a_n1992_n2088# 0.03241f
C412 source.n218 a_n1992_n2088# 0.017416f
C413 source.n219 a_n1992_n2088# 0.041164f
C414 source.n220 a_n1992_n2088# 0.01844f
C415 source.n221 a_n1992_n2088# 0.03241f
C416 source.n222 a_n1992_n2088# 0.017416f
C417 source.n223 a_n1992_n2088# 0.041164f
C418 source.n224 a_n1992_n2088# 0.01844f
C419 source.n225 a_n1992_n2088# 0.138691f
C420 source.t38 a_n1992_n2088# 0.067092f
C421 source.n226 a_n1992_n2088# 0.030873f
C422 source.n227 a_n1992_n2088# 0.024315f
C423 source.n228 a_n1992_n2088# 0.017416f
C424 source.n229 a_n1992_n2088# 0.771158f
C425 source.n230 a_n1992_n2088# 0.03241f
C426 source.n231 a_n1992_n2088# 0.017416f
C427 source.n232 a_n1992_n2088# 0.01844f
C428 source.n233 a_n1992_n2088# 0.041164f
C429 source.n234 a_n1992_n2088# 0.041164f
C430 source.n235 a_n1992_n2088# 0.01844f
C431 source.n236 a_n1992_n2088# 0.017416f
C432 source.n237 a_n1992_n2088# 0.03241f
C433 source.n238 a_n1992_n2088# 0.03241f
C434 source.n239 a_n1992_n2088# 0.017416f
C435 source.n240 a_n1992_n2088# 0.01844f
C436 source.n241 a_n1992_n2088# 0.041164f
C437 source.n242 a_n1992_n2088# 0.089113f
C438 source.n243 a_n1992_n2088# 0.01844f
C439 source.n244 a_n1992_n2088# 0.017416f
C440 source.n245 a_n1992_n2088# 0.074914f
C441 source.n246 a_n1992_n2088# 0.049862f
C442 source.n247 a_n1992_n2088# 0.128961f
C443 source.t4 a_n1992_n2088# 0.153667f
C444 source.t15 a_n1992_n2088# 0.153667f
C445 source.n248 a_n1992_n2088# 1.19676f
C446 source.n249 a_n1992_n2088# 0.40825f
C447 source.t16 a_n1992_n2088# 0.153667f
C448 source.t6 a_n1992_n2088# 0.153667f
C449 source.n250 a_n1992_n2088# 1.19676f
C450 source.n251 a_n1992_n2088# 0.40825f
C451 source.t9 a_n1992_n2088# 0.153667f
C452 source.t5 a_n1992_n2088# 0.153667f
C453 source.n252 a_n1992_n2088# 1.19676f
C454 source.n253 a_n1992_n2088# 0.40825f
C455 source.t7 a_n1992_n2088# 0.153667f
C456 source.t13 a_n1992_n2088# 0.153667f
C457 source.n254 a_n1992_n2088# 1.19676f
C458 source.n255 a_n1992_n2088# 0.40825f
C459 source.n256 a_n1992_n2088# 0.045555f
C460 source.n257 a_n1992_n2088# 0.03241f
C461 source.n258 a_n1992_n2088# 0.017416f
C462 source.n259 a_n1992_n2088# 0.041164f
C463 source.n260 a_n1992_n2088# 0.01844f
C464 source.n261 a_n1992_n2088# 0.03241f
C465 source.n262 a_n1992_n2088# 0.017416f
C466 source.n263 a_n1992_n2088# 0.041164f
C467 source.n264 a_n1992_n2088# 0.01844f
C468 source.n265 a_n1992_n2088# 0.138691f
C469 source.t0 a_n1992_n2088# 0.067092f
C470 source.n266 a_n1992_n2088# 0.030873f
C471 source.n267 a_n1992_n2088# 0.024315f
C472 source.n268 a_n1992_n2088# 0.017416f
C473 source.n269 a_n1992_n2088# 0.771158f
C474 source.n270 a_n1992_n2088# 0.03241f
C475 source.n271 a_n1992_n2088# 0.017416f
C476 source.n272 a_n1992_n2088# 0.01844f
C477 source.n273 a_n1992_n2088# 0.041164f
C478 source.n274 a_n1992_n2088# 0.041164f
C479 source.n275 a_n1992_n2088# 0.01844f
C480 source.n276 a_n1992_n2088# 0.017416f
C481 source.n277 a_n1992_n2088# 0.03241f
C482 source.n278 a_n1992_n2088# 0.03241f
C483 source.n279 a_n1992_n2088# 0.017416f
C484 source.n280 a_n1992_n2088# 0.01844f
C485 source.n281 a_n1992_n2088# 0.041164f
C486 source.n282 a_n1992_n2088# 0.089113f
C487 source.n283 a_n1992_n2088# 0.01844f
C488 source.n284 a_n1992_n2088# 0.017416f
C489 source.n285 a_n1992_n2088# 0.074914f
C490 source.n286 a_n1992_n2088# 0.049862f
C491 source.n287 a_n1992_n2088# 0.30831f
C492 source.n288 a_n1992_n2088# 1.32397f
C493 plus.n0 a_n1992_n2088# 0.052188f
C494 plus.t15 a_n1992_n2088# 0.223038f
C495 plus.t4 a_n1992_n2088# 0.223038f
C496 plus.t11 a_n1992_n2088# 0.223038f
C497 plus.n1 a_n1992_n2088# 0.10506f
C498 plus.n2 a_n1992_n2088# 0.052188f
C499 plus.t18 a_n1992_n2088# 0.223038f
C500 plus.t12 a_n1992_n2088# 0.223038f
C501 plus.n3 a_n1992_n2088# 0.10506f
C502 plus.n4 a_n1992_n2088# 0.052188f
C503 plus.t0 a_n1992_n2088# 0.223038f
C504 plus.t13 a_n1992_n2088# 0.223038f
C505 plus.t1 a_n1992_n2088# 0.223038f
C506 plus.n5 a_n1992_n2088# 0.10506f
C507 plus.t5 a_n1992_n2088# 0.230589f
C508 plus.n6 a_n1992_n2088# 0.121014f
C509 plus.n7 a_n1992_n2088# 0.119419f
C510 plus.n8 a_n1992_n2088# 0.019886f
C511 plus.n9 a_n1992_n2088# 0.10506f
C512 plus.n10 a_n1992_n2088# 0.019886f
C513 plus.n11 a_n1992_n2088# 0.10506f
C514 plus.n12 a_n1992_n2088# 0.019886f
C515 plus.n13 a_n1992_n2088# 0.052188f
C516 plus.n14 a_n1992_n2088# 0.052188f
C517 plus.n15 a_n1992_n2088# 0.0186f
C518 plus.n16 a_n1992_n2088# 0.0186f
C519 plus.n17 a_n1992_n2088# 0.10506f
C520 plus.n18 a_n1992_n2088# 0.019886f
C521 plus.n19 a_n1992_n2088# 0.052188f
C522 plus.n20 a_n1992_n2088# 0.052188f
C523 plus.n21 a_n1992_n2088# 0.019886f
C524 plus.n22 a_n1992_n2088# 0.10506f
C525 plus.n23 a_n1992_n2088# 0.019886f
C526 plus.n24 a_n1992_n2088# 0.10506f
C527 plus.t3 a_n1992_n2088# 0.230589f
C528 plus.n25 a_n1992_n2088# 0.120935f
C529 plus.n26 a_n1992_n2088# 0.446773f
C530 plus.n27 a_n1992_n2088# 0.052188f
C531 plus.t6 a_n1992_n2088# 0.230589f
C532 plus.t9 a_n1992_n2088# 0.223038f
C533 plus.t19 a_n1992_n2088# 0.223038f
C534 plus.t7 a_n1992_n2088# 0.223038f
C535 plus.n28 a_n1992_n2088# 0.10506f
C536 plus.n29 a_n1992_n2088# 0.052188f
C537 plus.t10 a_n1992_n2088# 0.223038f
C538 plus.t17 a_n1992_n2088# 0.223038f
C539 plus.n30 a_n1992_n2088# 0.10506f
C540 plus.n31 a_n1992_n2088# 0.052188f
C541 plus.t16 a_n1992_n2088# 0.223038f
C542 plus.t2 a_n1992_n2088# 0.223038f
C543 plus.t8 a_n1992_n2088# 0.223038f
C544 plus.n32 a_n1992_n2088# 0.10506f
C545 plus.t14 a_n1992_n2088# 0.230589f
C546 plus.n33 a_n1992_n2088# 0.121014f
C547 plus.n34 a_n1992_n2088# 0.119419f
C548 plus.n35 a_n1992_n2088# 0.019886f
C549 plus.n36 a_n1992_n2088# 0.10506f
C550 plus.n37 a_n1992_n2088# 0.019886f
C551 plus.n38 a_n1992_n2088# 0.10506f
C552 plus.n39 a_n1992_n2088# 0.019886f
C553 plus.n40 a_n1992_n2088# 0.052188f
C554 plus.n41 a_n1992_n2088# 0.052188f
C555 plus.n42 a_n1992_n2088# 0.0186f
C556 plus.n43 a_n1992_n2088# 0.0186f
C557 plus.n44 a_n1992_n2088# 0.10506f
C558 plus.n45 a_n1992_n2088# 0.019886f
C559 plus.n46 a_n1992_n2088# 0.052188f
C560 plus.n47 a_n1992_n2088# 0.052188f
C561 plus.n48 a_n1992_n2088# 0.019886f
C562 plus.n49 a_n1992_n2088# 0.10506f
C563 plus.n50 a_n1992_n2088# 0.019886f
C564 plus.n51 a_n1992_n2088# 0.10506f
C565 plus.n52 a_n1992_n2088# 0.120935f
C566 plus.n53 a_n1992_n2088# 1.3751f
.ends

