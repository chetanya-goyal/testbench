* NGSPICE file created from diffpair417.ext - technology: sky130A

.subckt diffpair417 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t25 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X1 drain_right.t14 minus.t1 source.t15 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X2 source.t27 minus.t2 drain_right.t13 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X3 source.t26 minus.t3 drain_right.t12 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X4 a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X5 source.t13 plus.t0 drain_left.t15 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X6 drain_left.t14 plus.t1 source.t6 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X7 drain_right.t11 minus.t4 source.t28 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X8 drain_right.t10 minus.t5 source.t23 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X9 a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X10 drain_right.t9 minus.t6 source.t24 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X11 drain_right.t8 minus.t7 source.t19 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X12 source.t16 minus.t8 drain_right.t7 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X13 source.t14 minus.t9 drain_right.t6 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X14 source.t29 minus.t10 drain_right.t5 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X15 drain_left.t13 plus.t2 source.t5 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X16 source.t30 plus.t3 drain_left.t12 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X17 source.t22 minus.t11 drain_right.t4 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X18 a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X19 drain_right.t3 minus.t12 source.t21 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X20 drain_right.t2 minus.t13 source.t18 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X21 source.t31 plus.t4 drain_left.t11 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X22 source.t3 plus.t5 drain_left.t10 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X23 source.t12 plus.t6 drain_left.t9 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X24 source.t1 plus.t7 drain_left.t8 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X25 drain_left.t7 plus.t8 source.t8 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X26 drain_left.t6 plus.t9 source.t10 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X27 drain_left.t5 plus.t10 source.t4 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X28 drain_left.t4 plus.t11 source.t7 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X29 source.t20 minus.t14 drain_right.t1 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X30 source.t17 minus.t15 drain_right.t0 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X31 drain_left.t3 plus.t12 source.t9 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X32 a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X33 drain_left.t2 plus.t13 source.t0 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X34 source.t11 plus.t14 drain_left.t1 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X35 source.t2 plus.t15 drain_left.t0 a_n1670_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 minus.n17 minus.t15 1654.5
R1 minus.n4 minus.t12 1654.5
R2 minus.n36 minus.t6 1654.5
R3 minus.n23 minus.t3 1654.5
R4 minus.n16 minus.t1 1602.65
R5 minus.n14 minus.t8 1602.65
R6 minus.n1 minus.t13 1602.65
R7 minus.n9 minus.t14 1602.65
R8 minus.n7 minus.t0 1602.65
R9 minus.n3 minus.t9 1602.65
R10 minus.n35 minus.t10 1602.65
R11 minus.n33 minus.t7 1602.65
R12 minus.n20 minus.t11 1602.65
R13 minus.n28 minus.t4 1602.65
R14 minus.n26 minus.t2 1602.65
R15 minus.n22 minus.t5 1602.65
R16 minus.n5 minus.n4 161.489
R17 minus.n24 minus.n23 161.489
R18 minus.n18 minus.n17 161.3
R19 minus.n15 minus.n0 161.3
R20 minus.n13 minus.n12 161.3
R21 minus.n11 minus.n10 161.3
R22 minus.n8 minus.n2 161.3
R23 minus.n6 minus.n5 161.3
R24 minus.n37 minus.n36 161.3
R25 minus.n34 minus.n19 161.3
R26 minus.n32 minus.n31 161.3
R27 minus.n30 minus.n29 161.3
R28 minus.n27 minus.n21 161.3
R29 minus.n25 minus.n24 161.3
R30 minus.n16 minus.n15 47.4702
R31 minus.n6 minus.n3 47.4702
R32 minus.n25 minus.n22 47.4702
R33 minus.n35 minus.n34 47.4702
R34 minus.n14 minus.n13 43.0884
R35 minus.n8 minus.n7 43.0884
R36 minus.n27 minus.n26 43.0884
R37 minus.n33 minus.n32 43.0884
R38 minus.n10 minus.n1 38.7066
R39 minus.n10 minus.n9 38.7066
R40 minus.n29 minus.n28 38.7066
R41 minus.n29 minus.n20 38.7066
R42 minus.n38 minus.n18 35.4134
R43 minus.n13 minus.n1 34.3247
R44 minus.n9 minus.n8 34.3247
R45 minus.n28 minus.n27 34.3247
R46 minus.n32 minus.n20 34.3247
R47 minus.n15 minus.n14 29.9429
R48 minus.n7 minus.n6 29.9429
R49 minus.n26 minus.n25 29.9429
R50 minus.n34 minus.n33 29.9429
R51 minus.n17 minus.n16 25.5611
R52 minus.n4 minus.n3 25.5611
R53 minus.n23 minus.n22 25.5611
R54 minus.n36 minus.n35 25.5611
R55 minus.n38 minus.n37 6.46641
R56 minus.n18 minus.n0 0.189894
R57 minus.n12 minus.n0 0.189894
R58 minus.n12 minus.n11 0.189894
R59 minus.n11 minus.n2 0.189894
R60 minus.n5 minus.n2 0.189894
R61 minus.n24 minus.n21 0.189894
R62 minus.n30 minus.n21 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n19 0.189894
R65 minus.n37 minus.n19 0.189894
R66 minus minus.n38 0.188
R67 source.n546 source.n486 289.615
R68 source.n474 source.n414 289.615
R69 source.n408 source.n348 289.615
R70 source.n336 source.n276 289.615
R71 source.n60 source.n0 289.615
R72 source.n132 source.n72 289.615
R73 source.n198 source.n138 289.615
R74 source.n270 source.n210 289.615
R75 source.n506 source.n505 185
R76 source.n511 source.n510 185
R77 source.n513 source.n512 185
R78 source.n502 source.n501 185
R79 source.n519 source.n518 185
R80 source.n521 source.n520 185
R81 source.n498 source.n497 185
R82 source.n528 source.n527 185
R83 source.n529 source.n496 185
R84 source.n531 source.n530 185
R85 source.n494 source.n493 185
R86 source.n537 source.n536 185
R87 source.n539 source.n538 185
R88 source.n490 source.n489 185
R89 source.n545 source.n544 185
R90 source.n547 source.n546 185
R91 source.n434 source.n433 185
R92 source.n439 source.n438 185
R93 source.n441 source.n440 185
R94 source.n430 source.n429 185
R95 source.n447 source.n446 185
R96 source.n449 source.n448 185
R97 source.n426 source.n425 185
R98 source.n456 source.n455 185
R99 source.n457 source.n424 185
R100 source.n459 source.n458 185
R101 source.n422 source.n421 185
R102 source.n465 source.n464 185
R103 source.n467 source.n466 185
R104 source.n418 source.n417 185
R105 source.n473 source.n472 185
R106 source.n475 source.n474 185
R107 source.n368 source.n367 185
R108 source.n373 source.n372 185
R109 source.n375 source.n374 185
R110 source.n364 source.n363 185
R111 source.n381 source.n380 185
R112 source.n383 source.n382 185
R113 source.n360 source.n359 185
R114 source.n390 source.n389 185
R115 source.n391 source.n358 185
R116 source.n393 source.n392 185
R117 source.n356 source.n355 185
R118 source.n399 source.n398 185
R119 source.n401 source.n400 185
R120 source.n352 source.n351 185
R121 source.n407 source.n406 185
R122 source.n409 source.n408 185
R123 source.n296 source.n295 185
R124 source.n301 source.n300 185
R125 source.n303 source.n302 185
R126 source.n292 source.n291 185
R127 source.n309 source.n308 185
R128 source.n311 source.n310 185
R129 source.n288 source.n287 185
R130 source.n318 source.n317 185
R131 source.n319 source.n286 185
R132 source.n321 source.n320 185
R133 source.n284 source.n283 185
R134 source.n327 source.n326 185
R135 source.n329 source.n328 185
R136 source.n280 source.n279 185
R137 source.n335 source.n334 185
R138 source.n337 source.n336 185
R139 source.n61 source.n60 185
R140 source.n59 source.n58 185
R141 source.n4 source.n3 185
R142 source.n53 source.n52 185
R143 source.n51 source.n50 185
R144 source.n8 source.n7 185
R145 source.n45 source.n44 185
R146 source.n43 source.n10 185
R147 source.n42 source.n41 185
R148 source.n13 source.n11 185
R149 source.n36 source.n35 185
R150 source.n34 source.n33 185
R151 source.n17 source.n16 185
R152 source.n28 source.n27 185
R153 source.n26 source.n25 185
R154 source.n21 source.n20 185
R155 source.n133 source.n132 185
R156 source.n131 source.n130 185
R157 source.n76 source.n75 185
R158 source.n125 source.n124 185
R159 source.n123 source.n122 185
R160 source.n80 source.n79 185
R161 source.n117 source.n116 185
R162 source.n115 source.n82 185
R163 source.n114 source.n113 185
R164 source.n85 source.n83 185
R165 source.n108 source.n107 185
R166 source.n106 source.n105 185
R167 source.n89 source.n88 185
R168 source.n100 source.n99 185
R169 source.n98 source.n97 185
R170 source.n93 source.n92 185
R171 source.n199 source.n198 185
R172 source.n197 source.n196 185
R173 source.n142 source.n141 185
R174 source.n191 source.n190 185
R175 source.n189 source.n188 185
R176 source.n146 source.n145 185
R177 source.n183 source.n182 185
R178 source.n181 source.n148 185
R179 source.n180 source.n179 185
R180 source.n151 source.n149 185
R181 source.n174 source.n173 185
R182 source.n172 source.n171 185
R183 source.n155 source.n154 185
R184 source.n166 source.n165 185
R185 source.n164 source.n163 185
R186 source.n159 source.n158 185
R187 source.n271 source.n270 185
R188 source.n269 source.n268 185
R189 source.n214 source.n213 185
R190 source.n263 source.n262 185
R191 source.n261 source.n260 185
R192 source.n218 source.n217 185
R193 source.n255 source.n254 185
R194 source.n253 source.n220 185
R195 source.n252 source.n251 185
R196 source.n223 source.n221 185
R197 source.n246 source.n245 185
R198 source.n244 source.n243 185
R199 source.n227 source.n226 185
R200 source.n238 source.n237 185
R201 source.n236 source.n235 185
R202 source.n231 source.n230 185
R203 source.n507 source.t24 149.524
R204 source.n435 source.t26 149.524
R205 source.n369 source.t9 149.524
R206 source.n297 source.t3 149.524
R207 source.n22 source.t0 149.524
R208 source.n94 source.t30 149.524
R209 source.n160 source.t21 149.524
R210 source.n232 source.t17 149.524
R211 source.n511 source.n505 104.615
R212 source.n512 source.n511 104.615
R213 source.n512 source.n501 104.615
R214 source.n519 source.n501 104.615
R215 source.n520 source.n519 104.615
R216 source.n520 source.n497 104.615
R217 source.n528 source.n497 104.615
R218 source.n529 source.n528 104.615
R219 source.n530 source.n529 104.615
R220 source.n530 source.n493 104.615
R221 source.n537 source.n493 104.615
R222 source.n538 source.n537 104.615
R223 source.n538 source.n489 104.615
R224 source.n545 source.n489 104.615
R225 source.n546 source.n545 104.615
R226 source.n439 source.n433 104.615
R227 source.n440 source.n439 104.615
R228 source.n440 source.n429 104.615
R229 source.n447 source.n429 104.615
R230 source.n448 source.n447 104.615
R231 source.n448 source.n425 104.615
R232 source.n456 source.n425 104.615
R233 source.n457 source.n456 104.615
R234 source.n458 source.n457 104.615
R235 source.n458 source.n421 104.615
R236 source.n465 source.n421 104.615
R237 source.n466 source.n465 104.615
R238 source.n466 source.n417 104.615
R239 source.n473 source.n417 104.615
R240 source.n474 source.n473 104.615
R241 source.n373 source.n367 104.615
R242 source.n374 source.n373 104.615
R243 source.n374 source.n363 104.615
R244 source.n381 source.n363 104.615
R245 source.n382 source.n381 104.615
R246 source.n382 source.n359 104.615
R247 source.n390 source.n359 104.615
R248 source.n391 source.n390 104.615
R249 source.n392 source.n391 104.615
R250 source.n392 source.n355 104.615
R251 source.n399 source.n355 104.615
R252 source.n400 source.n399 104.615
R253 source.n400 source.n351 104.615
R254 source.n407 source.n351 104.615
R255 source.n408 source.n407 104.615
R256 source.n301 source.n295 104.615
R257 source.n302 source.n301 104.615
R258 source.n302 source.n291 104.615
R259 source.n309 source.n291 104.615
R260 source.n310 source.n309 104.615
R261 source.n310 source.n287 104.615
R262 source.n318 source.n287 104.615
R263 source.n319 source.n318 104.615
R264 source.n320 source.n319 104.615
R265 source.n320 source.n283 104.615
R266 source.n327 source.n283 104.615
R267 source.n328 source.n327 104.615
R268 source.n328 source.n279 104.615
R269 source.n335 source.n279 104.615
R270 source.n336 source.n335 104.615
R271 source.n60 source.n59 104.615
R272 source.n59 source.n3 104.615
R273 source.n52 source.n3 104.615
R274 source.n52 source.n51 104.615
R275 source.n51 source.n7 104.615
R276 source.n44 source.n7 104.615
R277 source.n44 source.n43 104.615
R278 source.n43 source.n42 104.615
R279 source.n42 source.n11 104.615
R280 source.n35 source.n11 104.615
R281 source.n35 source.n34 104.615
R282 source.n34 source.n16 104.615
R283 source.n27 source.n16 104.615
R284 source.n27 source.n26 104.615
R285 source.n26 source.n20 104.615
R286 source.n132 source.n131 104.615
R287 source.n131 source.n75 104.615
R288 source.n124 source.n75 104.615
R289 source.n124 source.n123 104.615
R290 source.n123 source.n79 104.615
R291 source.n116 source.n79 104.615
R292 source.n116 source.n115 104.615
R293 source.n115 source.n114 104.615
R294 source.n114 source.n83 104.615
R295 source.n107 source.n83 104.615
R296 source.n107 source.n106 104.615
R297 source.n106 source.n88 104.615
R298 source.n99 source.n88 104.615
R299 source.n99 source.n98 104.615
R300 source.n98 source.n92 104.615
R301 source.n198 source.n197 104.615
R302 source.n197 source.n141 104.615
R303 source.n190 source.n141 104.615
R304 source.n190 source.n189 104.615
R305 source.n189 source.n145 104.615
R306 source.n182 source.n145 104.615
R307 source.n182 source.n181 104.615
R308 source.n181 source.n180 104.615
R309 source.n180 source.n149 104.615
R310 source.n173 source.n149 104.615
R311 source.n173 source.n172 104.615
R312 source.n172 source.n154 104.615
R313 source.n165 source.n154 104.615
R314 source.n165 source.n164 104.615
R315 source.n164 source.n158 104.615
R316 source.n270 source.n269 104.615
R317 source.n269 source.n213 104.615
R318 source.n262 source.n213 104.615
R319 source.n262 source.n261 104.615
R320 source.n261 source.n217 104.615
R321 source.n254 source.n217 104.615
R322 source.n254 source.n253 104.615
R323 source.n253 source.n252 104.615
R324 source.n252 source.n221 104.615
R325 source.n245 source.n221 104.615
R326 source.n245 source.n244 104.615
R327 source.n244 source.n226 104.615
R328 source.n237 source.n226 104.615
R329 source.n237 source.n236 104.615
R330 source.n236 source.n230 104.615
R331 source.t24 source.n505 52.3082
R332 source.t26 source.n433 52.3082
R333 source.t9 source.n367 52.3082
R334 source.t3 source.n295 52.3082
R335 source.t0 source.n20 52.3082
R336 source.t30 source.n92 52.3082
R337 source.t21 source.n158 52.3082
R338 source.t17 source.n230 52.3082
R339 source.n67 source.n66 42.8739
R340 source.n69 source.n68 42.8739
R341 source.n71 source.n70 42.8739
R342 source.n205 source.n204 42.8739
R343 source.n207 source.n206 42.8739
R344 source.n209 source.n208 42.8739
R345 source.n485 source.n484 42.8737
R346 source.n483 source.n482 42.8737
R347 source.n481 source.n480 42.8737
R348 source.n347 source.n346 42.8737
R349 source.n345 source.n344 42.8737
R350 source.n343 source.n342 42.8737
R351 source.n551 source.n550 29.8581
R352 source.n479 source.n478 29.8581
R353 source.n413 source.n412 29.8581
R354 source.n341 source.n340 29.8581
R355 source.n65 source.n64 29.8581
R356 source.n137 source.n136 29.8581
R357 source.n203 source.n202 29.8581
R358 source.n275 source.n274 29.8581
R359 source.n341 source.n275 21.7446
R360 source.n552 source.n65 16.2532
R361 source.n531 source.n496 13.1884
R362 source.n459 source.n424 13.1884
R363 source.n393 source.n358 13.1884
R364 source.n321 source.n286 13.1884
R365 source.n45 source.n10 13.1884
R366 source.n117 source.n82 13.1884
R367 source.n183 source.n148 13.1884
R368 source.n255 source.n220 13.1884
R369 source.n527 source.n526 12.8005
R370 source.n532 source.n494 12.8005
R371 source.n455 source.n454 12.8005
R372 source.n460 source.n422 12.8005
R373 source.n389 source.n388 12.8005
R374 source.n394 source.n356 12.8005
R375 source.n317 source.n316 12.8005
R376 source.n322 source.n284 12.8005
R377 source.n46 source.n8 12.8005
R378 source.n41 source.n12 12.8005
R379 source.n118 source.n80 12.8005
R380 source.n113 source.n84 12.8005
R381 source.n184 source.n146 12.8005
R382 source.n179 source.n150 12.8005
R383 source.n256 source.n218 12.8005
R384 source.n251 source.n222 12.8005
R385 source.n525 source.n498 12.0247
R386 source.n536 source.n535 12.0247
R387 source.n453 source.n426 12.0247
R388 source.n464 source.n463 12.0247
R389 source.n387 source.n360 12.0247
R390 source.n398 source.n397 12.0247
R391 source.n315 source.n288 12.0247
R392 source.n326 source.n325 12.0247
R393 source.n50 source.n49 12.0247
R394 source.n40 source.n13 12.0247
R395 source.n122 source.n121 12.0247
R396 source.n112 source.n85 12.0247
R397 source.n188 source.n187 12.0247
R398 source.n178 source.n151 12.0247
R399 source.n260 source.n259 12.0247
R400 source.n250 source.n223 12.0247
R401 source.n522 source.n521 11.249
R402 source.n539 source.n492 11.249
R403 source.n450 source.n449 11.249
R404 source.n467 source.n420 11.249
R405 source.n384 source.n383 11.249
R406 source.n401 source.n354 11.249
R407 source.n312 source.n311 11.249
R408 source.n329 source.n282 11.249
R409 source.n53 source.n6 11.249
R410 source.n37 source.n36 11.249
R411 source.n125 source.n78 11.249
R412 source.n109 source.n108 11.249
R413 source.n191 source.n144 11.249
R414 source.n175 source.n174 11.249
R415 source.n263 source.n216 11.249
R416 source.n247 source.n246 11.249
R417 source.n518 source.n500 10.4732
R418 source.n540 source.n490 10.4732
R419 source.n446 source.n428 10.4732
R420 source.n468 source.n418 10.4732
R421 source.n380 source.n362 10.4732
R422 source.n402 source.n352 10.4732
R423 source.n308 source.n290 10.4732
R424 source.n330 source.n280 10.4732
R425 source.n54 source.n4 10.4732
R426 source.n33 source.n15 10.4732
R427 source.n126 source.n76 10.4732
R428 source.n105 source.n87 10.4732
R429 source.n192 source.n142 10.4732
R430 source.n171 source.n153 10.4732
R431 source.n264 source.n214 10.4732
R432 source.n243 source.n225 10.4732
R433 source.n507 source.n506 10.2747
R434 source.n435 source.n434 10.2747
R435 source.n369 source.n368 10.2747
R436 source.n297 source.n296 10.2747
R437 source.n22 source.n21 10.2747
R438 source.n94 source.n93 10.2747
R439 source.n160 source.n159 10.2747
R440 source.n232 source.n231 10.2747
R441 source.n517 source.n502 9.69747
R442 source.n544 source.n543 9.69747
R443 source.n445 source.n430 9.69747
R444 source.n472 source.n471 9.69747
R445 source.n379 source.n364 9.69747
R446 source.n406 source.n405 9.69747
R447 source.n307 source.n292 9.69747
R448 source.n334 source.n333 9.69747
R449 source.n58 source.n57 9.69747
R450 source.n32 source.n17 9.69747
R451 source.n130 source.n129 9.69747
R452 source.n104 source.n89 9.69747
R453 source.n196 source.n195 9.69747
R454 source.n170 source.n155 9.69747
R455 source.n268 source.n267 9.69747
R456 source.n242 source.n227 9.69747
R457 source.n550 source.n549 9.45567
R458 source.n478 source.n477 9.45567
R459 source.n412 source.n411 9.45567
R460 source.n340 source.n339 9.45567
R461 source.n64 source.n63 9.45567
R462 source.n136 source.n135 9.45567
R463 source.n202 source.n201 9.45567
R464 source.n274 source.n273 9.45567
R465 source.n549 source.n548 9.3005
R466 source.n488 source.n487 9.3005
R467 source.n543 source.n542 9.3005
R468 source.n541 source.n540 9.3005
R469 source.n492 source.n491 9.3005
R470 source.n535 source.n534 9.3005
R471 source.n533 source.n532 9.3005
R472 source.n509 source.n508 9.3005
R473 source.n504 source.n503 9.3005
R474 source.n515 source.n514 9.3005
R475 source.n517 source.n516 9.3005
R476 source.n500 source.n499 9.3005
R477 source.n523 source.n522 9.3005
R478 source.n525 source.n524 9.3005
R479 source.n526 source.n495 9.3005
R480 source.n477 source.n476 9.3005
R481 source.n416 source.n415 9.3005
R482 source.n471 source.n470 9.3005
R483 source.n469 source.n468 9.3005
R484 source.n420 source.n419 9.3005
R485 source.n463 source.n462 9.3005
R486 source.n461 source.n460 9.3005
R487 source.n437 source.n436 9.3005
R488 source.n432 source.n431 9.3005
R489 source.n443 source.n442 9.3005
R490 source.n445 source.n444 9.3005
R491 source.n428 source.n427 9.3005
R492 source.n451 source.n450 9.3005
R493 source.n453 source.n452 9.3005
R494 source.n454 source.n423 9.3005
R495 source.n411 source.n410 9.3005
R496 source.n350 source.n349 9.3005
R497 source.n405 source.n404 9.3005
R498 source.n403 source.n402 9.3005
R499 source.n354 source.n353 9.3005
R500 source.n397 source.n396 9.3005
R501 source.n395 source.n394 9.3005
R502 source.n371 source.n370 9.3005
R503 source.n366 source.n365 9.3005
R504 source.n377 source.n376 9.3005
R505 source.n379 source.n378 9.3005
R506 source.n362 source.n361 9.3005
R507 source.n385 source.n384 9.3005
R508 source.n387 source.n386 9.3005
R509 source.n388 source.n357 9.3005
R510 source.n339 source.n338 9.3005
R511 source.n278 source.n277 9.3005
R512 source.n333 source.n332 9.3005
R513 source.n331 source.n330 9.3005
R514 source.n282 source.n281 9.3005
R515 source.n325 source.n324 9.3005
R516 source.n323 source.n322 9.3005
R517 source.n299 source.n298 9.3005
R518 source.n294 source.n293 9.3005
R519 source.n305 source.n304 9.3005
R520 source.n307 source.n306 9.3005
R521 source.n290 source.n289 9.3005
R522 source.n313 source.n312 9.3005
R523 source.n315 source.n314 9.3005
R524 source.n316 source.n285 9.3005
R525 source.n24 source.n23 9.3005
R526 source.n19 source.n18 9.3005
R527 source.n30 source.n29 9.3005
R528 source.n32 source.n31 9.3005
R529 source.n15 source.n14 9.3005
R530 source.n38 source.n37 9.3005
R531 source.n40 source.n39 9.3005
R532 source.n12 source.n9 9.3005
R533 source.n63 source.n62 9.3005
R534 source.n2 source.n1 9.3005
R535 source.n57 source.n56 9.3005
R536 source.n55 source.n54 9.3005
R537 source.n6 source.n5 9.3005
R538 source.n49 source.n48 9.3005
R539 source.n47 source.n46 9.3005
R540 source.n96 source.n95 9.3005
R541 source.n91 source.n90 9.3005
R542 source.n102 source.n101 9.3005
R543 source.n104 source.n103 9.3005
R544 source.n87 source.n86 9.3005
R545 source.n110 source.n109 9.3005
R546 source.n112 source.n111 9.3005
R547 source.n84 source.n81 9.3005
R548 source.n135 source.n134 9.3005
R549 source.n74 source.n73 9.3005
R550 source.n129 source.n128 9.3005
R551 source.n127 source.n126 9.3005
R552 source.n78 source.n77 9.3005
R553 source.n121 source.n120 9.3005
R554 source.n119 source.n118 9.3005
R555 source.n162 source.n161 9.3005
R556 source.n157 source.n156 9.3005
R557 source.n168 source.n167 9.3005
R558 source.n170 source.n169 9.3005
R559 source.n153 source.n152 9.3005
R560 source.n176 source.n175 9.3005
R561 source.n178 source.n177 9.3005
R562 source.n150 source.n147 9.3005
R563 source.n201 source.n200 9.3005
R564 source.n140 source.n139 9.3005
R565 source.n195 source.n194 9.3005
R566 source.n193 source.n192 9.3005
R567 source.n144 source.n143 9.3005
R568 source.n187 source.n186 9.3005
R569 source.n185 source.n184 9.3005
R570 source.n234 source.n233 9.3005
R571 source.n229 source.n228 9.3005
R572 source.n240 source.n239 9.3005
R573 source.n242 source.n241 9.3005
R574 source.n225 source.n224 9.3005
R575 source.n248 source.n247 9.3005
R576 source.n250 source.n249 9.3005
R577 source.n222 source.n219 9.3005
R578 source.n273 source.n272 9.3005
R579 source.n212 source.n211 9.3005
R580 source.n267 source.n266 9.3005
R581 source.n265 source.n264 9.3005
R582 source.n216 source.n215 9.3005
R583 source.n259 source.n258 9.3005
R584 source.n257 source.n256 9.3005
R585 source.n514 source.n513 8.92171
R586 source.n547 source.n488 8.92171
R587 source.n442 source.n441 8.92171
R588 source.n475 source.n416 8.92171
R589 source.n376 source.n375 8.92171
R590 source.n409 source.n350 8.92171
R591 source.n304 source.n303 8.92171
R592 source.n337 source.n278 8.92171
R593 source.n61 source.n2 8.92171
R594 source.n29 source.n28 8.92171
R595 source.n133 source.n74 8.92171
R596 source.n101 source.n100 8.92171
R597 source.n199 source.n140 8.92171
R598 source.n167 source.n166 8.92171
R599 source.n271 source.n212 8.92171
R600 source.n239 source.n238 8.92171
R601 source.n510 source.n504 8.14595
R602 source.n548 source.n486 8.14595
R603 source.n438 source.n432 8.14595
R604 source.n476 source.n414 8.14595
R605 source.n372 source.n366 8.14595
R606 source.n410 source.n348 8.14595
R607 source.n300 source.n294 8.14595
R608 source.n338 source.n276 8.14595
R609 source.n62 source.n0 8.14595
R610 source.n25 source.n19 8.14595
R611 source.n134 source.n72 8.14595
R612 source.n97 source.n91 8.14595
R613 source.n200 source.n138 8.14595
R614 source.n163 source.n157 8.14595
R615 source.n272 source.n210 8.14595
R616 source.n235 source.n229 8.14595
R617 source.n509 source.n506 7.3702
R618 source.n437 source.n434 7.3702
R619 source.n371 source.n368 7.3702
R620 source.n299 source.n296 7.3702
R621 source.n24 source.n21 7.3702
R622 source.n96 source.n93 7.3702
R623 source.n162 source.n159 7.3702
R624 source.n234 source.n231 7.3702
R625 source.n510 source.n509 5.81868
R626 source.n550 source.n486 5.81868
R627 source.n438 source.n437 5.81868
R628 source.n478 source.n414 5.81868
R629 source.n372 source.n371 5.81868
R630 source.n412 source.n348 5.81868
R631 source.n300 source.n299 5.81868
R632 source.n340 source.n276 5.81868
R633 source.n64 source.n0 5.81868
R634 source.n25 source.n24 5.81868
R635 source.n136 source.n72 5.81868
R636 source.n97 source.n96 5.81868
R637 source.n202 source.n138 5.81868
R638 source.n163 source.n162 5.81868
R639 source.n274 source.n210 5.81868
R640 source.n235 source.n234 5.81868
R641 source.n552 source.n551 5.49188
R642 source.n513 source.n504 5.04292
R643 source.n548 source.n547 5.04292
R644 source.n441 source.n432 5.04292
R645 source.n476 source.n475 5.04292
R646 source.n375 source.n366 5.04292
R647 source.n410 source.n409 5.04292
R648 source.n303 source.n294 5.04292
R649 source.n338 source.n337 5.04292
R650 source.n62 source.n61 5.04292
R651 source.n28 source.n19 5.04292
R652 source.n134 source.n133 5.04292
R653 source.n100 source.n91 5.04292
R654 source.n200 source.n199 5.04292
R655 source.n166 source.n157 5.04292
R656 source.n272 source.n271 5.04292
R657 source.n238 source.n229 5.04292
R658 source.n514 source.n502 4.26717
R659 source.n544 source.n488 4.26717
R660 source.n442 source.n430 4.26717
R661 source.n472 source.n416 4.26717
R662 source.n376 source.n364 4.26717
R663 source.n406 source.n350 4.26717
R664 source.n304 source.n292 4.26717
R665 source.n334 source.n278 4.26717
R666 source.n58 source.n2 4.26717
R667 source.n29 source.n17 4.26717
R668 source.n130 source.n74 4.26717
R669 source.n101 source.n89 4.26717
R670 source.n196 source.n140 4.26717
R671 source.n167 source.n155 4.26717
R672 source.n268 source.n212 4.26717
R673 source.n239 source.n227 4.26717
R674 source.n518 source.n517 3.49141
R675 source.n543 source.n490 3.49141
R676 source.n446 source.n445 3.49141
R677 source.n471 source.n418 3.49141
R678 source.n380 source.n379 3.49141
R679 source.n405 source.n352 3.49141
R680 source.n308 source.n307 3.49141
R681 source.n333 source.n280 3.49141
R682 source.n57 source.n4 3.49141
R683 source.n33 source.n32 3.49141
R684 source.n129 source.n76 3.49141
R685 source.n105 source.n104 3.49141
R686 source.n195 source.n142 3.49141
R687 source.n171 source.n170 3.49141
R688 source.n267 source.n214 3.49141
R689 source.n243 source.n242 3.49141
R690 source.n508 source.n507 2.84303
R691 source.n436 source.n435 2.84303
R692 source.n370 source.n369 2.84303
R693 source.n298 source.n297 2.84303
R694 source.n23 source.n22 2.84303
R695 source.n95 source.n94 2.84303
R696 source.n161 source.n160 2.84303
R697 source.n233 source.n232 2.84303
R698 source.n521 source.n500 2.71565
R699 source.n540 source.n539 2.71565
R700 source.n449 source.n428 2.71565
R701 source.n468 source.n467 2.71565
R702 source.n383 source.n362 2.71565
R703 source.n402 source.n401 2.71565
R704 source.n311 source.n290 2.71565
R705 source.n330 source.n329 2.71565
R706 source.n54 source.n53 2.71565
R707 source.n36 source.n15 2.71565
R708 source.n126 source.n125 2.71565
R709 source.n108 source.n87 2.71565
R710 source.n192 source.n191 2.71565
R711 source.n174 source.n153 2.71565
R712 source.n264 source.n263 2.71565
R713 source.n246 source.n225 2.71565
R714 source.n522 source.n498 1.93989
R715 source.n536 source.n492 1.93989
R716 source.n450 source.n426 1.93989
R717 source.n464 source.n420 1.93989
R718 source.n384 source.n360 1.93989
R719 source.n398 source.n354 1.93989
R720 source.n312 source.n288 1.93989
R721 source.n326 source.n282 1.93989
R722 source.n50 source.n6 1.93989
R723 source.n37 source.n13 1.93989
R724 source.n122 source.n78 1.93989
R725 source.n109 source.n85 1.93989
R726 source.n188 source.n144 1.93989
R727 source.n175 source.n151 1.93989
R728 source.n260 source.n216 1.93989
R729 source.n247 source.n223 1.93989
R730 source.n484 source.t19 1.6505
R731 source.n484 source.t29 1.6505
R732 source.n482 source.t28 1.6505
R733 source.n482 source.t22 1.6505
R734 source.n480 source.t23 1.6505
R735 source.n480 source.t27 1.6505
R736 source.n346 source.t4 1.6505
R737 source.n346 source.t2 1.6505
R738 source.n344 source.t7 1.6505
R739 source.n344 source.t12 1.6505
R740 source.n342 source.t10 1.6505
R741 source.n342 source.t31 1.6505
R742 source.n66 source.t5 1.6505
R743 source.n66 source.t13 1.6505
R744 source.n68 source.t8 1.6505
R745 source.n68 source.t1 1.6505
R746 source.n70 source.t6 1.6505
R747 source.n70 source.t11 1.6505
R748 source.n204 source.t25 1.6505
R749 source.n204 source.t14 1.6505
R750 source.n206 source.t18 1.6505
R751 source.n206 source.t20 1.6505
R752 source.n208 source.t15 1.6505
R753 source.n208 source.t16 1.6505
R754 source.n527 source.n525 1.16414
R755 source.n535 source.n494 1.16414
R756 source.n455 source.n453 1.16414
R757 source.n463 source.n422 1.16414
R758 source.n389 source.n387 1.16414
R759 source.n397 source.n356 1.16414
R760 source.n317 source.n315 1.16414
R761 source.n325 source.n284 1.16414
R762 source.n49 source.n8 1.16414
R763 source.n41 source.n40 1.16414
R764 source.n121 source.n80 1.16414
R765 source.n113 source.n112 1.16414
R766 source.n187 source.n146 1.16414
R767 source.n179 source.n178 1.16414
R768 source.n259 source.n218 1.16414
R769 source.n251 source.n250 1.16414
R770 source.n203 source.n137 0.470328
R771 source.n479 source.n413 0.470328
R772 source.n275 source.n209 0.457397
R773 source.n209 source.n207 0.457397
R774 source.n207 source.n205 0.457397
R775 source.n205 source.n203 0.457397
R776 source.n137 source.n71 0.457397
R777 source.n71 source.n69 0.457397
R778 source.n69 source.n67 0.457397
R779 source.n67 source.n65 0.457397
R780 source.n343 source.n341 0.457397
R781 source.n345 source.n343 0.457397
R782 source.n347 source.n345 0.457397
R783 source.n413 source.n347 0.457397
R784 source.n481 source.n479 0.457397
R785 source.n483 source.n481 0.457397
R786 source.n485 source.n483 0.457397
R787 source.n551 source.n485 0.457397
R788 source.n526 source.n496 0.388379
R789 source.n532 source.n531 0.388379
R790 source.n454 source.n424 0.388379
R791 source.n460 source.n459 0.388379
R792 source.n388 source.n358 0.388379
R793 source.n394 source.n393 0.388379
R794 source.n316 source.n286 0.388379
R795 source.n322 source.n321 0.388379
R796 source.n46 source.n45 0.388379
R797 source.n12 source.n10 0.388379
R798 source.n118 source.n117 0.388379
R799 source.n84 source.n82 0.388379
R800 source.n184 source.n183 0.388379
R801 source.n150 source.n148 0.388379
R802 source.n256 source.n255 0.388379
R803 source.n222 source.n220 0.388379
R804 source source.n552 0.188
R805 source.n508 source.n503 0.155672
R806 source.n515 source.n503 0.155672
R807 source.n516 source.n515 0.155672
R808 source.n516 source.n499 0.155672
R809 source.n523 source.n499 0.155672
R810 source.n524 source.n523 0.155672
R811 source.n524 source.n495 0.155672
R812 source.n533 source.n495 0.155672
R813 source.n534 source.n533 0.155672
R814 source.n534 source.n491 0.155672
R815 source.n541 source.n491 0.155672
R816 source.n542 source.n541 0.155672
R817 source.n542 source.n487 0.155672
R818 source.n549 source.n487 0.155672
R819 source.n436 source.n431 0.155672
R820 source.n443 source.n431 0.155672
R821 source.n444 source.n443 0.155672
R822 source.n444 source.n427 0.155672
R823 source.n451 source.n427 0.155672
R824 source.n452 source.n451 0.155672
R825 source.n452 source.n423 0.155672
R826 source.n461 source.n423 0.155672
R827 source.n462 source.n461 0.155672
R828 source.n462 source.n419 0.155672
R829 source.n469 source.n419 0.155672
R830 source.n470 source.n469 0.155672
R831 source.n470 source.n415 0.155672
R832 source.n477 source.n415 0.155672
R833 source.n370 source.n365 0.155672
R834 source.n377 source.n365 0.155672
R835 source.n378 source.n377 0.155672
R836 source.n378 source.n361 0.155672
R837 source.n385 source.n361 0.155672
R838 source.n386 source.n385 0.155672
R839 source.n386 source.n357 0.155672
R840 source.n395 source.n357 0.155672
R841 source.n396 source.n395 0.155672
R842 source.n396 source.n353 0.155672
R843 source.n403 source.n353 0.155672
R844 source.n404 source.n403 0.155672
R845 source.n404 source.n349 0.155672
R846 source.n411 source.n349 0.155672
R847 source.n298 source.n293 0.155672
R848 source.n305 source.n293 0.155672
R849 source.n306 source.n305 0.155672
R850 source.n306 source.n289 0.155672
R851 source.n313 source.n289 0.155672
R852 source.n314 source.n313 0.155672
R853 source.n314 source.n285 0.155672
R854 source.n323 source.n285 0.155672
R855 source.n324 source.n323 0.155672
R856 source.n324 source.n281 0.155672
R857 source.n331 source.n281 0.155672
R858 source.n332 source.n331 0.155672
R859 source.n332 source.n277 0.155672
R860 source.n339 source.n277 0.155672
R861 source.n63 source.n1 0.155672
R862 source.n56 source.n1 0.155672
R863 source.n56 source.n55 0.155672
R864 source.n55 source.n5 0.155672
R865 source.n48 source.n5 0.155672
R866 source.n48 source.n47 0.155672
R867 source.n47 source.n9 0.155672
R868 source.n39 source.n9 0.155672
R869 source.n39 source.n38 0.155672
R870 source.n38 source.n14 0.155672
R871 source.n31 source.n14 0.155672
R872 source.n31 source.n30 0.155672
R873 source.n30 source.n18 0.155672
R874 source.n23 source.n18 0.155672
R875 source.n135 source.n73 0.155672
R876 source.n128 source.n73 0.155672
R877 source.n128 source.n127 0.155672
R878 source.n127 source.n77 0.155672
R879 source.n120 source.n77 0.155672
R880 source.n120 source.n119 0.155672
R881 source.n119 source.n81 0.155672
R882 source.n111 source.n81 0.155672
R883 source.n111 source.n110 0.155672
R884 source.n110 source.n86 0.155672
R885 source.n103 source.n86 0.155672
R886 source.n103 source.n102 0.155672
R887 source.n102 source.n90 0.155672
R888 source.n95 source.n90 0.155672
R889 source.n201 source.n139 0.155672
R890 source.n194 source.n139 0.155672
R891 source.n194 source.n193 0.155672
R892 source.n193 source.n143 0.155672
R893 source.n186 source.n143 0.155672
R894 source.n186 source.n185 0.155672
R895 source.n185 source.n147 0.155672
R896 source.n177 source.n147 0.155672
R897 source.n177 source.n176 0.155672
R898 source.n176 source.n152 0.155672
R899 source.n169 source.n152 0.155672
R900 source.n169 source.n168 0.155672
R901 source.n168 source.n156 0.155672
R902 source.n161 source.n156 0.155672
R903 source.n273 source.n211 0.155672
R904 source.n266 source.n211 0.155672
R905 source.n266 source.n265 0.155672
R906 source.n265 source.n215 0.155672
R907 source.n258 source.n215 0.155672
R908 source.n258 source.n257 0.155672
R909 source.n257 source.n219 0.155672
R910 source.n249 source.n219 0.155672
R911 source.n249 source.n248 0.155672
R912 source.n248 source.n224 0.155672
R913 source.n241 source.n224 0.155672
R914 source.n241 source.n240 0.155672
R915 source.n240 source.n228 0.155672
R916 source.n233 source.n228 0.155672
R917 drain_right.n5 drain_right.n3 60.0094
R918 drain_right.n2 drain_right.n0 60.0094
R919 drain_right.n9 drain_right.n7 60.0094
R920 drain_right.n9 drain_right.n8 59.5527
R921 drain_right.n11 drain_right.n10 59.5527
R922 drain_right.n13 drain_right.n12 59.5527
R923 drain_right.n5 drain_right.n4 59.5525
R924 drain_right.n2 drain_right.n1 59.5525
R925 drain_right drain_right.n6 29.7837
R926 drain_right drain_right.n13 6.11011
R927 drain_right.n3 drain_right.t5 1.6505
R928 drain_right.n3 drain_right.t9 1.6505
R929 drain_right.n4 drain_right.t4 1.6505
R930 drain_right.n4 drain_right.t8 1.6505
R931 drain_right.n1 drain_right.t13 1.6505
R932 drain_right.n1 drain_right.t11 1.6505
R933 drain_right.n0 drain_right.t12 1.6505
R934 drain_right.n0 drain_right.t10 1.6505
R935 drain_right.n7 drain_right.t6 1.6505
R936 drain_right.n7 drain_right.t3 1.6505
R937 drain_right.n8 drain_right.t1 1.6505
R938 drain_right.n8 drain_right.t15 1.6505
R939 drain_right.n10 drain_right.t7 1.6505
R940 drain_right.n10 drain_right.t2 1.6505
R941 drain_right.n12 drain_right.t0 1.6505
R942 drain_right.n12 drain_right.t14 1.6505
R943 drain_right.n13 drain_right.n11 0.457397
R944 drain_right.n11 drain_right.n9 0.457397
R945 drain_right.n6 drain_right.n5 0.173602
R946 drain_right.n6 drain_right.n2 0.173602
R947 plus.n4 plus.t3 1654.5
R948 plus.n17 plus.t13 1654.5
R949 plus.n23 plus.t12 1654.5
R950 plus.n36 plus.t5 1654.5
R951 plus.n3 plus.t1 1602.65
R952 plus.n7 plus.t14 1602.65
R953 plus.n9 plus.t8 1602.65
R954 plus.n1 plus.t7 1602.65
R955 plus.n14 plus.t2 1602.65
R956 plus.n16 plus.t0 1602.65
R957 plus.n22 plus.t15 1602.65
R958 plus.n26 plus.t10 1602.65
R959 plus.n28 plus.t6 1602.65
R960 plus.n20 plus.t11 1602.65
R961 plus.n33 plus.t4 1602.65
R962 plus.n35 plus.t9 1602.65
R963 plus.n5 plus.n4 161.489
R964 plus.n24 plus.n23 161.489
R965 plus.n6 plus.n5 161.3
R966 plus.n8 plus.n2 161.3
R967 plus.n11 plus.n10 161.3
R968 plus.n13 plus.n12 161.3
R969 plus.n15 plus.n0 161.3
R970 plus.n18 plus.n17 161.3
R971 plus.n25 plus.n24 161.3
R972 plus.n27 plus.n21 161.3
R973 plus.n30 plus.n29 161.3
R974 plus.n32 plus.n31 161.3
R975 plus.n34 plus.n19 161.3
R976 plus.n37 plus.n36 161.3
R977 plus.n6 plus.n3 47.4702
R978 plus.n16 plus.n15 47.4702
R979 plus.n35 plus.n34 47.4702
R980 plus.n25 plus.n22 47.4702
R981 plus.n8 plus.n7 43.0884
R982 plus.n14 plus.n13 43.0884
R983 plus.n33 plus.n32 43.0884
R984 plus.n27 plus.n26 43.0884
R985 plus.n10 plus.n9 38.7066
R986 plus.n10 plus.n1 38.7066
R987 plus.n29 plus.n20 38.7066
R988 plus.n29 plus.n28 38.7066
R989 plus.n9 plus.n8 34.3247
R990 plus.n13 plus.n1 34.3247
R991 plus.n32 plus.n20 34.3247
R992 plus.n28 plus.n27 34.3247
R993 plus.n7 plus.n6 29.9429
R994 plus.n15 plus.n14 29.9429
R995 plus.n34 plus.n33 29.9429
R996 plus.n26 plus.n25 29.9429
R997 plus plus.n37 29.2945
R998 plus.n4 plus.n3 25.5611
R999 plus.n17 plus.n16 25.5611
R1000 plus.n36 plus.n35 25.5611
R1001 plus.n23 plus.n22 25.5611
R1002 plus plus.n18 12.1103
R1003 plus.n5 plus.n2 0.189894
R1004 plus.n11 plus.n2 0.189894
R1005 plus.n12 plus.n11 0.189894
R1006 plus.n12 plus.n0 0.189894
R1007 plus.n18 plus.n0 0.189894
R1008 plus.n37 plus.n19 0.189894
R1009 plus.n31 plus.n19 0.189894
R1010 plus.n31 plus.n30 0.189894
R1011 plus.n30 plus.n21 0.189894
R1012 plus.n24 plus.n21 0.189894
R1013 drain_left.n9 drain_left.n7 60.0096
R1014 drain_left.n5 drain_left.n3 60.0094
R1015 drain_left.n2 drain_left.n0 60.0094
R1016 drain_left.n11 drain_left.n10 59.5527
R1017 drain_left.n9 drain_left.n8 59.5527
R1018 drain_left.n5 drain_left.n4 59.5525
R1019 drain_left.n2 drain_left.n1 59.5525
R1020 drain_left.n13 drain_left.n12 59.5525
R1021 drain_left drain_left.n6 30.3369
R1022 drain_left drain_left.n13 6.11011
R1023 drain_left.n3 drain_left.t0 1.6505
R1024 drain_left.n3 drain_left.t3 1.6505
R1025 drain_left.n4 drain_left.t9 1.6505
R1026 drain_left.n4 drain_left.t5 1.6505
R1027 drain_left.n1 drain_left.t11 1.6505
R1028 drain_left.n1 drain_left.t4 1.6505
R1029 drain_left.n0 drain_left.t10 1.6505
R1030 drain_left.n0 drain_left.t6 1.6505
R1031 drain_left.n12 drain_left.t15 1.6505
R1032 drain_left.n12 drain_left.t2 1.6505
R1033 drain_left.n10 drain_left.t8 1.6505
R1034 drain_left.n10 drain_left.t13 1.6505
R1035 drain_left.n8 drain_left.t1 1.6505
R1036 drain_left.n8 drain_left.t7 1.6505
R1037 drain_left.n7 drain_left.t12 1.6505
R1038 drain_left.n7 drain_left.t14 1.6505
R1039 drain_left.n11 drain_left.n9 0.457397
R1040 drain_left.n13 drain_left.n11 0.457397
R1041 drain_left.n6 drain_left.n5 0.173602
R1042 drain_left.n6 drain_left.n2 0.173602
C0 drain_right minus 4.42496f
C1 drain_left source 36.6909f
C2 plus source 4.0303f
C3 drain_left plus 4.58593f
C4 source minus 4.01626f
C5 drain_right source 36.6906f
C6 drain_left minus 0.170856f
C7 drain_right drain_left 0.846053f
C8 plus minus 5.23723f
C9 drain_right plus 0.314737f
C10 drain_right a_n1670_n3288# 6.78189f
C11 drain_left a_n1670_n3288# 7.05679f
C12 source a_n1670_n3288# 8.541806f
C13 minus a_n1670_n3288# 6.472262f
C14 plus a_n1670_n3288# 8.53483f
C15 drain_left.t10 a_n1670_n3288# 0.366405f
C16 drain_left.t6 a_n1670_n3288# 0.366405f
C17 drain_left.n0 a_n1670_n3288# 3.26389f
C18 drain_left.t11 a_n1670_n3288# 0.366405f
C19 drain_left.t4 a_n1670_n3288# 0.366405f
C20 drain_left.n1 a_n1670_n3288# 3.26044f
C21 drain_left.n2 a_n1670_n3288# 0.858053f
C22 drain_left.t0 a_n1670_n3288# 0.366405f
C23 drain_left.t3 a_n1670_n3288# 0.366405f
C24 drain_left.n3 a_n1670_n3288# 3.26389f
C25 drain_left.t9 a_n1670_n3288# 0.366405f
C26 drain_left.t5 a_n1670_n3288# 0.366405f
C27 drain_left.n4 a_n1670_n3288# 3.26044f
C28 drain_left.n5 a_n1670_n3288# 0.858053f
C29 drain_left.n6 a_n1670_n3288# 1.81155f
C30 drain_left.t12 a_n1670_n3288# 0.366405f
C31 drain_left.t14 a_n1670_n3288# 0.366405f
C32 drain_left.n7 a_n1670_n3288# 3.26391f
C33 drain_left.t1 a_n1670_n3288# 0.366405f
C34 drain_left.t7 a_n1670_n3288# 0.366405f
C35 drain_left.n8 a_n1670_n3288# 3.26045f
C36 drain_left.n9 a_n1670_n3288# 0.888185f
C37 drain_left.t8 a_n1670_n3288# 0.366405f
C38 drain_left.t13 a_n1670_n3288# 0.366405f
C39 drain_left.n10 a_n1670_n3288# 3.26045f
C40 drain_left.n11 a_n1670_n3288# 0.438038f
C41 drain_left.t15 a_n1670_n3288# 0.366405f
C42 drain_left.t2 a_n1670_n3288# 0.366405f
C43 drain_left.n12 a_n1670_n3288# 3.26044f
C44 drain_left.n13 a_n1670_n3288# 0.754275f
C45 plus.n0 a_n1670_n3288# 0.054862f
C46 plus.t0 a_n1670_n3288# 0.372075f
C47 plus.t2 a_n1670_n3288# 0.372075f
C48 plus.t7 a_n1670_n3288# 0.372075f
C49 plus.n1 a_n1670_n3288# 0.153237f
C50 plus.n2 a_n1670_n3288# 0.054862f
C51 plus.t8 a_n1670_n3288# 0.372075f
C52 plus.t14 a_n1670_n3288# 0.372075f
C53 plus.t1 a_n1670_n3288# 0.372075f
C54 plus.n3 a_n1670_n3288# 0.153237f
C55 plus.t3 a_n1670_n3288# 0.376936f
C56 plus.n4 a_n1670_n3288# 0.169532f
C57 plus.n5 a_n1670_n3288# 0.123512f
C58 plus.n6 a_n1670_n3288# 0.019214f
C59 plus.n7 a_n1670_n3288# 0.153237f
C60 plus.n8 a_n1670_n3288# 0.019214f
C61 plus.n9 a_n1670_n3288# 0.153237f
C62 plus.n10 a_n1670_n3288# 0.019214f
C63 plus.n11 a_n1670_n3288# 0.054862f
C64 plus.n12 a_n1670_n3288# 0.054862f
C65 plus.n13 a_n1670_n3288# 0.019214f
C66 plus.n14 a_n1670_n3288# 0.153237f
C67 plus.n15 a_n1670_n3288# 0.019214f
C68 plus.n16 a_n1670_n3288# 0.153237f
C69 plus.t13 a_n1670_n3288# 0.376936f
C70 plus.n17 a_n1670_n3288# 0.169452f
C71 plus.n18 a_n1670_n3288# 0.609416f
C72 plus.n19 a_n1670_n3288# 0.054862f
C73 plus.t5 a_n1670_n3288# 0.376936f
C74 plus.t9 a_n1670_n3288# 0.372075f
C75 plus.t4 a_n1670_n3288# 0.372075f
C76 plus.t11 a_n1670_n3288# 0.372075f
C77 plus.n20 a_n1670_n3288# 0.153237f
C78 plus.n21 a_n1670_n3288# 0.054862f
C79 plus.t6 a_n1670_n3288# 0.372075f
C80 plus.t10 a_n1670_n3288# 0.372075f
C81 plus.t15 a_n1670_n3288# 0.372075f
C82 plus.n22 a_n1670_n3288# 0.153237f
C83 plus.t12 a_n1670_n3288# 0.376936f
C84 plus.n23 a_n1670_n3288# 0.169532f
C85 plus.n24 a_n1670_n3288# 0.123512f
C86 plus.n25 a_n1670_n3288# 0.019214f
C87 plus.n26 a_n1670_n3288# 0.153237f
C88 plus.n27 a_n1670_n3288# 0.019214f
C89 plus.n28 a_n1670_n3288# 0.153237f
C90 plus.n29 a_n1670_n3288# 0.019214f
C91 plus.n30 a_n1670_n3288# 0.054862f
C92 plus.n31 a_n1670_n3288# 0.054862f
C93 plus.n32 a_n1670_n3288# 0.019214f
C94 plus.n33 a_n1670_n3288# 0.153237f
C95 plus.n34 a_n1670_n3288# 0.019214f
C96 plus.n35 a_n1670_n3288# 0.153237f
C97 plus.n36 a_n1670_n3288# 0.169452f
C98 plus.n37 a_n1670_n3288# 1.58025f
C99 drain_right.t12 a_n1670_n3288# 0.36597f
C100 drain_right.t10 a_n1670_n3288# 0.36597f
C101 drain_right.n0 a_n1670_n3288# 3.26002f
C102 drain_right.t13 a_n1670_n3288# 0.36597f
C103 drain_right.t11 a_n1670_n3288# 0.36597f
C104 drain_right.n1 a_n1670_n3288# 3.25657f
C105 drain_right.n2 a_n1670_n3288# 0.857035f
C106 drain_right.t5 a_n1670_n3288# 0.36597f
C107 drain_right.t9 a_n1670_n3288# 0.36597f
C108 drain_right.n3 a_n1670_n3288# 3.26002f
C109 drain_right.t4 a_n1670_n3288# 0.36597f
C110 drain_right.t8 a_n1670_n3288# 0.36597f
C111 drain_right.n4 a_n1670_n3288# 3.25657f
C112 drain_right.n5 a_n1670_n3288# 0.857034f
C113 drain_right.n6 a_n1670_n3288# 1.72912f
C114 drain_right.t6 a_n1670_n3288# 0.36597f
C115 drain_right.t3 a_n1670_n3288# 0.36597f
C116 drain_right.n7 a_n1670_n3288# 3.26002f
C117 drain_right.t1 a_n1670_n3288# 0.36597f
C118 drain_right.t15 a_n1670_n3288# 0.36597f
C119 drain_right.n8 a_n1670_n3288# 3.25658f
C120 drain_right.n9 a_n1670_n3288# 0.887144f
C121 drain_right.t7 a_n1670_n3288# 0.36597f
C122 drain_right.t2 a_n1670_n3288# 0.36597f
C123 drain_right.n10 a_n1670_n3288# 3.25658f
C124 drain_right.n11 a_n1670_n3288# 0.437518f
C125 drain_right.t0 a_n1670_n3288# 0.36597f
C126 drain_right.t14 a_n1670_n3288# 0.36597f
C127 drain_right.n12 a_n1670_n3288# 3.25658f
C128 drain_right.n13 a_n1670_n3288# 0.753367f
C129 source.n0 a_n1670_n3288# 0.0426f
C130 source.n1 a_n1670_n3288# 0.03216f
C131 source.n2 a_n1670_n3288# 0.017282f
C132 source.n3 a_n1670_n3288# 0.040847f
C133 source.n4 a_n1670_n3288# 0.018298f
C134 source.n5 a_n1670_n3288# 0.03216f
C135 source.n6 a_n1670_n3288# 0.017282f
C136 source.n7 a_n1670_n3288# 0.040847f
C137 source.n8 a_n1670_n3288# 0.018298f
C138 source.n9 a_n1670_n3288# 0.03216f
C139 source.n10 a_n1670_n3288# 0.01779f
C140 source.n11 a_n1670_n3288# 0.040847f
C141 source.n12 a_n1670_n3288# 0.017282f
C142 source.n13 a_n1670_n3288# 0.018298f
C143 source.n14 a_n1670_n3288# 0.03216f
C144 source.n15 a_n1670_n3288# 0.017282f
C145 source.n16 a_n1670_n3288# 0.040847f
C146 source.n17 a_n1670_n3288# 0.018298f
C147 source.n18 a_n1670_n3288# 0.03216f
C148 source.n19 a_n1670_n3288# 0.017282f
C149 source.n20 a_n1670_n3288# 0.030636f
C150 source.n21 a_n1670_n3288# 0.028876f
C151 source.t0 a_n1670_n3288# 0.068988f
C152 source.n22 a_n1670_n3288# 0.231872f
C153 source.n23 a_n1670_n3288# 1.62243f
C154 source.n24 a_n1670_n3288# 0.017282f
C155 source.n25 a_n1670_n3288# 0.018298f
C156 source.n26 a_n1670_n3288# 0.040847f
C157 source.n27 a_n1670_n3288# 0.040847f
C158 source.n28 a_n1670_n3288# 0.018298f
C159 source.n29 a_n1670_n3288# 0.017282f
C160 source.n30 a_n1670_n3288# 0.03216f
C161 source.n31 a_n1670_n3288# 0.03216f
C162 source.n32 a_n1670_n3288# 0.017282f
C163 source.n33 a_n1670_n3288# 0.018298f
C164 source.n34 a_n1670_n3288# 0.040847f
C165 source.n35 a_n1670_n3288# 0.040847f
C166 source.n36 a_n1670_n3288# 0.018298f
C167 source.n37 a_n1670_n3288# 0.017282f
C168 source.n38 a_n1670_n3288# 0.03216f
C169 source.n39 a_n1670_n3288# 0.03216f
C170 source.n40 a_n1670_n3288# 0.017282f
C171 source.n41 a_n1670_n3288# 0.018298f
C172 source.n42 a_n1670_n3288# 0.040847f
C173 source.n43 a_n1670_n3288# 0.040847f
C174 source.n44 a_n1670_n3288# 0.040847f
C175 source.n45 a_n1670_n3288# 0.01779f
C176 source.n46 a_n1670_n3288# 0.017282f
C177 source.n47 a_n1670_n3288# 0.03216f
C178 source.n48 a_n1670_n3288# 0.03216f
C179 source.n49 a_n1670_n3288# 0.017282f
C180 source.n50 a_n1670_n3288# 0.018298f
C181 source.n51 a_n1670_n3288# 0.040847f
C182 source.n52 a_n1670_n3288# 0.040847f
C183 source.n53 a_n1670_n3288# 0.018298f
C184 source.n54 a_n1670_n3288# 0.017282f
C185 source.n55 a_n1670_n3288# 0.03216f
C186 source.n56 a_n1670_n3288# 0.03216f
C187 source.n57 a_n1670_n3288# 0.017282f
C188 source.n58 a_n1670_n3288# 0.018298f
C189 source.n59 a_n1670_n3288# 0.040847f
C190 source.n60 a_n1670_n3288# 0.083823f
C191 source.n61 a_n1670_n3288# 0.018298f
C192 source.n62 a_n1670_n3288# 0.017282f
C193 source.n63 a_n1670_n3288# 0.069065f
C194 source.n64 a_n1670_n3288# 0.046261f
C195 source.n65 a_n1670_n3288# 1.27963f
C196 source.t5 a_n1670_n3288# 0.304969f
C197 source.t13 a_n1670_n3288# 0.304969f
C198 source.n66 a_n1670_n3288# 2.61115f
C199 source.n67 a_n1670_n3288# 0.423493f
C200 source.t8 a_n1670_n3288# 0.304969f
C201 source.t1 a_n1670_n3288# 0.304969f
C202 source.n68 a_n1670_n3288# 2.61115f
C203 source.n69 a_n1670_n3288# 0.423493f
C204 source.t6 a_n1670_n3288# 0.304969f
C205 source.t11 a_n1670_n3288# 0.304969f
C206 source.n70 a_n1670_n3288# 2.61115f
C207 source.n71 a_n1670_n3288# 0.423493f
C208 source.n72 a_n1670_n3288# 0.0426f
C209 source.n73 a_n1670_n3288# 0.03216f
C210 source.n74 a_n1670_n3288# 0.017282f
C211 source.n75 a_n1670_n3288# 0.040847f
C212 source.n76 a_n1670_n3288# 0.018298f
C213 source.n77 a_n1670_n3288# 0.03216f
C214 source.n78 a_n1670_n3288# 0.017282f
C215 source.n79 a_n1670_n3288# 0.040847f
C216 source.n80 a_n1670_n3288# 0.018298f
C217 source.n81 a_n1670_n3288# 0.03216f
C218 source.n82 a_n1670_n3288# 0.01779f
C219 source.n83 a_n1670_n3288# 0.040847f
C220 source.n84 a_n1670_n3288# 0.017282f
C221 source.n85 a_n1670_n3288# 0.018298f
C222 source.n86 a_n1670_n3288# 0.03216f
C223 source.n87 a_n1670_n3288# 0.017282f
C224 source.n88 a_n1670_n3288# 0.040847f
C225 source.n89 a_n1670_n3288# 0.018298f
C226 source.n90 a_n1670_n3288# 0.03216f
C227 source.n91 a_n1670_n3288# 0.017282f
C228 source.n92 a_n1670_n3288# 0.030636f
C229 source.n93 a_n1670_n3288# 0.028876f
C230 source.t30 a_n1670_n3288# 0.068988f
C231 source.n94 a_n1670_n3288# 0.231872f
C232 source.n95 a_n1670_n3288# 1.62243f
C233 source.n96 a_n1670_n3288# 0.017282f
C234 source.n97 a_n1670_n3288# 0.018298f
C235 source.n98 a_n1670_n3288# 0.040847f
C236 source.n99 a_n1670_n3288# 0.040847f
C237 source.n100 a_n1670_n3288# 0.018298f
C238 source.n101 a_n1670_n3288# 0.017282f
C239 source.n102 a_n1670_n3288# 0.03216f
C240 source.n103 a_n1670_n3288# 0.03216f
C241 source.n104 a_n1670_n3288# 0.017282f
C242 source.n105 a_n1670_n3288# 0.018298f
C243 source.n106 a_n1670_n3288# 0.040847f
C244 source.n107 a_n1670_n3288# 0.040847f
C245 source.n108 a_n1670_n3288# 0.018298f
C246 source.n109 a_n1670_n3288# 0.017282f
C247 source.n110 a_n1670_n3288# 0.03216f
C248 source.n111 a_n1670_n3288# 0.03216f
C249 source.n112 a_n1670_n3288# 0.017282f
C250 source.n113 a_n1670_n3288# 0.018298f
C251 source.n114 a_n1670_n3288# 0.040847f
C252 source.n115 a_n1670_n3288# 0.040847f
C253 source.n116 a_n1670_n3288# 0.040847f
C254 source.n117 a_n1670_n3288# 0.01779f
C255 source.n118 a_n1670_n3288# 0.017282f
C256 source.n119 a_n1670_n3288# 0.03216f
C257 source.n120 a_n1670_n3288# 0.03216f
C258 source.n121 a_n1670_n3288# 0.017282f
C259 source.n122 a_n1670_n3288# 0.018298f
C260 source.n123 a_n1670_n3288# 0.040847f
C261 source.n124 a_n1670_n3288# 0.040847f
C262 source.n125 a_n1670_n3288# 0.018298f
C263 source.n126 a_n1670_n3288# 0.017282f
C264 source.n127 a_n1670_n3288# 0.03216f
C265 source.n128 a_n1670_n3288# 0.03216f
C266 source.n129 a_n1670_n3288# 0.017282f
C267 source.n130 a_n1670_n3288# 0.018298f
C268 source.n131 a_n1670_n3288# 0.040847f
C269 source.n132 a_n1670_n3288# 0.083823f
C270 source.n133 a_n1670_n3288# 0.018298f
C271 source.n134 a_n1670_n3288# 0.017282f
C272 source.n135 a_n1670_n3288# 0.069065f
C273 source.n136 a_n1670_n3288# 0.046261f
C274 source.n137 a_n1670_n3288# 0.120532f
C275 source.n138 a_n1670_n3288# 0.0426f
C276 source.n139 a_n1670_n3288# 0.03216f
C277 source.n140 a_n1670_n3288# 0.017282f
C278 source.n141 a_n1670_n3288# 0.040847f
C279 source.n142 a_n1670_n3288# 0.018298f
C280 source.n143 a_n1670_n3288# 0.03216f
C281 source.n144 a_n1670_n3288# 0.017282f
C282 source.n145 a_n1670_n3288# 0.040847f
C283 source.n146 a_n1670_n3288# 0.018298f
C284 source.n147 a_n1670_n3288# 0.03216f
C285 source.n148 a_n1670_n3288# 0.01779f
C286 source.n149 a_n1670_n3288# 0.040847f
C287 source.n150 a_n1670_n3288# 0.017282f
C288 source.n151 a_n1670_n3288# 0.018298f
C289 source.n152 a_n1670_n3288# 0.03216f
C290 source.n153 a_n1670_n3288# 0.017282f
C291 source.n154 a_n1670_n3288# 0.040847f
C292 source.n155 a_n1670_n3288# 0.018298f
C293 source.n156 a_n1670_n3288# 0.03216f
C294 source.n157 a_n1670_n3288# 0.017282f
C295 source.n158 a_n1670_n3288# 0.030636f
C296 source.n159 a_n1670_n3288# 0.028876f
C297 source.t21 a_n1670_n3288# 0.068988f
C298 source.n160 a_n1670_n3288# 0.231872f
C299 source.n161 a_n1670_n3288# 1.62243f
C300 source.n162 a_n1670_n3288# 0.017282f
C301 source.n163 a_n1670_n3288# 0.018298f
C302 source.n164 a_n1670_n3288# 0.040847f
C303 source.n165 a_n1670_n3288# 0.040847f
C304 source.n166 a_n1670_n3288# 0.018298f
C305 source.n167 a_n1670_n3288# 0.017282f
C306 source.n168 a_n1670_n3288# 0.03216f
C307 source.n169 a_n1670_n3288# 0.03216f
C308 source.n170 a_n1670_n3288# 0.017282f
C309 source.n171 a_n1670_n3288# 0.018298f
C310 source.n172 a_n1670_n3288# 0.040847f
C311 source.n173 a_n1670_n3288# 0.040847f
C312 source.n174 a_n1670_n3288# 0.018298f
C313 source.n175 a_n1670_n3288# 0.017282f
C314 source.n176 a_n1670_n3288# 0.03216f
C315 source.n177 a_n1670_n3288# 0.03216f
C316 source.n178 a_n1670_n3288# 0.017282f
C317 source.n179 a_n1670_n3288# 0.018298f
C318 source.n180 a_n1670_n3288# 0.040847f
C319 source.n181 a_n1670_n3288# 0.040847f
C320 source.n182 a_n1670_n3288# 0.040847f
C321 source.n183 a_n1670_n3288# 0.01779f
C322 source.n184 a_n1670_n3288# 0.017282f
C323 source.n185 a_n1670_n3288# 0.03216f
C324 source.n186 a_n1670_n3288# 0.03216f
C325 source.n187 a_n1670_n3288# 0.017282f
C326 source.n188 a_n1670_n3288# 0.018298f
C327 source.n189 a_n1670_n3288# 0.040847f
C328 source.n190 a_n1670_n3288# 0.040847f
C329 source.n191 a_n1670_n3288# 0.018298f
C330 source.n192 a_n1670_n3288# 0.017282f
C331 source.n193 a_n1670_n3288# 0.03216f
C332 source.n194 a_n1670_n3288# 0.03216f
C333 source.n195 a_n1670_n3288# 0.017282f
C334 source.n196 a_n1670_n3288# 0.018298f
C335 source.n197 a_n1670_n3288# 0.040847f
C336 source.n198 a_n1670_n3288# 0.083823f
C337 source.n199 a_n1670_n3288# 0.018298f
C338 source.n200 a_n1670_n3288# 0.017282f
C339 source.n201 a_n1670_n3288# 0.069065f
C340 source.n202 a_n1670_n3288# 0.046261f
C341 source.n203 a_n1670_n3288# 0.120532f
C342 source.t25 a_n1670_n3288# 0.304969f
C343 source.t14 a_n1670_n3288# 0.304969f
C344 source.n204 a_n1670_n3288# 2.61115f
C345 source.n205 a_n1670_n3288# 0.423493f
C346 source.t18 a_n1670_n3288# 0.304969f
C347 source.t20 a_n1670_n3288# 0.304969f
C348 source.n206 a_n1670_n3288# 2.61115f
C349 source.n207 a_n1670_n3288# 0.423493f
C350 source.t15 a_n1670_n3288# 0.304969f
C351 source.t16 a_n1670_n3288# 0.304969f
C352 source.n208 a_n1670_n3288# 2.61115f
C353 source.n209 a_n1670_n3288# 0.423493f
C354 source.n210 a_n1670_n3288# 0.0426f
C355 source.n211 a_n1670_n3288# 0.03216f
C356 source.n212 a_n1670_n3288# 0.017282f
C357 source.n213 a_n1670_n3288# 0.040847f
C358 source.n214 a_n1670_n3288# 0.018298f
C359 source.n215 a_n1670_n3288# 0.03216f
C360 source.n216 a_n1670_n3288# 0.017282f
C361 source.n217 a_n1670_n3288# 0.040847f
C362 source.n218 a_n1670_n3288# 0.018298f
C363 source.n219 a_n1670_n3288# 0.03216f
C364 source.n220 a_n1670_n3288# 0.01779f
C365 source.n221 a_n1670_n3288# 0.040847f
C366 source.n222 a_n1670_n3288# 0.017282f
C367 source.n223 a_n1670_n3288# 0.018298f
C368 source.n224 a_n1670_n3288# 0.03216f
C369 source.n225 a_n1670_n3288# 0.017282f
C370 source.n226 a_n1670_n3288# 0.040847f
C371 source.n227 a_n1670_n3288# 0.018298f
C372 source.n228 a_n1670_n3288# 0.03216f
C373 source.n229 a_n1670_n3288# 0.017282f
C374 source.n230 a_n1670_n3288# 0.030636f
C375 source.n231 a_n1670_n3288# 0.028876f
C376 source.t17 a_n1670_n3288# 0.068988f
C377 source.n232 a_n1670_n3288# 0.231872f
C378 source.n233 a_n1670_n3288# 1.62243f
C379 source.n234 a_n1670_n3288# 0.017282f
C380 source.n235 a_n1670_n3288# 0.018298f
C381 source.n236 a_n1670_n3288# 0.040847f
C382 source.n237 a_n1670_n3288# 0.040847f
C383 source.n238 a_n1670_n3288# 0.018298f
C384 source.n239 a_n1670_n3288# 0.017282f
C385 source.n240 a_n1670_n3288# 0.03216f
C386 source.n241 a_n1670_n3288# 0.03216f
C387 source.n242 a_n1670_n3288# 0.017282f
C388 source.n243 a_n1670_n3288# 0.018298f
C389 source.n244 a_n1670_n3288# 0.040847f
C390 source.n245 a_n1670_n3288# 0.040847f
C391 source.n246 a_n1670_n3288# 0.018298f
C392 source.n247 a_n1670_n3288# 0.017282f
C393 source.n248 a_n1670_n3288# 0.03216f
C394 source.n249 a_n1670_n3288# 0.03216f
C395 source.n250 a_n1670_n3288# 0.017282f
C396 source.n251 a_n1670_n3288# 0.018298f
C397 source.n252 a_n1670_n3288# 0.040847f
C398 source.n253 a_n1670_n3288# 0.040847f
C399 source.n254 a_n1670_n3288# 0.040847f
C400 source.n255 a_n1670_n3288# 0.01779f
C401 source.n256 a_n1670_n3288# 0.017282f
C402 source.n257 a_n1670_n3288# 0.03216f
C403 source.n258 a_n1670_n3288# 0.03216f
C404 source.n259 a_n1670_n3288# 0.017282f
C405 source.n260 a_n1670_n3288# 0.018298f
C406 source.n261 a_n1670_n3288# 0.040847f
C407 source.n262 a_n1670_n3288# 0.040847f
C408 source.n263 a_n1670_n3288# 0.018298f
C409 source.n264 a_n1670_n3288# 0.017282f
C410 source.n265 a_n1670_n3288# 0.03216f
C411 source.n266 a_n1670_n3288# 0.03216f
C412 source.n267 a_n1670_n3288# 0.017282f
C413 source.n268 a_n1670_n3288# 0.018298f
C414 source.n269 a_n1670_n3288# 0.040847f
C415 source.n270 a_n1670_n3288# 0.083823f
C416 source.n271 a_n1670_n3288# 0.018298f
C417 source.n272 a_n1670_n3288# 0.017282f
C418 source.n273 a_n1670_n3288# 0.069065f
C419 source.n274 a_n1670_n3288# 0.046261f
C420 source.n275 a_n1670_n3288# 1.78212f
C421 source.n276 a_n1670_n3288# 0.0426f
C422 source.n277 a_n1670_n3288# 0.03216f
C423 source.n278 a_n1670_n3288# 0.017282f
C424 source.n279 a_n1670_n3288# 0.040847f
C425 source.n280 a_n1670_n3288# 0.018298f
C426 source.n281 a_n1670_n3288# 0.03216f
C427 source.n282 a_n1670_n3288# 0.017282f
C428 source.n283 a_n1670_n3288# 0.040847f
C429 source.n284 a_n1670_n3288# 0.018298f
C430 source.n285 a_n1670_n3288# 0.03216f
C431 source.n286 a_n1670_n3288# 0.01779f
C432 source.n287 a_n1670_n3288# 0.040847f
C433 source.n288 a_n1670_n3288# 0.018298f
C434 source.n289 a_n1670_n3288# 0.03216f
C435 source.n290 a_n1670_n3288# 0.017282f
C436 source.n291 a_n1670_n3288# 0.040847f
C437 source.n292 a_n1670_n3288# 0.018298f
C438 source.n293 a_n1670_n3288# 0.03216f
C439 source.n294 a_n1670_n3288# 0.017282f
C440 source.n295 a_n1670_n3288# 0.030636f
C441 source.n296 a_n1670_n3288# 0.028876f
C442 source.t3 a_n1670_n3288# 0.068988f
C443 source.n297 a_n1670_n3288# 0.231872f
C444 source.n298 a_n1670_n3288# 1.62243f
C445 source.n299 a_n1670_n3288# 0.017282f
C446 source.n300 a_n1670_n3288# 0.018298f
C447 source.n301 a_n1670_n3288# 0.040847f
C448 source.n302 a_n1670_n3288# 0.040847f
C449 source.n303 a_n1670_n3288# 0.018298f
C450 source.n304 a_n1670_n3288# 0.017282f
C451 source.n305 a_n1670_n3288# 0.03216f
C452 source.n306 a_n1670_n3288# 0.03216f
C453 source.n307 a_n1670_n3288# 0.017282f
C454 source.n308 a_n1670_n3288# 0.018298f
C455 source.n309 a_n1670_n3288# 0.040847f
C456 source.n310 a_n1670_n3288# 0.040847f
C457 source.n311 a_n1670_n3288# 0.018298f
C458 source.n312 a_n1670_n3288# 0.017282f
C459 source.n313 a_n1670_n3288# 0.03216f
C460 source.n314 a_n1670_n3288# 0.03216f
C461 source.n315 a_n1670_n3288# 0.017282f
C462 source.n316 a_n1670_n3288# 0.017282f
C463 source.n317 a_n1670_n3288# 0.018298f
C464 source.n318 a_n1670_n3288# 0.040847f
C465 source.n319 a_n1670_n3288# 0.040847f
C466 source.n320 a_n1670_n3288# 0.040847f
C467 source.n321 a_n1670_n3288# 0.01779f
C468 source.n322 a_n1670_n3288# 0.017282f
C469 source.n323 a_n1670_n3288# 0.03216f
C470 source.n324 a_n1670_n3288# 0.03216f
C471 source.n325 a_n1670_n3288# 0.017282f
C472 source.n326 a_n1670_n3288# 0.018298f
C473 source.n327 a_n1670_n3288# 0.040847f
C474 source.n328 a_n1670_n3288# 0.040847f
C475 source.n329 a_n1670_n3288# 0.018298f
C476 source.n330 a_n1670_n3288# 0.017282f
C477 source.n331 a_n1670_n3288# 0.03216f
C478 source.n332 a_n1670_n3288# 0.03216f
C479 source.n333 a_n1670_n3288# 0.017282f
C480 source.n334 a_n1670_n3288# 0.018298f
C481 source.n335 a_n1670_n3288# 0.040847f
C482 source.n336 a_n1670_n3288# 0.083823f
C483 source.n337 a_n1670_n3288# 0.018298f
C484 source.n338 a_n1670_n3288# 0.017282f
C485 source.n339 a_n1670_n3288# 0.069065f
C486 source.n340 a_n1670_n3288# 0.046261f
C487 source.n341 a_n1670_n3288# 1.78212f
C488 source.t10 a_n1670_n3288# 0.304969f
C489 source.t31 a_n1670_n3288# 0.304969f
C490 source.n342 a_n1670_n3288# 2.61113f
C491 source.n343 a_n1670_n3288# 0.423508f
C492 source.t7 a_n1670_n3288# 0.304969f
C493 source.t12 a_n1670_n3288# 0.304969f
C494 source.n344 a_n1670_n3288# 2.61113f
C495 source.n345 a_n1670_n3288# 0.423508f
C496 source.t4 a_n1670_n3288# 0.304969f
C497 source.t2 a_n1670_n3288# 0.304969f
C498 source.n346 a_n1670_n3288# 2.61113f
C499 source.n347 a_n1670_n3288# 0.423508f
C500 source.n348 a_n1670_n3288# 0.0426f
C501 source.n349 a_n1670_n3288# 0.03216f
C502 source.n350 a_n1670_n3288# 0.017282f
C503 source.n351 a_n1670_n3288# 0.040847f
C504 source.n352 a_n1670_n3288# 0.018298f
C505 source.n353 a_n1670_n3288# 0.03216f
C506 source.n354 a_n1670_n3288# 0.017282f
C507 source.n355 a_n1670_n3288# 0.040847f
C508 source.n356 a_n1670_n3288# 0.018298f
C509 source.n357 a_n1670_n3288# 0.03216f
C510 source.n358 a_n1670_n3288# 0.01779f
C511 source.n359 a_n1670_n3288# 0.040847f
C512 source.n360 a_n1670_n3288# 0.018298f
C513 source.n361 a_n1670_n3288# 0.03216f
C514 source.n362 a_n1670_n3288# 0.017282f
C515 source.n363 a_n1670_n3288# 0.040847f
C516 source.n364 a_n1670_n3288# 0.018298f
C517 source.n365 a_n1670_n3288# 0.03216f
C518 source.n366 a_n1670_n3288# 0.017282f
C519 source.n367 a_n1670_n3288# 0.030636f
C520 source.n368 a_n1670_n3288# 0.028876f
C521 source.t9 a_n1670_n3288# 0.068988f
C522 source.n369 a_n1670_n3288# 0.231872f
C523 source.n370 a_n1670_n3288# 1.62243f
C524 source.n371 a_n1670_n3288# 0.017282f
C525 source.n372 a_n1670_n3288# 0.018298f
C526 source.n373 a_n1670_n3288# 0.040847f
C527 source.n374 a_n1670_n3288# 0.040847f
C528 source.n375 a_n1670_n3288# 0.018298f
C529 source.n376 a_n1670_n3288# 0.017282f
C530 source.n377 a_n1670_n3288# 0.03216f
C531 source.n378 a_n1670_n3288# 0.03216f
C532 source.n379 a_n1670_n3288# 0.017282f
C533 source.n380 a_n1670_n3288# 0.018298f
C534 source.n381 a_n1670_n3288# 0.040847f
C535 source.n382 a_n1670_n3288# 0.040847f
C536 source.n383 a_n1670_n3288# 0.018298f
C537 source.n384 a_n1670_n3288# 0.017282f
C538 source.n385 a_n1670_n3288# 0.03216f
C539 source.n386 a_n1670_n3288# 0.03216f
C540 source.n387 a_n1670_n3288# 0.017282f
C541 source.n388 a_n1670_n3288# 0.017282f
C542 source.n389 a_n1670_n3288# 0.018298f
C543 source.n390 a_n1670_n3288# 0.040847f
C544 source.n391 a_n1670_n3288# 0.040847f
C545 source.n392 a_n1670_n3288# 0.040847f
C546 source.n393 a_n1670_n3288# 0.01779f
C547 source.n394 a_n1670_n3288# 0.017282f
C548 source.n395 a_n1670_n3288# 0.03216f
C549 source.n396 a_n1670_n3288# 0.03216f
C550 source.n397 a_n1670_n3288# 0.017282f
C551 source.n398 a_n1670_n3288# 0.018298f
C552 source.n399 a_n1670_n3288# 0.040847f
C553 source.n400 a_n1670_n3288# 0.040847f
C554 source.n401 a_n1670_n3288# 0.018298f
C555 source.n402 a_n1670_n3288# 0.017282f
C556 source.n403 a_n1670_n3288# 0.03216f
C557 source.n404 a_n1670_n3288# 0.03216f
C558 source.n405 a_n1670_n3288# 0.017282f
C559 source.n406 a_n1670_n3288# 0.018298f
C560 source.n407 a_n1670_n3288# 0.040847f
C561 source.n408 a_n1670_n3288# 0.083823f
C562 source.n409 a_n1670_n3288# 0.018298f
C563 source.n410 a_n1670_n3288# 0.017282f
C564 source.n411 a_n1670_n3288# 0.069065f
C565 source.n412 a_n1670_n3288# 0.046261f
C566 source.n413 a_n1670_n3288# 0.120532f
C567 source.n414 a_n1670_n3288# 0.0426f
C568 source.n415 a_n1670_n3288# 0.03216f
C569 source.n416 a_n1670_n3288# 0.017282f
C570 source.n417 a_n1670_n3288# 0.040847f
C571 source.n418 a_n1670_n3288# 0.018298f
C572 source.n419 a_n1670_n3288# 0.03216f
C573 source.n420 a_n1670_n3288# 0.017282f
C574 source.n421 a_n1670_n3288# 0.040847f
C575 source.n422 a_n1670_n3288# 0.018298f
C576 source.n423 a_n1670_n3288# 0.03216f
C577 source.n424 a_n1670_n3288# 0.01779f
C578 source.n425 a_n1670_n3288# 0.040847f
C579 source.n426 a_n1670_n3288# 0.018298f
C580 source.n427 a_n1670_n3288# 0.03216f
C581 source.n428 a_n1670_n3288# 0.017282f
C582 source.n429 a_n1670_n3288# 0.040847f
C583 source.n430 a_n1670_n3288# 0.018298f
C584 source.n431 a_n1670_n3288# 0.03216f
C585 source.n432 a_n1670_n3288# 0.017282f
C586 source.n433 a_n1670_n3288# 0.030636f
C587 source.n434 a_n1670_n3288# 0.028876f
C588 source.t26 a_n1670_n3288# 0.068988f
C589 source.n435 a_n1670_n3288# 0.231872f
C590 source.n436 a_n1670_n3288# 1.62243f
C591 source.n437 a_n1670_n3288# 0.017282f
C592 source.n438 a_n1670_n3288# 0.018298f
C593 source.n439 a_n1670_n3288# 0.040847f
C594 source.n440 a_n1670_n3288# 0.040847f
C595 source.n441 a_n1670_n3288# 0.018298f
C596 source.n442 a_n1670_n3288# 0.017282f
C597 source.n443 a_n1670_n3288# 0.03216f
C598 source.n444 a_n1670_n3288# 0.03216f
C599 source.n445 a_n1670_n3288# 0.017282f
C600 source.n446 a_n1670_n3288# 0.018298f
C601 source.n447 a_n1670_n3288# 0.040847f
C602 source.n448 a_n1670_n3288# 0.040847f
C603 source.n449 a_n1670_n3288# 0.018298f
C604 source.n450 a_n1670_n3288# 0.017282f
C605 source.n451 a_n1670_n3288# 0.03216f
C606 source.n452 a_n1670_n3288# 0.03216f
C607 source.n453 a_n1670_n3288# 0.017282f
C608 source.n454 a_n1670_n3288# 0.017282f
C609 source.n455 a_n1670_n3288# 0.018298f
C610 source.n456 a_n1670_n3288# 0.040847f
C611 source.n457 a_n1670_n3288# 0.040847f
C612 source.n458 a_n1670_n3288# 0.040847f
C613 source.n459 a_n1670_n3288# 0.01779f
C614 source.n460 a_n1670_n3288# 0.017282f
C615 source.n461 a_n1670_n3288# 0.03216f
C616 source.n462 a_n1670_n3288# 0.03216f
C617 source.n463 a_n1670_n3288# 0.017282f
C618 source.n464 a_n1670_n3288# 0.018298f
C619 source.n465 a_n1670_n3288# 0.040847f
C620 source.n466 a_n1670_n3288# 0.040847f
C621 source.n467 a_n1670_n3288# 0.018298f
C622 source.n468 a_n1670_n3288# 0.017282f
C623 source.n469 a_n1670_n3288# 0.03216f
C624 source.n470 a_n1670_n3288# 0.03216f
C625 source.n471 a_n1670_n3288# 0.017282f
C626 source.n472 a_n1670_n3288# 0.018298f
C627 source.n473 a_n1670_n3288# 0.040847f
C628 source.n474 a_n1670_n3288# 0.083823f
C629 source.n475 a_n1670_n3288# 0.018298f
C630 source.n476 a_n1670_n3288# 0.017282f
C631 source.n477 a_n1670_n3288# 0.069065f
C632 source.n478 a_n1670_n3288# 0.046261f
C633 source.n479 a_n1670_n3288# 0.120532f
C634 source.t23 a_n1670_n3288# 0.304969f
C635 source.t27 a_n1670_n3288# 0.304969f
C636 source.n480 a_n1670_n3288# 2.61113f
C637 source.n481 a_n1670_n3288# 0.423508f
C638 source.t28 a_n1670_n3288# 0.304969f
C639 source.t22 a_n1670_n3288# 0.304969f
C640 source.n482 a_n1670_n3288# 2.61113f
C641 source.n483 a_n1670_n3288# 0.423508f
C642 source.t19 a_n1670_n3288# 0.304969f
C643 source.t29 a_n1670_n3288# 0.304969f
C644 source.n484 a_n1670_n3288# 2.61113f
C645 source.n485 a_n1670_n3288# 0.423508f
C646 source.n486 a_n1670_n3288# 0.0426f
C647 source.n487 a_n1670_n3288# 0.03216f
C648 source.n488 a_n1670_n3288# 0.017282f
C649 source.n489 a_n1670_n3288# 0.040847f
C650 source.n490 a_n1670_n3288# 0.018298f
C651 source.n491 a_n1670_n3288# 0.03216f
C652 source.n492 a_n1670_n3288# 0.017282f
C653 source.n493 a_n1670_n3288# 0.040847f
C654 source.n494 a_n1670_n3288# 0.018298f
C655 source.n495 a_n1670_n3288# 0.03216f
C656 source.n496 a_n1670_n3288# 0.01779f
C657 source.n497 a_n1670_n3288# 0.040847f
C658 source.n498 a_n1670_n3288# 0.018298f
C659 source.n499 a_n1670_n3288# 0.03216f
C660 source.n500 a_n1670_n3288# 0.017282f
C661 source.n501 a_n1670_n3288# 0.040847f
C662 source.n502 a_n1670_n3288# 0.018298f
C663 source.n503 a_n1670_n3288# 0.03216f
C664 source.n504 a_n1670_n3288# 0.017282f
C665 source.n505 a_n1670_n3288# 0.030636f
C666 source.n506 a_n1670_n3288# 0.028876f
C667 source.t24 a_n1670_n3288# 0.068988f
C668 source.n507 a_n1670_n3288# 0.231872f
C669 source.n508 a_n1670_n3288# 1.62243f
C670 source.n509 a_n1670_n3288# 0.017282f
C671 source.n510 a_n1670_n3288# 0.018298f
C672 source.n511 a_n1670_n3288# 0.040847f
C673 source.n512 a_n1670_n3288# 0.040847f
C674 source.n513 a_n1670_n3288# 0.018298f
C675 source.n514 a_n1670_n3288# 0.017282f
C676 source.n515 a_n1670_n3288# 0.03216f
C677 source.n516 a_n1670_n3288# 0.03216f
C678 source.n517 a_n1670_n3288# 0.017282f
C679 source.n518 a_n1670_n3288# 0.018298f
C680 source.n519 a_n1670_n3288# 0.040847f
C681 source.n520 a_n1670_n3288# 0.040847f
C682 source.n521 a_n1670_n3288# 0.018298f
C683 source.n522 a_n1670_n3288# 0.017282f
C684 source.n523 a_n1670_n3288# 0.03216f
C685 source.n524 a_n1670_n3288# 0.03216f
C686 source.n525 a_n1670_n3288# 0.017282f
C687 source.n526 a_n1670_n3288# 0.017282f
C688 source.n527 a_n1670_n3288# 0.018298f
C689 source.n528 a_n1670_n3288# 0.040847f
C690 source.n529 a_n1670_n3288# 0.040847f
C691 source.n530 a_n1670_n3288# 0.040847f
C692 source.n531 a_n1670_n3288# 0.01779f
C693 source.n532 a_n1670_n3288# 0.017282f
C694 source.n533 a_n1670_n3288# 0.03216f
C695 source.n534 a_n1670_n3288# 0.03216f
C696 source.n535 a_n1670_n3288# 0.017282f
C697 source.n536 a_n1670_n3288# 0.018298f
C698 source.n537 a_n1670_n3288# 0.040847f
C699 source.n538 a_n1670_n3288# 0.040847f
C700 source.n539 a_n1670_n3288# 0.018298f
C701 source.n540 a_n1670_n3288# 0.017282f
C702 source.n541 a_n1670_n3288# 0.03216f
C703 source.n542 a_n1670_n3288# 0.03216f
C704 source.n543 a_n1670_n3288# 0.017282f
C705 source.n544 a_n1670_n3288# 0.018298f
C706 source.n545 a_n1670_n3288# 0.040847f
C707 source.n546 a_n1670_n3288# 0.083823f
C708 source.n547 a_n1670_n3288# 0.018298f
C709 source.n548 a_n1670_n3288# 0.017282f
C710 source.n549 a_n1670_n3288# 0.069065f
C711 source.n550 a_n1670_n3288# 0.046261f
C712 source.n551 a_n1670_n3288# 0.294915f
C713 source.n552 a_n1670_n3288# 2.01257f
C714 minus.n0 a_n1670_n3288# 0.053636f
C715 minus.t15 a_n1670_n3288# 0.36851f
C716 minus.t1 a_n1670_n3288# 0.363758f
C717 minus.t8 a_n1670_n3288# 0.363758f
C718 minus.t13 a_n1670_n3288# 0.363758f
C719 minus.n1 a_n1670_n3288# 0.149812f
C720 minus.n2 a_n1670_n3288# 0.053636f
C721 minus.t14 a_n1670_n3288# 0.363758f
C722 minus.t0 a_n1670_n3288# 0.363758f
C723 minus.t9 a_n1670_n3288# 0.363758f
C724 minus.n3 a_n1670_n3288# 0.149812f
C725 minus.t12 a_n1670_n3288# 0.36851f
C726 minus.n4 a_n1670_n3288# 0.165743f
C727 minus.n5 a_n1670_n3288# 0.120751f
C728 minus.n6 a_n1670_n3288# 0.018785f
C729 minus.n7 a_n1670_n3288# 0.149812f
C730 minus.n8 a_n1670_n3288# 0.018785f
C731 minus.n9 a_n1670_n3288# 0.149812f
C732 minus.n10 a_n1670_n3288# 0.018785f
C733 minus.n11 a_n1670_n3288# 0.053636f
C734 minus.n12 a_n1670_n3288# 0.053636f
C735 minus.n13 a_n1670_n3288# 0.018785f
C736 minus.n14 a_n1670_n3288# 0.149812f
C737 minus.n15 a_n1670_n3288# 0.018785f
C738 minus.n16 a_n1670_n3288# 0.149812f
C739 minus.n17 a_n1670_n3288# 0.165664f
C740 minus.n18 a_n1670_n3288# 1.83032f
C741 minus.n19 a_n1670_n3288# 0.053636f
C742 minus.t10 a_n1670_n3288# 0.363758f
C743 minus.t7 a_n1670_n3288# 0.363758f
C744 minus.t11 a_n1670_n3288# 0.363758f
C745 minus.n20 a_n1670_n3288# 0.149812f
C746 minus.n21 a_n1670_n3288# 0.053636f
C747 minus.t4 a_n1670_n3288# 0.363758f
C748 minus.t2 a_n1670_n3288# 0.363758f
C749 minus.t5 a_n1670_n3288# 0.363758f
C750 minus.n22 a_n1670_n3288# 0.149812f
C751 minus.t3 a_n1670_n3288# 0.36851f
C752 minus.n23 a_n1670_n3288# 0.165743f
C753 minus.n24 a_n1670_n3288# 0.120751f
C754 minus.n25 a_n1670_n3288# 0.018785f
C755 minus.n26 a_n1670_n3288# 0.149812f
C756 minus.n27 a_n1670_n3288# 0.018785f
C757 minus.n28 a_n1670_n3288# 0.149812f
C758 minus.n29 a_n1670_n3288# 0.018785f
C759 minus.n30 a_n1670_n3288# 0.053636f
C760 minus.n31 a_n1670_n3288# 0.053636f
C761 minus.n32 a_n1670_n3288# 0.018785f
C762 minus.n33 a_n1670_n3288# 0.149812f
C763 minus.n34 a_n1670_n3288# 0.018785f
C764 minus.n35 a_n1670_n3288# 0.149812f
C765 minus.t6 a_n1670_n3288# 0.36851f
C766 minus.n36 a_n1670_n3288# 0.165664f
C767 minus.n37 a_n1670_n3288# 0.346407f
C768 minus.n38 a_n1670_n3288# 2.22991f
.ends

