* NGSPICE file created from diffpair653.ext - technology: sky130A

.subckt diffpair653 minus drain_right drain_left source plus
X0 source.t13 plus.t0 drain_left.t0 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X1 drain_right.t7 minus.t0 source.t14 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X2 a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.2
X3 drain_left.t6 plus.t1 source.t12 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X4 a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X5 source.t3 minus.t1 drain_right.t6 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X6 source.t0 minus.t2 drain_right.t5 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X7 source.t15 minus.t3 drain_right.t4 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X8 drain_right.t3 minus.t4 source.t1 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X9 drain_right.t2 minus.t5 source.t2 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X10 source.t11 plus.t2 drain_left.t7 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X11 a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X12 drain_right.t1 minus.t6 source.t5 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X13 drain_left.t5 plus.t3 source.t10 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X14 source.t9 plus.t4 drain_left.t3 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X15 source.t4 minus.t7 drain_right.t0 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X16 a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X17 source.t8 plus.t5 drain_left.t2 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X18 drain_left.t1 plus.t6 source.t7 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X19 drain_left.t4 plus.t7 source.t6 a_n1246_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
R0 plus.n1 plus.t2 3212.24
R1 plus.n5 plus.t3 3212.24
R2 plus.n8 plus.t6 3212.24
R3 plus.n12 plus.t4 3212.24
R4 plus.n2 plus.t1 3169.15
R5 plus.n4 plus.t5 3169.15
R6 plus.n9 plus.t0 3169.15
R7 plus.n11 plus.t7 3169.15
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 38.7066
R15 plus.n4 plus.n3 38.7066
R16 plus.n11 plus.n10 38.7066
R17 plus.n10 plus.n9 38.7066
R18 plus.n2 plus.n1 34.3247
R19 plus.n5 plus.n4 34.3247
R20 plus.n12 plus.n11 34.3247
R21 plus.n9 plus.n8 34.3247
R22 plus plus.n13 32.5899
R23 plus plus.n6 17.0119
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 drain_left.n5 drain_left.n3 59.1723
R27 drain_left.n2 drain_left.n1 58.8885
R28 drain_left.n2 drain_left.n0 58.8885
R29 drain_left.n5 drain_left.n4 58.7153
R30 drain_left drain_left.n2 38.8147
R31 drain_left drain_left.n5 6.11011
R32 drain_left.n1 drain_left.t0 0.7925
R33 drain_left.n1 drain_left.t1 0.7925
R34 drain_left.n0 drain_left.t3 0.7925
R35 drain_left.n0 drain_left.t4 0.7925
R36 drain_left.n4 drain_left.t2 0.7925
R37 drain_left.n4 drain_left.t5 0.7925
R38 drain_left.n3 drain_left.t7 0.7925
R39 drain_left.n3 drain_left.t6 0.7925
R40 source.n1122 source.n988 289.615
R41 source.n980 source.n846 289.615
R42 source.n840 source.n706 289.615
R43 source.n698 source.n564 289.615
R44 source.n134 source.n0 289.615
R45 source.n276 source.n142 289.615
R46 source.n416 source.n282 289.615
R47 source.n558 source.n424 289.615
R48 source.n1032 source.n1031 185
R49 source.n1037 source.n1036 185
R50 source.n1039 source.n1038 185
R51 source.n1028 source.n1027 185
R52 source.n1045 source.n1044 185
R53 source.n1047 source.n1046 185
R54 source.n1024 source.n1023 185
R55 source.n1054 source.n1053 185
R56 source.n1055 source.n1022 185
R57 source.n1057 source.n1056 185
R58 source.n1020 source.n1019 185
R59 source.n1063 source.n1062 185
R60 source.n1065 source.n1064 185
R61 source.n1016 source.n1015 185
R62 source.n1071 source.n1070 185
R63 source.n1073 source.n1072 185
R64 source.n1012 source.n1011 185
R65 source.n1079 source.n1078 185
R66 source.n1081 source.n1080 185
R67 source.n1008 source.n1007 185
R68 source.n1087 source.n1086 185
R69 source.n1089 source.n1088 185
R70 source.n1004 source.n1003 185
R71 source.n1095 source.n1094 185
R72 source.n1098 source.n1097 185
R73 source.n1096 source.n1000 185
R74 source.n1103 source.n999 185
R75 source.n1105 source.n1104 185
R76 source.n1107 source.n1106 185
R77 source.n996 source.n995 185
R78 source.n1113 source.n1112 185
R79 source.n1115 source.n1114 185
R80 source.n992 source.n991 185
R81 source.n1121 source.n1120 185
R82 source.n1123 source.n1122 185
R83 source.n890 source.n889 185
R84 source.n895 source.n894 185
R85 source.n897 source.n896 185
R86 source.n886 source.n885 185
R87 source.n903 source.n902 185
R88 source.n905 source.n904 185
R89 source.n882 source.n881 185
R90 source.n912 source.n911 185
R91 source.n913 source.n880 185
R92 source.n915 source.n914 185
R93 source.n878 source.n877 185
R94 source.n921 source.n920 185
R95 source.n923 source.n922 185
R96 source.n874 source.n873 185
R97 source.n929 source.n928 185
R98 source.n931 source.n930 185
R99 source.n870 source.n869 185
R100 source.n937 source.n936 185
R101 source.n939 source.n938 185
R102 source.n866 source.n865 185
R103 source.n945 source.n944 185
R104 source.n947 source.n946 185
R105 source.n862 source.n861 185
R106 source.n953 source.n952 185
R107 source.n956 source.n955 185
R108 source.n954 source.n858 185
R109 source.n961 source.n857 185
R110 source.n963 source.n962 185
R111 source.n965 source.n964 185
R112 source.n854 source.n853 185
R113 source.n971 source.n970 185
R114 source.n973 source.n972 185
R115 source.n850 source.n849 185
R116 source.n979 source.n978 185
R117 source.n981 source.n980 185
R118 source.n750 source.n749 185
R119 source.n755 source.n754 185
R120 source.n757 source.n756 185
R121 source.n746 source.n745 185
R122 source.n763 source.n762 185
R123 source.n765 source.n764 185
R124 source.n742 source.n741 185
R125 source.n772 source.n771 185
R126 source.n773 source.n740 185
R127 source.n775 source.n774 185
R128 source.n738 source.n737 185
R129 source.n781 source.n780 185
R130 source.n783 source.n782 185
R131 source.n734 source.n733 185
R132 source.n789 source.n788 185
R133 source.n791 source.n790 185
R134 source.n730 source.n729 185
R135 source.n797 source.n796 185
R136 source.n799 source.n798 185
R137 source.n726 source.n725 185
R138 source.n805 source.n804 185
R139 source.n807 source.n806 185
R140 source.n722 source.n721 185
R141 source.n813 source.n812 185
R142 source.n816 source.n815 185
R143 source.n814 source.n718 185
R144 source.n821 source.n717 185
R145 source.n823 source.n822 185
R146 source.n825 source.n824 185
R147 source.n714 source.n713 185
R148 source.n831 source.n830 185
R149 source.n833 source.n832 185
R150 source.n710 source.n709 185
R151 source.n839 source.n838 185
R152 source.n841 source.n840 185
R153 source.n608 source.n607 185
R154 source.n613 source.n612 185
R155 source.n615 source.n614 185
R156 source.n604 source.n603 185
R157 source.n621 source.n620 185
R158 source.n623 source.n622 185
R159 source.n600 source.n599 185
R160 source.n630 source.n629 185
R161 source.n631 source.n598 185
R162 source.n633 source.n632 185
R163 source.n596 source.n595 185
R164 source.n639 source.n638 185
R165 source.n641 source.n640 185
R166 source.n592 source.n591 185
R167 source.n647 source.n646 185
R168 source.n649 source.n648 185
R169 source.n588 source.n587 185
R170 source.n655 source.n654 185
R171 source.n657 source.n656 185
R172 source.n584 source.n583 185
R173 source.n663 source.n662 185
R174 source.n665 source.n664 185
R175 source.n580 source.n579 185
R176 source.n671 source.n670 185
R177 source.n674 source.n673 185
R178 source.n672 source.n576 185
R179 source.n679 source.n575 185
R180 source.n681 source.n680 185
R181 source.n683 source.n682 185
R182 source.n572 source.n571 185
R183 source.n689 source.n688 185
R184 source.n691 source.n690 185
R185 source.n568 source.n567 185
R186 source.n697 source.n696 185
R187 source.n699 source.n698 185
R188 source.n135 source.n134 185
R189 source.n133 source.n132 185
R190 source.n4 source.n3 185
R191 source.n127 source.n126 185
R192 source.n125 source.n124 185
R193 source.n8 source.n7 185
R194 source.n119 source.n118 185
R195 source.n117 source.n116 185
R196 source.n115 source.n11 185
R197 source.n15 source.n12 185
R198 source.n110 source.n109 185
R199 source.n108 source.n107 185
R200 source.n17 source.n16 185
R201 source.n102 source.n101 185
R202 source.n100 source.n99 185
R203 source.n21 source.n20 185
R204 source.n94 source.n93 185
R205 source.n92 source.n91 185
R206 source.n25 source.n24 185
R207 source.n86 source.n85 185
R208 source.n84 source.n83 185
R209 source.n29 source.n28 185
R210 source.n78 source.n77 185
R211 source.n76 source.n75 185
R212 source.n33 source.n32 185
R213 source.n70 source.n69 185
R214 source.n68 source.n35 185
R215 source.n67 source.n66 185
R216 source.n38 source.n36 185
R217 source.n61 source.n60 185
R218 source.n59 source.n58 185
R219 source.n42 source.n41 185
R220 source.n53 source.n52 185
R221 source.n51 source.n50 185
R222 source.n46 source.n45 185
R223 source.n277 source.n276 185
R224 source.n275 source.n274 185
R225 source.n146 source.n145 185
R226 source.n269 source.n268 185
R227 source.n267 source.n266 185
R228 source.n150 source.n149 185
R229 source.n261 source.n260 185
R230 source.n259 source.n258 185
R231 source.n257 source.n153 185
R232 source.n157 source.n154 185
R233 source.n252 source.n251 185
R234 source.n250 source.n249 185
R235 source.n159 source.n158 185
R236 source.n244 source.n243 185
R237 source.n242 source.n241 185
R238 source.n163 source.n162 185
R239 source.n236 source.n235 185
R240 source.n234 source.n233 185
R241 source.n167 source.n166 185
R242 source.n228 source.n227 185
R243 source.n226 source.n225 185
R244 source.n171 source.n170 185
R245 source.n220 source.n219 185
R246 source.n218 source.n217 185
R247 source.n175 source.n174 185
R248 source.n212 source.n211 185
R249 source.n210 source.n177 185
R250 source.n209 source.n208 185
R251 source.n180 source.n178 185
R252 source.n203 source.n202 185
R253 source.n201 source.n200 185
R254 source.n184 source.n183 185
R255 source.n195 source.n194 185
R256 source.n193 source.n192 185
R257 source.n188 source.n187 185
R258 source.n417 source.n416 185
R259 source.n415 source.n414 185
R260 source.n286 source.n285 185
R261 source.n409 source.n408 185
R262 source.n407 source.n406 185
R263 source.n290 source.n289 185
R264 source.n401 source.n400 185
R265 source.n399 source.n398 185
R266 source.n397 source.n293 185
R267 source.n297 source.n294 185
R268 source.n392 source.n391 185
R269 source.n390 source.n389 185
R270 source.n299 source.n298 185
R271 source.n384 source.n383 185
R272 source.n382 source.n381 185
R273 source.n303 source.n302 185
R274 source.n376 source.n375 185
R275 source.n374 source.n373 185
R276 source.n307 source.n306 185
R277 source.n368 source.n367 185
R278 source.n366 source.n365 185
R279 source.n311 source.n310 185
R280 source.n360 source.n359 185
R281 source.n358 source.n357 185
R282 source.n315 source.n314 185
R283 source.n352 source.n351 185
R284 source.n350 source.n317 185
R285 source.n349 source.n348 185
R286 source.n320 source.n318 185
R287 source.n343 source.n342 185
R288 source.n341 source.n340 185
R289 source.n324 source.n323 185
R290 source.n335 source.n334 185
R291 source.n333 source.n332 185
R292 source.n328 source.n327 185
R293 source.n559 source.n558 185
R294 source.n557 source.n556 185
R295 source.n428 source.n427 185
R296 source.n551 source.n550 185
R297 source.n549 source.n548 185
R298 source.n432 source.n431 185
R299 source.n543 source.n542 185
R300 source.n541 source.n540 185
R301 source.n539 source.n435 185
R302 source.n439 source.n436 185
R303 source.n534 source.n533 185
R304 source.n532 source.n531 185
R305 source.n441 source.n440 185
R306 source.n526 source.n525 185
R307 source.n524 source.n523 185
R308 source.n445 source.n444 185
R309 source.n518 source.n517 185
R310 source.n516 source.n515 185
R311 source.n449 source.n448 185
R312 source.n510 source.n509 185
R313 source.n508 source.n507 185
R314 source.n453 source.n452 185
R315 source.n502 source.n501 185
R316 source.n500 source.n499 185
R317 source.n457 source.n456 185
R318 source.n494 source.n493 185
R319 source.n492 source.n459 185
R320 source.n491 source.n490 185
R321 source.n462 source.n460 185
R322 source.n485 source.n484 185
R323 source.n483 source.n482 185
R324 source.n466 source.n465 185
R325 source.n477 source.n476 185
R326 source.n475 source.n474 185
R327 source.n470 source.n469 185
R328 source.n1033 source.t1 149.524
R329 source.n891 source.t0 149.524
R330 source.n751 source.t7 149.524
R331 source.n609 source.t9 149.524
R332 source.n47 source.t10 149.524
R333 source.n189 source.t11 149.524
R334 source.n329 source.t5 149.524
R335 source.n471 source.t4 149.524
R336 source.n1037 source.n1031 104.615
R337 source.n1038 source.n1037 104.615
R338 source.n1038 source.n1027 104.615
R339 source.n1045 source.n1027 104.615
R340 source.n1046 source.n1045 104.615
R341 source.n1046 source.n1023 104.615
R342 source.n1054 source.n1023 104.615
R343 source.n1055 source.n1054 104.615
R344 source.n1056 source.n1055 104.615
R345 source.n1056 source.n1019 104.615
R346 source.n1063 source.n1019 104.615
R347 source.n1064 source.n1063 104.615
R348 source.n1064 source.n1015 104.615
R349 source.n1071 source.n1015 104.615
R350 source.n1072 source.n1071 104.615
R351 source.n1072 source.n1011 104.615
R352 source.n1079 source.n1011 104.615
R353 source.n1080 source.n1079 104.615
R354 source.n1080 source.n1007 104.615
R355 source.n1087 source.n1007 104.615
R356 source.n1088 source.n1087 104.615
R357 source.n1088 source.n1003 104.615
R358 source.n1095 source.n1003 104.615
R359 source.n1097 source.n1095 104.615
R360 source.n1097 source.n1096 104.615
R361 source.n1096 source.n999 104.615
R362 source.n1105 source.n999 104.615
R363 source.n1106 source.n1105 104.615
R364 source.n1106 source.n995 104.615
R365 source.n1113 source.n995 104.615
R366 source.n1114 source.n1113 104.615
R367 source.n1114 source.n991 104.615
R368 source.n1121 source.n991 104.615
R369 source.n1122 source.n1121 104.615
R370 source.n895 source.n889 104.615
R371 source.n896 source.n895 104.615
R372 source.n896 source.n885 104.615
R373 source.n903 source.n885 104.615
R374 source.n904 source.n903 104.615
R375 source.n904 source.n881 104.615
R376 source.n912 source.n881 104.615
R377 source.n913 source.n912 104.615
R378 source.n914 source.n913 104.615
R379 source.n914 source.n877 104.615
R380 source.n921 source.n877 104.615
R381 source.n922 source.n921 104.615
R382 source.n922 source.n873 104.615
R383 source.n929 source.n873 104.615
R384 source.n930 source.n929 104.615
R385 source.n930 source.n869 104.615
R386 source.n937 source.n869 104.615
R387 source.n938 source.n937 104.615
R388 source.n938 source.n865 104.615
R389 source.n945 source.n865 104.615
R390 source.n946 source.n945 104.615
R391 source.n946 source.n861 104.615
R392 source.n953 source.n861 104.615
R393 source.n955 source.n953 104.615
R394 source.n955 source.n954 104.615
R395 source.n954 source.n857 104.615
R396 source.n963 source.n857 104.615
R397 source.n964 source.n963 104.615
R398 source.n964 source.n853 104.615
R399 source.n971 source.n853 104.615
R400 source.n972 source.n971 104.615
R401 source.n972 source.n849 104.615
R402 source.n979 source.n849 104.615
R403 source.n980 source.n979 104.615
R404 source.n755 source.n749 104.615
R405 source.n756 source.n755 104.615
R406 source.n756 source.n745 104.615
R407 source.n763 source.n745 104.615
R408 source.n764 source.n763 104.615
R409 source.n764 source.n741 104.615
R410 source.n772 source.n741 104.615
R411 source.n773 source.n772 104.615
R412 source.n774 source.n773 104.615
R413 source.n774 source.n737 104.615
R414 source.n781 source.n737 104.615
R415 source.n782 source.n781 104.615
R416 source.n782 source.n733 104.615
R417 source.n789 source.n733 104.615
R418 source.n790 source.n789 104.615
R419 source.n790 source.n729 104.615
R420 source.n797 source.n729 104.615
R421 source.n798 source.n797 104.615
R422 source.n798 source.n725 104.615
R423 source.n805 source.n725 104.615
R424 source.n806 source.n805 104.615
R425 source.n806 source.n721 104.615
R426 source.n813 source.n721 104.615
R427 source.n815 source.n813 104.615
R428 source.n815 source.n814 104.615
R429 source.n814 source.n717 104.615
R430 source.n823 source.n717 104.615
R431 source.n824 source.n823 104.615
R432 source.n824 source.n713 104.615
R433 source.n831 source.n713 104.615
R434 source.n832 source.n831 104.615
R435 source.n832 source.n709 104.615
R436 source.n839 source.n709 104.615
R437 source.n840 source.n839 104.615
R438 source.n613 source.n607 104.615
R439 source.n614 source.n613 104.615
R440 source.n614 source.n603 104.615
R441 source.n621 source.n603 104.615
R442 source.n622 source.n621 104.615
R443 source.n622 source.n599 104.615
R444 source.n630 source.n599 104.615
R445 source.n631 source.n630 104.615
R446 source.n632 source.n631 104.615
R447 source.n632 source.n595 104.615
R448 source.n639 source.n595 104.615
R449 source.n640 source.n639 104.615
R450 source.n640 source.n591 104.615
R451 source.n647 source.n591 104.615
R452 source.n648 source.n647 104.615
R453 source.n648 source.n587 104.615
R454 source.n655 source.n587 104.615
R455 source.n656 source.n655 104.615
R456 source.n656 source.n583 104.615
R457 source.n663 source.n583 104.615
R458 source.n664 source.n663 104.615
R459 source.n664 source.n579 104.615
R460 source.n671 source.n579 104.615
R461 source.n673 source.n671 104.615
R462 source.n673 source.n672 104.615
R463 source.n672 source.n575 104.615
R464 source.n681 source.n575 104.615
R465 source.n682 source.n681 104.615
R466 source.n682 source.n571 104.615
R467 source.n689 source.n571 104.615
R468 source.n690 source.n689 104.615
R469 source.n690 source.n567 104.615
R470 source.n697 source.n567 104.615
R471 source.n698 source.n697 104.615
R472 source.n134 source.n133 104.615
R473 source.n133 source.n3 104.615
R474 source.n126 source.n3 104.615
R475 source.n126 source.n125 104.615
R476 source.n125 source.n7 104.615
R477 source.n118 source.n7 104.615
R478 source.n118 source.n117 104.615
R479 source.n117 source.n11 104.615
R480 source.n15 source.n11 104.615
R481 source.n109 source.n15 104.615
R482 source.n109 source.n108 104.615
R483 source.n108 source.n16 104.615
R484 source.n101 source.n16 104.615
R485 source.n101 source.n100 104.615
R486 source.n100 source.n20 104.615
R487 source.n93 source.n20 104.615
R488 source.n93 source.n92 104.615
R489 source.n92 source.n24 104.615
R490 source.n85 source.n24 104.615
R491 source.n85 source.n84 104.615
R492 source.n84 source.n28 104.615
R493 source.n77 source.n28 104.615
R494 source.n77 source.n76 104.615
R495 source.n76 source.n32 104.615
R496 source.n69 source.n32 104.615
R497 source.n69 source.n68 104.615
R498 source.n68 source.n67 104.615
R499 source.n67 source.n36 104.615
R500 source.n60 source.n36 104.615
R501 source.n60 source.n59 104.615
R502 source.n59 source.n41 104.615
R503 source.n52 source.n41 104.615
R504 source.n52 source.n51 104.615
R505 source.n51 source.n45 104.615
R506 source.n276 source.n275 104.615
R507 source.n275 source.n145 104.615
R508 source.n268 source.n145 104.615
R509 source.n268 source.n267 104.615
R510 source.n267 source.n149 104.615
R511 source.n260 source.n149 104.615
R512 source.n260 source.n259 104.615
R513 source.n259 source.n153 104.615
R514 source.n157 source.n153 104.615
R515 source.n251 source.n157 104.615
R516 source.n251 source.n250 104.615
R517 source.n250 source.n158 104.615
R518 source.n243 source.n158 104.615
R519 source.n243 source.n242 104.615
R520 source.n242 source.n162 104.615
R521 source.n235 source.n162 104.615
R522 source.n235 source.n234 104.615
R523 source.n234 source.n166 104.615
R524 source.n227 source.n166 104.615
R525 source.n227 source.n226 104.615
R526 source.n226 source.n170 104.615
R527 source.n219 source.n170 104.615
R528 source.n219 source.n218 104.615
R529 source.n218 source.n174 104.615
R530 source.n211 source.n174 104.615
R531 source.n211 source.n210 104.615
R532 source.n210 source.n209 104.615
R533 source.n209 source.n178 104.615
R534 source.n202 source.n178 104.615
R535 source.n202 source.n201 104.615
R536 source.n201 source.n183 104.615
R537 source.n194 source.n183 104.615
R538 source.n194 source.n193 104.615
R539 source.n193 source.n187 104.615
R540 source.n416 source.n415 104.615
R541 source.n415 source.n285 104.615
R542 source.n408 source.n285 104.615
R543 source.n408 source.n407 104.615
R544 source.n407 source.n289 104.615
R545 source.n400 source.n289 104.615
R546 source.n400 source.n399 104.615
R547 source.n399 source.n293 104.615
R548 source.n297 source.n293 104.615
R549 source.n391 source.n297 104.615
R550 source.n391 source.n390 104.615
R551 source.n390 source.n298 104.615
R552 source.n383 source.n298 104.615
R553 source.n383 source.n382 104.615
R554 source.n382 source.n302 104.615
R555 source.n375 source.n302 104.615
R556 source.n375 source.n374 104.615
R557 source.n374 source.n306 104.615
R558 source.n367 source.n306 104.615
R559 source.n367 source.n366 104.615
R560 source.n366 source.n310 104.615
R561 source.n359 source.n310 104.615
R562 source.n359 source.n358 104.615
R563 source.n358 source.n314 104.615
R564 source.n351 source.n314 104.615
R565 source.n351 source.n350 104.615
R566 source.n350 source.n349 104.615
R567 source.n349 source.n318 104.615
R568 source.n342 source.n318 104.615
R569 source.n342 source.n341 104.615
R570 source.n341 source.n323 104.615
R571 source.n334 source.n323 104.615
R572 source.n334 source.n333 104.615
R573 source.n333 source.n327 104.615
R574 source.n558 source.n557 104.615
R575 source.n557 source.n427 104.615
R576 source.n550 source.n427 104.615
R577 source.n550 source.n549 104.615
R578 source.n549 source.n431 104.615
R579 source.n542 source.n431 104.615
R580 source.n542 source.n541 104.615
R581 source.n541 source.n435 104.615
R582 source.n439 source.n435 104.615
R583 source.n533 source.n439 104.615
R584 source.n533 source.n532 104.615
R585 source.n532 source.n440 104.615
R586 source.n525 source.n440 104.615
R587 source.n525 source.n524 104.615
R588 source.n524 source.n444 104.615
R589 source.n517 source.n444 104.615
R590 source.n517 source.n516 104.615
R591 source.n516 source.n448 104.615
R592 source.n509 source.n448 104.615
R593 source.n509 source.n508 104.615
R594 source.n508 source.n452 104.615
R595 source.n501 source.n452 104.615
R596 source.n501 source.n500 104.615
R597 source.n500 source.n456 104.615
R598 source.n493 source.n456 104.615
R599 source.n493 source.n492 104.615
R600 source.n492 source.n491 104.615
R601 source.n491 source.n460 104.615
R602 source.n484 source.n460 104.615
R603 source.n484 source.n483 104.615
R604 source.n483 source.n465 104.615
R605 source.n476 source.n465 104.615
R606 source.n476 source.n475 104.615
R607 source.n475 source.n469 104.615
R608 source.t1 source.n1031 52.3082
R609 source.t0 source.n889 52.3082
R610 source.t7 source.n749 52.3082
R611 source.t9 source.n607 52.3082
R612 source.t10 source.n45 52.3082
R613 source.t11 source.n187 52.3082
R614 source.t5 source.n327 52.3082
R615 source.t4 source.n469 52.3082
R616 source.n987 source.n986 42.0366
R617 source.n705 source.n704 42.0366
R618 source.n141 source.n140 42.0366
R619 source.n423 source.n422 42.0366
R620 source.n703 source.n563 31.5931
R621 source.n1127 source.n1126 30.6338
R622 source.n985 source.n984 30.6338
R623 source.n845 source.n844 30.6338
R624 source.n703 source.n702 30.6338
R625 source.n139 source.n138 30.6338
R626 source.n281 source.n280 30.6338
R627 source.n421 source.n420 30.6338
R628 source.n563 source.n562 30.6338
R629 source.n1128 source.n139 26.1017
R630 source.n1057 source.n1022 13.1884
R631 source.n1104 source.n1103 13.1884
R632 source.n915 source.n880 13.1884
R633 source.n962 source.n961 13.1884
R634 source.n775 source.n740 13.1884
R635 source.n822 source.n821 13.1884
R636 source.n633 source.n598 13.1884
R637 source.n680 source.n679 13.1884
R638 source.n116 source.n115 13.1884
R639 source.n70 source.n35 13.1884
R640 source.n258 source.n257 13.1884
R641 source.n212 source.n177 13.1884
R642 source.n398 source.n397 13.1884
R643 source.n352 source.n317 13.1884
R644 source.n540 source.n539 13.1884
R645 source.n494 source.n459 13.1884
R646 source.n1053 source.n1052 12.8005
R647 source.n1058 source.n1020 12.8005
R648 source.n1102 source.n1000 12.8005
R649 source.n1107 source.n998 12.8005
R650 source.n911 source.n910 12.8005
R651 source.n916 source.n878 12.8005
R652 source.n960 source.n858 12.8005
R653 source.n965 source.n856 12.8005
R654 source.n771 source.n770 12.8005
R655 source.n776 source.n738 12.8005
R656 source.n820 source.n718 12.8005
R657 source.n825 source.n716 12.8005
R658 source.n629 source.n628 12.8005
R659 source.n634 source.n596 12.8005
R660 source.n678 source.n576 12.8005
R661 source.n683 source.n574 12.8005
R662 source.n119 source.n10 12.8005
R663 source.n114 source.n12 12.8005
R664 source.n71 source.n33 12.8005
R665 source.n66 source.n37 12.8005
R666 source.n261 source.n152 12.8005
R667 source.n256 source.n154 12.8005
R668 source.n213 source.n175 12.8005
R669 source.n208 source.n179 12.8005
R670 source.n401 source.n292 12.8005
R671 source.n396 source.n294 12.8005
R672 source.n353 source.n315 12.8005
R673 source.n348 source.n319 12.8005
R674 source.n543 source.n434 12.8005
R675 source.n538 source.n436 12.8005
R676 source.n495 source.n457 12.8005
R677 source.n490 source.n461 12.8005
R678 source.n1051 source.n1024 12.0247
R679 source.n1062 source.n1061 12.0247
R680 source.n1099 source.n1098 12.0247
R681 source.n1108 source.n996 12.0247
R682 source.n909 source.n882 12.0247
R683 source.n920 source.n919 12.0247
R684 source.n957 source.n956 12.0247
R685 source.n966 source.n854 12.0247
R686 source.n769 source.n742 12.0247
R687 source.n780 source.n779 12.0247
R688 source.n817 source.n816 12.0247
R689 source.n826 source.n714 12.0247
R690 source.n627 source.n600 12.0247
R691 source.n638 source.n637 12.0247
R692 source.n675 source.n674 12.0247
R693 source.n684 source.n572 12.0247
R694 source.n120 source.n8 12.0247
R695 source.n111 source.n110 12.0247
R696 source.n75 source.n74 12.0247
R697 source.n65 source.n38 12.0247
R698 source.n262 source.n150 12.0247
R699 source.n253 source.n252 12.0247
R700 source.n217 source.n216 12.0247
R701 source.n207 source.n180 12.0247
R702 source.n402 source.n290 12.0247
R703 source.n393 source.n392 12.0247
R704 source.n357 source.n356 12.0247
R705 source.n347 source.n320 12.0247
R706 source.n544 source.n432 12.0247
R707 source.n535 source.n534 12.0247
R708 source.n499 source.n498 12.0247
R709 source.n489 source.n462 12.0247
R710 source.n1048 source.n1047 11.249
R711 source.n1065 source.n1018 11.249
R712 source.n1094 source.n1002 11.249
R713 source.n1112 source.n1111 11.249
R714 source.n906 source.n905 11.249
R715 source.n923 source.n876 11.249
R716 source.n952 source.n860 11.249
R717 source.n970 source.n969 11.249
R718 source.n766 source.n765 11.249
R719 source.n783 source.n736 11.249
R720 source.n812 source.n720 11.249
R721 source.n830 source.n829 11.249
R722 source.n624 source.n623 11.249
R723 source.n641 source.n594 11.249
R724 source.n670 source.n578 11.249
R725 source.n688 source.n687 11.249
R726 source.n124 source.n123 11.249
R727 source.n107 source.n14 11.249
R728 source.n78 source.n31 11.249
R729 source.n62 source.n61 11.249
R730 source.n266 source.n265 11.249
R731 source.n249 source.n156 11.249
R732 source.n220 source.n173 11.249
R733 source.n204 source.n203 11.249
R734 source.n406 source.n405 11.249
R735 source.n389 source.n296 11.249
R736 source.n360 source.n313 11.249
R737 source.n344 source.n343 11.249
R738 source.n548 source.n547 11.249
R739 source.n531 source.n438 11.249
R740 source.n502 source.n455 11.249
R741 source.n486 source.n485 11.249
R742 source.n1044 source.n1026 10.4732
R743 source.n1066 source.n1016 10.4732
R744 source.n1093 source.n1004 10.4732
R745 source.n1115 source.n994 10.4732
R746 source.n902 source.n884 10.4732
R747 source.n924 source.n874 10.4732
R748 source.n951 source.n862 10.4732
R749 source.n973 source.n852 10.4732
R750 source.n762 source.n744 10.4732
R751 source.n784 source.n734 10.4732
R752 source.n811 source.n722 10.4732
R753 source.n833 source.n712 10.4732
R754 source.n620 source.n602 10.4732
R755 source.n642 source.n592 10.4732
R756 source.n669 source.n580 10.4732
R757 source.n691 source.n570 10.4732
R758 source.n127 source.n6 10.4732
R759 source.n106 source.n17 10.4732
R760 source.n79 source.n29 10.4732
R761 source.n58 source.n40 10.4732
R762 source.n269 source.n148 10.4732
R763 source.n248 source.n159 10.4732
R764 source.n221 source.n171 10.4732
R765 source.n200 source.n182 10.4732
R766 source.n409 source.n288 10.4732
R767 source.n388 source.n299 10.4732
R768 source.n361 source.n311 10.4732
R769 source.n340 source.n322 10.4732
R770 source.n551 source.n430 10.4732
R771 source.n530 source.n441 10.4732
R772 source.n503 source.n453 10.4732
R773 source.n482 source.n464 10.4732
R774 source.n1033 source.n1032 10.2747
R775 source.n891 source.n890 10.2747
R776 source.n751 source.n750 10.2747
R777 source.n609 source.n608 10.2747
R778 source.n47 source.n46 10.2747
R779 source.n189 source.n188 10.2747
R780 source.n329 source.n328 10.2747
R781 source.n471 source.n470 10.2747
R782 source.n1043 source.n1028 9.69747
R783 source.n1070 source.n1069 9.69747
R784 source.n1090 source.n1089 9.69747
R785 source.n1116 source.n992 9.69747
R786 source.n901 source.n886 9.69747
R787 source.n928 source.n927 9.69747
R788 source.n948 source.n947 9.69747
R789 source.n974 source.n850 9.69747
R790 source.n761 source.n746 9.69747
R791 source.n788 source.n787 9.69747
R792 source.n808 source.n807 9.69747
R793 source.n834 source.n710 9.69747
R794 source.n619 source.n604 9.69747
R795 source.n646 source.n645 9.69747
R796 source.n666 source.n665 9.69747
R797 source.n692 source.n568 9.69747
R798 source.n128 source.n4 9.69747
R799 source.n103 source.n102 9.69747
R800 source.n83 source.n82 9.69747
R801 source.n57 source.n42 9.69747
R802 source.n270 source.n146 9.69747
R803 source.n245 source.n244 9.69747
R804 source.n225 source.n224 9.69747
R805 source.n199 source.n184 9.69747
R806 source.n410 source.n286 9.69747
R807 source.n385 source.n384 9.69747
R808 source.n365 source.n364 9.69747
R809 source.n339 source.n324 9.69747
R810 source.n552 source.n428 9.69747
R811 source.n527 source.n526 9.69747
R812 source.n507 source.n506 9.69747
R813 source.n481 source.n466 9.69747
R814 source.n1126 source.n1125 9.45567
R815 source.n984 source.n983 9.45567
R816 source.n844 source.n843 9.45567
R817 source.n702 source.n701 9.45567
R818 source.n138 source.n137 9.45567
R819 source.n280 source.n279 9.45567
R820 source.n420 source.n419 9.45567
R821 source.n562 source.n561 9.45567
R822 source.n990 source.n989 9.3005
R823 source.n1119 source.n1118 9.3005
R824 source.n1117 source.n1116 9.3005
R825 source.n994 source.n993 9.3005
R826 source.n1111 source.n1110 9.3005
R827 source.n1109 source.n1108 9.3005
R828 source.n998 source.n997 9.3005
R829 source.n1077 source.n1076 9.3005
R830 source.n1075 source.n1074 9.3005
R831 source.n1014 source.n1013 9.3005
R832 source.n1069 source.n1068 9.3005
R833 source.n1067 source.n1066 9.3005
R834 source.n1018 source.n1017 9.3005
R835 source.n1061 source.n1060 9.3005
R836 source.n1059 source.n1058 9.3005
R837 source.n1035 source.n1034 9.3005
R838 source.n1030 source.n1029 9.3005
R839 source.n1041 source.n1040 9.3005
R840 source.n1043 source.n1042 9.3005
R841 source.n1026 source.n1025 9.3005
R842 source.n1049 source.n1048 9.3005
R843 source.n1051 source.n1050 9.3005
R844 source.n1052 source.n1021 9.3005
R845 source.n1010 source.n1009 9.3005
R846 source.n1083 source.n1082 9.3005
R847 source.n1085 source.n1084 9.3005
R848 source.n1006 source.n1005 9.3005
R849 source.n1091 source.n1090 9.3005
R850 source.n1093 source.n1092 9.3005
R851 source.n1002 source.n1001 9.3005
R852 source.n1100 source.n1099 9.3005
R853 source.n1102 source.n1101 9.3005
R854 source.n1125 source.n1124 9.3005
R855 source.n848 source.n847 9.3005
R856 source.n977 source.n976 9.3005
R857 source.n975 source.n974 9.3005
R858 source.n852 source.n851 9.3005
R859 source.n969 source.n968 9.3005
R860 source.n967 source.n966 9.3005
R861 source.n856 source.n855 9.3005
R862 source.n935 source.n934 9.3005
R863 source.n933 source.n932 9.3005
R864 source.n872 source.n871 9.3005
R865 source.n927 source.n926 9.3005
R866 source.n925 source.n924 9.3005
R867 source.n876 source.n875 9.3005
R868 source.n919 source.n918 9.3005
R869 source.n917 source.n916 9.3005
R870 source.n893 source.n892 9.3005
R871 source.n888 source.n887 9.3005
R872 source.n899 source.n898 9.3005
R873 source.n901 source.n900 9.3005
R874 source.n884 source.n883 9.3005
R875 source.n907 source.n906 9.3005
R876 source.n909 source.n908 9.3005
R877 source.n910 source.n879 9.3005
R878 source.n868 source.n867 9.3005
R879 source.n941 source.n940 9.3005
R880 source.n943 source.n942 9.3005
R881 source.n864 source.n863 9.3005
R882 source.n949 source.n948 9.3005
R883 source.n951 source.n950 9.3005
R884 source.n860 source.n859 9.3005
R885 source.n958 source.n957 9.3005
R886 source.n960 source.n959 9.3005
R887 source.n983 source.n982 9.3005
R888 source.n708 source.n707 9.3005
R889 source.n837 source.n836 9.3005
R890 source.n835 source.n834 9.3005
R891 source.n712 source.n711 9.3005
R892 source.n829 source.n828 9.3005
R893 source.n827 source.n826 9.3005
R894 source.n716 source.n715 9.3005
R895 source.n795 source.n794 9.3005
R896 source.n793 source.n792 9.3005
R897 source.n732 source.n731 9.3005
R898 source.n787 source.n786 9.3005
R899 source.n785 source.n784 9.3005
R900 source.n736 source.n735 9.3005
R901 source.n779 source.n778 9.3005
R902 source.n777 source.n776 9.3005
R903 source.n753 source.n752 9.3005
R904 source.n748 source.n747 9.3005
R905 source.n759 source.n758 9.3005
R906 source.n761 source.n760 9.3005
R907 source.n744 source.n743 9.3005
R908 source.n767 source.n766 9.3005
R909 source.n769 source.n768 9.3005
R910 source.n770 source.n739 9.3005
R911 source.n728 source.n727 9.3005
R912 source.n801 source.n800 9.3005
R913 source.n803 source.n802 9.3005
R914 source.n724 source.n723 9.3005
R915 source.n809 source.n808 9.3005
R916 source.n811 source.n810 9.3005
R917 source.n720 source.n719 9.3005
R918 source.n818 source.n817 9.3005
R919 source.n820 source.n819 9.3005
R920 source.n843 source.n842 9.3005
R921 source.n566 source.n565 9.3005
R922 source.n695 source.n694 9.3005
R923 source.n693 source.n692 9.3005
R924 source.n570 source.n569 9.3005
R925 source.n687 source.n686 9.3005
R926 source.n685 source.n684 9.3005
R927 source.n574 source.n573 9.3005
R928 source.n653 source.n652 9.3005
R929 source.n651 source.n650 9.3005
R930 source.n590 source.n589 9.3005
R931 source.n645 source.n644 9.3005
R932 source.n643 source.n642 9.3005
R933 source.n594 source.n593 9.3005
R934 source.n637 source.n636 9.3005
R935 source.n635 source.n634 9.3005
R936 source.n611 source.n610 9.3005
R937 source.n606 source.n605 9.3005
R938 source.n617 source.n616 9.3005
R939 source.n619 source.n618 9.3005
R940 source.n602 source.n601 9.3005
R941 source.n625 source.n624 9.3005
R942 source.n627 source.n626 9.3005
R943 source.n628 source.n597 9.3005
R944 source.n586 source.n585 9.3005
R945 source.n659 source.n658 9.3005
R946 source.n661 source.n660 9.3005
R947 source.n582 source.n581 9.3005
R948 source.n667 source.n666 9.3005
R949 source.n669 source.n668 9.3005
R950 source.n578 source.n577 9.3005
R951 source.n676 source.n675 9.3005
R952 source.n678 source.n677 9.3005
R953 source.n701 source.n700 9.3005
R954 source.n49 source.n48 9.3005
R955 source.n44 source.n43 9.3005
R956 source.n55 source.n54 9.3005
R957 source.n57 source.n56 9.3005
R958 source.n40 source.n39 9.3005
R959 source.n63 source.n62 9.3005
R960 source.n65 source.n64 9.3005
R961 source.n37 source.n34 9.3005
R962 source.n96 source.n95 9.3005
R963 source.n98 source.n97 9.3005
R964 source.n19 source.n18 9.3005
R965 source.n104 source.n103 9.3005
R966 source.n106 source.n105 9.3005
R967 source.n14 source.n13 9.3005
R968 source.n112 source.n111 9.3005
R969 source.n114 source.n113 9.3005
R970 source.n137 source.n136 9.3005
R971 source.n2 source.n1 9.3005
R972 source.n131 source.n130 9.3005
R973 source.n129 source.n128 9.3005
R974 source.n6 source.n5 9.3005
R975 source.n123 source.n122 9.3005
R976 source.n121 source.n120 9.3005
R977 source.n10 source.n9 9.3005
R978 source.n23 source.n22 9.3005
R979 source.n90 source.n89 9.3005
R980 source.n88 source.n87 9.3005
R981 source.n27 source.n26 9.3005
R982 source.n82 source.n81 9.3005
R983 source.n80 source.n79 9.3005
R984 source.n31 source.n30 9.3005
R985 source.n74 source.n73 9.3005
R986 source.n72 source.n71 9.3005
R987 source.n191 source.n190 9.3005
R988 source.n186 source.n185 9.3005
R989 source.n197 source.n196 9.3005
R990 source.n199 source.n198 9.3005
R991 source.n182 source.n181 9.3005
R992 source.n205 source.n204 9.3005
R993 source.n207 source.n206 9.3005
R994 source.n179 source.n176 9.3005
R995 source.n238 source.n237 9.3005
R996 source.n240 source.n239 9.3005
R997 source.n161 source.n160 9.3005
R998 source.n246 source.n245 9.3005
R999 source.n248 source.n247 9.3005
R1000 source.n156 source.n155 9.3005
R1001 source.n254 source.n253 9.3005
R1002 source.n256 source.n255 9.3005
R1003 source.n279 source.n278 9.3005
R1004 source.n144 source.n143 9.3005
R1005 source.n273 source.n272 9.3005
R1006 source.n271 source.n270 9.3005
R1007 source.n148 source.n147 9.3005
R1008 source.n265 source.n264 9.3005
R1009 source.n263 source.n262 9.3005
R1010 source.n152 source.n151 9.3005
R1011 source.n165 source.n164 9.3005
R1012 source.n232 source.n231 9.3005
R1013 source.n230 source.n229 9.3005
R1014 source.n169 source.n168 9.3005
R1015 source.n224 source.n223 9.3005
R1016 source.n222 source.n221 9.3005
R1017 source.n173 source.n172 9.3005
R1018 source.n216 source.n215 9.3005
R1019 source.n214 source.n213 9.3005
R1020 source.n331 source.n330 9.3005
R1021 source.n326 source.n325 9.3005
R1022 source.n337 source.n336 9.3005
R1023 source.n339 source.n338 9.3005
R1024 source.n322 source.n321 9.3005
R1025 source.n345 source.n344 9.3005
R1026 source.n347 source.n346 9.3005
R1027 source.n319 source.n316 9.3005
R1028 source.n378 source.n377 9.3005
R1029 source.n380 source.n379 9.3005
R1030 source.n301 source.n300 9.3005
R1031 source.n386 source.n385 9.3005
R1032 source.n388 source.n387 9.3005
R1033 source.n296 source.n295 9.3005
R1034 source.n394 source.n393 9.3005
R1035 source.n396 source.n395 9.3005
R1036 source.n419 source.n418 9.3005
R1037 source.n284 source.n283 9.3005
R1038 source.n413 source.n412 9.3005
R1039 source.n411 source.n410 9.3005
R1040 source.n288 source.n287 9.3005
R1041 source.n405 source.n404 9.3005
R1042 source.n403 source.n402 9.3005
R1043 source.n292 source.n291 9.3005
R1044 source.n305 source.n304 9.3005
R1045 source.n372 source.n371 9.3005
R1046 source.n370 source.n369 9.3005
R1047 source.n309 source.n308 9.3005
R1048 source.n364 source.n363 9.3005
R1049 source.n362 source.n361 9.3005
R1050 source.n313 source.n312 9.3005
R1051 source.n356 source.n355 9.3005
R1052 source.n354 source.n353 9.3005
R1053 source.n473 source.n472 9.3005
R1054 source.n468 source.n467 9.3005
R1055 source.n479 source.n478 9.3005
R1056 source.n481 source.n480 9.3005
R1057 source.n464 source.n463 9.3005
R1058 source.n487 source.n486 9.3005
R1059 source.n489 source.n488 9.3005
R1060 source.n461 source.n458 9.3005
R1061 source.n520 source.n519 9.3005
R1062 source.n522 source.n521 9.3005
R1063 source.n443 source.n442 9.3005
R1064 source.n528 source.n527 9.3005
R1065 source.n530 source.n529 9.3005
R1066 source.n438 source.n437 9.3005
R1067 source.n536 source.n535 9.3005
R1068 source.n538 source.n537 9.3005
R1069 source.n561 source.n560 9.3005
R1070 source.n426 source.n425 9.3005
R1071 source.n555 source.n554 9.3005
R1072 source.n553 source.n552 9.3005
R1073 source.n430 source.n429 9.3005
R1074 source.n547 source.n546 9.3005
R1075 source.n545 source.n544 9.3005
R1076 source.n434 source.n433 9.3005
R1077 source.n447 source.n446 9.3005
R1078 source.n514 source.n513 9.3005
R1079 source.n512 source.n511 9.3005
R1080 source.n451 source.n450 9.3005
R1081 source.n506 source.n505 9.3005
R1082 source.n504 source.n503 9.3005
R1083 source.n455 source.n454 9.3005
R1084 source.n498 source.n497 9.3005
R1085 source.n496 source.n495 9.3005
R1086 source.n1040 source.n1039 8.92171
R1087 source.n1073 source.n1014 8.92171
R1088 source.n1086 source.n1006 8.92171
R1089 source.n1120 source.n1119 8.92171
R1090 source.n898 source.n897 8.92171
R1091 source.n931 source.n872 8.92171
R1092 source.n944 source.n864 8.92171
R1093 source.n978 source.n977 8.92171
R1094 source.n758 source.n757 8.92171
R1095 source.n791 source.n732 8.92171
R1096 source.n804 source.n724 8.92171
R1097 source.n838 source.n837 8.92171
R1098 source.n616 source.n615 8.92171
R1099 source.n649 source.n590 8.92171
R1100 source.n662 source.n582 8.92171
R1101 source.n696 source.n695 8.92171
R1102 source.n132 source.n131 8.92171
R1103 source.n99 source.n19 8.92171
R1104 source.n86 source.n27 8.92171
R1105 source.n54 source.n53 8.92171
R1106 source.n274 source.n273 8.92171
R1107 source.n241 source.n161 8.92171
R1108 source.n228 source.n169 8.92171
R1109 source.n196 source.n195 8.92171
R1110 source.n414 source.n413 8.92171
R1111 source.n381 source.n301 8.92171
R1112 source.n368 source.n309 8.92171
R1113 source.n336 source.n335 8.92171
R1114 source.n556 source.n555 8.92171
R1115 source.n523 source.n443 8.92171
R1116 source.n510 source.n451 8.92171
R1117 source.n478 source.n477 8.92171
R1118 source.n1036 source.n1030 8.14595
R1119 source.n1074 source.n1012 8.14595
R1120 source.n1085 source.n1008 8.14595
R1121 source.n1123 source.n990 8.14595
R1122 source.n894 source.n888 8.14595
R1123 source.n932 source.n870 8.14595
R1124 source.n943 source.n866 8.14595
R1125 source.n981 source.n848 8.14595
R1126 source.n754 source.n748 8.14595
R1127 source.n792 source.n730 8.14595
R1128 source.n803 source.n726 8.14595
R1129 source.n841 source.n708 8.14595
R1130 source.n612 source.n606 8.14595
R1131 source.n650 source.n588 8.14595
R1132 source.n661 source.n584 8.14595
R1133 source.n699 source.n566 8.14595
R1134 source.n135 source.n2 8.14595
R1135 source.n98 source.n21 8.14595
R1136 source.n87 source.n25 8.14595
R1137 source.n50 source.n44 8.14595
R1138 source.n277 source.n144 8.14595
R1139 source.n240 source.n163 8.14595
R1140 source.n229 source.n167 8.14595
R1141 source.n192 source.n186 8.14595
R1142 source.n417 source.n284 8.14595
R1143 source.n380 source.n303 8.14595
R1144 source.n369 source.n307 8.14595
R1145 source.n332 source.n326 8.14595
R1146 source.n559 source.n426 8.14595
R1147 source.n522 source.n445 8.14595
R1148 source.n511 source.n449 8.14595
R1149 source.n474 source.n468 8.14595
R1150 source.n1035 source.n1032 7.3702
R1151 source.n1078 source.n1077 7.3702
R1152 source.n1082 source.n1081 7.3702
R1153 source.n1124 source.n988 7.3702
R1154 source.n893 source.n890 7.3702
R1155 source.n936 source.n935 7.3702
R1156 source.n940 source.n939 7.3702
R1157 source.n982 source.n846 7.3702
R1158 source.n753 source.n750 7.3702
R1159 source.n796 source.n795 7.3702
R1160 source.n800 source.n799 7.3702
R1161 source.n842 source.n706 7.3702
R1162 source.n611 source.n608 7.3702
R1163 source.n654 source.n653 7.3702
R1164 source.n658 source.n657 7.3702
R1165 source.n700 source.n564 7.3702
R1166 source.n136 source.n0 7.3702
R1167 source.n95 source.n94 7.3702
R1168 source.n91 source.n90 7.3702
R1169 source.n49 source.n46 7.3702
R1170 source.n278 source.n142 7.3702
R1171 source.n237 source.n236 7.3702
R1172 source.n233 source.n232 7.3702
R1173 source.n191 source.n188 7.3702
R1174 source.n418 source.n282 7.3702
R1175 source.n377 source.n376 7.3702
R1176 source.n373 source.n372 7.3702
R1177 source.n331 source.n328 7.3702
R1178 source.n560 source.n424 7.3702
R1179 source.n519 source.n518 7.3702
R1180 source.n515 source.n514 7.3702
R1181 source.n473 source.n470 7.3702
R1182 source.n1078 source.n1010 6.59444
R1183 source.n1081 source.n1010 6.59444
R1184 source.n1126 source.n988 6.59444
R1185 source.n936 source.n868 6.59444
R1186 source.n939 source.n868 6.59444
R1187 source.n984 source.n846 6.59444
R1188 source.n796 source.n728 6.59444
R1189 source.n799 source.n728 6.59444
R1190 source.n844 source.n706 6.59444
R1191 source.n654 source.n586 6.59444
R1192 source.n657 source.n586 6.59444
R1193 source.n702 source.n564 6.59444
R1194 source.n138 source.n0 6.59444
R1195 source.n94 source.n23 6.59444
R1196 source.n91 source.n23 6.59444
R1197 source.n280 source.n142 6.59444
R1198 source.n236 source.n165 6.59444
R1199 source.n233 source.n165 6.59444
R1200 source.n420 source.n282 6.59444
R1201 source.n376 source.n305 6.59444
R1202 source.n373 source.n305 6.59444
R1203 source.n562 source.n424 6.59444
R1204 source.n518 source.n447 6.59444
R1205 source.n515 source.n447 6.59444
R1206 source.n1036 source.n1035 5.81868
R1207 source.n1077 source.n1012 5.81868
R1208 source.n1082 source.n1008 5.81868
R1209 source.n1124 source.n1123 5.81868
R1210 source.n894 source.n893 5.81868
R1211 source.n935 source.n870 5.81868
R1212 source.n940 source.n866 5.81868
R1213 source.n982 source.n981 5.81868
R1214 source.n754 source.n753 5.81868
R1215 source.n795 source.n730 5.81868
R1216 source.n800 source.n726 5.81868
R1217 source.n842 source.n841 5.81868
R1218 source.n612 source.n611 5.81868
R1219 source.n653 source.n588 5.81868
R1220 source.n658 source.n584 5.81868
R1221 source.n700 source.n699 5.81868
R1222 source.n136 source.n135 5.81868
R1223 source.n95 source.n21 5.81868
R1224 source.n90 source.n25 5.81868
R1225 source.n50 source.n49 5.81868
R1226 source.n278 source.n277 5.81868
R1227 source.n237 source.n163 5.81868
R1228 source.n232 source.n167 5.81868
R1229 source.n192 source.n191 5.81868
R1230 source.n418 source.n417 5.81868
R1231 source.n377 source.n303 5.81868
R1232 source.n372 source.n307 5.81868
R1233 source.n332 source.n331 5.81868
R1234 source.n560 source.n559 5.81868
R1235 source.n519 source.n445 5.81868
R1236 source.n514 source.n449 5.81868
R1237 source.n474 source.n473 5.81868
R1238 source.n1128 source.n1127 5.49188
R1239 source.n1039 source.n1030 5.04292
R1240 source.n1074 source.n1073 5.04292
R1241 source.n1086 source.n1085 5.04292
R1242 source.n1120 source.n990 5.04292
R1243 source.n897 source.n888 5.04292
R1244 source.n932 source.n931 5.04292
R1245 source.n944 source.n943 5.04292
R1246 source.n978 source.n848 5.04292
R1247 source.n757 source.n748 5.04292
R1248 source.n792 source.n791 5.04292
R1249 source.n804 source.n803 5.04292
R1250 source.n838 source.n708 5.04292
R1251 source.n615 source.n606 5.04292
R1252 source.n650 source.n649 5.04292
R1253 source.n662 source.n661 5.04292
R1254 source.n696 source.n566 5.04292
R1255 source.n132 source.n2 5.04292
R1256 source.n99 source.n98 5.04292
R1257 source.n87 source.n86 5.04292
R1258 source.n53 source.n44 5.04292
R1259 source.n274 source.n144 5.04292
R1260 source.n241 source.n240 5.04292
R1261 source.n229 source.n228 5.04292
R1262 source.n195 source.n186 5.04292
R1263 source.n414 source.n284 5.04292
R1264 source.n381 source.n380 5.04292
R1265 source.n369 source.n368 5.04292
R1266 source.n335 source.n326 5.04292
R1267 source.n556 source.n426 5.04292
R1268 source.n523 source.n522 5.04292
R1269 source.n511 source.n510 5.04292
R1270 source.n477 source.n468 5.04292
R1271 source.n1040 source.n1028 4.26717
R1272 source.n1070 source.n1014 4.26717
R1273 source.n1089 source.n1006 4.26717
R1274 source.n1119 source.n992 4.26717
R1275 source.n898 source.n886 4.26717
R1276 source.n928 source.n872 4.26717
R1277 source.n947 source.n864 4.26717
R1278 source.n977 source.n850 4.26717
R1279 source.n758 source.n746 4.26717
R1280 source.n788 source.n732 4.26717
R1281 source.n807 source.n724 4.26717
R1282 source.n837 source.n710 4.26717
R1283 source.n616 source.n604 4.26717
R1284 source.n646 source.n590 4.26717
R1285 source.n665 source.n582 4.26717
R1286 source.n695 source.n568 4.26717
R1287 source.n131 source.n4 4.26717
R1288 source.n102 source.n19 4.26717
R1289 source.n83 source.n27 4.26717
R1290 source.n54 source.n42 4.26717
R1291 source.n273 source.n146 4.26717
R1292 source.n244 source.n161 4.26717
R1293 source.n225 source.n169 4.26717
R1294 source.n196 source.n184 4.26717
R1295 source.n413 source.n286 4.26717
R1296 source.n384 source.n301 4.26717
R1297 source.n365 source.n309 4.26717
R1298 source.n336 source.n324 4.26717
R1299 source.n555 source.n428 4.26717
R1300 source.n526 source.n443 4.26717
R1301 source.n507 source.n451 4.26717
R1302 source.n478 source.n466 4.26717
R1303 source.n1044 source.n1043 3.49141
R1304 source.n1069 source.n1016 3.49141
R1305 source.n1090 source.n1004 3.49141
R1306 source.n1116 source.n1115 3.49141
R1307 source.n902 source.n901 3.49141
R1308 source.n927 source.n874 3.49141
R1309 source.n948 source.n862 3.49141
R1310 source.n974 source.n973 3.49141
R1311 source.n762 source.n761 3.49141
R1312 source.n787 source.n734 3.49141
R1313 source.n808 source.n722 3.49141
R1314 source.n834 source.n833 3.49141
R1315 source.n620 source.n619 3.49141
R1316 source.n645 source.n592 3.49141
R1317 source.n666 source.n580 3.49141
R1318 source.n692 source.n691 3.49141
R1319 source.n128 source.n127 3.49141
R1320 source.n103 source.n17 3.49141
R1321 source.n82 source.n29 3.49141
R1322 source.n58 source.n57 3.49141
R1323 source.n270 source.n269 3.49141
R1324 source.n245 source.n159 3.49141
R1325 source.n224 source.n171 3.49141
R1326 source.n200 source.n199 3.49141
R1327 source.n410 source.n409 3.49141
R1328 source.n385 source.n299 3.49141
R1329 source.n364 source.n311 3.49141
R1330 source.n340 source.n339 3.49141
R1331 source.n552 source.n551 3.49141
R1332 source.n527 source.n441 3.49141
R1333 source.n506 source.n453 3.49141
R1334 source.n482 source.n481 3.49141
R1335 source.n48 source.n47 2.84303
R1336 source.n190 source.n189 2.84303
R1337 source.n330 source.n329 2.84303
R1338 source.n472 source.n471 2.84303
R1339 source.n1034 source.n1033 2.84303
R1340 source.n892 source.n891 2.84303
R1341 source.n752 source.n751 2.84303
R1342 source.n610 source.n609 2.84303
R1343 source.n1047 source.n1026 2.71565
R1344 source.n1066 source.n1065 2.71565
R1345 source.n1094 source.n1093 2.71565
R1346 source.n1112 source.n994 2.71565
R1347 source.n905 source.n884 2.71565
R1348 source.n924 source.n923 2.71565
R1349 source.n952 source.n951 2.71565
R1350 source.n970 source.n852 2.71565
R1351 source.n765 source.n744 2.71565
R1352 source.n784 source.n783 2.71565
R1353 source.n812 source.n811 2.71565
R1354 source.n830 source.n712 2.71565
R1355 source.n623 source.n602 2.71565
R1356 source.n642 source.n641 2.71565
R1357 source.n670 source.n669 2.71565
R1358 source.n688 source.n570 2.71565
R1359 source.n124 source.n6 2.71565
R1360 source.n107 source.n106 2.71565
R1361 source.n79 source.n78 2.71565
R1362 source.n61 source.n40 2.71565
R1363 source.n266 source.n148 2.71565
R1364 source.n249 source.n248 2.71565
R1365 source.n221 source.n220 2.71565
R1366 source.n203 source.n182 2.71565
R1367 source.n406 source.n288 2.71565
R1368 source.n389 source.n388 2.71565
R1369 source.n361 source.n360 2.71565
R1370 source.n343 source.n322 2.71565
R1371 source.n548 source.n430 2.71565
R1372 source.n531 source.n530 2.71565
R1373 source.n503 source.n502 2.71565
R1374 source.n485 source.n464 2.71565
R1375 source.n1048 source.n1024 1.93989
R1376 source.n1062 source.n1018 1.93989
R1377 source.n1098 source.n1002 1.93989
R1378 source.n1111 source.n996 1.93989
R1379 source.n906 source.n882 1.93989
R1380 source.n920 source.n876 1.93989
R1381 source.n956 source.n860 1.93989
R1382 source.n969 source.n854 1.93989
R1383 source.n766 source.n742 1.93989
R1384 source.n780 source.n736 1.93989
R1385 source.n816 source.n720 1.93989
R1386 source.n829 source.n714 1.93989
R1387 source.n624 source.n600 1.93989
R1388 source.n638 source.n594 1.93989
R1389 source.n674 source.n578 1.93989
R1390 source.n687 source.n572 1.93989
R1391 source.n123 source.n8 1.93989
R1392 source.n110 source.n14 1.93989
R1393 source.n75 source.n31 1.93989
R1394 source.n62 source.n38 1.93989
R1395 source.n265 source.n150 1.93989
R1396 source.n252 source.n156 1.93989
R1397 source.n217 source.n173 1.93989
R1398 source.n204 source.n180 1.93989
R1399 source.n405 source.n290 1.93989
R1400 source.n392 source.n296 1.93989
R1401 source.n357 source.n313 1.93989
R1402 source.n344 source.n320 1.93989
R1403 source.n547 source.n432 1.93989
R1404 source.n534 source.n438 1.93989
R1405 source.n499 source.n455 1.93989
R1406 source.n486 source.n462 1.93989
R1407 source.n1053 source.n1051 1.16414
R1408 source.n1061 source.n1020 1.16414
R1409 source.n1099 source.n1000 1.16414
R1410 source.n1108 source.n1107 1.16414
R1411 source.n911 source.n909 1.16414
R1412 source.n919 source.n878 1.16414
R1413 source.n957 source.n858 1.16414
R1414 source.n966 source.n965 1.16414
R1415 source.n771 source.n769 1.16414
R1416 source.n779 source.n738 1.16414
R1417 source.n817 source.n718 1.16414
R1418 source.n826 source.n825 1.16414
R1419 source.n629 source.n627 1.16414
R1420 source.n637 source.n596 1.16414
R1421 source.n675 source.n576 1.16414
R1422 source.n684 source.n683 1.16414
R1423 source.n120 source.n119 1.16414
R1424 source.n111 source.n12 1.16414
R1425 source.n74 source.n33 1.16414
R1426 source.n66 source.n65 1.16414
R1427 source.n262 source.n261 1.16414
R1428 source.n253 source.n154 1.16414
R1429 source.n216 source.n175 1.16414
R1430 source.n208 source.n207 1.16414
R1431 source.n402 source.n401 1.16414
R1432 source.n393 source.n294 1.16414
R1433 source.n356 source.n315 1.16414
R1434 source.n348 source.n347 1.16414
R1435 source.n544 source.n543 1.16414
R1436 source.n535 source.n436 1.16414
R1437 source.n498 source.n457 1.16414
R1438 source.n490 source.n489 1.16414
R1439 source.n986 source.t2 0.7925
R1440 source.n986 source.t3 0.7925
R1441 source.n704 source.t6 0.7925
R1442 source.n704 source.t13 0.7925
R1443 source.n140 source.t12 0.7925
R1444 source.n140 source.t8 0.7925
R1445 source.n422 source.t14 0.7925
R1446 source.n422 source.t15 0.7925
R1447 source.n421 source.n281 0.470328
R1448 source.n985 source.n845 0.470328
R1449 source.n563 source.n423 0.457397
R1450 source.n423 source.n421 0.457397
R1451 source.n281 source.n141 0.457397
R1452 source.n141 source.n139 0.457397
R1453 source.n705 source.n703 0.457397
R1454 source.n845 source.n705 0.457397
R1455 source.n987 source.n985 0.457397
R1456 source.n1127 source.n987 0.457397
R1457 source.n1052 source.n1022 0.388379
R1458 source.n1058 source.n1057 0.388379
R1459 source.n1103 source.n1102 0.388379
R1460 source.n1104 source.n998 0.388379
R1461 source.n910 source.n880 0.388379
R1462 source.n916 source.n915 0.388379
R1463 source.n961 source.n960 0.388379
R1464 source.n962 source.n856 0.388379
R1465 source.n770 source.n740 0.388379
R1466 source.n776 source.n775 0.388379
R1467 source.n821 source.n820 0.388379
R1468 source.n822 source.n716 0.388379
R1469 source.n628 source.n598 0.388379
R1470 source.n634 source.n633 0.388379
R1471 source.n679 source.n678 0.388379
R1472 source.n680 source.n574 0.388379
R1473 source.n116 source.n10 0.388379
R1474 source.n115 source.n114 0.388379
R1475 source.n71 source.n70 0.388379
R1476 source.n37 source.n35 0.388379
R1477 source.n258 source.n152 0.388379
R1478 source.n257 source.n256 0.388379
R1479 source.n213 source.n212 0.388379
R1480 source.n179 source.n177 0.388379
R1481 source.n398 source.n292 0.388379
R1482 source.n397 source.n396 0.388379
R1483 source.n353 source.n352 0.388379
R1484 source.n319 source.n317 0.388379
R1485 source.n540 source.n434 0.388379
R1486 source.n539 source.n538 0.388379
R1487 source.n495 source.n494 0.388379
R1488 source.n461 source.n459 0.388379
R1489 source source.n1128 0.188
R1490 source.n1034 source.n1029 0.155672
R1491 source.n1041 source.n1029 0.155672
R1492 source.n1042 source.n1041 0.155672
R1493 source.n1042 source.n1025 0.155672
R1494 source.n1049 source.n1025 0.155672
R1495 source.n1050 source.n1049 0.155672
R1496 source.n1050 source.n1021 0.155672
R1497 source.n1059 source.n1021 0.155672
R1498 source.n1060 source.n1059 0.155672
R1499 source.n1060 source.n1017 0.155672
R1500 source.n1067 source.n1017 0.155672
R1501 source.n1068 source.n1067 0.155672
R1502 source.n1068 source.n1013 0.155672
R1503 source.n1075 source.n1013 0.155672
R1504 source.n1076 source.n1075 0.155672
R1505 source.n1076 source.n1009 0.155672
R1506 source.n1083 source.n1009 0.155672
R1507 source.n1084 source.n1083 0.155672
R1508 source.n1084 source.n1005 0.155672
R1509 source.n1091 source.n1005 0.155672
R1510 source.n1092 source.n1091 0.155672
R1511 source.n1092 source.n1001 0.155672
R1512 source.n1100 source.n1001 0.155672
R1513 source.n1101 source.n1100 0.155672
R1514 source.n1101 source.n997 0.155672
R1515 source.n1109 source.n997 0.155672
R1516 source.n1110 source.n1109 0.155672
R1517 source.n1110 source.n993 0.155672
R1518 source.n1117 source.n993 0.155672
R1519 source.n1118 source.n1117 0.155672
R1520 source.n1118 source.n989 0.155672
R1521 source.n1125 source.n989 0.155672
R1522 source.n892 source.n887 0.155672
R1523 source.n899 source.n887 0.155672
R1524 source.n900 source.n899 0.155672
R1525 source.n900 source.n883 0.155672
R1526 source.n907 source.n883 0.155672
R1527 source.n908 source.n907 0.155672
R1528 source.n908 source.n879 0.155672
R1529 source.n917 source.n879 0.155672
R1530 source.n918 source.n917 0.155672
R1531 source.n918 source.n875 0.155672
R1532 source.n925 source.n875 0.155672
R1533 source.n926 source.n925 0.155672
R1534 source.n926 source.n871 0.155672
R1535 source.n933 source.n871 0.155672
R1536 source.n934 source.n933 0.155672
R1537 source.n934 source.n867 0.155672
R1538 source.n941 source.n867 0.155672
R1539 source.n942 source.n941 0.155672
R1540 source.n942 source.n863 0.155672
R1541 source.n949 source.n863 0.155672
R1542 source.n950 source.n949 0.155672
R1543 source.n950 source.n859 0.155672
R1544 source.n958 source.n859 0.155672
R1545 source.n959 source.n958 0.155672
R1546 source.n959 source.n855 0.155672
R1547 source.n967 source.n855 0.155672
R1548 source.n968 source.n967 0.155672
R1549 source.n968 source.n851 0.155672
R1550 source.n975 source.n851 0.155672
R1551 source.n976 source.n975 0.155672
R1552 source.n976 source.n847 0.155672
R1553 source.n983 source.n847 0.155672
R1554 source.n752 source.n747 0.155672
R1555 source.n759 source.n747 0.155672
R1556 source.n760 source.n759 0.155672
R1557 source.n760 source.n743 0.155672
R1558 source.n767 source.n743 0.155672
R1559 source.n768 source.n767 0.155672
R1560 source.n768 source.n739 0.155672
R1561 source.n777 source.n739 0.155672
R1562 source.n778 source.n777 0.155672
R1563 source.n778 source.n735 0.155672
R1564 source.n785 source.n735 0.155672
R1565 source.n786 source.n785 0.155672
R1566 source.n786 source.n731 0.155672
R1567 source.n793 source.n731 0.155672
R1568 source.n794 source.n793 0.155672
R1569 source.n794 source.n727 0.155672
R1570 source.n801 source.n727 0.155672
R1571 source.n802 source.n801 0.155672
R1572 source.n802 source.n723 0.155672
R1573 source.n809 source.n723 0.155672
R1574 source.n810 source.n809 0.155672
R1575 source.n810 source.n719 0.155672
R1576 source.n818 source.n719 0.155672
R1577 source.n819 source.n818 0.155672
R1578 source.n819 source.n715 0.155672
R1579 source.n827 source.n715 0.155672
R1580 source.n828 source.n827 0.155672
R1581 source.n828 source.n711 0.155672
R1582 source.n835 source.n711 0.155672
R1583 source.n836 source.n835 0.155672
R1584 source.n836 source.n707 0.155672
R1585 source.n843 source.n707 0.155672
R1586 source.n610 source.n605 0.155672
R1587 source.n617 source.n605 0.155672
R1588 source.n618 source.n617 0.155672
R1589 source.n618 source.n601 0.155672
R1590 source.n625 source.n601 0.155672
R1591 source.n626 source.n625 0.155672
R1592 source.n626 source.n597 0.155672
R1593 source.n635 source.n597 0.155672
R1594 source.n636 source.n635 0.155672
R1595 source.n636 source.n593 0.155672
R1596 source.n643 source.n593 0.155672
R1597 source.n644 source.n643 0.155672
R1598 source.n644 source.n589 0.155672
R1599 source.n651 source.n589 0.155672
R1600 source.n652 source.n651 0.155672
R1601 source.n652 source.n585 0.155672
R1602 source.n659 source.n585 0.155672
R1603 source.n660 source.n659 0.155672
R1604 source.n660 source.n581 0.155672
R1605 source.n667 source.n581 0.155672
R1606 source.n668 source.n667 0.155672
R1607 source.n668 source.n577 0.155672
R1608 source.n676 source.n577 0.155672
R1609 source.n677 source.n676 0.155672
R1610 source.n677 source.n573 0.155672
R1611 source.n685 source.n573 0.155672
R1612 source.n686 source.n685 0.155672
R1613 source.n686 source.n569 0.155672
R1614 source.n693 source.n569 0.155672
R1615 source.n694 source.n693 0.155672
R1616 source.n694 source.n565 0.155672
R1617 source.n701 source.n565 0.155672
R1618 source.n137 source.n1 0.155672
R1619 source.n130 source.n1 0.155672
R1620 source.n130 source.n129 0.155672
R1621 source.n129 source.n5 0.155672
R1622 source.n122 source.n5 0.155672
R1623 source.n122 source.n121 0.155672
R1624 source.n121 source.n9 0.155672
R1625 source.n113 source.n9 0.155672
R1626 source.n113 source.n112 0.155672
R1627 source.n112 source.n13 0.155672
R1628 source.n105 source.n13 0.155672
R1629 source.n105 source.n104 0.155672
R1630 source.n104 source.n18 0.155672
R1631 source.n97 source.n18 0.155672
R1632 source.n97 source.n96 0.155672
R1633 source.n96 source.n22 0.155672
R1634 source.n89 source.n22 0.155672
R1635 source.n89 source.n88 0.155672
R1636 source.n88 source.n26 0.155672
R1637 source.n81 source.n26 0.155672
R1638 source.n81 source.n80 0.155672
R1639 source.n80 source.n30 0.155672
R1640 source.n73 source.n30 0.155672
R1641 source.n73 source.n72 0.155672
R1642 source.n72 source.n34 0.155672
R1643 source.n64 source.n34 0.155672
R1644 source.n64 source.n63 0.155672
R1645 source.n63 source.n39 0.155672
R1646 source.n56 source.n39 0.155672
R1647 source.n56 source.n55 0.155672
R1648 source.n55 source.n43 0.155672
R1649 source.n48 source.n43 0.155672
R1650 source.n279 source.n143 0.155672
R1651 source.n272 source.n143 0.155672
R1652 source.n272 source.n271 0.155672
R1653 source.n271 source.n147 0.155672
R1654 source.n264 source.n147 0.155672
R1655 source.n264 source.n263 0.155672
R1656 source.n263 source.n151 0.155672
R1657 source.n255 source.n151 0.155672
R1658 source.n255 source.n254 0.155672
R1659 source.n254 source.n155 0.155672
R1660 source.n247 source.n155 0.155672
R1661 source.n247 source.n246 0.155672
R1662 source.n246 source.n160 0.155672
R1663 source.n239 source.n160 0.155672
R1664 source.n239 source.n238 0.155672
R1665 source.n238 source.n164 0.155672
R1666 source.n231 source.n164 0.155672
R1667 source.n231 source.n230 0.155672
R1668 source.n230 source.n168 0.155672
R1669 source.n223 source.n168 0.155672
R1670 source.n223 source.n222 0.155672
R1671 source.n222 source.n172 0.155672
R1672 source.n215 source.n172 0.155672
R1673 source.n215 source.n214 0.155672
R1674 source.n214 source.n176 0.155672
R1675 source.n206 source.n176 0.155672
R1676 source.n206 source.n205 0.155672
R1677 source.n205 source.n181 0.155672
R1678 source.n198 source.n181 0.155672
R1679 source.n198 source.n197 0.155672
R1680 source.n197 source.n185 0.155672
R1681 source.n190 source.n185 0.155672
R1682 source.n419 source.n283 0.155672
R1683 source.n412 source.n283 0.155672
R1684 source.n412 source.n411 0.155672
R1685 source.n411 source.n287 0.155672
R1686 source.n404 source.n287 0.155672
R1687 source.n404 source.n403 0.155672
R1688 source.n403 source.n291 0.155672
R1689 source.n395 source.n291 0.155672
R1690 source.n395 source.n394 0.155672
R1691 source.n394 source.n295 0.155672
R1692 source.n387 source.n295 0.155672
R1693 source.n387 source.n386 0.155672
R1694 source.n386 source.n300 0.155672
R1695 source.n379 source.n300 0.155672
R1696 source.n379 source.n378 0.155672
R1697 source.n378 source.n304 0.155672
R1698 source.n371 source.n304 0.155672
R1699 source.n371 source.n370 0.155672
R1700 source.n370 source.n308 0.155672
R1701 source.n363 source.n308 0.155672
R1702 source.n363 source.n362 0.155672
R1703 source.n362 source.n312 0.155672
R1704 source.n355 source.n312 0.155672
R1705 source.n355 source.n354 0.155672
R1706 source.n354 source.n316 0.155672
R1707 source.n346 source.n316 0.155672
R1708 source.n346 source.n345 0.155672
R1709 source.n345 source.n321 0.155672
R1710 source.n338 source.n321 0.155672
R1711 source.n338 source.n337 0.155672
R1712 source.n337 source.n325 0.155672
R1713 source.n330 source.n325 0.155672
R1714 source.n561 source.n425 0.155672
R1715 source.n554 source.n425 0.155672
R1716 source.n554 source.n553 0.155672
R1717 source.n553 source.n429 0.155672
R1718 source.n546 source.n429 0.155672
R1719 source.n546 source.n545 0.155672
R1720 source.n545 source.n433 0.155672
R1721 source.n537 source.n433 0.155672
R1722 source.n537 source.n536 0.155672
R1723 source.n536 source.n437 0.155672
R1724 source.n529 source.n437 0.155672
R1725 source.n529 source.n528 0.155672
R1726 source.n528 source.n442 0.155672
R1727 source.n521 source.n442 0.155672
R1728 source.n521 source.n520 0.155672
R1729 source.n520 source.n446 0.155672
R1730 source.n513 source.n446 0.155672
R1731 source.n513 source.n512 0.155672
R1732 source.n512 source.n450 0.155672
R1733 source.n505 source.n450 0.155672
R1734 source.n505 source.n504 0.155672
R1735 source.n504 source.n454 0.155672
R1736 source.n497 source.n454 0.155672
R1737 source.n497 source.n496 0.155672
R1738 source.n496 source.n458 0.155672
R1739 source.n488 source.n458 0.155672
R1740 source.n488 source.n487 0.155672
R1741 source.n487 source.n463 0.155672
R1742 source.n480 source.n463 0.155672
R1743 source.n480 source.n479 0.155672
R1744 source.n479 source.n467 0.155672
R1745 source.n472 source.n467 0.155672
R1746 minus.n5 minus.t7 3212.24
R1747 minus.n1 minus.t6 3212.24
R1748 minus.n12 minus.t4 3212.24
R1749 minus.n8 minus.t2 3212.24
R1750 minus.n4 minus.t0 3169.15
R1751 minus.n2 minus.t3 3169.15
R1752 minus.n11 minus.t1 3169.15
R1753 minus.n9 minus.t5 3169.15
R1754 minus.n1 minus.n0 161.489
R1755 minus.n8 minus.n7 161.489
R1756 minus.n6 minus.n5 161.3
R1757 minus.n3 minus.n0 161.3
R1758 minus.n13 minus.n12 161.3
R1759 minus.n10 minus.n7 161.3
R1760 minus.n14 minus.n6 43.6331
R1761 minus.n4 minus.n3 38.7066
R1762 minus.n3 minus.n2 38.7066
R1763 minus.n10 minus.n9 38.7066
R1764 minus.n11 minus.n10 38.7066
R1765 minus.n5 minus.n4 34.3247
R1766 minus.n2 minus.n1 34.3247
R1767 minus.n9 minus.n8 34.3247
R1768 minus.n12 minus.n11 34.3247
R1769 minus.n14 minus.n13 6.44368
R1770 minus.n6 minus.n0 0.189894
R1771 minus.n13 minus.n7 0.189894
R1772 minus minus.n14 0.188
R1773 drain_right.n5 drain_right.n3 59.1722
R1774 drain_right.n2 drain_right.n1 58.8885
R1775 drain_right.n2 drain_right.n0 58.8885
R1776 drain_right.n5 drain_right.n4 58.7154
R1777 drain_right drain_right.n2 38.2615
R1778 drain_right drain_right.n5 6.11011
R1779 drain_right.n1 drain_right.t6 0.7925
R1780 drain_right.n1 drain_right.t3 0.7925
R1781 drain_right.n0 drain_right.t5 0.7925
R1782 drain_right.n0 drain_right.t2 0.7925
R1783 drain_right.n3 drain_right.t4 0.7925
R1784 drain_right.n3 drain_right.t1 0.7925
R1785 drain_right.n4 drain_right.t0 0.7925
R1786 drain_right.n4 drain_right.t7 0.7925
C0 source drain_left 39.0398f
C1 drain_right source 39.0384f
C2 minus drain_left 0.17017f
C3 minus drain_right 5.10044f
C4 plus drain_left 5.21724f
C5 plus drain_right 0.269775f
C6 minus source 4.01737f
C7 plus source 4.03141f
C8 plus minus 7.11575f
C9 drain_right drain_left 0.58123f
C10 drain_right a_n1246_n5888# 9.00316f
C11 drain_left a_n1246_n5888# 9.19771f
C12 source a_n1246_n5888# 15.417097f
C13 minus a_n1246_n5888# 5.669911f
C14 plus a_n1246_n5888# 8.80105f
C15 drain_right.t5 a_n1246_n5888# 0.755784f
C16 drain_right.t2 a_n1246_n5888# 0.755784f
C17 drain_right.n0 a_n1246_n5888# 6.966609f
C18 drain_right.t6 a_n1246_n5888# 0.755784f
C19 drain_right.t3 a_n1246_n5888# 0.755784f
C20 drain_right.n1 a_n1246_n5888# 6.966609f
C21 drain_right.n2 a_n1246_n5888# 3.64191f
C22 drain_right.t4 a_n1246_n5888# 0.755784f
C23 drain_right.t1 a_n1246_n5888# 0.755784f
C24 drain_right.n3 a_n1246_n5888# 6.96884f
C25 drain_right.t0 a_n1246_n5888# 0.755784f
C26 drain_right.t7 a_n1246_n5888# 0.755784f
C27 drain_right.n4 a_n1246_n5888# 6.96537f
C28 drain_right.n5 a_n1246_n5888# 1.19707f
C29 minus.n0 a_n1246_n5888# 0.130515f
C30 minus.t7 a_n1246_n5888# 0.847462f
C31 minus.t0 a_n1246_n5888# 0.843266f
C32 minus.t3 a_n1246_n5888# 0.843266f
C33 minus.t6 a_n1246_n5888# 0.847462f
C34 minus.n1 a_n1246_n5888# 0.3297f
C35 minus.n2 a_n1246_n5888# 0.313005f
C36 minus.n3 a_n1246_n5888# 0.020993f
C37 minus.n4 a_n1246_n5888# 0.313005f
C38 minus.n5 a_n1246_n5888# 0.329617f
C39 minus.n6 a_n1246_n5888# 2.80465f
C40 minus.n7 a_n1246_n5888# 0.130515f
C41 minus.t1 a_n1246_n5888# 0.843266f
C42 minus.t5 a_n1246_n5888# 0.843266f
C43 minus.t2 a_n1246_n5888# 0.847462f
C44 minus.n8 a_n1246_n5888# 0.3297f
C45 minus.n9 a_n1246_n5888# 0.313005f
C46 minus.n10 a_n1246_n5888# 0.020993f
C47 minus.n11 a_n1246_n5888# 0.313005f
C48 minus.t4 a_n1246_n5888# 0.847462f
C49 minus.n12 a_n1246_n5888# 0.329617f
C50 minus.n13 a_n1246_n5888# 0.383901f
C51 minus.n14 a_n1246_n5888# 3.3355f
C52 source.n0 a_n1246_n5888# 0.036277f
C53 source.n1 a_n1246_n5888# 0.026315f
C54 source.n2 a_n1246_n5888# 0.01414f
C55 source.n3 a_n1246_n5888# 0.033423f
C56 source.n4 a_n1246_n5888# 0.014972f
C57 source.n5 a_n1246_n5888# 0.026315f
C58 source.n6 a_n1246_n5888# 0.01414f
C59 source.n7 a_n1246_n5888# 0.033423f
C60 source.n8 a_n1246_n5888# 0.014972f
C61 source.n9 a_n1246_n5888# 0.026315f
C62 source.n10 a_n1246_n5888# 0.01414f
C63 source.n11 a_n1246_n5888# 0.033423f
C64 source.n12 a_n1246_n5888# 0.014972f
C65 source.n13 a_n1246_n5888# 0.026315f
C66 source.n14 a_n1246_n5888# 0.01414f
C67 source.n15 a_n1246_n5888# 0.033423f
C68 source.n16 a_n1246_n5888# 0.033423f
C69 source.n17 a_n1246_n5888# 0.014972f
C70 source.n18 a_n1246_n5888# 0.026315f
C71 source.n19 a_n1246_n5888# 0.01414f
C72 source.n20 a_n1246_n5888# 0.033423f
C73 source.n21 a_n1246_n5888# 0.014972f
C74 source.n22 a_n1246_n5888# 0.026315f
C75 source.n23 a_n1246_n5888# 0.01414f
C76 source.n24 a_n1246_n5888# 0.033423f
C77 source.n25 a_n1246_n5888# 0.014972f
C78 source.n26 a_n1246_n5888# 0.026315f
C79 source.n27 a_n1246_n5888# 0.01414f
C80 source.n28 a_n1246_n5888# 0.033423f
C81 source.n29 a_n1246_n5888# 0.014972f
C82 source.n30 a_n1246_n5888# 0.026315f
C83 source.n31 a_n1246_n5888# 0.01414f
C84 source.n32 a_n1246_n5888# 0.033423f
C85 source.n33 a_n1246_n5888# 0.014972f
C86 source.n34 a_n1246_n5888# 0.026315f
C87 source.n35 a_n1246_n5888# 0.014556f
C88 source.n36 a_n1246_n5888# 0.033423f
C89 source.n37 a_n1246_n5888# 0.01414f
C90 source.n38 a_n1246_n5888# 0.014972f
C91 source.n39 a_n1246_n5888# 0.026315f
C92 source.n40 a_n1246_n5888# 0.01414f
C93 source.n41 a_n1246_n5888# 0.033423f
C94 source.n42 a_n1246_n5888# 0.014972f
C95 source.n43 a_n1246_n5888# 0.026315f
C96 source.n44 a_n1246_n5888# 0.01414f
C97 source.n45 a_n1246_n5888# 0.025067f
C98 source.n46 a_n1246_n5888# 0.023627f
C99 source.t10 a_n1246_n5888# 0.058291f
C100 source.n47 a_n1246_n5888# 0.32106f
C101 source.n48 a_n1246_n5888# 2.8491f
C102 source.n49 a_n1246_n5888# 0.01414f
C103 source.n50 a_n1246_n5888# 0.014972f
C104 source.n51 a_n1246_n5888# 0.033423f
C105 source.n52 a_n1246_n5888# 0.033423f
C106 source.n53 a_n1246_n5888# 0.014972f
C107 source.n54 a_n1246_n5888# 0.01414f
C108 source.n55 a_n1246_n5888# 0.026315f
C109 source.n56 a_n1246_n5888# 0.026315f
C110 source.n57 a_n1246_n5888# 0.01414f
C111 source.n58 a_n1246_n5888# 0.014972f
C112 source.n59 a_n1246_n5888# 0.033423f
C113 source.n60 a_n1246_n5888# 0.033423f
C114 source.n61 a_n1246_n5888# 0.014972f
C115 source.n62 a_n1246_n5888# 0.01414f
C116 source.n63 a_n1246_n5888# 0.026315f
C117 source.n64 a_n1246_n5888# 0.026315f
C118 source.n65 a_n1246_n5888# 0.01414f
C119 source.n66 a_n1246_n5888# 0.014972f
C120 source.n67 a_n1246_n5888# 0.033423f
C121 source.n68 a_n1246_n5888# 0.033423f
C122 source.n69 a_n1246_n5888# 0.033423f
C123 source.n70 a_n1246_n5888# 0.014556f
C124 source.n71 a_n1246_n5888# 0.01414f
C125 source.n72 a_n1246_n5888# 0.026315f
C126 source.n73 a_n1246_n5888# 0.026315f
C127 source.n74 a_n1246_n5888# 0.01414f
C128 source.n75 a_n1246_n5888# 0.014972f
C129 source.n76 a_n1246_n5888# 0.033423f
C130 source.n77 a_n1246_n5888# 0.033423f
C131 source.n78 a_n1246_n5888# 0.014972f
C132 source.n79 a_n1246_n5888# 0.01414f
C133 source.n80 a_n1246_n5888# 0.026315f
C134 source.n81 a_n1246_n5888# 0.026315f
C135 source.n82 a_n1246_n5888# 0.01414f
C136 source.n83 a_n1246_n5888# 0.014972f
C137 source.n84 a_n1246_n5888# 0.033423f
C138 source.n85 a_n1246_n5888# 0.033423f
C139 source.n86 a_n1246_n5888# 0.014972f
C140 source.n87 a_n1246_n5888# 0.01414f
C141 source.n88 a_n1246_n5888# 0.026315f
C142 source.n89 a_n1246_n5888# 0.026315f
C143 source.n90 a_n1246_n5888# 0.01414f
C144 source.n91 a_n1246_n5888# 0.014972f
C145 source.n92 a_n1246_n5888# 0.033423f
C146 source.n93 a_n1246_n5888# 0.033423f
C147 source.n94 a_n1246_n5888# 0.014972f
C148 source.n95 a_n1246_n5888# 0.01414f
C149 source.n96 a_n1246_n5888# 0.026315f
C150 source.n97 a_n1246_n5888# 0.026315f
C151 source.n98 a_n1246_n5888# 0.01414f
C152 source.n99 a_n1246_n5888# 0.014972f
C153 source.n100 a_n1246_n5888# 0.033423f
C154 source.n101 a_n1246_n5888# 0.033423f
C155 source.n102 a_n1246_n5888# 0.014972f
C156 source.n103 a_n1246_n5888# 0.01414f
C157 source.n104 a_n1246_n5888# 0.026315f
C158 source.n105 a_n1246_n5888# 0.026315f
C159 source.n106 a_n1246_n5888# 0.01414f
C160 source.n107 a_n1246_n5888# 0.014972f
C161 source.n108 a_n1246_n5888# 0.033423f
C162 source.n109 a_n1246_n5888# 0.033423f
C163 source.n110 a_n1246_n5888# 0.014972f
C164 source.n111 a_n1246_n5888# 0.01414f
C165 source.n112 a_n1246_n5888# 0.026315f
C166 source.n113 a_n1246_n5888# 0.026315f
C167 source.n114 a_n1246_n5888# 0.01414f
C168 source.n115 a_n1246_n5888# 0.014556f
C169 source.n116 a_n1246_n5888# 0.014556f
C170 source.n117 a_n1246_n5888# 0.033423f
C171 source.n118 a_n1246_n5888# 0.033423f
C172 source.n119 a_n1246_n5888# 0.014972f
C173 source.n120 a_n1246_n5888# 0.01414f
C174 source.n121 a_n1246_n5888# 0.026315f
C175 source.n122 a_n1246_n5888# 0.026315f
C176 source.n123 a_n1246_n5888# 0.01414f
C177 source.n124 a_n1246_n5888# 0.014972f
C178 source.n125 a_n1246_n5888# 0.033423f
C179 source.n126 a_n1246_n5888# 0.033423f
C180 source.n127 a_n1246_n5888# 0.014972f
C181 source.n128 a_n1246_n5888# 0.01414f
C182 source.n129 a_n1246_n5888# 0.026315f
C183 source.n130 a_n1246_n5888# 0.026315f
C184 source.n131 a_n1246_n5888# 0.01414f
C185 source.n132 a_n1246_n5888# 0.014972f
C186 source.n133 a_n1246_n5888# 0.033423f
C187 source.n134 a_n1246_n5888# 0.071098f
C188 source.n135 a_n1246_n5888# 0.014972f
C189 source.n136 a_n1246_n5888# 0.01414f
C190 source.n137 a_n1246_n5888# 0.057949f
C191 source.n138 a_n1246_n5888# 0.039563f
C192 source.n139 a_n1246_n5888# 2.0568f
C193 source.t12 a_n1246_n5888# 0.519865f
C194 source.t8 a_n1246_n5888# 0.519865f
C195 source.n140 a_n1246_n5888# 4.70485f
C196 source.n141 a_n1246_n5888# 0.350417f
C197 source.n142 a_n1246_n5888# 0.036277f
C198 source.n143 a_n1246_n5888# 0.026315f
C199 source.n144 a_n1246_n5888# 0.01414f
C200 source.n145 a_n1246_n5888# 0.033423f
C201 source.n146 a_n1246_n5888# 0.014972f
C202 source.n147 a_n1246_n5888# 0.026315f
C203 source.n148 a_n1246_n5888# 0.01414f
C204 source.n149 a_n1246_n5888# 0.033423f
C205 source.n150 a_n1246_n5888# 0.014972f
C206 source.n151 a_n1246_n5888# 0.026315f
C207 source.n152 a_n1246_n5888# 0.01414f
C208 source.n153 a_n1246_n5888# 0.033423f
C209 source.n154 a_n1246_n5888# 0.014972f
C210 source.n155 a_n1246_n5888# 0.026315f
C211 source.n156 a_n1246_n5888# 0.01414f
C212 source.n157 a_n1246_n5888# 0.033423f
C213 source.n158 a_n1246_n5888# 0.033423f
C214 source.n159 a_n1246_n5888# 0.014972f
C215 source.n160 a_n1246_n5888# 0.026315f
C216 source.n161 a_n1246_n5888# 0.01414f
C217 source.n162 a_n1246_n5888# 0.033423f
C218 source.n163 a_n1246_n5888# 0.014972f
C219 source.n164 a_n1246_n5888# 0.026315f
C220 source.n165 a_n1246_n5888# 0.01414f
C221 source.n166 a_n1246_n5888# 0.033423f
C222 source.n167 a_n1246_n5888# 0.014972f
C223 source.n168 a_n1246_n5888# 0.026315f
C224 source.n169 a_n1246_n5888# 0.01414f
C225 source.n170 a_n1246_n5888# 0.033423f
C226 source.n171 a_n1246_n5888# 0.014972f
C227 source.n172 a_n1246_n5888# 0.026315f
C228 source.n173 a_n1246_n5888# 0.01414f
C229 source.n174 a_n1246_n5888# 0.033423f
C230 source.n175 a_n1246_n5888# 0.014972f
C231 source.n176 a_n1246_n5888# 0.026315f
C232 source.n177 a_n1246_n5888# 0.014556f
C233 source.n178 a_n1246_n5888# 0.033423f
C234 source.n179 a_n1246_n5888# 0.01414f
C235 source.n180 a_n1246_n5888# 0.014972f
C236 source.n181 a_n1246_n5888# 0.026315f
C237 source.n182 a_n1246_n5888# 0.01414f
C238 source.n183 a_n1246_n5888# 0.033423f
C239 source.n184 a_n1246_n5888# 0.014972f
C240 source.n185 a_n1246_n5888# 0.026315f
C241 source.n186 a_n1246_n5888# 0.01414f
C242 source.n187 a_n1246_n5888# 0.025067f
C243 source.n188 a_n1246_n5888# 0.023627f
C244 source.t11 a_n1246_n5888# 0.058291f
C245 source.n189 a_n1246_n5888# 0.32106f
C246 source.n190 a_n1246_n5888# 2.8491f
C247 source.n191 a_n1246_n5888# 0.01414f
C248 source.n192 a_n1246_n5888# 0.014972f
C249 source.n193 a_n1246_n5888# 0.033423f
C250 source.n194 a_n1246_n5888# 0.033423f
C251 source.n195 a_n1246_n5888# 0.014972f
C252 source.n196 a_n1246_n5888# 0.01414f
C253 source.n197 a_n1246_n5888# 0.026315f
C254 source.n198 a_n1246_n5888# 0.026315f
C255 source.n199 a_n1246_n5888# 0.01414f
C256 source.n200 a_n1246_n5888# 0.014972f
C257 source.n201 a_n1246_n5888# 0.033423f
C258 source.n202 a_n1246_n5888# 0.033423f
C259 source.n203 a_n1246_n5888# 0.014972f
C260 source.n204 a_n1246_n5888# 0.01414f
C261 source.n205 a_n1246_n5888# 0.026315f
C262 source.n206 a_n1246_n5888# 0.026315f
C263 source.n207 a_n1246_n5888# 0.01414f
C264 source.n208 a_n1246_n5888# 0.014972f
C265 source.n209 a_n1246_n5888# 0.033423f
C266 source.n210 a_n1246_n5888# 0.033423f
C267 source.n211 a_n1246_n5888# 0.033423f
C268 source.n212 a_n1246_n5888# 0.014556f
C269 source.n213 a_n1246_n5888# 0.01414f
C270 source.n214 a_n1246_n5888# 0.026315f
C271 source.n215 a_n1246_n5888# 0.026315f
C272 source.n216 a_n1246_n5888# 0.01414f
C273 source.n217 a_n1246_n5888# 0.014972f
C274 source.n218 a_n1246_n5888# 0.033423f
C275 source.n219 a_n1246_n5888# 0.033423f
C276 source.n220 a_n1246_n5888# 0.014972f
C277 source.n221 a_n1246_n5888# 0.01414f
C278 source.n222 a_n1246_n5888# 0.026315f
C279 source.n223 a_n1246_n5888# 0.026315f
C280 source.n224 a_n1246_n5888# 0.01414f
C281 source.n225 a_n1246_n5888# 0.014972f
C282 source.n226 a_n1246_n5888# 0.033423f
C283 source.n227 a_n1246_n5888# 0.033423f
C284 source.n228 a_n1246_n5888# 0.014972f
C285 source.n229 a_n1246_n5888# 0.01414f
C286 source.n230 a_n1246_n5888# 0.026315f
C287 source.n231 a_n1246_n5888# 0.026315f
C288 source.n232 a_n1246_n5888# 0.01414f
C289 source.n233 a_n1246_n5888# 0.014972f
C290 source.n234 a_n1246_n5888# 0.033423f
C291 source.n235 a_n1246_n5888# 0.033423f
C292 source.n236 a_n1246_n5888# 0.014972f
C293 source.n237 a_n1246_n5888# 0.01414f
C294 source.n238 a_n1246_n5888# 0.026315f
C295 source.n239 a_n1246_n5888# 0.026315f
C296 source.n240 a_n1246_n5888# 0.01414f
C297 source.n241 a_n1246_n5888# 0.014972f
C298 source.n242 a_n1246_n5888# 0.033423f
C299 source.n243 a_n1246_n5888# 0.033423f
C300 source.n244 a_n1246_n5888# 0.014972f
C301 source.n245 a_n1246_n5888# 0.01414f
C302 source.n246 a_n1246_n5888# 0.026315f
C303 source.n247 a_n1246_n5888# 0.026315f
C304 source.n248 a_n1246_n5888# 0.01414f
C305 source.n249 a_n1246_n5888# 0.014972f
C306 source.n250 a_n1246_n5888# 0.033423f
C307 source.n251 a_n1246_n5888# 0.033423f
C308 source.n252 a_n1246_n5888# 0.014972f
C309 source.n253 a_n1246_n5888# 0.01414f
C310 source.n254 a_n1246_n5888# 0.026315f
C311 source.n255 a_n1246_n5888# 0.026315f
C312 source.n256 a_n1246_n5888# 0.01414f
C313 source.n257 a_n1246_n5888# 0.014556f
C314 source.n258 a_n1246_n5888# 0.014556f
C315 source.n259 a_n1246_n5888# 0.033423f
C316 source.n260 a_n1246_n5888# 0.033423f
C317 source.n261 a_n1246_n5888# 0.014972f
C318 source.n262 a_n1246_n5888# 0.01414f
C319 source.n263 a_n1246_n5888# 0.026315f
C320 source.n264 a_n1246_n5888# 0.026315f
C321 source.n265 a_n1246_n5888# 0.01414f
C322 source.n266 a_n1246_n5888# 0.014972f
C323 source.n267 a_n1246_n5888# 0.033423f
C324 source.n268 a_n1246_n5888# 0.033423f
C325 source.n269 a_n1246_n5888# 0.014972f
C326 source.n270 a_n1246_n5888# 0.01414f
C327 source.n271 a_n1246_n5888# 0.026315f
C328 source.n272 a_n1246_n5888# 0.026315f
C329 source.n273 a_n1246_n5888# 0.01414f
C330 source.n274 a_n1246_n5888# 0.014972f
C331 source.n275 a_n1246_n5888# 0.033423f
C332 source.n276 a_n1246_n5888# 0.071098f
C333 source.n277 a_n1246_n5888# 0.014972f
C334 source.n278 a_n1246_n5888# 0.01414f
C335 source.n279 a_n1246_n5888# 0.057949f
C336 source.n280 a_n1246_n5888# 0.039563f
C337 source.n281 a_n1246_n5888# 0.099432f
C338 source.n282 a_n1246_n5888# 0.036277f
C339 source.n283 a_n1246_n5888# 0.026315f
C340 source.n284 a_n1246_n5888# 0.01414f
C341 source.n285 a_n1246_n5888# 0.033423f
C342 source.n286 a_n1246_n5888# 0.014972f
C343 source.n287 a_n1246_n5888# 0.026315f
C344 source.n288 a_n1246_n5888# 0.01414f
C345 source.n289 a_n1246_n5888# 0.033423f
C346 source.n290 a_n1246_n5888# 0.014972f
C347 source.n291 a_n1246_n5888# 0.026315f
C348 source.n292 a_n1246_n5888# 0.01414f
C349 source.n293 a_n1246_n5888# 0.033423f
C350 source.n294 a_n1246_n5888# 0.014972f
C351 source.n295 a_n1246_n5888# 0.026315f
C352 source.n296 a_n1246_n5888# 0.01414f
C353 source.n297 a_n1246_n5888# 0.033423f
C354 source.n298 a_n1246_n5888# 0.033423f
C355 source.n299 a_n1246_n5888# 0.014972f
C356 source.n300 a_n1246_n5888# 0.026315f
C357 source.n301 a_n1246_n5888# 0.01414f
C358 source.n302 a_n1246_n5888# 0.033423f
C359 source.n303 a_n1246_n5888# 0.014972f
C360 source.n304 a_n1246_n5888# 0.026315f
C361 source.n305 a_n1246_n5888# 0.01414f
C362 source.n306 a_n1246_n5888# 0.033423f
C363 source.n307 a_n1246_n5888# 0.014972f
C364 source.n308 a_n1246_n5888# 0.026315f
C365 source.n309 a_n1246_n5888# 0.01414f
C366 source.n310 a_n1246_n5888# 0.033423f
C367 source.n311 a_n1246_n5888# 0.014972f
C368 source.n312 a_n1246_n5888# 0.026315f
C369 source.n313 a_n1246_n5888# 0.01414f
C370 source.n314 a_n1246_n5888# 0.033423f
C371 source.n315 a_n1246_n5888# 0.014972f
C372 source.n316 a_n1246_n5888# 0.026315f
C373 source.n317 a_n1246_n5888# 0.014556f
C374 source.n318 a_n1246_n5888# 0.033423f
C375 source.n319 a_n1246_n5888# 0.01414f
C376 source.n320 a_n1246_n5888# 0.014972f
C377 source.n321 a_n1246_n5888# 0.026315f
C378 source.n322 a_n1246_n5888# 0.01414f
C379 source.n323 a_n1246_n5888# 0.033423f
C380 source.n324 a_n1246_n5888# 0.014972f
C381 source.n325 a_n1246_n5888# 0.026315f
C382 source.n326 a_n1246_n5888# 0.01414f
C383 source.n327 a_n1246_n5888# 0.025067f
C384 source.n328 a_n1246_n5888# 0.023627f
C385 source.t5 a_n1246_n5888# 0.058291f
C386 source.n329 a_n1246_n5888# 0.32106f
C387 source.n330 a_n1246_n5888# 2.8491f
C388 source.n331 a_n1246_n5888# 0.01414f
C389 source.n332 a_n1246_n5888# 0.014972f
C390 source.n333 a_n1246_n5888# 0.033423f
C391 source.n334 a_n1246_n5888# 0.033423f
C392 source.n335 a_n1246_n5888# 0.014972f
C393 source.n336 a_n1246_n5888# 0.01414f
C394 source.n337 a_n1246_n5888# 0.026315f
C395 source.n338 a_n1246_n5888# 0.026315f
C396 source.n339 a_n1246_n5888# 0.01414f
C397 source.n340 a_n1246_n5888# 0.014972f
C398 source.n341 a_n1246_n5888# 0.033423f
C399 source.n342 a_n1246_n5888# 0.033423f
C400 source.n343 a_n1246_n5888# 0.014972f
C401 source.n344 a_n1246_n5888# 0.01414f
C402 source.n345 a_n1246_n5888# 0.026315f
C403 source.n346 a_n1246_n5888# 0.026315f
C404 source.n347 a_n1246_n5888# 0.01414f
C405 source.n348 a_n1246_n5888# 0.014972f
C406 source.n349 a_n1246_n5888# 0.033423f
C407 source.n350 a_n1246_n5888# 0.033423f
C408 source.n351 a_n1246_n5888# 0.033423f
C409 source.n352 a_n1246_n5888# 0.014556f
C410 source.n353 a_n1246_n5888# 0.01414f
C411 source.n354 a_n1246_n5888# 0.026315f
C412 source.n355 a_n1246_n5888# 0.026315f
C413 source.n356 a_n1246_n5888# 0.01414f
C414 source.n357 a_n1246_n5888# 0.014972f
C415 source.n358 a_n1246_n5888# 0.033423f
C416 source.n359 a_n1246_n5888# 0.033423f
C417 source.n360 a_n1246_n5888# 0.014972f
C418 source.n361 a_n1246_n5888# 0.01414f
C419 source.n362 a_n1246_n5888# 0.026315f
C420 source.n363 a_n1246_n5888# 0.026315f
C421 source.n364 a_n1246_n5888# 0.01414f
C422 source.n365 a_n1246_n5888# 0.014972f
C423 source.n366 a_n1246_n5888# 0.033423f
C424 source.n367 a_n1246_n5888# 0.033423f
C425 source.n368 a_n1246_n5888# 0.014972f
C426 source.n369 a_n1246_n5888# 0.01414f
C427 source.n370 a_n1246_n5888# 0.026315f
C428 source.n371 a_n1246_n5888# 0.026315f
C429 source.n372 a_n1246_n5888# 0.01414f
C430 source.n373 a_n1246_n5888# 0.014972f
C431 source.n374 a_n1246_n5888# 0.033423f
C432 source.n375 a_n1246_n5888# 0.033423f
C433 source.n376 a_n1246_n5888# 0.014972f
C434 source.n377 a_n1246_n5888# 0.01414f
C435 source.n378 a_n1246_n5888# 0.026315f
C436 source.n379 a_n1246_n5888# 0.026315f
C437 source.n380 a_n1246_n5888# 0.01414f
C438 source.n381 a_n1246_n5888# 0.014972f
C439 source.n382 a_n1246_n5888# 0.033423f
C440 source.n383 a_n1246_n5888# 0.033423f
C441 source.n384 a_n1246_n5888# 0.014972f
C442 source.n385 a_n1246_n5888# 0.01414f
C443 source.n386 a_n1246_n5888# 0.026315f
C444 source.n387 a_n1246_n5888# 0.026315f
C445 source.n388 a_n1246_n5888# 0.01414f
C446 source.n389 a_n1246_n5888# 0.014972f
C447 source.n390 a_n1246_n5888# 0.033423f
C448 source.n391 a_n1246_n5888# 0.033423f
C449 source.n392 a_n1246_n5888# 0.014972f
C450 source.n393 a_n1246_n5888# 0.01414f
C451 source.n394 a_n1246_n5888# 0.026315f
C452 source.n395 a_n1246_n5888# 0.026315f
C453 source.n396 a_n1246_n5888# 0.01414f
C454 source.n397 a_n1246_n5888# 0.014556f
C455 source.n398 a_n1246_n5888# 0.014556f
C456 source.n399 a_n1246_n5888# 0.033423f
C457 source.n400 a_n1246_n5888# 0.033423f
C458 source.n401 a_n1246_n5888# 0.014972f
C459 source.n402 a_n1246_n5888# 0.01414f
C460 source.n403 a_n1246_n5888# 0.026315f
C461 source.n404 a_n1246_n5888# 0.026315f
C462 source.n405 a_n1246_n5888# 0.01414f
C463 source.n406 a_n1246_n5888# 0.014972f
C464 source.n407 a_n1246_n5888# 0.033423f
C465 source.n408 a_n1246_n5888# 0.033423f
C466 source.n409 a_n1246_n5888# 0.014972f
C467 source.n410 a_n1246_n5888# 0.01414f
C468 source.n411 a_n1246_n5888# 0.026315f
C469 source.n412 a_n1246_n5888# 0.026315f
C470 source.n413 a_n1246_n5888# 0.01414f
C471 source.n414 a_n1246_n5888# 0.014972f
C472 source.n415 a_n1246_n5888# 0.033423f
C473 source.n416 a_n1246_n5888# 0.071098f
C474 source.n417 a_n1246_n5888# 0.014972f
C475 source.n418 a_n1246_n5888# 0.01414f
C476 source.n419 a_n1246_n5888# 0.057949f
C477 source.n420 a_n1246_n5888# 0.039563f
C478 source.n421 a_n1246_n5888# 0.099432f
C479 source.t14 a_n1246_n5888# 0.519865f
C480 source.t15 a_n1246_n5888# 0.519865f
C481 source.n422 a_n1246_n5888# 4.70485f
C482 source.n423 a_n1246_n5888# 0.350417f
C483 source.n424 a_n1246_n5888# 0.036277f
C484 source.n425 a_n1246_n5888# 0.026315f
C485 source.n426 a_n1246_n5888# 0.01414f
C486 source.n427 a_n1246_n5888# 0.033423f
C487 source.n428 a_n1246_n5888# 0.014972f
C488 source.n429 a_n1246_n5888# 0.026315f
C489 source.n430 a_n1246_n5888# 0.01414f
C490 source.n431 a_n1246_n5888# 0.033423f
C491 source.n432 a_n1246_n5888# 0.014972f
C492 source.n433 a_n1246_n5888# 0.026315f
C493 source.n434 a_n1246_n5888# 0.01414f
C494 source.n435 a_n1246_n5888# 0.033423f
C495 source.n436 a_n1246_n5888# 0.014972f
C496 source.n437 a_n1246_n5888# 0.026315f
C497 source.n438 a_n1246_n5888# 0.01414f
C498 source.n439 a_n1246_n5888# 0.033423f
C499 source.n440 a_n1246_n5888# 0.033423f
C500 source.n441 a_n1246_n5888# 0.014972f
C501 source.n442 a_n1246_n5888# 0.026315f
C502 source.n443 a_n1246_n5888# 0.01414f
C503 source.n444 a_n1246_n5888# 0.033423f
C504 source.n445 a_n1246_n5888# 0.014972f
C505 source.n446 a_n1246_n5888# 0.026315f
C506 source.n447 a_n1246_n5888# 0.01414f
C507 source.n448 a_n1246_n5888# 0.033423f
C508 source.n449 a_n1246_n5888# 0.014972f
C509 source.n450 a_n1246_n5888# 0.026315f
C510 source.n451 a_n1246_n5888# 0.01414f
C511 source.n452 a_n1246_n5888# 0.033423f
C512 source.n453 a_n1246_n5888# 0.014972f
C513 source.n454 a_n1246_n5888# 0.026315f
C514 source.n455 a_n1246_n5888# 0.01414f
C515 source.n456 a_n1246_n5888# 0.033423f
C516 source.n457 a_n1246_n5888# 0.014972f
C517 source.n458 a_n1246_n5888# 0.026315f
C518 source.n459 a_n1246_n5888# 0.014556f
C519 source.n460 a_n1246_n5888# 0.033423f
C520 source.n461 a_n1246_n5888# 0.01414f
C521 source.n462 a_n1246_n5888# 0.014972f
C522 source.n463 a_n1246_n5888# 0.026315f
C523 source.n464 a_n1246_n5888# 0.01414f
C524 source.n465 a_n1246_n5888# 0.033423f
C525 source.n466 a_n1246_n5888# 0.014972f
C526 source.n467 a_n1246_n5888# 0.026315f
C527 source.n468 a_n1246_n5888# 0.01414f
C528 source.n469 a_n1246_n5888# 0.025067f
C529 source.n470 a_n1246_n5888# 0.023627f
C530 source.t4 a_n1246_n5888# 0.058291f
C531 source.n471 a_n1246_n5888# 0.32106f
C532 source.n472 a_n1246_n5888# 2.8491f
C533 source.n473 a_n1246_n5888# 0.01414f
C534 source.n474 a_n1246_n5888# 0.014972f
C535 source.n475 a_n1246_n5888# 0.033423f
C536 source.n476 a_n1246_n5888# 0.033423f
C537 source.n477 a_n1246_n5888# 0.014972f
C538 source.n478 a_n1246_n5888# 0.01414f
C539 source.n479 a_n1246_n5888# 0.026315f
C540 source.n480 a_n1246_n5888# 0.026315f
C541 source.n481 a_n1246_n5888# 0.01414f
C542 source.n482 a_n1246_n5888# 0.014972f
C543 source.n483 a_n1246_n5888# 0.033423f
C544 source.n484 a_n1246_n5888# 0.033423f
C545 source.n485 a_n1246_n5888# 0.014972f
C546 source.n486 a_n1246_n5888# 0.01414f
C547 source.n487 a_n1246_n5888# 0.026315f
C548 source.n488 a_n1246_n5888# 0.026315f
C549 source.n489 a_n1246_n5888# 0.01414f
C550 source.n490 a_n1246_n5888# 0.014972f
C551 source.n491 a_n1246_n5888# 0.033423f
C552 source.n492 a_n1246_n5888# 0.033423f
C553 source.n493 a_n1246_n5888# 0.033423f
C554 source.n494 a_n1246_n5888# 0.014556f
C555 source.n495 a_n1246_n5888# 0.01414f
C556 source.n496 a_n1246_n5888# 0.026315f
C557 source.n497 a_n1246_n5888# 0.026315f
C558 source.n498 a_n1246_n5888# 0.01414f
C559 source.n499 a_n1246_n5888# 0.014972f
C560 source.n500 a_n1246_n5888# 0.033423f
C561 source.n501 a_n1246_n5888# 0.033423f
C562 source.n502 a_n1246_n5888# 0.014972f
C563 source.n503 a_n1246_n5888# 0.01414f
C564 source.n504 a_n1246_n5888# 0.026315f
C565 source.n505 a_n1246_n5888# 0.026315f
C566 source.n506 a_n1246_n5888# 0.01414f
C567 source.n507 a_n1246_n5888# 0.014972f
C568 source.n508 a_n1246_n5888# 0.033423f
C569 source.n509 a_n1246_n5888# 0.033423f
C570 source.n510 a_n1246_n5888# 0.014972f
C571 source.n511 a_n1246_n5888# 0.01414f
C572 source.n512 a_n1246_n5888# 0.026315f
C573 source.n513 a_n1246_n5888# 0.026315f
C574 source.n514 a_n1246_n5888# 0.01414f
C575 source.n515 a_n1246_n5888# 0.014972f
C576 source.n516 a_n1246_n5888# 0.033423f
C577 source.n517 a_n1246_n5888# 0.033423f
C578 source.n518 a_n1246_n5888# 0.014972f
C579 source.n519 a_n1246_n5888# 0.01414f
C580 source.n520 a_n1246_n5888# 0.026315f
C581 source.n521 a_n1246_n5888# 0.026315f
C582 source.n522 a_n1246_n5888# 0.01414f
C583 source.n523 a_n1246_n5888# 0.014972f
C584 source.n524 a_n1246_n5888# 0.033423f
C585 source.n525 a_n1246_n5888# 0.033423f
C586 source.n526 a_n1246_n5888# 0.014972f
C587 source.n527 a_n1246_n5888# 0.01414f
C588 source.n528 a_n1246_n5888# 0.026315f
C589 source.n529 a_n1246_n5888# 0.026315f
C590 source.n530 a_n1246_n5888# 0.01414f
C591 source.n531 a_n1246_n5888# 0.014972f
C592 source.n532 a_n1246_n5888# 0.033423f
C593 source.n533 a_n1246_n5888# 0.033423f
C594 source.n534 a_n1246_n5888# 0.014972f
C595 source.n535 a_n1246_n5888# 0.01414f
C596 source.n536 a_n1246_n5888# 0.026315f
C597 source.n537 a_n1246_n5888# 0.026315f
C598 source.n538 a_n1246_n5888# 0.01414f
C599 source.n539 a_n1246_n5888# 0.014556f
C600 source.n540 a_n1246_n5888# 0.014556f
C601 source.n541 a_n1246_n5888# 0.033423f
C602 source.n542 a_n1246_n5888# 0.033423f
C603 source.n543 a_n1246_n5888# 0.014972f
C604 source.n544 a_n1246_n5888# 0.01414f
C605 source.n545 a_n1246_n5888# 0.026315f
C606 source.n546 a_n1246_n5888# 0.026315f
C607 source.n547 a_n1246_n5888# 0.01414f
C608 source.n548 a_n1246_n5888# 0.014972f
C609 source.n549 a_n1246_n5888# 0.033423f
C610 source.n550 a_n1246_n5888# 0.033423f
C611 source.n551 a_n1246_n5888# 0.014972f
C612 source.n552 a_n1246_n5888# 0.01414f
C613 source.n553 a_n1246_n5888# 0.026315f
C614 source.n554 a_n1246_n5888# 0.026315f
C615 source.n555 a_n1246_n5888# 0.01414f
C616 source.n556 a_n1246_n5888# 0.014972f
C617 source.n557 a_n1246_n5888# 0.033423f
C618 source.n558 a_n1246_n5888# 0.071098f
C619 source.n559 a_n1246_n5888# 0.014972f
C620 source.n560 a_n1246_n5888# 0.01414f
C621 source.n561 a_n1246_n5888# 0.057949f
C622 source.n562 a_n1246_n5888# 0.039563f
C623 source.n563 a_n1246_n5888# 2.54032f
C624 source.n564 a_n1246_n5888# 0.036277f
C625 source.n565 a_n1246_n5888# 0.026315f
C626 source.n566 a_n1246_n5888# 0.01414f
C627 source.n567 a_n1246_n5888# 0.033423f
C628 source.n568 a_n1246_n5888# 0.014972f
C629 source.n569 a_n1246_n5888# 0.026315f
C630 source.n570 a_n1246_n5888# 0.01414f
C631 source.n571 a_n1246_n5888# 0.033423f
C632 source.n572 a_n1246_n5888# 0.014972f
C633 source.n573 a_n1246_n5888# 0.026315f
C634 source.n574 a_n1246_n5888# 0.01414f
C635 source.n575 a_n1246_n5888# 0.033423f
C636 source.n576 a_n1246_n5888# 0.014972f
C637 source.n577 a_n1246_n5888# 0.026315f
C638 source.n578 a_n1246_n5888# 0.01414f
C639 source.n579 a_n1246_n5888# 0.033423f
C640 source.n580 a_n1246_n5888# 0.014972f
C641 source.n581 a_n1246_n5888# 0.026315f
C642 source.n582 a_n1246_n5888# 0.01414f
C643 source.n583 a_n1246_n5888# 0.033423f
C644 source.n584 a_n1246_n5888# 0.014972f
C645 source.n585 a_n1246_n5888# 0.026315f
C646 source.n586 a_n1246_n5888# 0.01414f
C647 source.n587 a_n1246_n5888# 0.033423f
C648 source.n588 a_n1246_n5888# 0.014972f
C649 source.n589 a_n1246_n5888# 0.026315f
C650 source.n590 a_n1246_n5888# 0.01414f
C651 source.n591 a_n1246_n5888# 0.033423f
C652 source.n592 a_n1246_n5888# 0.014972f
C653 source.n593 a_n1246_n5888# 0.026315f
C654 source.n594 a_n1246_n5888# 0.01414f
C655 source.n595 a_n1246_n5888# 0.033423f
C656 source.n596 a_n1246_n5888# 0.014972f
C657 source.n597 a_n1246_n5888# 0.026315f
C658 source.n598 a_n1246_n5888# 0.014556f
C659 source.n599 a_n1246_n5888# 0.033423f
C660 source.n600 a_n1246_n5888# 0.014972f
C661 source.n601 a_n1246_n5888# 0.026315f
C662 source.n602 a_n1246_n5888# 0.01414f
C663 source.n603 a_n1246_n5888# 0.033423f
C664 source.n604 a_n1246_n5888# 0.014972f
C665 source.n605 a_n1246_n5888# 0.026315f
C666 source.n606 a_n1246_n5888# 0.01414f
C667 source.n607 a_n1246_n5888# 0.025067f
C668 source.n608 a_n1246_n5888# 0.023627f
C669 source.t9 a_n1246_n5888# 0.058291f
C670 source.n609 a_n1246_n5888# 0.32106f
C671 source.n610 a_n1246_n5888# 2.8491f
C672 source.n611 a_n1246_n5888# 0.01414f
C673 source.n612 a_n1246_n5888# 0.014972f
C674 source.n613 a_n1246_n5888# 0.033423f
C675 source.n614 a_n1246_n5888# 0.033423f
C676 source.n615 a_n1246_n5888# 0.014972f
C677 source.n616 a_n1246_n5888# 0.01414f
C678 source.n617 a_n1246_n5888# 0.026315f
C679 source.n618 a_n1246_n5888# 0.026315f
C680 source.n619 a_n1246_n5888# 0.01414f
C681 source.n620 a_n1246_n5888# 0.014972f
C682 source.n621 a_n1246_n5888# 0.033423f
C683 source.n622 a_n1246_n5888# 0.033423f
C684 source.n623 a_n1246_n5888# 0.014972f
C685 source.n624 a_n1246_n5888# 0.01414f
C686 source.n625 a_n1246_n5888# 0.026315f
C687 source.n626 a_n1246_n5888# 0.026315f
C688 source.n627 a_n1246_n5888# 0.01414f
C689 source.n628 a_n1246_n5888# 0.01414f
C690 source.n629 a_n1246_n5888# 0.014972f
C691 source.n630 a_n1246_n5888# 0.033423f
C692 source.n631 a_n1246_n5888# 0.033423f
C693 source.n632 a_n1246_n5888# 0.033423f
C694 source.n633 a_n1246_n5888# 0.014556f
C695 source.n634 a_n1246_n5888# 0.01414f
C696 source.n635 a_n1246_n5888# 0.026315f
C697 source.n636 a_n1246_n5888# 0.026315f
C698 source.n637 a_n1246_n5888# 0.01414f
C699 source.n638 a_n1246_n5888# 0.014972f
C700 source.n639 a_n1246_n5888# 0.033423f
C701 source.n640 a_n1246_n5888# 0.033423f
C702 source.n641 a_n1246_n5888# 0.014972f
C703 source.n642 a_n1246_n5888# 0.01414f
C704 source.n643 a_n1246_n5888# 0.026315f
C705 source.n644 a_n1246_n5888# 0.026315f
C706 source.n645 a_n1246_n5888# 0.01414f
C707 source.n646 a_n1246_n5888# 0.014972f
C708 source.n647 a_n1246_n5888# 0.033423f
C709 source.n648 a_n1246_n5888# 0.033423f
C710 source.n649 a_n1246_n5888# 0.014972f
C711 source.n650 a_n1246_n5888# 0.01414f
C712 source.n651 a_n1246_n5888# 0.026315f
C713 source.n652 a_n1246_n5888# 0.026315f
C714 source.n653 a_n1246_n5888# 0.01414f
C715 source.n654 a_n1246_n5888# 0.014972f
C716 source.n655 a_n1246_n5888# 0.033423f
C717 source.n656 a_n1246_n5888# 0.033423f
C718 source.n657 a_n1246_n5888# 0.014972f
C719 source.n658 a_n1246_n5888# 0.01414f
C720 source.n659 a_n1246_n5888# 0.026315f
C721 source.n660 a_n1246_n5888# 0.026315f
C722 source.n661 a_n1246_n5888# 0.01414f
C723 source.n662 a_n1246_n5888# 0.014972f
C724 source.n663 a_n1246_n5888# 0.033423f
C725 source.n664 a_n1246_n5888# 0.033423f
C726 source.n665 a_n1246_n5888# 0.014972f
C727 source.n666 a_n1246_n5888# 0.01414f
C728 source.n667 a_n1246_n5888# 0.026315f
C729 source.n668 a_n1246_n5888# 0.026315f
C730 source.n669 a_n1246_n5888# 0.01414f
C731 source.n670 a_n1246_n5888# 0.014972f
C732 source.n671 a_n1246_n5888# 0.033423f
C733 source.n672 a_n1246_n5888# 0.033423f
C734 source.n673 a_n1246_n5888# 0.033423f
C735 source.n674 a_n1246_n5888# 0.014972f
C736 source.n675 a_n1246_n5888# 0.01414f
C737 source.n676 a_n1246_n5888# 0.026315f
C738 source.n677 a_n1246_n5888# 0.026315f
C739 source.n678 a_n1246_n5888# 0.01414f
C740 source.n679 a_n1246_n5888# 0.014556f
C741 source.n680 a_n1246_n5888# 0.014556f
C742 source.n681 a_n1246_n5888# 0.033423f
C743 source.n682 a_n1246_n5888# 0.033423f
C744 source.n683 a_n1246_n5888# 0.014972f
C745 source.n684 a_n1246_n5888# 0.01414f
C746 source.n685 a_n1246_n5888# 0.026315f
C747 source.n686 a_n1246_n5888# 0.026315f
C748 source.n687 a_n1246_n5888# 0.01414f
C749 source.n688 a_n1246_n5888# 0.014972f
C750 source.n689 a_n1246_n5888# 0.033423f
C751 source.n690 a_n1246_n5888# 0.033423f
C752 source.n691 a_n1246_n5888# 0.014972f
C753 source.n692 a_n1246_n5888# 0.01414f
C754 source.n693 a_n1246_n5888# 0.026315f
C755 source.n694 a_n1246_n5888# 0.026315f
C756 source.n695 a_n1246_n5888# 0.01414f
C757 source.n696 a_n1246_n5888# 0.014972f
C758 source.n697 a_n1246_n5888# 0.033423f
C759 source.n698 a_n1246_n5888# 0.071098f
C760 source.n699 a_n1246_n5888# 0.014972f
C761 source.n700 a_n1246_n5888# 0.01414f
C762 source.n701 a_n1246_n5888# 0.057949f
C763 source.n702 a_n1246_n5888# 0.039563f
C764 source.n703 a_n1246_n5888# 2.54032f
C765 source.t6 a_n1246_n5888# 0.519865f
C766 source.t13 a_n1246_n5888# 0.519865f
C767 source.n704 a_n1246_n5888# 4.70485f
C768 source.n705 a_n1246_n5888# 0.350419f
C769 source.n706 a_n1246_n5888# 0.036277f
C770 source.n707 a_n1246_n5888# 0.026315f
C771 source.n708 a_n1246_n5888# 0.01414f
C772 source.n709 a_n1246_n5888# 0.033423f
C773 source.n710 a_n1246_n5888# 0.014972f
C774 source.n711 a_n1246_n5888# 0.026315f
C775 source.n712 a_n1246_n5888# 0.01414f
C776 source.n713 a_n1246_n5888# 0.033423f
C777 source.n714 a_n1246_n5888# 0.014972f
C778 source.n715 a_n1246_n5888# 0.026315f
C779 source.n716 a_n1246_n5888# 0.01414f
C780 source.n717 a_n1246_n5888# 0.033423f
C781 source.n718 a_n1246_n5888# 0.014972f
C782 source.n719 a_n1246_n5888# 0.026315f
C783 source.n720 a_n1246_n5888# 0.01414f
C784 source.n721 a_n1246_n5888# 0.033423f
C785 source.n722 a_n1246_n5888# 0.014972f
C786 source.n723 a_n1246_n5888# 0.026315f
C787 source.n724 a_n1246_n5888# 0.01414f
C788 source.n725 a_n1246_n5888# 0.033423f
C789 source.n726 a_n1246_n5888# 0.014972f
C790 source.n727 a_n1246_n5888# 0.026315f
C791 source.n728 a_n1246_n5888# 0.01414f
C792 source.n729 a_n1246_n5888# 0.033423f
C793 source.n730 a_n1246_n5888# 0.014972f
C794 source.n731 a_n1246_n5888# 0.026315f
C795 source.n732 a_n1246_n5888# 0.01414f
C796 source.n733 a_n1246_n5888# 0.033423f
C797 source.n734 a_n1246_n5888# 0.014972f
C798 source.n735 a_n1246_n5888# 0.026315f
C799 source.n736 a_n1246_n5888# 0.01414f
C800 source.n737 a_n1246_n5888# 0.033423f
C801 source.n738 a_n1246_n5888# 0.014972f
C802 source.n739 a_n1246_n5888# 0.026315f
C803 source.n740 a_n1246_n5888# 0.014556f
C804 source.n741 a_n1246_n5888# 0.033423f
C805 source.n742 a_n1246_n5888# 0.014972f
C806 source.n743 a_n1246_n5888# 0.026315f
C807 source.n744 a_n1246_n5888# 0.01414f
C808 source.n745 a_n1246_n5888# 0.033423f
C809 source.n746 a_n1246_n5888# 0.014972f
C810 source.n747 a_n1246_n5888# 0.026315f
C811 source.n748 a_n1246_n5888# 0.01414f
C812 source.n749 a_n1246_n5888# 0.025067f
C813 source.n750 a_n1246_n5888# 0.023627f
C814 source.t7 a_n1246_n5888# 0.058291f
C815 source.n751 a_n1246_n5888# 0.32106f
C816 source.n752 a_n1246_n5888# 2.8491f
C817 source.n753 a_n1246_n5888# 0.01414f
C818 source.n754 a_n1246_n5888# 0.014972f
C819 source.n755 a_n1246_n5888# 0.033423f
C820 source.n756 a_n1246_n5888# 0.033423f
C821 source.n757 a_n1246_n5888# 0.014972f
C822 source.n758 a_n1246_n5888# 0.01414f
C823 source.n759 a_n1246_n5888# 0.026315f
C824 source.n760 a_n1246_n5888# 0.026315f
C825 source.n761 a_n1246_n5888# 0.01414f
C826 source.n762 a_n1246_n5888# 0.014972f
C827 source.n763 a_n1246_n5888# 0.033423f
C828 source.n764 a_n1246_n5888# 0.033423f
C829 source.n765 a_n1246_n5888# 0.014972f
C830 source.n766 a_n1246_n5888# 0.01414f
C831 source.n767 a_n1246_n5888# 0.026315f
C832 source.n768 a_n1246_n5888# 0.026315f
C833 source.n769 a_n1246_n5888# 0.01414f
C834 source.n770 a_n1246_n5888# 0.01414f
C835 source.n771 a_n1246_n5888# 0.014972f
C836 source.n772 a_n1246_n5888# 0.033423f
C837 source.n773 a_n1246_n5888# 0.033423f
C838 source.n774 a_n1246_n5888# 0.033423f
C839 source.n775 a_n1246_n5888# 0.014556f
C840 source.n776 a_n1246_n5888# 0.01414f
C841 source.n777 a_n1246_n5888# 0.026315f
C842 source.n778 a_n1246_n5888# 0.026315f
C843 source.n779 a_n1246_n5888# 0.01414f
C844 source.n780 a_n1246_n5888# 0.014972f
C845 source.n781 a_n1246_n5888# 0.033423f
C846 source.n782 a_n1246_n5888# 0.033423f
C847 source.n783 a_n1246_n5888# 0.014972f
C848 source.n784 a_n1246_n5888# 0.01414f
C849 source.n785 a_n1246_n5888# 0.026315f
C850 source.n786 a_n1246_n5888# 0.026315f
C851 source.n787 a_n1246_n5888# 0.01414f
C852 source.n788 a_n1246_n5888# 0.014972f
C853 source.n789 a_n1246_n5888# 0.033423f
C854 source.n790 a_n1246_n5888# 0.033423f
C855 source.n791 a_n1246_n5888# 0.014972f
C856 source.n792 a_n1246_n5888# 0.01414f
C857 source.n793 a_n1246_n5888# 0.026315f
C858 source.n794 a_n1246_n5888# 0.026315f
C859 source.n795 a_n1246_n5888# 0.01414f
C860 source.n796 a_n1246_n5888# 0.014972f
C861 source.n797 a_n1246_n5888# 0.033423f
C862 source.n798 a_n1246_n5888# 0.033423f
C863 source.n799 a_n1246_n5888# 0.014972f
C864 source.n800 a_n1246_n5888# 0.01414f
C865 source.n801 a_n1246_n5888# 0.026315f
C866 source.n802 a_n1246_n5888# 0.026315f
C867 source.n803 a_n1246_n5888# 0.01414f
C868 source.n804 a_n1246_n5888# 0.014972f
C869 source.n805 a_n1246_n5888# 0.033423f
C870 source.n806 a_n1246_n5888# 0.033423f
C871 source.n807 a_n1246_n5888# 0.014972f
C872 source.n808 a_n1246_n5888# 0.01414f
C873 source.n809 a_n1246_n5888# 0.026315f
C874 source.n810 a_n1246_n5888# 0.026315f
C875 source.n811 a_n1246_n5888# 0.01414f
C876 source.n812 a_n1246_n5888# 0.014972f
C877 source.n813 a_n1246_n5888# 0.033423f
C878 source.n814 a_n1246_n5888# 0.033423f
C879 source.n815 a_n1246_n5888# 0.033423f
C880 source.n816 a_n1246_n5888# 0.014972f
C881 source.n817 a_n1246_n5888# 0.01414f
C882 source.n818 a_n1246_n5888# 0.026315f
C883 source.n819 a_n1246_n5888# 0.026315f
C884 source.n820 a_n1246_n5888# 0.01414f
C885 source.n821 a_n1246_n5888# 0.014556f
C886 source.n822 a_n1246_n5888# 0.014556f
C887 source.n823 a_n1246_n5888# 0.033423f
C888 source.n824 a_n1246_n5888# 0.033423f
C889 source.n825 a_n1246_n5888# 0.014972f
C890 source.n826 a_n1246_n5888# 0.01414f
C891 source.n827 a_n1246_n5888# 0.026315f
C892 source.n828 a_n1246_n5888# 0.026315f
C893 source.n829 a_n1246_n5888# 0.01414f
C894 source.n830 a_n1246_n5888# 0.014972f
C895 source.n831 a_n1246_n5888# 0.033423f
C896 source.n832 a_n1246_n5888# 0.033423f
C897 source.n833 a_n1246_n5888# 0.014972f
C898 source.n834 a_n1246_n5888# 0.01414f
C899 source.n835 a_n1246_n5888# 0.026315f
C900 source.n836 a_n1246_n5888# 0.026315f
C901 source.n837 a_n1246_n5888# 0.01414f
C902 source.n838 a_n1246_n5888# 0.014972f
C903 source.n839 a_n1246_n5888# 0.033423f
C904 source.n840 a_n1246_n5888# 0.071098f
C905 source.n841 a_n1246_n5888# 0.014972f
C906 source.n842 a_n1246_n5888# 0.01414f
C907 source.n843 a_n1246_n5888# 0.057949f
C908 source.n844 a_n1246_n5888# 0.039563f
C909 source.n845 a_n1246_n5888# 0.099432f
C910 source.n846 a_n1246_n5888# 0.036277f
C911 source.n847 a_n1246_n5888# 0.026315f
C912 source.n848 a_n1246_n5888# 0.01414f
C913 source.n849 a_n1246_n5888# 0.033423f
C914 source.n850 a_n1246_n5888# 0.014972f
C915 source.n851 a_n1246_n5888# 0.026315f
C916 source.n852 a_n1246_n5888# 0.01414f
C917 source.n853 a_n1246_n5888# 0.033423f
C918 source.n854 a_n1246_n5888# 0.014972f
C919 source.n855 a_n1246_n5888# 0.026315f
C920 source.n856 a_n1246_n5888# 0.01414f
C921 source.n857 a_n1246_n5888# 0.033423f
C922 source.n858 a_n1246_n5888# 0.014972f
C923 source.n859 a_n1246_n5888# 0.026315f
C924 source.n860 a_n1246_n5888# 0.01414f
C925 source.n861 a_n1246_n5888# 0.033423f
C926 source.n862 a_n1246_n5888# 0.014972f
C927 source.n863 a_n1246_n5888# 0.026315f
C928 source.n864 a_n1246_n5888# 0.01414f
C929 source.n865 a_n1246_n5888# 0.033423f
C930 source.n866 a_n1246_n5888# 0.014972f
C931 source.n867 a_n1246_n5888# 0.026315f
C932 source.n868 a_n1246_n5888# 0.01414f
C933 source.n869 a_n1246_n5888# 0.033423f
C934 source.n870 a_n1246_n5888# 0.014972f
C935 source.n871 a_n1246_n5888# 0.026315f
C936 source.n872 a_n1246_n5888# 0.01414f
C937 source.n873 a_n1246_n5888# 0.033423f
C938 source.n874 a_n1246_n5888# 0.014972f
C939 source.n875 a_n1246_n5888# 0.026315f
C940 source.n876 a_n1246_n5888# 0.01414f
C941 source.n877 a_n1246_n5888# 0.033423f
C942 source.n878 a_n1246_n5888# 0.014972f
C943 source.n879 a_n1246_n5888# 0.026315f
C944 source.n880 a_n1246_n5888# 0.014556f
C945 source.n881 a_n1246_n5888# 0.033423f
C946 source.n882 a_n1246_n5888# 0.014972f
C947 source.n883 a_n1246_n5888# 0.026315f
C948 source.n884 a_n1246_n5888# 0.01414f
C949 source.n885 a_n1246_n5888# 0.033423f
C950 source.n886 a_n1246_n5888# 0.014972f
C951 source.n887 a_n1246_n5888# 0.026315f
C952 source.n888 a_n1246_n5888# 0.01414f
C953 source.n889 a_n1246_n5888# 0.025067f
C954 source.n890 a_n1246_n5888# 0.023627f
C955 source.t0 a_n1246_n5888# 0.058291f
C956 source.n891 a_n1246_n5888# 0.32106f
C957 source.n892 a_n1246_n5888# 2.8491f
C958 source.n893 a_n1246_n5888# 0.01414f
C959 source.n894 a_n1246_n5888# 0.014972f
C960 source.n895 a_n1246_n5888# 0.033423f
C961 source.n896 a_n1246_n5888# 0.033423f
C962 source.n897 a_n1246_n5888# 0.014972f
C963 source.n898 a_n1246_n5888# 0.01414f
C964 source.n899 a_n1246_n5888# 0.026315f
C965 source.n900 a_n1246_n5888# 0.026315f
C966 source.n901 a_n1246_n5888# 0.01414f
C967 source.n902 a_n1246_n5888# 0.014972f
C968 source.n903 a_n1246_n5888# 0.033423f
C969 source.n904 a_n1246_n5888# 0.033423f
C970 source.n905 a_n1246_n5888# 0.014972f
C971 source.n906 a_n1246_n5888# 0.01414f
C972 source.n907 a_n1246_n5888# 0.026315f
C973 source.n908 a_n1246_n5888# 0.026315f
C974 source.n909 a_n1246_n5888# 0.01414f
C975 source.n910 a_n1246_n5888# 0.01414f
C976 source.n911 a_n1246_n5888# 0.014972f
C977 source.n912 a_n1246_n5888# 0.033423f
C978 source.n913 a_n1246_n5888# 0.033423f
C979 source.n914 a_n1246_n5888# 0.033423f
C980 source.n915 a_n1246_n5888# 0.014556f
C981 source.n916 a_n1246_n5888# 0.01414f
C982 source.n917 a_n1246_n5888# 0.026315f
C983 source.n918 a_n1246_n5888# 0.026315f
C984 source.n919 a_n1246_n5888# 0.01414f
C985 source.n920 a_n1246_n5888# 0.014972f
C986 source.n921 a_n1246_n5888# 0.033423f
C987 source.n922 a_n1246_n5888# 0.033423f
C988 source.n923 a_n1246_n5888# 0.014972f
C989 source.n924 a_n1246_n5888# 0.01414f
C990 source.n925 a_n1246_n5888# 0.026315f
C991 source.n926 a_n1246_n5888# 0.026315f
C992 source.n927 a_n1246_n5888# 0.01414f
C993 source.n928 a_n1246_n5888# 0.014972f
C994 source.n929 a_n1246_n5888# 0.033423f
C995 source.n930 a_n1246_n5888# 0.033423f
C996 source.n931 a_n1246_n5888# 0.014972f
C997 source.n932 a_n1246_n5888# 0.01414f
C998 source.n933 a_n1246_n5888# 0.026315f
C999 source.n934 a_n1246_n5888# 0.026315f
C1000 source.n935 a_n1246_n5888# 0.01414f
C1001 source.n936 a_n1246_n5888# 0.014972f
C1002 source.n937 a_n1246_n5888# 0.033423f
C1003 source.n938 a_n1246_n5888# 0.033423f
C1004 source.n939 a_n1246_n5888# 0.014972f
C1005 source.n940 a_n1246_n5888# 0.01414f
C1006 source.n941 a_n1246_n5888# 0.026315f
C1007 source.n942 a_n1246_n5888# 0.026315f
C1008 source.n943 a_n1246_n5888# 0.01414f
C1009 source.n944 a_n1246_n5888# 0.014972f
C1010 source.n945 a_n1246_n5888# 0.033423f
C1011 source.n946 a_n1246_n5888# 0.033423f
C1012 source.n947 a_n1246_n5888# 0.014972f
C1013 source.n948 a_n1246_n5888# 0.01414f
C1014 source.n949 a_n1246_n5888# 0.026315f
C1015 source.n950 a_n1246_n5888# 0.026315f
C1016 source.n951 a_n1246_n5888# 0.01414f
C1017 source.n952 a_n1246_n5888# 0.014972f
C1018 source.n953 a_n1246_n5888# 0.033423f
C1019 source.n954 a_n1246_n5888# 0.033423f
C1020 source.n955 a_n1246_n5888# 0.033423f
C1021 source.n956 a_n1246_n5888# 0.014972f
C1022 source.n957 a_n1246_n5888# 0.01414f
C1023 source.n958 a_n1246_n5888# 0.026315f
C1024 source.n959 a_n1246_n5888# 0.026315f
C1025 source.n960 a_n1246_n5888# 0.01414f
C1026 source.n961 a_n1246_n5888# 0.014556f
C1027 source.n962 a_n1246_n5888# 0.014556f
C1028 source.n963 a_n1246_n5888# 0.033423f
C1029 source.n964 a_n1246_n5888# 0.033423f
C1030 source.n965 a_n1246_n5888# 0.014972f
C1031 source.n966 a_n1246_n5888# 0.01414f
C1032 source.n967 a_n1246_n5888# 0.026315f
C1033 source.n968 a_n1246_n5888# 0.026315f
C1034 source.n969 a_n1246_n5888# 0.01414f
C1035 source.n970 a_n1246_n5888# 0.014972f
C1036 source.n971 a_n1246_n5888# 0.033423f
C1037 source.n972 a_n1246_n5888# 0.033423f
C1038 source.n973 a_n1246_n5888# 0.014972f
C1039 source.n974 a_n1246_n5888# 0.01414f
C1040 source.n975 a_n1246_n5888# 0.026315f
C1041 source.n976 a_n1246_n5888# 0.026315f
C1042 source.n977 a_n1246_n5888# 0.01414f
C1043 source.n978 a_n1246_n5888# 0.014972f
C1044 source.n979 a_n1246_n5888# 0.033423f
C1045 source.n980 a_n1246_n5888# 0.071098f
C1046 source.n981 a_n1246_n5888# 0.014972f
C1047 source.n982 a_n1246_n5888# 0.01414f
C1048 source.n983 a_n1246_n5888# 0.057949f
C1049 source.n984 a_n1246_n5888# 0.039563f
C1050 source.n985 a_n1246_n5888# 0.099432f
C1051 source.t2 a_n1246_n5888# 0.519865f
C1052 source.t3 a_n1246_n5888# 0.519865f
C1053 source.n986 a_n1246_n5888# 4.70485f
C1054 source.n987 a_n1246_n5888# 0.350419f
C1055 source.n988 a_n1246_n5888# 0.036277f
C1056 source.n989 a_n1246_n5888# 0.026315f
C1057 source.n990 a_n1246_n5888# 0.01414f
C1058 source.n991 a_n1246_n5888# 0.033423f
C1059 source.n992 a_n1246_n5888# 0.014972f
C1060 source.n993 a_n1246_n5888# 0.026315f
C1061 source.n994 a_n1246_n5888# 0.01414f
C1062 source.n995 a_n1246_n5888# 0.033423f
C1063 source.n996 a_n1246_n5888# 0.014972f
C1064 source.n997 a_n1246_n5888# 0.026315f
C1065 source.n998 a_n1246_n5888# 0.01414f
C1066 source.n999 a_n1246_n5888# 0.033423f
C1067 source.n1000 a_n1246_n5888# 0.014972f
C1068 source.n1001 a_n1246_n5888# 0.026315f
C1069 source.n1002 a_n1246_n5888# 0.01414f
C1070 source.n1003 a_n1246_n5888# 0.033423f
C1071 source.n1004 a_n1246_n5888# 0.014972f
C1072 source.n1005 a_n1246_n5888# 0.026315f
C1073 source.n1006 a_n1246_n5888# 0.01414f
C1074 source.n1007 a_n1246_n5888# 0.033423f
C1075 source.n1008 a_n1246_n5888# 0.014972f
C1076 source.n1009 a_n1246_n5888# 0.026315f
C1077 source.n1010 a_n1246_n5888# 0.01414f
C1078 source.n1011 a_n1246_n5888# 0.033423f
C1079 source.n1012 a_n1246_n5888# 0.014972f
C1080 source.n1013 a_n1246_n5888# 0.026315f
C1081 source.n1014 a_n1246_n5888# 0.01414f
C1082 source.n1015 a_n1246_n5888# 0.033423f
C1083 source.n1016 a_n1246_n5888# 0.014972f
C1084 source.n1017 a_n1246_n5888# 0.026315f
C1085 source.n1018 a_n1246_n5888# 0.01414f
C1086 source.n1019 a_n1246_n5888# 0.033423f
C1087 source.n1020 a_n1246_n5888# 0.014972f
C1088 source.n1021 a_n1246_n5888# 0.026315f
C1089 source.n1022 a_n1246_n5888# 0.014556f
C1090 source.n1023 a_n1246_n5888# 0.033423f
C1091 source.n1024 a_n1246_n5888# 0.014972f
C1092 source.n1025 a_n1246_n5888# 0.026315f
C1093 source.n1026 a_n1246_n5888# 0.01414f
C1094 source.n1027 a_n1246_n5888# 0.033423f
C1095 source.n1028 a_n1246_n5888# 0.014972f
C1096 source.n1029 a_n1246_n5888# 0.026315f
C1097 source.n1030 a_n1246_n5888# 0.01414f
C1098 source.n1031 a_n1246_n5888# 0.025067f
C1099 source.n1032 a_n1246_n5888# 0.023627f
C1100 source.t1 a_n1246_n5888# 0.058291f
C1101 source.n1033 a_n1246_n5888# 0.32106f
C1102 source.n1034 a_n1246_n5888# 2.8491f
C1103 source.n1035 a_n1246_n5888# 0.01414f
C1104 source.n1036 a_n1246_n5888# 0.014972f
C1105 source.n1037 a_n1246_n5888# 0.033423f
C1106 source.n1038 a_n1246_n5888# 0.033423f
C1107 source.n1039 a_n1246_n5888# 0.014972f
C1108 source.n1040 a_n1246_n5888# 0.01414f
C1109 source.n1041 a_n1246_n5888# 0.026315f
C1110 source.n1042 a_n1246_n5888# 0.026315f
C1111 source.n1043 a_n1246_n5888# 0.01414f
C1112 source.n1044 a_n1246_n5888# 0.014972f
C1113 source.n1045 a_n1246_n5888# 0.033423f
C1114 source.n1046 a_n1246_n5888# 0.033423f
C1115 source.n1047 a_n1246_n5888# 0.014972f
C1116 source.n1048 a_n1246_n5888# 0.01414f
C1117 source.n1049 a_n1246_n5888# 0.026315f
C1118 source.n1050 a_n1246_n5888# 0.026315f
C1119 source.n1051 a_n1246_n5888# 0.01414f
C1120 source.n1052 a_n1246_n5888# 0.01414f
C1121 source.n1053 a_n1246_n5888# 0.014972f
C1122 source.n1054 a_n1246_n5888# 0.033423f
C1123 source.n1055 a_n1246_n5888# 0.033423f
C1124 source.n1056 a_n1246_n5888# 0.033423f
C1125 source.n1057 a_n1246_n5888# 0.014556f
C1126 source.n1058 a_n1246_n5888# 0.01414f
C1127 source.n1059 a_n1246_n5888# 0.026315f
C1128 source.n1060 a_n1246_n5888# 0.026315f
C1129 source.n1061 a_n1246_n5888# 0.01414f
C1130 source.n1062 a_n1246_n5888# 0.014972f
C1131 source.n1063 a_n1246_n5888# 0.033423f
C1132 source.n1064 a_n1246_n5888# 0.033423f
C1133 source.n1065 a_n1246_n5888# 0.014972f
C1134 source.n1066 a_n1246_n5888# 0.01414f
C1135 source.n1067 a_n1246_n5888# 0.026315f
C1136 source.n1068 a_n1246_n5888# 0.026315f
C1137 source.n1069 a_n1246_n5888# 0.01414f
C1138 source.n1070 a_n1246_n5888# 0.014972f
C1139 source.n1071 a_n1246_n5888# 0.033423f
C1140 source.n1072 a_n1246_n5888# 0.033423f
C1141 source.n1073 a_n1246_n5888# 0.014972f
C1142 source.n1074 a_n1246_n5888# 0.01414f
C1143 source.n1075 a_n1246_n5888# 0.026315f
C1144 source.n1076 a_n1246_n5888# 0.026315f
C1145 source.n1077 a_n1246_n5888# 0.01414f
C1146 source.n1078 a_n1246_n5888# 0.014972f
C1147 source.n1079 a_n1246_n5888# 0.033423f
C1148 source.n1080 a_n1246_n5888# 0.033423f
C1149 source.n1081 a_n1246_n5888# 0.014972f
C1150 source.n1082 a_n1246_n5888# 0.01414f
C1151 source.n1083 a_n1246_n5888# 0.026315f
C1152 source.n1084 a_n1246_n5888# 0.026315f
C1153 source.n1085 a_n1246_n5888# 0.01414f
C1154 source.n1086 a_n1246_n5888# 0.014972f
C1155 source.n1087 a_n1246_n5888# 0.033423f
C1156 source.n1088 a_n1246_n5888# 0.033423f
C1157 source.n1089 a_n1246_n5888# 0.014972f
C1158 source.n1090 a_n1246_n5888# 0.01414f
C1159 source.n1091 a_n1246_n5888# 0.026315f
C1160 source.n1092 a_n1246_n5888# 0.026315f
C1161 source.n1093 a_n1246_n5888# 0.01414f
C1162 source.n1094 a_n1246_n5888# 0.014972f
C1163 source.n1095 a_n1246_n5888# 0.033423f
C1164 source.n1096 a_n1246_n5888# 0.033423f
C1165 source.n1097 a_n1246_n5888# 0.033423f
C1166 source.n1098 a_n1246_n5888# 0.014972f
C1167 source.n1099 a_n1246_n5888# 0.01414f
C1168 source.n1100 a_n1246_n5888# 0.026315f
C1169 source.n1101 a_n1246_n5888# 0.026315f
C1170 source.n1102 a_n1246_n5888# 0.01414f
C1171 source.n1103 a_n1246_n5888# 0.014556f
C1172 source.n1104 a_n1246_n5888# 0.014556f
C1173 source.n1105 a_n1246_n5888# 0.033423f
C1174 source.n1106 a_n1246_n5888# 0.033423f
C1175 source.n1107 a_n1246_n5888# 0.014972f
C1176 source.n1108 a_n1246_n5888# 0.01414f
C1177 source.n1109 a_n1246_n5888# 0.026315f
C1178 source.n1110 a_n1246_n5888# 0.026315f
C1179 source.n1111 a_n1246_n5888# 0.01414f
C1180 source.n1112 a_n1246_n5888# 0.014972f
C1181 source.n1113 a_n1246_n5888# 0.033423f
C1182 source.n1114 a_n1246_n5888# 0.033423f
C1183 source.n1115 a_n1246_n5888# 0.014972f
C1184 source.n1116 a_n1246_n5888# 0.01414f
C1185 source.n1117 a_n1246_n5888# 0.026315f
C1186 source.n1118 a_n1246_n5888# 0.026315f
C1187 source.n1119 a_n1246_n5888# 0.01414f
C1188 source.n1120 a_n1246_n5888# 0.014972f
C1189 source.n1121 a_n1246_n5888# 0.033423f
C1190 source.n1122 a_n1246_n5888# 0.071098f
C1191 source.n1123 a_n1246_n5888# 0.014972f
C1192 source.n1124 a_n1246_n5888# 0.01414f
C1193 source.n1125 a_n1246_n5888# 0.057949f
C1194 source.n1126 a_n1246_n5888# 0.039563f
C1195 source.n1127 a_n1246_n5888# 0.242118f
C1196 source.n1128 a_n1246_n5888# 2.80043f
C1197 drain_left.t3 a_n1246_n5888# 0.754936f
C1198 drain_left.t4 a_n1246_n5888# 0.754936f
C1199 drain_left.n0 a_n1246_n5888# 6.95879f
C1200 drain_left.t0 a_n1246_n5888# 0.754936f
C1201 drain_left.t1 a_n1246_n5888# 0.754936f
C1202 drain_left.n1 a_n1246_n5888# 6.95879f
C1203 drain_left.n2 a_n1246_n5888# 3.71768f
C1204 drain_left.t7 a_n1246_n5888# 0.754936f
C1205 drain_left.t6 a_n1246_n5888# 0.754936f
C1206 drain_left.n3 a_n1246_n5888# 6.96104f
C1207 drain_left.t2 a_n1246_n5888# 0.754936f
C1208 drain_left.t5 a_n1246_n5888# 0.754936f
C1209 drain_left.n4 a_n1246_n5888# 6.95754f
C1210 drain_left.n5 a_n1246_n5888# 1.19573f
C1211 plus.n0 a_n1246_n5888# 0.132311f
C1212 plus.t5 a_n1246_n5888# 0.854868f
C1213 plus.t1 a_n1246_n5888# 0.854868f
C1214 plus.t2 a_n1246_n5888# 0.859121f
C1215 plus.n1 a_n1246_n5888# 0.334236f
C1216 plus.n2 a_n1246_n5888# 0.317311f
C1217 plus.n3 a_n1246_n5888# 0.021282f
C1218 plus.n4 a_n1246_n5888# 0.317311f
C1219 plus.t3 a_n1246_n5888# 0.859121f
C1220 plus.n5 a_n1246_n5888# 0.334152f
C1221 plus.n6 a_n1246_n5888# 1.07699f
C1222 plus.n7 a_n1246_n5888# 0.132311f
C1223 plus.t4 a_n1246_n5888# 0.859121f
C1224 plus.t7 a_n1246_n5888# 0.854868f
C1225 plus.t0 a_n1246_n5888# 0.854868f
C1226 plus.t6 a_n1246_n5888# 0.859121f
C1227 plus.n8 a_n1246_n5888# 0.334236f
C1228 plus.n9 a_n1246_n5888# 0.317311f
C1229 plus.n10 a_n1246_n5888# 0.021282f
C1230 plus.n11 a_n1246_n5888# 0.317311f
C1231 plus.n12 a_n1246_n5888# 0.334152f
C1232 plus.n13 a_n1246_n5888# 2.1519f
.ends

