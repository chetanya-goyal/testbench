* NGSPICE file created from diffpair654.ext - technology: sky130A

.subckt diffpair654 minus drain_right drain_left source plus
X0 a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.2
X1 source.t19 plus.t0 drain_left.t7 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X2 drain_right.t9 minus.t0 source.t0 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X3 source.t18 plus.t1 drain_left.t6 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X4 drain_right.t8 minus.t1 source.t5 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X5 drain_right.t7 minus.t2 source.t3 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X6 source.t9 minus.t3 drain_right.t6 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X7 source.t2 minus.t4 drain_right.t5 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X8 source.t6 minus.t5 drain_right.t4 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X9 drain_left.t1 plus.t2 source.t17 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X10 drain_right.t3 minus.t6 source.t8 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X11 drain_right.t2 minus.t7 source.t7 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X12 drain_right.t1 minus.t8 source.t1 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X13 a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X14 a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X15 drain_left.t0 plus.t3 source.t16 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X16 source.t15 plus.t4 drain_left.t3 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X17 source.t14 plus.t5 drain_left.t2 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X18 source.t4 minus.t9 drain_right.t0 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X19 a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X20 drain_left.t5 plus.t6 source.t13 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X21 drain_left.t4 plus.t7 source.t12 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X22 drain_left.t9 plus.t8 source.t11 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X23 drain_left.t8 plus.t9 source.t10 a_n1352_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
R0 plus.n2 plus.t2 3214.43
R1 plus.n8 plus.t3 3214.43
R2 plus.n12 plus.t8 3214.43
R3 plus.n18 plus.t6 3214.43
R4 plus.n1 plus.t1 3169.15
R5 plus.n5 plus.t7 3169.15
R6 plus.n7 plus.t4 3169.15
R7 plus.n11 plus.t0 3169.15
R8 plus.n15 plus.t9 3169.15
R9 plus.n17 plus.t5 3169.15
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 40.8975
R19 plus.n7 plus.n6 40.8975
R20 plus.n17 plus.n16 40.8975
R21 plus.n14 plus.n11 40.8975
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 32.9971
R27 plus.n2 plus.n1 32.1338
R28 plus.n8 plus.n7 32.1338
R29 plus.n18 plus.n17 32.1338
R30 plus.n12 plus.n11 32.1338
R31 plus plus.n9 17.0175
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n134 drain_left.n0 289.615
R37 drain_left.n277 drain_left.n143 289.615
R38 drain_left.n44 drain_left.n43 185
R39 drain_left.n49 drain_left.n48 185
R40 drain_left.n51 drain_left.n50 185
R41 drain_left.n40 drain_left.n39 185
R42 drain_left.n57 drain_left.n56 185
R43 drain_left.n59 drain_left.n58 185
R44 drain_left.n36 drain_left.n35 185
R45 drain_left.n66 drain_left.n65 185
R46 drain_left.n67 drain_left.n34 185
R47 drain_left.n69 drain_left.n68 185
R48 drain_left.n32 drain_left.n31 185
R49 drain_left.n75 drain_left.n74 185
R50 drain_left.n77 drain_left.n76 185
R51 drain_left.n28 drain_left.n27 185
R52 drain_left.n83 drain_left.n82 185
R53 drain_left.n85 drain_left.n84 185
R54 drain_left.n24 drain_left.n23 185
R55 drain_left.n91 drain_left.n90 185
R56 drain_left.n93 drain_left.n92 185
R57 drain_left.n20 drain_left.n19 185
R58 drain_left.n99 drain_left.n98 185
R59 drain_left.n101 drain_left.n100 185
R60 drain_left.n16 drain_left.n15 185
R61 drain_left.n107 drain_left.n106 185
R62 drain_left.n110 drain_left.n109 185
R63 drain_left.n108 drain_left.n12 185
R64 drain_left.n115 drain_left.n11 185
R65 drain_left.n117 drain_left.n116 185
R66 drain_left.n119 drain_left.n118 185
R67 drain_left.n8 drain_left.n7 185
R68 drain_left.n125 drain_left.n124 185
R69 drain_left.n127 drain_left.n126 185
R70 drain_left.n4 drain_left.n3 185
R71 drain_left.n133 drain_left.n132 185
R72 drain_left.n135 drain_left.n134 185
R73 drain_left.n278 drain_left.n277 185
R74 drain_left.n276 drain_left.n275 185
R75 drain_left.n147 drain_left.n146 185
R76 drain_left.n270 drain_left.n269 185
R77 drain_left.n268 drain_left.n267 185
R78 drain_left.n151 drain_left.n150 185
R79 drain_left.n262 drain_left.n261 185
R80 drain_left.n260 drain_left.n259 185
R81 drain_left.n258 drain_left.n154 185
R82 drain_left.n158 drain_left.n155 185
R83 drain_left.n253 drain_left.n252 185
R84 drain_left.n251 drain_left.n250 185
R85 drain_left.n160 drain_left.n159 185
R86 drain_left.n245 drain_left.n244 185
R87 drain_left.n243 drain_left.n242 185
R88 drain_left.n164 drain_left.n163 185
R89 drain_left.n237 drain_left.n236 185
R90 drain_left.n235 drain_left.n234 185
R91 drain_left.n168 drain_left.n167 185
R92 drain_left.n229 drain_left.n228 185
R93 drain_left.n227 drain_left.n226 185
R94 drain_left.n172 drain_left.n171 185
R95 drain_left.n221 drain_left.n220 185
R96 drain_left.n219 drain_left.n218 185
R97 drain_left.n176 drain_left.n175 185
R98 drain_left.n213 drain_left.n212 185
R99 drain_left.n211 drain_left.n178 185
R100 drain_left.n210 drain_left.n209 185
R101 drain_left.n181 drain_left.n179 185
R102 drain_left.n204 drain_left.n203 185
R103 drain_left.n202 drain_left.n201 185
R104 drain_left.n185 drain_left.n184 185
R105 drain_left.n196 drain_left.n195 185
R106 drain_left.n194 drain_left.n193 185
R107 drain_left.n189 drain_left.n188 185
R108 drain_left.n45 drain_left.t5 149.524
R109 drain_left.n190 drain_left.t1 149.524
R110 drain_left.n49 drain_left.n43 104.615
R111 drain_left.n50 drain_left.n49 104.615
R112 drain_left.n50 drain_left.n39 104.615
R113 drain_left.n57 drain_left.n39 104.615
R114 drain_left.n58 drain_left.n57 104.615
R115 drain_left.n58 drain_left.n35 104.615
R116 drain_left.n66 drain_left.n35 104.615
R117 drain_left.n67 drain_left.n66 104.615
R118 drain_left.n68 drain_left.n67 104.615
R119 drain_left.n68 drain_left.n31 104.615
R120 drain_left.n75 drain_left.n31 104.615
R121 drain_left.n76 drain_left.n75 104.615
R122 drain_left.n76 drain_left.n27 104.615
R123 drain_left.n83 drain_left.n27 104.615
R124 drain_left.n84 drain_left.n83 104.615
R125 drain_left.n84 drain_left.n23 104.615
R126 drain_left.n91 drain_left.n23 104.615
R127 drain_left.n92 drain_left.n91 104.615
R128 drain_left.n92 drain_left.n19 104.615
R129 drain_left.n99 drain_left.n19 104.615
R130 drain_left.n100 drain_left.n99 104.615
R131 drain_left.n100 drain_left.n15 104.615
R132 drain_left.n107 drain_left.n15 104.615
R133 drain_left.n109 drain_left.n107 104.615
R134 drain_left.n109 drain_left.n108 104.615
R135 drain_left.n108 drain_left.n11 104.615
R136 drain_left.n117 drain_left.n11 104.615
R137 drain_left.n118 drain_left.n117 104.615
R138 drain_left.n118 drain_left.n7 104.615
R139 drain_left.n125 drain_left.n7 104.615
R140 drain_left.n126 drain_left.n125 104.615
R141 drain_left.n126 drain_left.n3 104.615
R142 drain_left.n133 drain_left.n3 104.615
R143 drain_left.n134 drain_left.n133 104.615
R144 drain_left.n277 drain_left.n276 104.615
R145 drain_left.n276 drain_left.n146 104.615
R146 drain_left.n269 drain_left.n146 104.615
R147 drain_left.n269 drain_left.n268 104.615
R148 drain_left.n268 drain_left.n150 104.615
R149 drain_left.n261 drain_left.n150 104.615
R150 drain_left.n261 drain_left.n260 104.615
R151 drain_left.n260 drain_left.n154 104.615
R152 drain_left.n158 drain_left.n154 104.615
R153 drain_left.n252 drain_left.n158 104.615
R154 drain_left.n252 drain_left.n251 104.615
R155 drain_left.n251 drain_left.n159 104.615
R156 drain_left.n244 drain_left.n159 104.615
R157 drain_left.n244 drain_left.n243 104.615
R158 drain_left.n243 drain_left.n163 104.615
R159 drain_left.n236 drain_left.n163 104.615
R160 drain_left.n236 drain_left.n235 104.615
R161 drain_left.n235 drain_left.n167 104.615
R162 drain_left.n228 drain_left.n167 104.615
R163 drain_left.n228 drain_left.n227 104.615
R164 drain_left.n227 drain_left.n171 104.615
R165 drain_left.n220 drain_left.n171 104.615
R166 drain_left.n220 drain_left.n219 104.615
R167 drain_left.n219 drain_left.n175 104.615
R168 drain_left.n212 drain_left.n175 104.615
R169 drain_left.n212 drain_left.n211 104.615
R170 drain_left.n211 drain_left.n210 104.615
R171 drain_left.n210 drain_left.n179 104.615
R172 drain_left.n203 drain_left.n179 104.615
R173 drain_left.n203 drain_left.n202 104.615
R174 drain_left.n202 drain_left.n184 104.615
R175 drain_left.n195 drain_left.n184 104.615
R176 drain_left.n195 drain_left.n194 104.615
R177 drain_left.n194 drain_left.n188 104.615
R178 drain_left.n142 drain_left.n141 59.0028
R179 drain_left.n140 drain_left.n139 58.7154
R180 drain_left.n283 drain_left.n282 58.7154
R181 drain_left.n285 drain_left.n284 58.7153
R182 drain_left.t5 drain_left.n43 52.3082
R183 drain_left.t1 drain_left.n188 52.3082
R184 drain_left.n140 drain_left.n138 47.7695
R185 drain_left.n283 drain_left.n281 47.7695
R186 drain_left drain_left.n142 39.1574
R187 drain_left.n69 drain_left.n34 13.1884
R188 drain_left.n116 drain_left.n115 13.1884
R189 drain_left.n259 drain_left.n258 13.1884
R190 drain_left.n213 drain_left.n178 13.1884
R191 drain_left.n65 drain_left.n64 12.8005
R192 drain_left.n70 drain_left.n32 12.8005
R193 drain_left.n114 drain_left.n12 12.8005
R194 drain_left.n119 drain_left.n10 12.8005
R195 drain_left.n262 drain_left.n153 12.8005
R196 drain_left.n257 drain_left.n155 12.8005
R197 drain_left.n214 drain_left.n176 12.8005
R198 drain_left.n209 drain_left.n180 12.8005
R199 drain_left.n63 drain_left.n36 12.0247
R200 drain_left.n74 drain_left.n73 12.0247
R201 drain_left.n111 drain_left.n110 12.0247
R202 drain_left.n120 drain_left.n8 12.0247
R203 drain_left.n263 drain_left.n151 12.0247
R204 drain_left.n254 drain_left.n253 12.0247
R205 drain_left.n218 drain_left.n217 12.0247
R206 drain_left.n208 drain_left.n181 12.0247
R207 drain_left.n60 drain_left.n59 11.249
R208 drain_left.n77 drain_left.n30 11.249
R209 drain_left.n106 drain_left.n14 11.249
R210 drain_left.n124 drain_left.n123 11.249
R211 drain_left.n267 drain_left.n266 11.249
R212 drain_left.n250 drain_left.n157 11.249
R213 drain_left.n221 drain_left.n174 11.249
R214 drain_left.n205 drain_left.n204 11.249
R215 drain_left.n56 drain_left.n38 10.4732
R216 drain_left.n78 drain_left.n28 10.4732
R217 drain_left.n105 drain_left.n16 10.4732
R218 drain_left.n127 drain_left.n6 10.4732
R219 drain_left.n270 drain_left.n149 10.4732
R220 drain_left.n249 drain_left.n160 10.4732
R221 drain_left.n222 drain_left.n172 10.4732
R222 drain_left.n201 drain_left.n183 10.4732
R223 drain_left.n45 drain_left.n44 10.2747
R224 drain_left.n190 drain_left.n189 10.2747
R225 drain_left.n55 drain_left.n40 9.69747
R226 drain_left.n82 drain_left.n81 9.69747
R227 drain_left.n102 drain_left.n101 9.69747
R228 drain_left.n128 drain_left.n4 9.69747
R229 drain_left.n271 drain_left.n147 9.69747
R230 drain_left.n246 drain_left.n245 9.69747
R231 drain_left.n226 drain_left.n225 9.69747
R232 drain_left.n200 drain_left.n185 9.69747
R233 drain_left.n138 drain_left.n137 9.45567
R234 drain_left.n281 drain_left.n280 9.45567
R235 drain_left.n2 drain_left.n1 9.3005
R236 drain_left.n131 drain_left.n130 9.3005
R237 drain_left.n129 drain_left.n128 9.3005
R238 drain_left.n6 drain_left.n5 9.3005
R239 drain_left.n123 drain_left.n122 9.3005
R240 drain_left.n121 drain_left.n120 9.3005
R241 drain_left.n10 drain_left.n9 9.3005
R242 drain_left.n89 drain_left.n88 9.3005
R243 drain_left.n87 drain_left.n86 9.3005
R244 drain_left.n26 drain_left.n25 9.3005
R245 drain_left.n81 drain_left.n80 9.3005
R246 drain_left.n79 drain_left.n78 9.3005
R247 drain_left.n30 drain_left.n29 9.3005
R248 drain_left.n73 drain_left.n72 9.3005
R249 drain_left.n71 drain_left.n70 9.3005
R250 drain_left.n47 drain_left.n46 9.3005
R251 drain_left.n42 drain_left.n41 9.3005
R252 drain_left.n53 drain_left.n52 9.3005
R253 drain_left.n55 drain_left.n54 9.3005
R254 drain_left.n38 drain_left.n37 9.3005
R255 drain_left.n61 drain_left.n60 9.3005
R256 drain_left.n63 drain_left.n62 9.3005
R257 drain_left.n64 drain_left.n33 9.3005
R258 drain_left.n22 drain_left.n21 9.3005
R259 drain_left.n95 drain_left.n94 9.3005
R260 drain_left.n97 drain_left.n96 9.3005
R261 drain_left.n18 drain_left.n17 9.3005
R262 drain_left.n103 drain_left.n102 9.3005
R263 drain_left.n105 drain_left.n104 9.3005
R264 drain_left.n14 drain_left.n13 9.3005
R265 drain_left.n112 drain_left.n111 9.3005
R266 drain_left.n114 drain_left.n113 9.3005
R267 drain_left.n137 drain_left.n136 9.3005
R268 drain_left.n192 drain_left.n191 9.3005
R269 drain_left.n187 drain_left.n186 9.3005
R270 drain_left.n198 drain_left.n197 9.3005
R271 drain_left.n200 drain_left.n199 9.3005
R272 drain_left.n183 drain_left.n182 9.3005
R273 drain_left.n206 drain_left.n205 9.3005
R274 drain_left.n208 drain_left.n207 9.3005
R275 drain_left.n180 drain_left.n177 9.3005
R276 drain_left.n239 drain_left.n238 9.3005
R277 drain_left.n241 drain_left.n240 9.3005
R278 drain_left.n162 drain_left.n161 9.3005
R279 drain_left.n247 drain_left.n246 9.3005
R280 drain_left.n249 drain_left.n248 9.3005
R281 drain_left.n157 drain_left.n156 9.3005
R282 drain_left.n255 drain_left.n254 9.3005
R283 drain_left.n257 drain_left.n256 9.3005
R284 drain_left.n280 drain_left.n279 9.3005
R285 drain_left.n145 drain_left.n144 9.3005
R286 drain_left.n274 drain_left.n273 9.3005
R287 drain_left.n272 drain_left.n271 9.3005
R288 drain_left.n149 drain_left.n148 9.3005
R289 drain_left.n266 drain_left.n265 9.3005
R290 drain_left.n264 drain_left.n263 9.3005
R291 drain_left.n153 drain_left.n152 9.3005
R292 drain_left.n166 drain_left.n165 9.3005
R293 drain_left.n233 drain_left.n232 9.3005
R294 drain_left.n231 drain_left.n230 9.3005
R295 drain_left.n170 drain_left.n169 9.3005
R296 drain_left.n225 drain_left.n224 9.3005
R297 drain_left.n223 drain_left.n222 9.3005
R298 drain_left.n174 drain_left.n173 9.3005
R299 drain_left.n217 drain_left.n216 9.3005
R300 drain_left.n215 drain_left.n214 9.3005
R301 drain_left.n52 drain_left.n51 8.92171
R302 drain_left.n85 drain_left.n26 8.92171
R303 drain_left.n98 drain_left.n18 8.92171
R304 drain_left.n132 drain_left.n131 8.92171
R305 drain_left.n275 drain_left.n274 8.92171
R306 drain_left.n242 drain_left.n162 8.92171
R307 drain_left.n229 drain_left.n170 8.92171
R308 drain_left.n197 drain_left.n196 8.92171
R309 drain_left.n48 drain_left.n42 8.14595
R310 drain_left.n86 drain_left.n24 8.14595
R311 drain_left.n97 drain_left.n20 8.14595
R312 drain_left.n135 drain_left.n2 8.14595
R313 drain_left.n278 drain_left.n145 8.14595
R314 drain_left.n241 drain_left.n164 8.14595
R315 drain_left.n230 drain_left.n168 8.14595
R316 drain_left.n193 drain_left.n187 8.14595
R317 drain_left.n47 drain_left.n44 7.3702
R318 drain_left.n90 drain_left.n89 7.3702
R319 drain_left.n94 drain_left.n93 7.3702
R320 drain_left.n136 drain_left.n0 7.3702
R321 drain_left.n279 drain_left.n143 7.3702
R322 drain_left.n238 drain_left.n237 7.3702
R323 drain_left.n234 drain_left.n233 7.3702
R324 drain_left.n192 drain_left.n189 7.3702
R325 drain_left.n90 drain_left.n22 6.59444
R326 drain_left.n93 drain_left.n22 6.59444
R327 drain_left.n138 drain_left.n0 6.59444
R328 drain_left.n281 drain_left.n143 6.59444
R329 drain_left.n237 drain_left.n166 6.59444
R330 drain_left.n234 drain_left.n166 6.59444
R331 drain_left drain_left.n285 6.11011
R332 drain_left.n48 drain_left.n47 5.81868
R333 drain_left.n89 drain_left.n24 5.81868
R334 drain_left.n94 drain_left.n20 5.81868
R335 drain_left.n136 drain_left.n135 5.81868
R336 drain_left.n279 drain_left.n278 5.81868
R337 drain_left.n238 drain_left.n164 5.81868
R338 drain_left.n233 drain_left.n168 5.81868
R339 drain_left.n193 drain_left.n192 5.81868
R340 drain_left.n51 drain_left.n42 5.04292
R341 drain_left.n86 drain_left.n85 5.04292
R342 drain_left.n98 drain_left.n97 5.04292
R343 drain_left.n132 drain_left.n2 5.04292
R344 drain_left.n275 drain_left.n145 5.04292
R345 drain_left.n242 drain_left.n241 5.04292
R346 drain_left.n230 drain_left.n229 5.04292
R347 drain_left.n196 drain_left.n187 5.04292
R348 drain_left.n52 drain_left.n40 4.26717
R349 drain_left.n82 drain_left.n26 4.26717
R350 drain_left.n101 drain_left.n18 4.26717
R351 drain_left.n131 drain_left.n4 4.26717
R352 drain_left.n274 drain_left.n147 4.26717
R353 drain_left.n245 drain_left.n162 4.26717
R354 drain_left.n226 drain_left.n170 4.26717
R355 drain_left.n197 drain_left.n185 4.26717
R356 drain_left.n56 drain_left.n55 3.49141
R357 drain_left.n81 drain_left.n28 3.49141
R358 drain_left.n102 drain_left.n16 3.49141
R359 drain_left.n128 drain_left.n127 3.49141
R360 drain_left.n271 drain_left.n270 3.49141
R361 drain_left.n246 drain_left.n160 3.49141
R362 drain_left.n225 drain_left.n172 3.49141
R363 drain_left.n201 drain_left.n200 3.49141
R364 drain_left.n191 drain_left.n190 2.84303
R365 drain_left.n46 drain_left.n45 2.84303
R366 drain_left.n59 drain_left.n38 2.71565
R367 drain_left.n78 drain_left.n77 2.71565
R368 drain_left.n106 drain_left.n105 2.71565
R369 drain_left.n124 drain_left.n6 2.71565
R370 drain_left.n267 drain_left.n149 2.71565
R371 drain_left.n250 drain_left.n249 2.71565
R372 drain_left.n222 drain_left.n221 2.71565
R373 drain_left.n204 drain_left.n183 2.71565
R374 drain_left.n60 drain_left.n36 1.93989
R375 drain_left.n74 drain_left.n30 1.93989
R376 drain_left.n110 drain_left.n14 1.93989
R377 drain_left.n123 drain_left.n8 1.93989
R378 drain_left.n266 drain_left.n151 1.93989
R379 drain_left.n253 drain_left.n157 1.93989
R380 drain_left.n218 drain_left.n174 1.93989
R381 drain_left.n205 drain_left.n181 1.93989
R382 drain_left.n65 drain_left.n63 1.16414
R383 drain_left.n73 drain_left.n32 1.16414
R384 drain_left.n111 drain_left.n12 1.16414
R385 drain_left.n120 drain_left.n119 1.16414
R386 drain_left.n263 drain_left.n262 1.16414
R387 drain_left.n254 drain_left.n155 1.16414
R388 drain_left.n217 drain_left.n176 1.16414
R389 drain_left.n209 drain_left.n208 1.16414
R390 drain_left.n141 drain_left.t7 0.7925
R391 drain_left.n141 drain_left.t9 0.7925
R392 drain_left.n139 drain_left.t2 0.7925
R393 drain_left.n139 drain_left.t8 0.7925
R394 drain_left.n284 drain_left.t3 0.7925
R395 drain_left.n284 drain_left.t0 0.7925
R396 drain_left.n282 drain_left.t6 0.7925
R397 drain_left.n282 drain_left.t4 0.7925
R398 drain_left.n285 drain_left.n283 0.457397
R399 drain_left.n64 drain_left.n34 0.388379
R400 drain_left.n70 drain_left.n69 0.388379
R401 drain_left.n115 drain_left.n114 0.388379
R402 drain_left.n116 drain_left.n10 0.388379
R403 drain_left.n259 drain_left.n153 0.388379
R404 drain_left.n258 drain_left.n257 0.388379
R405 drain_left.n214 drain_left.n213 0.388379
R406 drain_left.n180 drain_left.n178 0.388379
R407 drain_left.n46 drain_left.n41 0.155672
R408 drain_left.n53 drain_left.n41 0.155672
R409 drain_left.n54 drain_left.n53 0.155672
R410 drain_left.n54 drain_left.n37 0.155672
R411 drain_left.n61 drain_left.n37 0.155672
R412 drain_left.n62 drain_left.n61 0.155672
R413 drain_left.n62 drain_left.n33 0.155672
R414 drain_left.n71 drain_left.n33 0.155672
R415 drain_left.n72 drain_left.n71 0.155672
R416 drain_left.n72 drain_left.n29 0.155672
R417 drain_left.n79 drain_left.n29 0.155672
R418 drain_left.n80 drain_left.n79 0.155672
R419 drain_left.n80 drain_left.n25 0.155672
R420 drain_left.n87 drain_left.n25 0.155672
R421 drain_left.n88 drain_left.n87 0.155672
R422 drain_left.n88 drain_left.n21 0.155672
R423 drain_left.n95 drain_left.n21 0.155672
R424 drain_left.n96 drain_left.n95 0.155672
R425 drain_left.n96 drain_left.n17 0.155672
R426 drain_left.n103 drain_left.n17 0.155672
R427 drain_left.n104 drain_left.n103 0.155672
R428 drain_left.n104 drain_left.n13 0.155672
R429 drain_left.n112 drain_left.n13 0.155672
R430 drain_left.n113 drain_left.n112 0.155672
R431 drain_left.n113 drain_left.n9 0.155672
R432 drain_left.n121 drain_left.n9 0.155672
R433 drain_left.n122 drain_left.n121 0.155672
R434 drain_left.n122 drain_left.n5 0.155672
R435 drain_left.n129 drain_left.n5 0.155672
R436 drain_left.n130 drain_left.n129 0.155672
R437 drain_left.n130 drain_left.n1 0.155672
R438 drain_left.n137 drain_left.n1 0.155672
R439 drain_left.n280 drain_left.n144 0.155672
R440 drain_left.n273 drain_left.n144 0.155672
R441 drain_left.n273 drain_left.n272 0.155672
R442 drain_left.n272 drain_left.n148 0.155672
R443 drain_left.n265 drain_left.n148 0.155672
R444 drain_left.n265 drain_left.n264 0.155672
R445 drain_left.n264 drain_left.n152 0.155672
R446 drain_left.n256 drain_left.n152 0.155672
R447 drain_left.n256 drain_left.n255 0.155672
R448 drain_left.n255 drain_left.n156 0.155672
R449 drain_left.n248 drain_left.n156 0.155672
R450 drain_left.n248 drain_left.n247 0.155672
R451 drain_left.n247 drain_left.n161 0.155672
R452 drain_left.n240 drain_left.n161 0.155672
R453 drain_left.n240 drain_left.n239 0.155672
R454 drain_left.n239 drain_left.n165 0.155672
R455 drain_left.n232 drain_left.n165 0.155672
R456 drain_left.n232 drain_left.n231 0.155672
R457 drain_left.n231 drain_left.n169 0.155672
R458 drain_left.n224 drain_left.n169 0.155672
R459 drain_left.n224 drain_left.n223 0.155672
R460 drain_left.n223 drain_left.n173 0.155672
R461 drain_left.n216 drain_left.n173 0.155672
R462 drain_left.n216 drain_left.n215 0.155672
R463 drain_left.n215 drain_left.n177 0.155672
R464 drain_left.n207 drain_left.n177 0.155672
R465 drain_left.n207 drain_left.n206 0.155672
R466 drain_left.n206 drain_left.n182 0.155672
R467 drain_left.n199 drain_left.n182 0.155672
R468 drain_left.n199 drain_left.n198 0.155672
R469 drain_left.n198 drain_left.n186 0.155672
R470 drain_left.n191 drain_left.n186 0.155672
R471 drain_left.n142 drain_left.n140 0.0593781
R472 source.n570 source.n436 289.615
R473 source.n426 source.n292 289.615
R474 source.n134 source.n0 289.615
R475 source.n278 source.n144 289.615
R476 source.n480 source.n479 185
R477 source.n485 source.n484 185
R478 source.n487 source.n486 185
R479 source.n476 source.n475 185
R480 source.n493 source.n492 185
R481 source.n495 source.n494 185
R482 source.n472 source.n471 185
R483 source.n502 source.n501 185
R484 source.n503 source.n470 185
R485 source.n505 source.n504 185
R486 source.n468 source.n467 185
R487 source.n511 source.n510 185
R488 source.n513 source.n512 185
R489 source.n464 source.n463 185
R490 source.n519 source.n518 185
R491 source.n521 source.n520 185
R492 source.n460 source.n459 185
R493 source.n527 source.n526 185
R494 source.n529 source.n528 185
R495 source.n456 source.n455 185
R496 source.n535 source.n534 185
R497 source.n537 source.n536 185
R498 source.n452 source.n451 185
R499 source.n543 source.n542 185
R500 source.n546 source.n545 185
R501 source.n544 source.n448 185
R502 source.n551 source.n447 185
R503 source.n553 source.n552 185
R504 source.n555 source.n554 185
R505 source.n444 source.n443 185
R506 source.n561 source.n560 185
R507 source.n563 source.n562 185
R508 source.n440 source.n439 185
R509 source.n569 source.n568 185
R510 source.n571 source.n570 185
R511 source.n336 source.n335 185
R512 source.n341 source.n340 185
R513 source.n343 source.n342 185
R514 source.n332 source.n331 185
R515 source.n349 source.n348 185
R516 source.n351 source.n350 185
R517 source.n328 source.n327 185
R518 source.n358 source.n357 185
R519 source.n359 source.n326 185
R520 source.n361 source.n360 185
R521 source.n324 source.n323 185
R522 source.n367 source.n366 185
R523 source.n369 source.n368 185
R524 source.n320 source.n319 185
R525 source.n375 source.n374 185
R526 source.n377 source.n376 185
R527 source.n316 source.n315 185
R528 source.n383 source.n382 185
R529 source.n385 source.n384 185
R530 source.n312 source.n311 185
R531 source.n391 source.n390 185
R532 source.n393 source.n392 185
R533 source.n308 source.n307 185
R534 source.n399 source.n398 185
R535 source.n402 source.n401 185
R536 source.n400 source.n304 185
R537 source.n407 source.n303 185
R538 source.n409 source.n408 185
R539 source.n411 source.n410 185
R540 source.n300 source.n299 185
R541 source.n417 source.n416 185
R542 source.n419 source.n418 185
R543 source.n296 source.n295 185
R544 source.n425 source.n424 185
R545 source.n427 source.n426 185
R546 source.n135 source.n134 185
R547 source.n133 source.n132 185
R548 source.n4 source.n3 185
R549 source.n127 source.n126 185
R550 source.n125 source.n124 185
R551 source.n8 source.n7 185
R552 source.n119 source.n118 185
R553 source.n117 source.n116 185
R554 source.n115 source.n11 185
R555 source.n15 source.n12 185
R556 source.n110 source.n109 185
R557 source.n108 source.n107 185
R558 source.n17 source.n16 185
R559 source.n102 source.n101 185
R560 source.n100 source.n99 185
R561 source.n21 source.n20 185
R562 source.n94 source.n93 185
R563 source.n92 source.n91 185
R564 source.n25 source.n24 185
R565 source.n86 source.n85 185
R566 source.n84 source.n83 185
R567 source.n29 source.n28 185
R568 source.n78 source.n77 185
R569 source.n76 source.n75 185
R570 source.n33 source.n32 185
R571 source.n70 source.n69 185
R572 source.n68 source.n35 185
R573 source.n67 source.n66 185
R574 source.n38 source.n36 185
R575 source.n61 source.n60 185
R576 source.n59 source.n58 185
R577 source.n42 source.n41 185
R578 source.n53 source.n52 185
R579 source.n51 source.n50 185
R580 source.n46 source.n45 185
R581 source.n279 source.n278 185
R582 source.n277 source.n276 185
R583 source.n148 source.n147 185
R584 source.n271 source.n270 185
R585 source.n269 source.n268 185
R586 source.n152 source.n151 185
R587 source.n263 source.n262 185
R588 source.n261 source.n260 185
R589 source.n259 source.n155 185
R590 source.n159 source.n156 185
R591 source.n254 source.n253 185
R592 source.n252 source.n251 185
R593 source.n161 source.n160 185
R594 source.n246 source.n245 185
R595 source.n244 source.n243 185
R596 source.n165 source.n164 185
R597 source.n238 source.n237 185
R598 source.n236 source.n235 185
R599 source.n169 source.n168 185
R600 source.n230 source.n229 185
R601 source.n228 source.n227 185
R602 source.n173 source.n172 185
R603 source.n222 source.n221 185
R604 source.n220 source.n219 185
R605 source.n177 source.n176 185
R606 source.n214 source.n213 185
R607 source.n212 source.n179 185
R608 source.n211 source.n210 185
R609 source.n182 source.n180 185
R610 source.n205 source.n204 185
R611 source.n203 source.n202 185
R612 source.n186 source.n185 185
R613 source.n197 source.n196 185
R614 source.n195 source.n194 185
R615 source.n190 source.n189 185
R616 source.n481 source.t8 149.524
R617 source.n337 source.t11 149.524
R618 source.n47 source.t16 149.524
R619 source.n191 source.t7 149.524
R620 source.n485 source.n479 104.615
R621 source.n486 source.n485 104.615
R622 source.n486 source.n475 104.615
R623 source.n493 source.n475 104.615
R624 source.n494 source.n493 104.615
R625 source.n494 source.n471 104.615
R626 source.n502 source.n471 104.615
R627 source.n503 source.n502 104.615
R628 source.n504 source.n503 104.615
R629 source.n504 source.n467 104.615
R630 source.n511 source.n467 104.615
R631 source.n512 source.n511 104.615
R632 source.n512 source.n463 104.615
R633 source.n519 source.n463 104.615
R634 source.n520 source.n519 104.615
R635 source.n520 source.n459 104.615
R636 source.n527 source.n459 104.615
R637 source.n528 source.n527 104.615
R638 source.n528 source.n455 104.615
R639 source.n535 source.n455 104.615
R640 source.n536 source.n535 104.615
R641 source.n536 source.n451 104.615
R642 source.n543 source.n451 104.615
R643 source.n545 source.n543 104.615
R644 source.n545 source.n544 104.615
R645 source.n544 source.n447 104.615
R646 source.n553 source.n447 104.615
R647 source.n554 source.n553 104.615
R648 source.n554 source.n443 104.615
R649 source.n561 source.n443 104.615
R650 source.n562 source.n561 104.615
R651 source.n562 source.n439 104.615
R652 source.n569 source.n439 104.615
R653 source.n570 source.n569 104.615
R654 source.n341 source.n335 104.615
R655 source.n342 source.n341 104.615
R656 source.n342 source.n331 104.615
R657 source.n349 source.n331 104.615
R658 source.n350 source.n349 104.615
R659 source.n350 source.n327 104.615
R660 source.n358 source.n327 104.615
R661 source.n359 source.n358 104.615
R662 source.n360 source.n359 104.615
R663 source.n360 source.n323 104.615
R664 source.n367 source.n323 104.615
R665 source.n368 source.n367 104.615
R666 source.n368 source.n319 104.615
R667 source.n375 source.n319 104.615
R668 source.n376 source.n375 104.615
R669 source.n376 source.n315 104.615
R670 source.n383 source.n315 104.615
R671 source.n384 source.n383 104.615
R672 source.n384 source.n311 104.615
R673 source.n391 source.n311 104.615
R674 source.n392 source.n391 104.615
R675 source.n392 source.n307 104.615
R676 source.n399 source.n307 104.615
R677 source.n401 source.n399 104.615
R678 source.n401 source.n400 104.615
R679 source.n400 source.n303 104.615
R680 source.n409 source.n303 104.615
R681 source.n410 source.n409 104.615
R682 source.n410 source.n299 104.615
R683 source.n417 source.n299 104.615
R684 source.n418 source.n417 104.615
R685 source.n418 source.n295 104.615
R686 source.n425 source.n295 104.615
R687 source.n426 source.n425 104.615
R688 source.n134 source.n133 104.615
R689 source.n133 source.n3 104.615
R690 source.n126 source.n3 104.615
R691 source.n126 source.n125 104.615
R692 source.n125 source.n7 104.615
R693 source.n118 source.n7 104.615
R694 source.n118 source.n117 104.615
R695 source.n117 source.n11 104.615
R696 source.n15 source.n11 104.615
R697 source.n109 source.n15 104.615
R698 source.n109 source.n108 104.615
R699 source.n108 source.n16 104.615
R700 source.n101 source.n16 104.615
R701 source.n101 source.n100 104.615
R702 source.n100 source.n20 104.615
R703 source.n93 source.n20 104.615
R704 source.n93 source.n92 104.615
R705 source.n92 source.n24 104.615
R706 source.n85 source.n24 104.615
R707 source.n85 source.n84 104.615
R708 source.n84 source.n28 104.615
R709 source.n77 source.n28 104.615
R710 source.n77 source.n76 104.615
R711 source.n76 source.n32 104.615
R712 source.n69 source.n32 104.615
R713 source.n69 source.n68 104.615
R714 source.n68 source.n67 104.615
R715 source.n67 source.n36 104.615
R716 source.n60 source.n36 104.615
R717 source.n60 source.n59 104.615
R718 source.n59 source.n41 104.615
R719 source.n52 source.n41 104.615
R720 source.n52 source.n51 104.615
R721 source.n51 source.n45 104.615
R722 source.n278 source.n277 104.615
R723 source.n277 source.n147 104.615
R724 source.n270 source.n147 104.615
R725 source.n270 source.n269 104.615
R726 source.n269 source.n151 104.615
R727 source.n262 source.n151 104.615
R728 source.n262 source.n261 104.615
R729 source.n261 source.n155 104.615
R730 source.n159 source.n155 104.615
R731 source.n253 source.n159 104.615
R732 source.n253 source.n252 104.615
R733 source.n252 source.n160 104.615
R734 source.n245 source.n160 104.615
R735 source.n245 source.n244 104.615
R736 source.n244 source.n164 104.615
R737 source.n237 source.n164 104.615
R738 source.n237 source.n236 104.615
R739 source.n236 source.n168 104.615
R740 source.n229 source.n168 104.615
R741 source.n229 source.n228 104.615
R742 source.n228 source.n172 104.615
R743 source.n221 source.n172 104.615
R744 source.n221 source.n220 104.615
R745 source.n220 source.n176 104.615
R746 source.n213 source.n176 104.615
R747 source.n213 source.n212 104.615
R748 source.n212 source.n211 104.615
R749 source.n211 source.n180 104.615
R750 source.n204 source.n180 104.615
R751 source.n204 source.n203 104.615
R752 source.n203 source.n185 104.615
R753 source.n196 source.n185 104.615
R754 source.n196 source.n195 104.615
R755 source.n195 source.n189 104.615
R756 source.t8 source.n479 52.3082
R757 source.t11 source.n335 52.3082
R758 source.t16 source.n45 52.3082
R759 source.t7 source.n189 52.3082
R760 source.n435 source.n434 42.0366
R761 source.n433 source.n432 42.0366
R762 source.n291 source.n290 42.0366
R763 source.n289 source.n288 42.0366
R764 source.n141 source.n140 42.0366
R765 source.n143 source.n142 42.0366
R766 source.n285 source.n284 42.0366
R767 source.n287 source.n286 42.0366
R768 source.n289 source.n287 32.05
R769 source.n575 source.n574 30.6338
R770 source.n431 source.n430 30.6338
R771 source.n139 source.n138 30.6338
R772 source.n283 source.n282 30.6338
R773 source.n576 source.n139 26.1017
R774 source.n505 source.n470 13.1884
R775 source.n552 source.n551 13.1884
R776 source.n361 source.n326 13.1884
R777 source.n408 source.n407 13.1884
R778 source.n116 source.n115 13.1884
R779 source.n70 source.n35 13.1884
R780 source.n260 source.n259 13.1884
R781 source.n214 source.n179 13.1884
R782 source.n501 source.n500 12.8005
R783 source.n506 source.n468 12.8005
R784 source.n550 source.n448 12.8005
R785 source.n555 source.n446 12.8005
R786 source.n357 source.n356 12.8005
R787 source.n362 source.n324 12.8005
R788 source.n406 source.n304 12.8005
R789 source.n411 source.n302 12.8005
R790 source.n119 source.n10 12.8005
R791 source.n114 source.n12 12.8005
R792 source.n71 source.n33 12.8005
R793 source.n66 source.n37 12.8005
R794 source.n263 source.n154 12.8005
R795 source.n258 source.n156 12.8005
R796 source.n215 source.n177 12.8005
R797 source.n210 source.n181 12.8005
R798 source.n499 source.n472 12.0247
R799 source.n510 source.n509 12.0247
R800 source.n547 source.n546 12.0247
R801 source.n556 source.n444 12.0247
R802 source.n355 source.n328 12.0247
R803 source.n366 source.n365 12.0247
R804 source.n403 source.n402 12.0247
R805 source.n412 source.n300 12.0247
R806 source.n120 source.n8 12.0247
R807 source.n111 source.n110 12.0247
R808 source.n75 source.n74 12.0247
R809 source.n65 source.n38 12.0247
R810 source.n264 source.n152 12.0247
R811 source.n255 source.n254 12.0247
R812 source.n219 source.n218 12.0247
R813 source.n209 source.n182 12.0247
R814 source.n496 source.n495 11.249
R815 source.n513 source.n466 11.249
R816 source.n542 source.n450 11.249
R817 source.n560 source.n559 11.249
R818 source.n352 source.n351 11.249
R819 source.n369 source.n322 11.249
R820 source.n398 source.n306 11.249
R821 source.n416 source.n415 11.249
R822 source.n124 source.n123 11.249
R823 source.n107 source.n14 11.249
R824 source.n78 source.n31 11.249
R825 source.n62 source.n61 11.249
R826 source.n268 source.n267 11.249
R827 source.n251 source.n158 11.249
R828 source.n222 source.n175 11.249
R829 source.n206 source.n205 11.249
R830 source.n492 source.n474 10.4732
R831 source.n514 source.n464 10.4732
R832 source.n541 source.n452 10.4732
R833 source.n563 source.n442 10.4732
R834 source.n348 source.n330 10.4732
R835 source.n370 source.n320 10.4732
R836 source.n397 source.n308 10.4732
R837 source.n419 source.n298 10.4732
R838 source.n127 source.n6 10.4732
R839 source.n106 source.n17 10.4732
R840 source.n79 source.n29 10.4732
R841 source.n58 source.n40 10.4732
R842 source.n271 source.n150 10.4732
R843 source.n250 source.n161 10.4732
R844 source.n223 source.n173 10.4732
R845 source.n202 source.n184 10.4732
R846 source.n481 source.n480 10.2747
R847 source.n337 source.n336 10.2747
R848 source.n47 source.n46 10.2747
R849 source.n191 source.n190 10.2747
R850 source.n491 source.n476 9.69747
R851 source.n518 source.n517 9.69747
R852 source.n538 source.n537 9.69747
R853 source.n564 source.n440 9.69747
R854 source.n347 source.n332 9.69747
R855 source.n374 source.n373 9.69747
R856 source.n394 source.n393 9.69747
R857 source.n420 source.n296 9.69747
R858 source.n128 source.n4 9.69747
R859 source.n103 source.n102 9.69747
R860 source.n83 source.n82 9.69747
R861 source.n57 source.n42 9.69747
R862 source.n272 source.n148 9.69747
R863 source.n247 source.n246 9.69747
R864 source.n227 source.n226 9.69747
R865 source.n201 source.n186 9.69747
R866 source.n574 source.n573 9.45567
R867 source.n430 source.n429 9.45567
R868 source.n138 source.n137 9.45567
R869 source.n282 source.n281 9.45567
R870 source.n438 source.n437 9.3005
R871 source.n567 source.n566 9.3005
R872 source.n565 source.n564 9.3005
R873 source.n442 source.n441 9.3005
R874 source.n559 source.n558 9.3005
R875 source.n557 source.n556 9.3005
R876 source.n446 source.n445 9.3005
R877 source.n525 source.n524 9.3005
R878 source.n523 source.n522 9.3005
R879 source.n462 source.n461 9.3005
R880 source.n517 source.n516 9.3005
R881 source.n515 source.n514 9.3005
R882 source.n466 source.n465 9.3005
R883 source.n509 source.n508 9.3005
R884 source.n507 source.n506 9.3005
R885 source.n483 source.n482 9.3005
R886 source.n478 source.n477 9.3005
R887 source.n489 source.n488 9.3005
R888 source.n491 source.n490 9.3005
R889 source.n474 source.n473 9.3005
R890 source.n497 source.n496 9.3005
R891 source.n499 source.n498 9.3005
R892 source.n500 source.n469 9.3005
R893 source.n458 source.n457 9.3005
R894 source.n531 source.n530 9.3005
R895 source.n533 source.n532 9.3005
R896 source.n454 source.n453 9.3005
R897 source.n539 source.n538 9.3005
R898 source.n541 source.n540 9.3005
R899 source.n450 source.n449 9.3005
R900 source.n548 source.n547 9.3005
R901 source.n550 source.n549 9.3005
R902 source.n573 source.n572 9.3005
R903 source.n294 source.n293 9.3005
R904 source.n423 source.n422 9.3005
R905 source.n421 source.n420 9.3005
R906 source.n298 source.n297 9.3005
R907 source.n415 source.n414 9.3005
R908 source.n413 source.n412 9.3005
R909 source.n302 source.n301 9.3005
R910 source.n381 source.n380 9.3005
R911 source.n379 source.n378 9.3005
R912 source.n318 source.n317 9.3005
R913 source.n373 source.n372 9.3005
R914 source.n371 source.n370 9.3005
R915 source.n322 source.n321 9.3005
R916 source.n365 source.n364 9.3005
R917 source.n363 source.n362 9.3005
R918 source.n339 source.n338 9.3005
R919 source.n334 source.n333 9.3005
R920 source.n345 source.n344 9.3005
R921 source.n347 source.n346 9.3005
R922 source.n330 source.n329 9.3005
R923 source.n353 source.n352 9.3005
R924 source.n355 source.n354 9.3005
R925 source.n356 source.n325 9.3005
R926 source.n314 source.n313 9.3005
R927 source.n387 source.n386 9.3005
R928 source.n389 source.n388 9.3005
R929 source.n310 source.n309 9.3005
R930 source.n395 source.n394 9.3005
R931 source.n397 source.n396 9.3005
R932 source.n306 source.n305 9.3005
R933 source.n404 source.n403 9.3005
R934 source.n406 source.n405 9.3005
R935 source.n429 source.n428 9.3005
R936 source.n49 source.n48 9.3005
R937 source.n44 source.n43 9.3005
R938 source.n55 source.n54 9.3005
R939 source.n57 source.n56 9.3005
R940 source.n40 source.n39 9.3005
R941 source.n63 source.n62 9.3005
R942 source.n65 source.n64 9.3005
R943 source.n37 source.n34 9.3005
R944 source.n96 source.n95 9.3005
R945 source.n98 source.n97 9.3005
R946 source.n19 source.n18 9.3005
R947 source.n104 source.n103 9.3005
R948 source.n106 source.n105 9.3005
R949 source.n14 source.n13 9.3005
R950 source.n112 source.n111 9.3005
R951 source.n114 source.n113 9.3005
R952 source.n137 source.n136 9.3005
R953 source.n2 source.n1 9.3005
R954 source.n131 source.n130 9.3005
R955 source.n129 source.n128 9.3005
R956 source.n6 source.n5 9.3005
R957 source.n123 source.n122 9.3005
R958 source.n121 source.n120 9.3005
R959 source.n10 source.n9 9.3005
R960 source.n23 source.n22 9.3005
R961 source.n90 source.n89 9.3005
R962 source.n88 source.n87 9.3005
R963 source.n27 source.n26 9.3005
R964 source.n82 source.n81 9.3005
R965 source.n80 source.n79 9.3005
R966 source.n31 source.n30 9.3005
R967 source.n74 source.n73 9.3005
R968 source.n72 source.n71 9.3005
R969 source.n193 source.n192 9.3005
R970 source.n188 source.n187 9.3005
R971 source.n199 source.n198 9.3005
R972 source.n201 source.n200 9.3005
R973 source.n184 source.n183 9.3005
R974 source.n207 source.n206 9.3005
R975 source.n209 source.n208 9.3005
R976 source.n181 source.n178 9.3005
R977 source.n240 source.n239 9.3005
R978 source.n242 source.n241 9.3005
R979 source.n163 source.n162 9.3005
R980 source.n248 source.n247 9.3005
R981 source.n250 source.n249 9.3005
R982 source.n158 source.n157 9.3005
R983 source.n256 source.n255 9.3005
R984 source.n258 source.n257 9.3005
R985 source.n281 source.n280 9.3005
R986 source.n146 source.n145 9.3005
R987 source.n275 source.n274 9.3005
R988 source.n273 source.n272 9.3005
R989 source.n150 source.n149 9.3005
R990 source.n267 source.n266 9.3005
R991 source.n265 source.n264 9.3005
R992 source.n154 source.n153 9.3005
R993 source.n167 source.n166 9.3005
R994 source.n234 source.n233 9.3005
R995 source.n232 source.n231 9.3005
R996 source.n171 source.n170 9.3005
R997 source.n226 source.n225 9.3005
R998 source.n224 source.n223 9.3005
R999 source.n175 source.n174 9.3005
R1000 source.n218 source.n217 9.3005
R1001 source.n216 source.n215 9.3005
R1002 source.n488 source.n487 8.92171
R1003 source.n521 source.n462 8.92171
R1004 source.n534 source.n454 8.92171
R1005 source.n568 source.n567 8.92171
R1006 source.n344 source.n343 8.92171
R1007 source.n377 source.n318 8.92171
R1008 source.n390 source.n310 8.92171
R1009 source.n424 source.n423 8.92171
R1010 source.n132 source.n131 8.92171
R1011 source.n99 source.n19 8.92171
R1012 source.n86 source.n27 8.92171
R1013 source.n54 source.n53 8.92171
R1014 source.n276 source.n275 8.92171
R1015 source.n243 source.n163 8.92171
R1016 source.n230 source.n171 8.92171
R1017 source.n198 source.n197 8.92171
R1018 source.n484 source.n478 8.14595
R1019 source.n522 source.n460 8.14595
R1020 source.n533 source.n456 8.14595
R1021 source.n571 source.n438 8.14595
R1022 source.n340 source.n334 8.14595
R1023 source.n378 source.n316 8.14595
R1024 source.n389 source.n312 8.14595
R1025 source.n427 source.n294 8.14595
R1026 source.n135 source.n2 8.14595
R1027 source.n98 source.n21 8.14595
R1028 source.n87 source.n25 8.14595
R1029 source.n50 source.n44 8.14595
R1030 source.n279 source.n146 8.14595
R1031 source.n242 source.n165 8.14595
R1032 source.n231 source.n169 8.14595
R1033 source.n194 source.n188 8.14595
R1034 source.n483 source.n480 7.3702
R1035 source.n526 source.n525 7.3702
R1036 source.n530 source.n529 7.3702
R1037 source.n572 source.n436 7.3702
R1038 source.n339 source.n336 7.3702
R1039 source.n382 source.n381 7.3702
R1040 source.n386 source.n385 7.3702
R1041 source.n428 source.n292 7.3702
R1042 source.n136 source.n0 7.3702
R1043 source.n95 source.n94 7.3702
R1044 source.n91 source.n90 7.3702
R1045 source.n49 source.n46 7.3702
R1046 source.n280 source.n144 7.3702
R1047 source.n239 source.n238 7.3702
R1048 source.n235 source.n234 7.3702
R1049 source.n193 source.n190 7.3702
R1050 source.n526 source.n458 6.59444
R1051 source.n529 source.n458 6.59444
R1052 source.n574 source.n436 6.59444
R1053 source.n382 source.n314 6.59444
R1054 source.n385 source.n314 6.59444
R1055 source.n430 source.n292 6.59444
R1056 source.n138 source.n0 6.59444
R1057 source.n94 source.n23 6.59444
R1058 source.n91 source.n23 6.59444
R1059 source.n282 source.n144 6.59444
R1060 source.n238 source.n167 6.59444
R1061 source.n235 source.n167 6.59444
R1062 source.n484 source.n483 5.81868
R1063 source.n525 source.n460 5.81868
R1064 source.n530 source.n456 5.81868
R1065 source.n572 source.n571 5.81868
R1066 source.n340 source.n339 5.81868
R1067 source.n381 source.n316 5.81868
R1068 source.n386 source.n312 5.81868
R1069 source.n428 source.n427 5.81868
R1070 source.n136 source.n135 5.81868
R1071 source.n95 source.n21 5.81868
R1072 source.n90 source.n25 5.81868
R1073 source.n50 source.n49 5.81868
R1074 source.n280 source.n279 5.81868
R1075 source.n239 source.n165 5.81868
R1076 source.n234 source.n169 5.81868
R1077 source.n194 source.n193 5.81868
R1078 source.n576 source.n575 5.49188
R1079 source.n487 source.n478 5.04292
R1080 source.n522 source.n521 5.04292
R1081 source.n534 source.n533 5.04292
R1082 source.n568 source.n438 5.04292
R1083 source.n343 source.n334 5.04292
R1084 source.n378 source.n377 5.04292
R1085 source.n390 source.n389 5.04292
R1086 source.n424 source.n294 5.04292
R1087 source.n132 source.n2 5.04292
R1088 source.n99 source.n98 5.04292
R1089 source.n87 source.n86 5.04292
R1090 source.n53 source.n44 5.04292
R1091 source.n276 source.n146 5.04292
R1092 source.n243 source.n242 5.04292
R1093 source.n231 source.n230 5.04292
R1094 source.n197 source.n188 5.04292
R1095 source.n488 source.n476 4.26717
R1096 source.n518 source.n462 4.26717
R1097 source.n537 source.n454 4.26717
R1098 source.n567 source.n440 4.26717
R1099 source.n344 source.n332 4.26717
R1100 source.n374 source.n318 4.26717
R1101 source.n393 source.n310 4.26717
R1102 source.n423 source.n296 4.26717
R1103 source.n131 source.n4 4.26717
R1104 source.n102 source.n19 4.26717
R1105 source.n83 source.n27 4.26717
R1106 source.n54 source.n42 4.26717
R1107 source.n275 source.n148 4.26717
R1108 source.n246 source.n163 4.26717
R1109 source.n227 source.n171 4.26717
R1110 source.n198 source.n186 4.26717
R1111 source.n492 source.n491 3.49141
R1112 source.n517 source.n464 3.49141
R1113 source.n538 source.n452 3.49141
R1114 source.n564 source.n563 3.49141
R1115 source.n348 source.n347 3.49141
R1116 source.n373 source.n320 3.49141
R1117 source.n394 source.n308 3.49141
R1118 source.n420 source.n419 3.49141
R1119 source.n128 source.n127 3.49141
R1120 source.n103 source.n17 3.49141
R1121 source.n82 source.n29 3.49141
R1122 source.n58 source.n57 3.49141
R1123 source.n272 source.n271 3.49141
R1124 source.n247 source.n161 3.49141
R1125 source.n226 source.n173 3.49141
R1126 source.n202 source.n201 3.49141
R1127 source.n48 source.n47 2.84303
R1128 source.n192 source.n191 2.84303
R1129 source.n482 source.n481 2.84303
R1130 source.n338 source.n337 2.84303
R1131 source.n495 source.n474 2.71565
R1132 source.n514 source.n513 2.71565
R1133 source.n542 source.n541 2.71565
R1134 source.n560 source.n442 2.71565
R1135 source.n351 source.n330 2.71565
R1136 source.n370 source.n369 2.71565
R1137 source.n398 source.n397 2.71565
R1138 source.n416 source.n298 2.71565
R1139 source.n124 source.n6 2.71565
R1140 source.n107 source.n106 2.71565
R1141 source.n79 source.n78 2.71565
R1142 source.n61 source.n40 2.71565
R1143 source.n268 source.n150 2.71565
R1144 source.n251 source.n250 2.71565
R1145 source.n223 source.n222 2.71565
R1146 source.n205 source.n184 2.71565
R1147 source.n496 source.n472 1.93989
R1148 source.n510 source.n466 1.93989
R1149 source.n546 source.n450 1.93989
R1150 source.n559 source.n444 1.93989
R1151 source.n352 source.n328 1.93989
R1152 source.n366 source.n322 1.93989
R1153 source.n402 source.n306 1.93989
R1154 source.n415 source.n300 1.93989
R1155 source.n123 source.n8 1.93989
R1156 source.n110 source.n14 1.93989
R1157 source.n75 source.n31 1.93989
R1158 source.n62 source.n38 1.93989
R1159 source.n267 source.n152 1.93989
R1160 source.n254 source.n158 1.93989
R1161 source.n219 source.n175 1.93989
R1162 source.n206 source.n182 1.93989
R1163 source.n501 source.n499 1.16414
R1164 source.n509 source.n468 1.16414
R1165 source.n547 source.n448 1.16414
R1166 source.n556 source.n555 1.16414
R1167 source.n357 source.n355 1.16414
R1168 source.n365 source.n324 1.16414
R1169 source.n403 source.n304 1.16414
R1170 source.n412 source.n411 1.16414
R1171 source.n120 source.n119 1.16414
R1172 source.n111 source.n12 1.16414
R1173 source.n74 source.n33 1.16414
R1174 source.n66 source.n65 1.16414
R1175 source.n264 source.n263 1.16414
R1176 source.n255 source.n156 1.16414
R1177 source.n218 source.n177 1.16414
R1178 source.n210 source.n209 1.16414
R1179 source.n434 source.t5 0.7925
R1180 source.n434 source.t2 0.7925
R1181 source.n432 source.t3 0.7925
R1182 source.n432 source.t6 0.7925
R1183 source.n290 source.t10 0.7925
R1184 source.n290 source.t19 0.7925
R1185 source.n288 source.t13 0.7925
R1186 source.n288 source.t14 0.7925
R1187 source.n140 source.t12 0.7925
R1188 source.n140 source.t15 0.7925
R1189 source.n142 source.t17 0.7925
R1190 source.n142 source.t18 0.7925
R1191 source.n284 source.t0 0.7925
R1192 source.n284 source.t9 0.7925
R1193 source.n286 source.t1 0.7925
R1194 source.n286 source.t4 0.7925
R1195 source.n283 source.n143 0.698776
R1196 source.n433 source.n431 0.698776
R1197 source.n287 source.n285 0.457397
R1198 source.n285 source.n283 0.457397
R1199 source.n143 source.n141 0.457397
R1200 source.n141 source.n139 0.457397
R1201 source.n291 source.n289 0.457397
R1202 source.n431 source.n291 0.457397
R1203 source.n435 source.n433 0.457397
R1204 source.n575 source.n435 0.457397
R1205 source.n500 source.n470 0.388379
R1206 source.n506 source.n505 0.388379
R1207 source.n551 source.n550 0.388379
R1208 source.n552 source.n446 0.388379
R1209 source.n356 source.n326 0.388379
R1210 source.n362 source.n361 0.388379
R1211 source.n407 source.n406 0.388379
R1212 source.n408 source.n302 0.388379
R1213 source.n116 source.n10 0.388379
R1214 source.n115 source.n114 0.388379
R1215 source.n71 source.n70 0.388379
R1216 source.n37 source.n35 0.388379
R1217 source.n260 source.n154 0.388379
R1218 source.n259 source.n258 0.388379
R1219 source.n215 source.n214 0.388379
R1220 source.n181 source.n179 0.388379
R1221 source source.n576 0.188
R1222 source.n482 source.n477 0.155672
R1223 source.n489 source.n477 0.155672
R1224 source.n490 source.n489 0.155672
R1225 source.n490 source.n473 0.155672
R1226 source.n497 source.n473 0.155672
R1227 source.n498 source.n497 0.155672
R1228 source.n498 source.n469 0.155672
R1229 source.n507 source.n469 0.155672
R1230 source.n508 source.n507 0.155672
R1231 source.n508 source.n465 0.155672
R1232 source.n515 source.n465 0.155672
R1233 source.n516 source.n515 0.155672
R1234 source.n516 source.n461 0.155672
R1235 source.n523 source.n461 0.155672
R1236 source.n524 source.n523 0.155672
R1237 source.n524 source.n457 0.155672
R1238 source.n531 source.n457 0.155672
R1239 source.n532 source.n531 0.155672
R1240 source.n532 source.n453 0.155672
R1241 source.n539 source.n453 0.155672
R1242 source.n540 source.n539 0.155672
R1243 source.n540 source.n449 0.155672
R1244 source.n548 source.n449 0.155672
R1245 source.n549 source.n548 0.155672
R1246 source.n549 source.n445 0.155672
R1247 source.n557 source.n445 0.155672
R1248 source.n558 source.n557 0.155672
R1249 source.n558 source.n441 0.155672
R1250 source.n565 source.n441 0.155672
R1251 source.n566 source.n565 0.155672
R1252 source.n566 source.n437 0.155672
R1253 source.n573 source.n437 0.155672
R1254 source.n338 source.n333 0.155672
R1255 source.n345 source.n333 0.155672
R1256 source.n346 source.n345 0.155672
R1257 source.n346 source.n329 0.155672
R1258 source.n353 source.n329 0.155672
R1259 source.n354 source.n353 0.155672
R1260 source.n354 source.n325 0.155672
R1261 source.n363 source.n325 0.155672
R1262 source.n364 source.n363 0.155672
R1263 source.n364 source.n321 0.155672
R1264 source.n371 source.n321 0.155672
R1265 source.n372 source.n371 0.155672
R1266 source.n372 source.n317 0.155672
R1267 source.n379 source.n317 0.155672
R1268 source.n380 source.n379 0.155672
R1269 source.n380 source.n313 0.155672
R1270 source.n387 source.n313 0.155672
R1271 source.n388 source.n387 0.155672
R1272 source.n388 source.n309 0.155672
R1273 source.n395 source.n309 0.155672
R1274 source.n396 source.n395 0.155672
R1275 source.n396 source.n305 0.155672
R1276 source.n404 source.n305 0.155672
R1277 source.n405 source.n404 0.155672
R1278 source.n405 source.n301 0.155672
R1279 source.n413 source.n301 0.155672
R1280 source.n414 source.n413 0.155672
R1281 source.n414 source.n297 0.155672
R1282 source.n421 source.n297 0.155672
R1283 source.n422 source.n421 0.155672
R1284 source.n422 source.n293 0.155672
R1285 source.n429 source.n293 0.155672
R1286 source.n137 source.n1 0.155672
R1287 source.n130 source.n1 0.155672
R1288 source.n130 source.n129 0.155672
R1289 source.n129 source.n5 0.155672
R1290 source.n122 source.n5 0.155672
R1291 source.n122 source.n121 0.155672
R1292 source.n121 source.n9 0.155672
R1293 source.n113 source.n9 0.155672
R1294 source.n113 source.n112 0.155672
R1295 source.n112 source.n13 0.155672
R1296 source.n105 source.n13 0.155672
R1297 source.n105 source.n104 0.155672
R1298 source.n104 source.n18 0.155672
R1299 source.n97 source.n18 0.155672
R1300 source.n97 source.n96 0.155672
R1301 source.n96 source.n22 0.155672
R1302 source.n89 source.n22 0.155672
R1303 source.n89 source.n88 0.155672
R1304 source.n88 source.n26 0.155672
R1305 source.n81 source.n26 0.155672
R1306 source.n81 source.n80 0.155672
R1307 source.n80 source.n30 0.155672
R1308 source.n73 source.n30 0.155672
R1309 source.n73 source.n72 0.155672
R1310 source.n72 source.n34 0.155672
R1311 source.n64 source.n34 0.155672
R1312 source.n64 source.n63 0.155672
R1313 source.n63 source.n39 0.155672
R1314 source.n56 source.n39 0.155672
R1315 source.n56 source.n55 0.155672
R1316 source.n55 source.n43 0.155672
R1317 source.n48 source.n43 0.155672
R1318 source.n281 source.n145 0.155672
R1319 source.n274 source.n145 0.155672
R1320 source.n274 source.n273 0.155672
R1321 source.n273 source.n149 0.155672
R1322 source.n266 source.n149 0.155672
R1323 source.n266 source.n265 0.155672
R1324 source.n265 source.n153 0.155672
R1325 source.n257 source.n153 0.155672
R1326 source.n257 source.n256 0.155672
R1327 source.n256 source.n157 0.155672
R1328 source.n249 source.n157 0.155672
R1329 source.n249 source.n248 0.155672
R1330 source.n248 source.n162 0.155672
R1331 source.n241 source.n162 0.155672
R1332 source.n241 source.n240 0.155672
R1333 source.n240 source.n166 0.155672
R1334 source.n233 source.n166 0.155672
R1335 source.n233 source.n232 0.155672
R1336 source.n232 source.n170 0.155672
R1337 source.n225 source.n170 0.155672
R1338 source.n225 source.n224 0.155672
R1339 source.n224 source.n174 0.155672
R1340 source.n217 source.n174 0.155672
R1341 source.n217 source.n216 0.155672
R1342 source.n216 source.n178 0.155672
R1343 source.n208 source.n178 0.155672
R1344 source.n208 source.n207 0.155672
R1345 source.n207 source.n183 0.155672
R1346 source.n200 source.n183 0.155672
R1347 source.n200 source.n199 0.155672
R1348 source.n199 source.n187 0.155672
R1349 source.n192 source.n187 0.155672
R1350 minus.n8 minus.t8 3214.43
R1351 minus.n2 minus.t7 3214.43
R1352 minus.n18 minus.t6 3214.43
R1353 minus.n12 minus.t2 3214.43
R1354 minus.n7 minus.t9 3169.15
R1355 minus.n5 minus.t0 3169.15
R1356 minus.n1 minus.t3 3169.15
R1357 minus.n17 minus.t4 3169.15
R1358 minus.n15 minus.t1 3169.15
R1359 minus.n11 minus.t5 3169.15
R1360 minus.n3 minus.n2 161.489
R1361 minus.n13 minus.n12 161.489
R1362 minus.n9 minus.n8 161.3
R1363 minus.n6 minus.n0 161.3
R1364 minus.n4 minus.n3 161.3
R1365 minus.n19 minus.n18 161.3
R1366 minus.n16 minus.n10 161.3
R1367 minus.n14 minus.n13 161.3
R1368 minus.n20 minus.n9 44.0403
R1369 minus.n7 minus.n6 40.8975
R1370 minus.n4 minus.n1 40.8975
R1371 minus.n14 minus.n11 40.8975
R1372 minus.n17 minus.n16 40.8975
R1373 minus.n6 minus.n5 36.5157
R1374 minus.n5 minus.n4 36.5157
R1375 minus.n15 minus.n14 36.5157
R1376 minus.n16 minus.n15 36.5157
R1377 minus.n8 minus.n7 32.1338
R1378 minus.n2 minus.n1 32.1338
R1379 minus.n12 minus.n11 32.1338
R1380 minus.n18 minus.n17 32.1338
R1381 minus.n20 minus.n19 6.44936
R1382 minus.n9 minus.n0 0.189894
R1383 minus.n3 minus.n0 0.189894
R1384 minus.n13 minus.n10 0.189894
R1385 minus.n19 minus.n10 0.189894
R1386 minus minus.n20 0.188
R1387 drain_right.n134 drain_right.n0 289.615
R1388 drain_right.n280 drain_right.n146 289.615
R1389 drain_right.n44 drain_right.n43 185
R1390 drain_right.n49 drain_right.n48 185
R1391 drain_right.n51 drain_right.n50 185
R1392 drain_right.n40 drain_right.n39 185
R1393 drain_right.n57 drain_right.n56 185
R1394 drain_right.n59 drain_right.n58 185
R1395 drain_right.n36 drain_right.n35 185
R1396 drain_right.n66 drain_right.n65 185
R1397 drain_right.n67 drain_right.n34 185
R1398 drain_right.n69 drain_right.n68 185
R1399 drain_right.n32 drain_right.n31 185
R1400 drain_right.n75 drain_right.n74 185
R1401 drain_right.n77 drain_right.n76 185
R1402 drain_right.n28 drain_right.n27 185
R1403 drain_right.n83 drain_right.n82 185
R1404 drain_right.n85 drain_right.n84 185
R1405 drain_right.n24 drain_right.n23 185
R1406 drain_right.n91 drain_right.n90 185
R1407 drain_right.n93 drain_right.n92 185
R1408 drain_right.n20 drain_right.n19 185
R1409 drain_right.n99 drain_right.n98 185
R1410 drain_right.n101 drain_right.n100 185
R1411 drain_right.n16 drain_right.n15 185
R1412 drain_right.n107 drain_right.n106 185
R1413 drain_right.n110 drain_right.n109 185
R1414 drain_right.n108 drain_right.n12 185
R1415 drain_right.n115 drain_right.n11 185
R1416 drain_right.n117 drain_right.n116 185
R1417 drain_right.n119 drain_right.n118 185
R1418 drain_right.n8 drain_right.n7 185
R1419 drain_right.n125 drain_right.n124 185
R1420 drain_right.n127 drain_right.n126 185
R1421 drain_right.n4 drain_right.n3 185
R1422 drain_right.n133 drain_right.n132 185
R1423 drain_right.n135 drain_right.n134 185
R1424 drain_right.n281 drain_right.n280 185
R1425 drain_right.n279 drain_right.n278 185
R1426 drain_right.n150 drain_right.n149 185
R1427 drain_right.n273 drain_right.n272 185
R1428 drain_right.n271 drain_right.n270 185
R1429 drain_right.n154 drain_right.n153 185
R1430 drain_right.n265 drain_right.n264 185
R1431 drain_right.n263 drain_right.n262 185
R1432 drain_right.n261 drain_right.n157 185
R1433 drain_right.n161 drain_right.n158 185
R1434 drain_right.n256 drain_right.n255 185
R1435 drain_right.n254 drain_right.n253 185
R1436 drain_right.n163 drain_right.n162 185
R1437 drain_right.n248 drain_right.n247 185
R1438 drain_right.n246 drain_right.n245 185
R1439 drain_right.n167 drain_right.n166 185
R1440 drain_right.n240 drain_right.n239 185
R1441 drain_right.n238 drain_right.n237 185
R1442 drain_right.n171 drain_right.n170 185
R1443 drain_right.n232 drain_right.n231 185
R1444 drain_right.n230 drain_right.n229 185
R1445 drain_right.n175 drain_right.n174 185
R1446 drain_right.n224 drain_right.n223 185
R1447 drain_right.n222 drain_right.n221 185
R1448 drain_right.n179 drain_right.n178 185
R1449 drain_right.n216 drain_right.n215 185
R1450 drain_right.n214 drain_right.n181 185
R1451 drain_right.n213 drain_right.n212 185
R1452 drain_right.n184 drain_right.n182 185
R1453 drain_right.n207 drain_right.n206 185
R1454 drain_right.n205 drain_right.n204 185
R1455 drain_right.n188 drain_right.n187 185
R1456 drain_right.n199 drain_right.n198 185
R1457 drain_right.n197 drain_right.n196 185
R1458 drain_right.n192 drain_right.n191 185
R1459 drain_right.n45 drain_right.t7 149.524
R1460 drain_right.n193 drain_right.t1 149.524
R1461 drain_right.n49 drain_right.n43 104.615
R1462 drain_right.n50 drain_right.n49 104.615
R1463 drain_right.n50 drain_right.n39 104.615
R1464 drain_right.n57 drain_right.n39 104.615
R1465 drain_right.n58 drain_right.n57 104.615
R1466 drain_right.n58 drain_right.n35 104.615
R1467 drain_right.n66 drain_right.n35 104.615
R1468 drain_right.n67 drain_right.n66 104.615
R1469 drain_right.n68 drain_right.n67 104.615
R1470 drain_right.n68 drain_right.n31 104.615
R1471 drain_right.n75 drain_right.n31 104.615
R1472 drain_right.n76 drain_right.n75 104.615
R1473 drain_right.n76 drain_right.n27 104.615
R1474 drain_right.n83 drain_right.n27 104.615
R1475 drain_right.n84 drain_right.n83 104.615
R1476 drain_right.n84 drain_right.n23 104.615
R1477 drain_right.n91 drain_right.n23 104.615
R1478 drain_right.n92 drain_right.n91 104.615
R1479 drain_right.n92 drain_right.n19 104.615
R1480 drain_right.n99 drain_right.n19 104.615
R1481 drain_right.n100 drain_right.n99 104.615
R1482 drain_right.n100 drain_right.n15 104.615
R1483 drain_right.n107 drain_right.n15 104.615
R1484 drain_right.n109 drain_right.n107 104.615
R1485 drain_right.n109 drain_right.n108 104.615
R1486 drain_right.n108 drain_right.n11 104.615
R1487 drain_right.n117 drain_right.n11 104.615
R1488 drain_right.n118 drain_right.n117 104.615
R1489 drain_right.n118 drain_right.n7 104.615
R1490 drain_right.n125 drain_right.n7 104.615
R1491 drain_right.n126 drain_right.n125 104.615
R1492 drain_right.n126 drain_right.n3 104.615
R1493 drain_right.n133 drain_right.n3 104.615
R1494 drain_right.n134 drain_right.n133 104.615
R1495 drain_right.n280 drain_right.n279 104.615
R1496 drain_right.n279 drain_right.n149 104.615
R1497 drain_right.n272 drain_right.n149 104.615
R1498 drain_right.n272 drain_right.n271 104.615
R1499 drain_right.n271 drain_right.n153 104.615
R1500 drain_right.n264 drain_right.n153 104.615
R1501 drain_right.n264 drain_right.n263 104.615
R1502 drain_right.n263 drain_right.n157 104.615
R1503 drain_right.n161 drain_right.n157 104.615
R1504 drain_right.n255 drain_right.n161 104.615
R1505 drain_right.n255 drain_right.n254 104.615
R1506 drain_right.n254 drain_right.n162 104.615
R1507 drain_right.n247 drain_right.n162 104.615
R1508 drain_right.n247 drain_right.n246 104.615
R1509 drain_right.n246 drain_right.n166 104.615
R1510 drain_right.n239 drain_right.n166 104.615
R1511 drain_right.n239 drain_right.n238 104.615
R1512 drain_right.n238 drain_right.n170 104.615
R1513 drain_right.n231 drain_right.n170 104.615
R1514 drain_right.n231 drain_right.n230 104.615
R1515 drain_right.n230 drain_right.n174 104.615
R1516 drain_right.n223 drain_right.n174 104.615
R1517 drain_right.n223 drain_right.n222 104.615
R1518 drain_right.n222 drain_right.n178 104.615
R1519 drain_right.n215 drain_right.n178 104.615
R1520 drain_right.n215 drain_right.n214 104.615
R1521 drain_right.n214 drain_right.n213 104.615
R1522 drain_right.n213 drain_right.n182 104.615
R1523 drain_right.n206 drain_right.n182 104.615
R1524 drain_right.n206 drain_right.n205 104.615
R1525 drain_right.n205 drain_right.n187 104.615
R1526 drain_right.n198 drain_right.n187 104.615
R1527 drain_right.n198 drain_right.n197 104.615
R1528 drain_right.n197 drain_right.n191 104.615
R1529 drain_right.n145 drain_right.n143 59.1722
R1530 drain_right.n142 drain_right.n141 59.0028
R1531 drain_right.n140 drain_right.n139 58.7154
R1532 drain_right.n145 drain_right.n144 58.7154
R1533 drain_right.t7 drain_right.n43 52.3082
R1534 drain_right.t1 drain_right.n191 52.3082
R1535 drain_right.n140 drain_right.n138 47.7695
R1536 drain_right.n285 drain_right.n284 47.3126
R1537 drain_right drain_right.n142 38.6041
R1538 drain_right.n69 drain_right.n34 13.1884
R1539 drain_right.n116 drain_right.n115 13.1884
R1540 drain_right.n262 drain_right.n261 13.1884
R1541 drain_right.n216 drain_right.n181 13.1884
R1542 drain_right.n65 drain_right.n64 12.8005
R1543 drain_right.n70 drain_right.n32 12.8005
R1544 drain_right.n114 drain_right.n12 12.8005
R1545 drain_right.n119 drain_right.n10 12.8005
R1546 drain_right.n265 drain_right.n156 12.8005
R1547 drain_right.n260 drain_right.n158 12.8005
R1548 drain_right.n217 drain_right.n179 12.8005
R1549 drain_right.n212 drain_right.n183 12.8005
R1550 drain_right.n63 drain_right.n36 12.0247
R1551 drain_right.n74 drain_right.n73 12.0247
R1552 drain_right.n111 drain_right.n110 12.0247
R1553 drain_right.n120 drain_right.n8 12.0247
R1554 drain_right.n266 drain_right.n154 12.0247
R1555 drain_right.n257 drain_right.n256 12.0247
R1556 drain_right.n221 drain_right.n220 12.0247
R1557 drain_right.n211 drain_right.n184 12.0247
R1558 drain_right.n60 drain_right.n59 11.249
R1559 drain_right.n77 drain_right.n30 11.249
R1560 drain_right.n106 drain_right.n14 11.249
R1561 drain_right.n124 drain_right.n123 11.249
R1562 drain_right.n270 drain_right.n269 11.249
R1563 drain_right.n253 drain_right.n160 11.249
R1564 drain_right.n224 drain_right.n177 11.249
R1565 drain_right.n208 drain_right.n207 11.249
R1566 drain_right.n56 drain_right.n38 10.4732
R1567 drain_right.n78 drain_right.n28 10.4732
R1568 drain_right.n105 drain_right.n16 10.4732
R1569 drain_right.n127 drain_right.n6 10.4732
R1570 drain_right.n273 drain_right.n152 10.4732
R1571 drain_right.n252 drain_right.n163 10.4732
R1572 drain_right.n225 drain_right.n175 10.4732
R1573 drain_right.n204 drain_right.n186 10.4732
R1574 drain_right.n45 drain_right.n44 10.2747
R1575 drain_right.n193 drain_right.n192 10.2747
R1576 drain_right.n55 drain_right.n40 9.69747
R1577 drain_right.n82 drain_right.n81 9.69747
R1578 drain_right.n102 drain_right.n101 9.69747
R1579 drain_right.n128 drain_right.n4 9.69747
R1580 drain_right.n274 drain_right.n150 9.69747
R1581 drain_right.n249 drain_right.n248 9.69747
R1582 drain_right.n229 drain_right.n228 9.69747
R1583 drain_right.n203 drain_right.n188 9.69747
R1584 drain_right.n138 drain_right.n137 9.45567
R1585 drain_right.n284 drain_right.n283 9.45567
R1586 drain_right.n2 drain_right.n1 9.3005
R1587 drain_right.n131 drain_right.n130 9.3005
R1588 drain_right.n129 drain_right.n128 9.3005
R1589 drain_right.n6 drain_right.n5 9.3005
R1590 drain_right.n123 drain_right.n122 9.3005
R1591 drain_right.n121 drain_right.n120 9.3005
R1592 drain_right.n10 drain_right.n9 9.3005
R1593 drain_right.n89 drain_right.n88 9.3005
R1594 drain_right.n87 drain_right.n86 9.3005
R1595 drain_right.n26 drain_right.n25 9.3005
R1596 drain_right.n81 drain_right.n80 9.3005
R1597 drain_right.n79 drain_right.n78 9.3005
R1598 drain_right.n30 drain_right.n29 9.3005
R1599 drain_right.n73 drain_right.n72 9.3005
R1600 drain_right.n71 drain_right.n70 9.3005
R1601 drain_right.n47 drain_right.n46 9.3005
R1602 drain_right.n42 drain_right.n41 9.3005
R1603 drain_right.n53 drain_right.n52 9.3005
R1604 drain_right.n55 drain_right.n54 9.3005
R1605 drain_right.n38 drain_right.n37 9.3005
R1606 drain_right.n61 drain_right.n60 9.3005
R1607 drain_right.n63 drain_right.n62 9.3005
R1608 drain_right.n64 drain_right.n33 9.3005
R1609 drain_right.n22 drain_right.n21 9.3005
R1610 drain_right.n95 drain_right.n94 9.3005
R1611 drain_right.n97 drain_right.n96 9.3005
R1612 drain_right.n18 drain_right.n17 9.3005
R1613 drain_right.n103 drain_right.n102 9.3005
R1614 drain_right.n105 drain_right.n104 9.3005
R1615 drain_right.n14 drain_right.n13 9.3005
R1616 drain_right.n112 drain_right.n111 9.3005
R1617 drain_right.n114 drain_right.n113 9.3005
R1618 drain_right.n137 drain_right.n136 9.3005
R1619 drain_right.n195 drain_right.n194 9.3005
R1620 drain_right.n190 drain_right.n189 9.3005
R1621 drain_right.n201 drain_right.n200 9.3005
R1622 drain_right.n203 drain_right.n202 9.3005
R1623 drain_right.n186 drain_right.n185 9.3005
R1624 drain_right.n209 drain_right.n208 9.3005
R1625 drain_right.n211 drain_right.n210 9.3005
R1626 drain_right.n183 drain_right.n180 9.3005
R1627 drain_right.n242 drain_right.n241 9.3005
R1628 drain_right.n244 drain_right.n243 9.3005
R1629 drain_right.n165 drain_right.n164 9.3005
R1630 drain_right.n250 drain_right.n249 9.3005
R1631 drain_right.n252 drain_right.n251 9.3005
R1632 drain_right.n160 drain_right.n159 9.3005
R1633 drain_right.n258 drain_right.n257 9.3005
R1634 drain_right.n260 drain_right.n259 9.3005
R1635 drain_right.n283 drain_right.n282 9.3005
R1636 drain_right.n148 drain_right.n147 9.3005
R1637 drain_right.n277 drain_right.n276 9.3005
R1638 drain_right.n275 drain_right.n274 9.3005
R1639 drain_right.n152 drain_right.n151 9.3005
R1640 drain_right.n269 drain_right.n268 9.3005
R1641 drain_right.n267 drain_right.n266 9.3005
R1642 drain_right.n156 drain_right.n155 9.3005
R1643 drain_right.n169 drain_right.n168 9.3005
R1644 drain_right.n236 drain_right.n235 9.3005
R1645 drain_right.n234 drain_right.n233 9.3005
R1646 drain_right.n173 drain_right.n172 9.3005
R1647 drain_right.n228 drain_right.n227 9.3005
R1648 drain_right.n226 drain_right.n225 9.3005
R1649 drain_right.n177 drain_right.n176 9.3005
R1650 drain_right.n220 drain_right.n219 9.3005
R1651 drain_right.n218 drain_right.n217 9.3005
R1652 drain_right.n52 drain_right.n51 8.92171
R1653 drain_right.n85 drain_right.n26 8.92171
R1654 drain_right.n98 drain_right.n18 8.92171
R1655 drain_right.n132 drain_right.n131 8.92171
R1656 drain_right.n278 drain_right.n277 8.92171
R1657 drain_right.n245 drain_right.n165 8.92171
R1658 drain_right.n232 drain_right.n173 8.92171
R1659 drain_right.n200 drain_right.n199 8.92171
R1660 drain_right.n48 drain_right.n42 8.14595
R1661 drain_right.n86 drain_right.n24 8.14595
R1662 drain_right.n97 drain_right.n20 8.14595
R1663 drain_right.n135 drain_right.n2 8.14595
R1664 drain_right.n281 drain_right.n148 8.14595
R1665 drain_right.n244 drain_right.n167 8.14595
R1666 drain_right.n233 drain_right.n171 8.14595
R1667 drain_right.n196 drain_right.n190 8.14595
R1668 drain_right.n47 drain_right.n44 7.3702
R1669 drain_right.n90 drain_right.n89 7.3702
R1670 drain_right.n94 drain_right.n93 7.3702
R1671 drain_right.n136 drain_right.n0 7.3702
R1672 drain_right.n282 drain_right.n146 7.3702
R1673 drain_right.n241 drain_right.n240 7.3702
R1674 drain_right.n237 drain_right.n236 7.3702
R1675 drain_right.n195 drain_right.n192 7.3702
R1676 drain_right.n90 drain_right.n22 6.59444
R1677 drain_right.n93 drain_right.n22 6.59444
R1678 drain_right.n138 drain_right.n0 6.59444
R1679 drain_right.n284 drain_right.n146 6.59444
R1680 drain_right.n240 drain_right.n169 6.59444
R1681 drain_right.n237 drain_right.n169 6.59444
R1682 drain_right drain_right.n285 5.88166
R1683 drain_right.n48 drain_right.n47 5.81868
R1684 drain_right.n89 drain_right.n24 5.81868
R1685 drain_right.n94 drain_right.n20 5.81868
R1686 drain_right.n136 drain_right.n135 5.81868
R1687 drain_right.n282 drain_right.n281 5.81868
R1688 drain_right.n241 drain_right.n167 5.81868
R1689 drain_right.n236 drain_right.n171 5.81868
R1690 drain_right.n196 drain_right.n195 5.81868
R1691 drain_right.n51 drain_right.n42 5.04292
R1692 drain_right.n86 drain_right.n85 5.04292
R1693 drain_right.n98 drain_right.n97 5.04292
R1694 drain_right.n132 drain_right.n2 5.04292
R1695 drain_right.n278 drain_right.n148 5.04292
R1696 drain_right.n245 drain_right.n244 5.04292
R1697 drain_right.n233 drain_right.n232 5.04292
R1698 drain_right.n199 drain_right.n190 5.04292
R1699 drain_right.n52 drain_right.n40 4.26717
R1700 drain_right.n82 drain_right.n26 4.26717
R1701 drain_right.n101 drain_right.n18 4.26717
R1702 drain_right.n131 drain_right.n4 4.26717
R1703 drain_right.n277 drain_right.n150 4.26717
R1704 drain_right.n248 drain_right.n165 4.26717
R1705 drain_right.n229 drain_right.n173 4.26717
R1706 drain_right.n200 drain_right.n188 4.26717
R1707 drain_right.n56 drain_right.n55 3.49141
R1708 drain_right.n81 drain_right.n28 3.49141
R1709 drain_right.n102 drain_right.n16 3.49141
R1710 drain_right.n128 drain_right.n127 3.49141
R1711 drain_right.n274 drain_right.n273 3.49141
R1712 drain_right.n249 drain_right.n163 3.49141
R1713 drain_right.n228 drain_right.n175 3.49141
R1714 drain_right.n204 drain_right.n203 3.49141
R1715 drain_right.n194 drain_right.n193 2.84303
R1716 drain_right.n46 drain_right.n45 2.84303
R1717 drain_right.n59 drain_right.n38 2.71565
R1718 drain_right.n78 drain_right.n77 2.71565
R1719 drain_right.n106 drain_right.n105 2.71565
R1720 drain_right.n124 drain_right.n6 2.71565
R1721 drain_right.n270 drain_right.n152 2.71565
R1722 drain_right.n253 drain_right.n252 2.71565
R1723 drain_right.n225 drain_right.n224 2.71565
R1724 drain_right.n207 drain_right.n186 2.71565
R1725 drain_right.n60 drain_right.n36 1.93989
R1726 drain_right.n74 drain_right.n30 1.93989
R1727 drain_right.n110 drain_right.n14 1.93989
R1728 drain_right.n123 drain_right.n8 1.93989
R1729 drain_right.n269 drain_right.n154 1.93989
R1730 drain_right.n256 drain_right.n160 1.93989
R1731 drain_right.n221 drain_right.n177 1.93989
R1732 drain_right.n208 drain_right.n184 1.93989
R1733 drain_right.n65 drain_right.n63 1.16414
R1734 drain_right.n73 drain_right.n32 1.16414
R1735 drain_right.n111 drain_right.n12 1.16414
R1736 drain_right.n120 drain_right.n119 1.16414
R1737 drain_right.n266 drain_right.n265 1.16414
R1738 drain_right.n257 drain_right.n158 1.16414
R1739 drain_right.n220 drain_right.n179 1.16414
R1740 drain_right.n212 drain_right.n211 1.16414
R1741 drain_right.n141 drain_right.t5 0.7925
R1742 drain_right.n141 drain_right.t3 0.7925
R1743 drain_right.n139 drain_right.t4 0.7925
R1744 drain_right.n139 drain_right.t8 0.7925
R1745 drain_right.n143 drain_right.t6 0.7925
R1746 drain_right.n143 drain_right.t2 0.7925
R1747 drain_right.n144 drain_right.t0 0.7925
R1748 drain_right.n144 drain_right.t9 0.7925
R1749 drain_right.n285 drain_right.n145 0.457397
R1750 drain_right.n64 drain_right.n34 0.388379
R1751 drain_right.n70 drain_right.n69 0.388379
R1752 drain_right.n115 drain_right.n114 0.388379
R1753 drain_right.n116 drain_right.n10 0.388379
R1754 drain_right.n262 drain_right.n156 0.388379
R1755 drain_right.n261 drain_right.n260 0.388379
R1756 drain_right.n217 drain_right.n216 0.388379
R1757 drain_right.n183 drain_right.n181 0.388379
R1758 drain_right.n46 drain_right.n41 0.155672
R1759 drain_right.n53 drain_right.n41 0.155672
R1760 drain_right.n54 drain_right.n53 0.155672
R1761 drain_right.n54 drain_right.n37 0.155672
R1762 drain_right.n61 drain_right.n37 0.155672
R1763 drain_right.n62 drain_right.n61 0.155672
R1764 drain_right.n62 drain_right.n33 0.155672
R1765 drain_right.n71 drain_right.n33 0.155672
R1766 drain_right.n72 drain_right.n71 0.155672
R1767 drain_right.n72 drain_right.n29 0.155672
R1768 drain_right.n79 drain_right.n29 0.155672
R1769 drain_right.n80 drain_right.n79 0.155672
R1770 drain_right.n80 drain_right.n25 0.155672
R1771 drain_right.n87 drain_right.n25 0.155672
R1772 drain_right.n88 drain_right.n87 0.155672
R1773 drain_right.n88 drain_right.n21 0.155672
R1774 drain_right.n95 drain_right.n21 0.155672
R1775 drain_right.n96 drain_right.n95 0.155672
R1776 drain_right.n96 drain_right.n17 0.155672
R1777 drain_right.n103 drain_right.n17 0.155672
R1778 drain_right.n104 drain_right.n103 0.155672
R1779 drain_right.n104 drain_right.n13 0.155672
R1780 drain_right.n112 drain_right.n13 0.155672
R1781 drain_right.n113 drain_right.n112 0.155672
R1782 drain_right.n113 drain_right.n9 0.155672
R1783 drain_right.n121 drain_right.n9 0.155672
R1784 drain_right.n122 drain_right.n121 0.155672
R1785 drain_right.n122 drain_right.n5 0.155672
R1786 drain_right.n129 drain_right.n5 0.155672
R1787 drain_right.n130 drain_right.n129 0.155672
R1788 drain_right.n130 drain_right.n1 0.155672
R1789 drain_right.n137 drain_right.n1 0.155672
R1790 drain_right.n283 drain_right.n147 0.155672
R1791 drain_right.n276 drain_right.n147 0.155672
R1792 drain_right.n276 drain_right.n275 0.155672
R1793 drain_right.n275 drain_right.n151 0.155672
R1794 drain_right.n268 drain_right.n151 0.155672
R1795 drain_right.n268 drain_right.n267 0.155672
R1796 drain_right.n267 drain_right.n155 0.155672
R1797 drain_right.n259 drain_right.n155 0.155672
R1798 drain_right.n259 drain_right.n258 0.155672
R1799 drain_right.n258 drain_right.n159 0.155672
R1800 drain_right.n251 drain_right.n159 0.155672
R1801 drain_right.n251 drain_right.n250 0.155672
R1802 drain_right.n250 drain_right.n164 0.155672
R1803 drain_right.n243 drain_right.n164 0.155672
R1804 drain_right.n243 drain_right.n242 0.155672
R1805 drain_right.n242 drain_right.n168 0.155672
R1806 drain_right.n235 drain_right.n168 0.155672
R1807 drain_right.n235 drain_right.n234 0.155672
R1808 drain_right.n234 drain_right.n172 0.155672
R1809 drain_right.n227 drain_right.n172 0.155672
R1810 drain_right.n227 drain_right.n226 0.155672
R1811 drain_right.n226 drain_right.n176 0.155672
R1812 drain_right.n219 drain_right.n176 0.155672
R1813 drain_right.n219 drain_right.n218 0.155672
R1814 drain_right.n218 drain_right.n180 0.155672
R1815 drain_right.n210 drain_right.n180 0.155672
R1816 drain_right.n210 drain_right.n209 0.155672
R1817 drain_right.n209 drain_right.n185 0.155672
R1818 drain_right.n202 drain_right.n185 0.155672
R1819 drain_right.n202 drain_right.n201 0.155672
R1820 drain_right.n201 drain_right.n189 0.155672
R1821 drain_right.n194 drain_right.n189 0.155672
R1822 drain_right.n142 drain_right.n140 0.0593781
C0 drain_right source 49.6435f
C1 drain_left minus 0.170748f
C2 minus plus 7.24796f
C3 minus source 4.95088f
C4 drain_right minus 5.99873f
C5 drain_left plus 6.12049f
C6 drain_left source 49.6672f
C7 drain_right drain_left 0.66859f
C8 source plus 4.96638f
C9 drain_right plus 0.286116f
C10 drain_right a_n1352_n5888# 11.114849f
C11 drain_left a_n1352_n5888# 11.33943f
C12 source a_n1352_n5888# 10.408701f
C13 minus a_n1352_n5888# 6.089818f
C14 plus a_n1352_n5888# 9.16081f
C15 drain_right.n0 a_n1352_n5888# 0.046548f
C16 drain_right.n1 a_n1352_n5888# 0.033764f
C17 drain_right.n2 a_n1352_n5888# 0.018143f
C18 drain_right.n3 a_n1352_n5888# 0.042885f
C19 drain_right.n4 a_n1352_n5888# 0.019211f
C20 drain_right.n5 a_n1352_n5888# 0.033764f
C21 drain_right.n6 a_n1352_n5888# 0.018143f
C22 drain_right.n7 a_n1352_n5888# 0.042885f
C23 drain_right.n8 a_n1352_n5888# 0.019211f
C24 drain_right.n9 a_n1352_n5888# 0.033764f
C25 drain_right.n10 a_n1352_n5888# 0.018143f
C26 drain_right.n11 a_n1352_n5888# 0.042885f
C27 drain_right.n12 a_n1352_n5888# 0.019211f
C28 drain_right.n13 a_n1352_n5888# 0.033764f
C29 drain_right.n14 a_n1352_n5888# 0.018143f
C30 drain_right.n15 a_n1352_n5888# 0.042885f
C31 drain_right.n16 a_n1352_n5888# 0.019211f
C32 drain_right.n17 a_n1352_n5888# 0.033764f
C33 drain_right.n18 a_n1352_n5888# 0.018143f
C34 drain_right.n19 a_n1352_n5888# 0.042885f
C35 drain_right.n20 a_n1352_n5888# 0.019211f
C36 drain_right.n21 a_n1352_n5888# 0.033764f
C37 drain_right.n22 a_n1352_n5888# 0.018143f
C38 drain_right.n23 a_n1352_n5888# 0.042885f
C39 drain_right.n24 a_n1352_n5888# 0.019211f
C40 drain_right.n25 a_n1352_n5888# 0.033764f
C41 drain_right.n26 a_n1352_n5888# 0.018143f
C42 drain_right.n27 a_n1352_n5888# 0.042885f
C43 drain_right.n28 a_n1352_n5888# 0.019211f
C44 drain_right.n29 a_n1352_n5888# 0.033764f
C45 drain_right.n30 a_n1352_n5888# 0.018143f
C46 drain_right.n31 a_n1352_n5888# 0.042885f
C47 drain_right.n32 a_n1352_n5888# 0.019211f
C48 drain_right.n33 a_n1352_n5888# 0.033764f
C49 drain_right.n34 a_n1352_n5888# 0.018677f
C50 drain_right.n35 a_n1352_n5888# 0.042885f
C51 drain_right.n36 a_n1352_n5888# 0.019211f
C52 drain_right.n37 a_n1352_n5888# 0.033764f
C53 drain_right.n38 a_n1352_n5888# 0.018143f
C54 drain_right.n39 a_n1352_n5888# 0.042885f
C55 drain_right.n40 a_n1352_n5888# 0.019211f
C56 drain_right.n41 a_n1352_n5888# 0.033764f
C57 drain_right.n42 a_n1352_n5888# 0.018143f
C58 drain_right.n43 a_n1352_n5888# 0.032164f
C59 drain_right.n44 a_n1352_n5888# 0.030316f
C60 drain_right.t7 a_n1352_n5888# 0.074794f
C61 drain_right.n45 a_n1352_n5888# 0.411954f
C62 drain_right.n46 a_n1352_n5888# 3.65569f
C63 drain_right.n47 a_n1352_n5888# 0.018143f
C64 drain_right.n48 a_n1352_n5888# 0.019211f
C65 drain_right.n49 a_n1352_n5888# 0.042885f
C66 drain_right.n50 a_n1352_n5888# 0.042885f
C67 drain_right.n51 a_n1352_n5888# 0.019211f
C68 drain_right.n52 a_n1352_n5888# 0.018143f
C69 drain_right.n53 a_n1352_n5888# 0.033764f
C70 drain_right.n54 a_n1352_n5888# 0.033764f
C71 drain_right.n55 a_n1352_n5888# 0.018143f
C72 drain_right.n56 a_n1352_n5888# 0.019211f
C73 drain_right.n57 a_n1352_n5888# 0.042885f
C74 drain_right.n58 a_n1352_n5888# 0.042885f
C75 drain_right.n59 a_n1352_n5888# 0.019211f
C76 drain_right.n60 a_n1352_n5888# 0.018143f
C77 drain_right.n61 a_n1352_n5888# 0.033764f
C78 drain_right.n62 a_n1352_n5888# 0.033764f
C79 drain_right.n63 a_n1352_n5888# 0.018143f
C80 drain_right.n64 a_n1352_n5888# 0.018143f
C81 drain_right.n65 a_n1352_n5888# 0.019211f
C82 drain_right.n66 a_n1352_n5888# 0.042885f
C83 drain_right.n67 a_n1352_n5888# 0.042885f
C84 drain_right.n68 a_n1352_n5888# 0.042885f
C85 drain_right.n69 a_n1352_n5888# 0.018677f
C86 drain_right.n70 a_n1352_n5888# 0.018143f
C87 drain_right.n71 a_n1352_n5888# 0.033764f
C88 drain_right.n72 a_n1352_n5888# 0.033764f
C89 drain_right.n73 a_n1352_n5888# 0.018143f
C90 drain_right.n74 a_n1352_n5888# 0.019211f
C91 drain_right.n75 a_n1352_n5888# 0.042885f
C92 drain_right.n76 a_n1352_n5888# 0.042885f
C93 drain_right.n77 a_n1352_n5888# 0.019211f
C94 drain_right.n78 a_n1352_n5888# 0.018143f
C95 drain_right.n79 a_n1352_n5888# 0.033764f
C96 drain_right.n80 a_n1352_n5888# 0.033764f
C97 drain_right.n81 a_n1352_n5888# 0.018143f
C98 drain_right.n82 a_n1352_n5888# 0.019211f
C99 drain_right.n83 a_n1352_n5888# 0.042885f
C100 drain_right.n84 a_n1352_n5888# 0.042885f
C101 drain_right.n85 a_n1352_n5888# 0.019211f
C102 drain_right.n86 a_n1352_n5888# 0.018143f
C103 drain_right.n87 a_n1352_n5888# 0.033764f
C104 drain_right.n88 a_n1352_n5888# 0.033764f
C105 drain_right.n89 a_n1352_n5888# 0.018143f
C106 drain_right.n90 a_n1352_n5888# 0.019211f
C107 drain_right.n91 a_n1352_n5888# 0.042885f
C108 drain_right.n92 a_n1352_n5888# 0.042885f
C109 drain_right.n93 a_n1352_n5888# 0.019211f
C110 drain_right.n94 a_n1352_n5888# 0.018143f
C111 drain_right.n95 a_n1352_n5888# 0.033764f
C112 drain_right.n96 a_n1352_n5888# 0.033764f
C113 drain_right.n97 a_n1352_n5888# 0.018143f
C114 drain_right.n98 a_n1352_n5888# 0.019211f
C115 drain_right.n99 a_n1352_n5888# 0.042885f
C116 drain_right.n100 a_n1352_n5888# 0.042885f
C117 drain_right.n101 a_n1352_n5888# 0.019211f
C118 drain_right.n102 a_n1352_n5888# 0.018143f
C119 drain_right.n103 a_n1352_n5888# 0.033764f
C120 drain_right.n104 a_n1352_n5888# 0.033764f
C121 drain_right.n105 a_n1352_n5888# 0.018143f
C122 drain_right.n106 a_n1352_n5888# 0.019211f
C123 drain_right.n107 a_n1352_n5888# 0.042885f
C124 drain_right.n108 a_n1352_n5888# 0.042885f
C125 drain_right.n109 a_n1352_n5888# 0.042885f
C126 drain_right.n110 a_n1352_n5888# 0.019211f
C127 drain_right.n111 a_n1352_n5888# 0.018143f
C128 drain_right.n112 a_n1352_n5888# 0.033764f
C129 drain_right.n113 a_n1352_n5888# 0.033764f
C130 drain_right.n114 a_n1352_n5888# 0.018143f
C131 drain_right.n115 a_n1352_n5888# 0.018677f
C132 drain_right.n116 a_n1352_n5888# 0.018677f
C133 drain_right.n117 a_n1352_n5888# 0.042885f
C134 drain_right.n118 a_n1352_n5888# 0.042885f
C135 drain_right.n119 a_n1352_n5888# 0.019211f
C136 drain_right.n120 a_n1352_n5888# 0.018143f
C137 drain_right.n121 a_n1352_n5888# 0.033764f
C138 drain_right.n122 a_n1352_n5888# 0.033764f
C139 drain_right.n123 a_n1352_n5888# 0.018143f
C140 drain_right.n124 a_n1352_n5888# 0.019211f
C141 drain_right.n125 a_n1352_n5888# 0.042885f
C142 drain_right.n126 a_n1352_n5888# 0.042885f
C143 drain_right.n127 a_n1352_n5888# 0.019211f
C144 drain_right.n128 a_n1352_n5888# 0.018143f
C145 drain_right.n129 a_n1352_n5888# 0.033764f
C146 drain_right.n130 a_n1352_n5888# 0.033764f
C147 drain_right.n131 a_n1352_n5888# 0.018143f
C148 drain_right.n132 a_n1352_n5888# 0.019211f
C149 drain_right.n133 a_n1352_n5888# 0.042885f
C150 drain_right.n134 a_n1352_n5888# 0.091227f
C151 drain_right.n135 a_n1352_n5888# 0.019211f
C152 drain_right.n136 a_n1352_n5888# 0.018143f
C153 drain_right.n137 a_n1352_n5888# 0.074355f
C154 drain_right.n138 a_n1352_n5888# 0.075185f
C155 drain_right.t4 a_n1352_n5888# 0.667041f
C156 drain_right.t8 a_n1352_n5888# 0.667041f
C157 drain_right.n139 a_n1352_n5888# 6.1475f
C158 drain_right.n140 a_n1352_n5888# 0.466352f
C159 drain_right.t5 a_n1352_n5888# 0.667041f
C160 drain_right.t3 a_n1352_n5888# 0.667041f
C161 drain_right.n141 a_n1352_n5888# 6.14937f
C162 drain_right.n142 a_n1352_n5888# 2.88316f
C163 drain_right.t6 a_n1352_n5888# 0.667041f
C164 drain_right.t2 a_n1352_n5888# 0.667041f
C165 drain_right.n143 a_n1352_n5888# 6.15056f
C166 drain_right.t0 a_n1352_n5888# 0.667041f
C167 drain_right.t9 a_n1352_n5888# 0.667041f
C168 drain_right.n144 a_n1352_n5888# 6.1475f
C169 drain_right.n145 a_n1352_n5888# 0.780184f
C170 drain_right.n146 a_n1352_n5888# 0.046548f
C171 drain_right.n147 a_n1352_n5888# 0.033764f
C172 drain_right.n148 a_n1352_n5888# 0.018143f
C173 drain_right.n149 a_n1352_n5888# 0.042885f
C174 drain_right.n150 a_n1352_n5888# 0.019211f
C175 drain_right.n151 a_n1352_n5888# 0.033764f
C176 drain_right.n152 a_n1352_n5888# 0.018143f
C177 drain_right.n153 a_n1352_n5888# 0.042885f
C178 drain_right.n154 a_n1352_n5888# 0.019211f
C179 drain_right.n155 a_n1352_n5888# 0.033764f
C180 drain_right.n156 a_n1352_n5888# 0.018143f
C181 drain_right.n157 a_n1352_n5888# 0.042885f
C182 drain_right.n158 a_n1352_n5888# 0.019211f
C183 drain_right.n159 a_n1352_n5888# 0.033764f
C184 drain_right.n160 a_n1352_n5888# 0.018143f
C185 drain_right.n161 a_n1352_n5888# 0.042885f
C186 drain_right.n162 a_n1352_n5888# 0.042885f
C187 drain_right.n163 a_n1352_n5888# 0.019211f
C188 drain_right.n164 a_n1352_n5888# 0.033764f
C189 drain_right.n165 a_n1352_n5888# 0.018143f
C190 drain_right.n166 a_n1352_n5888# 0.042885f
C191 drain_right.n167 a_n1352_n5888# 0.019211f
C192 drain_right.n168 a_n1352_n5888# 0.033764f
C193 drain_right.n169 a_n1352_n5888# 0.018143f
C194 drain_right.n170 a_n1352_n5888# 0.042885f
C195 drain_right.n171 a_n1352_n5888# 0.019211f
C196 drain_right.n172 a_n1352_n5888# 0.033764f
C197 drain_right.n173 a_n1352_n5888# 0.018143f
C198 drain_right.n174 a_n1352_n5888# 0.042885f
C199 drain_right.n175 a_n1352_n5888# 0.019211f
C200 drain_right.n176 a_n1352_n5888# 0.033764f
C201 drain_right.n177 a_n1352_n5888# 0.018143f
C202 drain_right.n178 a_n1352_n5888# 0.042885f
C203 drain_right.n179 a_n1352_n5888# 0.019211f
C204 drain_right.n180 a_n1352_n5888# 0.033764f
C205 drain_right.n181 a_n1352_n5888# 0.018677f
C206 drain_right.n182 a_n1352_n5888# 0.042885f
C207 drain_right.n183 a_n1352_n5888# 0.018143f
C208 drain_right.n184 a_n1352_n5888# 0.019211f
C209 drain_right.n185 a_n1352_n5888# 0.033764f
C210 drain_right.n186 a_n1352_n5888# 0.018143f
C211 drain_right.n187 a_n1352_n5888# 0.042885f
C212 drain_right.n188 a_n1352_n5888# 0.019211f
C213 drain_right.n189 a_n1352_n5888# 0.033764f
C214 drain_right.n190 a_n1352_n5888# 0.018143f
C215 drain_right.n191 a_n1352_n5888# 0.032164f
C216 drain_right.n192 a_n1352_n5888# 0.030316f
C217 drain_right.t1 a_n1352_n5888# 0.074794f
C218 drain_right.n193 a_n1352_n5888# 0.411954f
C219 drain_right.n194 a_n1352_n5888# 3.65569f
C220 drain_right.n195 a_n1352_n5888# 0.018143f
C221 drain_right.n196 a_n1352_n5888# 0.019211f
C222 drain_right.n197 a_n1352_n5888# 0.042885f
C223 drain_right.n198 a_n1352_n5888# 0.042885f
C224 drain_right.n199 a_n1352_n5888# 0.019211f
C225 drain_right.n200 a_n1352_n5888# 0.018143f
C226 drain_right.n201 a_n1352_n5888# 0.033764f
C227 drain_right.n202 a_n1352_n5888# 0.033764f
C228 drain_right.n203 a_n1352_n5888# 0.018143f
C229 drain_right.n204 a_n1352_n5888# 0.019211f
C230 drain_right.n205 a_n1352_n5888# 0.042885f
C231 drain_right.n206 a_n1352_n5888# 0.042885f
C232 drain_right.n207 a_n1352_n5888# 0.019211f
C233 drain_right.n208 a_n1352_n5888# 0.018143f
C234 drain_right.n209 a_n1352_n5888# 0.033764f
C235 drain_right.n210 a_n1352_n5888# 0.033764f
C236 drain_right.n211 a_n1352_n5888# 0.018143f
C237 drain_right.n212 a_n1352_n5888# 0.019211f
C238 drain_right.n213 a_n1352_n5888# 0.042885f
C239 drain_right.n214 a_n1352_n5888# 0.042885f
C240 drain_right.n215 a_n1352_n5888# 0.042885f
C241 drain_right.n216 a_n1352_n5888# 0.018677f
C242 drain_right.n217 a_n1352_n5888# 0.018143f
C243 drain_right.n218 a_n1352_n5888# 0.033764f
C244 drain_right.n219 a_n1352_n5888# 0.033764f
C245 drain_right.n220 a_n1352_n5888# 0.018143f
C246 drain_right.n221 a_n1352_n5888# 0.019211f
C247 drain_right.n222 a_n1352_n5888# 0.042885f
C248 drain_right.n223 a_n1352_n5888# 0.042885f
C249 drain_right.n224 a_n1352_n5888# 0.019211f
C250 drain_right.n225 a_n1352_n5888# 0.018143f
C251 drain_right.n226 a_n1352_n5888# 0.033764f
C252 drain_right.n227 a_n1352_n5888# 0.033764f
C253 drain_right.n228 a_n1352_n5888# 0.018143f
C254 drain_right.n229 a_n1352_n5888# 0.019211f
C255 drain_right.n230 a_n1352_n5888# 0.042885f
C256 drain_right.n231 a_n1352_n5888# 0.042885f
C257 drain_right.n232 a_n1352_n5888# 0.019211f
C258 drain_right.n233 a_n1352_n5888# 0.018143f
C259 drain_right.n234 a_n1352_n5888# 0.033764f
C260 drain_right.n235 a_n1352_n5888# 0.033764f
C261 drain_right.n236 a_n1352_n5888# 0.018143f
C262 drain_right.n237 a_n1352_n5888# 0.019211f
C263 drain_right.n238 a_n1352_n5888# 0.042885f
C264 drain_right.n239 a_n1352_n5888# 0.042885f
C265 drain_right.n240 a_n1352_n5888# 0.019211f
C266 drain_right.n241 a_n1352_n5888# 0.018143f
C267 drain_right.n242 a_n1352_n5888# 0.033764f
C268 drain_right.n243 a_n1352_n5888# 0.033764f
C269 drain_right.n244 a_n1352_n5888# 0.018143f
C270 drain_right.n245 a_n1352_n5888# 0.019211f
C271 drain_right.n246 a_n1352_n5888# 0.042885f
C272 drain_right.n247 a_n1352_n5888# 0.042885f
C273 drain_right.n248 a_n1352_n5888# 0.019211f
C274 drain_right.n249 a_n1352_n5888# 0.018143f
C275 drain_right.n250 a_n1352_n5888# 0.033764f
C276 drain_right.n251 a_n1352_n5888# 0.033764f
C277 drain_right.n252 a_n1352_n5888# 0.018143f
C278 drain_right.n253 a_n1352_n5888# 0.019211f
C279 drain_right.n254 a_n1352_n5888# 0.042885f
C280 drain_right.n255 a_n1352_n5888# 0.042885f
C281 drain_right.n256 a_n1352_n5888# 0.019211f
C282 drain_right.n257 a_n1352_n5888# 0.018143f
C283 drain_right.n258 a_n1352_n5888# 0.033764f
C284 drain_right.n259 a_n1352_n5888# 0.033764f
C285 drain_right.n260 a_n1352_n5888# 0.018143f
C286 drain_right.n261 a_n1352_n5888# 0.018677f
C287 drain_right.n262 a_n1352_n5888# 0.018677f
C288 drain_right.n263 a_n1352_n5888# 0.042885f
C289 drain_right.n264 a_n1352_n5888# 0.042885f
C290 drain_right.n265 a_n1352_n5888# 0.019211f
C291 drain_right.n266 a_n1352_n5888# 0.018143f
C292 drain_right.n267 a_n1352_n5888# 0.033764f
C293 drain_right.n268 a_n1352_n5888# 0.033764f
C294 drain_right.n269 a_n1352_n5888# 0.018143f
C295 drain_right.n270 a_n1352_n5888# 0.019211f
C296 drain_right.n271 a_n1352_n5888# 0.042885f
C297 drain_right.n272 a_n1352_n5888# 0.042885f
C298 drain_right.n273 a_n1352_n5888# 0.019211f
C299 drain_right.n274 a_n1352_n5888# 0.018143f
C300 drain_right.n275 a_n1352_n5888# 0.033764f
C301 drain_right.n276 a_n1352_n5888# 0.033764f
C302 drain_right.n277 a_n1352_n5888# 0.018143f
C303 drain_right.n278 a_n1352_n5888# 0.019211f
C304 drain_right.n279 a_n1352_n5888# 0.042885f
C305 drain_right.n280 a_n1352_n5888# 0.091227f
C306 drain_right.n281 a_n1352_n5888# 0.019211f
C307 drain_right.n282 a_n1352_n5888# 0.018143f
C308 drain_right.n283 a_n1352_n5888# 0.074355f
C309 drain_right.n284 a_n1352_n5888# 0.074108f
C310 drain_right.n285 a_n1352_n5888# 0.387042f
C311 minus.n0 a_n1352_n5888# 0.058153f
C312 minus.t8 a_n1352_n5888# 0.822402f
C313 minus.t9 a_n1352_n5888# 0.81812f
C314 minus.t0 a_n1352_n5888# 0.81812f
C315 minus.t3 a_n1352_n5888# 0.81812f
C316 minus.n1 a_n1352_n5888# 0.303671f
C317 minus.t7 a_n1352_n5888# 0.822402f
C318 minus.n2 a_n1352_n5888# 0.320196f
C319 minus.n3 a_n1352_n5888# 0.127698f
C320 minus.n4 a_n1352_n5888# 0.020367f
C321 minus.n5 a_n1352_n5888# 0.303671f
C322 minus.n6 a_n1352_n5888# 0.020367f
C323 minus.n7 a_n1352_n5888# 0.303671f
C324 minus.n8 a_n1352_n5888# 0.320114f
C325 minus.n9 a_n1352_n5888# 2.75816f
C326 minus.n10 a_n1352_n5888# 0.058153f
C327 minus.t4 a_n1352_n5888# 0.81812f
C328 minus.t1 a_n1352_n5888# 0.81812f
C329 minus.t5 a_n1352_n5888# 0.81812f
C330 minus.n11 a_n1352_n5888# 0.303671f
C331 minus.t2 a_n1352_n5888# 0.822402f
C332 minus.n12 a_n1352_n5888# 0.320196f
C333 minus.n13 a_n1352_n5888# 0.127698f
C334 minus.n14 a_n1352_n5888# 0.020367f
C335 minus.n15 a_n1352_n5888# 0.303671f
C336 minus.n16 a_n1352_n5888# 0.020367f
C337 minus.n17 a_n1352_n5888# 0.303671f
C338 minus.t6 a_n1352_n5888# 0.822402f
C339 minus.n18 a_n1352_n5888# 0.320114f
C340 minus.n19 a_n1352_n5888# 0.373236f
C341 minus.n20 a_n1352_n5888# 3.27627f
C342 source.n0 a_n1352_n5888# 0.046845f
C343 source.n1 a_n1352_n5888# 0.03398f
C344 source.n2 a_n1352_n5888# 0.01826f
C345 source.n3 a_n1352_n5888# 0.043159f
C346 source.n4 a_n1352_n5888# 0.019334f
C347 source.n5 a_n1352_n5888# 0.03398f
C348 source.n6 a_n1352_n5888# 0.01826f
C349 source.n7 a_n1352_n5888# 0.043159f
C350 source.n8 a_n1352_n5888# 0.019334f
C351 source.n9 a_n1352_n5888# 0.03398f
C352 source.n10 a_n1352_n5888# 0.01826f
C353 source.n11 a_n1352_n5888# 0.043159f
C354 source.n12 a_n1352_n5888# 0.019334f
C355 source.n13 a_n1352_n5888# 0.03398f
C356 source.n14 a_n1352_n5888# 0.01826f
C357 source.n15 a_n1352_n5888# 0.043159f
C358 source.n16 a_n1352_n5888# 0.043159f
C359 source.n17 a_n1352_n5888# 0.019334f
C360 source.n18 a_n1352_n5888# 0.03398f
C361 source.n19 a_n1352_n5888# 0.01826f
C362 source.n20 a_n1352_n5888# 0.043159f
C363 source.n21 a_n1352_n5888# 0.019334f
C364 source.n22 a_n1352_n5888# 0.03398f
C365 source.n23 a_n1352_n5888# 0.01826f
C366 source.n24 a_n1352_n5888# 0.043159f
C367 source.n25 a_n1352_n5888# 0.019334f
C368 source.n26 a_n1352_n5888# 0.03398f
C369 source.n27 a_n1352_n5888# 0.01826f
C370 source.n28 a_n1352_n5888# 0.043159f
C371 source.n29 a_n1352_n5888# 0.019334f
C372 source.n30 a_n1352_n5888# 0.03398f
C373 source.n31 a_n1352_n5888# 0.01826f
C374 source.n32 a_n1352_n5888# 0.043159f
C375 source.n33 a_n1352_n5888# 0.019334f
C376 source.n34 a_n1352_n5888# 0.03398f
C377 source.n35 a_n1352_n5888# 0.018797f
C378 source.n36 a_n1352_n5888# 0.043159f
C379 source.n37 a_n1352_n5888# 0.01826f
C380 source.n38 a_n1352_n5888# 0.019334f
C381 source.n39 a_n1352_n5888# 0.03398f
C382 source.n40 a_n1352_n5888# 0.01826f
C383 source.n41 a_n1352_n5888# 0.043159f
C384 source.n42 a_n1352_n5888# 0.019334f
C385 source.n43 a_n1352_n5888# 0.03398f
C386 source.n44 a_n1352_n5888# 0.01826f
C387 source.n45 a_n1352_n5888# 0.032369f
C388 source.n46 a_n1352_n5888# 0.03051f
C389 source.t16 a_n1352_n5888# 0.075272f
C390 source.n47 a_n1352_n5888# 0.414589f
C391 source.n48 a_n1352_n5888# 3.67907f
C392 source.n49 a_n1352_n5888# 0.01826f
C393 source.n50 a_n1352_n5888# 0.019334f
C394 source.n51 a_n1352_n5888# 0.043159f
C395 source.n52 a_n1352_n5888# 0.043159f
C396 source.n53 a_n1352_n5888# 0.019334f
C397 source.n54 a_n1352_n5888# 0.01826f
C398 source.n55 a_n1352_n5888# 0.03398f
C399 source.n56 a_n1352_n5888# 0.03398f
C400 source.n57 a_n1352_n5888# 0.01826f
C401 source.n58 a_n1352_n5888# 0.019334f
C402 source.n59 a_n1352_n5888# 0.043159f
C403 source.n60 a_n1352_n5888# 0.043159f
C404 source.n61 a_n1352_n5888# 0.019334f
C405 source.n62 a_n1352_n5888# 0.01826f
C406 source.n63 a_n1352_n5888# 0.03398f
C407 source.n64 a_n1352_n5888# 0.03398f
C408 source.n65 a_n1352_n5888# 0.01826f
C409 source.n66 a_n1352_n5888# 0.019334f
C410 source.n67 a_n1352_n5888# 0.043159f
C411 source.n68 a_n1352_n5888# 0.043159f
C412 source.n69 a_n1352_n5888# 0.043159f
C413 source.n70 a_n1352_n5888# 0.018797f
C414 source.n71 a_n1352_n5888# 0.01826f
C415 source.n72 a_n1352_n5888# 0.03398f
C416 source.n73 a_n1352_n5888# 0.03398f
C417 source.n74 a_n1352_n5888# 0.01826f
C418 source.n75 a_n1352_n5888# 0.019334f
C419 source.n76 a_n1352_n5888# 0.043159f
C420 source.n77 a_n1352_n5888# 0.043159f
C421 source.n78 a_n1352_n5888# 0.019334f
C422 source.n79 a_n1352_n5888# 0.01826f
C423 source.n80 a_n1352_n5888# 0.03398f
C424 source.n81 a_n1352_n5888# 0.03398f
C425 source.n82 a_n1352_n5888# 0.01826f
C426 source.n83 a_n1352_n5888# 0.019334f
C427 source.n84 a_n1352_n5888# 0.043159f
C428 source.n85 a_n1352_n5888# 0.043159f
C429 source.n86 a_n1352_n5888# 0.019334f
C430 source.n87 a_n1352_n5888# 0.01826f
C431 source.n88 a_n1352_n5888# 0.03398f
C432 source.n89 a_n1352_n5888# 0.03398f
C433 source.n90 a_n1352_n5888# 0.01826f
C434 source.n91 a_n1352_n5888# 0.019334f
C435 source.n92 a_n1352_n5888# 0.043159f
C436 source.n93 a_n1352_n5888# 0.043159f
C437 source.n94 a_n1352_n5888# 0.019334f
C438 source.n95 a_n1352_n5888# 0.01826f
C439 source.n96 a_n1352_n5888# 0.03398f
C440 source.n97 a_n1352_n5888# 0.03398f
C441 source.n98 a_n1352_n5888# 0.01826f
C442 source.n99 a_n1352_n5888# 0.019334f
C443 source.n100 a_n1352_n5888# 0.043159f
C444 source.n101 a_n1352_n5888# 0.043159f
C445 source.n102 a_n1352_n5888# 0.019334f
C446 source.n103 a_n1352_n5888# 0.01826f
C447 source.n104 a_n1352_n5888# 0.03398f
C448 source.n105 a_n1352_n5888# 0.03398f
C449 source.n106 a_n1352_n5888# 0.01826f
C450 source.n107 a_n1352_n5888# 0.019334f
C451 source.n108 a_n1352_n5888# 0.043159f
C452 source.n109 a_n1352_n5888# 0.043159f
C453 source.n110 a_n1352_n5888# 0.019334f
C454 source.n111 a_n1352_n5888# 0.01826f
C455 source.n112 a_n1352_n5888# 0.03398f
C456 source.n113 a_n1352_n5888# 0.03398f
C457 source.n114 a_n1352_n5888# 0.01826f
C458 source.n115 a_n1352_n5888# 0.018797f
C459 source.n116 a_n1352_n5888# 0.018797f
C460 source.n117 a_n1352_n5888# 0.043159f
C461 source.n118 a_n1352_n5888# 0.043159f
C462 source.n119 a_n1352_n5888# 0.019334f
C463 source.n120 a_n1352_n5888# 0.01826f
C464 source.n121 a_n1352_n5888# 0.03398f
C465 source.n122 a_n1352_n5888# 0.03398f
C466 source.n123 a_n1352_n5888# 0.01826f
C467 source.n124 a_n1352_n5888# 0.019334f
C468 source.n125 a_n1352_n5888# 0.043159f
C469 source.n126 a_n1352_n5888# 0.043159f
C470 source.n127 a_n1352_n5888# 0.019334f
C471 source.n128 a_n1352_n5888# 0.01826f
C472 source.n129 a_n1352_n5888# 0.03398f
C473 source.n130 a_n1352_n5888# 0.03398f
C474 source.n131 a_n1352_n5888# 0.01826f
C475 source.n132 a_n1352_n5888# 0.019334f
C476 source.n133 a_n1352_n5888# 0.043159f
C477 source.n134 a_n1352_n5888# 0.09181f
C478 source.n135 a_n1352_n5888# 0.019334f
C479 source.n136 a_n1352_n5888# 0.01826f
C480 source.n137 a_n1352_n5888# 0.07483f
C481 source.n138 a_n1352_n5888# 0.051088f
C482 source.n139 a_n1352_n5888# 2.65597f
C483 source.t12 a_n1352_n5888# 0.671308f
C484 source.t15 a_n1352_n5888# 0.671308f
C485 source.n140 a_n1352_n5888# 6.07543f
C486 source.n141 a_n1352_n5888# 0.452497f
C487 source.t17 a_n1352_n5888# 0.671308f
C488 source.t18 a_n1352_n5888# 0.671308f
C489 source.n142 a_n1352_n5888# 6.07543f
C490 source.n143 a_n1352_n5888# 0.478926f
C491 source.n144 a_n1352_n5888# 0.046845f
C492 source.n145 a_n1352_n5888# 0.03398f
C493 source.n146 a_n1352_n5888# 0.01826f
C494 source.n147 a_n1352_n5888# 0.043159f
C495 source.n148 a_n1352_n5888# 0.019334f
C496 source.n149 a_n1352_n5888# 0.03398f
C497 source.n150 a_n1352_n5888# 0.01826f
C498 source.n151 a_n1352_n5888# 0.043159f
C499 source.n152 a_n1352_n5888# 0.019334f
C500 source.n153 a_n1352_n5888# 0.03398f
C501 source.n154 a_n1352_n5888# 0.01826f
C502 source.n155 a_n1352_n5888# 0.043159f
C503 source.n156 a_n1352_n5888# 0.019334f
C504 source.n157 a_n1352_n5888# 0.03398f
C505 source.n158 a_n1352_n5888# 0.01826f
C506 source.n159 a_n1352_n5888# 0.043159f
C507 source.n160 a_n1352_n5888# 0.043159f
C508 source.n161 a_n1352_n5888# 0.019334f
C509 source.n162 a_n1352_n5888# 0.03398f
C510 source.n163 a_n1352_n5888# 0.01826f
C511 source.n164 a_n1352_n5888# 0.043159f
C512 source.n165 a_n1352_n5888# 0.019334f
C513 source.n166 a_n1352_n5888# 0.03398f
C514 source.n167 a_n1352_n5888# 0.01826f
C515 source.n168 a_n1352_n5888# 0.043159f
C516 source.n169 a_n1352_n5888# 0.019334f
C517 source.n170 a_n1352_n5888# 0.03398f
C518 source.n171 a_n1352_n5888# 0.01826f
C519 source.n172 a_n1352_n5888# 0.043159f
C520 source.n173 a_n1352_n5888# 0.019334f
C521 source.n174 a_n1352_n5888# 0.03398f
C522 source.n175 a_n1352_n5888# 0.01826f
C523 source.n176 a_n1352_n5888# 0.043159f
C524 source.n177 a_n1352_n5888# 0.019334f
C525 source.n178 a_n1352_n5888# 0.03398f
C526 source.n179 a_n1352_n5888# 0.018797f
C527 source.n180 a_n1352_n5888# 0.043159f
C528 source.n181 a_n1352_n5888# 0.01826f
C529 source.n182 a_n1352_n5888# 0.019334f
C530 source.n183 a_n1352_n5888# 0.03398f
C531 source.n184 a_n1352_n5888# 0.01826f
C532 source.n185 a_n1352_n5888# 0.043159f
C533 source.n186 a_n1352_n5888# 0.019334f
C534 source.n187 a_n1352_n5888# 0.03398f
C535 source.n188 a_n1352_n5888# 0.01826f
C536 source.n189 a_n1352_n5888# 0.032369f
C537 source.n190 a_n1352_n5888# 0.03051f
C538 source.t7 a_n1352_n5888# 0.075272f
C539 source.n191 a_n1352_n5888# 0.414589f
C540 source.n192 a_n1352_n5888# 3.67907f
C541 source.n193 a_n1352_n5888# 0.01826f
C542 source.n194 a_n1352_n5888# 0.019334f
C543 source.n195 a_n1352_n5888# 0.043159f
C544 source.n196 a_n1352_n5888# 0.043159f
C545 source.n197 a_n1352_n5888# 0.019334f
C546 source.n198 a_n1352_n5888# 0.01826f
C547 source.n199 a_n1352_n5888# 0.03398f
C548 source.n200 a_n1352_n5888# 0.03398f
C549 source.n201 a_n1352_n5888# 0.01826f
C550 source.n202 a_n1352_n5888# 0.019334f
C551 source.n203 a_n1352_n5888# 0.043159f
C552 source.n204 a_n1352_n5888# 0.043159f
C553 source.n205 a_n1352_n5888# 0.019334f
C554 source.n206 a_n1352_n5888# 0.01826f
C555 source.n207 a_n1352_n5888# 0.03398f
C556 source.n208 a_n1352_n5888# 0.03398f
C557 source.n209 a_n1352_n5888# 0.01826f
C558 source.n210 a_n1352_n5888# 0.019334f
C559 source.n211 a_n1352_n5888# 0.043159f
C560 source.n212 a_n1352_n5888# 0.043159f
C561 source.n213 a_n1352_n5888# 0.043159f
C562 source.n214 a_n1352_n5888# 0.018797f
C563 source.n215 a_n1352_n5888# 0.01826f
C564 source.n216 a_n1352_n5888# 0.03398f
C565 source.n217 a_n1352_n5888# 0.03398f
C566 source.n218 a_n1352_n5888# 0.01826f
C567 source.n219 a_n1352_n5888# 0.019334f
C568 source.n220 a_n1352_n5888# 0.043159f
C569 source.n221 a_n1352_n5888# 0.043159f
C570 source.n222 a_n1352_n5888# 0.019334f
C571 source.n223 a_n1352_n5888# 0.01826f
C572 source.n224 a_n1352_n5888# 0.03398f
C573 source.n225 a_n1352_n5888# 0.03398f
C574 source.n226 a_n1352_n5888# 0.01826f
C575 source.n227 a_n1352_n5888# 0.019334f
C576 source.n228 a_n1352_n5888# 0.043159f
C577 source.n229 a_n1352_n5888# 0.043159f
C578 source.n230 a_n1352_n5888# 0.019334f
C579 source.n231 a_n1352_n5888# 0.01826f
C580 source.n232 a_n1352_n5888# 0.03398f
C581 source.n233 a_n1352_n5888# 0.03398f
C582 source.n234 a_n1352_n5888# 0.01826f
C583 source.n235 a_n1352_n5888# 0.019334f
C584 source.n236 a_n1352_n5888# 0.043159f
C585 source.n237 a_n1352_n5888# 0.043159f
C586 source.n238 a_n1352_n5888# 0.019334f
C587 source.n239 a_n1352_n5888# 0.01826f
C588 source.n240 a_n1352_n5888# 0.03398f
C589 source.n241 a_n1352_n5888# 0.03398f
C590 source.n242 a_n1352_n5888# 0.01826f
C591 source.n243 a_n1352_n5888# 0.019334f
C592 source.n244 a_n1352_n5888# 0.043159f
C593 source.n245 a_n1352_n5888# 0.043159f
C594 source.n246 a_n1352_n5888# 0.019334f
C595 source.n247 a_n1352_n5888# 0.01826f
C596 source.n248 a_n1352_n5888# 0.03398f
C597 source.n249 a_n1352_n5888# 0.03398f
C598 source.n250 a_n1352_n5888# 0.01826f
C599 source.n251 a_n1352_n5888# 0.019334f
C600 source.n252 a_n1352_n5888# 0.043159f
C601 source.n253 a_n1352_n5888# 0.043159f
C602 source.n254 a_n1352_n5888# 0.019334f
C603 source.n255 a_n1352_n5888# 0.01826f
C604 source.n256 a_n1352_n5888# 0.03398f
C605 source.n257 a_n1352_n5888# 0.03398f
C606 source.n258 a_n1352_n5888# 0.01826f
C607 source.n259 a_n1352_n5888# 0.018797f
C608 source.n260 a_n1352_n5888# 0.018797f
C609 source.n261 a_n1352_n5888# 0.043159f
C610 source.n262 a_n1352_n5888# 0.043159f
C611 source.n263 a_n1352_n5888# 0.019334f
C612 source.n264 a_n1352_n5888# 0.01826f
C613 source.n265 a_n1352_n5888# 0.03398f
C614 source.n266 a_n1352_n5888# 0.03398f
C615 source.n267 a_n1352_n5888# 0.01826f
C616 source.n268 a_n1352_n5888# 0.019334f
C617 source.n269 a_n1352_n5888# 0.043159f
C618 source.n270 a_n1352_n5888# 0.043159f
C619 source.n271 a_n1352_n5888# 0.019334f
C620 source.n272 a_n1352_n5888# 0.01826f
C621 source.n273 a_n1352_n5888# 0.03398f
C622 source.n274 a_n1352_n5888# 0.03398f
C623 source.n275 a_n1352_n5888# 0.01826f
C624 source.n276 a_n1352_n5888# 0.019334f
C625 source.n277 a_n1352_n5888# 0.043159f
C626 source.n278 a_n1352_n5888# 0.09181f
C627 source.n279 a_n1352_n5888# 0.019334f
C628 source.n280 a_n1352_n5888# 0.01826f
C629 source.n281 a_n1352_n5888# 0.07483f
C630 source.n282 a_n1352_n5888# 0.051088f
C631 source.n283 a_n1352_n5888# 0.153411f
C632 source.t0 a_n1352_n5888# 0.671308f
C633 source.t9 a_n1352_n5888# 0.671308f
C634 source.n284 a_n1352_n5888# 6.07543f
C635 source.n285 a_n1352_n5888# 0.452497f
C636 source.t1 a_n1352_n5888# 0.671308f
C637 source.t4 a_n1352_n5888# 0.671308f
C638 source.n286 a_n1352_n5888# 6.07543f
C639 source.n287 a_n1352_n5888# 3.65588f
C640 source.t13 a_n1352_n5888# 0.671308f
C641 source.t14 a_n1352_n5888# 0.671308f
C642 source.n288 a_n1352_n5888# 6.07543f
C643 source.n289 a_n1352_n5888# 3.65588f
C644 source.t10 a_n1352_n5888# 0.671308f
C645 source.t19 a_n1352_n5888# 0.671308f
C646 source.n290 a_n1352_n5888# 6.07543f
C647 source.n291 a_n1352_n5888# 0.4525f
C648 source.n292 a_n1352_n5888# 0.046845f
C649 source.n293 a_n1352_n5888# 0.03398f
C650 source.n294 a_n1352_n5888# 0.01826f
C651 source.n295 a_n1352_n5888# 0.043159f
C652 source.n296 a_n1352_n5888# 0.019334f
C653 source.n297 a_n1352_n5888# 0.03398f
C654 source.n298 a_n1352_n5888# 0.01826f
C655 source.n299 a_n1352_n5888# 0.043159f
C656 source.n300 a_n1352_n5888# 0.019334f
C657 source.n301 a_n1352_n5888# 0.03398f
C658 source.n302 a_n1352_n5888# 0.01826f
C659 source.n303 a_n1352_n5888# 0.043159f
C660 source.n304 a_n1352_n5888# 0.019334f
C661 source.n305 a_n1352_n5888# 0.03398f
C662 source.n306 a_n1352_n5888# 0.01826f
C663 source.n307 a_n1352_n5888# 0.043159f
C664 source.n308 a_n1352_n5888# 0.019334f
C665 source.n309 a_n1352_n5888# 0.03398f
C666 source.n310 a_n1352_n5888# 0.01826f
C667 source.n311 a_n1352_n5888# 0.043159f
C668 source.n312 a_n1352_n5888# 0.019334f
C669 source.n313 a_n1352_n5888# 0.03398f
C670 source.n314 a_n1352_n5888# 0.01826f
C671 source.n315 a_n1352_n5888# 0.043159f
C672 source.n316 a_n1352_n5888# 0.019334f
C673 source.n317 a_n1352_n5888# 0.03398f
C674 source.n318 a_n1352_n5888# 0.01826f
C675 source.n319 a_n1352_n5888# 0.043159f
C676 source.n320 a_n1352_n5888# 0.019334f
C677 source.n321 a_n1352_n5888# 0.03398f
C678 source.n322 a_n1352_n5888# 0.01826f
C679 source.n323 a_n1352_n5888# 0.043159f
C680 source.n324 a_n1352_n5888# 0.019334f
C681 source.n325 a_n1352_n5888# 0.03398f
C682 source.n326 a_n1352_n5888# 0.018797f
C683 source.n327 a_n1352_n5888# 0.043159f
C684 source.n328 a_n1352_n5888# 0.019334f
C685 source.n329 a_n1352_n5888# 0.03398f
C686 source.n330 a_n1352_n5888# 0.01826f
C687 source.n331 a_n1352_n5888# 0.043159f
C688 source.n332 a_n1352_n5888# 0.019334f
C689 source.n333 a_n1352_n5888# 0.03398f
C690 source.n334 a_n1352_n5888# 0.01826f
C691 source.n335 a_n1352_n5888# 0.032369f
C692 source.n336 a_n1352_n5888# 0.03051f
C693 source.t11 a_n1352_n5888# 0.075272f
C694 source.n337 a_n1352_n5888# 0.414589f
C695 source.n338 a_n1352_n5888# 3.67907f
C696 source.n339 a_n1352_n5888# 0.01826f
C697 source.n340 a_n1352_n5888# 0.019334f
C698 source.n341 a_n1352_n5888# 0.043159f
C699 source.n342 a_n1352_n5888# 0.043159f
C700 source.n343 a_n1352_n5888# 0.019334f
C701 source.n344 a_n1352_n5888# 0.01826f
C702 source.n345 a_n1352_n5888# 0.03398f
C703 source.n346 a_n1352_n5888# 0.03398f
C704 source.n347 a_n1352_n5888# 0.01826f
C705 source.n348 a_n1352_n5888# 0.019334f
C706 source.n349 a_n1352_n5888# 0.043159f
C707 source.n350 a_n1352_n5888# 0.043159f
C708 source.n351 a_n1352_n5888# 0.019334f
C709 source.n352 a_n1352_n5888# 0.01826f
C710 source.n353 a_n1352_n5888# 0.03398f
C711 source.n354 a_n1352_n5888# 0.03398f
C712 source.n355 a_n1352_n5888# 0.01826f
C713 source.n356 a_n1352_n5888# 0.01826f
C714 source.n357 a_n1352_n5888# 0.019334f
C715 source.n358 a_n1352_n5888# 0.043159f
C716 source.n359 a_n1352_n5888# 0.043159f
C717 source.n360 a_n1352_n5888# 0.043159f
C718 source.n361 a_n1352_n5888# 0.018797f
C719 source.n362 a_n1352_n5888# 0.01826f
C720 source.n363 a_n1352_n5888# 0.03398f
C721 source.n364 a_n1352_n5888# 0.03398f
C722 source.n365 a_n1352_n5888# 0.01826f
C723 source.n366 a_n1352_n5888# 0.019334f
C724 source.n367 a_n1352_n5888# 0.043159f
C725 source.n368 a_n1352_n5888# 0.043159f
C726 source.n369 a_n1352_n5888# 0.019334f
C727 source.n370 a_n1352_n5888# 0.01826f
C728 source.n371 a_n1352_n5888# 0.03398f
C729 source.n372 a_n1352_n5888# 0.03398f
C730 source.n373 a_n1352_n5888# 0.01826f
C731 source.n374 a_n1352_n5888# 0.019334f
C732 source.n375 a_n1352_n5888# 0.043159f
C733 source.n376 a_n1352_n5888# 0.043159f
C734 source.n377 a_n1352_n5888# 0.019334f
C735 source.n378 a_n1352_n5888# 0.01826f
C736 source.n379 a_n1352_n5888# 0.03398f
C737 source.n380 a_n1352_n5888# 0.03398f
C738 source.n381 a_n1352_n5888# 0.01826f
C739 source.n382 a_n1352_n5888# 0.019334f
C740 source.n383 a_n1352_n5888# 0.043159f
C741 source.n384 a_n1352_n5888# 0.043159f
C742 source.n385 a_n1352_n5888# 0.019334f
C743 source.n386 a_n1352_n5888# 0.01826f
C744 source.n387 a_n1352_n5888# 0.03398f
C745 source.n388 a_n1352_n5888# 0.03398f
C746 source.n389 a_n1352_n5888# 0.01826f
C747 source.n390 a_n1352_n5888# 0.019334f
C748 source.n391 a_n1352_n5888# 0.043159f
C749 source.n392 a_n1352_n5888# 0.043159f
C750 source.n393 a_n1352_n5888# 0.019334f
C751 source.n394 a_n1352_n5888# 0.01826f
C752 source.n395 a_n1352_n5888# 0.03398f
C753 source.n396 a_n1352_n5888# 0.03398f
C754 source.n397 a_n1352_n5888# 0.01826f
C755 source.n398 a_n1352_n5888# 0.019334f
C756 source.n399 a_n1352_n5888# 0.043159f
C757 source.n400 a_n1352_n5888# 0.043159f
C758 source.n401 a_n1352_n5888# 0.043159f
C759 source.n402 a_n1352_n5888# 0.019334f
C760 source.n403 a_n1352_n5888# 0.01826f
C761 source.n404 a_n1352_n5888# 0.03398f
C762 source.n405 a_n1352_n5888# 0.03398f
C763 source.n406 a_n1352_n5888# 0.01826f
C764 source.n407 a_n1352_n5888# 0.018797f
C765 source.n408 a_n1352_n5888# 0.018797f
C766 source.n409 a_n1352_n5888# 0.043159f
C767 source.n410 a_n1352_n5888# 0.043159f
C768 source.n411 a_n1352_n5888# 0.019334f
C769 source.n412 a_n1352_n5888# 0.01826f
C770 source.n413 a_n1352_n5888# 0.03398f
C771 source.n414 a_n1352_n5888# 0.03398f
C772 source.n415 a_n1352_n5888# 0.01826f
C773 source.n416 a_n1352_n5888# 0.019334f
C774 source.n417 a_n1352_n5888# 0.043159f
C775 source.n418 a_n1352_n5888# 0.043159f
C776 source.n419 a_n1352_n5888# 0.019334f
C777 source.n420 a_n1352_n5888# 0.01826f
C778 source.n421 a_n1352_n5888# 0.03398f
C779 source.n422 a_n1352_n5888# 0.03398f
C780 source.n423 a_n1352_n5888# 0.01826f
C781 source.n424 a_n1352_n5888# 0.019334f
C782 source.n425 a_n1352_n5888# 0.043159f
C783 source.n426 a_n1352_n5888# 0.09181f
C784 source.n427 a_n1352_n5888# 0.019334f
C785 source.n428 a_n1352_n5888# 0.01826f
C786 source.n429 a_n1352_n5888# 0.07483f
C787 source.n430 a_n1352_n5888# 0.051088f
C788 source.n431 a_n1352_n5888# 0.153411f
C789 source.t3 a_n1352_n5888# 0.671308f
C790 source.t6 a_n1352_n5888# 0.671308f
C791 source.n432 a_n1352_n5888# 6.07543f
C792 source.n433 a_n1352_n5888# 0.478929f
C793 source.t5 a_n1352_n5888# 0.671308f
C794 source.t2 a_n1352_n5888# 0.671308f
C795 source.n434 a_n1352_n5888# 6.07543f
C796 source.n435 a_n1352_n5888# 0.4525f
C797 source.n436 a_n1352_n5888# 0.046845f
C798 source.n437 a_n1352_n5888# 0.03398f
C799 source.n438 a_n1352_n5888# 0.01826f
C800 source.n439 a_n1352_n5888# 0.043159f
C801 source.n440 a_n1352_n5888# 0.019334f
C802 source.n441 a_n1352_n5888# 0.03398f
C803 source.n442 a_n1352_n5888# 0.01826f
C804 source.n443 a_n1352_n5888# 0.043159f
C805 source.n444 a_n1352_n5888# 0.019334f
C806 source.n445 a_n1352_n5888# 0.03398f
C807 source.n446 a_n1352_n5888# 0.01826f
C808 source.n447 a_n1352_n5888# 0.043159f
C809 source.n448 a_n1352_n5888# 0.019334f
C810 source.n449 a_n1352_n5888# 0.03398f
C811 source.n450 a_n1352_n5888# 0.01826f
C812 source.n451 a_n1352_n5888# 0.043159f
C813 source.n452 a_n1352_n5888# 0.019334f
C814 source.n453 a_n1352_n5888# 0.03398f
C815 source.n454 a_n1352_n5888# 0.01826f
C816 source.n455 a_n1352_n5888# 0.043159f
C817 source.n456 a_n1352_n5888# 0.019334f
C818 source.n457 a_n1352_n5888# 0.03398f
C819 source.n458 a_n1352_n5888# 0.01826f
C820 source.n459 a_n1352_n5888# 0.043159f
C821 source.n460 a_n1352_n5888# 0.019334f
C822 source.n461 a_n1352_n5888# 0.03398f
C823 source.n462 a_n1352_n5888# 0.01826f
C824 source.n463 a_n1352_n5888# 0.043159f
C825 source.n464 a_n1352_n5888# 0.019334f
C826 source.n465 a_n1352_n5888# 0.03398f
C827 source.n466 a_n1352_n5888# 0.01826f
C828 source.n467 a_n1352_n5888# 0.043159f
C829 source.n468 a_n1352_n5888# 0.019334f
C830 source.n469 a_n1352_n5888# 0.03398f
C831 source.n470 a_n1352_n5888# 0.018797f
C832 source.n471 a_n1352_n5888# 0.043159f
C833 source.n472 a_n1352_n5888# 0.019334f
C834 source.n473 a_n1352_n5888# 0.03398f
C835 source.n474 a_n1352_n5888# 0.01826f
C836 source.n475 a_n1352_n5888# 0.043159f
C837 source.n476 a_n1352_n5888# 0.019334f
C838 source.n477 a_n1352_n5888# 0.03398f
C839 source.n478 a_n1352_n5888# 0.01826f
C840 source.n479 a_n1352_n5888# 0.032369f
C841 source.n480 a_n1352_n5888# 0.03051f
C842 source.t8 a_n1352_n5888# 0.075272f
C843 source.n481 a_n1352_n5888# 0.414589f
C844 source.n482 a_n1352_n5888# 3.67907f
C845 source.n483 a_n1352_n5888# 0.01826f
C846 source.n484 a_n1352_n5888# 0.019334f
C847 source.n485 a_n1352_n5888# 0.043159f
C848 source.n486 a_n1352_n5888# 0.043159f
C849 source.n487 a_n1352_n5888# 0.019334f
C850 source.n488 a_n1352_n5888# 0.01826f
C851 source.n489 a_n1352_n5888# 0.03398f
C852 source.n490 a_n1352_n5888# 0.03398f
C853 source.n491 a_n1352_n5888# 0.01826f
C854 source.n492 a_n1352_n5888# 0.019334f
C855 source.n493 a_n1352_n5888# 0.043159f
C856 source.n494 a_n1352_n5888# 0.043159f
C857 source.n495 a_n1352_n5888# 0.019334f
C858 source.n496 a_n1352_n5888# 0.01826f
C859 source.n497 a_n1352_n5888# 0.03398f
C860 source.n498 a_n1352_n5888# 0.03398f
C861 source.n499 a_n1352_n5888# 0.01826f
C862 source.n500 a_n1352_n5888# 0.01826f
C863 source.n501 a_n1352_n5888# 0.019334f
C864 source.n502 a_n1352_n5888# 0.043159f
C865 source.n503 a_n1352_n5888# 0.043159f
C866 source.n504 a_n1352_n5888# 0.043159f
C867 source.n505 a_n1352_n5888# 0.018797f
C868 source.n506 a_n1352_n5888# 0.01826f
C869 source.n507 a_n1352_n5888# 0.03398f
C870 source.n508 a_n1352_n5888# 0.03398f
C871 source.n509 a_n1352_n5888# 0.01826f
C872 source.n510 a_n1352_n5888# 0.019334f
C873 source.n511 a_n1352_n5888# 0.043159f
C874 source.n512 a_n1352_n5888# 0.043159f
C875 source.n513 a_n1352_n5888# 0.019334f
C876 source.n514 a_n1352_n5888# 0.01826f
C877 source.n515 a_n1352_n5888# 0.03398f
C878 source.n516 a_n1352_n5888# 0.03398f
C879 source.n517 a_n1352_n5888# 0.01826f
C880 source.n518 a_n1352_n5888# 0.019334f
C881 source.n519 a_n1352_n5888# 0.043159f
C882 source.n520 a_n1352_n5888# 0.043159f
C883 source.n521 a_n1352_n5888# 0.019334f
C884 source.n522 a_n1352_n5888# 0.01826f
C885 source.n523 a_n1352_n5888# 0.03398f
C886 source.n524 a_n1352_n5888# 0.03398f
C887 source.n525 a_n1352_n5888# 0.01826f
C888 source.n526 a_n1352_n5888# 0.019334f
C889 source.n527 a_n1352_n5888# 0.043159f
C890 source.n528 a_n1352_n5888# 0.043159f
C891 source.n529 a_n1352_n5888# 0.019334f
C892 source.n530 a_n1352_n5888# 0.01826f
C893 source.n531 a_n1352_n5888# 0.03398f
C894 source.n532 a_n1352_n5888# 0.03398f
C895 source.n533 a_n1352_n5888# 0.01826f
C896 source.n534 a_n1352_n5888# 0.019334f
C897 source.n535 a_n1352_n5888# 0.043159f
C898 source.n536 a_n1352_n5888# 0.043159f
C899 source.n537 a_n1352_n5888# 0.019334f
C900 source.n538 a_n1352_n5888# 0.01826f
C901 source.n539 a_n1352_n5888# 0.03398f
C902 source.n540 a_n1352_n5888# 0.03398f
C903 source.n541 a_n1352_n5888# 0.01826f
C904 source.n542 a_n1352_n5888# 0.019334f
C905 source.n543 a_n1352_n5888# 0.043159f
C906 source.n544 a_n1352_n5888# 0.043159f
C907 source.n545 a_n1352_n5888# 0.043159f
C908 source.n546 a_n1352_n5888# 0.019334f
C909 source.n547 a_n1352_n5888# 0.01826f
C910 source.n548 a_n1352_n5888# 0.03398f
C911 source.n549 a_n1352_n5888# 0.03398f
C912 source.n550 a_n1352_n5888# 0.01826f
C913 source.n551 a_n1352_n5888# 0.018797f
C914 source.n552 a_n1352_n5888# 0.018797f
C915 source.n553 a_n1352_n5888# 0.043159f
C916 source.n554 a_n1352_n5888# 0.043159f
C917 source.n555 a_n1352_n5888# 0.019334f
C918 source.n556 a_n1352_n5888# 0.01826f
C919 source.n557 a_n1352_n5888# 0.03398f
C920 source.n558 a_n1352_n5888# 0.03398f
C921 source.n559 a_n1352_n5888# 0.01826f
C922 source.n560 a_n1352_n5888# 0.019334f
C923 source.n561 a_n1352_n5888# 0.043159f
C924 source.n562 a_n1352_n5888# 0.043159f
C925 source.n563 a_n1352_n5888# 0.019334f
C926 source.n564 a_n1352_n5888# 0.01826f
C927 source.n565 a_n1352_n5888# 0.03398f
C928 source.n566 a_n1352_n5888# 0.03398f
C929 source.n567 a_n1352_n5888# 0.01826f
C930 source.n568 a_n1352_n5888# 0.019334f
C931 source.n569 a_n1352_n5888# 0.043159f
C932 source.n570 a_n1352_n5888# 0.09181f
C933 source.n571 a_n1352_n5888# 0.019334f
C934 source.n572 a_n1352_n5888# 0.01826f
C935 source.n573 a_n1352_n5888# 0.07483f
C936 source.n574 a_n1352_n5888# 0.051088f
C937 source.n575 a_n1352_n5888# 0.31265f
C938 source.n576 a_n1352_n5888# 3.61622f
C939 drain_left.n0 a_n1352_n5888# 0.046604f
C940 drain_left.n1 a_n1352_n5888# 0.033805f
C941 drain_left.n2 a_n1352_n5888# 0.018166f
C942 drain_left.n3 a_n1352_n5888# 0.042937f
C943 drain_left.n4 a_n1352_n5888# 0.019234f
C944 drain_left.n5 a_n1352_n5888# 0.033805f
C945 drain_left.n6 a_n1352_n5888# 0.018166f
C946 drain_left.n7 a_n1352_n5888# 0.042937f
C947 drain_left.n8 a_n1352_n5888# 0.019234f
C948 drain_left.n9 a_n1352_n5888# 0.033805f
C949 drain_left.n10 a_n1352_n5888# 0.018166f
C950 drain_left.n11 a_n1352_n5888# 0.042937f
C951 drain_left.n12 a_n1352_n5888# 0.019234f
C952 drain_left.n13 a_n1352_n5888# 0.033805f
C953 drain_left.n14 a_n1352_n5888# 0.018166f
C954 drain_left.n15 a_n1352_n5888# 0.042937f
C955 drain_left.n16 a_n1352_n5888# 0.019234f
C956 drain_left.n17 a_n1352_n5888# 0.033805f
C957 drain_left.n18 a_n1352_n5888# 0.018166f
C958 drain_left.n19 a_n1352_n5888# 0.042937f
C959 drain_left.n20 a_n1352_n5888# 0.019234f
C960 drain_left.n21 a_n1352_n5888# 0.033805f
C961 drain_left.n22 a_n1352_n5888# 0.018166f
C962 drain_left.n23 a_n1352_n5888# 0.042937f
C963 drain_left.n24 a_n1352_n5888# 0.019234f
C964 drain_left.n25 a_n1352_n5888# 0.033805f
C965 drain_left.n26 a_n1352_n5888# 0.018166f
C966 drain_left.n27 a_n1352_n5888# 0.042937f
C967 drain_left.n28 a_n1352_n5888# 0.019234f
C968 drain_left.n29 a_n1352_n5888# 0.033805f
C969 drain_left.n30 a_n1352_n5888# 0.018166f
C970 drain_left.n31 a_n1352_n5888# 0.042937f
C971 drain_left.n32 a_n1352_n5888# 0.019234f
C972 drain_left.n33 a_n1352_n5888# 0.033805f
C973 drain_left.n34 a_n1352_n5888# 0.0187f
C974 drain_left.n35 a_n1352_n5888# 0.042937f
C975 drain_left.n36 a_n1352_n5888# 0.019234f
C976 drain_left.n37 a_n1352_n5888# 0.033805f
C977 drain_left.n38 a_n1352_n5888# 0.018166f
C978 drain_left.n39 a_n1352_n5888# 0.042937f
C979 drain_left.n40 a_n1352_n5888# 0.019234f
C980 drain_left.n41 a_n1352_n5888# 0.033805f
C981 drain_left.n42 a_n1352_n5888# 0.018166f
C982 drain_left.n43 a_n1352_n5888# 0.032203f
C983 drain_left.n44 a_n1352_n5888# 0.030353f
C984 drain_left.t5 a_n1352_n5888# 0.074885f
C985 drain_left.n45 a_n1352_n5888# 0.412456f
C986 drain_left.n46 a_n1352_n5888# 3.66014f
C987 drain_left.n47 a_n1352_n5888# 0.018166f
C988 drain_left.n48 a_n1352_n5888# 0.019234f
C989 drain_left.n49 a_n1352_n5888# 0.042937f
C990 drain_left.n50 a_n1352_n5888# 0.042937f
C991 drain_left.n51 a_n1352_n5888# 0.019234f
C992 drain_left.n52 a_n1352_n5888# 0.018166f
C993 drain_left.n53 a_n1352_n5888# 0.033805f
C994 drain_left.n54 a_n1352_n5888# 0.033805f
C995 drain_left.n55 a_n1352_n5888# 0.018166f
C996 drain_left.n56 a_n1352_n5888# 0.019234f
C997 drain_left.n57 a_n1352_n5888# 0.042937f
C998 drain_left.n58 a_n1352_n5888# 0.042937f
C999 drain_left.n59 a_n1352_n5888# 0.019234f
C1000 drain_left.n60 a_n1352_n5888# 0.018166f
C1001 drain_left.n61 a_n1352_n5888# 0.033805f
C1002 drain_left.n62 a_n1352_n5888# 0.033805f
C1003 drain_left.n63 a_n1352_n5888# 0.018166f
C1004 drain_left.n64 a_n1352_n5888# 0.018166f
C1005 drain_left.n65 a_n1352_n5888# 0.019234f
C1006 drain_left.n66 a_n1352_n5888# 0.042937f
C1007 drain_left.n67 a_n1352_n5888# 0.042937f
C1008 drain_left.n68 a_n1352_n5888# 0.042937f
C1009 drain_left.n69 a_n1352_n5888# 0.0187f
C1010 drain_left.n70 a_n1352_n5888# 0.018166f
C1011 drain_left.n71 a_n1352_n5888# 0.033805f
C1012 drain_left.n72 a_n1352_n5888# 0.033805f
C1013 drain_left.n73 a_n1352_n5888# 0.018166f
C1014 drain_left.n74 a_n1352_n5888# 0.019234f
C1015 drain_left.n75 a_n1352_n5888# 0.042937f
C1016 drain_left.n76 a_n1352_n5888# 0.042937f
C1017 drain_left.n77 a_n1352_n5888# 0.019234f
C1018 drain_left.n78 a_n1352_n5888# 0.018166f
C1019 drain_left.n79 a_n1352_n5888# 0.033805f
C1020 drain_left.n80 a_n1352_n5888# 0.033805f
C1021 drain_left.n81 a_n1352_n5888# 0.018166f
C1022 drain_left.n82 a_n1352_n5888# 0.019234f
C1023 drain_left.n83 a_n1352_n5888# 0.042937f
C1024 drain_left.n84 a_n1352_n5888# 0.042937f
C1025 drain_left.n85 a_n1352_n5888# 0.019234f
C1026 drain_left.n86 a_n1352_n5888# 0.018166f
C1027 drain_left.n87 a_n1352_n5888# 0.033805f
C1028 drain_left.n88 a_n1352_n5888# 0.033805f
C1029 drain_left.n89 a_n1352_n5888# 0.018166f
C1030 drain_left.n90 a_n1352_n5888# 0.019234f
C1031 drain_left.n91 a_n1352_n5888# 0.042937f
C1032 drain_left.n92 a_n1352_n5888# 0.042937f
C1033 drain_left.n93 a_n1352_n5888# 0.019234f
C1034 drain_left.n94 a_n1352_n5888# 0.018166f
C1035 drain_left.n95 a_n1352_n5888# 0.033805f
C1036 drain_left.n96 a_n1352_n5888# 0.033805f
C1037 drain_left.n97 a_n1352_n5888# 0.018166f
C1038 drain_left.n98 a_n1352_n5888# 0.019234f
C1039 drain_left.n99 a_n1352_n5888# 0.042937f
C1040 drain_left.n100 a_n1352_n5888# 0.042937f
C1041 drain_left.n101 a_n1352_n5888# 0.019234f
C1042 drain_left.n102 a_n1352_n5888# 0.018166f
C1043 drain_left.n103 a_n1352_n5888# 0.033805f
C1044 drain_left.n104 a_n1352_n5888# 0.033805f
C1045 drain_left.n105 a_n1352_n5888# 0.018166f
C1046 drain_left.n106 a_n1352_n5888# 0.019234f
C1047 drain_left.n107 a_n1352_n5888# 0.042937f
C1048 drain_left.n108 a_n1352_n5888# 0.042937f
C1049 drain_left.n109 a_n1352_n5888# 0.042937f
C1050 drain_left.n110 a_n1352_n5888# 0.019234f
C1051 drain_left.n111 a_n1352_n5888# 0.018166f
C1052 drain_left.n112 a_n1352_n5888# 0.033805f
C1053 drain_left.n113 a_n1352_n5888# 0.033805f
C1054 drain_left.n114 a_n1352_n5888# 0.018166f
C1055 drain_left.n115 a_n1352_n5888# 0.0187f
C1056 drain_left.n116 a_n1352_n5888# 0.0187f
C1057 drain_left.n117 a_n1352_n5888# 0.042937f
C1058 drain_left.n118 a_n1352_n5888# 0.042937f
C1059 drain_left.n119 a_n1352_n5888# 0.019234f
C1060 drain_left.n120 a_n1352_n5888# 0.018166f
C1061 drain_left.n121 a_n1352_n5888# 0.033805f
C1062 drain_left.n122 a_n1352_n5888# 0.033805f
C1063 drain_left.n123 a_n1352_n5888# 0.018166f
C1064 drain_left.n124 a_n1352_n5888# 0.019234f
C1065 drain_left.n125 a_n1352_n5888# 0.042937f
C1066 drain_left.n126 a_n1352_n5888# 0.042937f
C1067 drain_left.n127 a_n1352_n5888# 0.019234f
C1068 drain_left.n128 a_n1352_n5888# 0.018166f
C1069 drain_left.n129 a_n1352_n5888# 0.033805f
C1070 drain_left.n130 a_n1352_n5888# 0.033805f
C1071 drain_left.n131 a_n1352_n5888# 0.018166f
C1072 drain_left.n132 a_n1352_n5888# 0.019234f
C1073 drain_left.n133 a_n1352_n5888# 0.042937f
C1074 drain_left.n134 a_n1352_n5888# 0.091338f
C1075 drain_left.n135 a_n1352_n5888# 0.019234f
C1076 drain_left.n136 a_n1352_n5888# 0.018166f
C1077 drain_left.n137 a_n1352_n5888# 0.074445f
C1078 drain_left.n138 a_n1352_n5888# 0.075277f
C1079 drain_left.t2 a_n1352_n5888# 0.667854f
C1080 drain_left.t8 a_n1352_n5888# 0.667854f
C1081 drain_left.n139 a_n1352_n5888# 6.15499f
C1082 drain_left.n140 a_n1352_n5888# 0.466921f
C1083 drain_left.t7 a_n1352_n5888# 0.667854f
C1084 drain_left.t9 a_n1352_n5888# 0.667854f
C1085 drain_left.n141 a_n1352_n5888# 6.15686f
C1086 drain_left.n142 a_n1352_n5888# 2.95722f
C1087 drain_left.n143 a_n1352_n5888# 0.046604f
C1088 drain_left.n144 a_n1352_n5888# 0.033805f
C1089 drain_left.n145 a_n1352_n5888# 0.018166f
C1090 drain_left.n146 a_n1352_n5888# 0.042937f
C1091 drain_left.n147 a_n1352_n5888# 0.019234f
C1092 drain_left.n148 a_n1352_n5888# 0.033805f
C1093 drain_left.n149 a_n1352_n5888# 0.018166f
C1094 drain_left.n150 a_n1352_n5888# 0.042937f
C1095 drain_left.n151 a_n1352_n5888# 0.019234f
C1096 drain_left.n152 a_n1352_n5888# 0.033805f
C1097 drain_left.n153 a_n1352_n5888# 0.018166f
C1098 drain_left.n154 a_n1352_n5888# 0.042937f
C1099 drain_left.n155 a_n1352_n5888# 0.019234f
C1100 drain_left.n156 a_n1352_n5888# 0.033805f
C1101 drain_left.n157 a_n1352_n5888# 0.018166f
C1102 drain_left.n158 a_n1352_n5888# 0.042937f
C1103 drain_left.n159 a_n1352_n5888# 0.042937f
C1104 drain_left.n160 a_n1352_n5888# 0.019234f
C1105 drain_left.n161 a_n1352_n5888# 0.033805f
C1106 drain_left.n162 a_n1352_n5888# 0.018166f
C1107 drain_left.n163 a_n1352_n5888# 0.042937f
C1108 drain_left.n164 a_n1352_n5888# 0.019234f
C1109 drain_left.n165 a_n1352_n5888# 0.033805f
C1110 drain_left.n166 a_n1352_n5888# 0.018166f
C1111 drain_left.n167 a_n1352_n5888# 0.042937f
C1112 drain_left.n168 a_n1352_n5888# 0.019234f
C1113 drain_left.n169 a_n1352_n5888# 0.033805f
C1114 drain_left.n170 a_n1352_n5888# 0.018166f
C1115 drain_left.n171 a_n1352_n5888# 0.042937f
C1116 drain_left.n172 a_n1352_n5888# 0.019234f
C1117 drain_left.n173 a_n1352_n5888# 0.033805f
C1118 drain_left.n174 a_n1352_n5888# 0.018166f
C1119 drain_left.n175 a_n1352_n5888# 0.042937f
C1120 drain_left.n176 a_n1352_n5888# 0.019234f
C1121 drain_left.n177 a_n1352_n5888# 0.033805f
C1122 drain_left.n178 a_n1352_n5888# 0.0187f
C1123 drain_left.n179 a_n1352_n5888# 0.042937f
C1124 drain_left.n180 a_n1352_n5888# 0.018166f
C1125 drain_left.n181 a_n1352_n5888# 0.019234f
C1126 drain_left.n182 a_n1352_n5888# 0.033805f
C1127 drain_left.n183 a_n1352_n5888# 0.018166f
C1128 drain_left.n184 a_n1352_n5888# 0.042937f
C1129 drain_left.n185 a_n1352_n5888# 0.019234f
C1130 drain_left.n186 a_n1352_n5888# 0.033805f
C1131 drain_left.n187 a_n1352_n5888# 0.018166f
C1132 drain_left.n188 a_n1352_n5888# 0.032203f
C1133 drain_left.n189 a_n1352_n5888# 0.030353f
C1134 drain_left.t1 a_n1352_n5888# 0.074885f
C1135 drain_left.n190 a_n1352_n5888# 0.412456f
C1136 drain_left.n191 a_n1352_n5888# 3.66014f
C1137 drain_left.n192 a_n1352_n5888# 0.018166f
C1138 drain_left.n193 a_n1352_n5888# 0.019234f
C1139 drain_left.n194 a_n1352_n5888# 0.042937f
C1140 drain_left.n195 a_n1352_n5888# 0.042937f
C1141 drain_left.n196 a_n1352_n5888# 0.019234f
C1142 drain_left.n197 a_n1352_n5888# 0.018166f
C1143 drain_left.n198 a_n1352_n5888# 0.033805f
C1144 drain_left.n199 a_n1352_n5888# 0.033805f
C1145 drain_left.n200 a_n1352_n5888# 0.018166f
C1146 drain_left.n201 a_n1352_n5888# 0.019234f
C1147 drain_left.n202 a_n1352_n5888# 0.042937f
C1148 drain_left.n203 a_n1352_n5888# 0.042937f
C1149 drain_left.n204 a_n1352_n5888# 0.019234f
C1150 drain_left.n205 a_n1352_n5888# 0.018166f
C1151 drain_left.n206 a_n1352_n5888# 0.033805f
C1152 drain_left.n207 a_n1352_n5888# 0.033805f
C1153 drain_left.n208 a_n1352_n5888# 0.018166f
C1154 drain_left.n209 a_n1352_n5888# 0.019234f
C1155 drain_left.n210 a_n1352_n5888# 0.042937f
C1156 drain_left.n211 a_n1352_n5888# 0.042937f
C1157 drain_left.n212 a_n1352_n5888# 0.042937f
C1158 drain_left.n213 a_n1352_n5888# 0.0187f
C1159 drain_left.n214 a_n1352_n5888# 0.018166f
C1160 drain_left.n215 a_n1352_n5888# 0.033805f
C1161 drain_left.n216 a_n1352_n5888# 0.033805f
C1162 drain_left.n217 a_n1352_n5888# 0.018166f
C1163 drain_left.n218 a_n1352_n5888# 0.019234f
C1164 drain_left.n219 a_n1352_n5888# 0.042937f
C1165 drain_left.n220 a_n1352_n5888# 0.042937f
C1166 drain_left.n221 a_n1352_n5888# 0.019234f
C1167 drain_left.n222 a_n1352_n5888# 0.018166f
C1168 drain_left.n223 a_n1352_n5888# 0.033805f
C1169 drain_left.n224 a_n1352_n5888# 0.033805f
C1170 drain_left.n225 a_n1352_n5888# 0.018166f
C1171 drain_left.n226 a_n1352_n5888# 0.019234f
C1172 drain_left.n227 a_n1352_n5888# 0.042937f
C1173 drain_left.n228 a_n1352_n5888# 0.042937f
C1174 drain_left.n229 a_n1352_n5888# 0.019234f
C1175 drain_left.n230 a_n1352_n5888# 0.018166f
C1176 drain_left.n231 a_n1352_n5888# 0.033805f
C1177 drain_left.n232 a_n1352_n5888# 0.033805f
C1178 drain_left.n233 a_n1352_n5888# 0.018166f
C1179 drain_left.n234 a_n1352_n5888# 0.019234f
C1180 drain_left.n235 a_n1352_n5888# 0.042937f
C1181 drain_left.n236 a_n1352_n5888# 0.042937f
C1182 drain_left.n237 a_n1352_n5888# 0.019234f
C1183 drain_left.n238 a_n1352_n5888# 0.018166f
C1184 drain_left.n239 a_n1352_n5888# 0.033805f
C1185 drain_left.n240 a_n1352_n5888# 0.033805f
C1186 drain_left.n241 a_n1352_n5888# 0.018166f
C1187 drain_left.n242 a_n1352_n5888# 0.019234f
C1188 drain_left.n243 a_n1352_n5888# 0.042937f
C1189 drain_left.n244 a_n1352_n5888# 0.042937f
C1190 drain_left.n245 a_n1352_n5888# 0.019234f
C1191 drain_left.n246 a_n1352_n5888# 0.018166f
C1192 drain_left.n247 a_n1352_n5888# 0.033805f
C1193 drain_left.n248 a_n1352_n5888# 0.033805f
C1194 drain_left.n249 a_n1352_n5888# 0.018166f
C1195 drain_left.n250 a_n1352_n5888# 0.019234f
C1196 drain_left.n251 a_n1352_n5888# 0.042937f
C1197 drain_left.n252 a_n1352_n5888# 0.042937f
C1198 drain_left.n253 a_n1352_n5888# 0.019234f
C1199 drain_left.n254 a_n1352_n5888# 0.018166f
C1200 drain_left.n255 a_n1352_n5888# 0.033805f
C1201 drain_left.n256 a_n1352_n5888# 0.033805f
C1202 drain_left.n257 a_n1352_n5888# 0.018166f
C1203 drain_left.n258 a_n1352_n5888# 0.0187f
C1204 drain_left.n259 a_n1352_n5888# 0.0187f
C1205 drain_left.n260 a_n1352_n5888# 0.042937f
C1206 drain_left.n261 a_n1352_n5888# 0.042937f
C1207 drain_left.n262 a_n1352_n5888# 0.019234f
C1208 drain_left.n263 a_n1352_n5888# 0.018166f
C1209 drain_left.n264 a_n1352_n5888# 0.033805f
C1210 drain_left.n265 a_n1352_n5888# 0.033805f
C1211 drain_left.n266 a_n1352_n5888# 0.018166f
C1212 drain_left.n267 a_n1352_n5888# 0.019234f
C1213 drain_left.n268 a_n1352_n5888# 0.042937f
C1214 drain_left.n269 a_n1352_n5888# 0.042937f
C1215 drain_left.n270 a_n1352_n5888# 0.019234f
C1216 drain_left.n271 a_n1352_n5888# 0.018166f
C1217 drain_left.n272 a_n1352_n5888# 0.033805f
C1218 drain_left.n273 a_n1352_n5888# 0.033805f
C1219 drain_left.n274 a_n1352_n5888# 0.018166f
C1220 drain_left.n275 a_n1352_n5888# 0.019234f
C1221 drain_left.n276 a_n1352_n5888# 0.042937f
C1222 drain_left.n277 a_n1352_n5888# 0.091338f
C1223 drain_left.n278 a_n1352_n5888# 0.019234f
C1224 drain_left.n279 a_n1352_n5888# 0.018166f
C1225 drain_left.n280 a_n1352_n5888# 0.074445f
C1226 drain_left.n281 a_n1352_n5888# 0.075277f
C1227 drain_left.t6 a_n1352_n5888# 0.667854f
C1228 drain_left.t4 a_n1352_n5888# 0.667854f
C1229 drain_left.n282 a_n1352_n5888# 6.15499f
C1230 drain_left.n283 a_n1352_n5888# 0.496964f
C1231 drain_left.t3 a_n1352_n5888# 0.667854f
C1232 drain_left.t0 a_n1352_n5888# 0.667854f
C1233 drain_left.n284 a_n1352_n5888# 6.15498f
C1234 drain_left.n285 a_n1352_n5888# 0.661973f
C1235 plus.n0 a_n1352_n5888# 0.058853f
C1236 plus.t4 a_n1352_n5888# 0.827965f
C1237 plus.t7 a_n1352_n5888# 0.827965f
C1238 plus.t1 a_n1352_n5888# 0.827965f
C1239 plus.n1 a_n1352_n5888# 0.307326f
C1240 plus.t2 a_n1352_n5888# 0.832299f
C1241 plus.n2 a_n1352_n5888# 0.324049f
C1242 plus.n3 a_n1352_n5888# 0.129234f
C1243 plus.n4 a_n1352_n5888# 0.020612f
C1244 plus.n5 a_n1352_n5888# 0.307326f
C1245 plus.n6 a_n1352_n5888# 0.020612f
C1246 plus.n7 a_n1352_n5888# 0.307326f
C1247 plus.t3 a_n1352_n5888# 0.832299f
C1248 plus.n8 a_n1352_n5888# 0.323966f
C1249 plus.n9 a_n1352_n5888# 1.04385f
C1250 plus.n10 a_n1352_n5888# 0.058853f
C1251 plus.t6 a_n1352_n5888# 0.832299f
C1252 plus.t5 a_n1352_n5888# 0.827965f
C1253 plus.t9 a_n1352_n5888# 0.827965f
C1254 plus.t0 a_n1352_n5888# 0.827965f
C1255 plus.n11 a_n1352_n5888# 0.307326f
C1256 plus.t8 a_n1352_n5888# 0.832299f
C1257 plus.n12 a_n1352_n5888# 0.324049f
C1258 plus.n13 a_n1352_n5888# 0.129234f
C1259 plus.n14 a_n1352_n5888# 0.020612f
C1260 plus.n15 a_n1352_n5888# 0.307326f
C1261 plus.n16 a_n1352_n5888# 0.020612f
C1262 plus.n17 a_n1352_n5888# 0.307326f
C1263 plus.n18 a_n1352_n5888# 0.323966f
C1264 plus.n19 a_n1352_n5888# 2.1165f
.ends

