* NGSPICE file created from diffpair127.ext - technology: sky130A

.subckt diffpair127 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t26 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 drain_right.t14 minus.t1 source.t28 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X2 drain_right.t13 minus.t2 source.t19 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 source.t6 plus.t0 drain_left.t15 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X4 source.t2 plus.t1 drain_left.t14 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X5 source.t30 minus.t3 drain_right.t12 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X6 source.t14 plus.t2 drain_left.t13 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X7 source.t15 plus.t3 drain_left.t12 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X8 source.t24 minus.t4 drain_right.t11 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X9 drain_left.t11 plus.t4 source.t3 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X10 drain_right.t10 minus.t5 source.t29 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X12 drain_right.t9 minus.t6 source.t23 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X13 source.t25 minus.t7 drain_right.t8 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X14 drain_left.t10 plus.t5 source.t9 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X15 drain_left.t9 plus.t6 source.t12 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X16 source.t1 plus.t7 drain_left.t8 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X17 source.t16 minus.t8 drain_right.t7 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X18 source.t31 minus.t9 drain_right.t6 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X19 a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X20 a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X21 drain_right.t5 minus.t10 source.t22 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X22 drain_right.t4 minus.t11 source.t18 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X23 source.t11 plus.t8 drain_left.t7 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X24 a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X25 drain_left.t6 plus.t9 source.t4 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X26 source.t17 minus.t12 drain_right.t3 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X27 source.t20 minus.t13 drain_right.t2 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X28 drain_left.t5 plus.t10 source.t13 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X29 source.t21 minus.t14 drain_right.t1 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X30 source.t0 plus.t11 drain_left.t4 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X31 drain_right.t0 minus.t15 source.t27 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X32 drain_left.t3 plus.t12 source.t8 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X33 source.t10 plus.t13 drain_left.t2 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X34 drain_left.t1 plus.t14 source.t5 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X35 drain_left.t0 plus.t15 source.t7 a_n2210_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
R0 minus.n5 minus.t10 195.948
R1 minus.n27 minus.t14 195.948
R2 minus.n6 minus.t3 174.966
R3 minus.n8 minus.t6 174.966
R4 minus.n12 minus.t13 174.966
R5 minus.n13 minus.t5 174.966
R6 minus.n1 minus.t8 174.966
R7 minus.n19 minus.t1 174.966
R8 minus.n20 minus.t9 174.966
R9 minus.n28 minus.t0 174.966
R10 minus.n30 minus.t12 174.966
R11 minus.n34 minus.t15 174.966
R12 minus.n35 minus.t7 174.966
R13 minus.n23 minus.t2 174.966
R14 minus.n41 minus.t4 174.966
R15 minus.n42 minus.t11 174.966
R16 minus.n21 minus.n20 161.3
R17 minus.n19 minus.n0 161.3
R18 minus.n18 minus.n17 161.3
R19 minus.n16 minus.n1 161.3
R20 minus.n15 minus.n14 161.3
R21 minus.n13 minus.n2 161.3
R22 minus.n12 minus.n11 161.3
R23 minus.n10 minus.n3 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n43 minus.n42 161.3
R27 minus.n41 minus.n22 161.3
R28 minus.n40 minus.n39 161.3
R29 minus.n38 minus.n23 161.3
R30 minus.n37 minus.n36 161.3
R31 minus.n35 minus.n24 161.3
R32 minus.n34 minus.n33 161.3
R33 minus.n32 minus.n25 161.3
R34 minus.n31 minus.n30 161.3
R35 minus.n29 minus.n26 161.3
R36 minus.n5 minus.n4 70.4033
R37 minus.n27 minus.n26 70.4033
R38 minus.n13 minus.n12 48.2005
R39 minus.n20 minus.n19 48.2005
R40 minus.n35 minus.n34 48.2005
R41 minus.n42 minus.n41 48.2005
R42 minus.n8 minus.n7 37.246
R43 minus.n18 minus.n1 37.246
R44 minus.n30 minus.n29 37.246
R45 minus.n40 minus.n23 37.246
R46 minus.n8 minus.n3 35.7853
R47 minus.n14 minus.n1 35.7853
R48 minus.n30 minus.n25 35.7853
R49 minus.n36 minus.n23 35.7853
R50 minus.n44 minus.n21 29.9778
R51 minus.n6 minus.n5 20.9576
R52 minus.n28 minus.n27 20.9576
R53 minus.n12 minus.n3 12.4157
R54 minus.n14 minus.n13 12.4157
R55 minus.n34 minus.n25 12.4157
R56 minus.n36 minus.n35 12.4157
R57 minus.n7 minus.n6 10.955
R58 minus.n19 minus.n18 10.955
R59 minus.n29 minus.n28 10.955
R60 minus.n41 minus.n40 10.955
R61 minus.n44 minus.n43 6.56111
R62 minus.n21 minus.n0 0.189894
R63 minus.n17 minus.n0 0.189894
R64 minus.n17 minus.n16 0.189894
R65 minus.n16 minus.n15 0.189894
R66 minus.n15 minus.n2 0.189894
R67 minus.n11 minus.n2 0.189894
R68 minus.n11 minus.n10 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n31 minus.n26 0.189894
R72 minus.n32 minus.n31 0.189894
R73 minus.n33 minus.n32 0.189894
R74 minus.n33 minus.n24 0.189894
R75 minus.n37 minus.n24 0.189894
R76 minus.n38 minus.n37 0.189894
R77 minus.n39 minus.n38 0.189894
R78 minus.n39 minus.n22 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 source.n82 source.n80 289.615
R82 source.n68 source.n66 289.615
R83 source.n60 source.n58 289.615
R84 source.n46 source.n44 289.615
R85 source.n2 source.n0 289.615
R86 source.n16 source.n14 289.615
R87 source.n24 source.n22 289.615
R88 source.n38 source.n36 289.615
R89 source.n83 source.n82 185
R90 source.n69 source.n68 185
R91 source.n61 source.n60 185
R92 source.n47 source.n46 185
R93 source.n3 source.n2 185
R94 source.n17 source.n16 185
R95 source.n25 source.n24 185
R96 source.n39 source.n38 185
R97 source.t18 source.n81 167.117
R98 source.t21 source.n67 167.117
R99 source.t5 source.n59 167.117
R100 source.t11 source.n45 167.117
R101 source.t8 source.n1 167.117
R102 source.t14 source.n15 167.117
R103 source.t22 source.n23 167.117
R104 source.t31 source.n37 167.117
R105 source.n9 source.n8 84.1169
R106 source.n11 source.n10 84.1169
R107 source.n13 source.n12 84.1169
R108 source.n31 source.n30 84.1169
R109 source.n33 source.n32 84.1169
R110 source.n35 source.n34 84.1169
R111 source.n79 source.n78 84.1168
R112 source.n77 source.n76 84.1168
R113 source.n75 source.n74 84.1168
R114 source.n57 source.n56 84.1168
R115 source.n55 source.n54 84.1168
R116 source.n53 source.n52 84.1168
R117 source.n82 source.t18 52.3082
R118 source.n68 source.t21 52.3082
R119 source.n60 source.t5 52.3082
R120 source.n46 source.t11 52.3082
R121 source.n2 source.t8 52.3082
R122 source.n16 source.t14 52.3082
R123 source.n24 source.t22 52.3082
R124 source.n38 source.t31 52.3082
R125 source.n87 source.n86 31.4096
R126 source.n73 source.n72 31.4096
R127 source.n65 source.n64 31.4096
R128 source.n51 source.n50 31.4096
R129 source.n7 source.n6 31.4096
R130 source.n21 source.n20 31.4096
R131 source.n29 source.n28 31.4096
R132 source.n43 source.n42 31.4096
R133 source.n51 source.n43 14.4275
R134 source.n78 source.t19 9.9005
R135 source.n78 source.t24 9.9005
R136 source.n76 source.t27 9.9005
R137 source.n76 source.t25 9.9005
R138 source.n74 source.t26 9.9005
R139 source.n74 source.t17 9.9005
R140 source.n56 source.t13 9.9005
R141 source.n56 source.t2 9.9005
R142 source.n54 source.t12 9.9005
R143 source.n54 source.t15 9.9005
R144 source.n52 source.t3 9.9005
R145 source.n52 source.t6 9.9005
R146 source.n8 source.t7 9.9005
R147 source.n8 source.t1 9.9005
R148 source.n10 source.t9 9.9005
R149 source.n10 source.t0 9.9005
R150 source.n12 source.t4 9.9005
R151 source.n12 source.t10 9.9005
R152 source.n30 source.t23 9.9005
R153 source.n30 source.t30 9.9005
R154 source.n32 source.t29 9.9005
R155 source.n32 source.t20 9.9005
R156 source.n34 source.t28 9.9005
R157 source.n34 source.t16 9.9005
R158 source.n83 source.n81 9.71174
R159 source.n69 source.n67 9.71174
R160 source.n61 source.n59 9.71174
R161 source.n47 source.n45 9.71174
R162 source.n3 source.n1 9.71174
R163 source.n17 source.n15 9.71174
R164 source.n25 source.n23 9.71174
R165 source.n39 source.n37 9.71174
R166 source.n86 source.n85 9.45567
R167 source.n72 source.n71 9.45567
R168 source.n64 source.n63 9.45567
R169 source.n50 source.n49 9.45567
R170 source.n6 source.n5 9.45567
R171 source.n20 source.n19 9.45567
R172 source.n28 source.n27 9.45567
R173 source.n42 source.n41 9.45567
R174 source.n85 source.n84 9.3005
R175 source.n71 source.n70 9.3005
R176 source.n63 source.n62 9.3005
R177 source.n49 source.n48 9.3005
R178 source.n5 source.n4 9.3005
R179 source.n19 source.n18 9.3005
R180 source.n27 source.n26 9.3005
R181 source.n41 source.n40 9.3005
R182 source.n88 source.n7 8.8068
R183 source.n86 source.n80 8.14595
R184 source.n72 source.n66 8.14595
R185 source.n64 source.n58 8.14595
R186 source.n50 source.n44 8.14595
R187 source.n6 source.n0 8.14595
R188 source.n20 source.n14 8.14595
R189 source.n28 source.n22 8.14595
R190 source.n42 source.n36 8.14595
R191 source.n84 source.n83 7.3702
R192 source.n70 source.n69 7.3702
R193 source.n62 source.n61 7.3702
R194 source.n48 source.n47 7.3702
R195 source.n4 source.n3 7.3702
R196 source.n18 source.n17 7.3702
R197 source.n26 source.n25 7.3702
R198 source.n40 source.n39 7.3702
R199 source.n84 source.n80 5.81868
R200 source.n70 source.n66 5.81868
R201 source.n62 source.n58 5.81868
R202 source.n48 source.n44 5.81868
R203 source.n4 source.n0 5.81868
R204 source.n18 source.n14 5.81868
R205 source.n26 source.n22 5.81868
R206 source.n40 source.n36 5.81868
R207 source.n88 source.n87 5.62119
R208 source.n85 source.n81 3.44771
R209 source.n71 source.n67 3.44771
R210 source.n63 source.n59 3.44771
R211 source.n49 source.n45 3.44771
R212 source.n5 source.n1 3.44771
R213 source.n19 source.n15 3.44771
R214 source.n27 source.n23 3.44771
R215 source.n41 source.n37 3.44771
R216 source.n43 source.n35 0.716017
R217 source.n35 source.n33 0.716017
R218 source.n33 source.n31 0.716017
R219 source.n31 source.n29 0.716017
R220 source.n21 source.n13 0.716017
R221 source.n13 source.n11 0.716017
R222 source.n11 source.n9 0.716017
R223 source.n9 source.n7 0.716017
R224 source.n53 source.n51 0.716017
R225 source.n55 source.n53 0.716017
R226 source.n57 source.n55 0.716017
R227 source.n65 source.n57 0.716017
R228 source.n75 source.n73 0.716017
R229 source.n77 source.n75 0.716017
R230 source.n79 source.n77 0.716017
R231 source.n87 source.n79 0.716017
R232 source.n29 source.n21 0.470328
R233 source.n73 source.n65 0.470328
R234 source source.n88 0.188
R235 drain_right.n9 drain_right.n7 101.511
R236 drain_right.n5 drain_right.n3 101.511
R237 drain_right.n2 drain_right.n0 101.511
R238 drain_right.n9 drain_right.n8 100.796
R239 drain_right.n11 drain_right.n10 100.796
R240 drain_right.n13 drain_right.n12 100.796
R241 drain_right.n5 drain_right.n4 100.796
R242 drain_right.n2 drain_right.n1 100.796
R243 drain_right drain_right.n6 23.8889
R244 drain_right.n3 drain_right.t11 9.9005
R245 drain_right.n3 drain_right.t4 9.9005
R246 drain_right.n4 drain_right.t8 9.9005
R247 drain_right.n4 drain_right.t13 9.9005
R248 drain_right.n1 drain_right.t3 9.9005
R249 drain_right.n1 drain_right.t0 9.9005
R250 drain_right.n0 drain_right.t1 9.9005
R251 drain_right.n0 drain_right.t15 9.9005
R252 drain_right.n7 drain_right.t12 9.9005
R253 drain_right.n7 drain_right.t5 9.9005
R254 drain_right.n8 drain_right.t2 9.9005
R255 drain_right.n8 drain_right.t9 9.9005
R256 drain_right.n10 drain_right.t7 9.9005
R257 drain_right.n10 drain_right.t10 9.9005
R258 drain_right.n12 drain_right.t6 9.9005
R259 drain_right.n12 drain_right.t14 9.9005
R260 drain_right drain_right.n13 6.36873
R261 drain_right.n13 drain_right.n11 0.716017
R262 drain_right.n11 drain_right.n9 0.716017
R263 drain_right.n6 drain_right.n5 0.302913
R264 drain_right.n6 drain_right.n2 0.302913
R265 plus.n5 plus.t2 195.948
R266 plus.n27 plus.t14 195.948
R267 plus.n20 plus.t12 174.966
R268 plus.n19 plus.t7 174.966
R269 plus.n1 plus.t15 174.966
R270 plus.n13 plus.t11 174.966
R271 plus.n12 plus.t5 174.966
R272 plus.n4 plus.t13 174.966
R273 plus.n6 plus.t9 174.966
R274 plus.n42 plus.t8 174.966
R275 plus.n41 plus.t4 174.966
R276 plus.n23 plus.t0 174.966
R277 plus.n35 plus.t6 174.966
R278 plus.n34 plus.t3 174.966
R279 plus.n26 plus.t10 174.966
R280 plus.n28 plus.t1 174.966
R281 plus.n8 plus.n7 161.3
R282 plus.n9 plus.n4 161.3
R283 plus.n11 plus.n10 161.3
R284 plus.n12 plus.n3 161.3
R285 plus.n13 plus.n2 161.3
R286 plus.n15 plus.n14 161.3
R287 plus.n16 plus.n1 161.3
R288 plus.n18 plus.n17 161.3
R289 plus.n19 plus.n0 161.3
R290 plus.n21 plus.n20 161.3
R291 plus.n30 plus.n29 161.3
R292 plus.n31 plus.n26 161.3
R293 plus.n33 plus.n32 161.3
R294 plus.n34 plus.n25 161.3
R295 plus.n35 plus.n24 161.3
R296 plus.n37 plus.n36 161.3
R297 plus.n38 plus.n23 161.3
R298 plus.n40 plus.n39 161.3
R299 plus.n41 plus.n22 161.3
R300 plus.n43 plus.n42 161.3
R301 plus.n8 plus.n5 70.4033
R302 plus.n30 plus.n27 70.4033
R303 plus.n20 plus.n19 48.2005
R304 plus.n13 plus.n12 48.2005
R305 plus.n42 plus.n41 48.2005
R306 plus.n35 plus.n34 48.2005
R307 plus.n18 plus.n1 37.246
R308 plus.n7 plus.n4 37.246
R309 plus.n40 plus.n23 37.246
R310 plus.n29 plus.n26 37.246
R311 plus.n14 plus.n1 35.7853
R312 plus.n11 plus.n4 35.7853
R313 plus.n36 plus.n23 35.7853
R314 plus.n33 plus.n26 35.7853
R315 plus plus.n43 27.6467
R316 plus.n6 plus.n5 20.9576
R317 plus.n28 plus.n27 20.9576
R318 plus.n14 plus.n13 12.4157
R319 plus.n12 plus.n11 12.4157
R320 plus.n36 plus.n35 12.4157
R321 plus.n34 plus.n33 12.4157
R322 plus.n19 plus.n18 10.955
R323 plus.n7 plus.n6 10.955
R324 plus.n41 plus.n40 10.955
R325 plus.n29 plus.n28 10.955
R326 plus plus.n21 8.41717
R327 plus.n9 plus.n8 0.189894
R328 plus.n10 plus.n9 0.189894
R329 plus.n10 plus.n3 0.189894
R330 plus.n3 plus.n2 0.189894
R331 plus.n15 plus.n2 0.189894
R332 plus.n16 plus.n15 0.189894
R333 plus.n17 plus.n16 0.189894
R334 plus.n17 plus.n0 0.189894
R335 plus.n21 plus.n0 0.189894
R336 plus.n43 plus.n22 0.189894
R337 plus.n39 plus.n22 0.189894
R338 plus.n39 plus.n38 0.189894
R339 plus.n38 plus.n37 0.189894
R340 plus.n37 plus.n24 0.189894
R341 plus.n25 plus.n24 0.189894
R342 plus.n32 plus.n25 0.189894
R343 plus.n32 plus.n31 0.189894
R344 plus.n31 plus.n30 0.189894
R345 drain_left.n9 drain_left.n7 101.511
R346 drain_left.n5 drain_left.n3 101.511
R347 drain_left.n2 drain_left.n0 101.511
R348 drain_left.n13 drain_left.n12 100.796
R349 drain_left.n11 drain_left.n10 100.796
R350 drain_left.n9 drain_left.n8 100.796
R351 drain_left.n5 drain_left.n4 100.796
R352 drain_left.n2 drain_left.n1 100.796
R353 drain_left drain_left.n6 24.4422
R354 drain_left.n3 drain_left.t14 9.9005
R355 drain_left.n3 drain_left.t1 9.9005
R356 drain_left.n4 drain_left.t12 9.9005
R357 drain_left.n4 drain_left.t5 9.9005
R358 drain_left.n1 drain_left.t15 9.9005
R359 drain_left.n1 drain_left.t9 9.9005
R360 drain_left.n0 drain_left.t7 9.9005
R361 drain_left.n0 drain_left.t11 9.9005
R362 drain_left.n12 drain_left.t8 9.9005
R363 drain_left.n12 drain_left.t3 9.9005
R364 drain_left.n10 drain_left.t4 9.9005
R365 drain_left.n10 drain_left.t0 9.9005
R366 drain_left.n8 drain_left.t2 9.9005
R367 drain_left.n8 drain_left.t10 9.9005
R368 drain_left.n7 drain_left.t13 9.9005
R369 drain_left.n7 drain_left.t6 9.9005
R370 drain_left drain_left.n13 6.36873
R371 drain_left.n11 drain_left.n9 0.716017
R372 drain_left.n13 drain_left.n11 0.716017
R373 drain_left.n6 drain_left.n5 0.302913
R374 drain_left.n6 drain_left.n2 0.302913
C0 minus drain_left 0.178338f
C1 plus source 2.27177f
C2 source drain_right 6.52188f
C3 plus drain_right 0.379534f
C4 drain_left source 6.52068f
C5 plus drain_left 2.07241f
C6 drain_left drain_right 1.15071f
C7 minus source 2.2578f
C8 plus minus 4.06267f
C9 minus drain_right 1.85533f
C10 drain_right a_n2210_n1288# 4.10513f
C11 drain_left a_n2210_n1288# 4.80744f
C12 source a_n2210_n1288# 3.248483f
C13 minus a_n2210_n1288# 7.925713f
C14 plus a_n2210_n1288# 9.247581f
C15 drain_left.t7 a_n2210_n1288# 0.044906f
C16 drain_left.t11 a_n2210_n1288# 0.044906f
C17 drain_left.n0 a_n2210_n1288# 0.284648f
C18 drain_left.t15 a_n2210_n1288# 0.044906f
C19 drain_left.t9 a_n2210_n1288# 0.044906f
C20 drain_left.n1 a_n2210_n1288# 0.282111f
C21 drain_left.n2 a_n2210_n1288# 0.670237f
C22 drain_left.t14 a_n2210_n1288# 0.044906f
C23 drain_left.t1 a_n2210_n1288# 0.044906f
C24 drain_left.n3 a_n2210_n1288# 0.284648f
C25 drain_left.t12 a_n2210_n1288# 0.044906f
C26 drain_left.t5 a_n2210_n1288# 0.044906f
C27 drain_left.n4 a_n2210_n1288# 0.282111f
C28 drain_left.n5 a_n2210_n1288# 0.670237f
C29 drain_left.n6 a_n2210_n1288# 0.926404f
C30 drain_left.t13 a_n2210_n1288# 0.044906f
C31 drain_left.t6 a_n2210_n1288# 0.044906f
C32 drain_left.n7 a_n2210_n1288# 0.284649f
C33 drain_left.t2 a_n2210_n1288# 0.044906f
C34 drain_left.t10 a_n2210_n1288# 0.044906f
C35 drain_left.n8 a_n2210_n1288# 0.282112f
C36 drain_left.n9 a_n2210_n1288# 0.705878f
C37 drain_left.t4 a_n2210_n1288# 0.044906f
C38 drain_left.t0 a_n2210_n1288# 0.044906f
C39 drain_left.n10 a_n2210_n1288# 0.282112f
C40 drain_left.n11 a_n2210_n1288# 0.348485f
C41 drain_left.t8 a_n2210_n1288# 0.044906f
C42 drain_left.t3 a_n2210_n1288# 0.044906f
C43 drain_left.n12 a_n2210_n1288# 0.282112f
C44 drain_left.n13 a_n2210_n1288# 0.592593f
C45 plus.n0 a_n2210_n1288# 0.048947f
C46 plus.t12 a_n2210_n1288# 0.151576f
C47 plus.t7 a_n2210_n1288# 0.151576f
C48 plus.t15 a_n2210_n1288# 0.151576f
C49 plus.n1 a_n2210_n1288# 0.114316f
C50 plus.n2 a_n2210_n1288# 0.048947f
C51 plus.t11 a_n2210_n1288# 0.151576f
C52 plus.t5 a_n2210_n1288# 0.151576f
C53 plus.n3 a_n2210_n1288# 0.048947f
C54 plus.t13 a_n2210_n1288# 0.151576f
C55 plus.n4 a_n2210_n1288# 0.114316f
C56 plus.t2 a_n2210_n1288# 0.163275f
C57 plus.n5 a_n2210_n1288# 0.097844f
C58 plus.t9 a_n2210_n1288# 0.151576f
C59 plus.n6 a_n2210_n1288# 0.111449f
C60 plus.n7 a_n2210_n1288# 0.011107f
C61 plus.n8 a_n2210_n1288# 0.15584f
C62 plus.n9 a_n2210_n1288# 0.048947f
C63 plus.n10 a_n2210_n1288# 0.048947f
C64 plus.n11 a_n2210_n1288# 0.011107f
C65 plus.n12 a_n2210_n1288# 0.111751f
C66 plus.n13 a_n2210_n1288# 0.111751f
C67 plus.n14 a_n2210_n1288# 0.011107f
C68 plus.n15 a_n2210_n1288# 0.048947f
C69 plus.n16 a_n2210_n1288# 0.048947f
C70 plus.n17 a_n2210_n1288# 0.048947f
C71 plus.n18 a_n2210_n1288# 0.011107f
C72 plus.n19 a_n2210_n1288# 0.111449f
C73 plus.n20 a_n2210_n1288# 0.109186f
C74 plus.n21 a_n2210_n1288# 0.357326f
C75 plus.n22 a_n2210_n1288# 0.048947f
C76 plus.t8 a_n2210_n1288# 0.151576f
C77 plus.t4 a_n2210_n1288# 0.151576f
C78 plus.t0 a_n2210_n1288# 0.151576f
C79 plus.n23 a_n2210_n1288# 0.114316f
C80 plus.n24 a_n2210_n1288# 0.048947f
C81 plus.t6 a_n2210_n1288# 0.151576f
C82 plus.n25 a_n2210_n1288# 0.048947f
C83 plus.t3 a_n2210_n1288# 0.151576f
C84 plus.t10 a_n2210_n1288# 0.151576f
C85 plus.n26 a_n2210_n1288# 0.114316f
C86 plus.t14 a_n2210_n1288# 0.163275f
C87 plus.n27 a_n2210_n1288# 0.097844f
C88 plus.t1 a_n2210_n1288# 0.151576f
C89 plus.n28 a_n2210_n1288# 0.111449f
C90 plus.n29 a_n2210_n1288# 0.011107f
C91 plus.n30 a_n2210_n1288# 0.15584f
C92 plus.n31 a_n2210_n1288# 0.048947f
C93 plus.n32 a_n2210_n1288# 0.048947f
C94 plus.n33 a_n2210_n1288# 0.011107f
C95 plus.n34 a_n2210_n1288# 0.111751f
C96 plus.n35 a_n2210_n1288# 0.111751f
C97 plus.n36 a_n2210_n1288# 0.011107f
C98 plus.n37 a_n2210_n1288# 0.048947f
C99 plus.n38 a_n2210_n1288# 0.048947f
C100 plus.n39 a_n2210_n1288# 0.048947f
C101 plus.n40 a_n2210_n1288# 0.011107f
C102 plus.n41 a_n2210_n1288# 0.111449f
C103 plus.n42 a_n2210_n1288# 0.109186f
C104 plus.n43 a_n2210_n1288# 1.21403f
C105 drain_right.t1 a_n2210_n1288# 0.034385f
C106 drain_right.t15 a_n2210_n1288# 0.034385f
C107 drain_right.n0 a_n2210_n1288# 0.217958f
C108 drain_right.t3 a_n2210_n1288# 0.034385f
C109 drain_right.t0 a_n2210_n1288# 0.034385f
C110 drain_right.n1 a_n2210_n1288# 0.216015f
C111 drain_right.n2 a_n2210_n1288# 0.513207f
C112 drain_right.t11 a_n2210_n1288# 0.034385f
C113 drain_right.t4 a_n2210_n1288# 0.034385f
C114 drain_right.n3 a_n2210_n1288# 0.217958f
C115 drain_right.t8 a_n2210_n1288# 0.034385f
C116 drain_right.t13 a_n2210_n1288# 0.034385f
C117 drain_right.n4 a_n2210_n1288# 0.216015f
C118 drain_right.n5 a_n2210_n1288# 0.513207f
C119 drain_right.n6 a_n2210_n1288# 0.666887f
C120 drain_right.t12 a_n2210_n1288# 0.034385f
C121 drain_right.t5 a_n2210_n1288# 0.034385f
C122 drain_right.n7 a_n2210_n1288# 0.217959f
C123 drain_right.t2 a_n2210_n1288# 0.034385f
C124 drain_right.t9 a_n2210_n1288# 0.034385f
C125 drain_right.n8 a_n2210_n1288# 0.216016f
C126 drain_right.n9 a_n2210_n1288# 0.540498f
C127 drain_right.t7 a_n2210_n1288# 0.034385f
C128 drain_right.t10 a_n2210_n1288# 0.034385f
C129 drain_right.n10 a_n2210_n1288# 0.216016f
C130 drain_right.n11 a_n2210_n1288# 0.266839f
C131 drain_right.t6 a_n2210_n1288# 0.034385f
C132 drain_right.t14 a_n2210_n1288# 0.034385f
C133 drain_right.n12 a_n2210_n1288# 0.216016f
C134 drain_right.n13 a_n2210_n1288# 0.453754f
C135 source.n0 a_n2210_n1288# 0.045168f
C136 source.n1 a_n2210_n1288# 0.099939f
C137 source.t8 a_n2210_n1288# 0.074999f
C138 source.n2 a_n2210_n1288# 0.078217f
C139 source.n3 a_n2210_n1288# 0.025214f
C140 source.n4 a_n2210_n1288# 0.016629f
C141 source.n5 a_n2210_n1288# 0.220291f
C142 source.n6 a_n2210_n1288# 0.049514f
C143 source.n7 a_n2210_n1288# 0.497743f
C144 source.t7 a_n2210_n1288# 0.048909f
C145 source.t1 a_n2210_n1288# 0.048909f
C146 source.n8 a_n2210_n1288# 0.261467f
C147 source.n9 a_n2210_n1288# 0.383289f
C148 source.t9 a_n2210_n1288# 0.048909f
C149 source.t0 a_n2210_n1288# 0.048909f
C150 source.n10 a_n2210_n1288# 0.261467f
C151 source.n11 a_n2210_n1288# 0.383289f
C152 source.t4 a_n2210_n1288# 0.048909f
C153 source.t10 a_n2210_n1288# 0.048909f
C154 source.n12 a_n2210_n1288# 0.261467f
C155 source.n13 a_n2210_n1288# 0.383289f
C156 source.n14 a_n2210_n1288# 0.045168f
C157 source.n15 a_n2210_n1288# 0.099939f
C158 source.t14 a_n2210_n1288# 0.074999f
C159 source.n16 a_n2210_n1288# 0.078217f
C160 source.n17 a_n2210_n1288# 0.025214f
C161 source.n18 a_n2210_n1288# 0.016629f
C162 source.n19 a_n2210_n1288# 0.220291f
C163 source.n20 a_n2210_n1288# 0.049514f
C164 source.n21 a_n2210_n1288# 0.143673f
C165 source.n22 a_n2210_n1288# 0.045168f
C166 source.n23 a_n2210_n1288# 0.099939f
C167 source.t22 a_n2210_n1288# 0.074999f
C168 source.n24 a_n2210_n1288# 0.078217f
C169 source.n25 a_n2210_n1288# 0.025214f
C170 source.n26 a_n2210_n1288# 0.016629f
C171 source.n27 a_n2210_n1288# 0.220291f
C172 source.n28 a_n2210_n1288# 0.049514f
C173 source.n29 a_n2210_n1288# 0.143673f
C174 source.t23 a_n2210_n1288# 0.048909f
C175 source.t30 a_n2210_n1288# 0.048909f
C176 source.n30 a_n2210_n1288# 0.261467f
C177 source.n31 a_n2210_n1288# 0.383289f
C178 source.t29 a_n2210_n1288# 0.048909f
C179 source.t20 a_n2210_n1288# 0.048909f
C180 source.n32 a_n2210_n1288# 0.261467f
C181 source.n33 a_n2210_n1288# 0.383289f
C182 source.t28 a_n2210_n1288# 0.048909f
C183 source.t16 a_n2210_n1288# 0.048909f
C184 source.n34 a_n2210_n1288# 0.261467f
C185 source.n35 a_n2210_n1288# 0.383289f
C186 source.n36 a_n2210_n1288# 0.045168f
C187 source.n37 a_n2210_n1288# 0.099939f
C188 source.t31 a_n2210_n1288# 0.074999f
C189 source.n38 a_n2210_n1288# 0.078217f
C190 source.n39 a_n2210_n1288# 0.025214f
C191 source.n40 a_n2210_n1288# 0.016629f
C192 source.n41 a_n2210_n1288# 0.220291f
C193 source.n42 a_n2210_n1288# 0.049514f
C194 source.n43 a_n2210_n1288# 0.790134f
C195 source.n44 a_n2210_n1288# 0.045168f
C196 source.n45 a_n2210_n1288# 0.099939f
C197 source.t11 a_n2210_n1288# 0.074999f
C198 source.n46 a_n2210_n1288# 0.078217f
C199 source.n47 a_n2210_n1288# 0.025214f
C200 source.n48 a_n2210_n1288# 0.016629f
C201 source.n49 a_n2210_n1288# 0.220291f
C202 source.n50 a_n2210_n1288# 0.049514f
C203 source.n51 a_n2210_n1288# 0.790134f
C204 source.t3 a_n2210_n1288# 0.048909f
C205 source.t6 a_n2210_n1288# 0.048909f
C206 source.n52 a_n2210_n1288# 0.261466f
C207 source.n53 a_n2210_n1288# 0.38329f
C208 source.t12 a_n2210_n1288# 0.048909f
C209 source.t15 a_n2210_n1288# 0.048909f
C210 source.n54 a_n2210_n1288# 0.261466f
C211 source.n55 a_n2210_n1288# 0.38329f
C212 source.t13 a_n2210_n1288# 0.048909f
C213 source.t2 a_n2210_n1288# 0.048909f
C214 source.n56 a_n2210_n1288# 0.261466f
C215 source.n57 a_n2210_n1288# 0.38329f
C216 source.n58 a_n2210_n1288# 0.045168f
C217 source.n59 a_n2210_n1288# 0.099939f
C218 source.t5 a_n2210_n1288# 0.074999f
C219 source.n60 a_n2210_n1288# 0.078217f
C220 source.n61 a_n2210_n1288# 0.025214f
C221 source.n62 a_n2210_n1288# 0.016629f
C222 source.n63 a_n2210_n1288# 0.220291f
C223 source.n64 a_n2210_n1288# 0.049514f
C224 source.n65 a_n2210_n1288# 0.143673f
C225 source.n66 a_n2210_n1288# 0.045168f
C226 source.n67 a_n2210_n1288# 0.099939f
C227 source.t21 a_n2210_n1288# 0.074999f
C228 source.n68 a_n2210_n1288# 0.078217f
C229 source.n69 a_n2210_n1288# 0.025214f
C230 source.n70 a_n2210_n1288# 0.016629f
C231 source.n71 a_n2210_n1288# 0.220291f
C232 source.n72 a_n2210_n1288# 0.049514f
C233 source.n73 a_n2210_n1288# 0.143673f
C234 source.t26 a_n2210_n1288# 0.048909f
C235 source.t17 a_n2210_n1288# 0.048909f
C236 source.n74 a_n2210_n1288# 0.261466f
C237 source.n75 a_n2210_n1288# 0.38329f
C238 source.t27 a_n2210_n1288# 0.048909f
C239 source.t25 a_n2210_n1288# 0.048909f
C240 source.n76 a_n2210_n1288# 0.261466f
C241 source.n77 a_n2210_n1288# 0.38329f
C242 source.t19 a_n2210_n1288# 0.048909f
C243 source.t24 a_n2210_n1288# 0.048909f
C244 source.n78 a_n2210_n1288# 0.261466f
C245 source.n79 a_n2210_n1288# 0.38329f
C246 source.n80 a_n2210_n1288# 0.045168f
C247 source.n81 a_n2210_n1288# 0.099939f
C248 source.t18 a_n2210_n1288# 0.074999f
C249 source.n82 a_n2210_n1288# 0.078217f
C250 source.n83 a_n2210_n1288# 0.025214f
C251 source.n84 a_n2210_n1288# 0.016629f
C252 source.n85 a_n2210_n1288# 0.220291f
C253 source.n86 a_n2210_n1288# 0.049514f
C254 source.n87 a_n2210_n1288# 0.332027f
C255 source.n88 a_n2210_n1288# 0.772509f
C256 minus.n0 a_n2210_n1288# 0.03643f
C257 minus.t8 a_n2210_n1288# 0.112814f
C258 minus.n1 a_n2210_n1288# 0.085083f
C259 minus.n2 a_n2210_n1288# 0.03643f
C260 minus.n3 a_n2210_n1288# 0.008267f
C261 minus.t13 a_n2210_n1288# 0.112814f
C262 minus.n4 a_n2210_n1288# 0.115988f
C263 minus.t3 a_n2210_n1288# 0.112814f
C264 minus.t10 a_n2210_n1288# 0.121521f
C265 minus.n5 a_n2210_n1288# 0.072823f
C266 minus.n6 a_n2210_n1288# 0.082949f
C267 minus.n7 a_n2210_n1288# 0.008267f
C268 minus.t6 a_n2210_n1288# 0.112814f
C269 minus.n8 a_n2210_n1288# 0.085083f
C270 minus.n9 a_n2210_n1288# 0.03643f
C271 minus.n10 a_n2210_n1288# 0.03643f
C272 minus.n11 a_n2210_n1288# 0.03643f
C273 minus.n12 a_n2210_n1288# 0.083173f
C274 minus.t5 a_n2210_n1288# 0.112814f
C275 minus.n13 a_n2210_n1288# 0.083173f
C276 minus.n14 a_n2210_n1288# 0.008267f
C277 minus.n15 a_n2210_n1288# 0.03643f
C278 minus.n16 a_n2210_n1288# 0.03643f
C279 minus.n17 a_n2210_n1288# 0.03643f
C280 minus.n18 a_n2210_n1288# 0.008267f
C281 minus.t1 a_n2210_n1288# 0.112814f
C282 minus.n19 a_n2210_n1288# 0.082949f
C283 minus.t9 a_n2210_n1288# 0.112814f
C284 minus.n20 a_n2210_n1288# 0.081264f
C285 minus.n21 a_n2210_n1288# 0.948577f
C286 minus.n22 a_n2210_n1288# 0.03643f
C287 minus.t2 a_n2210_n1288# 0.112814f
C288 minus.n23 a_n2210_n1288# 0.085083f
C289 minus.n24 a_n2210_n1288# 0.03643f
C290 minus.n25 a_n2210_n1288# 0.008267f
C291 minus.n26 a_n2210_n1288# 0.115988f
C292 minus.t14 a_n2210_n1288# 0.121521f
C293 minus.n27 a_n2210_n1288# 0.072823f
C294 minus.t0 a_n2210_n1288# 0.112814f
C295 minus.n28 a_n2210_n1288# 0.082949f
C296 minus.n29 a_n2210_n1288# 0.008267f
C297 minus.t12 a_n2210_n1288# 0.112814f
C298 minus.n30 a_n2210_n1288# 0.085083f
C299 minus.n31 a_n2210_n1288# 0.03643f
C300 minus.n32 a_n2210_n1288# 0.03643f
C301 minus.n33 a_n2210_n1288# 0.03643f
C302 minus.t15 a_n2210_n1288# 0.112814f
C303 minus.n34 a_n2210_n1288# 0.083173f
C304 minus.t7 a_n2210_n1288# 0.112814f
C305 minus.n35 a_n2210_n1288# 0.083173f
C306 minus.n36 a_n2210_n1288# 0.008267f
C307 minus.n37 a_n2210_n1288# 0.03643f
C308 minus.n38 a_n2210_n1288# 0.03643f
C309 minus.n39 a_n2210_n1288# 0.03643f
C310 minus.n40 a_n2210_n1288# 0.008267f
C311 minus.t4 a_n2210_n1288# 0.112814f
C312 minus.n41 a_n2210_n1288# 0.082949f
C313 minus.t11 a_n2210_n1288# 0.112814f
C314 minus.n42 a_n2210_n1288# 0.081264f
C315 minus.n43 a_n2210_n1288# 0.243401f
C316 minus.n44 a_n2210_n1288# 1.16767f
.ends

