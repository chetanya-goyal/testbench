* NGSPICE file created from diffpair173.ext - technology: sky130A

.subckt diffpair173 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t9 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X1 drain_right.t7 minus.t0 source.t1 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X2 a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X3 a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X4 drain_right.t6 minus.t1 source.t14 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X5 drain_left.t6 plus.t1 source.t8 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X6 source.t4 minus.t2 drain_right.t5 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X7 a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X8 drain_left.t5 plus.t2 source.t6 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X9 source.t0 minus.t3 drain_right.t4 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X10 source.t13 plus.t3 drain_left.t4 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X11 drain_right.t3 minus.t4 source.t15 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X12 source.t12 plus.t4 drain_left.t3 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X13 source.t11 plus.t5 drain_left.t2 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X14 drain_right.t2 minus.t5 source.t2 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X15 drain_left.t1 plus.t6 source.t10 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X16 source.t3 minus.t6 drain_right.t1 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X17 a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X18 source.t7 plus.t7 drain_left.t0 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X19 source.t5 minus.t7 drain_right.t0 a_n1246_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n1 plus.t3 561.239
R1 plus.n5 plus.t6 561.239
R2 plus.n8 plus.t2 561.239
R3 plus.n12 plus.t4 561.239
R4 plus.n2 plus.t1 518.15
R5 plus.n4 plus.t7 518.15
R6 plus.n9 plus.t5 518.15
R7 plus.n11 plus.t0 518.15
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 38.7066
R15 plus.n4 plus.n3 38.7066
R16 plus.n11 plus.n10 38.7066
R17 plus.n10 plus.n9 38.7066
R18 plus.n2 plus.n1 34.3247
R19 plus.n5 plus.n4 34.3247
R20 plus.n12 plus.n11 34.3247
R21 plus.n9 plus.n8 34.3247
R22 plus plus.n13 24.2566
R23 plus plus.n6 8.67853
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n0 source.t10 69.6943
R27 source.n3 source.t13 69.6943
R28 source.n4 source.t2 69.6943
R29 source.n7 source.t3 69.6943
R30 source.n15 source.t14 69.6942
R31 source.n12 source.t4 69.6942
R32 source.n11 source.t6 69.6942
R33 source.n8 source.t12 69.6942
R34 source.n2 source.n1 63.0943
R35 source.n6 source.n5 63.0943
R36 source.n14 source.n13 63.0942
R37 source.n10 source.n9 63.0942
R38 source.n8 source.n7 14.9264
R39 source.n16 source.n0 9.43506
R40 source.n13 source.t15 6.6005
R41 source.n13 source.t5 6.6005
R42 source.n9 source.t9 6.6005
R43 source.n9 source.t11 6.6005
R44 source.n1 source.t8 6.6005
R45 source.n1 source.t7 6.6005
R46 source.n5 source.t1 6.6005
R47 source.n5 source.t0 6.6005
R48 source.n16 source.n15 5.49188
R49 source.n4 source.n3 0.470328
R50 source.n12 source.n11 0.470328
R51 source.n7 source.n6 0.457397
R52 source.n6 source.n4 0.457397
R53 source.n3 source.n2 0.457397
R54 source.n2 source.n0 0.457397
R55 source.n10 source.n8 0.457397
R56 source.n11 source.n10 0.457397
R57 source.n14 source.n12 0.457397
R58 source.n15 source.n14 0.457397
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 80.23
R61 drain_left.n2 drain_left.n1 79.9461
R62 drain_left.n2 drain_left.n0 79.9461
R63 drain_left.n5 drain_left.n4 79.7731
R64 drain_left drain_left.n2 22.148
R65 drain_left.n1 drain_left.t2 6.6005
R66 drain_left.n1 drain_left.t5 6.6005
R67 drain_left.n0 drain_left.t3 6.6005
R68 drain_left.n0 drain_left.t7 6.6005
R69 drain_left.n4 drain_left.t0 6.6005
R70 drain_left.n4 drain_left.t1 6.6005
R71 drain_left.n3 drain_left.t4 6.6005
R72 drain_left.n3 drain_left.t6 6.6005
R73 drain_left drain_left.n5 6.11011
R74 minus.n5 minus.t6 561.239
R75 minus.n1 minus.t5 561.239
R76 minus.n12 minus.t1 561.239
R77 minus.n8 minus.t2 561.239
R78 minus.n4 minus.t0 518.15
R79 minus.n2 minus.t3 518.15
R80 minus.n11 minus.t7 518.15
R81 minus.n9 minus.t4 518.15
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 38.7066
R89 minus.n3 minus.n2 38.7066
R90 minus.n10 minus.n9 38.7066
R91 minus.n11 minus.n10 38.7066
R92 minus.n5 minus.n4 34.3247
R93 minus.n2 minus.n1 34.3247
R94 minus.n9 minus.n8 34.3247
R95 minus.n12 minus.n11 34.3247
R96 minus.n14 minus.n6 26.9664
R97 minus.n14 minus.n13 6.44368
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 80.23
R102 drain_right.n2 drain_right.n1 79.9461
R103 drain_right.n2 drain_right.n0 79.9461
R104 drain_right.n5 drain_right.n4 79.7731
R105 drain_right drain_right.n2 21.5948
R106 drain_right.n1 drain_right.t0 6.6005
R107 drain_right.n1 drain_right.t6 6.6005
R108 drain_right.n0 drain_right.t5 6.6005
R109 drain_right.n0 drain_right.t3 6.6005
R110 drain_right.n3 drain_right.t4 6.6005
R111 drain_right.n3 drain_right.t2 6.6005
R112 drain_right.n4 drain_right.t1 6.6005
R113 drain_right.n4 drain_right.t7 6.6005
R114 drain_right drain_right.n5 6.11011
C0 drain_left minus 0.175091f
C1 source plus 0.893519f
C2 source minus 0.879521f
C3 minus plus 3.04816f
C4 drain_right drain_left 0.58123f
C5 drain_right source 6.23565f
C6 drain_right plus 0.275117f
C7 drain_right minus 0.918078f
C8 source drain_left 6.23707f
C9 drain_left plus 1.03489f
C10 drain_right a_n1246_n1488# 3.4243f
C11 drain_left a_n1246_n1488# 3.58316f
C12 source a_n1246_n1488# 3.394763f
C13 minus a_n1246_n1488# 4.086458f
C14 plus a_n1246_n1488# 4.84625f
C15 drain_right.t5 a_n1246_n1488# 0.069038f
C16 drain_right.t3 a_n1246_n1488# 0.069038f
C17 drain_right.n0 a_n1246_n1488# 0.498563f
C18 drain_right.t0 a_n1246_n1488# 0.069038f
C19 drain_right.t6 a_n1246_n1488# 0.069038f
C20 drain_right.n1 a_n1246_n1488# 0.498563f
C21 drain_right.n2 a_n1246_n1488# 1.25668f
C22 drain_right.t4 a_n1246_n1488# 0.069038f
C23 drain_right.t2 a_n1246_n1488# 0.069038f
C24 drain_right.n3 a_n1246_n1488# 0.499782f
C25 drain_right.t1 a_n1246_n1488# 0.069038f
C26 drain_right.t7 a_n1246_n1488# 0.069038f
C27 drain_right.n4 a_n1246_n1488# 0.497899f
C28 drain_right.n5 a_n1246_n1488# 0.885896f
C29 minus.n0 a_n1246_n1488# 0.07732f
C30 minus.t6 a_n1246_n1488# 0.064722f
C31 minus.t0 a_n1246_n1488# 0.0617f
C32 minus.t3 a_n1246_n1488# 0.0617f
C33 minus.t5 a_n1246_n1488# 0.064722f
C34 minus.n1 a_n1246_n1488# 0.048829f
C35 minus.n2 a_n1246_n1488# 0.039475f
C36 minus.n3 a_n1246_n1488# 0.012437f
C37 minus.n4 a_n1246_n1488# 0.039475f
C38 minus.n5 a_n1246_n1488# 0.04878f
C39 minus.n6 a_n1246_n1488# 0.763972f
C40 minus.n7 a_n1246_n1488# 0.07732f
C41 minus.t7 a_n1246_n1488# 0.0617f
C42 minus.t4 a_n1246_n1488# 0.0617f
C43 minus.t2 a_n1246_n1488# 0.064722f
C44 minus.n8 a_n1246_n1488# 0.048829f
C45 minus.n9 a_n1246_n1488# 0.039475f
C46 minus.n10 a_n1246_n1488# 0.012437f
C47 minus.n11 a_n1246_n1488# 0.039475f
C48 minus.t1 a_n1246_n1488# 0.064722f
C49 minus.n12 a_n1246_n1488# 0.04878f
C50 minus.n13 a_n1246_n1488# 0.227431f
C51 minus.n14 a_n1246_n1488# 0.946964f
C52 drain_left.t3 a_n1246_n1488# 0.067793f
C53 drain_left.t7 a_n1246_n1488# 0.067793f
C54 drain_left.n0 a_n1246_n1488# 0.489568f
C55 drain_left.t2 a_n1246_n1488# 0.067793f
C56 drain_left.t5 a_n1246_n1488# 0.067793f
C57 drain_left.n1 a_n1246_n1488# 0.489568f
C58 drain_left.n2 a_n1246_n1488# 1.29111f
C59 drain_left.t4 a_n1246_n1488# 0.067793f
C60 drain_left.t6 a_n1246_n1488# 0.067793f
C61 drain_left.n3 a_n1246_n1488# 0.490765f
C62 drain_left.t0 a_n1246_n1488# 0.067793f
C63 drain_left.t1 a_n1246_n1488# 0.067793f
C64 drain_left.n4 a_n1246_n1488# 0.488916f
C65 drain_left.n5 a_n1246_n1488# 0.869912f
C66 source.t10 a_n1246_n1488# 0.501719f
C67 source.n0 a_n1246_n1488# 0.672036f
C68 source.t8 a_n1246_n1488# 0.06042f
C69 source.t7 a_n1246_n1488# 0.06042f
C70 source.n1 a_n1246_n1488# 0.383099f
C71 source.n2 a_n1246_n1488# 0.297062f
C72 source.t13 a_n1246_n1488# 0.501719f
C73 source.n3 a_n1246_n1488# 0.344287f
C74 source.t2 a_n1246_n1488# 0.501719f
C75 source.n4 a_n1246_n1488# 0.344287f
C76 source.t1 a_n1246_n1488# 0.06042f
C77 source.t0 a_n1246_n1488# 0.06042f
C78 source.n5 a_n1246_n1488# 0.383099f
C79 source.n6 a_n1246_n1488# 0.297062f
C80 source.t3 a_n1246_n1488# 0.501719f
C81 source.n7 a_n1246_n1488# 0.936015f
C82 source.t12 a_n1246_n1488# 0.501717f
C83 source.n8 a_n1246_n1488# 0.936017f
C84 source.t9 a_n1246_n1488# 0.06042f
C85 source.t11 a_n1246_n1488# 0.06042f
C86 source.n9 a_n1246_n1488# 0.383096f
C87 source.n10 a_n1246_n1488# 0.297065f
C88 source.t6 a_n1246_n1488# 0.501717f
C89 source.n11 a_n1246_n1488# 0.344289f
C90 source.t4 a_n1246_n1488# 0.501717f
C91 source.n12 a_n1246_n1488# 0.344289f
C92 source.t15 a_n1246_n1488# 0.06042f
C93 source.t5 a_n1246_n1488# 0.06042f
C94 source.n13 a_n1246_n1488# 0.383096f
C95 source.n14 a_n1246_n1488# 0.297065f
C96 source.t14 a_n1246_n1488# 0.501717f
C97 source.n15 a_n1246_n1488# 0.482484f
C98 source.n16 a_n1246_n1488# 0.73564f
C99 plus.n0 a_n1246_n1488# 0.079216f
C100 plus.t7 a_n1246_n1488# 0.063213f
C101 plus.t1 a_n1246_n1488# 0.063213f
C102 plus.t3 a_n1246_n1488# 0.066309f
C103 plus.n1 a_n1246_n1488# 0.050026f
C104 plus.n2 a_n1246_n1488# 0.040443f
C105 plus.n3 a_n1246_n1488# 0.012742f
C106 plus.n4 a_n1246_n1488# 0.040443f
C107 plus.t6 a_n1246_n1488# 0.066309f
C108 plus.n5 a_n1246_n1488# 0.049976f
C109 plus.n6 a_n1246_n1488# 0.26667f
C110 plus.n7 a_n1246_n1488# 0.079216f
C111 plus.t4 a_n1246_n1488# 0.066309f
C112 plus.t0 a_n1246_n1488# 0.063213f
C113 plus.t5 a_n1246_n1488# 0.063213f
C114 plus.t2 a_n1246_n1488# 0.066309f
C115 plus.n8 a_n1246_n1488# 0.050026f
C116 plus.n9 a_n1246_n1488# 0.040443f
C117 plus.n10 a_n1246_n1488# 0.012742f
C118 plus.n11 a_n1246_n1488# 0.040443f
C119 plus.n12 a_n1246_n1488# 0.049976f
C120 plus.n13 a_n1246_n1488# 0.740342f
.ends

