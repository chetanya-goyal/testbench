* NGSPICE file created from diffpair380.ext - technology: sky130A

.subckt diffpair380 minus drain_right drain_left source plus
X0 drain_right minus source a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.7
X1 a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X2 a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X3 drain_left plus source a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.7
X4 drain_right minus source a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.7
X5 drain_left plus source a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.7
X6 a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X7 a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# a_n1128_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
.ends

