* NGSPICE file created from diffpair337.ext - technology: sky130A

.subckt diffpair337 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t4 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 source.t30 minus.t1 drain_right.t13 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 drain_right.t6 minus.t2 source.t29 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X3 drain_right.t15 minus.t3 source.t28 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 drain_right.t8 minus.t4 source.t27 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 drain_right.t1 minus.t5 source.t26 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X6 drain_right.t2 minus.t6 source.t25 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X7 a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X8 drain_right.t7 minus.t7 source.t24 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X9 a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X10 source.t4 plus.t0 drain_left.t15 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X11 drain_left.t14 plus.t1 source.t15 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X12 source.t23 minus.t8 drain_right.t5 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X13 source.t22 minus.t9 drain_right.t14 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X14 source.t21 minus.t10 drain_right.t10 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X15 source.t20 minus.t11 drain_right.t3 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X16 drain_left.t13 plus.t2 source.t14 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X17 source.t6 plus.t3 drain_left.t12 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X18 a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X19 source.t5 plus.t4 drain_left.t11 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X20 source.t7 plus.t5 drain_left.t10 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X21 source.t12 plus.t6 drain_left.t9 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X22 drain_right.t11 minus.t12 source.t19 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X23 drain_right.t0 minus.t13 source.t18 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X24 drain_left.t8 plus.t7 source.t0 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X25 drain_left.t7 plus.t8 source.t13 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X26 drain_left.t6 plus.t9 source.t1 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X27 drain_left.t5 plus.t10 source.t8 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X28 a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X29 source.t11 plus.t11 drain_left.t4 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X30 drain_left.t3 plus.t12 source.t3 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X31 source.t9 plus.t13 drain_left.t2 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X32 source.t17 minus.t14 drain_right.t9 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X33 source.t16 minus.t15 drain_right.t12 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X34 drain_left.t1 plus.t14 source.t2 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X35 source.t10 plus.t15 drain_left.t0 a_n1670_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n17 minus.t15 1293
R1 minus.n4 minus.t12 1293
R2 minus.n36 minus.t6 1293
R3 minus.n23 minus.t1 1293
R4 minus.n16 minus.t3 1241.15
R5 minus.n14 minus.t10 1241.15
R6 minus.n1 minus.t13 1241.15
R7 minus.n9 minus.t14 1241.15
R8 minus.n7 minus.t2 1241.15
R9 minus.n3 minus.t11 1241.15
R10 minus.n35 minus.t8 1241.15
R11 minus.n33 minus.t7 1241.15
R12 minus.n20 minus.t9 1241.15
R13 minus.n28 minus.t4 1241.15
R14 minus.n26 minus.t0 1241.15
R15 minus.n22 minus.t5 1241.15
R16 minus.n5 minus.n4 161.489
R17 minus.n24 minus.n23 161.489
R18 minus.n18 minus.n17 161.3
R19 minus.n15 minus.n0 161.3
R20 minus.n13 minus.n12 161.3
R21 minus.n11 minus.n10 161.3
R22 minus.n8 minus.n2 161.3
R23 minus.n6 minus.n5 161.3
R24 minus.n37 minus.n36 161.3
R25 minus.n34 minus.n19 161.3
R26 minus.n32 minus.n31 161.3
R27 minus.n30 minus.n29 161.3
R28 minus.n27 minus.n21 161.3
R29 minus.n25 minus.n24 161.3
R30 minus.n16 minus.n15 47.4702
R31 minus.n6 minus.n3 47.4702
R32 minus.n25 minus.n22 47.4702
R33 minus.n35 minus.n34 47.4702
R34 minus.n14 minus.n13 43.0884
R35 minus.n8 minus.n7 43.0884
R36 minus.n27 minus.n26 43.0884
R37 minus.n33 minus.n32 43.0884
R38 minus.n10 minus.n1 38.7066
R39 minus.n10 minus.n9 38.7066
R40 minus.n29 minus.n28 38.7066
R41 minus.n29 minus.n20 38.7066
R42 minus.n13 minus.n1 34.3247
R43 minus.n9 minus.n8 34.3247
R44 minus.n28 minus.n27 34.3247
R45 minus.n32 minus.n20 34.3247
R46 minus.n38 minus.n18 33.1407
R47 minus.n15 minus.n14 29.9429
R48 minus.n7 minus.n6 29.9429
R49 minus.n26 minus.n25 29.9429
R50 minus.n34 minus.n33 29.9429
R51 minus.n17 minus.n16 25.5611
R52 minus.n4 minus.n3 25.5611
R53 minus.n23 minus.n22 25.5611
R54 minus.n36 minus.n35 25.5611
R55 minus.n38 minus.n37 6.46641
R56 minus.n18 minus.n0 0.189894
R57 minus.n12 minus.n0 0.189894
R58 minus.n12 minus.n11 0.189894
R59 minus.n11 minus.n2 0.189894
R60 minus.n5 minus.n2 0.189894
R61 minus.n24 minus.n21 0.189894
R62 minus.n30 minus.n21 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n19 0.189894
R65 minus.n37 minus.n19 0.189894
R66 minus minus.n38 0.188
R67 drain_right.n9 drain_right.n7 65.9943
R68 drain_right.n5 drain_right.n3 65.9942
R69 drain_right.n2 drain_right.n0 65.9942
R70 drain_right.n9 drain_right.n8 65.5376
R71 drain_right.n11 drain_right.n10 65.5376
R72 drain_right.n13 drain_right.n12 65.5376
R73 drain_right.n5 drain_right.n4 65.5373
R74 drain_right.n2 drain_right.n1 65.5373
R75 drain_right drain_right.n6 27.5109
R76 drain_right drain_right.n13 6.11011
R77 drain_right.n3 drain_right.t5 2.2005
R78 drain_right.n3 drain_right.t2 2.2005
R79 drain_right.n4 drain_right.t14 2.2005
R80 drain_right.n4 drain_right.t7 2.2005
R81 drain_right.n1 drain_right.t4 2.2005
R82 drain_right.n1 drain_right.t8 2.2005
R83 drain_right.n0 drain_right.t13 2.2005
R84 drain_right.n0 drain_right.t1 2.2005
R85 drain_right.n7 drain_right.t3 2.2005
R86 drain_right.n7 drain_right.t11 2.2005
R87 drain_right.n8 drain_right.t9 2.2005
R88 drain_right.n8 drain_right.t6 2.2005
R89 drain_right.n10 drain_right.t10 2.2005
R90 drain_right.n10 drain_right.t0 2.2005
R91 drain_right.n12 drain_right.t12 2.2005
R92 drain_right.n12 drain_right.t15 2.2005
R93 drain_right.n13 drain_right.n11 0.457397
R94 drain_right.n11 drain_right.n9 0.457397
R95 drain_right.n6 drain_right.n5 0.173602
R96 drain_right.n6 drain_right.n2 0.173602
R97 source.n7 source.t6 51.0588
R98 source.n8 source.t19 51.0588
R99 source.n15 source.t16 51.0588
R100 source.n31 source.t25 51.0586
R101 source.n24 source.t30 51.0586
R102 source.n23 source.t1 51.0586
R103 source.n16 source.t5 51.0586
R104 source.n0 source.t2 51.0586
R105 source.n2 source.n1 48.8588
R106 source.n4 source.n3 48.8588
R107 source.n6 source.n5 48.8588
R108 source.n10 source.n9 48.8588
R109 source.n12 source.n11 48.8588
R110 source.n14 source.n13 48.8588
R111 source.n30 source.n29 48.8586
R112 source.n28 source.n27 48.8586
R113 source.n26 source.n25 48.8586
R114 source.n22 source.n21 48.8586
R115 source.n20 source.n19 48.8586
R116 source.n18 source.n17 48.8586
R117 source.n16 source.n15 19.4719
R118 source.n32 source.n0 13.9805
R119 source.n32 source.n31 5.49188
R120 source.n29 source.t24 2.2005
R121 source.n29 source.t23 2.2005
R122 source.n27 source.t27 2.2005
R123 source.n27 source.t22 2.2005
R124 source.n25 source.t26 2.2005
R125 source.n25 source.t31 2.2005
R126 source.n21 source.t8 2.2005
R127 source.n21 source.t9 2.2005
R128 source.n19 source.t13 2.2005
R129 source.n19 source.t7 2.2005
R130 source.n17 source.t0 2.2005
R131 source.n17 source.t12 2.2005
R132 source.n1 source.t14 2.2005
R133 source.n1 source.t4 2.2005
R134 source.n3 source.t3 2.2005
R135 source.n3 source.t11 2.2005
R136 source.n5 source.t15 2.2005
R137 source.n5 source.t10 2.2005
R138 source.n9 source.t29 2.2005
R139 source.n9 source.t20 2.2005
R140 source.n11 source.t18 2.2005
R141 source.n11 source.t17 2.2005
R142 source.n13 source.t28 2.2005
R143 source.n13 source.t21 2.2005
R144 source.n8 source.n7 0.470328
R145 source.n24 source.n23 0.470328
R146 source.n15 source.n14 0.457397
R147 source.n14 source.n12 0.457397
R148 source.n12 source.n10 0.457397
R149 source.n10 source.n8 0.457397
R150 source.n7 source.n6 0.457397
R151 source.n6 source.n4 0.457397
R152 source.n4 source.n2 0.457397
R153 source.n2 source.n0 0.457397
R154 source.n18 source.n16 0.457397
R155 source.n20 source.n18 0.457397
R156 source.n22 source.n20 0.457397
R157 source.n23 source.n22 0.457397
R158 source.n26 source.n24 0.457397
R159 source.n28 source.n26 0.457397
R160 source.n30 source.n28 0.457397
R161 source.n31 source.n30 0.457397
R162 source source.n32 0.188
R163 plus.n4 plus.t3 1293
R164 plus.n17 plus.t14 1293
R165 plus.n23 plus.t9 1293
R166 plus.n36 plus.t4 1293
R167 plus.n3 plus.t1 1241.15
R168 plus.n7 plus.t15 1241.15
R169 plus.n9 plus.t12 1241.15
R170 plus.n1 plus.t11 1241.15
R171 plus.n14 plus.t2 1241.15
R172 plus.n16 plus.t0 1241.15
R173 plus.n22 plus.t13 1241.15
R174 plus.n26 plus.t10 1241.15
R175 plus.n28 plus.t5 1241.15
R176 plus.n20 plus.t8 1241.15
R177 plus.n33 plus.t6 1241.15
R178 plus.n35 plus.t7 1241.15
R179 plus.n5 plus.n4 161.489
R180 plus.n24 plus.n23 161.489
R181 plus.n6 plus.n5 161.3
R182 plus.n8 plus.n2 161.3
R183 plus.n11 plus.n10 161.3
R184 plus.n13 plus.n12 161.3
R185 plus.n15 plus.n0 161.3
R186 plus.n18 plus.n17 161.3
R187 plus.n25 plus.n24 161.3
R188 plus.n27 plus.n21 161.3
R189 plus.n30 plus.n29 161.3
R190 plus.n32 plus.n31 161.3
R191 plus.n34 plus.n19 161.3
R192 plus.n37 plus.n36 161.3
R193 plus.n6 plus.n3 47.4702
R194 plus.n16 plus.n15 47.4702
R195 plus.n35 plus.n34 47.4702
R196 plus.n25 plus.n22 47.4702
R197 plus.n8 plus.n7 43.0884
R198 plus.n14 plus.n13 43.0884
R199 plus.n33 plus.n32 43.0884
R200 plus.n27 plus.n26 43.0884
R201 plus.n10 plus.n9 38.7066
R202 plus.n10 plus.n1 38.7066
R203 plus.n29 plus.n20 38.7066
R204 plus.n29 plus.n28 38.7066
R205 plus.n9 plus.n8 34.3247
R206 plus.n13 plus.n1 34.3247
R207 plus.n32 plus.n20 34.3247
R208 plus.n28 plus.n27 34.3247
R209 plus.n7 plus.n6 29.9429
R210 plus.n15 plus.n14 29.9429
R211 plus.n34 plus.n33 29.9429
R212 plus.n26 plus.n25 29.9429
R213 plus plus.n37 28.1581
R214 plus.n4 plus.n3 25.5611
R215 plus.n17 plus.n16 25.5611
R216 plus.n36 plus.n35 25.5611
R217 plus.n23 plus.n22 25.5611
R218 plus plus.n18 10.974
R219 plus.n5 plus.n2 0.189894
R220 plus.n11 plus.n2 0.189894
R221 plus.n12 plus.n11 0.189894
R222 plus.n12 plus.n0 0.189894
R223 plus.n18 plus.n0 0.189894
R224 plus.n37 plus.n19 0.189894
R225 plus.n31 plus.n19 0.189894
R226 plus.n31 plus.n30 0.189894
R227 plus.n30 plus.n21 0.189894
R228 plus.n24 plus.n21 0.189894
R229 drain_left.n9 drain_left.n7 65.9945
R230 drain_left.n5 drain_left.n3 65.9942
R231 drain_left.n2 drain_left.n0 65.9942
R232 drain_left.n11 drain_left.n10 65.5376
R233 drain_left.n9 drain_left.n8 65.5376
R234 drain_left.n13 drain_left.n12 65.5374
R235 drain_left.n5 drain_left.n4 65.5373
R236 drain_left.n2 drain_left.n1 65.5373
R237 drain_left drain_left.n6 28.0642
R238 drain_left drain_left.n13 6.11011
R239 drain_left.n3 drain_left.t2 2.2005
R240 drain_left.n3 drain_left.t6 2.2005
R241 drain_left.n4 drain_left.t10 2.2005
R242 drain_left.n4 drain_left.t5 2.2005
R243 drain_left.n1 drain_left.t9 2.2005
R244 drain_left.n1 drain_left.t7 2.2005
R245 drain_left.n0 drain_left.t11 2.2005
R246 drain_left.n0 drain_left.t8 2.2005
R247 drain_left.n12 drain_left.t15 2.2005
R248 drain_left.n12 drain_left.t1 2.2005
R249 drain_left.n10 drain_left.t4 2.2005
R250 drain_left.n10 drain_left.t13 2.2005
R251 drain_left.n8 drain_left.t0 2.2005
R252 drain_left.n8 drain_left.t3 2.2005
R253 drain_left.n7 drain_left.t12 2.2005
R254 drain_left.n7 drain_left.t14 2.2005
R255 drain_left.n11 drain_left.n9 0.457397
R256 drain_left.n13 drain_left.n11 0.457397
R257 drain_left.n6 drain_left.n5 0.173602
R258 drain_left.n6 drain_left.n2 0.173602
C0 drain_left drain_right 0.846053f
C1 drain_left source 28.1968f
C2 plus drain_right 0.314737f
C3 plus source 3.1789f
C4 minus drain_right 3.44236f
C5 source minus 3.16486f
C6 drain_left plus 3.60333f
C7 drain_left minus 0.170856f
C8 plus minus 4.68167f
C9 source drain_right 28.1965f
C10 drain_right a_n1670_n2688# 6.04632f
C11 drain_left a_n1670_n2688# 6.32178f
C12 source a_n1670_n2688# 6.943649f
C13 minus a_n1670_n2688# 6.270106f
C14 plus a_n1670_n2688# 8.12869f
C15 drain_left.t11 a_n1670_n2688# 0.271992f
C16 drain_left.t8 a_n1670_n2688# 0.271992f
C17 drain_left.n0 a_n1670_n2688# 2.38203f
C18 drain_left.t9 a_n1670_n2688# 0.271992f
C19 drain_left.t7 a_n1670_n2688# 0.271992f
C20 drain_left.n1 a_n1670_n2688# 2.37902f
C21 drain_left.n2 a_n1670_n2688# 0.820432f
C22 drain_left.t2 a_n1670_n2688# 0.271992f
C23 drain_left.t6 a_n1670_n2688# 0.271992f
C24 drain_left.n3 a_n1670_n2688# 2.38203f
C25 drain_left.t10 a_n1670_n2688# 0.271992f
C26 drain_left.t5 a_n1670_n2688# 0.271992f
C27 drain_left.n4 a_n1670_n2688# 2.37902f
C28 drain_left.n5 a_n1670_n2688# 0.820432f
C29 drain_left.n6 a_n1670_n2688# 1.53517f
C30 drain_left.t12 a_n1670_n2688# 0.271992f
C31 drain_left.t14 a_n1670_n2688# 0.271992f
C32 drain_left.n7 a_n1670_n2688# 2.38203f
C33 drain_left.t0 a_n1670_n2688# 0.271992f
C34 drain_left.t3 a_n1670_n2688# 0.271992f
C35 drain_left.n8 a_n1670_n2688# 2.37902f
C36 drain_left.n9 a_n1670_n2688# 0.850272f
C37 drain_left.t4 a_n1670_n2688# 0.271992f
C38 drain_left.t13 a_n1670_n2688# 0.271992f
C39 drain_left.n10 a_n1670_n2688# 2.37902f
C40 drain_left.n11 a_n1670_n2688# 0.418938f
C41 drain_left.t15 a_n1670_n2688# 0.271992f
C42 drain_left.t1 a_n1670_n2688# 0.271992f
C43 drain_left.n12 a_n1670_n2688# 2.37901f
C44 drain_left.n13 a_n1670_n2688# 0.731936f
C45 plus.n0 a_n1670_n2688# 0.055217f
C46 plus.t0 a_n1670_n2688# 0.281635f
C47 plus.t2 a_n1670_n2688# 0.281635f
C48 plus.t11 a_n1670_n2688# 0.281635f
C49 plus.n1 a_n1670_n2688# 0.12328f
C50 plus.n2 a_n1670_n2688# 0.055217f
C51 plus.t12 a_n1670_n2688# 0.281635f
C52 plus.t15 a_n1670_n2688# 0.281635f
C53 plus.t1 a_n1670_n2688# 0.281635f
C54 plus.n3 a_n1670_n2688# 0.12328f
C55 plus.t3 a_n1670_n2688# 0.286653f
C56 plus.n4 a_n1670_n2688# 0.139553f
C57 plus.n5 a_n1670_n2688# 0.124311f
C58 plus.n6 a_n1670_n2688# 0.019339f
C59 plus.n7 a_n1670_n2688# 0.12328f
C60 plus.n8 a_n1670_n2688# 0.019339f
C61 plus.n9 a_n1670_n2688# 0.12328f
C62 plus.n10 a_n1670_n2688# 0.019339f
C63 plus.n11 a_n1670_n2688# 0.055217f
C64 plus.n12 a_n1670_n2688# 0.055217f
C65 plus.n13 a_n1670_n2688# 0.019339f
C66 plus.n14 a_n1670_n2688# 0.12328f
C67 plus.n15 a_n1670_n2688# 0.019339f
C68 plus.n16 a_n1670_n2688# 0.12328f
C69 plus.t14 a_n1670_n2688# 0.286653f
C70 plus.n17 a_n1670_n2688# 0.139472f
C71 plus.n18 a_n1670_n2688# 0.537893f
C72 plus.n19 a_n1670_n2688# 0.055217f
C73 plus.t4 a_n1670_n2688# 0.286653f
C74 plus.t7 a_n1670_n2688# 0.281635f
C75 plus.t6 a_n1670_n2688# 0.281635f
C76 plus.t8 a_n1670_n2688# 0.281635f
C77 plus.n20 a_n1670_n2688# 0.12328f
C78 plus.n21 a_n1670_n2688# 0.055217f
C79 plus.t5 a_n1670_n2688# 0.281635f
C80 plus.t10 a_n1670_n2688# 0.281635f
C81 plus.t13 a_n1670_n2688# 0.281635f
C82 plus.n22 a_n1670_n2688# 0.12328f
C83 plus.t9 a_n1670_n2688# 0.286653f
C84 plus.n23 a_n1670_n2688# 0.139553f
C85 plus.n24 a_n1670_n2688# 0.124311f
C86 plus.n25 a_n1670_n2688# 0.019339f
C87 plus.n26 a_n1670_n2688# 0.12328f
C88 plus.n27 a_n1670_n2688# 0.019339f
C89 plus.n28 a_n1670_n2688# 0.12328f
C90 plus.n29 a_n1670_n2688# 0.019339f
C91 plus.n30 a_n1670_n2688# 0.055217f
C92 plus.n31 a_n1670_n2688# 0.055217f
C93 plus.n32 a_n1670_n2688# 0.019339f
C94 plus.n33 a_n1670_n2688# 0.12328f
C95 plus.n34 a_n1670_n2688# 0.019339f
C96 plus.n35 a_n1670_n2688# 0.12328f
C97 plus.n36 a_n1670_n2688# 0.139472f
C98 plus.n37 a_n1670_n2688# 1.47584f
C99 source.t2 a_n1670_n2688# 2.46343f
C100 source.n0 a_n1670_n2688# 1.40143f
C101 source.t14 a_n1670_n2688# 0.231016f
C102 source.t4 a_n1670_n2688# 0.231016f
C103 source.n1 a_n1670_n2688# 1.93391f
C104 source.n2 a_n1670_n2688# 0.398382f
C105 source.t3 a_n1670_n2688# 0.231016f
C106 source.t11 a_n1670_n2688# 0.231016f
C107 source.n3 a_n1670_n2688# 1.93391f
C108 source.n4 a_n1670_n2688# 0.398382f
C109 source.t15 a_n1670_n2688# 0.231016f
C110 source.t10 a_n1670_n2688# 0.231016f
C111 source.n5 a_n1670_n2688# 1.93391f
C112 source.n6 a_n1670_n2688# 0.398382f
C113 source.t6 a_n1670_n2688# 2.46343f
C114 source.n7 a_n1670_n2688# 0.500257f
C115 source.t19 a_n1670_n2688# 2.46343f
C116 source.n8 a_n1670_n2688# 0.500257f
C117 source.t29 a_n1670_n2688# 0.231016f
C118 source.t20 a_n1670_n2688# 0.231016f
C119 source.n9 a_n1670_n2688# 1.93391f
C120 source.n10 a_n1670_n2688# 0.398382f
C121 source.t18 a_n1670_n2688# 0.231016f
C122 source.t17 a_n1670_n2688# 0.231016f
C123 source.n11 a_n1670_n2688# 1.93391f
C124 source.n12 a_n1670_n2688# 0.398382f
C125 source.t28 a_n1670_n2688# 0.231016f
C126 source.t21 a_n1670_n2688# 0.231016f
C127 source.n13 a_n1670_n2688# 1.93391f
C128 source.n14 a_n1670_n2688# 0.398382f
C129 source.t16 a_n1670_n2688# 2.46343f
C130 source.n15 a_n1670_n2688# 1.87045f
C131 source.t5 a_n1670_n2688# 2.46343f
C132 source.n16 a_n1670_n2688# 1.87046f
C133 source.t0 a_n1670_n2688# 0.231016f
C134 source.t12 a_n1670_n2688# 0.231016f
C135 source.n17 a_n1670_n2688# 1.93391f
C136 source.n18 a_n1670_n2688# 0.398387f
C137 source.t13 a_n1670_n2688# 0.231016f
C138 source.t7 a_n1670_n2688# 0.231016f
C139 source.n19 a_n1670_n2688# 1.93391f
C140 source.n20 a_n1670_n2688# 0.398387f
C141 source.t8 a_n1670_n2688# 0.231016f
C142 source.t9 a_n1670_n2688# 0.231016f
C143 source.n21 a_n1670_n2688# 1.93391f
C144 source.n22 a_n1670_n2688# 0.398387f
C145 source.t1 a_n1670_n2688# 2.46343f
C146 source.n23 a_n1670_n2688# 0.500263f
C147 source.t30 a_n1670_n2688# 2.46343f
C148 source.n24 a_n1670_n2688# 0.500263f
C149 source.t26 a_n1670_n2688# 0.231016f
C150 source.t31 a_n1670_n2688# 0.231016f
C151 source.n25 a_n1670_n2688# 1.93391f
C152 source.n26 a_n1670_n2688# 0.398387f
C153 source.t27 a_n1670_n2688# 0.231016f
C154 source.t22 a_n1670_n2688# 0.231016f
C155 source.n27 a_n1670_n2688# 1.93391f
C156 source.n28 a_n1670_n2688# 0.398387f
C157 source.t24 a_n1670_n2688# 0.231016f
C158 source.t23 a_n1670_n2688# 0.231016f
C159 source.n29 a_n1670_n2688# 1.93391f
C160 source.n30 a_n1670_n2688# 0.398387f
C161 source.t25 a_n1670_n2688# 2.46343f
C162 source.n31 a_n1670_n2688# 0.676392f
C163 source.n32 a_n1670_n2688# 1.6862f
C164 drain_right.t13 a_n1670_n2688# 0.271559f
C165 drain_right.t1 a_n1670_n2688# 0.271559f
C166 drain_right.n0 a_n1670_n2688# 2.37823f
C167 drain_right.t4 a_n1670_n2688# 0.271559f
C168 drain_right.t8 a_n1670_n2688# 0.271559f
C169 drain_right.n1 a_n1670_n2688# 2.37523f
C170 drain_right.n2 a_n1670_n2688# 0.819125f
C171 drain_right.t5 a_n1670_n2688# 0.271559f
C172 drain_right.t2 a_n1670_n2688# 0.271559f
C173 drain_right.n3 a_n1670_n2688# 2.37823f
C174 drain_right.t14 a_n1670_n2688# 0.271559f
C175 drain_right.t7 a_n1670_n2688# 0.271559f
C176 drain_right.n4 a_n1670_n2688# 2.37523f
C177 drain_right.n5 a_n1670_n2688# 0.819125f
C178 drain_right.n6 a_n1670_n2688# 1.45389f
C179 drain_right.t3 a_n1670_n2688# 0.271559f
C180 drain_right.t11 a_n1670_n2688# 0.271559f
C181 drain_right.n7 a_n1670_n2688# 2.37823f
C182 drain_right.t9 a_n1670_n2688# 0.271559f
C183 drain_right.t6 a_n1670_n2688# 0.271559f
C184 drain_right.n8 a_n1670_n2688# 2.37524f
C185 drain_right.n9 a_n1670_n2688# 0.848928f
C186 drain_right.t10 a_n1670_n2688# 0.271559f
C187 drain_right.t0 a_n1670_n2688# 0.271559f
C188 drain_right.n10 a_n1670_n2688# 2.37524f
C189 drain_right.n11 a_n1670_n2688# 0.418271f
C190 drain_right.t12 a_n1670_n2688# 0.271559f
C191 drain_right.t15 a_n1670_n2688# 0.271559f
C192 drain_right.n12 a_n1670_n2688# 2.37524f
C193 drain_right.n13 a_n1670_n2688# 0.730761f
C194 minus.n0 a_n1670_n2688# 0.053735f
C195 minus.t15 a_n1670_n2688# 0.27896f
C196 minus.t3 a_n1670_n2688# 0.274075f
C197 minus.t10 a_n1670_n2688# 0.274075f
C198 minus.t13 a_n1670_n2688# 0.274075f
C199 minus.n1 a_n1670_n2688# 0.119971f
C200 minus.n2 a_n1670_n2688# 0.053735f
C201 minus.t14 a_n1670_n2688# 0.274075f
C202 minus.t2 a_n1670_n2688# 0.274075f
C203 minus.t11 a_n1670_n2688# 0.274075f
C204 minus.n3 a_n1670_n2688# 0.119971f
C205 minus.t12 a_n1670_n2688# 0.27896f
C206 minus.n4 a_n1670_n2688# 0.135807f
C207 minus.n5 a_n1670_n2688# 0.120975f
C208 minus.n6 a_n1670_n2688# 0.01882f
C209 minus.n7 a_n1670_n2688# 0.119971f
C210 minus.n8 a_n1670_n2688# 0.01882f
C211 minus.n9 a_n1670_n2688# 0.119971f
C212 minus.n10 a_n1670_n2688# 0.01882f
C213 minus.n11 a_n1670_n2688# 0.053735f
C214 minus.n12 a_n1670_n2688# 0.053735f
C215 minus.n13 a_n1670_n2688# 0.01882f
C216 minus.n14 a_n1670_n2688# 0.119971f
C217 minus.n15 a_n1670_n2688# 0.01882f
C218 minus.n16 a_n1670_n2688# 0.119971f
C219 minus.n17 a_n1670_n2688# 0.135728f
C220 minus.n18 a_n1670_n2688# 1.64859f
C221 minus.n19 a_n1670_n2688# 0.053735f
C222 minus.t8 a_n1670_n2688# 0.274075f
C223 minus.t7 a_n1670_n2688# 0.274075f
C224 minus.t9 a_n1670_n2688# 0.274075f
C225 minus.n20 a_n1670_n2688# 0.119971f
C226 minus.n21 a_n1670_n2688# 0.053735f
C227 minus.t4 a_n1670_n2688# 0.274075f
C228 minus.t0 a_n1670_n2688# 0.274075f
C229 minus.t5 a_n1670_n2688# 0.274075f
C230 minus.n22 a_n1670_n2688# 0.119971f
C231 minus.t1 a_n1670_n2688# 0.27896f
C232 minus.n23 a_n1670_n2688# 0.135807f
C233 minus.n24 a_n1670_n2688# 0.120975f
C234 minus.n25 a_n1670_n2688# 0.01882f
C235 minus.n26 a_n1670_n2688# 0.119971f
C236 minus.n27 a_n1670_n2688# 0.01882f
C237 minus.n28 a_n1670_n2688# 0.119971f
C238 minus.n29 a_n1670_n2688# 0.01882f
C239 minus.n30 a_n1670_n2688# 0.053735f
C240 minus.n31 a_n1670_n2688# 0.053735f
C241 minus.n32 a_n1670_n2688# 0.01882f
C242 minus.n33 a_n1670_n2688# 0.119971f
C243 minus.n34 a_n1670_n2688# 0.01882f
C244 minus.n35 a_n1670_n2688# 0.119971f
C245 minus.t6 a_n1670_n2688# 0.27896f
C246 minus.n36 a_n1670_n2688# 0.135728f
C247 minus.n37 a_n1670_n2688# 0.347047f
C248 minus.n38 a_n1670_n2688# 2.02158f
.ends

