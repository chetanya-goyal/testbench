* NGSPICE file created from diffpair461.ext - technology: sky130A

.subckt diffpair461 minus drain_right drain_left source plus
X0 a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X1 source minus drain_right a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X2 source minus drain_right a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X3 drain_right minus source a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X4 a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X5 source plus drain_left a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X6 a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X7 drain_right minus source a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X8 drain_left plus source a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X9 drain_left plus source a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X10 a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X11 source plus drain_left a_n1334_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
.ends

