* NGSPICE file created from diffpair591.ext - technology: sky130A

.subckt diffpair591 minus drain_right drain_left source plus
X0 drain_right minus source a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 source plus drain_left a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X2 drain_right minus source a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X3 source minus drain_right a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X4 a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X5 drain_left plus source a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X6 a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X7 source minus drain_right a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X8 a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X9 source plus drain_left a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X10 a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X11 drain_left plus source a_n1094_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
.ends

