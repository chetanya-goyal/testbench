* NGSPICE file created from diffpair198.ext - technology: sky130A

.subckt diffpair198 minus drain_right drain_left source plus
X0 source.t37 minus.t0 drain_right.t2 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 drain_right.t3 minus.t1 source.t36 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X2 drain_left.t19 plus.t0 source.t1 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X3 drain_left.t18 plus.t1 source.t4 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X4 source.t35 minus.t2 drain_right.t9 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X5 drain_right.t6 minus.t3 source.t34 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X6 drain_left.t17 plus.t2 source.t8 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X7 drain_right.t0 minus.t4 source.t33 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X8 drain_right.t7 minus.t5 source.t32 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X9 source.t31 minus.t6 drain_right.t4 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X10 source.t10 plus.t3 drain_left.t16 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X11 source.t14 plus.t4 drain_left.t15 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X12 drain_left.t14 plus.t5 source.t15 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X13 drain_right.t8 minus.t7 source.t30 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X14 source.t29 minus.t8 drain_right.t10 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X15 a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X16 source.t28 minus.t9 drain_right.t5 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X17 source.t38 plus.t6 drain_left.t13 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X18 source.t39 plus.t7 drain_left.t12 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X19 drain_left.t11 plus.t8 source.t3 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X20 drain_right.t1 minus.t10 source.t27 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X21 source.t26 minus.t11 drain_right.t12 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X22 drain_left.t10 plus.t9 source.t0 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X23 a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X24 source.t2 plus.t10 drain_left.t9 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X25 drain_right.t11 minus.t12 source.t25 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X26 drain_right.t13 minus.t13 source.t24 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X27 drain_left.t8 plus.t11 source.t13 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X28 source.t11 plus.t12 drain_left.t7 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X29 source.t23 minus.t14 drain_right.t14 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X30 source.t7 plus.t13 drain_left.t6 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X31 a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X32 drain_left.t5 plus.t14 source.t9 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X33 drain_left.t4 plus.t15 source.t12 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X34 drain_right.t15 minus.t15 source.t22 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X35 source.t21 minus.t16 drain_right.t16 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X36 source.t20 minus.t17 drain_right.t17 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X37 drain_right.t18 minus.t18 source.t19 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X38 a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X39 source.t18 minus.t19 drain_right.t19 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X40 source.t5 plus.t16 drain_left.t3 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X41 source.t6 plus.t17 drain_left.t2 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X42 source.t17 plus.t18 drain_left.t1 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X43 drain_left.t0 plus.t19 source.t16 a_n2102_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n27 minus.t8 394.365
R1 minus.n7 minus.t12 394.365
R2 minus.n56 minus.t18 394.365
R3 minus.n35 minus.t9 394.365
R4 minus.n26 minus.t5 345.433
R5 minus.n24 minus.t17 345.433
R6 minus.n3 minus.t7 345.433
R7 minus.n18 minus.t2 345.433
R8 minus.n16 minus.t15 345.433
R9 minus.n4 minus.t11 345.433
R10 minus.n10 minus.t4 345.433
R11 minus.n6 minus.t16 345.433
R12 minus.n55 minus.t0 345.433
R13 minus.n53 minus.t13 345.433
R14 minus.n47 minus.t14 345.433
R15 minus.n46 minus.t3 345.433
R16 minus.n44 minus.t6 345.433
R17 minus.n32 minus.t10 345.433
R18 minus.n38 minus.t19 345.433
R19 minus.n34 minus.t1 345.433
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 64.9975
R47 minus.n15 minus.n4 64.9975
R48 minus.n43 minus.n32 64.9975
R49 minus.n48 minus.n47 64.9975
R50 minus.n25 minus.n24 62.0763
R51 minus.n10 minus.n9 62.0763
R52 minus.n38 minus.n37 62.0763
R53 minus.n54 minus.n53 62.0763
R54 minus.n18 minus.n17 46.0096
R55 minus.n17 minus.n16 46.0096
R56 minus.n45 minus.n44 46.0096
R57 minus.n46 minus.n45 46.0096
R58 minus.n27 minus.n26 43.0884
R59 minus.n7 minus.n6 43.0884
R60 minus.n35 minus.n34 43.0884
R61 minus.n56 minus.n55 43.0884
R62 minus.n58 minus.n28 30.2808
R63 minus.n26 minus.n25 29.9429
R64 minus.n9 minus.n6 29.9429
R65 minus.n37 minus.n34 29.9429
R66 minus.n55 minus.n54 29.9429
R67 minus.n19 minus.n18 27.0217
R68 minus.n16 minus.n15 27.0217
R69 minus.n44 minus.n43 27.0217
R70 minus.n48 minus.n46 27.0217
R71 minus.n24 minus.n23 10.955
R72 minus.n11 minus.n10 10.955
R73 minus.n39 minus.n38 10.955
R74 minus.n53 minus.n52 10.955
R75 minus.n3 minus.n1 8.03383
R76 minus.n12 minus.n4 8.03383
R77 minus.n40 minus.n32 8.03383
R78 minus.n47 minus.n30 8.03383
R79 minus.n58 minus.n57 6.51565
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 drain_right.n10 drain_right.n8 80.3162
R100 drain_right.n6 drain_right.n4 80.3161
R101 drain_right.n2 drain_right.n0 80.3161
R102 drain_right.n10 drain_right.n9 79.7731
R103 drain_right.n12 drain_right.n11 79.7731
R104 drain_right.n14 drain_right.n13 79.7731
R105 drain_right.n16 drain_right.n15 79.7731
R106 drain_right.n7 drain_right.n3 79.773
R107 drain_right.n6 drain_right.n5 79.773
R108 drain_right.n2 drain_right.n1 79.773
R109 drain_right drain_right.n7 24.3405
R110 drain_right.n3 drain_right.t4 6.6005
R111 drain_right.n3 drain_right.t6 6.6005
R112 drain_right.n4 drain_right.t2 6.6005
R113 drain_right.n4 drain_right.t18 6.6005
R114 drain_right.n5 drain_right.t14 6.6005
R115 drain_right.n5 drain_right.t13 6.6005
R116 drain_right.n1 drain_right.t19 6.6005
R117 drain_right.n1 drain_right.t1 6.6005
R118 drain_right.n0 drain_right.t5 6.6005
R119 drain_right.n0 drain_right.t3 6.6005
R120 drain_right.n8 drain_right.t16 6.6005
R121 drain_right.n8 drain_right.t11 6.6005
R122 drain_right.n9 drain_right.t12 6.6005
R123 drain_right.n9 drain_right.t0 6.6005
R124 drain_right.n11 drain_right.t9 6.6005
R125 drain_right.n11 drain_right.t15 6.6005
R126 drain_right.n13 drain_right.t17 6.6005
R127 drain_right.n13 drain_right.t8 6.6005
R128 drain_right.n15 drain_right.t10 6.6005
R129 drain_right.n15 drain_right.t7 6.6005
R130 drain_right drain_right.n16 6.19632
R131 drain_right.n16 drain_right.n14 0.543603
R132 drain_right.n14 drain_right.n12 0.543603
R133 drain_right.n12 drain_right.n10 0.543603
R134 drain_right.n7 drain_right.n6 0.488257
R135 drain_right.n7 drain_right.n2 0.488257
R136 source.n0 source.t12 69.6943
R137 source.n9 source.t14 69.6943
R138 source.n10 source.t25 69.6943
R139 source.n19 source.t29 69.6943
R140 source.n39 source.t19 69.6942
R141 source.n30 source.t28 69.6942
R142 source.n29 source.t15 69.6942
R143 source.n20 source.t11 69.6942
R144 source.n2 source.n1 63.0943
R145 source.n4 source.n3 63.0943
R146 source.n6 source.n5 63.0943
R147 source.n8 source.n7 63.0943
R148 source.n12 source.n11 63.0943
R149 source.n14 source.n13 63.0943
R150 source.n16 source.n15 63.0943
R151 source.n18 source.n17 63.0943
R152 source.n38 source.n37 63.0942
R153 source.n36 source.n35 63.0942
R154 source.n34 source.n33 63.0942
R155 source.n32 source.n31 63.0942
R156 source.n28 source.n27 63.0942
R157 source.n26 source.n25 63.0942
R158 source.n24 source.n23 63.0942
R159 source.n22 source.n21 63.0942
R160 source.n20 source.n19 15.0126
R161 source.n40 source.n0 9.47816
R162 source.n37 source.t24 6.6005
R163 source.n37 source.t37 6.6005
R164 source.n35 source.t34 6.6005
R165 source.n35 source.t23 6.6005
R166 source.n33 source.t27 6.6005
R167 source.n33 source.t31 6.6005
R168 source.n31 source.t36 6.6005
R169 source.n31 source.t18 6.6005
R170 source.n27 source.t9 6.6005
R171 source.n27 source.t5 6.6005
R172 source.n25 source.t8 6.6005
R173 source.n25 source.t39 6.6005
R174 source.n23 source.t0 6.6005
R175 source.n23 source.t17 6.6005
R176 source.n21 source.t1 6.6005
R177 source.n21 source.t10 6.6005
R178 source.n1 source.t4 6.6005
R179 source.n1 source.t2 6.6005
R180 source.n3 source.t13 6.6005
R181 source.n3 source.t6 6.6005
R182 source.n5 source.t16 6.6005
R183 source.n5 source.t38 6.6005
R184 source.n7 source.t3 6.6005
R185 source.n7 source.t7 6.6005
R186 source.n11 source.t33 6.6005
R187 source.n11 source.t21 6.6005
R188 source.n13 source.t22 6.6005
R189 source.n13 source.t26 6.6005
R190 source.n15 source.t30 6.6005
R191 source.n15 source.t35 6.6005
R192 source.n17 source.t32 6.6005
R193 source.n17 source.t20 6.6005
R194 source.n40 source.n39 5.53498
R195 source.n19 source.n18 0.543603
R196 source.n18 source.n16 0.543603
R197 source.n16 source.n14 0.543603
R198 source.n14 source.n12 0.543603
R199 source.n12 source.n10 0.543603
R200 source.n9 source.n8 0.543603
R201 source.n8 source.n6 0.543603
R202 source.n6 source.n4 0.543603
R203 source.n4 source.n2 0.543603
R204 source.n2 source.n0 0.543603
R205 source.n22 source.n20 0.543603
R206 source.n24 source.n22 0.543603
R207 source.n26 source.n24 0.543603
R208 source.n28 source.n26 0.543603
R209 source.n29 source.n28 0.543603
R210 source.n32 source.n30 0.543603
R211 source.n34 source.n32 0.543603
R212 source.n36 source.n34 0.543603
R213 source.n38 source.n36 0.543603
R214 source.n39 source.n38 0.543603
R215 source.n10 source.n9 0.470328
R216 source.n30 source.n29 0.470328
R217 source source.n40 0.188
R218 plus.n6 plus.t4 394.365
R219 plus.n27 plus.t15 394.365
R220 plus.n36 plus.t5 394.365
R221 plus.n56 plus.t12 394.365
R222 plus.n5 plus.t8 345.433
R223 plus.n9 plus.t13 345.433
R224 plus.n3 plus.t19 345.433
R225 plus.n15 plus.t6 345.433
R226 plus.n17 plus.t11 345.433
R227 plus.n18 plus.t17 345.433
R228 plus.n24 plus.t1 345.433
R229 plus.n26 plus.t10 345.433
R230 plus.n35 plus.t16 345.433
R231 plus.n39 plus.t14 345.433
R232 plus.n33 plus.t7 345.433
R233 plus.n45 plus.t2 345.433
R234 plus.n47 plus.t18 345.433
R235 plus.n32 plus.t9 345.433
R236 plus.n53 plus.t3 345.433
R237 plus.n55 plus.t0 345.433
R238 plus.n7 plus.n6 161.489
R239 plus.n37 plus.n36 161.489
R240 plus.n8 plus.n7 161.3
R241 plus.n10 plus.n4 161.3
R242 plus.n12 plus.n11 161.3
R243 plus.n14 plus.n13 161.3
R244 plus.n16 plus.n2 161.3
R245 plus.n20 plus.n19 161.3
R246 plus.n21 plus.n1 161.3
R247 plus.n23 plus.n22 161.3
R248 plus.n25 plus.n0 161.3
R249 plus.n28 plus.n27 161.3
R250 plus.n38 plus.n37 161.3
R251 plus.n40 plus.n34 161.3
R252 plus.n42 plus.n41 161.3
R253 plus.n44 plus.n43 161.3
R254 plus.n46 plus.n31 161.3
R255 plus.n49 plus.n48 161.3
R256 plus.n50 plus.n30 161.3
R257 plus.n52 plus.n51 161.3
R258 plus.n54 plus.n29 161.3
R259 plus.n57 plus.n56 161.3
R260 plus.n11 plus.n10 73.0308
R261 plus.n23 plus.n1 73.0308
R262 plus.n52 plus.n30 73.0308
R263 plus.n41 plus.n40 73.0308
R264 plus.n14 plus.n3 64.9975
R265 plus.n19 plus.n18 64.9975
R266 plus.n48 plus.n32 64.9975
R267 plus.n44 plus.n33 64.9975
R268 plus.n9 plus.n8 62.0763
R269 plus.n25 plus.n24 62.0763
R270 plus.n54 plus.n53 62.0763
R271 plus.n39 plus.n38 62.0763
R272 plus.n16 plus.n15 46.0096
R273 plus.n17 plus.n16 46.0096
R274 plus.n47 plus.n46 46.0096
R275 plus.n46 plus.n45 46.0096
R276 plus.n6 plus.n5 43.0884
R277 plus.n27 plus.n26 43.0884
R278 plus.n56 plus.n55 43.0884
R279 plus.n36 plus.n35 43.0884
R280 plus.n8 plus.n5 29.9429
R281 plus.n26 plus.n25 29.9429
R282 plus.n55 plus.n54 29.9429
R283 plus.n38 plus.n35 29.9429
R284 plus plus.n57 27.571
R285 plus.n15 plus.n14 27.0217
R286 plus.n19 plus.n17 27.0217
R287 plus.n48 plus.n47 27.0217
R288 plus.n45 plus.n44 27.0217
R289 plus.n10 plus.n9 10.955
R290 plus.n24 plus.n23 10.955
R291 plus.n53 plus.n52 10.955
R292 plus.n40 plus.n39 10.955
R293 plus plus.n28 8.7505
R294 plus.n11 plus.n3 8.03383
R295 plus.n18 plus.n1 8.03383
R296 plus.n32 plus.n30 8.03383
R297 plus.n41 plus.n33 8.03383
R298 plus.n7 plus.n4 0.189894
R299 plus.n12 plus.n4 0.189894
R300 plus.n13 plus.n12 0.189894
R301 plus.n13 plus.n2 0.189894
R302 plus.n20 plus.n2 0.189894
R303 plus.n21 plus.n20 0.189894
R304 plus.n22 plus.n21 0.189894
R305 plus.n22 plus.n0 0.189894
R306 plus.n28 plus.n0 0.189894
R307 plus.n57 plus.n29 0.189894
R308 plus.n51 plus.n29 0.189894
R309 plus.n51 plus.n50 0.189894
R310 plus.n50 plus.n49 0.189894
R311 plus.n49 plus.n31 0.189894
R312 plus.n43 plus.n31 0.189894
R313 plus.n43 plus.n42 0.189894
R314 plus.n42 plus.n34 0.189894
R315 plus.n37 plus.n34 0.189894
R316 drain_left.n10 drain_left.n8 80.3162
R317 drain_left.n6 drain_left.n4 80.3161
R318 drain_left.n2 drain_left.n0 80.3161
R319 drain_left.n16 drain_left.n15 79.7731
R320 drain_left.n14 drain_left.n13 79.7731
R321 drain_left.n12 drain_left.n11 79.7731
R322 drain_left.n10 drain_left.n9 79.7731
R323 drain_left.n7 drain_left.n3 79.773
R324 drain_left.n6 drain_left.n5 79.773
R325 drain_left.n2 drain_left.n1 79.773
R326 drain_left drain_left.n7 24.8937
R327 drain_left.n3 drain_left.t1 6.6005
R328 drain_left.n3 drain_left.t17 6.6005
R329 drain_left.n4 drain_left.t3 6.6005
R330 drain_left.n4 drain_left.t14 6.6005
R331 drain_left.n5 drain_left.t12 6.6005
R332 drain_left.n5 drain_left.t5 6.6005
R333 drain_left.n1 drain_left.t16 6.6005
R334 drain_left.n1 drain_left.t10 6.6005
R335 drain_left.n0 drain_left.t7 6.6005
R336 drain_left.n0 drain_left.t19 6.6005
R337 drain_left.n15 drain_left.t9 6.6005
R338 drain_left.n15 drain_left.t4 6.6005
R339 drain_left.n13 drain_left.t2 6.6005
R340 drain_left.n13 drain_left.t18 6.6005
R341 drain_left.n11 drain_left.t13 6.6005
R342 drain_left.n11 drain_left.t8 6.6005
R343 drain_left.n9 drain_left.t6 6.6005
R344 drain_left.n9 drain_left.t0 6.6005
R345 drain_left.n8 drain_left.t15 6.6005
R346 drain_left.n8 drain_left.t11 6.6005
R347 drain_left drain_left.n16 6.19632
R348 drain_left.n12 drain_left.n10 0.543603
R349 drain_left.n14 drain_left.n12 0.543603
R350 drain_left.n16 drain_left.n14 0.543603
R351 drain_left.n7 drain_left.n6 0.488257
R352 drain_left.n7 drain_left.n2 0.488257
C0 drain_left minus 0.176821f
C1 plus minus 4.11459f
C2 drain_left source 11.8472f
C3 plus source 2.4731f
C4 minus source 2.4591f
C5 drain_left drain_right 1.10834f
C6 drain_right plus 0.366353f
C7 drain_right minus 2.2481f
C8 drain_right source 11.8477f
C9 drain_left plus 2.45404f
C10 drain_right a_n2102_n1488# 4.84687f
C11 drain_left a_n2102_n1488# 5.18622f
C12 source a_n2102_n1488# 3.797055f
C13 minus a_n2102_n1488# 7.526808f
C14 plus a_n2102_n1488# 8.96716f
C15 drain_left.t7 a_n2102_n1488# 0.077565f
C16 drain_left.t19 a_n2102_n1488# 0.077565f
C17 drain_left.n0 a_n2102_n1488# 0.562021f
C18 drain_left.t16 a_n2102_n1488# 0.077565f
C19 drain_left.t10 a_n2102_n1488# 0.077565f
C20 drain_left.n1 a_n2102_n1488# 0.559387f
C21 drain_left.n2 a_n2102_n1488# 0.759097f
C22 drain_left.t1 a_n2102_n1488# 0.077565f
C23 drain_left.t17 a_n2102_n1488# 0.077565f
C24 drain_left.n3 a_n2102_n1488# 0.559387f
C25 drain_left.t3 a_n2102_n1488# 0.077565f
C26 drain_left.t14 a_n2102_n1488# 0.077565f
C27 drain_left.n4 a_n2102_n1488# 0.562021f
C28 drain_left.t12 a_n2102_n1488# 0.077565f
C29 drain_left.t5 a_n2102_n1488# 0.077565f
C30 drain_left.n5 a_n2102_n1488# 0.559387f
C31 drain_left.n6 a_n2102_n1488# 0.759097f
C32 drain_left.n7 a_n2102_n1488# 1.39652f
C33 drain_left.t15 a_n2102_n1488# 0.077565f
C34 drain_left.t11 a_n2102_n1488# 0.077565f
C35 drain_left.n8 a_n2102_n1488# 0.562024f
C36 drain_left.t6 a_n2102_n1488# 0.077565f
C37 drain_left.t0 a_n2102_n1488# 0.077565f
C38 drain_left.n9 a_n2102_n1488# 0.55939f
C39 drain_left.n10 a_n2102_n1488# 0.763371f
C40 drain_left.t13 a_n2102_n1488# 0.077565f
C41 drain_left.t8 a_n2102_n1488# 0.077565f
C42 drain_left.n11 a_n2102_n1488# 0.55939f
C43 drain_left.n12 a_n2102_n1488# 0.376414f
C44 drain_left.t2 a_n2102_n1488# 0.077565f
C45 drain_left.t18 a_n2102_n1488# 0.077565f
C46 drain_left.n13 a_n2102_n1488# 0.55939f
C47 drain_left.n14 a_n2102_n1488# 0.376414f
C48 drain_left.t9 a_n2102_n1488# 0.077565f
C49 drain_left.t4 a_n2102_n1488# 0.077565f
C50 drain_left.n15 a_n2102_n1488# 0.55939f
C51 drain_left.n16 a_n2102_n1488# 0.648746f
C52 plus.n0 a_n2102_n1488# 0.051619f
C53 plus.t10 a_n2102_n1488# 0.134535f
C54 plus.t1 a_n2102_n1488# 0.134535f
C55 plus.n1 a_n2102_n1488# 0.018874f
C56 plus.n2 a_n2102_n1488# 0.051619f
C57 plus.t11 a_n2102_n1488# 0.134535f
C58 plus.t6 a_n2102_n1488# 0.134535f
C59 plus.t19 a_n2102_n1488# 0.134535f
C60 plus.n3 a_n2102_n1488# 0.078117f
C61 plus.n4 a_n2102_n1488# 0.051619f
C62 plus.t13 a_n2102_n1488# 0.134535f
C63 plus.t8 a_n2102_n1488# 0.134535f
C64 plus.n5 a_n2102_n1488# 0.078117f
C65 plus.t4 a_n2102_n1488# 0.144761f
C66 plus.n6 a_n2102_n1488# 0.093527f
C67 plus.n7 a_n2102_n1488# 0.118119f
C68 plus.n8 a_n2102_n1488# 0.021261f
C69 plus.n9 a_n2102_n1488# 0.078117f
C70 plus.n10 a_n2102_n1488# 0.019511f
C71 plus.n11 a_n2102_n1488# 0.018874f
C72 plus.n12 a_n2102_n1488# 0.051619f
C73 plus.n13 a_n2102_n1488# 0.051619f
C74 plus.n14 a_n2102_n1488# 0.021261f
C75 plus.n15 a_n2102_n1488# 0.078117f
C76 plus.n16 a_n2102_n1488# 0.021261f
C77 plus.n17 a_n2102_n1488# 0.078117f
C78 plus.t17 a_n2102_n1488# 0.134535f
C79 plus.n18 a_n2102_n1488# 0.078117f
C80 plus.n19 a_n2102_n1488# 0.021261f
C81 plus.n20 a_n2102_n1488# 0.051619f
C82 plus.n21 a_n2102_n1488# 0.051619f
C83 plus.n22 a_n2102_n1488# 0.051619f
C84 plus.n23 a_n2102_n1488# 0.019511f
C85 plus.n24 a_n2102_n1488# 0.078117f
C86 plus.n25 a_n2102_n1488# 0.021261f
C87 plus.n26 a_n2102_n1488# 0.078117f
C88 plus.t15 a_n2102_n1488# 0.144761f
C89 plus.n27 a_n2102_n1488# 0.093449f
C90 plus.n28 a_n2102_n1488# 0.387592f
C91 plus.n29 a_n2102_n1488# 0.051619f
C92 plus.t12 a_n2102_n1488# 0.144761f
C93 plus.t0 a_n2102_n1488# 0.134535f
C94 plus.t3 a_n2102_n1488# 0.134535f
C95 plus.n30 a_n2102_n1488# 0.018874f
C96 plus.n31 a_n2102_n1488# 0.051619f
C97 plus.t9 a_n2102_n1488# 0.134535f
C98 plus.n32 a_n2102_n1488# 0.078117f
C99 plus.t18 a_n2102_n1488# 0.134535f
C100 plus.t2 a_n2102_n1488# 0.134535f
C101 plus.t7 a_n2102_n1488# 0.134535f
C102 plus.n33 a_n2102_n1488# 0.078117f
C103 plus.n34 a_n2102_n1488# 0.051619f
C104 plus.t14 a_n2102_n1488# 0.134535f
C105 plus.t16 a_n2102_n1488# 0.134535f
C106 plus.n35 a_n2102_n1488# 0.078117f
C107 plus.t5 a_n2102_n1488# 0.144761f
C108 plus.n36 a_n2102_n1488# 0.093527f
C109 plus.n37 a_n2102_n1488# 0.118119f
C110 plus.n38 a_n2102_n1488# 0.021261f
C111 plus.n39 a_n2102_n1488# 0.078117f
C112 plus.n40 a_n2102_n1488# 0.019511f
C113 plus.n41 a_n2102_n1488# 0.018874f
C114 plus.n42 a_n2102_n1488# 0.051619f
C115 plus.n43 a_n2102_n1488# 0.051619f
C116 plus.n44 a_n2102_n1488# 0.021261f
C117 plus.n45 a_n2102_n1488# 0.078117f
C118 plus.n46 a_n2102_n1488# 0.021261f
C119 plus.n47 a_n2102_n1488# 0.078117f
C120 plus.n48 a_n2102_n1488# 0.021261f
C121 plus.n49 a_n2102_n1488# 0.051619f
C122 plus.n50 a_n2102_n1488# 0.051619f
C123 plus.n51 a_n2102_n1488# 0.051619f
C124 plus.n52 a_n2102_n1488# 0.019511f
C125 plus.n53 a_n2102_n1488# 0.078117f
C126 plus.n54 a_n2102_n1488# 0.021261f
C127 plus.n55 a_n2102_n1488# 0.078117f
C128 plus.n56 a_n2102_n1488# 0.093449f
C129 plus.n57 a_n2102_n1488# 1.28245f
C130 source.t12 a_n2102_n1488# 0.642782f
C131 source.n0 a_n2102_n1488# 0.876971f
C132 source.t4 a_n2102_n1488# 0.077408f
C133 source.t2 a_n2102_n1488# 0.077408f
C134 source.n1 a_n2102_n1488# 0.490811f
C135 source.n2 a_n2102_n1488# 0.398724f
C136 source.t13 a_n2102_n1488# 0.077408f
C137 source.t6 a_n2102_n1488# 0.077408f
C138 source.n3 a_n2102_n1488# 0.490811f
C139 source.n4 a_n2102_n1488# 0.398724f
C140 source.t16 a_n2102_n1488# 0.077408f
C141 source.t38 a_n2102_n1488# 0.077408f
C142 source.n5 a_n2102_n1488# 0.490811f
C143 source.n6 a_n2102_n1488# 0.398724f
C144 source.t3 a_n2102_n1488# 0.077408f
C145 source.t7 a_n2102_n1488# 0.077408f
C146 source.n7 a_n2102_n1488# 0.490811f
C147 source.n8 a_n2102_n1488# 0.398724f
C148 source.t14 a_n2102_n1488# 0.642782f
C149 source.n9 a_n2102_n1488# 0.450156f
C150 source.t25 a_n2102_n1488# 0.642782f
C151 source.n10 a_n2102_n1488# 0.450156f
C152 source.t33 a_n2102_n1488# 0.077408f
C153 source.t21 a_n2102_n1488# 0.077408f
C154 source.n11 a_n2102_n1488# 0.490811f
C155 source.n12 a_n2102_n1488# 0.398724f
C156 source.t22 a_n2102_n1488# 0.077408f
C157 source.t26 a_n2102_n1488# 0.077408f
C158 source.n13 a_n2102_n1488# 0.490811f
C159 source.n14 a_n2102_n1488# 0.398724f
C160 source.t30 a_n2102_n1488# 0.077408f
C161 source.t35 a_n2102_n1488# 0.077408f
C162 source.n15 a_n2102_n1488# 0.490811f
C163 source.n16 a_n2102_n1488# 0.398724f
C164 source.t32 a_n2102_n1488# 0.077408f
C165 source.t20 a_n2102_n1488# 0.077408f
C166 source.n17 a_n2102_n1488# 0.490811f
C167 source.n18 a_n2102_n1488# 0.398724f
C168 source.t29 a_n2102_n1488# 0.642782f
C169 source.n19 a_n2102_n1488# 1.21732f
C170 source.t11 a_n2102_n1488# 0.642779f
C171 source.n20 a_n2102_n1488# 1.21733f
C172 source.t1 a_n2102_n1488# 0.077408f
C173 source.t10 a_n2102_n1488# 0.077408f
C174 source.n21 a_n2102_n1488# 0.490808f
C175 source.n22 a_n2102_n1488# 0.398728f
C176 source.t0 a_n2102_n1488# 0.077408f
C177 source.t17 a_n2102_n1488# 0.077408f
C178 source.n23 a_n2102_n1488# 0.490808f
C179 source.n24 a_n2102_n1488# 0.398728f
C180 source.t8 a_n2102_n1488# 0.077408f
C181 source.t39 a_n2102_n1488# 0.077408f
C182 source.n25 a_n2102_n1488# 0.490808f
C183 source.n26 a_n2102_n1488# 0.398728f
C184 source.t9 a_n2102_n1488# 0.077408f
C185 source.t5 a_n2102_n1488# 0.077408f
C186 source.n27 a_n2102_n1488# 0.490808f
C187 source.n28 a_n2102_n1488# 0.398728f
C188 source.t15 a_n2102_n1488# 0.642779f
C189 source.n29 a_n2102_n1488# 0.45016f
C190 source.t28 a_n2102_n1488# 0.642779f
C191 source.n30 a_n2102_n1488# 0.45016f
C192 source.t36 a_n2102_n1488# 0.077408f
C193 source.t18 a_n2102_n1488# 0.077408f
C194 source.n31 a_n2102_n1488# 0.490808f
C195 source.n32 a_n2102_n1488# 0.398728f
C196 source.t27 a_n2102_n1488# 0.077408f
C197 source.t31 a_n2102_n1488# 0.077408f
C198 source.n33 a_n2102_n1488# 0.490808f
C199 source.n34 a_n2102_n1488# 0.398728f
C200 source.t34 a_n2102_n1488# 0.077408f
C201 source.t23 a_n2102_n1488# 0.077408f
C202 source.n35 a_n2102_n1488# 0.490808f
C203 source.n36 a_n2102_n1488# 0.398728f
C204 source.t24 a_n2102_n1488# 0.077408f
C205 source.t37 a_n2102_n1488# 0.077408f
C206 source.n37 a_n2102_n1488# 0.490808f
C207 source.n38 a_n2102_n1488# 0.398728f
C208 source.t19 a_n2102_n1488# 0.642779f
C209 source.n39 a_n2102_n1488# 0.63448f
C210 source.n40 a_n2102_n1488# 0.946426f
C211 drain_right.t5 a_n2102_n1488# 0.076623f
C212 drain_right.t3 a_n2102_n1488# 0.076623f
C213 drain_right.n0 a_n2102_n1488# 0.5552f
C214 drain_right.t19 a_n2102_n1488# 0.076623f
C215 drain_right.t1 a_n2102_n1488# 0.076623f
C216 drain_right.n1 a_n2102_n1488# 0.552597f
C217 drain_right.n2 a_n2102_n1488# 0.749883f
C218 drain_right.t4 a_n2102_n1488# 0.076623f
C219 drain_right.t6 a_n2102_n1488# 0.076623f
C220 drain_right.n3 a_n2102_n1488# 0.552597f
C221 drain_right.t2 a_n2102_n1488# 0.076623f
C222 drain_right.t18 a_n2102_n1488# 0.076623f
C223 drain_right.n4 a_n2102_n1488# 0.5552f
C224 drain_right.t14 a_n2102_n1488# 0.076623f
C225 drain_right.t13 a_n2102_n1488# 0.076623f
C226 drain_right.n5 a_n2102_n1488# 0.552597f
C227 drain_right.n6 a_n2102_n1488# 0.749883f
C228 drain_right.n7 a_n2102_n1488# 1.31574f
C229 drain_right.t16 a_n2102_n1488# 0.076623f
C230 drain_right.t11 a_n2102_n1488# 0.076623f
C231 drain_right.n8 a_n2102_n1488# 0.555202f
C232 drain_right.t12 a_n2102_n1488# 0.076623f
C233 drain_right.t0 a_n2102_n1488# 0.076623f
C234 drain_right.n9 a_n2102_n1488# 0.5526f
C235 drain_right.n10 a_n2102_n1488# 0.754106f
C236 drain_right.t9 a_n2102_n1488# 0.076623f
C237 drain_right.t15 a_n2102_n1488# 0.076623f
C238 drain_right.n11 a_n2102_n1488# 0.5526f
C239 drain_right.n12 a_n2102_n1488# 0.371845f
C240 drain_right.t17 a_n2102_n1488# 0.076623f
C241 drain_right.t8 a_n2102_n1488# 0.076623f
C242 drain_right.n13 a_n2102_n1488# 0.5526f
C243 drain_right.n14 a_n2102_n1488# 0.371845f
C244 drain_right.t10 a_n2102_n1488# 0.076623f
C245 drain_right.t7 a_n2102_n1488# 0.076623f
C246 drain_right.n15 a_n2102_n1488# 0.5526f
C247 drain_right.n16 a_n2102_n1488# 0.640872f
C248 minus.n0 a_n2102_n1488# 0.049352f
C249 minus.t8 a_n2102_n1488# 0.138401f
C250 minus.t5 a_n2102_n1488# 0.128624f
C251 minus.t17 a_n2102_n1488# 0.128624f
C252 minus.n1 a_n2102_n1488# 0.018045f
C253 minus.n2 a_n2102_n1488# 0.049352f
C254 minus.t7 a_n2102_n1488# 0.128624f
C255 minus.n3 a_n2102_n1488# 0.074685f
C256 minus.t2 a_n2102_n1488# 0.128624f
C257 minus.t15 a_n2102_n1488# 0.128624f
C258 minus.t11 a_n2102_n1488# 0.128624f
C259 minus.n4 a_n2102_n1488# 0.074685f
C260 minus.n5 a_n2102_n1488# 0.049352f
C261 minus.t4 a_n2102_n1488# 0.128624f
C262 minus.t16 a_n2102_n1488# 0.128624f
C263 minus.n6 a_n2102_n1488# 0.074685f
C264 minus.t12 a_n2102_n1488# 0.138401f
C265 minus.n7 a_n2102_n1488# 0.089418f
C266 minus.n8 a_n2102_n1488# 0.112929f
C267 minus.n9 a_n2102_n1488# 0.020327f
C268 minus.n10 a_n2102_n1488# 0.074685f
C269 minus.n11 a_n2102_n1488# 0.018654f
C270 minus.n12 a_n2102_n1488# 0.018045f
C271 minus.n13 a_n2102_n1488# 0.049352f
C272 minus.n14 a_n2102_n1488# 0.049352f
C273 minus.n15 a_n2102_n1488# 0.020327f
C274 minus.n16 a_n2102_n1488# 0.074685f
C275 minus.n17 a_n2102_n1488# 0.020327f
C276 minus.n18 a_n2102_n1488# 0.074685f
C277 minus.n19 a_n2102_n1488# 0.020327f
C278 minus.n20 a_n2102_n1488# 0.049352f
C279 minus.n21 a_n2102_n1488# 0.049352f
C280 minus.n22 a_n2102_n1488# 0.049352f
C281 minus.n23 a_n2102_n1488# 0.018654f
C282 minus.n24 a_n2102_n1488# 0.074685f
C283 minus.n25 a_n2102_n1488# 0.020327f
C284 minus.n26 a_n2102_n1488# 0.074685f
C285 minus.n27 a_n2102_n1488# 0.089344f
C286 minus.n28 a_n2102_n1488# 1.30509f
C287 minus.n29 a_n2102_n1488# 0.049352f
C288 minus.t0 a_n2102_n1488# 0.128624f
C289 minus.t13 a_n2102_n1488# 0.128624f
C290 minus.n30 a_n2102_n1488# 0.018045f
C291 minus.n31 a_n2102_n1488# 0.049352f
C292 minus.t3 a_n2102_n1488# 0.128624f
C293 minus.t6 a_n2102_n1488# 0.128624f
C294 minus.t10 a_n2102_n1488# 0.128624f
C295 minus.n32 a_n2102_n1488# 0.074685f
C296 minus.n33 a_n2102_n1488# 0.049352f
C297 minus.t19 a_n2102_n1488# 0.128624f
C298 minus.t1 a_n2102_n1488# 0.128624f
C299 minus.n34 a_n2102_n1488# 0.074685f
C300 minus.t9 a_n2102_n1488# 0.138401f
C301 minus.n35 a_n2102_n1488# 0.089418f
C302 minus.n36 a_n2102_n1488# 0.112929f
C303 minus.n37 a_n2102_n1488# 0.020327f
C304 minus.n38 a_n2102_n1488# 0.074685f
C305 minus.n39 a_n2102_n1488# 0.018654f
C306 minus.n40 a_n2102_n1488# 0.018045f
C307 minus.n41 a_n2102_n1488# 0.049352f
C308 minus.n42 a_n2102_n1488# 0.049352f
C309 minus.n43 a_n2102_n1488# 0.020327f
C310 minus.n44 a_n2102_n1488# 0.074685f
C311 minus.n45 a_n2102_n1488# 0.020327f
C312 minus.n46 a_n2102_n1488# 0.074685f
C313 minus.t14 a_n2102_n1488# 0.128624f
C314 minus.n47 a_n2102_n1488# 0.074685f
C315 minus.n48 a_n2102_n1488# 0.020327f
C316 minus.n49 a_n2102_n1488# 0.049352f
C317 minus.n50 a_n2102_n1488# 0.049352f
C318 minus.n51 a_n2102_n1488# 0.049352f
C319 minus.n52 a_n2102_n1488# 0.018654f
C320 minus.n53 a_n2102_n1488# 0.074685f
C321 minus.n54 a_n2102_n1488# 0.020327f
C322 minus.n55 a_n2102_n1488# 0.074685f
C323 minus.t18 a_n2102_n1488# 0.138401f
C324 minus.n56 a_n2102_n1488# 0.089344f
C325 minus.n57 a_n2102_n1488# 0.324466f
C326 minus.n58 a_n2102_n1488# 1.60841f
.ends

