* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t16 minus.t0 drain_right.t4 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 source.t5 plus.t0 drain_left.t9 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 drain_left.t8 plus.t1 source.t4 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X3 a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X4 drain_left.t7 plus.t2 source.t0 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X5 a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X6 drain_right.t5 minus.t1 source.t15 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X7 a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X8 drain_right.t6 minus.t2 source.t14 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X9 source.t13 minus.t3 drain_right.t0 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 source.t2 plus.t3 drain_left.t6 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X11 drain_right.t9 minus.t4 source.t12 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X12 drain_right.t1 minus.t5 source.t11 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X13 source.t10 minus.t6 drain_right.t8 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X14 drain_left.t5 plus.t4 source.t3 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X15 drain_left.t4 plus.t5 source.t6 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X16 drain_right.t2 minus.t7 source.t9 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X18 source.t1 plus.t6 drain_left.t3 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X19 source.t8 minus.t8 drain_right.t3 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X20 drain_left.t2 plus.t7 source.t17 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X21 source.t18 plus.t8 drain_left.t1 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X22 drain_right.t7 minus.t9 source.t7 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 drain_left.t0 plus.t9 source.t19 a_n1496_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
R0 minus.n9 minus.t5 734.686
R1 minus.n3 minus.t4 734.686
R2 minus.n20 minus.t1 734.686
R3 minus.n14 minus.t2 734.686
R4 minus.n6 minus.t7 690.867
R5 minus.n8 minus.t6 690.867
R6 minus.n2 minus.t3 690.867
R7 minus.n17 minus.t9 690.867
R8 minus.n19 minus.t8 690.867
R9 minus.n13 minus.t0 690.867
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 27.9835
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t6 90.3333
R42 drain_right.n7 drain_right.t1 89.7731
R43 drain_right.n6 drain_right.n4 80.3335
R44 drain_right.n3 drain_right.n2 80.1379
R45 drain_right.n6 drain_right.n5 79.7731
R46 drain_right.n1 drain_right.n0 79.773
R47 drain_right drain_right.n3 22.3771
R48 drain_right.n2 drain_right.t3 10.0005
R49 drain_right.n2 drain_right.t5 10.0005
R50 drain_right.n0 drain_right.t4 10.0005
R51 drain_right.n0 drain_right.t7 10.0005
R52 drain_right.n4 drain_right.t0 10.0005
R53 drain_right.n4 drain_right.t9 10.0005
R54 drain_right.n5 drain_right.t8 10.0005
R55 drain_right.n5 drain_right.t2 10.0005
R56 drain_right drain_right.n7 5.93339
R57 drain_right.n7 drain_right.n6 0.560845
R58 drain_right.n3 drain_right.n1 0.0852402
R59 source.n0 source.t19 73.0943
R60 source.n5 source.t12 73.0943
R61 source.n19 source.t15 73.0942
R62 source.n14 source.t4 73.0942
R63 source.n2 source.n1 63.0943
R64 source.n4 source.n3 63.0943
R65 source.n7 source.n6 63.0943
R66 source.n9 source.n8 63.0943
R67 source.n18 source.n17 63.0942
R68 source.n16 source.n15 63.0942
R69 source.n13 source.n12 63.0942
R70 source.n11 source.n10 63.0942
R71 source.n11 source.n9 15.5902
R72 source.n17 source.t7 10.0005
R73 source.n17 source.t8 10.0005
R74 source.n15 source.t14 10.0005
R75 source.n15 source.t16 10.0005
R76 source.n12 source.t3 10.0005
R77 source.n12 source.t5 10.0005
R78 source.n10 source.t0 10.0005
R79 source.n10 source.t2 10.0005
R80 source.n1 source.t17 10.0005
R81 source.n1 source.t1 10.0005
R82 source.n3 source.t6 10.0005
R83 source.n3 source.t18 10.0005
R84 source.n6 source.t9 10.0005
R85 source.n6 source.t13 10.0005
R86 source.n8 source.t11 10.0005
R87 source.n8 source.t10 10.0005
R88 source.n20 source.n0 9.48679
R89 source.n20 source.n19 5.5436
R90 source.n5 source.n4 0.7505
R91 source.n16 source.n14 0.7505
R92 source.n9 source.n7 0.560845
R93 source.n7 source.n5 0.560845
R94 source.n4 source.n2 0.560845
R95 source.n2 source.n0 0.560845
R96 source.n13 source.n11 0.560845
R97 source.n14 source.n13 0.560845
R98 source.n18 source.n16 0.560845
R99 source.n19 source.n18 0.560845
R100 source source.n20 0.188
R101 plus.n3 plus.t5 734.686
R102 plus.n9 plus.t9 734.686
R103 plus.n14 plus.t1 734.686
R104 plus.n20 plus.t2 734.686
R105 plus.n6 plus.t7 690.867
R106 plus.n2 plus.t8 690.867
R107 plus.n8 plus.t6 690.867
R108 plus.n17 plus.t4 690.867
R109 plus.n13 plus.t0 690.867
R110 plus.n19 plus.t3 690.867
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 25.2736
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 8.74861
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t4 90.3335
R142 drain_left.n1 drain_left.t7 90.3333
R143 drain_left.n3 drain_left.n2 80.1379
R144 drain_left.n7 drain_left.n6 79.7731
R145 drain_left.n5 drain_left.n4 79.7731
R146 drain_left.n1 drain_left.n0 79.773
R147 drain_left drain_left.n3 22.9304
R148 drain_left.n2 drain_left.t9 10.0005
R149 drain_left.n2 drain_left.t8 10.0005
R150 drain_left.n0 drain_left.t6 10.0005
R151 drain_left.n0 drain_left.t5 10.0005
R152 drain_left.n6 drain_left.t3 10.0005
R153 drain_left.n6 drain_left.t0 10.0005
R154 drain_left.n4 drain_left.t1 10.0005
R155 drain_left.n4 drain_left.t2 10.0005
R156 drain_left drain_left.n7 6.21356
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 source minus 0.900587f
C1 drain_right source 7.0048f
C2 plus drain_left 1.0608f
C3 drain_right minus 0.918547f
C4 source plus 0.914746f
C5 plus minus 3.34346f
C6 drain_right plus 0.302579f
C7 source drain_left 7.00838f
C8 minus drain_left 0.175926f
C9 drain_right drain_left 0.73287f
C10 drain_right a_n1496_n1488# 3.78252f
C11 drain_left a_n1496_n1488# 3.99639f
C12 source a_n1496_n1488# 2.868021f
C13 minus a_n1496_n1488# 4.787551f
C14 plus a_n1496_n1488# 5.605807f
C15 drain_left.t7 a_n1496_n1488# 0.522463f
C16 drain_left.t6 a_n1496_n1488# 0.079562f
C17 drain_left.t5 a_n1496_n1488# 0.079562f
C18 drain_left.n0 a_n1496_n1488# 0.432807f
C19 drain_left.n1 a_n1496_n1488# 0.509188f
C20 drain_left.t9 a_n1496_n1488# 0.079562f
C21 drain_left.t8 a_n1496_n1488# 0.079562f
C22 drain_left.n2 a_n1496_n1488# 0.433962f
C23 drain_left.n3 a_n1496_n1488# 0.844081f
C24 drain_left.t4 a_n1496_n1488# 0.522465f
C25 drain_left.t1 a_n1496_n1488# 0.079562f
C26 drain_left.t2 a_n1496_n1488# 0.079562f
C27 drain_left.n4 a_n1496_n1488# 0.432809f
C28 drain_left.n5 a_n1496_n1488# 0.53707f
C29 drain_left.t3 a_n1496_n1488# 0.079562f
C30 drain_left.t0 a_n1496_n1488# 0.079562f
C31 drain_left.n6 a_n1496_n1488# 0.432809f
C32 drain_left.n7 a_n1496_n1488# 0.44227f
C33 plus.n0 a_n1496_n1488# 0.036207f
C34 plus.t6 a_n1496_n1488# 0.047184f
C35 plus.t7 a_n1496_n1488# 0.047184f
C36 plus.n1 a_n1496_n1488# 0.01536f
C37 plus.t5 a_n1496_n1488# 0.049084f
C38 plus.t8 a_n1496_n1488# 0.047184f
C39 plus.n2 a_n1496_n1488# 0.032978f
C40 plus.n3 a_n1496_n1488# 0.04537f
C41 plus.n4 a_n1496_n1488# 0.077947f
C42 plus.n5 a_n1496_n1488# 0.036207f
C43 plus.n6 a_n1496_n1488# 0.044989f
C44 plus.n7 a_n1496_n1488# 0.01536f
C45 plus.n8 a_n1496_n1488# 0.032978f
C46 plus.t9 a_n1496_n1488# 0.049084f
C47 plus.n9 a_n1496_n1488# 0.045321f
C48 plus.n10 a_n1496_n1488# 0.2717f
C49 plus.n11 a_n1496_n1488# 0.036207f
C50 plus.t2 a_n1496_n1488# 0.049084f
C51 plus.t3 a_n1496_n1488# 0.047184f
C52 plus.t4 a_n1496_n1488# 0.047184f
C53 plus.n12 a_n1496_n1488# 0.01536f
C54 plus.t0 a_n1496_n1488# 0.047184f
C55 plus.n13 a_n1496_n1488# 0.032978f
C56 plus.t1 a_n1496_n1488# 0.049084f
C57 plus.n14 a_n1496_n1488# 0.04537f
C58 plus.n15 a_n1496_n1488# 0.077947f
C59 plus.n16 a_n1496_n1488# 0.036207f
C60 plus.n17 a_n1496_n1488# 0.044989f
C61 plus.n18 a_n1496_n1488# 0.01536f
C62 plus.n19 a_n1496_n1488# 0.032978f
C63 plus.n20 a_n1496_n1488# 0.045321f
C64 plus.n21 a_n1496_n1488# 0.787762f
C65 source.t19 a_n1496_n1488# 0.54608f
C66 source.n0 a_n1496_n1488# 0.720894f
C67 source.t17 a_n1496_n1488# 0.092717f
C68 source.t1 a_n1496_n1488# 0.092717f
C69 source.n1 a_n1496_n1488# 0.451046f
C70 source.n2 a_n1496_n1488# 0.318069f
C71 source.t6 a_n1496_n1488# 0.092717f
C72 source.t18 a_n1496_n1488# 0.092717f
C73 source.n3 a_n1496_n1488# 0.451046f
C74 source.n4 a_n1496_n1488# 0.333843f
C75 source.t12 a_n1496_n1488# 0.54608f
C76 source.n5 a_n1496_n1488# 0.405699f
C77 source.t9 a_n1496_n1488# 0.092717f
C78 source.t13 a_n1496_n1488# 0.092717f
C79 source.n6 a_n1496_n1488# 0.451046f
C80 source.n7 a_n1496_n1488# 0.318069f
C81 source.t11 a_n1496_n1488# 0.092717f
C82 source.t10 a_n1496_n1488# 0.092717f
C83 source.n8 a_n1496_n1488# 0.451046f
C84 source.n9 a_n1496_n1488# 0.965045f
C85 source.t0 a_n1496_n1488# 0.092717f
C86 source.t2 a_n1496_n1488# 0.092717f
C87 source.n10 a_n1496_n1488# 0.451043f
C88 source.n11 a_n1496_n1488# 0.965048f
C89 source.t3 a_n1496_n1488# 0.092717f
C90 source.t5 a_n1496_n1488# 0.092717f
C91 source.n12 a_n1496_n1488# 0.451043f
C92 source.n13 a_n1496_n1488# 0.318072f
C93 source.t4 a_n1496_n1488# 0.546077f
C94 source.n14 a_n1496_n1488# 0.405701f
C95 source.t14 a_n1496_n1488# 0.092717f
C96 source.t16 a_n1496_n1488# 0.092717f
C97 source.n15 a_n1496_n1488# 0.451043f
C98 source.n16 a_n1496_n1488# 0.333846f
C99 source.t7 a_n1496_n1488# 0.092717f
C100 source.t8 a_n1496_n1488# 0.092717f
C101 source.n17 a_n1496_n1488# 0.451043f
C102 source.n18 a_n1496_n1488# 0.318072f
C103 source.t15 a_n1496_n1488# 0.546077f
C104 source.n19 a_n1496_n1488# 0.529254f
C105 source.n20 a_n1496_n1488# 0.748804f
C106 drain_right.t6 a_n1496_n1488# 0.529012f
C107 drain_right.t4 a_n1496_n1488# 0.080559f
C108 drain_right.t7 a_n1496_n1488# 0.080559f
C109 drain_right.n0 a_n1496_n1488# 0.438231f
C110 drain_right.n1 a_n1496_n1488# 0.51557f
C111 drain_right.t3 a_n1496_n1488# 0.080559f
C112 drain_right.t5 a_n1496_n1488# 0.080559f
C113 drain_right.n2 a_n1496_n1488# 0.439401f
C114 drain_right.n3 a_n1496_n1488# 0.810024f
C115 drain_right.t0 a_n1496_n1488# 0.080559f
C116 drain_right.t9 a_n1496_n1488# 0.080559f
C117 drain_right.n4 a_n1496_n1488# 0.440113f
C118 drain_right.t8 a_n1496_n1488# 0.080559f
C119 drain_right.t2 a_n1496_n1488# 0.080559f
C120 drain_right.n5 a_n1496_n1488# 0.438233f
C121 drain_right.n6 a_n1496_n1488# 0.528189f
C122 drain_right.t1 a_n1496_n1488# 0.527245f
C123 drain_right.n7 a_n1496_n1488# 0.473114f
C124 minus.n0 a_n1496_n1488# 0.035422f
C125 minus.t5 a_n1496_n1488# 0.048019f
C126 minus.t6 a_n1496_n1488# 0.04616f
C127 minus.t7 a_n1496_n1488# 0.04616f
C128 minus.n1 a_n1496_n1488# 0.015026f
C129 minus.t3 a_n1496_n1488# 0.04616f
C130 minus.n2 a_n1496_n1488# 0.032262f
C131 minus.t4 a_n1496_n1488# 0.048019f
C132 minus.n3 a_n1496_n1488# 0.044385f
C133 minus.n4 a_n1496_n1488# 0.076255f
C134 minus.n5 a_n1496_n1488# 0.035422f
C135 minus.n6 a_n1496_n1488# 0.044013f
C136 minus.n7 a_n1496_n1488# 0.015026f
C137 minus.n8 a_n1496_n1488# 0.032262f
C138 minus.n9 a_n1496_n1488# 0.044337f
C139 minus.n10 a_n1496_n1488# 0.816941f
C140 minus.n11 a_n1496_n1488# 0.035422f
C141 minus.t8 a_n1496_n1488# 0.04616f
C142 minus.t9 a_n1496_n1488# 0.04616f
C143 minus.n12 a_n1496_n1488# 0.015026f
C144 minus.t2 a_n1496_n1488# 0.048019f
C145 minus.t0 a_n1496_n1488# 0.04616f
C146 minus.n13 a_n1496_n1488# 0.032262f
C147 minus.n14 a_n1496_n1488# 0.044385f
C148 minus.n15 a_n1496_n1488# 0.076255f
C149 minus.n16 a_n1496_n1488# 0.035422f
C150 minus.n17 a_n1496_n1488# 0.044013f
C151 minus.n18 a_n1496_n1488# 0.015026f
C152 minus.n19 a_n1496_n1488# 0.032262f
C153 minus.t1 a_n1496_n1488# 0.048019f
C154 minus.n20 a_n1496_n1488# 0.044337f
C155 minus.n21 a_n1496_n1488# 0.232724f
C156 minus.n22 a_n1496_n1488# 1.00923f
.ends

