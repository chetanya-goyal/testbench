* NGSPICE file created from diffpair281.ext - technology: sky130A

.subckt diffpair281 minus drain_right drain_left source plus
X0 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X1 source minus drain_right a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X2 source plus drain_left a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X3 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X4 drain_left plus source a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X5 source plus drain_left a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X6 drain_right minus source a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X7 drain_left plus source a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X8 drain_right minus source a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X9 source minus drain_right a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X10 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X11 a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# a_n1214_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
.ends

