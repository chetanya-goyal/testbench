* NGSPICE file created from diffpair419.ext - technology: sky130A

.subckt diffpair419 minus drain_right drain_left source plus
X0 a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X1 source.t30 plus.t0 drain_left.t15 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X2 drain_right.t23 minus.t0 source.t40 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X3 drain_right.t22 minus.t1 source.t46 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X4 source.t45 minus.t2 drain_right.t21 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X5 source.t42 minus.t3 drain_right.t20 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X6 source.t41 minus.t4 drain_right.t19 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X7 a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X8 source.t35 minus.t5 drain_right.t18 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X9 drain_right.t17 minus.t6 source.t5 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X10 source.t29 plus.t1 drain_left.t14 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X11 drain_left.t13 plus.t2 source.t28 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X12 drain_right.t16 minus.t7 source.t32 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X13 drain_right.t15 minus.t8 source.t36 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X14 drain_right.t14 minus.t9 source.t0 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X15 drain_right.t13 minus.t10 source.t1 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X16 drain_right.t12 minus.t11 source.t4 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X17 source.t31 minus.t12 drain_right.t11 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X18 source.t3 minus.t13 drain_right.t10 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X19 drain_left.t4 plus.t3 source.t27 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X20 source.t33 minus.t14 drain_right.t9 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X21 source.t38 minus.t15 drain_right.t8 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X22 drain_right.t7 minus.t16 source.t6 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X23 source.t43 minus.t17 drain_right.t6 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X24 source.t26 plus.t4 drain_left.t3 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X25 drain_left.t10 plus.t5 source.t25 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X26 source.t24 plus.t6 drain_left.t9 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X27 a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X28 source.t47 minus.t18 drain_right.t5 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X29 drain_left.t23 plus.t7 source.t23 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X30 a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X31 drain_right.t4 minus.t19 source.t37 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X32 drain_right.t3 minus.t20 source.t2 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X33 drain_right.t2 minus.t21 source.t44 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X34 drain_left.t22 plus.t8 source.t22 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X35 source.t21 plus.t9 drain_left.t8 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X36 source.t20 plus.t10 drain_left.t7 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X37 source.t19 plus.t11 drain_left.t6 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X38 source.t18 plus.t12 drain_left.t5 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X39 source.t17 plus.t13 drain_left.t17 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X40 drain_left.t16 plus.t14 source.t16 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X41 source.t15 plus.t15 drain_left.t12 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X42 drain_left.t11 plus.t16 source.t14 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X43 drain_left.t19 plus.t17 source.t13 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X44 drain_left.t18 plus.t18 source.t12 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X45 source.t34 minus.t22 drain_right.t1 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X46 source.t39 minus.t23 drain_right.t0 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X47 drain_left.t21 plus.t19 source.t11 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X48 drain_left.t20 plus.t20 source.t10 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X49 drain_left.t1 plus.t21 source.t9 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X50 source.t8 plus.t22 drain_left.t0 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X51 source.t7 plus.t23 drain_left.t2 a_n2094_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 plus.n6 plus.t6 1663.27
R1 plus.n29 plus.t20 1663.27
R2 plus.n37 plus.t19 1663.27
R3 plus.n60 plus.t15 1663.27
R4 plus.n7 plus.t2 1602.65
R5 plus.n5 plus.t22 1602.65
R6 plus.n12 plus.t14 1602.65
R7 plus.n14 plus.t13 1602.65
R8 plus.n3 plus.t5 1602.65
R9 plus.n19 plus.t1 1602.65
R10 plus.n21 plus.t21 1602.65
R11 plus.n1 plus.t11 1602.65
R12 plus.n26 plus.t3 1602.65
R13 plus.n28 plus.t0 1602.65
R14 plus.n38 plus.t23 1602.65
R15 plus.n36 plus.t17 1602.65
R16 plus.n43 plus.t12 1602.65
R17 plus.n45 plus.t18 1602.65
R18 plus.n34 plus.t9 1602.65
R19 plus.n50 plus.t16 1602.65
R20 plus.n52 plus.t10 1602.65
R21 plus.n32 plus.t7 1602.65
R22 plus.n57 plus.t4 1602.65
R23 plus.n59 plus.t8 1602.65
R24 plus.n9 plus.n6 161.489
R25 plus.n40 plus.n37 161.489
R26 plus.n9 plus.n8 161.3
R27 plus.n11 plus.n10 161.3
R28 plus.n13 plus.n4 161.3
R29 plus.n16 plus.n15 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n2 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n0 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n40 plus.n39 161.3
R37 plus.n42 plus.n41 161.3
R38 plus.n44 plus.n35 161.3
R39 plus.n47 plus.n46 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n33 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n31 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n8 plus.n7 56.2338
R47 plus.n28 plus.n27 56.2338
R48 plus.n59 plus.n58 56.2338
R49 plus.n39 plus.n38 56.2338
R50 plus.n11 plus.n5 51.852
R51 plus.n26 plus.n25 51.852
R52 plus.n57 plus.n56 51.852
R53 plus.n42 plus.n36 51.852
R54 plus.n13 plus.n12 47.4702
R55 plus.n22 plus.n1 47.4702
R56 plus.n53 plus.n32 47.4702
R57 plus.n44 plus.n43 47.4702
R58 plus.n15 plus.n14 43.0884
R59 plus.n21 plus.n20 43.0884
R60 plus.n52 plus.n51 43.0884
R61 plus.n46 plus.n45 43.0884
R62 plus.n18 plus.n3 38.7066
R63 plus.n19 plus.n18 38.7066
R64 plus.n50 plus.n49 38.7066
R65 plus.n49 plus.n34 38.7066
R66 plus.n15 plus.n3 34.3247
R67 plus.n20 plus.n19 34.3247
R68 plus.n51 plus.n50 34.3247
R69 plus.n46 plus.n34 34.3247
R70 plus plus.n61 30.9233
R71 plus.n14 plus.n13 29.9429
R72 plus.n22 plus.n21 29.9429
R73 plus.n53 plus.n52 29.9429
R74 plus.n45 plus.n44 29.9429
R75 plus.n12 plus.n11 25.5611
R76 plus.n25 plus.n1 25.5611
R77 plus.n56 plus.n32 25.5611
R78 plus.n43 plus.n42 25.5611
R79 plus.n8 plus.n5 21.1793
R80 plus.n27 plus.n26 21.1793
R81 plus.n58 plus.n57 21.1793
R82 plus.n39 plus.n36 21.1793
R83 plus.n7 plus.n6 16.7975
R84 plus.n29 plus.n28 16.7975
R85 plus.n60 plus.n59 16.7975
R86 plus.n38 plus.n37 16.7975
R87 plus plus.n30 12.1331
R88 plus.n10 plus.n9 0.189894
R89 plus.n10 plus.n4 0.189894
R90 plus.n16 plus.n4 0.189894
R91 plus.n17 plus.n16 0.189894
R92 plus.n17 plus.n2 0.189894
R93 plus.n23 plus.n2 0.189894
R94 plus.n24 plus.n23 0.189894
R95 plus.n24 plus.n0 0.189894
R96 plus.n30 plus.n0 0.189894
R97 plus.n61 plus.n31 0.189894
R98 plus.n55 plus.n31 0.189894
R99 plus.n55 plus.n54 0.189894
R100 plus.n54 plus.n33 0.189894
R101 plus.n48 plus.n33 0.189894
R102 plus.n48 plus.n47 0.189894
R103 plus.n47 plus.n35 0.189894
R104 plus.n41 plus.n35 0.189894
R105 plus.n41 plus.n40 0.189894
R106 drain_left.n13 drain_left.n11 60.0096
R107 drain_left.n7 drain_left.n5 60.0094
R108 drain_left.n2 drain_left.n0 60.0094
R109 drain_left.n19 drain_left.n18 59.5527
R110 drain_left.n17 drain_left.n16 59.5527
R111 drain_left.n15 drain_left.n14 59.5527
R112 drain_left.n13 drain_left.n12 59.5527
R113 drain_left.n7 drain_left.n6 59.5525
R114 drain_left.n9 drain_left.n8 59.5525
R115 drain_left.n4 drain_left.n3 59.5525
R116 drain_left.n2 drain_left.n1 59.5525
R117 drain_left.n21 drain_left.n20 59.5525
R118 drain_left drain_left.n10 31.7076
R119 drain_left drain_left.n21 6.11011
R120 drain_left.n5 drain_left.t2 1.6505
R121 drain_left.n5 drain_left.t21 1.6505
R122 drain_left.n6 drain_left.t5 1.6505
R123 drain_left.n6 drain_left.t19 1.6505
R124 drain_left.n8 drain_left.t8 1.6505
R125 drain_left.n8 drain_left.t18 1.6505
R126 drain_left.n3 drain_left.t7 1.6505
R127 drain_left.n3 drain_left.t11 1.6505
R128 drain_left.n1 drain_left.t3 1.6505
R129 drain_left.n1 drain_left.t23 1.6505
R130 drain_left.n0 drain_left.t12 1.6505
R131 drain_left.n0 drain_left.t22 1.6505
R132 drain_left.n20 drain_left.t15 1.6505
R133 drain_left.n20 drain_left.t20 1.6505
R134 drain_left.n18 drain_left.t6 1.6505
R135 drain_left.n18 drain_left.t4 1.6505
R136 drain_left.n16 drain_left.t14 1.6505
R137 drain_left.n16 drain_left.t1 1.6505
R138 drain_left.n14 drain_left.t17 1.6505
R139 drain_left.n14 drain_left.t10 1.6505
R140 drain_left.n12 drain_left.t0 1.6505
R141 drain_left.n12 drain_left.t16 1.6505
R142 drain_left.n11 drain_left.t9 1.6505
R143 drain_left.n11 drain_left.t13 1.6505
R144 drain_left.n9 drain_left.n7 0.457397
R145 drain_left.n4 drain_left.n2 0.457397
R146 drain_left.n15 drain_left.n13 0.457397
R147 drain_left.n17 drain_left.n15 0.457397
R148 drain_left.n19 drain_left.n17 0.457397
R149 drain_left.n21 drain_left.n19 0.457397
R150 drain_left.n10 drain_left.n9 0.173602
R151 drain_left.n10 drain_left.n4 0.173602
R152 source.n562 source.n502 289.615
R153 source.n486 source.n426 289.615
R154 source.n420 source.n360 289.615
R155 source.n344 source.n284 289.615
R156 source.n60 source.n0 289.615
R157 source.n136 source.n76 289.615
R158 source.n202 source.n142 289.615
R159 source.n278 source.n218 289.615
R160 source.n522 source.n521 185
R161 source.n527 source.n526 185
R162 source.n529 source.n528 185
R163 source.n518 source.n517 185
R164 source.n535 source.n534 185
R165 source.n537 source.n536 185
R166 source.n514 source.n513 185
R167 source.n544 source.n543 185
R168 source.n545 source.n512 185
R169 source.n547 source.n546 185
R170 source.n510 source.n509 185
R171 source.n553 source.n552 185
R172 source.n555 source.n554 185
R173 source.n506 source.n505 185
R174 source.n561 source.n560 185
R175 source.n563 source.n562 185
R176 source.n446 source.n445 185
R177 source.n451 source.n450 185
R178 source.n453 source.n452 185
R179 source.n442 source.n441 185
R180 source.n459 source.n458 185
R181 source.n461 source.n460 185
R182 source.n438 source.n437 185
R183 source.n468 source.n467 185
R184 source.n469 source.n436 185
R185 source.n471 source.n470 185
R186 source.n434 source.n433 185
R187 source.n477 source.n476 185
R188 source.n479 source.n478 185
R189 source.n430 source.n429 185
R190 source.n485 source.n484 185
R191 source.n487 source.n486 185
R192 source.n380 source.n379 185
R193 source.n385 source.n384 185
R194 source.n387 source.n386 185
R195 source.n376 source.n375 185
R196 source.n393 source.n392 185
R197 source.n395 source.n394 185
R198 source.n372 source.n371 185
R199 source.n402 source.n401 185
R200 source.n403 source.n370 185
R201 source.n405 source.n404 185
R202 source.n368 source.n367 185
R203 source.n411 source.n410 185
R204 source.n413 source.n412 185
R205 source.n364 source.n363 185
R206 source.n419 source.n418 185
R207 source.n421 source.n420 185
R208 source.n304 source.n303 185
R209 source.n309 source.n308 185
R210 source.n311 source.n310 185
R211 source.n300 source.n299 185
R212 source.n317 source.n316 185
R213 source.n319 source.n318 185
R214 source.n296 source.n295 185
R215 source.n326 source.n325 185
R216 source.n327 source.n294 185
R217 source.n329 source.n328 185
R218 source.n292 source.n291 185
R219 source.n335 source.n334 185
R220 source.n337 source.n336 185
R221 source.n288 source.n287 185
R222 source.n343 source.n342 185
R223 source.n345 source.n344 185
R224 source.n61 source.n60 185
R225 source.n59 source.n58 185
R226 source.n4 source.n3 185
R227 source.n53 source.n52 185
R228 source.n51 source.n50 185
R229 source.n8 source.n7 185
R230 source.n45 source.n44 185
R231 source.n43 source.n10 185
R232 source.n42 source.n41 185
R233 source.n13 source.n11 185
R234 source.n36 source.n35 185
R235 source.n34 source.n33 185
R236 source.n17 source.n16 185
R237 source.n28 source.n27 185
R238 source.n26 source.n25 185
R239 source.n21 source.n20 185
R240 source.n137 source.n136 185
R241 source.n135 source.n134 185
R242 source.n80 source.n79 185
R243 source.n129 source.n128 185
R244 source.n127 source.n126 185
R245 source.n84 source.n83 185
R246 source.n121 source.n120 185
R247 source.n119 source.n86 185
R248 source.n118 source.n117 185
R249 source.n89 source.n87 185
R250 source.n112 source.n111 185
R251 source.n110 source.n109 185
R252 source.n93 source.n92 185
R253 source.n104 source.n103 185
R254 source.n102 source.n101 185
R255 source.n97 source.n96 185
R256 source.n203 source.n202 185
R257 source.n201 source.n200 185
R258 source.n146 source.n145 185
R259 source.n195 source.n194 185
R260 source.n193 source.n192 185
R261 source.n150 source.n149 185
R262 source.n187 source.n186 185
R263 source.n185 source.n152 185
R264 source.n184 source.n183 185
R265 source.n155 source.n153 185
R266 source.n178 source.n177 185
R267 source.n176 source.n175 185
R268 source.n159 source.n158 185
R269 source.n170 source.n169 185
R270 source.n168 source.n167 185
R271 source.n163 source.n162 185
R272 source.n279 source.n278 185
R273 source.n277 source.n276 185
R274 source.n222 source.n221 185
R275 source.n271 source.n270 185
R276 source.n269 source.n268 185
R277 source.n226 source.n225 185
R278 source.n263 source.n262 185
R279 source.n261 source.n228 185
R280 source.n260 source.n259 185
R281 source.n231 source.n229 185
R282 source.n254 source.n253 185
R283 source.n252 source.n251 185
R284 source.n235 source.n234 185
R285 source.n246 source.n245 185
R286 source.n244 source.n243 185
R287 source.n239 source.n238 185
R288 source.n523 source.t5 149.524
R289 source.n447 source.t41 149.524
R290 source.n381 source.t11 149.524
R291 source.n305 source.t15 149.524
R292 source.n22 source.t10 149.524
R293 source.n98 source.t24 149.524
R294 source.n164 source.t2 149.524
R295 source.n240 source.t35 149.524
R296 source.n527 source.n521 104.615
R297 source.n528 source.n527 104.615
R298 source.n528 source.n517 104.615
R299 source.n535 source.n517 104.615
R300 source.n536 source.n535 104.615
R301 source.n536 source.n513 104.615
R302 source.n544 source.n513 104.615
R303 source.n545 source.n544 104.615
R304 source.n546 source.n545 104.615
R305 source.n546 source.n509 104.615
R306 source.n553 source.n509 104.615
R307 source.n554 source.n553 104.615
R308 source.n554 source.n505 104.615
R309 source.n561 source.n505 104.615
R310 source.n562 source.n561 104.615
R311 source.n451 source.n445 104.615
R312 source.n452 source.n451 104.615
R313 source.n452 source.n441 104.615
R314 source.n459 source.n441 104.615
R315 source.n460 source.n459 104.615
R316 source.n460 source.n437 104.615
R317 source.n468 source.n437 104.615
R318 source.n469 source.n468 104.615
R319 source.n470 source.n469 104.615
R320 source.n470 source.n433 104.615
R321 source.n477 source.n433 104.615
R322 source.n478 source.n477 104.615
R323 source.n478 source.n429 104.615
R324 source.n485 source.n429 104.615
R325 source.n486 source.n485 104.615
R326 source.n385 source.n379 104.615
R327 source.n386 source.n385 104.615
R328 source.n386 source.n375 104.615
R329 source.n393 source.n375 104.615
R330 source.n394 source.n393 104.615
R331 source.n394 source.n371 104.615
R332 source.n402 source.n371 104.615
R333 source.n403 source.n402 104.615
R334 source.n404 source.n403 104.615
R335 source.n404 source.n367 104.615
R336 source.n411 source.n367 104.615
R337 source.n412 source.n411 104.615
R338 source.n412 source.n363 104.615
R339 source.n419 source.n363 104.615
R340 source.n420 source.n419 104.615
R341 source.n309 source.n303 104.615
R342 source.n310 source.n309 104.615
R343 source.n310 source.n299 104.615
R344 source.n317 source.n299 104.615
R345 source.n318 source.n317 104.615
R346 source.n318 source.n295 104.615
R347 source.n326 source.n295 104.615
R348 source.n327 source.n326 104.615
R349 source.n328 source.n327 104.615
R350 source.n328 source.n291 104.615
R351 source.n335 source.n291 104.615
R352 source.n336 source.n335 104.615
R353 source.n336 source.n287 104.615
R354 source.n343 source.n287 104.615
R355 source.n344 source.n343 104.615
R356 source.n60 source.n59 104.615
R357 source.n59 source.n3 104.615
R358 source.n52 source.n3 104.615
R359 source.n52 source.n51 104.615
R360 source.n51 source.n7 104.615
R361 source.n44 source.n7 104.615
R362 source.n44 source.n43 104.615
R363 source.n43 source.n42 104.615
R364 source.n42 source.n11 104.615
R365 source.n35 source.n11 104.615
R366 source.n35 source.n34 104.615
R367 source.n34 source.n16 104.615
R368 source.n27 source.n16 104.615
R369 source.n27 source.n26 104.615
R370 source.n26 source.n20 104.615
R371 source.n136 source.n135 104.615
R372 source.n135 source.n79 104.615
R373 source.n128 source.n79 104.615
R374 source.n128 source.n127 104.615
R375 source.n127 source.n83 104.615
R376 source.n120 source.n83 104.615
R377 source.n120 source.n119 104.615
R378 source.n119 source.n118 104.615
R379 source.n118 source.n87 104.615
R380 source.n111 source.n87 104.615
R381 source.n111 source.n110 104.615
R382 source.n110 source.n92 104.615
R383 source.n103 source.n92 104.615
R384 source.n103 source.n102 104.615
R385 source.n102 source.n96 104.615
R386 source.n202 source.n201 104.615
R387 source.n201 source.n145 104.615
R388 source.n194 source.n145 104.615
R389 source.n194 source.n193 104.615
R390 source.n193 source.n149 104.615
R391 source.n186 source.n149 104.615
R392 source.n186 source.n185 104.615
R393 source.n185 source.n184 104.615
R394 source.n184 source.n153 104.615
R395 source.n177 source.n153 104.615
R396 source.n177 source.n176 104.615
R397 source.n176 source.n158 104.615
R398 source.n169 source.n158 104.615
R399 source.n169 source.n168 104.615
R400 source.n168 source.n162 104.615
R401 source.n278 source.n277 104.615
R402 source.n277 source.n221 104.615
R403 source.n270 source.n221 104.615
R404 source.n270 source.n269 104.615
R405 source.n269 source.n225 104.615
R406 source.n262 source.n225 104.615
R407 source.n262 source.n261 104.615
R408 source.n261 source.n260 104.615
R409 source.n260 source.n229 104.615
R410 source.n253 source.n229 104.615
R411 source.n253 source.n252 104.615
R412 source.n252 source.n234 104.615
R413 source.n245 source.n234 104.615
R414 source.n245 source.n244 104.615
R415 source.n244 source.n238 104.615
R416 source.t5 source.n521 52.3082
R417 source.t41 source.n445 52.3082
R418 source.t11 source.n379 52.3082
R419 source.t15 source.n303 52.3082
R420 source.t10 source.n20 52.3082
R421 source.t24 source.n96 52.3082
R422 source.t2 source.n162 52.3082
R423 source.t35 source.n238 52.3082
R424 source.n67 source.n66 42.8739
R425 source.n69 source.n68 42.8739
R426 source.n71 source.n70 42.8739
R427 source.n73 source.n72 42.8739
R428 source.n75 source.n74 42.8739
R429 source.n209 source.n208 42.8739
R430 source.n211 source.n210 42.8739
R431 source.n213 source.n212 42.8739
R432 source.n215 source.n214 42.8739
R433 source.n217 source.n216 42.8739
R434 source.n501 source.n500 42.8737
R435 source.n499 source.n498 42.8737
R436 source.n497 source.n496 42.8737
R437 source.n495 source.n494 42.8737
R438 source.n493 source.n492 42.8737
R439 source.n359 source.n358 42.8737
R440 source.n357 source.n356 42.8737
R441 source.n355 source.n354 42.8737
R442 source.n353 source.n352 42.8737
R443 source.n351 source.n350 42.8737
R444 source.n567 source.n566 29.8581
R445 source.n491 source.n490 29.8581
R446 source.n425 source.n424 29.8581
R447 source.n349 source.n348 29.8581
R448 source.n65 source.n64 29.8581
R449 source.n141 source.n140 29.8581
R450 source.n207 source.n206 29.8581
R451 source.n283 source.n282 29.8581
R452 source.n349 source.n283 21.7446
R453 source.n568 source.n65 16.2532
R454 source.n547 source.n512 13.1884
R455 source.n471 source.n436 13.1884
R456 source.n405 source.n370 13.1884
R457 source.n329 source.n294 13.1884
R458 source.n45 source.n10 13.1884
R459 source.n121 source.n86 13.1884
R460 source.n187 source.n152 13.1884
R461 source.n263 source.n228 13.1884
R462 source.n543 source.n542 12.8005
R463 source.n548 source.n510 12.8005
R464 source.n467 source.n466 12.8005
R465 source.n472 source.n434 12.8005
R466 source.n401 source.n400 12.8005
R467 source.n406 source.n368 12.8005
R468 source.n325 source.n324 12.8005
R469 source.n330 source.n292 12.8005
R470 source.n46 source.n8 12.8005
R471 source.n41 source.n12 12.8005
R472 source.n122 source.n84 12.8005
R473 source.n117 source.n88 12.8005
R474 source.n188 source.n150 12.8005
R475 source.n183 source.n154 12.8005
R476 source.n264 source.n226 12.8005
R477 source.n259 source.n230 12.8005
R478 source.n541 source.n514 12.0247
R479 source.n552 source.n551 12.0247
R480 source.n465 source.n438 12.0247
R481 source.n476 source.n475 12.0247
R482 source.n399 source.n372 12.0247
R483 source.n410 source.n409 12.0247
R484 source.n323 source.n296 12.0247
R485 source.n334 source.n333 12.0247
R486 source.n50 source.n49 12.0247
R487 source.n40 source.n13 12.0247
R488 source.n126 source.n125 12.0247
R489 source.n116 source.n89 12.0247
R490 source.n192 source.n191 12.0247
R491 source.n182 source.n155 12.0247
R492 source.n268 source.n267 12.0247
R493 source.n258 source.n231 12.0247
R494 source.n538 source.n537 11.249
R495 source.n555 source.n508 11.249
R496 source.n462 source.n461 11.249
R497 source.n479 source.n432 11.249
R498 source.n396 source.n395 11.249
R499 source.n413 source.n366 11.249
R500 source.n320 source.n319 11.249
R501 source.n337 source.n290 11.249
R502 source.n53 source.n6 11.249
R503 source.n37 source.n36 11.249
R504 source.n129 source.n82 11.249
R505 source.n113 source.n112 11.249
R506 source.n195 source.n148 11.249
R507 source.n179 source.n178 11.249
R508 source.n271 source.n224 11.249
R509 source.n255 source.n254 11.249
R510 source.n534 source.n516 10.4732
R511 source.n556 source.n506 10.4732
R512 source.n458 source.n440 10.4732
R513 source.n480 source.n430 10.4732
R514 source.n392 source.n374 10.4732
R515 source.n414 source.n364 10.4732
R516 source.n316 source.n298 10.4732
R517 source.n338 source.n288 10.4732
R518 source.n54 source.n4 10.4732
R519 source.n33 source.n15 10.4732
R520 source.n130 source.n80 10.4732
R521 source.n109 source.n91 10.4732
R522 source.n196 source.n146 10.4732
R523 source.n175 source.n157 10.4732
R524 source.n272 source.n222 10.4732
R525 source.n251 source.n233 10.4732
R526 source.n523 source.n522 10.2747
R527 source.n447 source.n446 10.2747
R528 source.n381 source.n380 10.2747
R529 source.n305 source.n304 10.2747
R530 source.n22 source.n21 10.2747
R531 source.n98 source.n97 10.2747
R532 source.n164 source.n163 10.2747
R533 source.n240 source.n239 10.2747
R534 source.n533 source.n518 9.69747
R535 source.n560 source.n559 9.69747
R536 source.n457 source.n442 9.69747
R537 source.n484 source.n483 9.69747
R538 source.n391 source.n376 9.69747
R539 source.n418 source.n417 9.69747
R540 source.n315 source.n300 9.69747
R541 source.n342 source.n341 9.69747
R542 source.n58 source.n57 9.69747
R543 source.n32 source.n17 9.69747
R544 source.n134 source.n133 9.69747
R545 source.n108 source.n93 9.69747
R546 source.n200 source.n199 9.69747
R547 source.n174 source.n159 9.69747
R548 source.n276 source.n275 9.69747
R549 source.n250 source.n235 9.69747
R550 source.n566 source.n565 9.45567
R551 source.n490 source.n489 9.45567
R552 source.n424 source.n423 9.45567
R553 source.n348 source.n347 9.45567
R554 source.n64 source.n63 9.45567
R555 source.n140 source.n139 9.45567
R556 source.n206 source.n205 9.45567
R557 source.n282 source.n281 9.45567
R558 source.n565 source.n564 9.3005
R559 source.n504 source.n503 9.3005
R560 source.n559 source.n558 9.3005
R561 source.n557 source.n556 9.3005
R562 source.n508 source.n507 9.3005
R563 source.n551 source.n550 9.3005
R564 source.n549 source.n548 9.3005
R565 source.n525 source.n524 9.3005
R566 source.n520 source.n519 9.3005
R567 source.n531 source.n530 9.3005
R568 source.n533 source.n532 9.3005
R569 source.n516 source.n515 9.3005
R570 source.n539 source.n538 9.3005
R571 source.n541 source.n540 9.3005
R572 source.n542 source.n511 9.3005
R573 source.n489 source.n488 9.3005
R574 source.n428 source.n427 9.3005
R575 source.n483 source.n482 9.3005
R576 source.n481 source.n480 9.3005
R577 source.n432 source.n431 9.3005
R578 source.n475 source.n474 9.3005
R579 source.n473 source.n472 9.3005
R580 source.n449 source.n448 9.3005
R581 source.n444 source.n443 9.3005
R582 source.n455 source.n454 9.3005
R583 source.n457 source.n456 9.3005
R584 source.n440 source.n439 9.3005
R585 source.n463 source.n462 9.3005
R586 source.n465 source.n464 9.3005
R587 source.n466 source.n435 9.3005
R588 source.n423 source.n422 9.3005
R589 source.n362 source.n361 9.3005
R590 source.n417 source.n416 9.3005
R591 source.n415 source.n414 9.3005
R592 source.n366 source.n365 9.3005
R593 source.n409 source.n408 9.3005
R594 source.n407 source.n406 9.3005
R595 source.n383 source.n382 9.3005
R596 source.n378 source.n377 9.3005
R597 source.n389 source.n388 9.3005
R598 source.n391 source.n390 9.3005
R599 source.n374 source.n373 9.3005
R600 source.n397 source.n396 9.3005
R601 source.n399 source.n398 9.3005
R602 source.n400 source.n369 9.3005
R603 source.n347 source.n346 9.3005
R604 source.n286 source.n285 9.3005
R605 source.n341 source.n340 9.3005
R606 source.n339 source.n338 9.3005
R607 source.n290 source.n289 9.3005
R608 source.n333 source.n332 9.3005
R609 source.n331 source.n330 9.3005
R610 source.n307 source.n306 9.3005
R611 source.n302 source.n301 9.3005
R612 source.n313 source.n312 9.3005
R613 source.n315 source.n314 9.3005
R614 source.n298 source.n297 9.3005
R615 source.n321 source.n320 9.3005
R616 source.n323 source.n322 9.3005
R617 source.n324 source.n293 9.3005
R618 source.n24 source.n23 9.3005
R619 source.n19 source.n18 9.3005
R620 source.n30 source.n29 9.3005
R621 source.n32 source.n31 9.3005
R622 source.n15 source.n14 9.3005
R623 source.n38 source.n37 9.3005
R624 source.n40 source.n39 9.3005
R625 source.n12 source.n9 9.3005
R626 source.n63 source.n62 9.3005
R627 source.n2 source.n1 9.3005
R628 source.n57 source.n56 9.3005
R629 source.n55 source.n54 9.3005
R630 source.n6 source.n5 9.3005
R631 source.n49 source.n48 9.3005
R632 source.n47 source.n46 9.3005
R633 source.n100 source.n99 9.3005
R634 source.n95 source.n94 9.3005
R635 source.n106 source.n105 9.3005
R636 source.n108 source.n107 9.3005
R637 source.n91 source.n90 9.3005
R638 source.n114 source.n113 9.3005
R639 source.n116 source.n115 9.3005
R640 source.n88 source.n85 9.3005
R641 source.n139 source.n138 9.3005
R642 source.n78 source.n77 9.3005
R643 source.n133 source.n132 9.3005
R644 source.n131 source.n130 9.3005
R645 source.n82 source.n81 9.3005
R646 source.n125 source.n124 9.3005
R647 source.n123 source.n122 9.3005
R648 source.n166 source.n165 9.3005
R649 source.n161 source.n160 9.3005
R650 source.n172 source.n171 9.3005
R651 source.n174 source.n173 9.3005
R652 source.n157 source.n156 9.3005
R653 source.n180 source.n179 9.3005
R654 source.n182 source.n181 9.3005
R655 source.n154 source.n151 9.3005
R656 source.n205 source.n204 9.3005
R657 source.n144 source.n143 9.3005
R658 source.n199 source.n198 9.3005
R659 source.n197 source.n196 9.3005
R660 source.n148 source.n147 9.3005
R661 source.n191 source.n190 9.3005
R662 source.n189 source.n188 9.3005
R663 source.n242 source.n241 9.3005
R664 source.n237 source.n236 9.3005
R665 source.n248 source.n247 9.3005
R666 source.n250 source.n249 9.3005
R667 source.n233 source.n232 9.3005
R668 source.n256 source.n255 9.3005
R669 source.n258 source.n257 9.3005
R670 source.n230 source.n227 9.3005
R671 source.n281 source.n280 9.3005
R672 source.n220 source.n219 9.3005
R673 source.n275 source.n274 9.3005
R674 source.n273 source.n272 9.3005
R675 source.n224 source.n223 9.3005
R676 source.n267 source.n266 9.3005
R677 source.n265 source.n264 9.3005
R678 source.n530 source.n529 8.92171
R679 source.n563 source.n504 8.92171
R680 source.n454 source.n453 8.92171
R681 source.n487 source.n428 8.92171
R682 source.n388 source.n387 8.92171
R683 source.n421 source.n362 8.92171
R684 source.n312 source.n311 8.92171
R685 source.n345 source.n286 8.92171
R686 source.n61 source.n2 8.92171
R687 source.n29 source.n28 8.92171
R688 source.n137 source.n78 8.92171
R689 source.n105 source.n104 8.92171
R690 source.n203 source.n144 8.92171
R691 source.n171 source.n170 8.92171
R692 source.n279 source.n220 8.92171
R693 source.n247 source.n246 8.92171
R694 source.n526 source.n520 8.14595
R695 source.n564 source.n502 8.14595
R696 source.n450 source.n444 8.14595
R697 source.n488 source.n426 8.14595
R698 source.n384 source.n378 8.14595
R699 source.n422 source.n360 8.14595
R700 source.n308 source.n302 8.14595
R701 source.n346 source.n284 8.14595
R702 source.n62 source.n0 8.14595
R703 source.n25 source.n19 8.14595
R704 source.n138 source.n76 8.14595
R705 source.n101 source.n95 8.14595
R706 source.n204 source.n142 8.14595
R707 source.n167 source.n161 8.14595
R708 source.n280 source.n218 8.14595
R709 source.n243 source.n237 8.14595
R710 source.n525 source.n522 7.3702
R711 source.n449 source.n446 7.3702
R712 source.n383 source.n380 7.3702
R713 source.n307 source.n304 7.3702
R714 source.n24 source.n21 7.3702
R715 source.n100 source.n97 7.3702
R716 source.n166 source.n163 7.3702
R717 source.n242 source.n239 7.3702
R718 source.n526 source.n525 5.81868
R719 source.n566 source.n502 5.81868
R720 source.n450 source.n449 5.81868
R721 source.n490 source.n426 5.81868
R722 source.n384 source.n383 5.81868
R723 source.n424 source.n360 5.81868
R724 source.n308 source.n307 5.81868
R725 source.n348 source.n284 5.81868
R726 source.n64 source.n0 5.81868
R727 source.n25 source.n24 5.81868
R728 source.n140 source.n76 5.81868
R729 source.n101 source.n100 5.81868
R730 source.n206 source.n142 5.81868
R731 source.n167 source.n166 5.81868
R732 source.n282 source.n218 5.81868
R733 source.n243 source.n242 5.81868
R734 source.n568 source.n567 5.49188
R735 source.n529 source.n520 5.04292
R736 source.n564 source.n563 5.04292
R737 source.n453 source.n444 5.04292
R738 source.n488 source.n487 5.04292
R739 source.n387 source.n378 5.04292
R740 source.n422 source.n421 5.04292
R741 source.n311 source.n302 5.04292
R742 source.n346 source.n345 5.04292
R743 source.n62 source.n61 5.04292
R744 source.n28 source.n19 5.04292
R745 source.n138 source.n137 5.04292
R746 source.n104 source.n95 5.04292
R747 source.n204 source.n203 5.04292
R748 source.n170 source.n161 5.04292
R749 source.n280 source.n279 5.04292
R750 source.n246 source.n237 5.04292
R751 source.n530 source.n518 4.26717
R752 source.n560 source.n504 4.26717
R753 source.n454 source.n442 4.26717
R754 source.n484 source.n428 4.26717
R755 source.n388 source.n376 4.26717
R756 source.n418 source.n362 4.26717
R757 source.n312 source.n300 4.26717
R758 source.n342 source.n286 4.26717
R759 source.n58 source.n2 4.26717
R760 source.n29 source.n17 4.26717
R761 source.n134 source.n78 4.26717
R762 source.n105 source.n93 4.26717
R763 source.n200 source.n144 4.26717
R764 source.n171 source.n159 4.26717
R765 source.n276 source.n220 4.26717
R766 source.n247 source.n235 4.26717
R767 source.n534 source.n533 3.49141
R768 source.n559 source.n506 3.49141
R769 source.n458 source.n457 3.49141
R770 source.n483 source.n430 3.49141
R771 source.n392 source.n391 3.49141
R772 source.n417 source.n364 3.49141
R773 source.n316 source.n315 3.49141
R774 source.n341 source.n288 3.49141
R775 source.n57 source.n4 3.49141
R776 source.n33 source.n32 3.49141
R777 source.n133 source.n80 3.49141
R778 source.n109 source.n108 3.49141
R779 source.n199 source.n146 3.49141
R780 source.n175 source.n174 3.49141
R781 source.n275 source.n222 3.49141
R782 source.n251 source.n250 3.49141
R783 source.n524 source.n523 2.84303
R784 source.n448 source.n447 2.84303
R785 source.n382 source.n381 2.84303
R786 source.n306 source.n305 2.84303
R787 source.n23 source.n22 2.84303
R788 source.n99 source.n98 2.84303
R789 source.n165 source.n164 2.84303
R790 source.n241 source.n240 2.84303
R791 source.n537 source.n516 2.71565
R792 source.n556 source.n555 2.71565
R793 source.n461 source.n440 2.71565
R794 source.n480 source.n479 2.71565
R795 source.n395 source.n374 2.71565
R796 source.n414 source.n413 2.71565
R797 source.n319 source.n298 2.71565
R798 source.n338 source.n337 2.71565
R799 source.n54 source.n53 2.71565
R800 source.n36 source.n15 2.71565
R801 source.n130 source.n129 2.71565
R802 source.n112 source.n91 2.71565
R803 source.n196 source.n195 2.71565
R804 source.n178 source.n157 2.71565
R805 source.n272 source.n271 2.71565
R806 source.n254 source.n233 2.71565
R807 source.n538 source.n514 1.93989
R808 source.n552 source.n508 1.93989
R809 source.n462 source.n438 1.93989
R810 source.n476 source.n432 1.93989
R811 source.n396 source.n372 1.93989
R812 source.n410 source.n366 1.93989
R813 source.n320 source.n296 1.93989
R814 source.n334 source.n290 1.93989
R815 source.n50 source.n6 1.93989
R816 source.n37 source.n13 1.93989
R817 source.n126 source.n82 1.93989
R818 source.n113 source.n89 1.93989
R819 source.n192 source.n148 1.93989
R820 source.n179 source.n155 1.93989
R821 source.n268 source.n224 1.93989
R822 source.n255 source.n231 1.93989
R823 source.n500 source.t32 1.6505
R824 source.n500 source.t45 1.6505
R825 source.n498 source.t1 1.6505
R826 source.n498 source.t33 1.6505
R827 source.n496 source.t4 1.6505
R828 source.n496 source.t43 1.6505
R829 source.n494 source.t36 1.6505
R830 source.n494 source.t47 1.6505
R831 source.n492 source.t0 1.6505
R832 source.n492 source.t42 1.6505
R833 source.n358 source.t13 1.6505
R834 source.n358 source.t7 1.6505
R835 source.n356 source.t12 1.6505
R836 source.n356 source.t18 1.6505
R837 source.n354 source.t14 1.6505
R838 source.n354 source.t21 1.6505
R839 source.n352 source.t23 1.6505
R840 source.n352 source.t20 1.6505
R841 source.n350 source.t22 1.6505
R842 source.n350 source.t26 1.6505
R843 source.n66 source.t27 1.6505
R844 source.n66 source.t30 1.6505
R845 source.n68 source.t9 1.6505
R846 source.n68 source.t19 1.6505
R847 source.n70 source.t25 1.6505
R848 source.n70 source.t29 1.6505
R849 source.n72 source.t16 1.6505
R850 source.n72 source.t17 1.6505
R851 source.n74 source.t28 1.6505
R852 source.n74 source.t8 1.6505
R853 source.n208 source.t40 1.6505
R854 source.n208 source.t3 1.6505
R855 source.n210 source.t44 1.6505
R856 source.n210 source.t34 1.6505
R857 source.n212 source.t46 1.6505
R858 source.n212 source.t31 1.6505
R859 source.n214 source.t37 1.6505
R860 source.n214 source.t39 1.6505
R861 source.n216 source.t6 1.6505
R862 source.n216 source.t38 1.6505
R863 source.n543 source.n541 1.16414
R864 source.n551 source.n510 1.16414
R865 source.n467 source.n465 1.16414
R866 source.n475 source.n434 1.16414
R867 source.n401 source.n399 1.16414
R868 source.n409 source.n368 1.16414
R869 source.n325 source.n323 1.16414
R870 source.n333 source.n292 1.16414
R871 source.n49 source.n8 1.16414
R872 source.n41 source.n40 1.16414
R873 source.n125 source.n84 1.16414
R874 source.n117 source.n116 1.16414
R875 source.n191 source.n150 1.16414
R876 source.n183 source.n182 1.16414
R877 source.n267 source.n226 1.16414
R878 source.n259 source.n258 1.16414
R879 source.n207 source.n141 0.470328
R880 source.n491 source.n425 0.470328
R881 source.n283 source.n217 0.457397
R882 source.n217 source.n215 0.457397
R883 source.n215 source.n213 0.457397
R884 source.n213 source.n211 0.457397
R885 source.n211 source.n209 0.457397
R886 source.n209 source.n207 0.457397
R887 source.n141 source.n75 0.457397
R888 source.n75 source.n73 0.457397
R889 source.n73 source.n71 0.457397
R890 source.n71 source.n69 0.457397
R891 source.n69 source.n67 0.457397
R892 source.n67 source.n65 0.457397
R893 source.n351 source.n349 0.457397
R894 source.n353 source.n351 0.457397
R895 source.n355 source.n353 0.457397
R896 source.n357 source.n355 0.457397
R897 source.n359 source.n357 0.457397
R898 source.n425 source.n359 0.457397
R899 source.n493 source.n491 0.457397
R900 source.n495 source.n493 0.457397
R901 source.n497 source.n495 0.457397
R902 source.n499 source.n497 0.457397
R903 source.n501 source.n499 0.457397
R904 source.n567 source.n501 0.457397
R905 source.n542 source.n512 0.388379
R906 source.n548 source.n547 0.388379
R907 source.n466 source.n436 0.388379
R908 source.n472 source.n471 0.388379
R909 source.n400 source.n370 0.388379
R910 source.n406 source.n405 0.388379
R911 source.n324 source.n294 0.388379
R912 source.n330 source.n329 0.388379
R913 source.n46 source.n45 0.388379
R914 source.n12 source.n10 0.388379
R915 source.n122 source.n121 0.388379
R916 source.n88 source.n86 0.388379
R917 source.n188 source.n187 0.388379
R918 source.n154 source.n152 0.388379
R919 source.n264 source.n263 0.388379
R920 source.n230 source.n228 0.388379
R921 source source.n568 0.188
R922 source.n524 source.n519 0.155672
R923 source.n531 source.n519 0.155672
R924 source.n532 source.n531 0.155672
R925 source.n532 source.n515 0.155672
R926 source.n539 source.n515 0.155672
R927 source.n540 source.n539 0.155672
R928 source.n540 source.n511 0.155672
R929 source.n549 source.n511 0.155672
R930 source.n550 source.n549 0.155672
R931 source.n550 source.n507 0.155672
R932 source.n557 source.n507 0.155672
R933 source.n558 source.n557 0.155672
R934 source.n558 source.n503 0.155672
R935 source.n565 source.n503 0.155672
R936 source.n448 source.n443 0.155672
R937 source.n455 source.n443 0.155672
R938 source.n456 source.n455 0.155672
R939 source.n456 source.n439 0.155672
R940 source.n463 source.n439 0.155672
R941 source.n464 source.n463 0.155672
R942 source.n464 source.n435 0.155672
R943 source.n473 source.n435 0.155672
R944 source.n474 source.n473 0.155672
R945 source.n474 source.n431 0.155672
R946 source.n481 source.n431 0.155672
R947 source.n482 source.n481 0.155672
R948 source.n482 source.n427 0.155672
R949 source.n489 source.n427 0.155672
R950 source.n382 source.n377 0.155672
R951 source.n389 source.n377 0.155672
R952 source.n390 source.n389 0.155672
R953 source.n390 source.n373 0.155672
R954 source.n397 source.n373 0.155672
R955 source.n398 source.n397 0.155672
R956 source.n398 source.n369 0.155672
R957 source.n407 source.n369 0.155672
R958 source.n408 source.n407 0.155672
R959 source.n408 source.n365 0.155672
R960 source.n415 source.n365 0.155672
R961 source.n416 source.n415 0.155672
R962 source.n416 source.n361 0.155672
R963 source.n423 source.n361 0.155672
R964 source.n306 source.n301 0.155672
R965 source.n313 source.n301 0.155672
R966 source.n314 source.n313 0.155672
R967 source.n314 source.n297 0.155672
R968 source.n321 source.n297 0.155672
R969 source.n322 source.n321 0.155672
R970 source.n322 source.n293 0.155672
R971 source.n331 source.n293 0.155672
R972 source.n332 source.n331 0.155672
R973 source.n332 source.n289 0.155672
R974 source.n339 source.n289 0.155672
R975 source.n340 source.n339 0.155672
R976 source.n340 source.n285 0.155672
R977 source.n347 source.n285 0.155672
R978 source.n63 source.n1 0.155672
R979 source.n56 source.n1 0.155672
R980 source.n56 source.n55 0.155672
R981 source.n55 source.n5 0.155672
R982 source.n48 source.n5 0.155672
R983 source.n48 source.n47 0.155672
R984 source.n47 source.n9 0.155672
R985 source.n39 source.n9 0.155672
R986 source.n39 source.n38 0.155672
R987 source.n38 source.n14 0.155672
R988 source.n31 source.n14 0.155672
R989 source.n31 source.n30 0.155672
R990 source.n30 source.n18 0.155672
R991 source.n23 source.n18 0.155672
R992 source.n139 source.n77 0.155672
R993 source.n132 source.n77 0.155672
R994 source.n132 source.n131 0.155672
R995 source.n131 source.n81 0.155672
R996 source.n124 source.n81 0.155672
R997 source.n124 source.n123 0.155672
R998 source.n123 source.n85 0.155672
R999 source.n115 source.n85 0.155672
R1000 source.n115 source.n114 0.155672
R1001 source.n114 source.n90 0.155672
R1002 source.n107 source.n90 0.155672
R1003 source.n107 source.n106 0.155672
R1004 source.n106 source.n94 0.155672
R1005 source.n99 source.n94 0.155672
R1006 source.n205 source.n143 0.155672
R1007 source.n198 source.n143 0.155672
R1008 source.n198 source.n197 0.155672
R1009 source.n197 source.n147 0.155672
R1010 source.n190 source.n147 0.155672
R1011 source.n190 source.n189 0.155672
R1012 source.n189 source.n151 0.155672
R1013 source.n181 source.n151 0.155672
R1014 source.n181 source.n180 0.155672
R1015 source.n180 source.n156 0.155672
R1016 source.n173 source.n156 0.155672
R1017 source.n173 source.n172 0.155672
R1018 source.n172 source.n160 0.155672
R1019 source.n165 source.n160 0.155672
R1020 source.n281 source.n219 0.155672
R1021 source.n274 source.n219 0.155672
R1022 source.n274 source.n273 0.155672
R1023 source.n273 source.n223 0.155672
R1024 source.n266 source.n223 0.155672
R1025 source.n266 source.n265 0.155672
R1026 source.n265 source.n227 0.155672
R1027 source.n257 source.n227 0.155672
R1028 source.n257 source.n256 0.155672
R1029 source.n256 source.n232 0.155672
R1030 source.n249 source.n232 0.155672
R1031 source.n249 source.n248 0.155672
R1032 source.n248 source.n236 0.155672
R1033 source.n241 source.n236 0.155672
R1034 minus.n29 minus.t5 1663.27
R1035 minus.n6 minus.t20 1663.27
R1036 minus.n60 minus.t6 1663.27
R1037 minus.n37 minus.t4 1663.27
R1038 minus.n28 minus.t16 1602.65
R1039 minus.n26 minus.t15 1602.65
R1040 minus.n1 minus.t19 1602.65
R1041 minus.n21 minus.t23 1602.65
R1042 minus.n19 minus.t1 1602.65
R1043 minus.n3 minus.t12 1602.65
R1044 minus.n14 minus.t21 1602.65
R1045 minus.n12 minus.t22 1602.65
R1046 minus.n5 minus.t0 1602.65
R1047 minus.n7 minus.t13 1602.65
R1048 minus.n59 minus.t2 1602.65
R1049 minus.n57 minus.t7 1602.65
R1050 minus.n32 minus.t14 1602.65
R1051 minus.n52 minus.t10 1602.65
R1052 minus.n50 minus.t17 1602.65
R1053 minus.n34 minus.t11 1602.65
R1054 minus.n45 minus.t18 1602.65
R1055 minus.n43 minus.t8 1602.65
R1056 minus.n36 minus.t3 1602.65
R1057 minus.n38 minus.t9 1602.65
R1058 minus.n9 minus.n6 161.489
R1059 minus.n40 minus.n37 161.489
R1060 minus.n30 minus.n29 161.3
R1061 minus.n27 minus.n0 161.3
R1062 minus.n25 minus.n24 161.3
R1063 minus.n23 minus.n22 161.3
R1064 minus.n20 minus.n2 161.3
R1065 minus.n18 minus.n17 161.3
R1066 minus.n16 minus.n15 161.3
R1067 minus.n13 minus.n4 161.3
R1068 minus.n11 minus.n10 161.3
R1069 minus.n9 minus.n8 161.3
R1070 minus.n61 minus.n60 161.3
R1071 minus.n58 minus.n31 161.3
R1072 minus.n56 minus.n55 161.3
R1073 minus.n54 minus.n53 161.3
R1074 minus.n51 minus.n33 161.3
R1075 minus.n49 minus.n48 161.3
R1076 minus.n47 minus.n46 161.3
R1077 minus.n44 minus.n35 161.3
R1078 minus.n42 minus.n41 161.3
R1079 minus.n40 minus.n39 161.3
R1080 minus.n28 minus.n27 56.2338
R1081 minus.n8 minus.n7 56.2338
R1082 minus.n39 minus.n38 56.2338
R1083 minus.n59 minus.n58 56.2338
R1084 minus.n26 minus.n25 51.852
R1085 minus.n11 minus.n5 51.852
R1086 minus.n42 minus.n36 51.852
R1087 minus.n57 minus.n56 51.852
R1088 minus.n22 minus.n1 47.4702
R1089 minus.n13 minus.n12 47.4702
R1090 minus.n44 minus.n43 47.4702
R1091 minus.n53 minus.n32 47.4702
R1092 minus.n21 minus.n20 43.0884
R1093 minus.n15 minus.n14 43.0884
R1094 minus.n46 minus.n45 43.0884
R1095 minus.n52 minus.n51 43.0884
R1096 minus.n19 minus.n18 38.7066
R1097 minus.n18 minus.n3 38.7066
R1098 minus.n49 minus.n34 38.7066
R1099 minus.n50 minus.n49 38.7066
R1100 minus.n62 minus.n30 37.0422
R1101 minus.n20 minus.n19 34.3247
R1102 minus.n15 minus.n3 34.3247
R1103 minus.n46 minus.n34 34.3247
R1104 minus.n51 minus.n50 34.3247
R1105 minus.n22 minus.n21 29.9429
R1106 minus.n14 minus.n13 29.9429
R1107 minus.n45 minus.n44 29.9429
R1108 minus.n53 minus.n52 29.9429
R1109 minus.n25 minus.n1 25.5611
R1110 minus.n12 minus.n11 25.5611
R1111 minus.n43 minus.n42 25.5611
R1112 minus.n56 minus.n32 25.5611
R1113 minus.n27 minus.n26 21.1793
R1114 minus.n8 minus.n5 21.1793
R1115 minus.n39 minus.n36 21.1793
R1116 minus.n58 minus.n57 21.1793
R1117 minus.n29 minus.n28 16.7975
R1118 minus.n7 minus.n6 16.7975
R1119 minus.n38 minus.n37 16.7975
R1120 minus.n60 minus.n59 16.7975
R1121 minus.n62 minus.n61 6.48914
R1122 minus.n30 minus.n0 0.189894
R1123 minus.n24 minus.n0 0.189894
R1124 minus.n24 minus.n23 0.189894
R1125 minus.n23 minus.n2 0.189894
R1126 minus.n17 minus.n2 0.189894
R1127 minus.n17 minus.n16 0.189894
R1128 minus.n16 minus.n4 0.189894
R1129 minus.n10 minus.n4 0.189894
R1130 minus.n10 minus.n9 0.189894
R1131 minus.n41 minus.n40 0.189894
R1132 minus.n41 minus.n35 0.189894
R1133 minus.n47 minus.n35 0.189894
R1134 minus.n48 minus.n47 0.189894
R1135 minus.n48 minus.n33 0.189894
R1136 minus.n54 minus.n33 0.189894
R1137 minus.n55 minus.n54 0.189894
R1138 minus.n55 minus.n31 0.189894
R1139 minus.n61 minus.n31 0.189894
R1140 minus minus.n62 0.188
R1141 drain_right.n7 drain_right.n5 60.0094
R1142 drain_right.n2 drain_right.n0 60.0094
R1143 drain_right.n13 drain_right.n11 60.0094
R1144 drain_right.n13 drain_right.n12 59.5527
R1145 drain_right.n15 drain_right.n14 59.5527
R1146 drain_right.n17 drain_right.n16 59.5527
R1147 drain_right.n19 drain_right.n18 59.5527
R1148 drain_right.n21 drain_right.n20 59.5527
R1149 drain_right.n7 drain_right.n6 59.5525
R1150 drain_right.n9 drain_right.n8 59.5525
R1151 drain_right.n4 drain_right.n3 59.5525
R1152 drain_right.n2 drain_right.n1 59.5525
R1153 drain_right drain_right.n10 31.1544
R1154 drain_right drain_right.n21 6.11011
R1155 drain_right.n5 drain_right.t21 1.6505
R1156 drain_right.n5 drain_right.t17 1.6505
R1157 drain_right.n6 drain_right.t9 1.6505
R1158 drain_right.n6 drain_right.t16 1.6505
R1159 drain_right.n8 drain_right.t6 1.6505
R1160 drain_right.n8 drain_right.t13 1.6505
R1161 drain_right.n3 drain_right.t5 1.6505
R1162 drain_right.n3 drain_right.t12 1.6505
R1163 drain_right.n1 drain_right.t20 1.6505
R1164 drain_right.n1 drain_right.t15 1.6505
R1165 drain_right.n0 drain_right.t19 1.6505
R1166 drain_right.n0 drain_right.t14 1.6505
R1167 drain_right.n11 drain_right.t10 1.6505
R1168 drain_right.n11 drain_right.t3 1.6505
R1169 drain_right.n12 drain_right.t1 1.6505
R1170 drain_right.n12 drain_right.t23 1.6505
R1171 drain_right.n14 drain_right.t11 1.6505
R1172 drain_right.n14 drain_right.t2 1.6505
R1173 drain_right.n16 drain_right.t0 1.6505
R1174 drain_right.n16 drain_right.t22 1.6505
R1175 drain_right.n18 drain_right.t8 1.6505
R1176 drain_right.n18 drain_right.t4 1.6505
R1177 drain_right.n20 drain_right.t18 1.6505
R1178 drain_right.n20 drain_right.t7 1.6505
R1179 drain_right.n9 drain_right.n7 0.457397
R1180 drain_right.n4 drain_right.n2 0.457397
R1181 drain_right.n21 drain_right.n19 0.457397
R1182 drain_right.n19 drain_right.n17 0.457397
R1183 drain_right.n17 drain_right.n15 0.457397
R1184 drain_right.n15 drain_right.n13 0.457397
R1185 drain_right.n10 drain_right.n9 0.173602
R1186 drain_right.n10 drain_right.n4 0.173602
C0 drain_left source 53.724102f
C1 drain_left plus 6.424f
C2 source minus 5.89859f
C3 plus minus 5.76611f
C4 drain_right source 53.7244f
C5 drain_right plus 0.359911f
C6 drain_left minus 0.171754f
C7 drain_right drain_left 1.11966f
C8 plus source 5.91263f
C9 drain_right minus 6.21886f
C10 drain_right a_n2094_n3288# 7.48597f
C11 drain_left a_n2094_n3288# 7.81381f
C12 source a_n2094_n3288# 8.699999f
C13 minus a_n2094_n3288# 8.14979f
C14 plus a_n2094_n3288# 10.26675f
C15 drain_right.t19 a_n2094_n3288# 0.370641f
C16 drain_right.t14 a_n2094_n3288# 0.370641f
C17 drain_right.n0 a_n2094_n3288# 3.30163f
C18 drain_right.t20 a_n2094_n3288# 0.370641f
C19 drain_right.t15 a_n2094_n3288# 0.370641f
C20 drain_right.n1 a_n2094_n3288# 3.29814f
C21 drain_right.n2 a_n2094_n3288# 0.898481f
C22 drain_right.t5 a_n2094_n3288# 0.370641f
C23 drain_right.t12 a_n2094_n3288# 0.370641f
C24 drain_right.n3 a_n2094_n3288# 3.29814f
C25 drain_right.n4 a_n2094_n3288# 0.412609f
C26 drain_right.t21 a_n2094_n3288# 0.370641f
C27 drain_right.t17 a_n2094_n3288# 0.370641f
C28 drain_right.n5 a_n2094_n3288# 3.30163f
C29 drain_right.t9 a_n2094_n3288# 0.370641f
C30 drain_right.t16 a_n2094_n3288# 0.370641f
C31 drain_right.n6 a_n2094_n3288# 3.29814f
C32 drain_right.n7 a_n2094_n3288# 0.898481f
C33 drain_right.t6 a_n2094_n3288# 0.370641f
C34 drain_right.t13 a_n2094_n3288# 0.370641f
C35 drain_right.n8 a_n2094_n3288# 3.29814f
C36 drain_right.n9 a_n2094_n3288# 0.412609f
C37 drain_right.n10 a_n2094_n3288# 1.92398f
C38 drain_right.t10 a_n2094_n3288# 0.370641f
C39 drain_right.t3 a_n2094_n3288# 0.370641f
C40 drain_right.n11 a_n2094_n3288# 3.30163f
C41 drain_right.t1 a_n2094_n3288# 0.370641f
C42 drain_right.t23 a_n2094_n3288# 0.370641f
C43 drain_right.n12 a_n2094_n3288# 3.29815f
C44 drain_right.n13 a_n2094_n3288# 0.898467f
C45 drain_right.t11 a_n2094_n3288# 0.370641f
C46 drain_right.t2 a_n2094_n3288# 0.370641f
C47 drain_right.n14 a_n2094_n3288# 3.29815f
C48 drain_right.n15 a_n2094_n3288# 0.443102f
C49 drain_right.t0 a_n2094_n3288# 0.370641f
C50 drain_right.t22 a_n2094_n3288# 0.370641f
C51 drain_right.n16 a_n2094_n3288# 3.29815f
C52 drain_right.n17 a_n2094_n3288# 0.443102f
C53 drain_right.t8 a_n2094_n3288# 0.370641f
C54 drain_right.t4 a_n2094_n3288# 0.370641f
C55 drain_right.n18 a_n2094_n3288# 3.29815f
C56 drain_right.n19 a_n2094_n3288# 0.443102f
C57 drain_right.t18 a_n2094_n3288# 0.370641f
C58 drain_right.t7 a_n2094_n3288# 0.370641f
C59 drain_right.n20 a_n2094_n3288# 3.29815f
C60 drain_right.n21 a_n2094_n3288# 0.762983f
C61 minus.n0 a_n2094_n3288# 0.051639f
C62 minus.t5 a_n2094_n3288# 0.355606f
C63 minus.t16 a_n2094_n3288# 0.350216f
C64 minus.t15 a_n2094_n3288# 0.350216f
C65 minus.t19 a_n2094_n3288# 0.350216f
C66 minus.n1 a_n2094_n3288# 0.144235f
C67 minus.n2 a_n2094_n3288# 0.051639f
C68 minus.t23 a_n2094_n3288# 0.350216f
C69 minus.t1 a_n2094_n3288# 0.350216f
C70 minus.t12 a_n2094_n3288# 0.350216f
C71 minus.n3 a_n2094_n3288# 0.144235f
C72 minus.n4 a_n2094_n3288# 0.051639f
C73 minus.t21 a_n2094_n3288# 0.350216f
C74 minus.t22 a_n2094_n3288# 0.350216f
C75 minus.t0 a_n2094_n3288# 0.350216f
C76 minus.n5 a_n2094_n3288# 0.144235f
C77 minus.t20 a_n2094_n3288# 0.355606f
C78 minus.n6 a_n2094_n3288# 0.160672f
C79 minus.t13 a_n2094_n3288# 0.350216f
C80 minus.n7 a_n2094_n3288# 0.144235f
C81 minus.n8 a_n2094_n3288# 0.018086f
C82 minus.n9 a_n2094_n3288# 0.120072f
C83 minus.n10 a_n2094_n3288# 0.051639f
C84 minus.n11 a_n2094_n3288# 0.018086f
C85 minus.n12 a_n2094_n3288# 0.144235f
C86 minus.n13 a_n2094_n3288# 0.018086f
C87 minus.n14 a_n2094_n3288# 0.144235f
C88 minus.n15 a_n2094_n3288# 0.018086f
C89 minus.n16 a_n2094_n3288# 0.051639f
C90 minus.n17 a_n2094_n3288# 0.051639f
C91 minus.n18 a_n2094_n3288# 0.018086f
C92 minus.n19 a_n2094_n3288# 0.144235f
C93 minus.n20 a_n2094_n3288# 0.018086f
C94 minus.n21 a_n2094_n3288# 0.144235f
C95 minus.n22 a_n2094_n3288# 0.018086f
C96 minus.n23 a_n2094_n3288# 0.051639f
C97 minus.n24 a_n2094_n3288# 0.051639f
C98 minus.n25 a_n2094_n3288# 0.018086f
C99 minus.n26 a_n2094_n3288# 0.144235f
C100 minus.n27 a_n2094_n3288# 0.018086f
C101 minus.n28 a_n2094_n3288# 0.144235f
C102 minus.n29 a_n2094_n3288# 0.160592f
C103 minus.n30 a_n2094_n3288# 1.89155f
C104 minus.n31 a_n2094_n3288# 0.051639f
C105 minus.t2 a_n2094_n3288# 0.350216f
C106 minus.t7 a_n2094_n3288# 0.350216f
C107 minus.t14 a_n2094_n3288# 0.350216f
C108 minus.n32 a_n2094_n3288# 0.144235f
C109 minus.n33 a_n2094_n3288# 0.051639f
C110 minus.t10 a_n2094_n3288# 0.350216f
C111 minus.t17 a_n2094_n3288# 0.350216f
C112 minus.t11 a_n2094_n3288# 0.350216f
C113 minus.n34 a_n2094_n3288# 0.144235f
C114 minus.n35 a_n2094_n3288# 0.051639f
C115 minus.t18 a_n2094_n3288# 0.350216f
C116 minus.t8 a_n2094_n3288# 0.350216f
C117 minus.t3 a_n2094_n3288# 0.350216f
C118 minus.n36 a_n2094_n3288# 0.144235f
C119 minus.t4 a_n2094_n3288# 0.355606f
C120 minus.n37 a_n2094_n3288# 0.160672f
C121 minus.t9 a_n2094_n3288# 0.350216f
C122 minus.n38 a_n2094_n3288# 0.144235f
C123 minus.n39 a_n2094_n3288# 0.018086f
C124 minus.n40 a_n2094_n3288# 0.120072f
C125 minus.n41 a_n2094_n3288# 0.051639f
C126 minus.n42 a_n2094_n3288# 0.018086f
C127 minus.n43 a_n2094_n3288# 0.144235f
C128 minus.n44 a_n2094_n3288# 0.018086f
C129 minus.n45 a_n2094_n3288# 0.144235f
C130 minus.n46 a_n2094_n3288# 0.018086f
C131 minus.n47 a_n2094_n3288# 0.051639f
C132 minus.n48 a_n2094_n3288# 0.051639f
C133 minus.n49 a_n2094_n3288# 0.018086f
C134 minus.n50 a_n2094_n3288# 0.144235f
C135 minus.n51 a_n2094_n3288# 0.018086f
C136 minus.n52 a_n2094_n3288# 0.144235f
C137 minus.n53 a_n2094_n3288# 0.018086f
C138 minus.n54 a_n2094_n3288# 0.051639f
C139 minus.n55 a_n2094_n3288# 0.051639f
C140 minus.n56 a_n2094_n3288# 0.018086f
C141 minus.n57 a_n2094_n3288# 0.144235f
C142 minus.n58 a_n2094_n3288# 0.018086f
C143 minus.n59 a_n2094_n3288# 0.144235f
C144 minus.t6 a_n2094_n3288# 0.355606f
C145 minus.n60 a_n2094_n3288# 0.160592f
C146 minus.n61 a_n2094_n3288# 0.336282f
C147 minus.n62 a_n2094_n3288# 2.29238f
C148 source.n0 a_n2094_n3288# 0.045931f
C149 source.n1 a_n2094_n3288# 0.034675f
C150 source.n2 a_n2094_n3288# 0.018633f
C151 source.n3 a_n2094_n3288# 0.044041f
C152 source.n4 a_n2094_n3288# 0.019729f
C153 source.n5 a_n2094_n3288# 0.034675f
C154 source.n6 a_n2094_n3288# 0.018633f
C155 source.n7 a_n2094_n3288# 0.044041f
C156 source.n8 a_n2094_n3288# 0.019729f
C157 source.n9 a_n2094_n3288# 0.034675f
C158 source.n10 a_n2094_n3288# 0.019181f
C159 source.n11 a_n2094_n3288# 0.044041f
C160 source.n12 a_n2094_n3288# 0.018633f
C161 source.n13 a_n2094_n3288# 0.019729f
C162 source.n14 a_n2094_n3288# 0.034675f
C163 source.n15 a_n2094_n3288# 0.018633f
C164 source.n16 a_n2094_n3288# 0.044041f
C165 source.n17 a_n2094_n3288# 0.019729f
C166 source.n18 a_n2094_n3288# 0.034675f
C167 source.n19 a_n2094_n3288# 0.018633f
C168 source.n20 a_n2094_n3288# 0.033031f
C169 source.n21 a_n2094_n3288# 0.031133f
C170 source.t10 a_n2094_n3288# 0.074382f
C171 source.n22 a_n2094_n3288# 0.25f
C172 source.n23 a_n2094_n3288# 1.74928f
C173 source.n24 a_n2094_n3288# 0.018633f
C174 source.n25 a_n2094_n3288# 0.019729f
C175 source.n26 a_n2094_n3288# 0.044041f
C176 source.n27 a_n2094_n3288# 0.044041f
C177 source.n28 a_n2094_n3288# 0.019729f
C178 source.n29 a_n2094_n3288# 0.018633f
C179 source.n30 a_n2094_n3288# 0.034675f
C180 source.n31 a_n2094_n3288# 0.034675f
C181 source.n32 a_n2094_n3288# 0.018633f
C182 source.n33 a_n2094_n3288# 0.019729f
C183 source.n34 a_n2094_n3288# 0.044041f
C184 source.n35 a_n2094_n3288# 0.044041f
C185 source.n36 a_n2094_n3288# 0.019729f
C186 source.n37 a_n2094_n3288# 0.018633f
C187 source.n38 a_n2094_n3288# 0.034675f
C188 source.n39 a_n2094_n3288# 0.034675f
C189 source.n40 a_n2094_n3288# 0.018633f
C190 source.n41 a_n2094_n3288# 0.019729f
C191 source.n42 a_n2094_n3288# 0.044041f
C192 source.n43 a_n2094_n3288# 0.044041f
C193 source.n44 a_n2094_n3288# 0.044041f
C194 source.n45 a_n2094_n3288# 0.019181f
C195 source.n46 a_n2094_n3288# 0.018633f
C196 source.n47 a_n2094_n3288# 0.034675f
C197 source.n48 a_n2094_n3288# 0.034675f
C198 source.n49 a_n2094_n3288# 0.018633f
C199 source.n50 a_n2094_n3288# 0.019729f
C200 source.n51 a_n2094_n3288# 0.044041f
C201 source.n52 a_n2094_n3288# 0.044041f
C202 source.n53 a_n2094_n3288# 0.019729f
C203 source.n54 a_n2094_n3288# 0.018633f
C204 source.n55 a_n2094_n3288# 0.034675f
C205 source.n56 a_n2094_n3288# 0.034675f
C206 source.n57 a_n2094_n3288# 0.018633f
C207 source.n58 a_n2094_n3288# 0.019729f
C208 source.n59 a_n2094_n3288# 0.044041f
C209 source.n60 a_n2094_n3288# 0.090376f
C210 source.n61 a_n2094_n3288# 0.019729f
C211 source.n62 a_n2094_n3288# 0.018633f
C212 source.n63 a_n2094_n3288# 0.074464f
C213 source.n64 a_n2094_n3288# 0.049878f
C214 source.n65 a_n2094_n3288# 1.37967f
C215 source.t27 a_n2094_n3288# 0.328811f
C216 source.t30 a_n2094_n3288# 0.328811f
C217 source.n66 a_n2094_n3288# 2.81529f
C218 source.n67 a_n2094_n3288# 0.456601f
C219 source.t9 a_n2094_n3288# 0.328811f
C220 source.t19 a_n2094_n3288# 0.328811f
C221 source.n68 a_n2094_n3288# 2.81529f
C222 source.n69 a_n2094_n3288# 0.456601f
C223 source.t25 a_n2094_n3288# 0.328811f
C224 source.t29 a_n2094_n3288# 0.328811f
C225 source.n70 a_n2094_n3288# 2.81529f
C226 source.n71 a_n2094_n3288# 0.456601f
C227 source.t16 a_n2094_n3288# 0.328811f
C228 source.t17 a_n2094_n3288# 0.328811f
C229 source.n72 a_n2094_n3288# 2.81529f
C230 source.n73 a_n2094_n3288# 0.456601f
C231 source.t28 a_n2094_n3288# 0.328811f
C232 source.t8 a_n2094_n3288# 0.328811f
C233 source.n74 a_n2094_n3288# 2.81529f
C234 source.n75 a_n2094_n3288# 0.456601f
C235 source.n76 a_n2094_n3288# 0.045931f
C236 source.n77 a_n2094_n3288# 0.034675f
C237 source.n78 a_n2094_n3288# 0.018633f
C238 source.n79 a_n2094_n3288# 0.044041f
C239 source.n80 a_n2094_n3288# 0.019729f
C240 source.n81 a_n2094_n3288# 0.034675f
C241 source.n82 a_n2094_n3288# 0.018633f
C242 source.n83 a_n2094_n3288# 0.044041f
C243 source.n84 a_n2094_n3288# 0.019729f
C244 source.n85 a_n2094_n3288# 0.034675f
C245 source.n86 a_n2094_n3288# 0.019181f
C246 source.n87 a_n2094_n3288# 0.044041f
C247 source.n88 a_n2094_n3288# 0.018633f
C248 source.n89 a_n2094_n3288# 0.019729f
C249 source.n90 a_n2094_n3288# 0.034675f
C250 source.n91 a_n2094_n3288# 0.018633f
C251 source.n92 a_n2094_n3288# 0.044041f
C252 source.n93 a_n2094_n3288# 0.019729f
C253 source.n94 a_n2094_n3288# 0.034675f
C254 source.n95 a_n2094_n3288# 0.018633f
C255 source.n96 a_n2094_n3288# 0.033031f
C256 source.n97 a_n2094_n3288# 0.031133f
C257 source.t24 a_n2094_n3288# 0.074382f
C258 source.n98 a_n2094_n3288# 0.25f
C259 source.n99 a_n2094_n3288# 1.74928f
C260 source.n100 a_n2094_n3288# 0.018633f
C261 source.n101 a_n2094_n3288# 0.019729f
C262 source.n102 a_n2094_n3288# 0.044041f
C263 source.n103 a_n2094_n3288# 0.044041f
C264 source.n104 a_n2094_n3288# 0.019729f
C265 source.n105 a_n2094_n3288# 0.018633f
C266 source.n106 a_n2094_n3288# 0.034675f
C267 source.n107 a_n2094_n3288# 0.034675f
C268 source.n108 a_n2094_n3288# 0.018633f
C269 source.n109 a_n2094_n3288# 0.019729f
C270 source.n110 a_n2094_n3288# 0.044041f
C271 source.n111 a_n2094_n3288# 0.044041f
C272 source.n112 a_n2094_n3288# 0.019729f
C273 source.n113 a_n2094_n3288# 0.018633f
C274 source.n114 a_n2094_n3288# 0.034675f
C275 source.n115 a_n2094_n3288# 0.034675f
C276 source.n116 a_n2094_n3288# 0.018633f
C277 source.n117 a_n2094_n3288# 0.019729f
C278 source.n118 a_n2094_n3288# 0.044041f
C279 source.n119 a_n2094_n3288# 0.044041f
C280 source.n120 a_n2094_n3288# 0.044041f
C281 source.n121 a_n2094_n3288# 0.019181f
C282 source.n122 a_n2094_n3288# 0.018633f
C283 source.n123 a_n2094_n3288# 0.034675f
C284 source.n124 a_n2094_n3288# 0.034675f
C285 source.n125 a_n2094_n3288# 0.018633f
C286 source.n126 a_n2094_n3288# 0.019729f
C287 source.n127 a_n2094_n3288# 0.044041f
C288 source.n128 a_n2094_n3288# 0.044041f
C289 source.n129 a_n2094_n3288# 0.019729f
C290 source.n130 a_n2094_n3288# 0.018633f
C291 source.n131 a_n2094_n3288# 0.034675f
C292 source.n132 a_n2094_n3288# 0.034675f
C293 source.n133 a_n2094_n3288# 0.018633f
C294 source.n134 a_n2094_n3288# 0.019729f
C295 source.n135 a_n2094_n3288# 0.044041f
C296 source.n136 a_n2094_n3288# 0.090376f
C297 source.n137 a_n2094_n3288# 0.019729f
C298 source.n138 a_n2094_n3288# 0.018633f
C299 source.n139 a_n2094_n3288# 0.074464f
C300 source.n140 a_n2094_n3288# 0.049878f
C301 source.n141 a_n2094_n3288# 0.129955f
C302 source.n142 a_n2094_n3288# 0.045931f
C303 source.n143 a_n2094_n3288# 0.034675f
C304 source.n144 a_n2094_n3288# 0.018633f
C305 source.n145 a_n2094_n3288# 0.044041f
C306 source.n146 a_n2094_n3288# 0.019729f
C307 source.n147 a_n2094_n3288# 0.034675f
C308 source.n148 a_n2094_n3288# 0.018633f
C309 source.n149 a_n2094_n3288# 0.044041f
C310 source.n150 a_n2094_n3288# 0.019729f
C311 source.n151 a_n2094_n3288# 0.034675f
C312 source.n152 a_n2094_n3288# 0.019181f
C313 source.n153 a_n2094_n3288# 0.044041f
C314 source.n154 a_n2094_n3288# 0.018633f
C315 source.n155 a_n2094_n3288# 0.019729f
C316 source.n156 a_n2094_n3288# 0.034675f
C317 source.n157 a_n2094_n3288# 0.018633f
C318 source.n158 a_n2094_n3288# 0.044041f
C319 source.n159 a_n2094_n3288# 0.019729f
C320 source.n160 a_n2094_n3288# 0.034675f
C321 source.n161 a_n2094_n3288# 0.018633f
C322 source.n162 a_n2094_n3288# 0.033031f
C323 source.n163 a_n2094_n3288# 0.031133f
C324 source.t2 a_n2094_n3288# 0.074382f
C325 source.n164 a_n2094_n3288# 0.25f
C326 source.n165 a_n2094_n3288# 1.74928f
C327 source.n166 a_n2094_n3288# 0.018633f
C328 source.n167 a_n2094_n3288# 0.019729f
C329 source.n168 a_n2094_n3288# 0.044041f
C330 source.n169 a_n2094_n3288# 0.044041f
C331 source.n170 a_n2094_n3288# 0.019729f
C332 source.n171 a_n2094_n3288# 0.018633f
C333 source.n172 a_n2094_n3288# 0.034675f
C334 source.n173 a_n2094_n3288# 0.034675f
C335 source.n174 a_n2094_n3288# 0.018633f
C336 source.n175 a_n2094_n3288# 0.019729f
C337 source.n176 a_n2094_n3288# 0.044041f
C338 source.n177 a_n2094_n3288# 0.044041f
C339 source.n178 a_n2094_n3288# 0.019729f
C340 source.n179 a_n2094_n3288# 0.018633f
C341 source.n180 a_n2094_n3288# 0.034675f
C342 source.n181 a_n2094_n3288# 0.034675f
C343 source.n182 a_n2094_n3288# 0.018633f
C344 source.n183 a_n2094_n3288# 0.019729f
C345 source.n184 a_n2094_n3288# 0.044041f
C346 source.n185 a_n2094_n3288# 0.044041f
C347 source.n186 a_n2094_n3288# 0.044041f
C348 source.n187 a_n2094_n3288# 0.019181f
C349 source.n188 a_n2094_n3288# 0.018633f
C350 source.n189 a_n2094_n3288# 0.034675f
C351 source.n190 a_n2094_n3288# 0.034675f
C352 source.n191 a_n2094_n3288# 0.018633f
C353 source.n192 a_n2094_n3288# 0.019729f
C354 source.n193 a_n2094_n3288# 0.044041f
C355 source.n194 a_n2094_n3288# 0.044041f
C356 source.n195 a_n2094_n3288# 0.019729f
C357 source.n196 a_n2094_n3288# 0.018633f
C358 source.n197 a_n2094_n3288# 0.034675f
C359 source.n198 a_n2094_n3288# 0.034675f
C360 source.n199 a_n2094_n3288# 0.018633f
C361 source.n200 a_n2094_n3288# 0.019729f
C362 source.n201 a_n2094_n3288# 0.044041f
C363 source.n202 a_n2094_n3288# 0.090376f
C364 source.n203 a_n2094_n3288# 0.019729f
C365 source.n204 a_n2094_n3288# 0.018633f
C366 source.n205 a_n2094_n3288# 0.074464f
C367 source.n206 a_n2094_n3288# 0.049878f
C368 source.n207 a_n2094_n3288# 0.129955f
C369 source.t40 a_n2094_n3288# 0.328811f
C370 source.t3 a_n2094_n3288# 0.328811f
C371 source.n208 a_n2094_n3288# 2.81529f
C372 source.n209 a_n2094_n3288# 0.456601f
C373 source.t44 a_n2094_n3288# 0.328811f
C374 source.t34 a_n2094_n3288# 0.328811f
C375 source.n210 a_n2094_n3288# 2.81529f
C376 source.n211 a_n2094_n3288# 0.456601f
C377 source.t46 a_n2094_n3288# 0.328811f
C378 source.t31 a_n2094_n3288# 0.328811f
C379 source.n212 a_n2094_n3288# 2.81529f
C380 source.n213 a_n2094_n3288# 0.456601f
C381 source.t37 a_n2094_n3288# 0.328811f
C382 source.t39 a_n2094_n3288# 0.328811f
C383 source.n214 a_n2094_n3288# 2.81529f
C384 source.n215 a_n2094_n3288# 0.456601f
C385 source.t6 a_n2094_n3288# 0.328811f
C386 source.t38 a_n2094_n3288# 0.328811f
C387 source.n216 a_n2094_n3288# 2.81529f
C388 source.n217 a_n2094_n3288# 0.456601f
C389 source.n218 a_n2094_n3288# 0.045931f
C390 source.n219 a_n2094_n3288# 0.034675f
C391 source.n220 a_n2094_n3288# 0.018633f
C392 source.n221 a_n2094_n3288# 0.044041f
C393 source.n222 a_n2094_n3288# 0.019729f
C394 source.n223 a_n2094_n3288# 0.034675f
C395 source.n224 a_n2094_n3288# 0.018633f
C396 source.n225 a_n2094_n3288# 0.044041f
C397 source.n226 a_n2094_n3288# 0.019729f
C398 source.n227 a_n2094_n3288# 0.034675f
C399 source.n228 a_n2094_n3288# 0.019181f
C400 source.n229 a_n2094_n3288# 0.044041f
C401 source.n230 a_n2094_n3288# 0.018633f
C402 source.n231 a_n2094_n3288# 0.019729f
C403 source.n232 a_n2094_n3288# 0.034675f
C404 source.n233 a_n2094_n3288# 0.018633f
C405 source.n234 a_n2094_n3288# 0.044041f
C406 source.n235 a_n2094_n3288# 0.019729f
C407 source.n236 a_n2094_n3288# 0.034675f
C408 source.n237 a_n2094_n3288# 0.018633f
C409 source.n238 a_n2094_n3288# 0.033031f
C410 source.n239 a_n2094_n3288# 0.031133f
C411 source.t35 a_n2094_n3288# 0.074382f
C412 source.n240 a_n2094_n3288# 0.25f
C413 source.n241 a_n2094_n3288# 1.74928f
C414 source.n242 a_n2094_n3288# 0.018633f
C415 source.n243 a_n2094_n3288# 0.019729f
C416 source.n244 a_n2094_n3288# 0.044041f
C417 source.n245 a_n2094_n3288# 0.044041f
C418 source.n246 a_n2094_n3288# 0.019729f
C419 source.n247 a_n2094_n3288# 0.018633f
C420 source.n248 a_n2094_n3288# 0.034675f
C421 source.n249 a_n2094_n3288# 0.034675f
C422 source.n250 a_n2094_n3288# 0.018633f
C423 source.n251 a_n2094_n3288# 0.019729f
C424 source.n252 a_n2094_n3288# 0.044041f
C425 source.n253 a_n2094_n3288# 0.044041f
C426 source.n254 a_n2094_n3288# 0.019729f
C427 source.n255 a_n2094_n3288# 0.018633f
C428 source.n256 a_n2094_n3288# 0.034675f
C429 source.n257 a_n2094_n3288# 0.034675f
C430 source.n258 a_n2094_n3288# 0.018633f
C431 source.n259 a_n2094_n3288# 0.019729f
C432 source.n260 a_n2094_n3288# 0.044041f
C433 source.n261 a_n2094_n3288# 0.044041f
C434 source.n262 a_n2094_n3288# 0.044041f
C435 source.n263 a_n2094_n3288# 0.019181f
C436 source.n264 a_n2094_n3288# 0.018633f
C437 source.n265 a_n2094_n3288# 0.034675f
C438 source.n266 a_n2094_n3288# 0.034675f
C439 source.n267 a_n2094_n3288# 0.018633f
C440 source.n268 a_n2094_n3288# 0.019729f
C441 source.n269 a_n2094_n3288# 0.044041f
C442 source.n270 a_n2094_n3288# 0.044041f
C443 source.n271 a_n2094_n3288# 0.019729f
C444 source.n272 a_n2094_n3288# 0.018633f
C445 source.n273 a_n2094_n3288# 0.034675f
C446 source.n274 a_n2094_n3288# 0.034675f
C447 source.n275 a_n2094_n3288# 0.018633f
C448 source.n276 a_n2094_n3288# 0.019729f
C449 source.n277 a_n2094_n3288# 0.044041f
C450 source.n278 a_n2094_n3288# 0.090376f
C451 source.n279 a_n2094_n3288# 0.019729f
C452 source.n280 a_n2094_n3288# 0.018633f
C453 source.n281 a_n2094_n3288# 0.074464f
C454 source.n282 a_n2094_n3288# 0.049878f
C455 source.n283 a_n2094_n3288# 1.92145f
C456 source.n284 a_n2094_n3288# 0.045931f
C457 source.n285 a_n2094_n3288# 0.034675f
C458 source.n286 a_n2094_n3288# 0.018633f
C459 source.n287 a_n2094_n3288# 0.044041f
C460 source.n288 a_n2094_n3288# 0.019729f
C461 source.n289 a_n2094_n3288# 0.034675f
C462 source.n290 a_n2094_n3288# 0.018633f
C463 source.n291 a_n2094_n3288# 0.044041f
C464 source.n292 a_n2094_n3288# 0.019729f
C465 source.n293 a_n2094_n3288# 0.034675f
C466 source.n294 a_n2094_n3288# 0.019181f
C467 source.n295 a_n2094_n3288# 0.044041f
C468 source.n296 a_n2094_n3288# 0.019729f
C469 source.n297 a_n2094_n3288# 0.034675f
C470 source.n298 a_n2094_n3288# 0.018633f
C471 source.n299 a_n2094_n3288# 0.044041f
C472 source.n300 a_n2094_n3288# 0.019729f
C473 source.n301 a_n2094_n3288# 0.034675f
C474 source.n302 a_n2094_n3288# 0.018633f
C475 source.n303 a_n2094_n3288# 0.033031f
C476 source.n304 a_n2094_n3288# 0.031133f
C477 source.t15 a_n2094_n3288# 0.074382f
C478 source.n305 a_n2094_n3288# 0.25f
C479 source.n306 a_n2094_n3288# 1.74928f
C480 source.n307 a_n2094_n3288# 0.018633f
C481 source.n308 a_n2094_n3288# 0.019729f
C482 source.n309 a_n2094_n3288# 0.044041f
C483 source.n310 a_n2094_n3288# 0.044041f
C484 source.n311 a_n2094_n3288# 0.019729f
C485 source.n312 a_n2094_n3288# 0.018633f
C486 source.n313 a_n2094_n3288# 0.034675f
C487 source.n314 a_n2094_n3288# 0.034675f
C488 source.n315 a_n2094_n3288# 0.018633f
C489 source.n316 a_n2094_n3288# 0.019729f
C490 source.n317 a_n2094_n3288# 0.044041f
C491 source.n318 a_n2094_n3288# 0.044041f
C492 source.n319 a_n2094_n3288# 0.019729f
C493 source.n320 a_n2094_n3288# 0.018633f
C494 source.n321 a_n2094_n3288# 0.034675f
C495 source.n322 a_n2094_n3288# 0.034675f
C496 source.n323 a_n2094_n3288# 0.018633f
C497 source.n324 a_n2094_n3288# 0.018633f
C498 source.n325 a_n2094_n3288# 0.019729f
C499 source.n326 a_n2094_n3288# 0.044041f
C500 source.n327 a_n2094_n3288# 0.044041f
C501 source.n328 a_n2094_n3288# 0.044041f
C502 source.n329 a_n2094_n3288# 0.019181f
C503 source.n330 a_n2094_n3288# 0.018633f
C504 source.n331 a_n2094_n3288# 0.034675f
C505 source.n332 a_n2094_n3288# 0.034675f
C506 source.n333 a_n2094_n3288# 0.018633f
C507 source.n334 a_n2094_n3288# 0.019729f
C508 source.n335 a_n2094_n3288# 0.044041f
C509 source.n336 a_n2094_n3288# 0.044041f
C510 source.n337 a_n2094_n3288# 0.019729f
C511 source.n338 a_n2094_n3288# 0.018633f
C512 source.n339 a_n2094_n3288# 0.034675f
C513 source.n340 a_n2094_n3288# 0.034675f
C514 source.n341 a_n2094_n3288# 0.018633f
C515 source.n342 a_n2094_n3288# 0.019729f
C516 source.n343 a_n2094_n3288# 0.044041f
C517 source.n344 a_n2094_n3288# 0.090376f
C518 source.n345 a_n2094_n3288# 0.019729f
C519 source.n346 a_n2094_n3288# 0.018633f
C520 source.n347 a_n2094_n3288# 0.074464f
C521 source.n348 a_n2094_n3288# 0.049878f
C522 source.n349 a_n2094_n3288# 1.92145f
C523 source.t22 a_n2094_n3288# 0.328811f
C524 source.t26 a_n2094_n3288# 0.328811f
C525 source.n350 a_n2094_n3288# 2.81527f
C526 source.n351 a_n2094_n3288# 0.456618f
C527 source.t23 a_n2094_n3288# 0.328811f
C528 source.t20 a_n2094_n3288# 0.328811f
C529 source.n352 a_n2094_n3288# 2.81527f
C530 source.n353 a_n2094_n3288# 0.456618f
C531 source.t14 a_n2094_n3288# 0.328811f
C532 source.t21 a_n2094_n3288# 0.328811f
C533 source.n354 a_n2094_n3288# 2.81527f
C534 source.n355 a_n2094_n3288# 0.456618f
C535 source.t12 a_n2094_n3288# 0.328811f
C536 source.t18 a_n2094_n3288# 0.328811f
C537 source.n356 a_n2094_n3288# 2.81527f
C538 source.n357 a_n2094_n3288# 0.456618f
C539 source.t13 a_n2094_n3288# 0.328811f
C540 source.t7 a_n2094_n3288# 0.328811f
C541 source.n358 a_n2094_n3288# 2.81527f
C542 source.n359 a_n2094_n3288# 0.456618f
C543 source.n360 a_n2094_n3288# 0.045931f
C544 source.n361 a_n2094_n3288# 0.034675f
C545 source.n362 a_n2094_n3288# 0.018633f
C546 source.n363 a_n2094_n3288# 0.044041f
C547 source.n364 a_n2094_n3288# 0.019729f
C548 source.n365 a_n2094_n3288# 0.034675f
C549 source.n366 a_n2094_n3288# 0.018633f
C550 source.n367 a_n2094_n3288# 0.044041f
C551 source.n368 a_n2094_n3288# 0.019729f
C552 source.n369 a_n2094_n3288# 0.034675f
C553 source.n370 a_n2094_n3288# 0.019181f
C554 source.n371 a_n2094_n3288# 0.044041f
C555 source.n372 a_n2094_n3288# 0.019729f
C556 source.n373 a_n2094_n3288# 0.034675f
C557 source.n374 a_n2094_n3288# 0.018633f
C558 source.n375 a_n2094_n3288# 0.044041f
C559 source.n376 a_n2094_n3288# 0.019729f
C560 source.n377 a_n2094_n3288# 0.034675f
C561 source.n378 a_n2094_n3288# 0.018633f
C562 source.n379 a_n2094_n3288# 0.033031f
C563 source.n380 a_n2094_n3288# 0.031133f
C564 source.t11 a_n2094_n3288# 0.074382f
C565 source.n381 a_n2094_n3288# 0.25f
C566 source.n382 a_n2094_n3288# 1.74928f
C567 source.n383 a_n2094_n3288# 0.018633f
C568 source.n384 a_n2094_n3288# 0.019729f
C569 source.n385 a_n2094_n3288# 0.044041f
C570 source.n386 a_n2094_n3288# 0.044041f
C571 source.n387 a_n2094_n3288# 0.019729f
C572 source.n388 a_n2094_n3288# 0.018633f
C573 source.n389 a_n2094_n3288# 0.034675f
C574 source.n390 a_n2094_n3288# 0.034675f
C575 source.n391 a_n2094_n3288# 0.018633f
C576 source.n392 a_n2094_n3288# 0.019729f
C577 source.n393 a_n2094_n3288# 0.044041f
C578 source.n394 a_n2094_n3288# 0.044041f
C579 source.n395 a_n2094_n3288# 0.019729f
C580 source.n396 a_n2094_n3288# 0.018633f
C581 source.n397 a_n2094_n3288# 0.034675f
C582 source.n398 a_n2094_n3288# 0.034675f
C583 source.n399 a_n2094_n3288# 0.018633f
C584 source.n400 a_n2094_n3288# 0.018633f
C585 source.n401 a_n2094_n3288# 0.019729f
C586 source.n402 a_n2094_n3288# 0.044041f
C587 source.n403 a_n2094_n3288# 0.044041f
C588 source.n404 a_n2094_n3288# 0.044041f
C589 source.n405 a_n2094_n3288# 0.019181f
C590 source.n406 a_n2094_n3288# 0.018633f
C591 source.n407 a_n2094_n3288# 0.034675f
C592 source.n408 a_n2094_n3288# 0.034675f
C593 source.n409 a_n2094_n3288# 0.018633f
C594 source.n410 a_n2094_n3288# 0.019729f
C595 source.n411 a_n2094_n3288# 0.044041f
C596 source.n412 a_n2094_n3288# 0.044041f
C597 source.n413 a_n2094_n3288# 0.019729f
C598 source.n414 a_n2094_n3288# 0.018633f
C599 source.n415 a_n2094_n3288# 0.034675f
C600 source.n416 a_n2094_n3288# 0.034675f
C601 source.n417 a_n2094_n3288# 0.018633f
C602 source.n418 a_n2094_n3288# 0.019729f
C603 source.n419 a_n2094_n3288# 0.044041f
C604 source.n420 a_n2094_n3288# 0.090376f
C605 source.n421 a_n2094_n3288# 0.019729f
C606 source.n422 a_n2094_n3288# 0.018633f
C607 source.n423 a_n2094_n3288# 0.074464f
C608 source.n424 a_n2094_n3288# 0.049878f
C609 source.n425 a_n2094_n3288# 0.129955f
C610 source.n426 a_n2094_n3288# 0.045931f
C611 source.n427 a_n2094_n3288# 0.034675f
C612 source.n428 a_n2094_n3288# 0.018633f
C613 source.n429 a_n2094_n3288# 0.044041f
C614 source.n430 a_n2094_n3288# 0.019729f
C615 source.n431 a_n2094_n3288# 0.034675f
C616 source.n432 a_n2094_n3288# 0.018633f
C617 source.n433 a_n2094_n3288# 0.044041f
C618 source.n434 a_n2094_n3288# 0.019729f
C619 source.n435 a_n2094_n3288# 0.034675f
C620 source.n436 a_n2094_n3288# 0.019181f
C621 source.n437 a_n2094_n3288# 0.044041f
C622 source.n438 a_n2094_n3288# 0.019729f
C623 source.n439 a_n2094_n3288# 0.034675f
C624 source.n440 a_n2094_n3288# 0.018633f
C625 source.n441 a_n2094_n3288# 0.044041f
C626 source.n442 a_n2094_n3288# 0.019729f
C627 source.n443 a_n2094_n3288# 0.034675f
C628 source.n444 a_n2094_n3288# 0.018633f
C629 source.n445 a_n2094_n3288# 0.033031f
C630 source.n446 a_n2094_n3288# 0.031133f
C631 source.t41 a_n2094_n3288# 0.074382f
C632 source.n447 a_n2094_n3288# 0.25f
C633 source.n448 a_n2094_n3288# 1.74928f
C634 source.n449 a_n2094_n3288# 0.018633f
C635 source.n450 a_n2094_n3288# 0.019729f
C636 source.n451 a_n2094_n3288# 0.044041f
C637 source.n452 a_n2094_n3288# 0.044041f
C638 source.n453 a_n2094_n3288# 0.019729f
C639 source.n454 a_n2094_n3288# 0.018633f
C640 source.n455 a_n2094_n3288# 0.034675f
C641 source.n456 a_n2094_n3288# 0.034675f
C642 source.n457 a_n2094_n3288# 0.018633f
C643 source.n458 a_n2094_n3288# 0.019729f
C644 source.n459 a_n2094_n3288# 0.044041f
C645 source.n460 a_n2094_n3288# 0.044041f
C646 source.n461 a_n2094_n3288# 0.019729f
C647 source.n462 a_n2094_n3288# 0.018633f
C648 source.n463 a_n2094_n3288# 0.034675f
C649 source.n464 a_n2094_n3288# 0.034675f
C650 source.n465 a_n2094_n3288# 0.018633f
C651 source.n466 a_n2094_n3288# 0.018633f
C652 source.n467 a_n2094_n3288# 0.019729f
C653 source.n468 a_n2094_n3288# 0.044041f
C654 source.n469 a_n2094_n3288# 0.044041f
C655 source.n470 a_n2094_n3288# 0.044041f
C656 source.n471 a_n2094_n3288# 0.019181f
C657 source.n472 a_n2094_n3288# 0.018633f
C658 source.n473 a_n2094_n3288# 0.034675f
C659 source.n474 a_n2094_n3288# 0.034675f
C660 source.n475 a_n2094_n3288# 0.018633f
C661 source.n476 a_n2094_n3288# 0.019729f
C662 source.n477 a_n2094_n3288# 0.044041f
C663 source.n478 a_n2094_n3288# 0.044041f
C664 source.n479 a_n2094_n3288# 0.019729f
C665 source.n480 a_n2094_n3288# 0.018633f
C666 source.n481 a_n2094_n3288# 0.034675f
C667 source.n482 a_n2094_n3288# 0.034675f
C668 source.n483 a_n2094_n3288# 0.018633f
C669 source.n484 a_n2094_n3288# 0.019729f
C670 source.n485 a_n2094_n3288# 0.044041f
C671 source.n486 a_n2094_n3288# 0.090376f
C672 source.n487 a_n2094_n3288# 0.019729f
C673 source.n488 a_n2094_n3288# 0.018633f
C674 source.n489 a_n2094_n3288# 0.074464f
C675 source.n490 a_n2094_n3288# 0.049878f
C676 source.n491 a_n2094_n3288# 0.129955f
C677 source.t0 a_n2094_n3288# 0.328811f
C678 source.t42 a_n2094_n3288# 0.328811f
C679 source.n492 a_n2094_n3288# 2.81527f
C680 source.n493 a_n2094_n3288# 0.456618f
C681 source.t36 a_n2094_n3288# 0.328811f
C682 source.t47 a_n2094_n3288# 0.328811f
C683 source.n494 a_n2094_n3288# 2.81527f
C684 source.n495 a_n2094_n3288# 0.456618f
C685 source.t4 a_n2094_n3288# 0.328811f
C686 source.t43 a_n2094_n3288# 0.328811f
C687 source.n496 a_n2094_n3288# 2.81527f
C688 source.n497 a_n2094_n3288# 0.456618f
C689 source.t1 a_n2094_n3288# 0.328811f
C690 source.t33 a_n2094_n3288# 0.328811f
C691 source.n498 a_n2094_n3288# 2.81527f
C692 source.n499 a_n2094_n3288# 0.456618f
C693 source.t32 a_n2094_n3288# 0.328811f
C694 source.t45 a_n2094_n3288# 0.328811f
C695 source.n500 a_n2094_n3288# 2.81527f
C696 source.n501 a_n2094_n3288# 0.456618f
C697 source.n502 a_n2094_n3288# 0.045931f
C698 source.n503 a_n2094_n3288# 0.034675f
C699 source.n504 a_n2094_n3288# 0.018633f
C700 source.n505 a_n2094_n3288# 0.044041f
C701 source.n506 a_n2094_n3288# 0.019729f
C702 source.n507 a_n2094_n3288# 0.034675f
C703 source.n508 a_n2094_n3288# 0.018633f
C704 source.n509 a_n2094_n3288# 0.044041f
C705 source.n510 a_n2094_n3288# 0.019729f
C706 source.n511 a_n2094_n3288# 0.034675f
C707 source.n512 a_n2094_n3288# 0.019181f
C708 source.n513 a_n2094_n3288# 0.044041f
C709 source.n514 a_n2094_n3288# 0.019729f
C710 source.n515 a_n2094_n3288# 0.034675f
C711 source.n516 a_n2094_n3288# 0.018633f
C712 source.n517 a_n2094_n3288# 0.044041f
C713 source.n518 a_n2094_n3288# 0.019729f
C714 source.n519 a_n2094_n3288# 0.034675f
C715 source.n520 a_n2094_n3288# 0.018633f
C716 source.n521 a_n2094_n3288# 0.033031f
C717 source.n522 a_n2094_n3288# 0.031133f
C718 source.t5 a_n2094_n3288# 0.074382f
C719 source.n523 a_n2094_n3288# 0.25f
C720 source.n524 a_n2094_n3288# 1.74928f
C721 source.n525 a_n2094_n3288# 0.018633f
C722 source.n526 a_n2094_n3288# 0.019729f
C723 source.n527 a_n2094_n3288# 0.044041f
C724 source.n528 a_n2094_n3288# 0.044041f
C725 source.n529 a_n2094_n3288# 0.019729f
C726 source.n530 a_n2094_n3288# 0.018633f
C727 source.n531 a_n2094_n3288# 0.034675f
C728 source.n532 a_n2094_n3288# 0.034675f
C729 source.n533 a_n2094_n3288# 0.018633f
C730 source.n534 a_n2094_n3288# 0.019729f
C731 source.n535 a_n2094_n3288# 0.044041f
C732 source.n536 a_n2094_n3288# 0.044041f
C733 source.n537 a_n2094_n3288# 0.019729f
C734 source.n538 a_n2094_n3288# 0.018633f
C735 source.n539 a_n2094_n3288# 0.034675f
C736 source.n540 a_n2094_n3288# 0.034675f
C737 source.n541 a_n2094_n3288# 0.018633f
C738 source.n542 a_n2094_n3288# 0.018633f
C739 source.n543 a_n2094_n3288# 0.019729f
C740 source.n544 a_n2094_n3288# 0.044041f
C741 source.n545 a_n2094_n3288# 0.044041f
C742 source.n546 a_n2094_n3288# 0.044041f
C743 source.n547 a_n2094_n3288# 0.019181f
C744 source.n548 a_n2094_n3288# 0.018633f
C745 source.n549 a_n2094_n3288# 0.034675f
C746 source.n550 a_n2094_n3288# 0.034675f
C747 source.n551 a_n2094_n3288# 0.018633f
C748 source.n552 a_n2094_n3288# 0.019729f
C749 source.n553 a_n2094_n3288# 0.044041f
C750 source.n554 a_n2094_n3288# 0.044041f
C751 source.n555 a_n2094_n3288# 0.019729f
C752 source.n556 a_n2094_n3288# 0.018633f
C753 source.n557 a_n2094_n3288# 0.034675f
C754 source.n558 a_n2094_n3288# 0.034675f
C755 source.n559 a_n2094_n3288# 0.018633f
C756 source.n560 a_n2094_n3288# 0.019729f
C757 source.n561 a_n2094_n3288# 0.044041f
C758 source.n562 a_n2094_n3288# 0.090376f
C759 source.n563 a_n2094_n3288# 0.019729f
C760 source.n564 a_n2094_n3288# 0.018633f
C761 source.n565 a_n2094_n3288# 0.074464f
C762 source.n566 a_n2094_n3288# 0.049878f
C763 source.n567 a_n2094_n3288# 0.317972f
C764 source.n568 a_n2094_n3288# 2.16991f
C765 drain_left.t12 a_n2094_n3288# 0.370932f
C766 drain_left.t22 a_n2094_n3288# 0.370932f
C767 drain_left.n0 a_n2094_n3288# 3.30422f
C768 drain_left.t3 a_n2094_n3288# 0.370932f
C769 drain_left.t23 a_n2094_n3288# 0.370932f
C770 drain_left.n1 a_n2094_n3288# 3.30072f
C771 drain_left.n2 a_n2094_n3288# 0.899186f
C772 drain_left.t7 a_n2094_n3288# 0.370932f
C773 drain_left.t11 a_n2094_n3288# 0.370932f
C774 drain_left.n3 a_n2094_n3288# 3.30072f
C775 drain_left.n4 a_n2094_n3288# 0.412932f
C776 drain_left.t2 a_n2094_n3288# 0.370932f
C777 drain_left.t21 a_n2094_n3288# 0.370932f
C778 drain_left.n5 a_n2094_n3288# 3.30422f
C779 drain_left.t5 a_n2094_n3288# 0.370932f
C780 drain_left.t19 a_n2094_n3288# 0.370932f
C781 drain_left.n6 a_n2094_n3288# 3.30072f
C782 drain_left.n7 a_n2094_n3288# 0.899186f
C783 drain_left.t8 a_n2094_n3288# 0.370932f
C784 drain_left.t18 a_n2094_n3288# 0.370932f
C785 drain_left.n8 a_n2094_n3288# 3.30072f
C786 drain_left.n9 a_n2094_n3288# 0.412932f
C787 drain_left.n10 a_n2094_n3288# 2.00625f
C788 drain_left.t9 a_n2094_n3288# 0.370932f
C789 drain_left.t13 a_n2094_n3288# 0.370932f
C790 drain_left.n11 a_n2094_n3288# 3.30423f
C791 drain_left.t0 a_n2094_n3288# 0.370932f
C792 drain_left.t16 a_n2094_n3288# 0.370932f
C793 drain_left.n12 a_n2094_n3288# 3.30074f
C794 drain_left.n13 a_n2094_n3288# 0.899159f
C795 drain_left.t17 a_n2094_n3288# 0.370932f
C796 drain_left.t10 a_n2094_n3288# 0.370932f
C797 drain_left.n14 a_n2094_n3288# 3.30074f
C798 drain_left.n15 a_n2094_n3288# 0.44345f
C799 drain_left.t14 a_n2094_n3288# 0.370932f
C800 drain_left.t1 a_n2094_n3288# 0.370932f
C801 drain_left.n16 a_n2094_n3288# 3.30074f
C802 drain_left.n17 a_n2094_n3288# 0.44345f
C803 drain_left.t6 a_n2094_n3288# 0.370932f
C804 drain_left.t4 a_n2094_n3288# 0.370932f
C805 drain_left.n18 a_n2094_n3288# 3.30074f
C806 drain_left.n19 a_n2094_n3288# 0.44345f
C807 drain_left.t15 a_n2094_n3288# 0.370932f
C808 drain_left.t20 a_n2094_n3288# 0.370932f
C809 drain_left.n20 a_n2094_n3288# 3.30072f
C810 drain_left.n21 a_n2094_n3288# 0.763595f
C811 plus.n0 a_n2094_n3288# 0.052523f
C812 plus.t0 a_n2094_n3288# 0.356207f
C813 plus.t3 a_n2094_n3288# 0.356207f
C814 plus.t11 a_n2094_n3288# 0.356207f
C815 plus.n1 a_n2094_n3288# 0.146702f
C816 plus.n2 a_n2094_n3288# 0.052523f
C817 plus.t21 a_n2094_n3288# 0.356207f
C818 plus.t1 a_n2094_n3288# 0.356207f
C819 plus.t5 a_n2094_n3288# 0.356207f
C820 plus.n3 a_n2094_n3288# 0.146702f
C821 plus.n4 a_n2094_n3288# 0.052523f
C822 plus.t13 a_n2094_n3288# 0.356207f
C823 plus.t14 a_n2094_n3288# 0.356207f
C824 plus.t22 a_n2094_n3288# 0.356207f
C825 plus.n5 a_n2094_n3288# 0.146702f
C826 plus.t6 a_n2094_n3288# 0.361689f
C827 plus.n6 a_n2094_n3288# 0.163421f
C828 plus.t2 a_n2094_n3288# 0.356207f
C829 plus.n7 a_n2094_n3288# 0.146702f
C830 plus.n8 a_n2094_n3288# 0.018395f
C831 plus.n9 a_n2094_n3288# 0.122126f
C832 plus.n10 a_n2094_n3288# 0.052523f
C833 plus.n11 a_n2094_n3288# 0.018395f
C834 plus.n12 a_n2094_n3288# 0.146702f
C835 plus.n13 a_n2094_n3288# 0.018395f
C836 plus.n14 a_n2094_n3288# 0.146702f
C837 plus.n15 a_n2094_n3288# 0.018395f
C838 plus.n16 a_n2094_n3288# 0.052523f
C839 plus.n17 a_n2094_n3288# 0.052523f
C840 plus.n18 a_n2094_n3288# 0.018395f
C841 plus.n19 a_n2094_n3288# 0.146702f
C842 plus.n20 a_n2094_n3288# 0.018395f
C843 plus.n21 a_n2094_n3288# 0.146702f
C844 plus.n22 a_n2094_n3288# 0.018395f
C845 plus.n23 a_n2094_n3288# 0.052523f
C846 plus.n24 a_n2094_n3288# 0.052523f
C847 plus.n25 a_n2094_n3288# 0.018395f
C848 plus.n26 a_n2094_n3288# 0.146702f
C849 plus.n27 a_n2094_n3288# 0.018395f
C850 plus.n28 a_n2094_n3288# 0.146702f
C851 plus.t20 a_n2094_n3288# 0.361689f
C852 plus.n29 a_n2094_n3288# 0.163339f
C853 plus.n30 a_n2094_n3288# 0.586283f
C854 plus.n31 a_n2094_n3288# 0.052523f
C855 plus.t15 a_n2094_n3288# 0.361689f
C856 plus.t8 a_n2094_n3288# 0.356207f
C857 plus.t4 a_n2094_n3288# 0.356207f
C858 plus.t7 a_n2094_n3288# 0.356207f
C859 plus.n32 a_n2094_n3288# 0.146702f
C860 plus.n33 a_n2094_n3288# 0.052523f
C861 plus.t10 a_n2094_n3288# 0.356207f
C862 plus.t16 a_n2094_n3288# 0.356207f
C863 plus.t9 a_n2094_n3288# 0.356207f
C864 plus.n34 a_n2094_n3288# 0.146702f
C865 plus.n35 a_n2094_n3288# 0.052523f
C866 plus.t18 a_n2094_n3288# 0.356207f
C867 plus.t12 a_n2094_n3288# 0.356207f
C868 plus.t17 a_n2094_n3288# 0.356207f
C869 plus.n36 a_n2094_n3288# 0.146702f
C870 plus.t19 a_n2094_n3288# 0.361689f
C871 plus.n37 a_n2094_n3288# 0.163421f
C872 plus.t23 a_n2094_n3288# 0.356207f
C873 plus.n38 a_n2094_n3288# 0.146702f
C874 plus.n39 a_n2094_n3288# 0.018395f
C875 plus.n40 a_n2094_n3288# 0.122126f
C876 plus.n41 a_n2094_n3288# 0.052523f
C877 plus.n42 a_n2094_n3288# 0.018395f
C878 plus.n43 a_n2094_n3288# 0.146702f
C879 plus.n44 a_n2094_n3288# 0.018395f
C880 plus.n45 a_n2094_n3288# 0.146702f
C881 plus.n46 a_n2094_n3288# 0.018395f
C882 plus.n47 a_n2094_n3288# 0.052523f
C883 plus.n48 a_n2094_n3288# 0.052523f
C884 plus.n49 a_n2094_n3288# 0.018395f
C885 plus.n50 a_n2094_n3288# 0.146702f
C886 plus.n51 a_n2094_n3288# 0.018395f
C887 plus.n52 a_n2094_n3288# 0.146702f
C888 plus.n53 a_n2094_n3288# 0.018395f
C889 plus.n54 a_n2094_n3288# 0.052523f
C890 plus.n55 a_n2094_n3288# 0.052523f
C891 plus.n56 a_n2094_n3288# 0.018395f
C892 plus.n57 a_n2094_n3288# 0.146702f
C893 plus.n58 a_n2094_n3288# 0.018395f
C894 plus.n59 a_n2094_n3288# 0.146702f
C895 plus.n60 a_n2094_n3288# 0.163339f
C896 plus.n61 a_n2094_n3288# 1.63009f
.ends

