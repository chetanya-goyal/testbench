* NGSPICE file created from diffpair593.ext - technology: sky130A

.subckt diffpair593 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t12 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 drain_left.t6 plus.t1 source.t11 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X2 drain_right.t7 minus.t0 source.t15 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X3 source.t0 minus.t1 drain_right.t6 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X4 source.t5 minus.t2 drain_right.t5 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X5 source.t13 plus.t2 drain_left.t5 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X6 a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X7 a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X8 a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X9 drain_left.t4 plus.t3 source.t6 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X10 source.t2 minus.t3 drain_right.t4 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X11 drain_right.t3 minus.t4 source.t3 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X12 source.t9 plus.t4 drain_left.t3 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X13 source.t10 plus.t5 drain_left.t2 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X14 source.t8 plus.t6 drain_left.t1 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X15 drain_right.t2 minus.t5 source.t4 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X16 drain_right.t1 minus.t6 source.t1 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X17 source.t14 minus.t7 drain_right.t0 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X18 a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X19 drain_left.t0 plus.t7 source.t7 a_n1346_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
R0 plus.n2 plus.t2 1739.58
R1 plus.n7 plus.t7 1739.58
R2 plus.n11 plus.t0 1739.58
R3 plus.n16 plus.t6 1739.58
R4 plus.n1 plus.t3 1711.1
R5 plus.n6 plus.t5 1711.1
R6 plus.n10 plus.t4 1711.1
R7 plus.n15 plus.t1 1711.1
R8 plus.n3 plus.n2 161.489
R9 plus.n12 plus.n11 161.489
R10 plus.n4 plus.n3 161.3
R11 plus.n5 plus.n0 161.3
R12 plus.n8 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n14 plus.n9 161.3
R15 plus.n17 plus.n16 161.3
R16 plus.n5 plus.n4 73.0308
R17 plus.n14 plus.n13 73.0308
R18 plus.n2 plus.n1 63.5369
R19 plus.n7 plus.n6 63.5369
R20 plus.n16 plus.n15 63.5369
R21 plus.n11 plus.n10 63.5369
R22 plus plus.n17 31.0937
R23 plus plus.n8 15.1369
R24 plus.n4 plus.n1 9.49444
R25 plus.n6 plus.n5 9.49444
R26 plus.n15 plus.n14 9.49444
R27 plus.n13 plus.n10 9.49444
R28 plus.n3 plus.n0 0.189894
R29 plus.n8 plus.n0 0.189894
R30 plus.n17 plus.n9 0.189894
R31 plus.n12 plus.n9 0.189894
R32 source.n0 source.t7 44.1297
R33 source.n3 source.t13 44.1296
R34 source.n4 source.t3 44.1296
R35 source.n7 source.t2 44.1296
R36 source.n15 source.t4 44.1295
R37 source.n12 source.t5 44.1295
R38 source.n11 source.t12 44.1295
R39 source.n8 source.t8 44.1295
R40 source.n2 source.n1 43.1397
R41 source.n6 source.n5 43.1397
R42 source.n14 source.n13 43.1396
R43 source.n10 source.n9 43.1396
R44 source.n8 source.n7 27.8914
R45 source.n16 source.n0 22.357
R46 source.n16 source.n15 5.53498
R47 source.n13 source.t1 0.9905
R48 source.n13 source.t0 0.9905
R49 source.n9 source.t11 0.9905
R50 source.n9 source.t9 0.9905
R51 source.n1 source.t6 0.9905
R52 source.n1 source.t10 0.9905
R53 source.n5 source.t15 0.9905
R54 source.n5 source.t14 0.9905
R55 source.n7 source.n6 0.543603
R56 source.n6 source.n4 0.543603
R57 source.n3 source.n2 0.543603
R58 source.n2 source.n0 0.543603
R59 source.n10 source.n8 0.543603
R60 source.n11 source.n10 0.543603
R61 source.n14 source.n12 0.543603
R62 source.n15 source.n14 0.543603
R63 source.n4 source.n3 0.470328
R64 source.n12 source.n11 0.470328
R65 source source.n16 0.188
R66 drain_left.n5 drain_left.n3 60.3616
R67 drain_left.n2 drain_left.n1 60.0346
R68 drain_left.n2 drain_left.n0 60.0346
R69 drain_left.n5 drain_left.n4 59.8185
R70 drain_left drain_left.n2 35.3285
R71 drain_left drain_left.n5 6.19632
R72 drain_left.n1 drain_left.t3 0.9905
R73 drain_left.n1 drain_left.t7 0.9905
R74 drain_left.n0 drain_left.t1 0.9905
R75 drain_left.n0 drain_left.t6 0.9905
R76 drain_left.n4 drain_left.t2 0.9905
R77 drain_left.n4 drain_left.t0 0.9905
R78 drain_left.n3 drain_left.t5 0.9905
R79 drain_left.n3 drain_left.t4 0.9905
R80 minus.n7 minus.t3 1739.58
R81 minus.n2 minus.t4 1739.58
R82 minus.n16 minus.t5 1739.58
R83 minus.n11 minus.t2 1739.58
R84 minus.n6 minus.t0 1711.1
R85 minus.n1 minus.t7 1711.1
R86 minus.n15 minus.t1 1711.1
R87 minus.n10 minus.t6 1711.1
R88 minus.n3 minus.n2 161.489
R89 minus.n12 minus.n11 161.489
R90 minus.n8 minus.n7 161.3
R91 minus.n5 minus.n0 161.3
R92 minus.n4 minus.n3 161.3
R93 minus.n17 minus.n16 161.3
R94 minus.n14 minus.n9 161.3
R95 minus.n13 minus.n12 161.3
R96 minus.n5 minus.n4 73.0308
R97 minus.n14 minus.n13 73.0308
R98 minus.n7 minus.n6 63.5369
R99 minus.n2 minus.n1 63.5369
R100 minus.n11 minus.n10 63.5369
R101 minus.n16 minus.n15 63.5369
R102 minus.n18 minus.n8 40.2429
R103 minus.n6 minus.n5 9.49444
R104 minus.n4 minus.n1 9.49444
R105 minus.n13 minus.n10 9.49444
R106 minus.n15 minus.n14 9.49444
R107 minus.n18 minus.n17 6.46262
R108 minus.n8 minus.n0 0.189894
R109 minus.n3 minus.n0 0.189894
R110 minus.n12 minus.n9 0.189894
R111 minus.n17 minus.n9 0.189894
R112 minus minus.n18 0.188
R113 drain_right.n5 drain_right.n3 60.3616
R114 drain_right.n2 drain_right.n1 60.0346
R115 drain_right.n2 drain_right.n0 60.0346
R116 drain_right.n5 drain_right.n4 59.8185
R117 drain_right drain_right.n2 34.7753
R118 drain_right drain_right.n5 6.19632
R119 drain_right.n1 drain_right.t6 0.9905
R120 drain_right.n1 drain_right.t2 0.9905
R121 drain_right.n0 drain_right.t5 0.9905
R122 drain_right.n0 drain_right.t1 0.9905
R123 drain_right.n3 drain_right.t0 0.9905
R124 drain_right.n3 drain_right.t3 0.9905
R125 drain_right.n4 drain_right.t4 0.9905
R126 drain_right.n4 drain_right.t7 0.9905
C0 drain_left source 26.3913f
C1 plus drain_right 0.280736f
C2 drain_right source 26.390501f
C3 drain_right drain_left 0.630082f
C4 plus minus 6.31364f
C5 source minus 4.59169f
C6 drain_left minus 0.170671f
C7 drain_right minus 5.36903f
C8 plus source 4.60573f
C9 plus drain_left 5.49623f
C10 drain_right a_n1346_n4888# 7.48655f
C11 drain_left a_n1346_n4888# 7.685009f
C12 source a_n1346_n4888# 12.910511f
C13 minus a_n1346_n4888# 5.725986f
C14 plus a_n1346_n4888# 8.30243f
C15 drain_right.t5 a_n1346_n4888# 0.532632f
C16 drain_right.t1 a_n1346_n4888# 0.532632f
C17 drain_right.n0 a_n1346_n4888# 4.87082f
C18 drain_right.t6 a_n1346_n4888# 0.532632f
C19 drain_right.t2 a_n1346_n4888# 0.532632f
C20 drain_right.n1 a_n1346_n4888# 4.87082f
C21 drain_right.n2 a_n1346_n4888# 2.83242f
C22 drain_right.t0 a_n1346_n4888# 0.532632f
C23 drain_right.t3 a_n1346_n4888# 0.532632f
C24 drain_right.n3 a_n1346_n4888# 4.87317f
C25 drain_right.t4 a_n1346_n4888# 0.532632f
C26 drain_right.t7 a_n1346_n4888# 0.532632f
C27 drain_right.n4 a_n1346_n4888# 4.86943f
C28 drain_right.n5 a_n1346_n4888# 1.09504f
C29 minus.n0 a_n1346_n4888# 0.055576f
C30 minus.t3 a_n1346_n4888# 0.94488f
C31 minus.t0 a_n1346_n4888# 0.939171f
C32 minus.t7 a_n1346_n4888# 0.939171f
C33 minus.n1 a_n1346_n4888# 0.348879f
C34 minus.t4 a_n1346_n4888# 0.94488f
C35 minus.n2 a_n1346_n4888# 0.365962f
C36 minus.n3 a_n1346_n4888# 0.117589f
C37 minus.n4 a_n1346_n4888# 0.020664f
C38 minus.n5 a_n1346_n4888# 0.020664f
C39 minus.n6 a_n1346_n4888# 0.348879f
C40 minus.n7 a_n1346_n4888# 0.36589f
C41 minus.n8 a_n1346_n4888# 2.30852f
C42 minus.n9 a_n1346_n4888# 0.055576f
C43 minus.t1 a_n1346_n4888# 0.939171f
C44 minus.t6 a_n1346_n4888# 0.939171f
C45 minus.n10 a_n1346_n4888# 0.348879f
C46 minus.t2 a_n1346_n4888# 0.94488f
C47 minus.n11 a_n1346_n4888# 0.365962f
C48 minus.n12 a_n1346_n4888# 0.117589f
C49 minus.n13 a_n1346_n4888# 0.020664f
C50 minus.n14 a_n1346_n4888# 0.020664f
C51 minus.n15 a_n1346_n4888# 0.348879f
C52 minus.t5 a_n1346_n4888# 0.94488f
C53 minus.n16 a_n1346_n4888# 0.36589f
C54 minus.n17 a_n1346_n4888# 0.358438f
C55 minus.n18 a_n1346_n4888# 2.77214f
C56 drain_left.t1 a_n1346_n4888# 0.532101f
C57 drain_left.t6 a_n1346_n4888# 0.532101f
C58 drain_left.n0 a_n1346_n4888# 4.86596f
C59 drain_left.t3 a_n1346_n4888# 0.532101f
C60 drain_left.t7 a_n1346_n4888# 0.532101f
C61 drain_left.n1 a_n1346_n4888# 4.86596f
C62 drain_left.n2 a_n1346_n4888# 2.90023f
C63 drain_left.t5 a_n1346_n4888# 0.532101f
C64 drain_left.t4 a_n1346_n4888# 0.532101f
C65 drain_left.n3 a_n1346_n4888# 4.86832f
C66 drain_left.t2 a_n1346_n4888# 0.532101f
C67 drain_left.t0 a_n1346_n4888# 0.532101f
C68 drain_left.n4 a_n1346_n4888# 4.86458f
C69 drain_left.n5 a_n1346_n4888# 1.09395f
C70 source.t7 a_n1346_n4888# 4.23942f
C71 source.n0 a_n1346_n4888# 1.80317f
C72 source.t6 a_n1346_n4888# 0.370956f
C73 source.t10 a_n1346_n4888# 0.370956f
C74 source.n1 a_n1346_n4888# 3.3165f
C75 source.n2 a_n1346_n4888# 0.323168f
C76 source.t13 a_n1346_n4888# 4.23943f
C77 source.n3 a_n1346_n4888# 0.406395f
C78 source.t3 a_n1346_n4888# 4.23943f
C79 source.n4 a_n1346_n4888# 0.406395f
C80 source.t15 a_n1346_n4888# 0.370956f
C81 source.t14 a_n1346_n4888# 0.370956f
C82 source.n5 a_n1346_n4888# 3.3165f
C83 source.n6 a_n1346_n4888# 0.323168f
C84 source.t2 a_n1346_n4888# 4.23943f
C85 source.n7 a_n1346_n4888# 2.21911f
C86 source.t8 a_n1346_n4888# 4.23941f
C87 source.n8 a_n1346_n4888# 2.21913f
C88 source.t11 a_n1346_n4888# 0.370956f
C89 source.t9 a_n1346_n4888# 0.370956f
C90 source.n9 a_n1346_n4888# 3.31651f
C91 source.n10 a_n1346_n4888# 0.323162f
C92 source.t12 a_n1346_n4888# 4.23941f
C93 source.n11 a_n1346_n4888# 0.406418f
C94 source.t5 a_n1346_n4888# 4.23941f
C95 source.n12 a_n1346_n4888# 0.406418f
C96 source.t1 a_n1346_n4888# 0.370956f
C97 source.t0 a_n1346_n4888# 0.370956f
C98 source.n13 a_n1346_n4888# 3.31651f
C99 source.n14 a_n1346_n4888# 0.323162f
C100 source.t4 a_n1346_n4888# 4.23941f
C101 source.n15 a_n1346_n4888# 0.538914f
C102 source.n16 a_n1346_n4888# 2.11286f
C103 plus.n0 a_n1346_n4888# 0.056305f
C104 plus.t5 a_n1346_n4888# 0.951493f
C105 plus.t3 a_n1346_n4888# 0.951493f
C106 plus.n1 a_n1346_n4888# 0.353457f
C107 plus.t2 a_n1346_n4888# 0.957277f
C108 plus.n2 a_n1346_n4888# 0.370764f
C109 plus.n3 a_n1346_n4888# 0.119132f
C110 plus.n4 a_n1346_n4888# 0.020935f
C111 plus.n5 a_n1346_n4888# 0.020935f
C112 plus.n6 a_n1346_n4888# 0.353457f
C113 plus.t7 a_n1346_n4888# 0.957277f
C114 plus.n7 a_n1346_n4888# 0.37069f
C115 plus.n8 a_n1346_n4888# 0.85011f
C116 plus.n9 a_n1346_n4888# 0.056305f
C117 plus.t6 a_n1346_n4888# 0.957277f
C118 plus.t1 a_n1346_n4888# 0.951493f
C119 plus.t4 a_n1346_n4888# 0.951493f
C120 plus.n10 a_n1346_n4888# 0.353457f
C121 plus.t0 a_n1346_n4888# 0.957277f
C122 plus.n11 a_n1346_n4888# 0.370764f
C123 plus.n12 a_n1346_n4888# 0.119132f
C124 plus.n13 a_n1346_n4888# 0.020935f
C125 plus.n14 a_n1346_n4888# 0.020935f
C126 plus.n15 a_n1346_n4888# 0.353457f
C127 plus.n16 a_n1346_n4888# 0.37069f
C128 plus.n17 a_n1346_n4888# 1.83591f
.ends

