* NGSPICE file created from diffpair515.ext - technology: sky130A

.subckt diffpair515 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t8 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X1 drain_left.t11 plus.t0 source.t9 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X2 drain_left.t10 plus.t1 source.t0 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X3 drain_right.t7 minus.t1 source.t22 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X4 a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X5 source.t8 plus.t2 drain_left.t9 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X6 source.t21 minus.t2 drain_right.t2 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X7 source.t20 minus.t3 drain_right.t0 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X8 a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X9 drain_left.t8 plus.t3 source.t11 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X10 source.t1 plus.t4 drain_left.t7 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X11 a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X12 a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X13 drain_left.t6 plus.t5 source.t2 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X14 source.t19 minus.t4 drain_right.t10 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X15 source.t18 minus.t5 drain_right.t3 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X16 drain_right.t1 minus.t6 source.t17 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X17 drain_left.t5 plus.t6 source.t3 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X18 source.t7 plus.t7 drain_left.t4 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X19 source.t10 plus.t8 drain_left.t3 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X20 source.t4 plus.t9 drain_left.t2 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X21 source.t6 plus.t10 drain_left.t1 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X22 drain_right.t9 minus.t7 source.t16 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 drain_right.t6 minus.t8 source.t15 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X24 drain_right.t5 minus.t9 source.t14 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X25 source.t13 minus.t10 drain_right.t11 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X26 drain_right.t4 minus.t11 source.t12 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X27 drain_left.t0 plus.t11 source.t5 a_n1598_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 minus.n13 minus.t0 1356.9
R1 minus.n2 minus.t6 1356.9
R2 minus.n28 minus.t11 1356.9
R3 minus.n17 minus.t3 1356.9
R4 minus.n12 minus.t7 1309.43
R5 minus.n10 minus.t4 1309.43
R6 minus.n3 minus.t1 1309.43
R7 minus.n4 minus.t10 1309.43
R8 minus.n27 minus.t5 1309.43
R9 minus.n25 minus.t8 1309.43
R10 minus.n19 minus.t2 1309.43
R11 minus.n18 minus.t9 1309.43
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n13 minus.n12 44.549
R31 minus.n4 minus.n2 44.549
R32 minus.n18 minus.n17 44.549
R33 minus.n28 minus.n27 44.549
R34 minus.n30 minus.n14 37.4588
R35 minus.n12 minus.n11 28.4823
R36 minus.n5 minus.n4 28.4823
R37 minus.n20 minus.n18 28.4823
R38 minus.n27 minus.n26 28.4823
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 61.4227
R54 drain_right.n3 drain_right.n2 61.3673
R55 drain_right.n3 drain_right.n0 61.3673
R56 drain_right.n6 drain_right.n5 60.8798
R57 drain_right.n8 drain_right.n7 60.8798
R58 drain_right.n3 drain_right.n1 60.8796
R59 drain_right drain_right.n3 31.8021
R60 drain_right drain_right.n8 6.19632
R61 drain_right.n1 drain_right.t2 1.3205
R62 drain_right.n1 drain_right.t6 1.3205
R63 drain_right.n2 drain_right.t3 1.3205
R64 drain_right.n2 drain_right.t4 1.3205
R65 drain_right.n0 drain_right.t0 1.3205
R66 drain_right.n0 drain_right.t5 1.3205
R67 drain_right.n4 drain_right.t11 1.3205
R68 drain_right.n4 drain_right.t1 1.3205
R69 drain_right.n5 drain_right.t10 1.3205
R70 drain_right.n5 drain_right.t7 1.3205
R71 drain_right.n7 drain_right.t8 1.3205
R72 drain_right.n7 drain_right.t9 1.3205
R73 drain_right.n8 drain_right.n6 0.543603
R74 source.n5 source.t8 45.521
R75 source.n6 source.t17 45.521
R76 source.n11 source.t23 45.521
R77 source.n23 source.t12 45.5208
R78 source.n18 source.t20 45.5208
R79 source.n17 source.t9 45.5208
R80 source.n12 source.t6 45.5208
R81 source.n0 source.t3 45.5208
R82 source.n2 source.n1 44.201
R83 source.n4 source.n3 44.201
R84 source.n8 source.n7 44.201
R85 source.n10 source.n9 44.201
R86 source.n22 source.n21 44.2008
R87 source.n20 source.n19 44.2008
R88 source.n16 source.n15 44.2008
R89 source.n14 source.n13 44.2008
R90 source.n12 source.n11 24.1036
R91 source.n24 source.n0 18.5691
R92 source.n24 source.n23 5.53498
R93 source.n21 source.t15 1.3205
R94 source.n21 source.t18 1.3205
R95 source.n19 source.t14 1.3205
R96 source.n19 source.t21 1.3205
R97 source.n15 source.t0 1.3205
R98 source.n15 source.t7 1.3205
R99 source.n13 source.t11 1.3205
R100 source.n13 source.t4 1.3205
R101 source.n1 source.t5 1.3205
R102 source.n1 source.t1 1.3205
R103 source.n3 source.t2 1.3205
R104 source.n3 source.t10 1.3205
R105 source.n7 source.t22 1.3205
R106 source.n7 source.t13 1.3205
R107 source.n9 source.t16 1.3205
R108 source.n9 source.t19 1.3205
R109 source.n11 source.n10 0.543603
R110 source.n10 source.n8 0.543603
R111 source.n8 source.n6 0.543603
R112 source.n5 source.n4 0.543603
R113 source.n4 source.n2 0.543603
R114 source.n2 source.n0 0.543603
R115 source.n14 source.n12 0.543603
R116 source.n16 source.n14 0.543603
R117 source.n17 source.n16 0.543603
R118 source.n20 source.n18 0.543603
R119 source.n22 source.n20 0.543603
R120 source.n23 source.n22 0.543603
R121 source.n6 source.n5 0.470328
R122 source.n18 source.n17 0.470328
R123 source source.n24 0.188
R124 plus.n2 plus.t2 1356.9
R125 plus.n13 plus.t6 1356.9
R126 plus.n17 plus.t0 1356.9
R127 plus.n28 plus.t10 1356.9
R128 plus.n3 plus.t5 1309.43
R129 plus.n4 plus.t8 1309.43
R130 plus.n10 plus.t11 1309.43
R131 plus.n12 plus.t4 1309.43
R132 plus.n19 plus.t7 1309.43
R133 plus.n18 plus.t1 1309.43
R134 plus.n25 plus.t9 1309.43
R135 plus.n27 plus.t3 1309.43
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 63.5369
R151 plus.n11 plus.n10 63.5369
R152 plus.n26 plus.n25 63.5369
R153 plus.n20 plus.n18 63.5369
R154 plus.n3 plus.n2 44.549
R155 plus.n13 plus.n12 44.549
R156 plus.n28 plus.n27 44.549
R157 plus.n19 plus.n17 44.549
R158 plus plus.n29 30.2036
R159 plus.n5 plus.n3 28.4823
R160 plus.n12 plus.n11 28.4823
R161 plus.n27 plus.n26 28.4823
R162 plus.n20 plus.n19 28.4823
R163 plus plus.n14 13.2922
R164 plus.n4 plus.n1 9.49444
R165 plus.n10 plus.n9 9.49444
R166 plus.n25 plus.n24 9.49444
R167 plus.n18 plus.n16 9.49444
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 61.4229
R177 drain_left.n3 drain_left.n2 61.3673
R178 drain_left.n3 drain_left.n0 61.3673
R179 drain_left.n6 drain_left.n5 60.8798
R180 drain_left.n8 drain_left.n7 60.8796
R181 drain_left.n3 drain_left.n1 60.8796
R182 drain_left drain_left.n3 32.3553
R183 drain_left drain_left.n8 6.19632
R184 drain_left.n1 drain_left.t2 1.3205
R185 drain_left.n1 drain_left.t10 1.3205
R186 drain_left.n2 drain_left.t4 1.3205
R187 drain_left.n2 drain_left.t11 1.3205
R188 drain_left.n0 drain_left.t1 1.3205
R189 drain_left.n0 drain_left.t8 1.3205
R190 drain_left.n7 drain_left.t7 1.3205
R191 drain_left.n7 drain_left.t5 1.3205
R192 drain_left.n5 drain_left.t3 1.3205
R193 drain_left.n5 drain_left.t0 1.3205
R194 drain_left.n4 drain_left.t9 1.3205
R195 drain_left.n4 drain_left.t6 1.3205
R196 drain_left.n8 drain_left.n6 0.543603
C0 minus plus 5.69908f
C1 source drain_right 28.826199f
C2 source minus 5.18261f
C3 source plus 5.19665f
C4 drain_right drain_left 0.785787f
C5 minus drain_left 0.170859f
C6 plus drain_left 5.84038f
C7 minus drain_right 5.68692f
C8 plus drain_right 0.30725f
C9 source drain_left 28.8265f
C10 drain_right a_n1598_n3888# 6.81141f
C11 drain_left a_n1598_n3888# 7.05815f
C12 source a_n1598_n3888# 10.258769f
C13 minus a_n1598_n3888# 6.401933f
C14 plus a_n1598_n3888# 8.58194f
C15 drain_left.t1 a_n1598_n3888# 0.400428f
C16 drain_left.t8 a_n1598_n3888# 0.400428f
C17 drain_left.n0 a_n1598_n3888# 3.62261f
C18 drain_left.t2 a_n1598_n3888# 0.400428f
C19 drain_left.t10 a_n1598_n3888# 0.400428f
C20 drain_left.n1 a_n1598_n3888# 3.6194f
C21 drain_left.t4 a_n1598_n3888# 0.400428f
C22 drain_left.t11 a_n1598_n3888# 0.400428f
C23 drain_left.n2 a_n1598_n3888# 3.62261f
C24 drain_left.n3 a_n1598_n3888# 2.94965f
C25 drain_left.t9 a_n1598_n3888# 0.400428f
C26 drain_left.t6 a_n1598_n3888# 0.400428f
C27 drain_left.n4 a_n1598_n3888# 3.62301f
C28 drain_left.t3 a_n1598_n3888# 0.400428f
C29 drain_left.t0 a_n1598_n3888# 0.400428f
C30 drain_left.n5 a_n1598_n3888# 3.6194f
C31 drain_left.n6 a_n1598_n3888# 0.799841f
C32 drain_left.t7 a_n1598_n3888# 0.400428f
C33 drain_left.t5 a_n1598_n3888# 0.400428f
C34 drain_left.n7 a_n1598_n3888# 3.61939f
C35 drain_left.n8 a_n1598_n3888# 0.676121f
C36 plus.n0 a_n1598_n3888# 0.053167f
C37 plus.t4 a_n1598_n3888# 0.674969f
C38 plus.t11 a_n1598_n3888# 0.674969f
C39 plus.n1 a_n1598_n3888# 0.019768f
C40 plus.t2 a_n1598_n3888# 0.684182f
C41 plus.n2 a_n1598_n3888# 0.276122f
C42 plus.t5 a_n1598_n3888# 0.674969f
C43 plus.n3 a_n1598_n3888# 0.25926f
C44 plus.t8 a_n1598_n3888# 0.674969f
C45 plus.n4 a_n1598_n3888# 0.25926f
C46 plus.n5 a_n1598_n3888# 0.021899f
C47 plus.n6 a_n1598_n3888# 0.121006f
C48 plus.n7 a_n1598_n3888# 0.053167f
C49 plus.n8 a_n1598_n3888# 0.053167f
C50 plus.n9 a_n1598_n3888# 0.019768f
C51 plus.n10 a_n1598_n3888# 0.25926f
C52 plus.n11 a_n1598_n3888# 0.021899f
C53 plus.n12 a_n1598_n3888# 0.25926f
C54 plus.t6 a_n1598_n3888# 0.684182f
C55 plus.n13 a_n1598_n3888# 0.276043f
C56 plus.n14 a_n1598_n3888# 0.673353f
C57 plus.n15 a_n1598_n3888# 0.053167f
C58 plus.t10 a_n1598_n3888# 0.684182f
C59 plus.t3 a_n1598_n3888# 0.674969f
C60 plus.t9 a_n1598_n3888# 0.674969f
C61 plus.n16 a_n1598_n3888# 0.019768f
C62 plus.t0 a_n1598_n3888# 0.684182f
C63 plus.n17 a_n1598_n3888# 0.276122f
C64 plus.t1 a_n1598_n3888# 0.674969f
C65 plus.n18 a_n1598_n3888# 0.25926f
C66 plus.t7 a_n1598_n3888# 0.674969f
C67 plus.n19 a_n1598_n3888# 0.25926f
C68 plus.n20 a_n1598_n3888# 0.021899f
C69 plus.n21 a_n1598_n3888# 0.121006f
C70 plus.n22 a_n1598_n3888# 0.053167f
C71 plus.n23 a_n1598_n3888# 0.053167f
C72 plus.n24 a_n1598_n3888# 0.019768f
C73 plus.n25 a_n1598_n3888# 0.25926f
C74 plus.n26 a_n1598_n3888# 0.021899f
C75 plus.n27 a_n1598_n3888# 0.25926f
C76 plus.n28 a_n1598_n3888# 0.276043f
C77 plus.n29 a_n1598_n3888# 1.6269f
C78 source.t3 a_n1598_n3888# 3.50922f
C79 source.n0 a_n1598_n3888# 1.6254f
C80 source.t5 a_n1598_n3888# 0.313139f
C81 source.t1 a_n1598_n3888# 0.313139f
C82 source.n1 a_n1598_n3888# 2.75066f
C83 source.n2 a_n1598_n3888# 0.352677f
C84 source.t2 a_n1598_n3888# 0.313139f
C85 source.t10 a_n1598_n3888# 0.313139f
C86 source.n3 a_n1598_n3888# 2.75066f
C87 source.n4 a_n1598_n3888# 0.352677f
C88 source.t8 a_n1598_n3888# 3.50923f
C89 source.n5 a_n1598_n3888# 0.441887f
C90 source.t17 a_n1598_n3888# 3.50923f
C91 source.n6 a_n1598_n3888# 0.441887f
C92 source.t22 a_n1598_n3888# 0.313139f
C93 source.t13 a_n1598_n3888# 0.313139f
C94 source.n7 a_n1598_n3888# 2.75066f
C95 source.n8 a_n1598_n3888# 0.352677f
C96 source.t16 a_n1598_n3888# 0.313139f
C97 source.t19 a_n1598_n3888# 0.313139f
C98 source.n9 a_n1598_n3888# 2.75066f
C99 source.n10 a_n1598_n3888# 0.352677f
C100 source.t23 a_n1598_n3888# 3.50923f
C101 source.n11 a_n1598_n3888# 2.06462f
C102 source.t6 a_n1598_n3888# 3.50922f
C103 source.n12 a_n1598_n3888# 2.06462f
C104 source.t11 a_n1598_n3888# 0.313139f
C105 source.t4 a_n1598_n3888# 0.313139f
C106 source.n13 a_n1598_n3888# 2.75066f
C107 source.n14 a_n1598_n3888# 0.35268f
C108 source.t0 a_n1598_n3888# 0.313139f
C109 source.t7 a_n1598_n3888# 0.313139f
C110 source.n15 a_n1598_n3888# 2.75066f
C111 source.n16 a_n1598_n3888# 0.35268f
C112 source.t9 a_n1598_n3888# 3.50922f
C113 source.n17 a_n1598_n3888# 0.441891f
C114 source.t20 a_n1598_n3888# 3.50922f
C115 source.n18 a_n1598_n3888# 0.441891f
C116 source.t14 a_n1598_n3888# 0.313139f
C117 source.t21 a_n1598_n3888# 0.313139f
C118 source.n19 a_n1598_n3888# 2.75066f
C119 source.n20 a_n1598_n3888# 0.35268f
C120 source.t15 a_n1598_n3888# 0.313139f
C121 source.t18 a_n1598_n3888# 0.313139f
C122 source.n21 a_n1598_n3888# 2.75066f
C123 source.n22 a_n1598_n3888# 0.35268f
C124 source.t12 a_n1598_n3888# 3.50922f
C125 source.n23 a_n1598_n3888# 0.591018f
C126 source.n24 a_n1598_n3888# 1.93161f
C127 drain_right.t0 a_n1598_n3888# 0.400801f
C128 drain_right.t5 a_n1598_n3888# 0.400801f
C129 drain_right.n0 a_n1598_n3888# 3.62599f
C130 drain_right.t2 a_n1598_n3888# 0.400801f
C131 drain_right.t6 a_n1598_n3888# 0.400801f
C132 drain_right.n1 a_n1598_n3888# 3.62277f
C133 drain_right.t3 a_n1598_n3888# 0.400801f
C134 drain_right.t4 a_n1598_n3888# 0.400801f
C135 drain_right.n2 a_n1598_n3888# 3.62599f
C136 drain_right.n3 a_n1598_n3888# 2.88172f
C137 drain_right.t11 a_n1598_n3888# 0.400801f
C138 drain_right.t1 a_n1598_n3888# 0.400801f
C139 drain_right.n4 a_n1598_n3888# 3.62638f
C140 drain_right.t10 a_n1598_n3888# 0.400801f
C141 drain_right.t7 a_n1598_n3888# 0.400801f
C142 drain_right.n5 a_n1598_n3888# 3.62278f
C143 drain_right.n6 a_n1598_n3888# 0.8006f
C144 drain_right.t8 a_n1598_n3888# 0.400801f
C145 drain_right.t9 a_n1598_n3888# 0.400801f
C146 drain_right.n7 a_n1598_n3888# 3.62278f
C147 drain_right.n8 a_n1598_n3888# 0.676738f
C148 minus.n0 a_n1598_n3888# 0.052511f
C149 minus.t0 a_n1598_n3888# 0.675735f
C150 minus.t7 a_n1598_n3888# 0.666636f
C151 minus.t4 a_n1598_n3888# 0.666636f
C152 minus.n1 a_n1598_n3888# 0.019524f
C153 minus.t6 a_n1598_n3888# 0.675735f
C154 minus.n2 a_n1598_n3888# 0.272713f
C155 minus.t1 a_n1598_n3888# 0.666636f
C156 minus.n3 a_n1598_n3888# 0.256059f
C157 minus.t10 a_n1598_n3888# 0.666636f
C158 minus.n4 a_n1598_n3888# 0.256059f
C159 minus.n5 a_n1598_n3888# 0.021628f
C160 minus.n6 a_n1598_n3888# 0.119512f
C161 minus.n7 a_n1598_n3888# 0.052511f
C162 minus.n8 a_n1598_n3888# 0.052511f
C163 minus.n9 a_n1598_n3888# 0.019524f
C164 minus.n10 a_n1598_n3888# 0.256059f
C165 minus.n11 a_n1598_n3888# 0.021628f
C166 minus.n12 a_n1598_n3888# 0.256059f
C167 minus.n13 a_n1598_n3888# 0.272634f
C168 minus.n14 a_n1598_n3888# 1.9579f
C169 minus.n15 a_n1598_n3888# 0.052511f
C170 minus.t5 a_n1598_n3888# 0.666636f
C171 minus.t8 a_n1598_n3888# 0.666636f
C172 minus.n16 a_n1598_n3888# 0.019524f
C173 minus.t3 a_n1598_n3888# 0.675735f
C174 minus.n17 a_n1598_n3888# 0.272713f
C175 minus.t9 a_n1598_n3888# 0.666636f
C176 minus.n18 a_n1598_n3888# 0.256059f
C177 minus.t2 a_n1598_n3888# 0.666636f
C178 minus.n19 a_n1598_n3888# 0.256059f
C179 minus.n20 a_n1598_n3888# 0.021628f
C180 minus.n21 a_n1598_n3888# 0.119512f
C181 minus.n22 a_n1598_n3888# 0.052511f
C182 minus.n23 a_n1598_n3888# 0.052511f
C183 minus.n24 a_n1598_n3888# 0.019524f
C184 minus.n25 a_n1598_n3888# 0.256059f
C185 minus.n26 a_n1598_n3888# 0.021628f
C186 minus.n27 a_n1598_n3888# 0.256059f
C187 minus.t11 a_n1598_n3888# 0.675735f
C188 minus.n28 a_n1598_n3888# 0.272634f
C189 minus.n29 a_n1598_n3888# 0.34477f
C190 minus.n30 a_n1598_n3888# 2.36896f
.ends

