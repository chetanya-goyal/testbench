* NGSPICE file created from diffpair87.ext - technology: sky130A

.subckt diffpair87 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t21 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 source.t10 minus.t0 drain_right.t15 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 source.t0 minus.t1 drain_right.t14 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 source.t27 plus.t1 drain_left.t14 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 drain_left.t13 plus.t2 source.t25 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X5 source.t30 plus.t3 drain_left.t12 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X6 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X7 drain_right.t13 minus.t2 source.t13 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X8 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X9 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X10 drain_left.t11 plus.t4 source.t28 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 source.t2 minus.t3 drain_right.t12 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X12 source.t7 minus.t4 drain_right.t11 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 drain_right.t10 minus.t5 source.t3 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X14 drain_right.t9 minus.t6 source.t5 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 source.t19 plus.t5 drain_left.t10 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 source.t14 minus.t7 drain_right.t8 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_right.t7 minus.t8 source.t6 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X18 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X19 drain_right.t6 minus.t9 source.t8 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X20 source.t26 plus.t6 drain_left.t9 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X21 drain_left.t8 plus.t7 source.t22 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X22 source.t23 plus.t8 drain_left.t7 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_right.t5 minus.t10 source.t11 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X24 drain_right.t4 minus.t11 source.t4 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X25 source.t1 minus.t12 drain_right.t3 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X26 source.t15 minus.t13 drain_right.t2 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X27 drain_left.t6 plus.t9 source.t17 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X28 source.t9 minus.t14 drain_right.t1 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X29 drain_left.t5 plus.t10 source.t24 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X30 source.t29 plus.t11 drain_left.t4 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X31 source.t31 plus.t12 drain_left.t3 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X32 drain_right.t0 minus.t15 source.t12 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X33 drain_left.t2 plus.t13 source.t20 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X34 drain_left.t1 plus.t14 source.t18 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X35 source.t16 plus.t15 drain_left.t0 a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 plus.n5 plus.t8 570.367
R1 plus.n21 plus.t7 570.367
R2 plus.n28 plus.t10 570.367
R3 plus.n44 plus.t3 570.367
R4 plus.n6 plus.t14 530.201
R5 plus.n3 plus.t12 530.201
R6 plus.n12 plus.t9 530.201
R7 plus.n14 plus.t15 530.201
R8 plus.n1 plus.t13 530.201
R9 plus.n20 plus.t11 530.201
R10 plus.n29 plus.t6 530.201
R11 plus.n26 plus.t2 530.201
R12 plus.n35 plus.t1 530.201
R13 plus.n37 plus.t0 530.201
R14 plus.n24 plus.t5 530.201
R15 plus.n43 plus.t4 530.201
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 69.3793
R39 plus.n15 plus.n1 69.3793
R40 plus.n38 plus.n24 69.3793
R41 plus.n34 plus.n26 69.3793
R42 plus.n6 plus.n5 54.7732
R43 plus.n21 plus.n20 54.7732
R44 plus.n44 plus.n43 54.7732
R45 plus.n29 plus.n28 54.7732
R46 plus.n13 plus.n12 47.4702
R47 plus.n14 plus.n13 47.4702
R48 plus.n37 plus.n36 47.4702
R49 plus.n36 plus.n35 47.4702
R50 plus plus.n45 26.3627
R51 plus.n12 plus.n11 25.5611
R52 plus.n15 plus.n14 25.5611
R53 plus.n38 plus.n37 25.5611
R54 plus.n35 plus.n34 25.5611
R55 plus.n7 plus.n6 18.2581
R56 plus.n20 plus.n19 18.2581
R57 plus.n43 plus.n42 18.2581
R58 plus.n30 plus.n29 18.2581
R59 plus plus.n22 8.36035
R60 plus.n8 plus.n3 3.65202
R61 plus.n18 plus.n1 3.65202
R62 plus.n41 plus.n24 3.65202
R63 plus.n31 plus.n26 3.65202
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 source.n0 source.t22 99.1169
R79 source.n7 source.t23 99.1169
R80 source.n8 source.t3 99.1169
R81 source.n15 source.t1 99.1169
R82 source.n31 source.t6 99.1168
R83 source.n24 source.t0 99.1168
R84 source.n23 source.t24 99.1168
R85 source.n16 source.t30 99.1168
R86 source.n2 source.n1 84.1169
R87 source.n4 source.n3 84.1169
R88 source.n6 source.n5 84.1169
R89 source.n10 source.n9 84.1169
R90 source.n12 source.n11 84.1169
R91 source.n14 source.n13 84.1169
R92 source.n30 source.n29 84.1168
R93 source.n28 source.n27 84.1168
R94 source.n26 source.n25 84.1168
R95 source.n22 source.n21 84.1168
R96 source.n20 source.n19 84.1168
R97 source.n18 source.n17 84.1168
R98 source.n29 source.t12 15.0005
R99 source.n29 source.t15 15.0005
R100 source.n27 source.t13 15.0005
R101 source.n27 source.t10 15.0005
R102 source.n25 source.t8 15.0005
R103 source.n25 source.t7 15.0005
R104 source.n21 source.t25 15.0005
R105 source.n21 source.t26 15.0005
R106 source.n19 source.t21 15.0005
R107 source.n19 source.t27 15.0005
R108 source.n17 source.t28 15.0005
R109 source.n17 source.t19 15.0005
R110 source.n1 source.t20 15.0005
R111 source.n1 source.t29 15.0005
R112 source.n3 source.t17 15.0005
R113 source.n3 source.t16 15.0005
R114 source.n5 source.t18 15.0005
R115 source.n5 source.t31 15.0005
R116 source.n9 source.t11 15.0005
R117 source.n9 source.t2 15.0005
R118 source.n11 source.t5 15.0005
R119 source.n11 source.t14 15.0005
R120 source.n13 source.t4 15.0005
R121 source.n13 source.t9 15.0005
R122 source.n16 source.n15 14.2723
R123 source.n32 source.n0 8.72921
R124 source.n32 source.n31 5.5436
R125 source.n15 source.n14 0.560845
R126 source.n14 source.n12 0.560845
R127 source.n12 source.n10 0.560845
R128 source.n10 source.n8 0.560845
R129 source.n7 source.n6 0.560845
R130 source.n6 source.n4 0.560845
R131 source.n4 source.n2 0.560845
R132 source.n2 source.n0 0.560845
R133 source.n18 source.n16 0.560845
R134 source.n20 source.n18 0.560845
R135 source.n22 source.n20 0.560845
R136 source.n23 source.n22 0.560845
R137 source.n26 source.n24 0.560845
R138 source.n28 source.n26 0.560845
R139 source.n30 source.n28 0.560845
R140 source.n31 source.n30 0.560845
R141 source.n8 source.n7 0.470328
R142 source.n24 source.n23 0.470328
R143 source source.n32 0.188
R144 drain_left.n9 drain_left.n7 101.356
R145 drain_left.n5 drain_left.n3 101.356
R146 drain_left.n2 drain_left.n0 101.356
R147 drain_left.n13 drain_left.n12 100.796
R148 drain_left.n11 drain_left.n10 100.796
R149 drain_left.n9 drain_left.n8 100.796
R150 drain_left.n5 drain_left.n4 100.796
R151 drain_left.n2 drain_left.n1 100.796
R152 drain_left drain_left.n6 23.4336
R153 drain_left.n3 drain_left.t9 15.0005
R154 drain_left.n3 drain_left.t5 15.0005
R155 drain_left.n4 drain_left.t14 15.0005
R156 drain_left.n4 drain_left.t13 15.0005
R157 drain_left.n1 drain_left.t10 15.0005
R158 drain_left.n1 drain_left.t15 15.0005
R159 drain_left.n0 drain_left.t12 15.0005
R160 drain_left.n0 drain_left.t11 15.0005
R161 drain_left.n12 drain_left.t4 15.0005
R162 drain_left.n12 drain_left.t8 15.0005
R163 drain_left.n10 drain_left.t0 15.0005
R164 drain_left.n10 drain_left.t2 15.0005
R165 drain_left.n8 drain_left.t3 15.0005
R166 drain_left.n8 drain_left.t6 15.0005
R167 drain_left.n7 drain_left.t7 15.0005
R168 drain_left.n7 drain_left.t1 15.0005
R169 drain_left drain_left.n13 6.21356
R170 drain_left.n11 drain_left.n9 0.560845
R171 drain_left.n13 drain_left.n11 0.560845
R172 drain_left.n6 drain_left.n5 0.225326
R173 drain_left.n6 drain_left.n2 0.225326
R174 minus.n21 minus.t12 570.367
R175 minus.n5 minus.t5 570.367
R176 minus.n44 minus.t8 570.367
R177 minus.n28 minus.t1 570.367
R178 minus.n20 minus.t11 530.201
R179 minus.n1 minus.t14 530.201
R180 minus.n14 minus.t6 530.201
R181 minus.n12 minus.t7 530.201
R182 minus.n3 minus.t10 530.201
R183 minus.n6 minus.t3 530.201
R184 minus.n43 minus.t13 530.201
R185 minus.n24 minus.t15 530.201
R186 minus.n37 minus.t0 530.201
R187 minus.n35 minus.t2 530.201
R188 minus.n26 minus.t4 530.201
R189 minus.n29 minus.t9 530.201
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 69.3793
R213 minus.n11 minus.n3 69.3793
R214 minus.n34 minus.n26 69.3793
R215 minus.n38 minus.n24 69.3793
R216 minus.n21 minus.n20 54.7732
R217 minus.n6 minus.n5 54.7732
R218 minus.n29 minus.n28 54.7732
R219 minus.n44 minus.n43 54.7732
R220 minus.n14 minus.n13 47.4702
R221 minus.n13 minus.n12 47.4702
R222 minus.n36 minus.n35 47.4702
R223 minus.n37 minus.n36 47.4702
R224 minus.n46 minus.n22 28.6937
R225 minus.n15 minus.n14 25.5611
R226 minus.n12 minus.n11 25.5611
R227 minus.n35 minus.n34 25.5611
R228 minus.n38 minus.n37 25.5611
R229 minus.n20 minus.n19 18.2581
R230 minus.n7 minus.n6 18.2581
R231 minus.n30 minus.n29 18.2581
R232 minus.n43 minus.n42 18.2581
R233 minus.n46 minus.n45 6.50429
R234 minus.n18 minus.n1 3.65202
R235 minus.n8 minus.n3 3.65202
R236 minus.n31 minus.n26 3.65202
R237 minus.n41 minus.n24 3.65202
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 101.356
R254 drain_right.n5 drain_right.n3 101.356
R255 drain_right.n2 drain_right.n0 101.356
R256 drain_right.n9 drain_right.n8 100.796
R257 drain_right.n11 drain_right.n10 100.796
R258 drain_right.n13 drain_right.n12 100.796
R259 drain_right.n5 drain_right.n4 100.796
R260 drain_right.n2 drain_right.n1 100.796
R261 drain_right drain_right.n6 22.8803
R262 drain_right.n3 drain_right.t2 15.0005
R263 drain_right.n3 drain_right.t7 15.0005
R264 drain_right.n4 drain_right.t15 15.0005
R265 drain_right.n4 drain_right.t0 15.0005
R266 drain_right.n1 drain_right.t11 15.0005
R267 drain_right.n1 drain_right.t13 15.0005
R268 drain_right.n0 drain_right.t14 15.0005
R269 drain_right.n0 drain_right.t6 15.0005
R270 drain_right.n7 drain_right.t12 15.0005
R271 drain_right.n7 drain_right.t10 15.0005
R272 drain_right.n8 drain_right.t8 15.0005
R273 drain_right.n8 drain_right.t5 15.0005
R274 drain_right.n10 drain_right.t1 15.0005
R275 drain_right.n10 drain_right.t9 15.0005
R276 drain_right.n12 drain_right.t3 15.0005
R277 drain_right.n12 drain_right.t4 15.0005
R278 drain_right drain_right.n13 6.21356
R279 drain_right.n13 drain_right.n11 0.560845
R280 drain_right.n11 drain_right.n9 0.560845
R281 drain_right.n6 drain_right.n5 0.225326
R282 drain_right.n6 drain_right.n2 0.225326
C0 drain_left minus 0.177f
C1 drain_right source 7.58582f
C2 plus source 1.13446f
C3 minus source 1.1205f
C4 drain_right plus 0.344074f
C5 drain_left source 7.585471f
C6 drain_right minus 1.01594f
C7 drain_right drain_left 0.96779f
C8 plus minus 3.64866f
C9 plus drain_left 1.1995f
C10 drain_right a_n1886_n1288# 3.8982f
C11 drain_left a_n1886_n1288# 4.15351f
C12 source a_n1886_n1288# 3.210594f
C13 minus a_n1886_n1288# 6.167137f
C14 plus a_n1886_n1288# 6.92527f
C15 drain_right.t14 a_n1886_n1288# 0.058741f
C16 drain_right.t6 a_n1886_n1288# 0.058741f
C17 drain_right.n0 a_n1886_n1288# 0.285087f
C18 drain_right.t11 a_n1886_n1288# 0.058741f
C19 drain_right.t13 a_n1886_n1288# 0.058741f
C20 drain_right.n1 a_n1886_n1288# 0.283505f
C21 drain_right.n2 a_n1886_n1288# 0.536978f
C22 drain_right.t2 a_n1886_n1288# 0.058741f
C23 drain_right.t7 a_n1886_n1288# 0.058741f
C24 drain_right.n3 a_n1886_n1288# 0.285087f
C25 drain_right.t15 a_n1886_n1288# 0.058741f
C26 drain_right.t0 a_n1886_n1288# 0.058741f
C27 drain_right.n4 a_n1886_n1288# 0.283505f
C28 drain_right.n5 a_n1886_n1288# 0.536978f
C29 drain_right.n6 a_n1886_n1288# 0.662748f
C30 drain_right.t12 a_n1886_n1288# 0.058741f
C31 drain_right.t10 a_n1886_n1288# 0.058741f
C32 drain_right.n7 a_n1886_n1288# 0.285088f
C33 drain_right.t8 a_n1886_n1288# 0.058741f
C34 drain_right.t5 a_n1886_n1288# 0.058741f
C35 drain_right.n8 a_n1886_n1288# 0.283506f
C36 drain_right.n9 a_n1886_n1288# 0.560967f
C37 drain_right.t1 a_n1886_n1288# 0.058741f
C38 drain_right.t9 a_n1886_n1288# 0.058741f
C39 drain_right.n10 a_n1886_n1288# 0.283506f
C40 drain_right.n11 a_n1886_n1288# 0.276334f
C41 drain_right.t3 a_n1886_n1288# 0.058741f
C42 drain_right.t4 a_n1886_n1288# 0.058741f
C43 drain_right.n12 a_n1886_n1288# 0.283506f
C44 drain_right.n13 a_n1886_n1288# 0.481189f
C45 minus.n0 a_n1886_n1288# 0.032477f
C46 minus.t12 a_n1886_n1288# 0.030327f
C47 minus.t11 a_n1886_n1288# 0.02867f
C48 minus.t14 a_n1886_n1288# 0.02867f
C49 minus.n1 a_n1886_n1288# 0.02503f
C50 minus.n2 a_n1886_n1288# 0.032477f
C51 minus.t6 a_n1886_n1288# 0.02867f
C52 minus.t7 a_n1886_n1288# 0.02867f
C53 minus.t10 a_n1886_n1288# 0.02867f
C54 minus.n3 a_n1886_n1288# 0.02503f
C55 minus.n4 a_n1886_n1288# 0.068917f
C56 minus.t3 a_n1886_n1288# 0.02867f
C57 minus.t5 a_n1886_n1288# 0.030327f
C58 minus.n5 a_n1886_n1288# 0.035691f
C59 minus.n6 a_n1886_n1288# 0.02503f
C60 minus.n7 a_n1886_n1288# 0.013277f
C61 minus.n8 a_n1886_n1288# 0.011274f
C62 minus.n9 a_n1886_n1288# 0.032477f
C63 minus.n10 a_n1886_n1288# 0.032477f
C64 minus.n11 a_n1886_n1288# 0.013777f
C65 minus.n12 a_n1886_n1288# 0.02503f
C66 minus.n13 a_n1886_n1288# 0.013777f
C67 minus.n14 a_n1886_n1288# 0.02503f
C68 minus.n15 a_n1886_n1288# 0.013777f
C69 minus.n16 a_n1886_n1288# 0.032477f
C70 minus.n17 a_n1886_n1288# 0.032477f
C71 minus.n18 a_n1886_n1288# 0.011274f
C72 minus.n19 a_n1886_n1288# 0.013277f
C73 minus.n20 a_n1886_n1288# 0.02503f
C74 minus.n21 a_n1886_n1288# 0.035648f
C75 minus.n22 a_n1886_n1288# 0.782475f
C76 minus.n23 a_n1886_n1288# 0.032477f
C77 minus.t13 a_n1886_n1288# 0.02867f
C78 minus.t15 a_n1886_n1288# 0.02867f
C79 minus.n24 a_n1886_n1288# 0.02503f
C80 minus.n25 a_n1886_n1288# 0.032477f
C81 minus.t0 a_n1886_n1288# 0.02867f
C82 minus.t2 a_n1886_n1288# 0.02867f
C83 minus.t4 a_n1886_n1288# 0.02867f
C84 minus.n26 a_n1886_n1288# 0.02503f
C85 minus.n27 a_n1886_n1288# 0.068917f
C86 minus.t9 a_n1886_n1288# 0.02867f
C87 minus.t1 a_n1886_n1288# 0.030327f
C88 minus.n28 a_n1886_n1288# 0.035691f
C89 minus.n29 a_n1886_n1288# 0.02503f
C90 minus.n30 a_n1886_n1288# 0.013277f
C91 minus.n31 a_n1886_n1288# 0.011274f
C92 minus.n32 a_n1886_n1288# 0.032477f
C93 minus.n33 a_n1886_n1288# 0.032477f
C94 minus.n34 a_n1886_n1288# 0.013777f
C95 minus.n35 a_n1886_n1288# 0.02503f
C96 minus.n36 a_n1886_n1288# 0.013777f
C97 minus.n37 a_n1886_n1288# 0.02503f
C98 minus.n38 a_n1886_n1288# 0.013777f
C99 minus.n39 a_n1886_n1288# 0.032477f
C100 minus.n40 a_n1886_n1288# 0.032477f
C101 minus.n41 a_n1886_n1288# 0.011274f
C102 minus.n42 a_n1886_n1288# 0.013277f
C103 minus.n43 a_n1886_n1288# 0.02503f
C104 minus.t8 a_n1886_n1288# 0.030327f
C105 minus.n44 a_n1886_n1288# 0.035648f
C106 minus.n45 a_n1886_n1288# 0.212657f
C107 minus.n46 a_n1886_n1288# 0.966721f
C108 drain_left.t12 a_n1886_n1288# 0.058009f
C109 drain_left.t11 a_n1886_n1288# 0.058009f
C110 drain_left.n0 a_n1886_n1288# 0.281532f
C111 drain_left.t10 a_n1886_n1288# 0.058009f
C112 drain_left.t15 a_n1886_n1288# 0.058009f
C113 drain_left.n1 a_n1886_n1288# 0.27997f
C114 drain_left.n2 a_n1886_n1288# 0.530283f
C115 drain_left.t9 a_n1886_n1288# 0.058009f
C116 drain_left.t5 a_n1886_n1288# 0.058009f
C117 drain_left.n3 a_n1886_n1288# 0.281532f
C118 drain_left.t14 a_n1886_n1288# 0.058009f
C119 drain_left.t13 a_n1886_n1288# 0.058009f
C120 drain_left.n4 a_n1886_n1288# 0.27997f
C121 drain_left.n5 a_n1886_n1288# 0.530283f
C122 drain_left.n6 a_n1886_n1288# 0.70192f
C123 drain_left.t7 a_n1886_n1288# 0.058009f
C124 drain_left.t1 a_n1886_n1288# 0.058009f
C125 drain_left.n7 a_n1886_n1288# 0.281533f
C126 drain_left.t3 a_n1886_n1288# 0.058009f
C127 drain_left.t6 a_n1886_n1288# 0.058009f
C128 drain_left.n8 a_n1886_n1288# 0.279971f
C129 drain_left.n9 a_n1886_n1288# 0.553972f
C130 drain_left.t0 a_n1886_n1288# 0.058009f
C131 drain_left.t2 a_n1886_n1288# 0.058009f
C132 drain_left.n10 a_n1886_n1288# 0.279971f
C133 drain_left.n11 a_n1886_n1288# 0.272889f
C134 drain_left.t4 a_n1886_n1288# 0.058009f
C135 drain_left.t8 a_n1886_n1288# 0.058009f
C136 drain_left.n12 a_n1886_n1288# 0.279971f
C137 drain_left.n13 a_n1886_n1288# 0.475189f
C138 source.t22 a_n1886_n1288# 0.317012f
C139 source.n0 a_n1886_n1288# 0.604216f
C140 source.t20 a_n1886_n1288# 0.060379f
C141 source.t29 a_n1886_n1288# 0.060379f
C142 source.n1 a_n1886_n1288# 0.254094f
C143 source.n2 a_n1886_n1288# 0.287079f
C144 source.t17 a_n1886_n1288# 0.060379f
C145 source.t16 a_n1886_n1288# 0.060379f
C146 source.n3 a_n1886_n1288# 0.254094f
C147 source.n4 a_n1886_n1288# 0.287079f
C148 source.t18 a_n1886_n1288# 0.060379f
C149 source.t31 a_n1886_n1288# 0.060379f
C150 source.n5 a_n1886_n1288# 0.254094f
C151 source.n6 a_n1886_n1288# 0.287079f
C152 source.t23 a_n1886_n1288# 0.317012f
C153 source.n7 a_n1886_n1288# 0.325489f
C154 source.t3 a_n1886_n1288# 0.317012f
C155 source.n8 a_n1886_n1288# 0.325489f
C156 source.t11 a_n1886_n1288# 0.060379f
C157 source.t2 a_n1886_n1288# 0.060379f
C158 source.n9 a_n1886_n1288# 0.254094f
C159 source.n10 a_n1886_n1288# 0.287079f
C160 source.t5 a_n1886_n1288# 0.060379f
C161 source.t14 a_n1886_n1288# 0.060379f
C162 source.n11 a_n1886_n1288# 0.254094f
C163 source.n12 a_n1886_n1288# 0.287079f
C164 source.t4 a_n1886_n1288# 0.060379f
C165 source.t9 a_n1886_n1288# 0.060379f
C166 source.n13 a_n1886_n1288# 0.254094f
C167 source.n14 a_n1886_n1288# 0.287079f
C168 source.t1 a_n1886_n1288# 0.317012f
C169 source.n15 a_n1886_n1288# 0.839601f
C170 source.t30 a_n1886_n1288# 0.317011f
C171 source.n16 a_n1886_n1288# 0.839602f
C172 source.t28 a_n1886_n1288# 0.060379f
C173 source.t19 a_n1886_n1288# 0.060379f
C174 source.n17 a_n1886_n1288# 0.254093f
C175 source.n18 a_n1886_n1288# 0.287081f
C176 source.t21 a_n1886_n1288# 0.060379f
C177 source.t27 a_n1886_n1288# 0.060379f
C178 source.n19 a_n1886_n1288# 0.254093f
C179 source.n20 a_n1886_n1288# 0.287081f
C180 source.t25 a_n1886_n1288# 0.060379f
C181 source.t26 a_n1886_n1288# 0.060379f
C182 source.n21 a_n1886_n1288# 0.254093f
C183 source.n22 a_n1886_n1288# 0.287081f
C184 source.t24 a_n1886_n1288# 0.317011f
C185 source.n23 a_n1886_n1288# 0.32549f
C186 source.t0 a_n1886_n1288# 0.317011f
C187 source.n24 a_n1886_n1288# 0.32549f
C188 source.t8 a_n1886_n1288# 0.060379f
C189 source.t7 a_n1886_n1288# 0.060379f
C190 source.n25 a_n1886_n1288# 0.254093f
C191 source.n26 a_n1886_n1288# 0.287081f
C192 source.t13 a_n1886_n1288# 0.060379f
C193 source.t10 a_n1886_n1288# 0.060379f
C194 source.n27 a_n1886_n1288# 0.254093f
C195 source.n28 a_n1886_n1288# 0.287081f
C196 source.t12 a_n1886_n1288# 0.060379f
C197 source.t15 a_n1886_n1288# 0.060379f
C198 source.n29 a_n1886_n1288# 0.254093f
C199 source.n30 a_n1886_n1288# 0.287081f
C200 source.t6 a_n1886_n1288# 0.317011f
C201 source.n31 a_n1886_n1288# 0.468943f
C202 source.n32 a_n1886_n1288# 0.623978f
C203 plus.n0 a_n1886_n1288# 0.033081f
C204 plus.t11 a_n1886_n1288# 0.029203f
C205 plus.t13 a_n1886_n1288# 0.029203f
C206 plus.n1 a_n1886_n1288# 0.025495f
C207 plus.n2 a_n1886_n1288# 0.033081f
C208 plus.t15 a_n1886_n1288# 0.029203f
C209 plus.t9 a_n1886_n1288# 0.029203f
C210 plus.t12 a_n1886_n1288# 0.029203f
C211 plus.n3 a_n1886_n1288# 0.025495f
C212 plus.n4 a_n1886_n1288# 0.070198f
C213 plus.t14 a_n1886_n1288# 0.029203f
C214 plus.t8 a_n1886_n1288# 0.030891f
C215 plus.n5 a_n1886_n1288# 0.036354f
C216 plus.n6 a_n1886_n1288# 0.025495f
C217 plus.n7 a_n1886_n1288# 0.013524f
C218 plus.n8 a_n1886_n1288# 0.011484f
C219 plus.n9 a_n1886_n1288# 0.033081f
C220 plus.n10 a_n1886_n1288# 0.033081f
C221 plus.n11 a_n1886_n1288# 0.014033f
C222 plus.n12 a_n1886_n1288# 0.025495f
C223 plus.n13 a_n1886_n1288# 0.014033f
C224 plus.n14 a_n1886_n1288# 0.025495f
C225 plus.n15 a_n1886_n1288# 0.014033f
C226 plus.n16 a_n1886_n1288# 0.033081f
C227 plus.n17 a_n1886_n1288# 0.033081f
C228 plus.n18 a_n1886_n1288# 0.011484f
C229 plus.n19 a_n1886_n1288# 0.013524f
C230 plus.n20 a_n1886_n1288# 0.025495f
C231 plus.t7 a_n1886_n1288# 0.030891f
C232 plus.n21 a_n1886_n1288# 0.036311f
C233 plus.n22 a_n1886_n1288# 0.236845f
C234 plus.n23 a_n1886_n1288# 0.033081f
C235 plus.t3 a_n1886_n1288# 0.030891f
C236 plus.t4 a_n1886_n1288# 0.029203f
C237 plus.t5 a_n1886_n1288# 0.029203f
C238 plus.n24 a_n1886_n1288# 0.025495f
C239 plus.n25 a_n1886_n1288# 0.033081f
C240 plus.t0 a_n1886_n1288# 0.029203f
C241 plus.t1 a_n1886_n1288# 0.029203f
C242 plus.t2 a_n1886_n1288# 0.029203f
C243 plus.n26 a_n1886_n1288# 0.025495f
C244 plus.n27 a_n1886_n1288# 0.070198f
C245 plus.t6 a_n1886_n1288# 0.029203f
C246 plus.t10 a_n1886_n1288# 0.030891f
C247 plus.n28 a_n1886_n1288# 0.036354f
C248 plus.n29 a_n1886_n1288# 0.025495f
C249 plus.n30 a_n1886_n1288# 0.013524f
C250 plus.n31 a_n1886_n1288# 0.011484f
C251 plus.n32 a_n1886_n1288# 0.033081f
C252 plus.n33 a_n1886_n1288# 0.033081f
C253 plus.n34 a_n1886_n1288# 0.014033f
C254 plus.n35 a_n1886_n1288# 0.025495f
C255 plus.n36 a_n1886_n1288# 0.014033f
C256 plus.n37 a_n1886_n1288# 0.025495f
C257 plus.n38 a_n1886_n1288# 0.014033f
C258 plus.n39 a_n1886_n1288# 0.033081f
C259 plus.n40 a_n1886_n1288# 0.033081f
C260 plus.n41 a_n1886_n1288# 0.011484f
C261 plus.n42 a_n1886_n1288# 0.013524f
C262 plus.n43 a_n1886_n1288# 0.025495f
C263 plus.n44 a_n1886_n1288# 0.036311f
C264 plus.n45 a_n1886_n1288# 0.76069f
.ends

