* NGSPICE file created from diffpair610.ext - technology: sky130A

.subckt diffpair610 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t3 a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.6
X1 drain_left.t1 plus.t0 source.t1 a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.6
X2 drain_right.t0 minus.t1 source.t2 a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.6
X3 drain_left.t0 plus.t1 source.t0 a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.6
X4 a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X5 a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X6 a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X7 a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# a_n1088_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
R0 minus.n0 minus.t0 1069.48
R1 minus.n0 minus.t1 1036.66
R2 minus minus.n0 0.188
R3 source.n0 source.t1 44.1297
R4 source.n1 source.t3 44.1296
R5 source.n3 source.t2 44.1295
R6 source.n2 source.t0 44.1295
R7 source.n2 source.n1 28.9669
R8 source.n4 source.n0 22.5014
R9 source.n4 source.n3 5.66429
R10 source.n1 source.n0 0.87119
R11 source.n3 source.n2 0.87119
R12 source source.n4 0.188
R13 drain_right drain_right.t0 94.8446
R14 drain_right drain_right.t1 66.862
R15 plus plus.t1 1060.33
R16 plus plus.t0 1045.34
R17 drain_left drain_left.t0 95.3978
R18 drain_left drain_left.t1 67.2629
C0 source plus 2.11396f
C1 drain_right source 9.153701f
C2 drain_left plus 3.09556f
C3 drain_right drain_left 0.454995f
C4 minus plus 5.97848f
C5 drain_right minus 2.99931f
C6 drain_right plus 0.258094f
C7 source drain_left 9.16801f
C8 source minus 2.09904f
C9 drain_left minus 0.171812f
C10 drain_right a_n1088_n4892# 9.02569f
C11 drain_left a_n1088_n4892# 9.191879f
C12 source a_n1088_n4892# 9.470078f
C13 minus a_n1088_n4892# 4.571388f
C14 plus a_n1088_n4892# 11.209311f
C15 drain_left.t0 a_n1088_n4892# 4.42168f
C16 drain_left.t1 a_n1088_n4892# 3.92799f
C17 plus.t0 a_n1088_n4892# 2.17394f
C18 plus.t1 a_n1088_n4892# 2.22328f
C19 drain_right.t0 a_n1088_n4892# 4.39387f
C20 drain_right.t1 a_n1088_n4892# 3.92091f
C21 source.t1 a_n1088_n4892# 3.65762f
C22 source.n0 a_n1088_n4892# 1.58801f
C23 source.t3 a_n1088_n4892# 3.65762f
C24 source.n1 a_n1088_n4892# 2.00641f
C25 source.t0 a_n1088_n4892# 3.6576f
C26 source.n2 a_n1088_n4892# 2.00643f
C27 source.t2 a_n1088_n4892# 3.6576f
C28 source.n3 a_n1088_n4892# 0.499703f
C29 source.n4 a_n1088_n4892# 1.83491f
C30 minus.t0 a_n1088_n4892# 2.21926f
C31 minus.t1 a_n1088_n4892# 2.11574f
C32 minus.n0 a_n1088_n4892# 6.72647f
.ends

