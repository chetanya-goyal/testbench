* NGSPICE file created from diffpair297.ext - technology: sky130A

.subckt diffpair297 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t13 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X1 drain_left.t10 plus.t1 source.t30 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X2 source.t29 plus.t2 drain_left.t3 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X3 drain_left.t8 plus.t3 source.t28 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X4 source.t15 minus.t0 drain_right.t15 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X5 source.t3 minus.t1 drain_right.t14 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X6 drain_right.t13 minus.t2 source.t9 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X7 drain_right.t12 minus.t3 source.t13 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X8 source.t2 minus.t4 drain_right.t11 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X9 source.t10 minus.t5 drain_right.t10 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X10 drain_left.t6 plus.t4 source.t27 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X11 drain_left.t2 plus.t5 source.t26 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X12 drain_right.t9 minus.t6 source.t0 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X13 source.t25 plus.t6 drain_left.t12 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X14 source.t14 minus.t7 drain_right.t8 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X15 drain_right.t7 minus.t8 source.t1 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X16 drain_left.t7 plus.t7 source.t24 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X17 drain_right.t6 minus.t9 source.t7 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X18 source.t23 plus.t8 drain_left.t5 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X19 source.t22 plus.t9 drain_left.t14 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X20 a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.6
X21 drain_left.t0 plus.t10 source.t21 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X22 source.t11 minus.t10 drain_right.t5 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X23 source.t20 plus.t11 drain_left.t1 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X24 drain_right.t4 minus.t11 source.t5 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X25 drain_right.t3 minus.t12 source.t6 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X26 drain_left.t15 plus.t12 source.t19 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X27 source.t18 plus.t13 drain_left.t11 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X28 a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X29 drain_left.t9 plus.t14 source.t17 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X30 source.t12 minus.t13 drain_right.t2 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X31 drain_right.t1 minus.t14 source.t4 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X32 source.t16 plus.t15 drain_left.t4 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X33 a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X34 source.t8 minus.t15 drain_right.t0 a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X35 a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# a_n2390_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
R0 plus.n6 plus.t13 327.454
R1 plus.n30 plus.t7 327.454
R2 plus.n22 plus.t1 306.473
R3 plus.n21 plus.t2 306.473
R4 plus.n1 plus.t3 306.473
R5 plus.n15 plus.t6 306.473
R6 plus.n3 plus.t10 306.473
R7 plus.n9 plus.t11 306.473
R8 plus.n5 plus.t12 306.473
R9 plus.n46 plus.t9 306.473
R10 plus.n45 plus.t5 306.473
R11 plus.n25 plus.t15 306.473
R12 plus.n39 plus.t14 306.473
R13 plus.n27 plus.t8 306.473
R14 plus.n33 plus.t4 306.473
R15 plus.n29 plus.t0 306.473
R16 plus.n8 plus.n7 161.3
R17 plus.n9 plus.n4 161.3
R18 plus.n11 plus.n10 161.3
R19 plus.n12 plus.n3 161.3
R20 plus.n14 plus.n13 161.3
R21 plus.n15 plus.n2 161.3
R22 plus.n17 plus.n16 161.3
R23 plus.n18 plus.n1 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n21 plus.n0 161.3
R26 plus.n23 plus.n22 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n33 plus.n28 161.3
R29 plus.n35 plus.n34 161.3
R30 plus.n36 plus.n27 161.3
R31 plus.n38 plus.n37 161.3
R32 plus.n39 plus.n26 161.3
R33 plus.n41 plus.n40 161.3
R34 plus.n42 plus.n25 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n45 plus.n24 161.3
R37 plus.n47 plus.n46 161.3
R38 plus.n7 plus.n6 70.4033
R39 plus.n31 plus.n30 70.4033
R40 plus.n22 plus.n21 48.2005
R41 plus.n46 plus.n45 48.2005
R42 plus.n20 plus.n1 44.549
R43 plus.n9 plus.n8 44.549
R44 plus.n44 plus.n25 44.549
R45 plus.n33 plus.n32 44.549
R46 plus.n16 plus.n15 34.3247
R47 plus.n10 plus.n3 34.3247
R48 plus.n40 plus.n39 34.3247
R49 plus.n34 plus.n27 34.3247
R50 plus plus.n47 29.9384
R51 plus.n14 plus.n3 24.1005
R52 plus.n15 plus.n14 24.1005
R53 plus.n39 plus.n38 24.1005
R54 plus.n38 plus.n27 24.1005
R55 plus.n6 plus.n5 20.9576
R56 plus.n30 plus.n29 20.9576
R57 plus.n16 plus.n1 13.8763
R58 plus.n10 plus.n9 13.8763
R59 plus.n40 plus.n25 13.8763
R60 plus.n34 plus.n33 13.8763
R61 plus plus.n23 10.027
R62 plus.n21 plus.n20 3.65202
R63 plus.n8 plus.n5 3.65202
R64 plus.n45 plus.n44 3.65202
R65 plus.n32 plus.n29 3.65202
R66 plus.n7 plus.n4 0.189894
R67 plus.n11 plus.n4 0.189894
R68 plus.n12 plus.n11 0.189894
R69 plus.n13 plus.n12 0.189894
R70 plus.n13 plus.n2 0.189894
R71 plus.n17 plus.n2 0.189894
R72 plus.n18 plus.n17 0.189894
R73 plus.n19 plus.n18 0.189894
R74 plus.n19 plus.n0 0.189894
R75 plus.n23 plus.n0 0.189894
R76 plus.n47 plus.n24 0.189894
R77 plus.n43 plus.n24 0.189894
R78 plus.n43 plus.n42 0.189894
R79 plus.n42 plus.n41 0.189894
R80 plus.n41 plus.n26 0.189894
R81 plus.n37 plus.n26 0.189894
R82 plus.n37 plus.n36 0.189894
R83 plus.n36 plus.n35 0.189894
R84 plus.n35 plus.n28 0.189894
R85 plus.n31 plus.n28 0.189894
R86 drain_left.n9 drain_left.n7 67.9925
R87 drain_left.n5 drain_left.n3 67.9924
R88 drain_left.n2 drain_left.n0 67.9924
R89 drain_left.n11 drain_left.n10 67.1908
R90 drain_left.n9 drain_left.n8 67.1908
R91 drain_left.n13 drain_left.n12 67.1907
R92 drain_left.n5 drain_left.n4 67.1907
R93 drain_left.n2 drain_left.n1 67.1907
R94 drain_left drain_left.n6 28.0328
R95 drain_left drain_left.n13 6.45494
R96 drain_left.n3 drain_left.t13 3.3005
R97 drain_left.n3 drain_left.t7 3.3005
R98 drain_left.n4 drain_left.t5 3.3005
R99 drain_left.n4 drain_left.t6 3.3005
R100 drain_left.n1 drain_left.t4 3.3005
R101 drain_left.n1 drain_left.t9 3.3005
R102 drain_left.n0 drain_left.t14 3.3005
R103 drain_left.n0 drain_left.t2 3.3005
R104 drain_left.n12 drain_left.t3 3.3005
R105 drain_left.n12 drain_left.t10 3.3005
R106 drain_left.n10 drain_left.t12 3.3005
R107 drain_left.n10 drain_left.t8 3.3005
R108 drain_left.n8 drain_left.t1 3.3005
R109 drain_left.n8 drain_left.t0 3.3005
R110 drain_left.n7 drain_left.t11 3.3005
R111 drain_left.n7 drain_left.t15 3.3005
R112 drain_left.n11 drain_left.n9 0.802224
R113 drain_left.n13 drain_left.n11 0.802224
R114 drain_left.n6 drain_left.n5 0.346016
R115 drain_left.n6 drain_left.n2 0.346016
R116 source.n274 source.n248 289.615
R117 source.n236 source.n210 289.615
R118 source.n204 source.n178 289.615
R119 source.n166 source.n140 289.615
R120 source.n26 source.n0 289.615
R121 source.n64 source.n38 289.615
R122 source.n96 source.n70 289.615
R123 source.n134 source.n108 289.615
R124 source.n259 source.n258 185
R125 source.n256 source.n255 185
R126 source.n265 source.n264 185
R127 source.n267 source.n266 185
R128 source.n252 source.n251 185
R129 source.n273 source.n272 185
R130 source.n275 source.n274 185
R131 source.n221 source.n220 185
R132 source.n218 source.n217 185
R133 source.n227 source.n226 185
R134 source.n229 source.n228 185
R135 source.n214 source.n213 185
R136 source.n235 source.n234 185
R137 source.n237 source.n236 185
R138 source.n189 source.n188 185
R139 source.n186 source.n185 185
R140 source.n195 source.n194 185
R141 source.n197 source.n196 185
R142 source.n182 source.n181 185
R143 source.n203 source.n202 185
R144 source.n205 source.n204 185
R145 source.n151 source.n150 185
R146 source.n148 source.n147 185
R147 source.n157 source.n156 185
R148 source.n159 source.n158 185
R149 source.n144 source.n143 185
R150 source.n165 source.n164 185
R151 source.n167 source.n166 185
R152 source.n27 source.n26 185
R153 source.n25 source.n24 185
R154 source.n4 source.n3 185
R155 source.n19 source.n18 185
R156 source.n17 source.n16 185
R157 source.n8 source.n7 185
R158 source.n11 source.n10 185
R159 source.n65 source.n64 185
R160 source.n63 source.n62 185
R161 source.n42 source.n41 185
R162 source.n57 source.n56 185
R163 source.n55 source.n54 185
R164 source.n46 source.n45 185
R165 source.n49 source.n48 185
R166 source.n97 source.n96 185
R167 source.n95 source.n94 185
R168 source.n74 source.n73 185
R169 source.n89 source.n88 185
R170 source.n87 source.n86 185
R171 source.n78 source.n77 185
R172 source.n81 source.n80 185
R173 source.n135 source.n134 185
R174 source.n133 source.n132 185
R175 source.n112 source.n111 185
R176 source.n127 source.n126 185
R177 source.n125 source.n124 185
R178 source.n116 source.n115 185
R179 source.n119 source.n118 185
R180 source.t0 source.n257 147.661
R181 source.t2 source.n219 147.661
R182 source.t24 source.n187 147.661
R183 source.t22 source.n149 147.661
R184 source.t30 source.n9 147.661
R185 source.t18 source.n47 147.661
R186 source.t5 source.n79 147.661
R187 source.t15 source.n117 147.661
R188 source.n258 source.n255 104.615
R189 source.n265 source.n255 104.615
R190 source.n266 source.n265 104.615
R191 source.n266 source.n251 104.615
R192 source.n273 source.n251 104.615
R193 source.n274 source.n273 104.615
R194 source.n220 source.n217 104.615
R195 source.n227 source.n217 104.615
R196 source.n228 source.n227 104.615
R197 source.n228 source.n213 104.615
R198 source.n235 source.n213 104.615
R199 source.n236 source.n235 104.615
R200 source.n188 source.n185 104.615
R201 source.n195 source.n185 104.615
R202 source.n196 source.n195 104.615
R203 source.n196 source.n181 104.615
R204 source.n203 source.n181 104.615
R205 source.n204 source.n203 104.615
R206 source.n150 source.n147 104.615
R207 source.n157 source.n147 104.615
R208 source.n158 source.n157 104.615
R209 source.n158 source.n143 104.615
R210 source.n165 source.n143 104.615
R211 source.n166 source.n165 104.615
R212 source.n26 source.n25 104.615
R213 source.n25 source.n3 104.615
R214 source.n18 source.n3 104.615
R215 source.n18 source.n17 104.615
R216 source.n17 source.n7 104.615
R217 source.n10 source.n7 104.615
R218 source.n64 source.n63 104.615
R219 source.n63 source.n41 104.615
R220 source.n56 source.n41 104.615
R221 source.n56 source.n55 104.615
R222 source.n55 source.n45 104.615
R223 source.n48 source.n45 104.615
R224 source.n96 source.n95 104.615
R225 source.n95 source.n73 104.615
R226 source.n88 source.n73 104.615
R227 source.n88 source.n87 104.615
R228 source.n87 source.n77 104.615
R229 source.n80 source.n77 104.615
R230 source.n134 source.n133 104.615
R231 source.n133 source.n111 104.615
R232 source.n126 source.n111 104.615
R233 source.n126 source.n125 104.615
R234 source.n125 source.n115 104.615
R235 source.n118 source.n115 104.615
R236 source.n258 source.t0 52.3082
R237 source.n220 source.t2 52.3082
R238 source.n188 source.t24 52.3082
R239 source.n150 source.t22 52.3082
R240 source.n10 source.t30 52.3082
R241 source.n48 source.t18 52.3082
R242 source.n80 source.t5 52.3082
R243 source.n118 source.t15 52.3082
R244 source.n33 source.n32 50.512
R245 source.n35 source.n34 50.512
R246 source.n37 source.n36 50.512
R247 source.n103 source.n102 50.512
R248 source.n105 source.n104 50.512
R249 source.n107 source.n106 50.512
R250 source.n247 source.n246 50.5119
R251 source.n245 source.n244 50.5119
R252 source.n243 source.n242 50.5119
R253 source.n177 source.n176 50.5119
R254 source.n175 source.n174 50.5119
R255 source.n173 source.n172 50.5119
R256 source.n279 source.n278 32.1853
R257 source.n241 source.n240 32.1853
R258 source.n209 source.n208 32.1853
R259 source.n171 source.n170 32.1853
R260 source.n31 source.n30 32.1853
R261 source.n69 source.n68 32.1853
R262 source.n101 source.n100 32.1853
R263 source.n139 source.n138 32.1853
R264 source.n171 source.n139 17.544
R265 source.n259 source.n257 15.6674
R266 source.n221 source.n219 15.6674
R267 source.n189 source.n187 15.6674
R268 source.n151 source.n149 15.6674
R269 source.n11 source.n9 15.6674
R270 source.n49 source.n47 15.6674
R271 source.n81 source.n79 15.6674
R272 source.n119 source.n117 15.6674
R273 source.n260 source.n256 12.8005
R274 source.n222 source.n218 12.8005
R275 source.n190 source.n186 12.8005
R276 source.n152 source.n148 12.8005
R277 source.n12 source.n8 12.8005
R278 source.n50 source.n46 12.8005
R279 source.n82 source.n78 12.8005
R280 source.n120 source.n116 12.8005
R281 source.n264 source.n263 12.0247
R282 source.n226 source.n225 12.0247
R283 source.n194 source.n193 12.0247
R284 source.n156 source.n155 12.0247
R285 source.n16 source.n15 12.0247
R286 source.n54 source.n53 12.0247
R287 source.n86 source.n85 12.0247
R288 source.n124 source.n123 12.0247
R289 source.n280 source.n31 11.8802
R290 source.n267 source.n254 11.249
R291 source.n229 source.n216 11.249
R292 source.n197 source.n184 11.249
R293 source.n159 source.n146 11.249
R294 source.n19 source.n6 11.249
R295 source.n57 source.n44 11.249
R296 source.n89 source.n76 11.249
R297 source.n127 source.n114 11.249
R298 source.n268 source.n252 10.4732
R299 source.n230 source.n214 10.4732
R300 source.n198 source.n182 10.4732
R301 source.n160 source.n144 10.4732
R302 source.n20 source.n4 10.4732
R303 source.n58 source.n42 10.4732
R304 source.n90 source.n74 10.4732
R305 source.n128 source.n112 10.4732
R306 source.n272 source.n271 9.69747
R307 source.n234 source.n233 9.69747
R308 source.n202 source.n201 9.69747
R309 source.n164 source.n163 9.69747
R310 source.n24 source.n23 9.69747
R311 source.n62 source.n61 9.69747
R312 source.n94 source.n93 9.69747
R313 source.n132 source.n131 9.69747
R314 source.n278 source.n277 9.45567
R315 source.n240 source.n239 9.45567
R316 source.n208 source.n207 9.45567
R317 source.n170 source.n169 9.45567
R318 source.n30 source.n29 9.45567
R319 source.n68 source.n67 9.45567
R320 source.n100 source.n99 9.45567
R321 source.n138 source.n137 9.45567
R322 source.n277 source.n276 9.3005
R323 source.n250 source.n249 9.3005
R324 source.n271 source.n270 9.3005
R325 source.n269 source.n268 9.3005
R326 source.n254 source.n253 9.3005
R327 source.n263 source.n262 9.3005
R328 source.n261 source.n260 9.3005
R329 source.n239 source.n238 9.3005
R330 source.n212 source.n211 9.3005
R331 source.n233 source.n232 9.3005
R332 source.n231 source.n230 9.3005
R333 source.n216 source.n215 9.3005
R334 source.n225 source.n224 9.3005
R335 source.n223 source.n222 9.3005
R336 source.n207 source.n206 9.3005
R337 source.n180 source.n179 9.3005
R338 source.n201 source.n200 9.3005
R339 source.n199 source.n198 9.3005
R340 source.n184 source.n183 9.3005
R341 source.n193 source.n192 9.3005
R342 source.n191 source.n190 9.3005
R343 source.n169 source.n168 9.3005
R344 source.n142 source.n141 9.3005
R345 source.n163 source.n162 9.3005
R346 source.n161 source.n160 9.3005
R347 source.n146 source.n145 9.3005
R348 source.n155 source.n154 9.3005
R349 source.n153 source.n152 9.3005
R350 source.n29 source.n28 9.3005
R351 source.n2 source.n1 9.3005
R352 source.n23 source.n22 9.3005
R353 source.n21 source.n20 9.3005
R354 source.n6 source.n5 9.3005
R355 source.n15 source.n14 9.3005
R356 source.n13 source.n12 9.3005
R357 source.n67 source.n66 9.3005
R358 source.n40 source.n39 9.3005
R359 source.n61 source.n60 9.3005
R360 source.n59 source.n58 9.3005
R361 source.n44 source.n43 9.3005
R362 source.n53 source.n52 9.3005
R363 source.n51 source.n50 9.3005
R364 source.n99 source.n98 9.3005
R365 source.n72 source.n71 9.3005
R366 source.n93 source.n92 9.3005
R367 source.n91 source.n90 9.3005
R368 source.n76 source.n75 9.3005
R369 source.n85 source.n84 9.3005
R370 source.n83 source.n82 9.3005
R371 source.n137 source.n136 9.3005
R372 source.n110 source.n109 9.3005
R373 source.n131 source.n130 9.3005
R374 source.n129 source.n128 9.3005
R375 source.n114 source.n113 9.3005
R376 source.n123 source.n122 9.3005
R377 source.n121 source.n120 9.3005
R378 source.n275 source.n250 8.92171
R379 source.n237 source.n212 8.92171
R380 source.n205 source.n180 8.92171
R381 source.n167 source.n142 8.92171
R382 source.n27 source.n2 8.92171
R383 source.n65 source.n40 8.92171
R384 source.n97 source.n72 8.92171
R385 source.n135 source.n110 8.92171
R386 source.n276 source.n248 8.14595
R387 source.n238 source.n210 8.14595
R388 source.n206 source.n178 8.14595
R389 source.n168 source.n140 8.14595
R390 source.n28 source.n0 8.14595
R391 source.n66 source.n38 8.14595
R392 source.n98 source.n70 8.14595
R393 source.n136 source.n108 8.14595
R394 source.n278 source.n248 5.81868
R395 source.n240 source.n210 5.81868
R396 source.n208 source.n178 5.81868
R397 source.n170 source.n140 5.81868
R398 source.n30 source.n0 5.81868
R399 source.n68 source.n38 5.81868
R400 source.n100 source.n70 5.81868
R401 source.n138 source.n108 5.81868
R402 source.n280 source.n279 5.66429
R403 source.n276 source.n275 5.04292
R404 source.n238 source.n237 5.04292
R405 source.n206 source.n205 5.04292
R406 source.n168 source.n167 5.04292
R407 source.n28 source.n27 5.04292
R408 source.n66 source.n65 5.04292
R409 source.n98 source.n97 5.04292
R410 source.n136 source.n135 5.04292
R411 source.n261 source.n257 4.38594
R412 source.n223 source.n219 4.38594
R413 source.n191 source.n187 4.38594
R414 source.n153 source.n149 4.38594
R415 source.n13 source.n9 4.38594
R416 source.n51 source.n47 4.38594
R417 source.n83 source.n79 4.38594
R418 source.n121 source.n117 4.38594
R419 source.n272 source.n250 4.26717
R420 source.n234 source.n212 4.26717
R421 source.n202 source.n180 4.26717
R422 source.n164 source.n142 4.26717
R423 source.n24 source.n2 4.26717
R424 source.n62 source.n40 4.26717
R425 source.n94 source.n72 4.26717
R426 source.n132 source.n110 4.26717
R427 source.n271 source.n252 3.49141
R428 source.n233 source.n214 3.49141
R429 source.n201 source.n182 3.49141
R430 source.n163 source.n144 3.49141
R431 source.n23 source.n4 3.49141
R432 source.n61 source.n42 3.49141
R433 source.n93 source.n74 3.49141
R434 source.n131 source.n112 3.49141
R435 source.n246 source.t6 3.3005
R436 source.n246 source.t3 3.3005
R437 source.n244 source.t1 3.3005
R438 source.n244 source.t12 3.3005
R439 source.n242 source.t4 3.3005
R440 source.n242 source.t8 3.3005
R441 source.n176 source.t27 3.3005
R442 source.n176 source.t31 3.3005
R443 source.n174 source.t17 3.3005
R444 source.n174 source.t23 3.3005
R445 source.n172 source.t26 3.3005
R446 source.n172 source.t16 3.3005
R447 source.n32 source.t28 3.3005
R448 source.n32 source.t29 3.3005
R449 source.n34 source.t21 3.3005
R450 source.n34 source.t25 3.3005
R451 source.n36 source.t19 3.3005
R452 source.n36 source.t20 3.3005
R453 source.n102 source.t7 3.3005
R454 source.n102 source.t11 3.3005
R455 source.n104 source.t9 3.3005
R456 source.n104 source.t14 3.3005
R457 source.n106 source.t13 3.3005
R458 source.n106 source.t10 3.3005
R459 source.n268 source.n267 2.71565
R460 source.n230 source.n229 2.71565
R461 source.n198 source.n197 2.71565
R462 source.n160 source.n159 2.71565
R463 source.n20 source.n19 2.71565
R464 source.n58 source.n57 2.71565
R465 source.n90 source.n89 2.71565
R466 source.n128 source.n127 2.71565
R467 source.n264 source.n254 1.93989
R468 source.n226 source.n216 1.93989
R469 source.n194 source.n184 1.93989
R470 source.n156 source.n146 1.93989
R471 source.n16 source.n6 1.93989
R472 source.n54 source.n44 1.93989
R473 source.n86 source.n76 1.93989
R474 source.n124 source.n114 1.93989
R475 source.n263 source.n256 1.16414
R476 source.n225 source.n218 1.16414
R477 source.n193 source.n186 1.16414
R478 source.n155 source.n148 1.16414
R479 source.n15 source.n8 1.16414
R480 source.n53 source.n46 1.16414
R481 source.n85 source.n78 1.16414
R482 source.n123 source.n116 1.16414
R483 source.n139 source.n107 0.802224
R484 source.n107 source.n105 0.802224
R485 source.n105 source.n103 0.802224
R486 source.n103 source.n101 0.802224
R487 source.n69 source.n37 0.802224
R488 source.n37 source.n35 0.802224
R489 source.n35 source.n33 0.802224
R490 source.n33 source.n31 0.802224
R491 source.n173 source.n171 0.802224
R492 source.n175 source.n173 0.802224
R493 source.n177 source.n175 0.802224
R494 source.n209 source.n177 0.802224
R495 source.n243 source.n241 0.802224
R496 source.n245 source.n243 0.802224
R497 source.n247 source.n245 0.802224
R498 source.n279 source.n247 0.802224
R499 source.n101 source.n69 0.470328
R500 source.n241 source.n209 0.470328
R501 source.n260 source.n259 0.388379
R502 source.n222 source.n221 0.388379
R503 source.n190 source.n189 0.388379
R504 source.n152 source.n151 0.388379
R505 source.n12 source.n11 0.388379
R506 source.n50 source.n49 0.388379
R507 source.n82 source.n81 0.388379
R508 source.n120 source.n119 0.388379
R509 source source.n280 0.188
R510 source.n262 source.n261 0.155672
R511 source.n262 source.n253 0.155672
R512 source.n269 source.n253 0.155672
R513 source.n270 source.n269 0.155672
R514 source.n270 source.n249 0.155672
R515 source.n277 source.n249 0.155672
R516 source.n224 source.n223 0.155672
R517 source.n224 source.n215 0.155672
R518 source.n231 source.n215 0.155672
R519 source.n232 source.n231 0.155672
R520 source.n232 source.n211 0.155672
R521 source.n239 source.n211 0.155672
R522 source.n192 source.n191 0.155672
R523 source.n192 source.n183 0.155672
R524 source.n199 source.n183 0.155672
R525 source.n200 source.n199 0.155672
R526 source.n200 source.n179 0.155672
R527 source.n207 source.n179 0.155672
R528 source.n154 source.n153 0.155672
R529 source.n154 source.n145 0.155672
R530 source.n161 source.n145 0.155672
R531 source.n162 source.n161 0.155672
R532 source.n162 source.n141 0.155672
R533 source.n169 source.n141 0.155672
R534 source.n29 source.n1 0.155672
R535 source.n22 source.n1 0.155672
R536 source.n22 source.n21 0.155672
R537 source.n21 source.n5 0.155672
R538 source.n14 source.n5 0.155672
R539 source.n14 source.n13 0.155672
R540 source.n67 source.n39 0.155672
R541 source.n60 source.n39 0.155672
R542 source.n60 source.n59 0.155672
R543 source.n59 source.n43 0.155672
R544 source.n52 source.n43 0.155672
R545 source.n52 source.n51 0.155672
R546 source.n99 source.n71 0.155672
R547 source.n92 source.n71 0.155672
R548 source.n92 source.n91 0.155672
R549 source.n91 source.n75 0.155672
R550 source.n84 source.n75 0.155672
R551 source.n84 source.n83 0.155672
R552 source.n137 source.n109 0.155672
R553 source.n130 source.n109 0.155672
R554 source.n130 source.n129 0.155672
R555 source.n129 source.n113 0.155672
R556 source.n122 source.n113 0.155672
R557 source.n122 source.n121 0.155672
R558 minus.n6 minus.t11 327.454
R559 minus.n30 minus.t4 327.454
R560 minus.n5 minus.t10 306.473
R561 minus.n9 minus.t9 306.473
R562 minus.n3 minus.t7 306.473
R563 minus.n15 minus.t2 306.473
R564 minus.n1 minus.t5 306.473
R565 minus.n21 minus.t3 306.473
R566 minus.n22 minus.t0 306.473
R567 minus.n29 minus.t14 306.473
R568 minus.n33 minus.t15 306.473
R569 minus.n27 minus.t8 306.473
R570 minus.n39 minus.t13 306.473
R571 minus.n25 minus.t12 306.473
R572 minus.n45 minus.t1 306.473
R573 minus.n46 minus.t6 306.473
R574 minus.n23 minus.n22 161.3
R575 minus.n21 minus.n0 161.3
R576 minus.n20 minus.n19 161.3
R577 minus.n18 minus.n1 161.3
R578 minus.n17 minus.n16 161.3
R579 minus.n15 minus.n2 161.3
R580 minus.n14 minus.n13 161.3
R581 minus.n12 minus.n3 161.3
R582 minus.n11 minus.n10 161.3
R583 minus.n9 minus.n4 161.3
R584 minus.n8 minus.n7 161.3
R585 minus.n47 minus.n46 161.3
R586 minus.n45 minus.n24 161.3
R587 minus.n44 minus.n43 161.3
R588 minus.n42 minus.n25 161.3
R589 minus.n41 minus.n40 161.3
R590 minus.n39 minus.n26 161.3
R591 minus.n38 minus.n37 161.3
R592 minus.n36 minus.n27 161.3
R593 minus.n35 minus.n34 161.3
R594 minus.n33 minus.n28 161.3
R595 minus.n32 minus.n31 161.3
R596 minus.n7 minus.n6 70.4033
R597 minus.n31 minus.n30 70.4033
R598 minus.n22 minus.n21 48.2005
R599 minus.n46 minus.n45 48.2005
R600 minus.n9 minus.n8 44.549
R601 minus.n20 minus.n1 44.549
R602 minus.n33 minus.n32 44.549
R603 minus.n44 minus.n25 44.549
R604 minus.n10 minus.n3 34.3247
R605 minus.n16 minus.n15 34.3247
R606 minus.n34 minus.n27 34.3247
R607 minus.n40 minus.n39 34.3247
R608 minus.n48 minus.n23 33.7846
R609 minus.n15 minus.n14 24.1005
R610 minus.n14 minus.n3 24.1005
R611 minus.n38 minus.n27 24.1005
R612 minus.n39 minus.n38 24.1005
R613 minus.n6 minus.n5 20.9576
R614 minus.n30 minus.n29 20.9576
R615 minus.n10 minus.n9 13.8763
R616 minus.n16 minus.n1 13.8763
R617 minus.n34 minus.n33 13.8763
R618 minus.n40 minus.n25 13.8763
R619 minus.n48 minus.n47 6.6558
R620 minus.n8 minus.n5 3.65202
R621 minus.n21 minus.n20 3.65202
R622 minus.n32 minus.n29 3.65202
R623 minus.n45 minus.n44 3.65202
R624 minus.n23 minus.n0 0.189894
R625 minus.n19 minus.n0 0.189894
R626 minus.n19 minus.n18 0.189894
R627 minus.n18 minus.n17 0.189894
R628 minus.n17 minus.n2 0.189894
R629 minus.n13 minus.n2 0.189894
R630 minus.n13 minus.n12 0.189894
R631 minus.n12 minus.n11 0.189894
R632 minus.n11 minus.n4 0.189894
R633 minus.n7 minus.n4 0.189894
R634 minus.n31 minus.n28 0.189894
R635 minus.n35 minus.n28 0.189894
R636 minus.n36 minus.n35 0.189894
R637 minus.n37 minus.n36 0.189894
R638 minus.n37 minus.n26 0.189894
R639 minus.n41 minus.n26 0.189894
R640 minus.n42 minus.n41 0.189894
R641 minus.n43 minus.n42 0.189894
R642 minus.n43 minus.n24 0.189894
R643 minus.n47 minus.n24 0.189894
R644 minus minus.n48 0.188
R645 drain_right.n5 drain_right.n3 67.9924
R646 drain_right.n2 drain_right.n0 67.9924
R647 drain_right.n9 drain_right.n7 67.9924
R648 drain_right.n9 drain_right.n8 67.1908
R649 drain_right.n11 drain_right.n10 67.1908
R650 drain_right.n13 drain_right.n12 67.1908
R651 drain_right.n5 drain_right.n4 67.1907
R652 drain_right.n2 drain_right.n1 67.1907
R653 drain_right drain_right.n6 27.4796
R654 drain_right drain_right.n13 6.45494
R655 drain_right.n3 drain_right.t14 3.3005
R656 drain_right.n3 drain_right.t9 3.3005
R657 drain_right.n4 drain_right.t2 3.3005
R658 drain_right.n4 drain_right.t3 3.3005
R659 drain_right.n1 drain_right.t0 3.3005
R660 drain_right.n1 drain_right.t7 3.3005
R661 drain_right.n0 drain_right.t11 3.3005
R662 drain_right.n0 drain_right.t1 3.3005
R663 drain_right.n7 drain_right.t5 3.3005
R664 drain_right.n7 drain_right.t4 3.3005
R665 drain_right.n8 drain_right.t8 3.3005
R666 drain_right.n8 drain_right.t6 3.3005
R667 drain_right.n10 drain_right.t10 3.3005
R668 drain_right.n10 drain_right.t13 3.3005
R669 drain_right.n12 drain_right.t15 3.3005
R670 drain_right.n12 drain_right.t12 3.3005
R671 drain_right.n13 drain_right.n11 0.802224
R672 drain_right.n11 drain_right.n9 0.802224
R673 drain_right.n6 drain_right.n5 0.346016
R674 drain_right.n6 drain_right.n2 0.346016
C0 source drain_left 12.3496f
C1 drain_left plus 5.20197f
C2 minus drain_right 4.96607f
C3 source minus 5.24444f
C4 minus plus 5.01313f
C5 drain_left minus 0.172752f
C6 source drain_right 12.351299f
C7 drain_right plus 0.391974f
C8 drain_left drain_right 1.24373f
C9 source plus 5.25846f
C10 drain_right a_n2390_n2088# 5.502571f
C11 drain_left a_n2390_n2088# 5.83464f
C12 source a_n2390_n2088# 5.603483f
C13 minus a_n2390_n2088# 8.97676f
C14 plus a_n2390_n2088# 10.48641f
C15 drain_right.t11 a_n2390_n2088# 0.132302f
C16 drain_right.t1 a_n2390_n2088# 0.132302f
C17 drain_right.n0 a_n2390_n2088# 1.1079f
C18 drain_right.t0 a_n2390_n2088# 0.132302f
C19 drain_right.t7 a_n2390_n2088# 0.132302f
C20 drain_right.n1 a_n2390_n2088# 1.1034f
C21 drain_right.n2 a_n2390_n2088# 0.708879f
C22 drain_right.t14 a_n2390_n2088# 0.132302f
C23 drain_right.t9 a_n2390_n2088# 0.132302f
C24 drain_right.n3 a_n2390_n2088# 1.1079f
C25 drain_right.t2 a_n2390_n2088# 0.132302f
C26 drain_right.t3 a_n2390_n2088# 0.132302f
C27 drain_right.n4 a_n2390_n2088# 1.1034f
C28 drain_right.n5 a_n2390_n2088# 0.708879f
C29 drain_right.n6 a_n2390_n2088# 1.12128f
C30 drain_right.t5 a_n2390_n2088# 0.132302f
C31 drain_right.t4 a_n2390_n2088# 0.132302f
C32 drain_right.n7 a_n2390_n2088# 1.1079f
C33 drain_right.t8 a_n2390_n2088# 0.132302f
C34 drain_right.t6 a_n2390_n2088# 0.132302f
C35 drain_right.n8 a_n2390_n2088# 1.1034f
C36 drain_right.n9 a_n2390_n2088# 0.74802f
C37 drain_right.t10 a_n2390_n2088# 0.132302f
C38 drain_right.t13 a_n2390_n2088# 0.132302f
C39 drain_right.n10 a_n2390_n2088# 1.1034f
C40 drain_right.n11 a_n2390_n2088# 0.370639f
C41 drain_right.t15 a_n2390_n2088# 0.132302f
C42 drain_right.t12 a_n2390_n2088# 0.132302f
C43 drain_right.n12 a_n2390_n2088# 1.1034f
C44 drain_right.n13 a_n2390_n2088# 0.613957f
C45 minus.n0 a_n2390_n2088# 0.043354f
C46 minus.t5 a_n2390_n2088# 0.4527f
C47 minus.n1 a_n2390_n2088# 0.213152f
C48 minus.n2 a_n2390_n2088# 0.043354f
C49 minus.t7 a_n2390_n2088# 0.4527f
C50 minus.n3 a_n2390_n2088# 0.213152f
C51 minus.n4 a_n2390_n2088# 0.043354f
C52 minus.t10 a_n2390_n2088# 0.4527f
C53 minus.n5 a_n2390_n2088# 0.211949f
C54 minus.t11 a_n2390_n2088# 0.466242f
C55 minus.n6 a_n2390_n2088# 0.198085f
C56 minus.n7 a_n2390_n2088# 0.146019f
C57 minus.n8 a_n2390_n2088# 0.009838f
C58 minus.t9 a_n2390_n2088# 0.4527f
C59 minus.n9 a_n2390_n2088# 0.213152f
C60 minus.n10 a_n2390_n2088# 0.009838f
C61 minus.n11 a_n2390_n2088# 0.043354f
C62 minus.n12 a_n2390_n2088# 0.043354f
C63 minus.n13 a_n2390_n2088# 0.043354f
C64 minus.n14 a_n2390_n2088# 0.009838f
C65 minus.t2 a_n2390_n2088# 0.4527f
C66 minus.n15 a_n2390_n2088# 0.213152f
C67 minus.n16 a_n2390_n2088# 0.009838f
C68 minus.n17 a_n2390_n2088# 0.043354f
C69 minus.n18 a_n2390_n2088# 0.043354f
C70 minus.n19 a_n2390_n2088# 0.043354f
C71 minus.n20 a_n2390_n2088# 0.009838f
C72 minus.t3 a_n2390_n2088# 0.4527f
C73 minus.n21 a_n2390_n2088# 0.211949f
C74 minus.t0 a_n2390_n2088# 0.4527f
C75 minus.n22 a_n2390_n2088# 0.211281f
C76 minus.n23 a_n2390_n2088# 1.37904f
C77 minus.n24 a_n2390_n2088# 0.043354f
C78 minus.t12 a_n2390_n2088# 0.4527f
C79 minus.n25 a_n2390_n2088# 0.213152f
C80 minus.n26 a_n2390_n2088# 0.043354f
C81 minus.t8 a_n2390_n2088# 0.4527f
C82 minus.n27 a_n2390_n2088# 0.213152f
C83 minus.n28 a_n2390_n2088# 0.043354f
C84 minus.t14 a_n2390_n2088# 0.4527f
C85 minus.n29 a_n2390_n2088# 0.211949f
C86 minus.t4 a_n2390_n2088# 0.466242f
C87 minus.n30 a_n2390_n2088# 0.198085f
C88 minus.n31 a_n2390_n2088# 0.146019f
C89 minus.n32 a_n2390_n2088# 0.009838f
C90 minus.t15 a_n2390_n2088# 0.4527f
C91 minus.n33 a_n2390_n2088# 0.213152f
C92 minus.n34 a_n2390_n2088# 0.009838f
C93 minus.n35 a_n2390_n2088# 0.043354f
C94 minus.n36 a_n2390_n2088# 0.043354f
C95 minus.n37 a_n2390_n2088# 0.043354f
C96 minus.n38 a_n2390_n2088# 0.009838f
C97 minus.t13 a_n2390_n2088# 0.4527f
C98 minus.n39 a_n2390_n2088# 0.213152f
C99 minus.n40 a_n2390_n2088# 0.009838f
C100 minus.n41 a_n2390_n2088# 0.043354f
C101 minus.n42 a_n2390_n2088# 0.043354f
C102 minus.n43 a_n2390_n2088# 0.043354f
C103 minus.n44 a_n2390_n2088# 0.009838f
C104 minus.t1 a_n2390_n2088# 0.4527f
C105 minus.n45 a_n2390_n2088# 0.211949f
C106 minus.t6 a_n2390_n2088# 0.4527f
C107 minus.n46 a_n2390_n2088# 0.211281f
C108 minus.n47 a_n2390_n2088# 0.299234f
C109 minus.n48 a_n2390_n2088# 1.68045f
C110 source.n0 a_n2390_n2088# 0.035966f
C111 source.n1 a_n2390_n2088# 0.025588f
C112 source.n2 a_n2390_n2088# 0.01375f
C113 source.n3 a_n2390_n2088# 0.032499f
C114 source.n4 a_n2390_n2088# 0.014558f
C115 source.n5 a_n2390_n2088# 0.025588f
C116 source.n6 a_n2390_n2088# 0.01375f
C117 source.n7 a_n2390_n2088# 0.032499f
C118 source.n8 a_n2390_n2088# 0.014558f
C119 source.n9 a_n2390_n2088# 0.109497f
C120 source.t30 a_n2390_n2088# 0.05297f
C121 source.n10 a_n2390_n2088# 0.024374f
C122 source.n11 a_n2390_n2088# 0.019197f
C123 source.n12 a_n2390_n2088# 0.01375f
C124 source.n13 a_n2390_n2088# 0.608832f
C125 source.n14 a_n2390_n2088# 0.025588f
C126 source.n15 a_n2390_n2088# 0.01375f
C127 source.n16 a_n2390_n2088# 0.014558f
C128 source.n17 a_n2390_n2088# 0.032499f
C129 source.n18 a_n2390_n2088# 0.032499f
C130 source.n19 a_n2390_n2088# 0.014558f
C131 source.n20 a_n2390_n2088# 0.01375f
C132 source.n21 a_n2390_n2088# 0.025588f
C133 source.n22 a_n2390_n2088# 0.025588f
C134 source.n23 a_n2390_n2088# 0.01375f
C135 source.n24 a_n2390_n2088# 0.014558f
C136 source.n25 a_n2390_n2088# 0.032499f
C137 source.n26 a_n2390_n2088# 0.070355f
C138 source.n27 a_n2390_n2088# 0.014558f
C139 source.n28 a_n2390_n2088# 0.01375f
C140 source.n29 a_n2390_n2088# 0.059145f
C141 source.n30 a_n2390_n2088# 0.039367f
C142 source.n31 a_n2390_n2088# 0.656292f
C143 source.t28 a_n2390_n2088# 0.121321f
C144 source.t29 a_n2390_n2088# 0.121321f
C145 source.n32 a_n2390_n2088# 0.944855f
C146 source.n33 a_n2390_n2088# 0.372062f
C147 source.t21 a_n2390_n2088# 0.121321f
C148 source.t25 a_n2390_n2088# 0.121321f
C149 source.n34 a_n2390_n2088# 0.944855f
C150 source.n35 a_n2390_n2088# 0.372062f
C151 source.t19 a_n2390_n2088# 0.121321f
C152 source.t20 a_n2390_n2088# 0.121321f
C153 source.n36 a_n2390_n2088# 0.944855f
C154 source.n37 a_n2390_n2088# 0.372062f
C155 source.n38 a_n2390_n2088# 0.035966f
C156 source.n39 a_n2390_n2088# 0.025588f
C157 source.n40 a_n2390_n2088# 0.01375f
C158 source.n41 a_n2390_n2088# 0.032499f
C159 source.n42 a_n2390_n2088# 0.014558f
C160 source.n43 a_n2390_n2088# 0.025588f
C161 source.n44 a_n2390_n2088# 0.01375f
C162 source.n45 a_n2390_n2088# 0.032499f
C163 source.n46 a_n2390_n2088# 0.014558f
C164 source.n47 a_n2390_n2088# 0.109497f
C165 source.t18 a_n2390_n2088# 0.05297f
C166 source.n48 a_n2390_n2088# 0.024374f
C167 source.n49 a_n2390_n2088# 0.019197f
C168 source.n50 a_n2390_n2088# 0.01375f
C169 source.n51 a_n2390_n2088# 0.608832f
C170 source.n52 a_n2390_n2088# 0.025588f
C171 source.n53 a_n2390_n2088# 0.01375f
C172 source.n54 a_n2390_n2088# 0.014558f
C173 source.n55 a_n2390_n2088# 0.032499f
C174 source.n56 a_n2390_n2088# 0.032499f
C175 source.n57 a_n2390_n2088# 0.014558f
C176 source.n58 a_n2390_n2088# 0.01375f
C177 source.n59 a_n2390_n2088# 0.025588f
C178 source.n60 a_n2390_n2088# 0.025588f
C179 source.n61 a_n2390_n2088# 0.01375f
C180 source.n62 a_n2390_n2088# 0.014558f
C181 source.n63 a_n2390_n2088# 0.032499f
C182 source.n64 a_n2390_n2088# 0.070355f
C183 source.n65 a_n2390_n2088# 0.014558f
C184 source.n66 a_n2390_n2088# 0.01375f
C185 source.n67 a_n2390_n2088# 0.059145f
C186 source.n68 a_n2390_n2088# 0.039367f
C187 source.n69 a_n2390_n2088# 0.126692f
C188 source.n70 a_n2390_n2088# 0.035966f
C189 source.n71 a_n2390_n2088# 0.025588f
C190 source.n72 a_n2390_n2088# 0.01375f
C191 source.n73 a_n2390_n2088# 0.032499f
C192 source.n74 a_n2390_n2088# 0.014558f
C193 source.n75 a_n2390_n2088# 0.025588f
C194 source.n76 a_n2390_n2088# 0.01375f
C195 source.n77 a_n2390_n2088# 0.032499f
C196 source.n78 a_n2390_n2088# 0.014558f
C197 source.n79 a_n2390_n2088# 0.109497f
C198 source.t5 a_n2390_n2088# 0.05297f
C199 source.n80 a_n2390_n2088# 0.024374f
C200 source.n81 a_n2390_n2088# 0.019197f
C201 source.n82 a_n2390_n2088# 0.01375f
C202 source.n83 a_n2390_n2088# 0.608832f
C203 source.n84 a_n2390_n2088# 0.025588f
C204 source.n85 a_n2390_n2088# 0.01375f
C205 source.n86 a_n2390_n2088# 0.014558f
C206 source.n87 a_n2390_n2088# 0.032499f
C207 source.n88 a_n2390_n2088# 0.032499f
C208 source.n89 a_n2390_n2088# 0.014558f
C209 source.n90 a_n2390_n2088# 0.01375f
C210 source.n91 a_n2390_n2088# 0.025588f
C211 source.n92 a_n2390_n2088# 0.025588f
C212 source.n93 a_n2390_n2088# 0.01375f
C213 source.n94 a_n2390_n2088# 0.014558f
C214 source.n95 a_n2390_n2088# 0.032499f
C215 source.n96 a_n2390_n2088# 0.070355f
C216 source.n97 a_n2390_n2088# 0.014558f
C217 source.n98 a_n2390_n2088# 0.01375f
C218 source.n99 a_n2390_n2088# 0.059145f
C219 source.n100 a_n2390_n2088# 0.039367f
C220 source.n101 a_n2390_n2088# 0.126692f
C221 source.t7 a_n2390_n2088# 0.121321f
C222 source.t11 a_n2390_n2088# 0.121321f
C223 source.n102 a_n2390_n2088# 0.944855f
C224 source.n103 a_n2390_n2088# 0.372062f
C225 source.t9 a_n2390_n2088# 0.121321f
C226 source.t14 a_n2390_n2088# 0.121321f
C227 source.n104 a_n2390_n2088# 0.944855f
C228 source.n105 a_n2390_n2088# 0.372062f
C229 source.t13 a_n2390_n2088# 0.121321f
C230 source.t10 a_n2390_n2088# 0.121321f
C231 source.n106 a_n2390_n2088# 0.944855f
C232 source.n107 a_n2390_n2088# 0.372062f
C233 source.n108 a_n2390_n2088# 0.035966f
C234 source.n109 a_n2390_n2088# 0.025588f
C235 source.n110 a_n2390_n2088# 0.01375f
C236 source.n111 a_n2390_n2088# 0.032499f
C237 source.n112 a_n2390_n2088# 0.014558f
C238 source.n113 a_n2390_n2088# 0.025588f
C239 source.n114 a_n2390_n2088# 0.01375f
C240 source.n115 a_n2390_n2088# 0.032499f
C241 source.n116 a_n2390_n2088# 0.014558f
C242 source.n117 a_n2390_n2088# 0.109497f
C243 source.t15 a_n2390_n2088# 0.05297f
C244 source.n118 a_n2390_n2088# 0.024374f
C245 source.n119 a_n2390_n2088# 0.019197f
C246 source.n120 a_n2390_n2088# 0.01375f
C247 source.n121 a_n2390_n2088# 0.608832f
C248 source.n122 a_n2390_n2088# 0.025588f
C249 source.n123 a_n2390_n2088# 0.01375f
C250 source.n124 a_n2390_n2088# 0.014558f
C251 source.n125 a_n2390_n2088# 0.032499f
C252 source.n126 a_n2390_n2088# 0.032499f
C253 source.n127 a_n2390_n2088# 0.014558f
C254 source.n128 a_n2390_n2088# 0.01375f
C255 source.n129 a_n2390_n2088# 0.025588f
C256 source.n130 a_n2390_n2088# 0.025588f
C257 source.n131 a_n2390_n2088# 0.01375f
C258 source.n132 a_n2390_n2088# 0.014558f
C259 source.n133 a_n2390_n2088# 0.032499f
C260 source.n134 a_n2390_n2088# 0.070355f
C261 source.n135 a_n2390_n2088# 0.014558f
C262 source.n136 a_n2390_n2088# 0.01375f
C263 source.n137 a_n2390_n2088# 0.059145f
C264 source.n138 a_n2390_n2088# 0.039367f
C265 source.n139 a_n2390_n2088# 0.991843f
C266 source.n140 a_n2390_n2088# 0.035966f
C267 source.n141 a_n2390_n2088# 0.025588f
C268 source.n142 a_n2390_n2088# 0.01375f
C269 source.n143 a_n2390_n2088# 0.032499f
C270 source.n144 a_n2390_n2088# 0.014558f
C271 source.n145 a_n2390_n2088# 0.025588f
C272 source.n146 a_n2390_n2088# 0.01375f
C273 source.n147 a_n2390_n2088# 0.032499f
C274 source.n148 a_n2390_n2088# 0.014558f
C275 source.n149 a_n2390_n2088# 0.109497f
C276 source.t22 a_n2390_n2088# 0.05297f
C277 source.n150 a_n2390_n2088# 0.024374f
C278 source.n151 a_n2390_n2088# 0.019197f
C279 source.n152 a_n2390_n2088# 0.01375f
C280 source.n153 a_n2390_n2088# 0.608832f
C281 source.n154 a_n2390_n2088# 0.025588f
C282 source.n155 a_n2390_n2088# 0.01375f
C283 source.n156 a_n2390_n2088# 0.014558f
C284 source.n157 a_n2390_n2088# 0.032499f
C285 source.n158 a_n2390_n2088# 0.032499f
C286 source.n159 a_n2390_n2088# 0.014558f
C287 source.n160 a_n2390_n2088# 0.01375f
C288 source.n161 a_n2390_n2088# 0.025588f
C289 source.n162 a_n2390_n2088# 0.025588f
C290 source.n163 a_n2390_n2088# 0.01375f
C291 source.n164 a_n2390_n2088# 0.014558f
C292 source.n165 a_n2390_n2088# 0.032499f
C293 source.n166 a_n2390_n2088# 0.070355f
C294 source.n167 a_n2390_n2088# 0.014558f
C295 source.n168 a_n2390_n2088# 0.01375f
C296 source.n169 a_n2390_n2088# 0.059145f
C297 source.n170 a_n2390_n2088# 0.039367f
C298 source.n171 a_n2390_n2088# 0.991843f
C299 source.t26 a_n2390_n2088# 0.121321f
C300 source.t16 a_n2390_n2088# 0.121321f
C301 source.n172 a_n2390_n2088# 0.944849f
C302 source.n173 a_n2390_n2088# 0.372069f
C303 source.t17 a_n2390_n2088# 0.121321f
C304 source.t23 a_n2390_n2088# 0.121321f
C305 source.n174 a_n2390_n2088# 0.944849f
C306 source.n175 a_n2390_n2088# 0.372069f
C307 source.t27 a_n2390_n2088# 0.121321f
C308 source.t31 a_n2390_n2088# 0.121321f
C309 source.n176 a_n2390_n2088# 0.944849f
C310 source.n177 a_n2390_n2088# 0.372069f
C311 source.n178 a_n2390_n2088# 0.035966f
C312 source.n179 a_n2390_n2088# 0.025588f
C313 source.n180 a_n2390_n2088# 0.01375f
C314 source.n181 a_n2390_n2088# 0.032499f
C315 source.n182 a_n2390_n2088# 0.014558f
C316 source.n183 a_n2390_n2088# 0.025588f
C317 source.n184 a_n2390_n2088# 0.01375f
C318 source.n185 a_n2390_n2088# 0.032499f
C319 source.n186 a_n2390_n2088# 0.014558f
C320 source.n187 a_n2390_n2088# 0.109497f
C321 source.t24 a_n2390_n2088# 0.05297f
C322 source.n188 a_n2390_n2088# 0.024374f
C323 source.n189 a_n2390_n2088# 0.019197f
C324 source.n190 a_n2390_n2088# 0.01375f
C325 source.n191 a_n2390_n2088# 0.608832f
C326 source.n192 a_n2390_n2088# 0.025588f
C327 source.n193 a_n2390_n2088# 0.01375f
C328 source.n194 a_n2390_n2088# 0.014558f
C329 source.n195 a_n2390_n2088# 0.032499f
C330 source.n196 a_n2390_n2088# 0.032499f
C331 source.n197 a_n2390_n2088# 0.014558f
C332 source.n198 a_n2390_n2088# 0.01375f
C333 source.n199 a_n2390_n2088# 0.025588f
C334 source.n200 a_n2390_n2088# 0.025588f
C335 source.n201 a_n2390_n2088# 0.01375f
C336 source.n202 a_n2390_n2088# 0.014558f
C337 source.n203 a_n2390_n2088# 0.032499f
C338 source.n204 a_n2390_n2088# 0.070355f
C339 source.n205 a_n2390_n2088# 0.014558f
C340 source.n206 a_n2390_n2088# 0.01375f
C341 source.n207 a_n2390_n2088# 0.059145f
C342 source.n208 a_n2390_n2088# 0.039367f
C343 source.n209 a_n2390_n2088# 0.126692f
C344 source.n210 a_n2390_n2088# 0.035966f
C345 source.n211 a_n2390_n2088# 0.025588f
C346 source.n212 a_n2390_n2088# 0.01375f
C347 source.n213 a_n2390_n2088# 0.032499f
C348 source.n214 a_n2390_n2088# 0.014558f
C349 source.n215 a_n2390_n2088# 0.025588f
C350 source.n216 a_n2390_n2088# 0.01375f
C351 source.n217 a_n2390_n2088# 0.032499f
C352 source.n218 a_n2390_n2088# 0.014558f
C353 source.n219 a_n2390_n2088# 0.109497f
C354 source.t2 a_n2390_n2088# 0.05297f
C355 source.n220 a_n2390_n2088# 0.024374f
C356 source.n221 a_n2390_n2088# 0.019197f
C357 source.n222 a_n2390_n2088# 0.01375f
C358 source.n223 a_n2390_n2088# 0.608832f
C359 source.n224 a_n2390_n2088# 0.025588f
C360 source.n225 a_n2390_n2088# 0.01375f
C361 source.n226 a_n2390_n2088# 0.014558f
C362 source.n227 a_n2390_n2088# 0.032499f
C363 source.n228 a_n2390_n2088# 0.032499f
C364 source.n229 a_n2390_n2088# 0.014558f
C365 source.n230 a_n2390_n2088# 0.01375f
C366 source.n231 a_n2390_n2088# 0.025588f
C367 source.n232 a_n2390_n2088# 0.025588f
C368 source.n233 a_n2390_n2088# 0.01375f
C369 source.n234 a_n2390_n2088# 0.014558f
C370 source.n235 a_n2390_n2088# 0.032499f
C371 source.n236 a_n2390_n2088# 0.070355f
C372 source.n237 a_n2390_n2088# 0.014558f
C373 source.n238 a_n2390_n2088# 0.01375f
C374 source.n239 a_n2390_n2088# 0.059145f
C375 source.n240 a_n2390_n2088# 0.039367f
C376 source.n241 a_n2390_n2088# 0.126692f
C377 source.t4 a_n2390_n2088# 0.121321f
C378 source.t8 a_n2390_n2088# 0.121321f
C379 source.n242 a_n2390_n2088# 0.944849f
C380 source.n243 a_n2390_n2088# 0.372069f
C381 source.t1 a_n2390_n2088# 0.121321f
C382 source.t12 a_n2390_n2088# 0.121321f
C383 source.n244 a_n2390_n2088# 0.944849f
C384 source.n245 a_n2390_n2088# 0.372069f
C385 source.t6 a_n2390_n2088# 0.121321f
C386 source.t3 a_n2390_n2088# 0.121321f
C387 source.n246 a_n2390_n2088# 0.944849f
C388 source.n247 a_n2390_n2088# 0.372069f
C389 source.n248 a_n2390_n2088# 0.035966f
C390 source.n249 a_n2390_n2088# 0.025588f
C391 source.n250 a_n2390_n2088# 0.01375f
C392 source.n251 a_n2390_n2088# 0.032499f
C393 source.n252 a_n2390_n2088# 0.014558f
C394 source.n253 a_n2390_n2088# 0.025588f
C395 source.n254 a_n2390_n2088# 0.01375f
C396 source.n255 a_n2390_n2088# 0.032499f
C397 source.n256 a_n2390_n2088# 0.014558f
C398 source.n257 a_n2390_n2088# 0.109497f
C399 source.t0 a_n2390_n2088# 0.05297f
C400 source.n258 a_n2390_n2088# 0.024374f
C401 source.n259 a_n2390_n2088# 0.019197f
C402 source.n260 a_n2390_n2088# 0.01375f
C403 source.n261 a_n2390_n2088# 0.608832f
C404 source.n262 a_n2390_n2088# 0.025588f
C405 source.n263 a_n2390_n2088# 0.01375f
C406 source.n264 a_n2390_n2088# 0.014558f
C407 source.n265 a_n2390_n2088# 0.032499f
C408 source.n266 a_n2390_n2088# 0.032499f
C409 source.n267 a_n2390_n2088# 0.014558f
C410 source.n268 a_n2390_n2088# 0.01375f
C411 source.n269 a_n2390_n2088# 0.025588f
C412 source.n270 a_n2390_n2088# 0.025588f
C413 source.n271 a_n2390_n2088# 0.01375f
C414 source.n272 a_n2390_n2088# 0.014558f
C415 source.n273 a_n2390_n2088# 0.032499f
C416 source.n274 a_n2390_n2088# 0.070355f
C417 source.n275 a_n2390_n2088# 0.014558f
C418 source.n276 a_n2390_n2088# 0.01375f
C419 source.n277 a_n2390_n2088# 0.059145f
C420 source.n278 a_n2390_n2088# 0.039367f
C421 source.n279 a_n2390_n2088# 0.288031f
C422 source.n280 a_n2390_n2088# 1.05756f
C423 drain_left.t14 a_n2390_n2088# 0.132233f
C424 drain_left.t2 a_n2390_n2088# 0.132233f
C425 drain_left.n0 a_n2390_n2088# 1.10732f
C426 drain_left.t4 a_n2390_n2088# 0.132233f
C427 drain_left.t9 a_n2390_n2088# 0.132233f
C428 drain_left.n1 a_n2390_n2088# 1.10282f
C429 drain_left.n2 a_n2390_n2088# 0.708508f
C430 drain_left.t13 a_n2390_n2088# 0.132233f
C431 drain_left.t7 a_n2390_n2088# 0.132233f
C432 drain_left.n3 a_n2390_n2088# 1.10732f
C433 drain_left.t5 a_n2390_n2088# 0.132233f
C434 drain_left.t6 a_n2390_n2088# 0.132233f
C435 drain_left.n4 a_n2390_n2088# 1.10282f
C436 drain_left.n5 a_n2390_n2088# 0.708508f
C437 drain_left.n6 a_n2390_n2088# 1.17682f
C438 drain_left.t11 a_n2390_n2088# 0.132233f
C439 drain_left.t15 a_n2390_n2088# 0.132233f
C440 drain_left.n7 a_n2390_n2088# 1.10733f
C441 drain_left.t1 a_n2390_n2088# 0.132233f
C442 drain_left.t0 a_n2390_n2088# 0.132233f
C443 drain_left.n8 a_n2390_n2088# 1.10283f
C444 drain_left.n9 a_n2390_n2088# 0.747623f
C445 drain_left.t12 a_n2390_n2088# 0.132233f
C446 drain_left.t8 a_n2390_n2088# 0.132233f
C447 drain_left.n10 a_n2390_n2088# 1.10283f
C448 drain_left.n11 a_n2390_n2088# 0.370445f
C449 drain_left.t3 a_n2390_n2088# 0.132233f
C450 drain_left.t10 a_n2390_n2088# 0.132233f
C451 drain_left.n12 a_n2390_n2088# 1.10282f
C452 drain_left.n13 a_n2390_n2088# 0.613641f
C453 plus.n0 a_n2390_n2088# 0.044466f
C454 plus.t1 a_n2390_n2088# 0.464313f
C455 plus.t2 a_n2390_n2088# 0.464313f
C456 plus.t3 a_n2390_n2088# 0.464313f
C457 plus.n1 a_n2390_n2088# 0.21862f
C458 plus.n2 a_n2390_n2088# 0.044466f
C459 plus.t6 a_n2390_n2088# 0.464313f
C460 plus.t10 a_n2390_n2088# 0.464313f
C461 plus.n3 a_n2390_n2088# 0.21862f
C462 plus.n4 a_n2390_n2088# 0.044466f
C463 plus.t11 a_n2390_n2088# 0.464313f
C464 plus.t12 a_n2390_n2088# 0.464313f
C465 plus.n5 a_n2390_n2088# 0.217386f
C466 plus.t13 a_n2390_n2088# 0.478202f
C467 plus.n6 a_n2390_n2088# 0.203167f
C468 plus.n7 a_n2390_n2088# 0.149765f
C469 plus.n8 a_n2390_n2088# 0.01009f
C470 plus.n9 a_n2390_n2088# 0.21862f
C471 plus.n10 a_n2390_n2088# 0.01009f
C472 plus.n11 a_n2390_n2088# 0.044466f
C473 plus.n12 a_n2390_n2088# 0.044466f
C474 plus.n13 a_n2390_n2088# 0.044466f
C475 plus.n14 a_n2390_n2088# 0.01009f
C476 plus.n15 a_n2390_n2088# 0.21862f
C477 plus.n16 a_n2390_n2088# 0.01009f
C478 plus.n17 a_n2390_n2088# 0.044466f
C479 plus.n18 a_n2390_n2088# 0.044466f
C480 plus.n19 a_n2390_n2088# 0.044466f
C481 plus.n20 a_n2390_n2088# 0.01009f
C482 plus.n21 a_n2390_n2088# 0.217386f
C483 plus.n22 a_n2390_n2088# 0.216701f
C484 plus.n23 a_n2390_n2088# 0.39796f
C485 plus.n24 a_n2390_n2088# 0.044466f
C486 plus.t9 a_n2390_n2088# 0.464313f
C487 plus.t5 a_n2390_n2088# 0.464313f
C488 plus.t15 a_n2390_n2088# 0.464313f
C489 plus.n25 a_n2390_n2088# 0.21862f
C490 plus.n26 a_n2390_n2088# 0.044466f
C491 plus.t14 a_n2390_n2088# 0.464313f
C492 plus.t8 a_n2390_n2088# 0.464313f
C493 plus.n27 a_n2390_n2088# 0.21862f
C494 plus.n28 a_n2390_n2088# 0.044466f
C495 plus.t4 a_n2390_n2088# 0.464313f
C496 plus.t0 a_n2390_n2088# 0.464313f
C497 plus.n29 a_n2390_n2088# 0.217386f
C498 plus.t7 a_n2390_n2088# 0.478202f
C499 plus.n30 a_n2390_n2088# 0.203167f
C500 plus.n31 a_n2390_n2088# 0.149765f
C501 plus.n32 a_n2390_n2088# 0.01009f
C502 plus.n33 a_n2390_n2088# 0.21862f
C503 plus.n34 a_n2390_n2088# 0.01009f
C504 plus.n35 a_n2390_n2088# 0.044466f
C505 plus.n36 a_n2390_n2088# 0.044466f
C506 plus.n37 a_n2390_n2088# 0.044466f
C507 plus.n38 a_n2390_n2088# 0.01009f
C508 plus.n39 a_n2390_n2088# 0.21862f
C509 plus.n40 a_n2390_n2088# 0.01009f
C510 plus.n41 a_n2390_n2088# 0.044466f
C511 plus.n42 a_n2390_n2088# 0.044466f
C512 plus.n43 a_n2390_n2088# 0.044466f
C513 plus.n44 a_n2390_n2088# 0.01009f
C514 plus.n45 a_n2390_n2088# 0.217386f
C515 plus.n46 a_n2390_n2088# 0.216701f
C516 plus.n47 a_n2390_n2088# 1.28015f
.ends

