* NGSPICE file created from diffpair568.ext - technology: sky130A

.subckt diffpair568 minus drain_right drain_left source plus
X0 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X1 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X4 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X5 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X6 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X7 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X8 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X9 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X10 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X13 a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X14 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X16 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X18 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X20 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X23 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X24 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X25 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X26 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X28 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X29 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X30 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X31 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X32 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X33 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X34 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X35 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X36 drain_right minus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X37 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X38 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X39 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X40 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X41 drain_left plus source a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X42 source minus drain_right a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X43 source plus drain_left a_n2146_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
.ends

