* NGSPICE file created from diffpair606.ext - technology: sky130A

.subckt diffpair606 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t19 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t22 plus.t1 drain_left.t12 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 drain_right.t13 minus.t0 source.t3 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X3 a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X4 a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X5 source.t9 minus.t1 drain_right.t12 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t25 plus.t2 drain_left.t11 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X7 drain_left.t10 plus.t3 source.t14 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 drain_left.t9 plus.t4 source.t17 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X9 source.t0 minus.t2 drain_right.t11 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 drain_right.t10 minus.t3 source.t13 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X11 drain_right.t9 minus.t4 source.t2 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X12 drain_right.t8 minus.t5 source.t7 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X13 drain_right.t7 minus.t6 source.t10 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X14 source.t20 plus.t5 drain_left.t8 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 drain_left.t7 plus.t6 source.t24 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X16 a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X17 drain_left.t6 plus.t7 source.t18 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X18 a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X19 drain_left.t5 plus.t8 source.t26 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X20 source.t5 minus.t7 drain_right.t6 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X21 source.t16 plus.t9 drain_left.t4 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X22 source.t6 minus.t8 drain_right.t5 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 drain_right.t4 minus.t9 source.t11 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X24 drain_right.t3 minus.t10 source.t4 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X25 source.t23 plus.t10 drain_left.t3 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X26 drain_right.t2 minus.t11 source.t8 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X27 source.t12 minus.t12 drain_right.t1 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X28 source.t1 minus.t13 drain_right.t0 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X29 drain_left.t2 plus.t11 source.t27 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X30 drain_left.t1 plus.t12 source.t15 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X31 source.t21 plus.t13 drain_left.t0 a_n2044_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
R0 plus.n4 plus.t4 1063.55
R1 plus.n20 plus.t0 1063.55
R2 plus.n14 plus.t8 1042.57
R3 plus.n13 plus.t13 1042.57
R4 plus.n1 plus.t11 1042.57
R5 plus.n8 plus.t5 1042.57
R6 plus.n7 plus.t12 1042.57
R7 plus.n3 plus.t10 1042.57
R8 plus.n30 plus.t6 1042.57
R9 plus.n29 plus.t9 1042.57
R10 plus.n17 plus.t3 1042.57
R11 plus.n24 plus.t2 1042.57
R12 plus.n23 plus.t7 1042.57
R13 plus.n19 plus.t1 1042.57
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n2 161.3
R16 plus.n10 plus.n1 161.3
R17 plus.n12 plus.n11 161.3
R18 plus.n13 plus.n0 161.3
R19 plus.n15 plus.n14 161.3
R20 plus.n22 plus.n21 161.3
R21 plus.n23 plus.n18 161.3
R22 plus.n26 plus.n17 161.3
R23 plus.n28 plus.n27 161.3
R24 plus.n29 plus.n16 161.3
R25 plus.n31 plus.n30 161.3
R26 plus.n9 plus.n8 80.6037
R27 plus.n25 plus.n24 80.6037
R28 plus.n5 plus.n4 70.4033
R29 plus.n21 plus.n20 70.4033
R30 plus.n14 plus.n13 48.2005
R31 plus.n8 plus.n1 48.2005
R32 plus.n8 plus.n7 48.2005
R33 plus.n30 plus.n29 48.2005
R34 plus.n24 plus.n17 48.2005
R35 plus.n24 plus.n23 48.2005
R36 plus plus.n31 33.8683
R37 plus.n12 plus.n1 24.8308
R38 plus.n7 plus.n6 24.8308
R39 plus.n28 plus.n17 24.8308
R40 plus.n23 plus.n22 24.8308
R41 plus.n13 plus.n12 23.3702
R42 plus.n6 plus.n3 23.3702
R43 plus.n29 plus.n28 23.3702
R44 plus.n22 plus.n19 23.3702
R45 plus.n4 plus.n3 20.9576
R46 plus.n20 plus.n19 20.9576
R47 plus plus.n15 15.2675
R48 plus.n9 plus.n2 0.285035
R49 plus.n10 plus.n9 0.285035
R50 plus.n26 plus.n25 0.285035
R51 plus.n25 plus.n18 0.285035
R52 plus.n5 plus.n2 0.189894
R53 plus.n11 plus.n10 0.189894
R54 plus.n11 plus.n0 0.189894
R55 plus.n15 plus.n0 0.189894
R56 plus.n31 plus.n16 0.189894
R57 plus.n27 plus.n16 0.189894
R58 plus.n27 plus.n26 0.189894
R59 plus.n21 plus.n18 0.189894
R60 source.n0 source.t26 44.1297
R61 source.n7 source.t11 44.1296
R62 source.n27 source.t8 44.1295
R63 source.n20 source.t19 44.1295
R64 source.n2 source.n1 43.1397
R65 source.n4 source.n3 43.1397
R66 source.n6 source.n5 43.1397
R67 source.n9 source.n8 43.1397
R68 source.n11 source.n10 43.1397
R69 source.n13 source.n12 43.1397
R70 source.n26 source.n25 43.1396
R71 source.n24 source.n23 43.1396
R72 source.n22 source.n21 43.1396
R73 source.n19 source.n18 43.1396
R74 source.n17 source.n16 43.1396
R75 source.n15 source.n14 43.1396
R76 source.n15 source.n13 28.7794
R77 source.n28 source.n0 22.4432
R78 source.n28 source.n27 5.62119
R79 source.n25 source.t10 0.9905
R80 source.n25 source.t12 0.9905
R81 source.n23 source.t4 0.9905
R82 source.n23 source.t6 0.9905
R83 source.n21 source.t13 0.9905
R84 source.n21 source.t0 0.9905
R85 source.n18 source.t18 0.9905
R86 source.n18 source.t22 0.9905
R87 source.n16 source.t14 0.9905
R88 source.n16 source.t25 0.9905
R89 source.n14 source.t24 0.9905
R90 source.n14 source.t16 0.9905
R91 source.n1 source.t27 0.9905
R92 source.n1 source.t21 0.9905
R93 source.n3 source.t15 0.9905
R94 source.n3 source.t20 0.9905
R95 source.n5 source.t17 0.9905
R96 source.n5 source.t23 0.9905
R97 source.n8 source.t7 0.9905
R98 source.n8 source.t9 0.9905
R99 source.n10 source.t2 0.9905
R100 source.n10 source.t1 0.9905
R101 source.n12 source.t3 0.9905
R102 source.n12 source.t5 0.9905
R103 source.n7 source.n6 0.828086
R104 source.n22 source.n20 0.828086
R105 source.n13 source.n11 0.716017
R106 source.n11 source.n9 0.716017
R107 source.n9 source.n7 0.716017
R108 source.n6 source.n4 0.716017
R109 source.n4 source.n2 0.716017
R110 source.n2 source.n0 0.716017
R111 source.n17 source.n15 0.716017
R112 source.n19 source.n17 0.716017
R113 source.n20 source.n19 0.716017
R114 source.n24 source.n22 0.716017
R115 source.n26 source.n24 0.716017
R116 source.n27 source.n26 0.716017
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t9 61.5239
R119 drain_left.n1 drain_left.t7 61.5238
R120 drain_left.n4 drain_left.n2 60.5339
R121 drain_left.n11 drain_left.n10 59.8185
R122 drain_left.n9 drain_left.n8 59.8185
R123 drain_left.n7 drain_left.n6 59.8185
R124 drain_left.n4 drain_left.n3 59.8184
R125 drain_left.n1 drain_left.n0 59.8184
R126 drain_left drain_left.n5 37.5419
R127 drain_left drain_left.n11 6.36873
R128 drain_left.n2 drain_left.t12 0.9905
R129 drain_left.n2 drain_left.t13 0.9905
R130 drain_left.n3 drain_left.t11 0.9905
R131 drain_left.n3 drain_left.t6 0.9905
R132 drain_left.n0 drain_left.t4 0.9905
R133 drain_left.n0 drain_left.t10 0.9905
R134 drain_left.n10 drain_left.t0 0.9905
R135 drain_left.n10 drain_left.t5 0.9905
R136 drain_left.n8 drain_left.t8 0.9905
R137 drain_left.n8 drain_left.t2 0.9905
R138 drain_left.n6 drain_left.t3 0.9905
R139 drain_left.n6 drain_left.t1 0.9905
R140 drain_left.n9 drain_left.n7 0.716017
R141 drain_left.n11 drain_left.n9 0.716017
R142 drain_left.n5 drain_left.n1 0.481792
R143 drain_left.n5 drain_left.n4 0.124033
R144 minus.n4 minus.t9 1063.55
R145 minus.n20 minus.t3 1063.55
R146 minus.n3 minus.t1 1042.57
R147 minus.n7 minus.t5 1042.57
R148 minus.n8 minus.t13 1042.57
R149 minus.n1 minus.t4 1042.57
R150 minus.n13 minus.t7 1042.57
R151 minus.n14 minus.t0 1042.57
R152 minus.n19 minus.t2 1042.57
R153 minus.n23 minus.t10 1042.57
R154 minus.n24 minus.t8 1042.57
R155 minus.n17 minus.t6 1042.57
R156 minus.n29 minus.t12 1042.57
R157 minus.n30 minus.t11 1042.57
R158 minus.n15 minus.n14 161.3
R159 minus.n13 minus.n0 161.3
R160 minus.n12 minus.n11 161.3
R161 minus.n10 minus.n1 161.3
R162 minus.n7 minus.n2 161.3
R163 minus.n6 minus.n5 161.3
R164 minus.n31 minus.n30 161.3
R165 minus.n29 minus.n16 161.3
R166 minus.n28 minus.n27 161.3
R167 minus.n26 minus.n17 161.3
R168 minus.n23 minus.n18 161.3
R169 minus.n22 minus.n21 161.3
R170 minus.n9 minus.n8 80.6037
R171 minus.n25 minus.n24 80.6037
R172 minus.n5 minus.n4 70.4033
R173 minus.n21 minus.n20 70.4033
R174 minus.n8 minus.n7 48.2005
R175 minus.n8 minus.n1 48.2005
R176 minus.n14 minus.n13 48.2005
R177 minus.n24 minus.n23 48.2005
R178 minus.n24 minus.n17 48.2005
R179 minus.n30 minus.n29 48.2005
R180 minus.n32 minus.n15 43.0175
R181 minus.n7 minus.n6 24.8308
R182 minus.n12 minus.n1 24.8308
R183 minus.n23 minus.n22 24.8308
R184 minus.n28 minus.n17 24.8308
R185 minus.n6 minus.n3 23.3702
R186 minus.n13 minus.n12 23.3702
R187 minus.n22 minus.n19 23.3702
R188 minus.n29 minus.n28 23.3702
R189 minus.n4 minus.n3 20.9576
R190 minus.n20 minus.n19 20.9576
R191 minus.n32 minus.n31 6.5933
R192 minus.n10 minus.n9 0.285035
R193 minus.n9 minus.n2 0.285035
R194 minus.n25 minus.n18 0.285035
R195 minus.n26 minus.n25 0.285035
R196 minus.n15 minus.n0 0.189894
R197 minus.n11 minus.n0 0.189894
R198 minus.n11 minus.n10 0.189894
R199 minus.n5 minus.n2 0.189894
R200 minus.n21 minus.n18 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n16 0.189894
R203 minus.n31 minus.n16 0.189894
R204 minus minus.n32 0.188
R205 drain_right.n1 drain_right.t10 61.5238
R206 drain_right.n11 drain_right.t13 60.8084
R207 drain_right.n8 drain_right.n6 60.534
R208 drain_right.n4 drain_right.n2 60.5339
R209 drain_right.n8 drain_right.n7 59.8185
R210 drain_right.n10 drain_right.n9 59.8185
R211 drain_right.n4 drain_right.n3 59.8184
R212 drain_right.n1 drain_right.n0 59.8184
R213 drain_right drain_right.n5 36.9887
R214 drain_right drain_right.n11 6.01097
R215 drain_right.n2 drain_right.t1 0.9905
R216 drain_right.n2 drain_right.t2 0.9905
R217 drain_right.n3 drain_right.t5 0.9905
R218 drain_right.n3 drain_right.t7 0.9905
R219 drain_right.n0 drain_right.t11 0.9905
R220 drain_right.n0 drain_right.t3 0.9905
R221 drain_right.n6 drain_right.t12 0.9905
R222 drain_right.n6 drain_right.t4 0.9905
R223 drain_right.n7 drain_right.t0 0.9905
R224 drain_right.n7 drain_right.t8 0.9905
R225 drain_right.n9 drain_right.t6 0.9905
R226 drain_right.n9 drain_right.t9 0.9905
R227 drain_right.n11 drain_right.n10 0.716017
R228 drain_right.n10 drain_right.n8 0.716017
R229 drain_right.n5 drain_right.n1 0.481792
R230 drain_right.n5 drain_right.n4 0.124033
C0 drain_left drain_right 1.06216f
C1 source drain_right 34.5693f
C2 minus drain_right 12.036099f
C3 plus drain_right 0.35873f
C4 source drain_left 34.5834f
C5 minus drain_left 0.172393f
C6 drain_left plus 12.2317f
C7 source minus 11.550099f
C8 source plus 11.5651f
C9 minus plus 7.17731f
C10 drain_right a_n2044_n4888# 9.63162f
C11 drain_left a_n2044_n4888# 9.94373f
C12 source a_n2044_n4888# 9.273215f
C13 minus a_n2044_n4888# 8.578952f
C14 plus a_n2044_n4888# 10.886609f
C15 drain_right.t10 a_n2044_n4888# 4.95966f
C16 drain_right.t11 a_n2044_n4888# 0.423803f
C17 drain_right.t3 a_n2044_n4888# 0.423803f
C18 drain_right.n0 a_n2044_n4888# 3.8745f
C19 drain_right.n1 a_n2044_n4888# 0.700554f
C20 drain_right.t1 a_n2044_n4888# 0.423803f
C21 drain_right.t2 a_n2044_n4888# 0.423803f
C22 drain_right.n2 a_n2044_n4888# 3.87876f
C23 drain_right.t5 a_n2044_n4888# 0.423803f
C24 drain_right.t7 a_n2044_n4888# 0.423803f
C25 drain_right.n3 a_n2044_n4888# 3.8745f
C26 drain_right.n4 a_n2044_n4888# 0.660277f
C27 drain_right.n5 a_n2044_n4888# 1.85029f
C28 drain_right.t12 a_n2044_n4888# 0.423803f
C29 drain_right.t4 a_n2044_n4888# 0.423803f
C30 drain_right.n6 a_n2044_n4888# 3.87876f
C31 drain_right.t0 a_n2044_n4888# 0.423803f
C32 drain_right.t8 a_n2044_n4888# 0.423803f
C33 drain_right.n7 a_n2044_n4888# 3.87449f
C34 drain_right.n8 a_n2044_n4888# 0.706406f
C35 drain_right.t6 a_n2044_n4888# 0.423803f
C36 drain_right.t9 a_n2044_n4888# 0.423803f
C37 drain_right.n9 a_n2044_n4888# 3.87449f
C38 drain_right.n10 a_n2044_n4888# 0.349934f
C39 drain_right.t13 a_n2044_n4888# 4.95533f
C40 drain_right.n11 a_n2044_n4888# 0.609033f
C41 minus.n0 a_n2044_n4888# 0.045687f
C42 minus.t4 a_n2044_n4888# 1.29382f
C43 minus.n1 a_n2044_n4888# 0.490814f
C44 minus.n2 a_n2044_n4888# 0.060964f
C45 minus.t1 a_n2044_n4888# 1.29382f
C46 minus.n3 a_n2044_n4888# 0.490533f
C47 minus.t9 a_n2044_n4888# 1.30341f
C48 minus.n4 a_n2044_n4888# 0.476787f
C49 minus.n5 a_n2044_n4888# 0.150231f
C50 minus.n6 a_n2044_n4888# 0.010367f
C51 minus.t5 a_n2044_n4888# 1.29382f
C52 minus.n7 a_n2044_n4888# 0.490814f
C53 minus.t13 a_n2044_n4888# 1.29382f
C54 minus.n8 a_n2044_n4888# 0.496393f
C55 minus.n9 a_n2044_n4888# 0.060821f
C56 minus.n10 a_n2044_n4888# 0.060964f
C57 minus.n11 a_n2044_n4888# 0.045687f
C58 minus.n12 a_n2044_n4888# 0.010367f
C59 minus.t7 a_n2044_n4888# 1.29382f
C60 minus.n13 a_n2044_n4888# 0.490533f
C61 minus.t0 a_n2044_n4888# 1.29382f
C62 minus.n14 a_n2044_n4888# 0.486026f
C63 minus.n15 a_n2044_n4888# 2.09836f
C64 minus.n16 a_n2044_n4888# 0.045687f
C65 minus.t6 a_n2044_n4888# 1.29382f
C66 minus.n17 a_n2044_n4888# 0.490814f
C67 minus.n18 a_n2044_n4888# 0.060964f
C68 minus.t2 a_n2044_n4888# 1.29382f
C69 minus.n19 a_n2044_n4888# 0.490533f
C70 minus.t3 a_n2044_n4888# 1.30341f
C71 minus.n20 a_n2044_n4888# 0.476787f
C72 minus.n21 a_n2044_n4888# 0.150231f
C73 minus.n22 a_n2044_n4888# 0.010367f
C74 minus.t10 a_n2044_n4888# 1.29382f
C75 minus.n23 a_n2044_n4888# 0.490814f
C76 minus.t8 a_n2044_n4888# 1.29382f
C77 minus.n24 a_n2044_n4888# 0.496393f
C78 minus.n25 a_n2044_n4888# 0.060821f
C79 minus.n26 a_n2044_n4888# 0.060964f
C80 minus.n27 a_n2044_n4888# 0.045687f
C81 minus.n28 a_n2044_n4888# 0.010367f
C82 minus.t12 a_n2044_n4888# 1.29382f
C83 minus.n29 a_n2044_n4888# 0.490533f
C84 minus.t11 a_n2044_n4888# 1.29382f
C85 minus.n30 a_n2044_n4888# 0.486026f
C86 minus.n31 a_n2044_n4888# 0.308691f
C87 minus.n32 a_n2044_n4888# 2.49637f
C88 drain_left.t7 a_n2044_n4888# 4.969759f
C89 drain_left.t4 a_n2044_n4888# 0.424666f
C90 drain_left.t10 a_n2044_n4888# 0.424666f
C91 drain_left.n0 a_n2044_n4888# 3.88239f
C92 drain_left.n1 a_n2044_n4888# 0.701981f
C93 drain_left.t12 a_n2044_n4888# 0.424666f
C94 drain_left.t13 a_n2044_n4888# 0.424666f
C95 drain_left.n2 a_n2044_n4888# 3.88666f
C96 drain_left.t11 a_n2044_n4888# 0.424666f
C97 drain_left.t6 a_n2044_n4888# 0.424666f
C98 drain_left.n3 a_n2044_n4888# 3.88239f
C99 drain_left.n4 a_n2044_n4888# 0.661621f
C100 drain_left.n5 a_n2044_n4888# 1.90983f
C101 drain_left.t9 a_n2044_n4888# 4.96978f
C102 drain_left.t3 a_n2044_n4888# 0.424666f
C103 drain_left.t1 a_n2044_n4888# 0.424666f
C104 drain_left.n6 a_n2044_n4888# 3.88238f
C105 drain_left.n7 a_n2044_n4888# 0.720952f
C106 drain_left.t8 a_n2044_n4888# 0.424666f
C107 drain_left.t2 a_n2044_n4888# 0.424666f
C108 drain_left.n8 a_n2044_n4888# 3.88238f
C109 drain_left.n9 a_n2044_n4888# 0.350647f
C110 drain_left.t0 a_n2044_n4888# 0.424666f
C111 drain_left.t5 a_n2044_n4888# 0.424666f
C112 drain_left.n10 a_n2044_n4888# 3.88238f
C113 drain_left.n11 a_n2044_n4888# 0.581496f
C114 source.t26 a_n2044_n4888# 4.95671f
C115 source.n0 a_n2044_n4888# 2.13229f
C116 source.t27 a_n2044_n4888# 0.433719f
C117 source.t21 a_n2044_n4888# 0.433719f
C118 source.n1 a_n2044_n4888# 3.87764f
C119 source.n2 a_n2044_n4888# 0.408339f
C120 source.t15 a_n2044_n4888# 0.433719f
C121 source.t20 a_n2044_n4888# 0.433719f
C122 source.n3 a_n2044_n4888# 3.87764f
C123 source.n4 a_n2044_n4888# 0.408339f
C124 source.t17 a_n2044_n4888# 0.433719f
C125 source.t23 a_n2044_n4888# 0.433719f
C126 source.n5 a_n2044_n4888# 3.87764f
C127 source.n6 a_n2044_n4888# 0.418248f
C128 source.t11 a_n2044_n4888# 4.95672f
C129 source.n7 a_n2044_n4888# 0.522036f
C130 source.t7 a_n2044_n4888# 0.433719f
C131 source.t9 a_n2044_n4888# 0.433719f
C132 source.n8 a_n2044_n4888# 3.87764f
C133 source.n9 a_n2044_n4888# 0.408339f
C134 source.t2 a_n2044_n4888# 0.433719f
C135 source.t1 a_n2044_n4888# 0.433719f
C136 source.n10 a_n2044_n4888# 3.87764f
C137 source.n11 a_n2044_n4888# 0.408339f
C138 source.t3 a_n2044_n4888# 0.433719f
C139 source.t5 a_n2044_n4888# 0.433719f
C140 source.n12 a_n2044_n4888# 3.87764f
C141 source.n13 a_n2044_n4888# 2.58455f
C142 source.t24 a_n2044_n4888# 0.433719f
C143 source.t16 a_n2044_n4888# 0.433719f
C144 source.n14 a_n2044_n4888# 3.87764f
C145 source.n15 a_n2044_n4888# 2.58454f
C146 source.t14 a_n2044_n4888# 0.433719f
C147 source.t25 a_n2044_n4888# 0.433719f
C148 source.n16 a_n2044_n4888# 3.87764f
C149 source.n17 a_n2044_n4888# 0.408331f
C150 source.t18 a_n2044_n4888# 0.433719f
C151 source.t22 a_n2044_n4888# 0.433719f
C152 source.n18 a_n2044_n4888# 3.87764f
C153 source.n19 a_n2044_n4888# 0.408331f
C154 source.t19 a_n2044_n4888# 4.95669f
C155 source.n20 a_n2044_n4888# 0.522063f
C156 source.t13 a_n2044_n4888# 0.433719f
C157 source.t0 a_n2044_n4888# 0.433719f
C158 source.n21 a_n2044_n4888# 3.87764f
C159 source.n22 a_n2044_n4888# 0.418241f
C160 source.t4 a_n2044_n4888# 0.433719f
C161 source.t6 a_n2044_n4888# 0.433719f
C162 source.n23 a_n2044_n4888# 3.87764f
C163 source.n24 a_n2044_n4888# 0.408331f
C164 source.t10 a_n2044_n4888# 0.433719f
C165 source.t12 a_n2044_n4888# 0.433719f
C166 source.n25 a_n2044_n4888# 3.87764f
C167 source.n26 a_n2044_n4888# 0.408331f
C168 source.t8 a_n2044_n4888# 4.95669f
C169 source.n27 a_n2044_n4888# 0.657457f
C170 source.n28 a_n2044_n4888# 2.47994f
C171 plus.n0 a_n2044_n4888# 0.046122f
C172 plus.t8 a_n2044_n4888# 1.30614f
C173 plus.t13 a_n2044_n4888# 1.30614f
C174 plus.t11 a_n2044_n4888# 1.30614f
C175 plus.n1 a_n2044_n4888# 0.495488f
C176 plus.n2 a_n2044_n4888# 0.061545f
C177 plus.t5 a_n2044_n4888# 1.30614f
C178 plus.t12 a_n2044_n4888# 1.30614f
C179 plus.t10 a_n2044_n4888# 1.30614f
C180 plus.n3 a_n2044_n4888# 0.495203f
C181 plus.t4 a_n2044_n4888# 1.31582f
C182 plus.n4 a_n2044_n4888# 0.481327f
C183 plus.n5 a_n2044_n4888# 0.151662f
C184 plus.n6 a_n2044_n4888# 0.010466f
C185 plus.n7 a_n2044_n4888# 0.495488f
C186 plus.n8 a_n2044_n4888# 0.50112f
C187 plus.n9 a_n2044_n4888# 0.0614f
C188 plus.n10 a_n2044_n4888# 0.061545f
C189 plus.n11 a_n2044_n4888# 0.046122f
C190 plus.n12 a_n2044_n4888# 0.010466f
C191 plus.n13 a_n2044_n4888# 0.495203f
C192 plus.n14 a_n2044_n4888# 0.490654f
C193 plus.n15 a_n2044_n4888# 0.710218f
C194 plus.n16 a_n2044_n4888# 0.046122f
C195 plus.t6 a_n2044_n4888# 1.30614f
C196 plus.t9 a_n2044_n4888# 1.30614f
C197 plus.t3 a_n2044_n4888# 1.30614f
C198 plus.n17 a_n2044_n4888# 0.495488f
C199 plus.n18 a_n2044_n4888# 0.061545f
C200 plus.t2 a_n2044_n4888# 1.30614f
C201 plus.t7 a_n2044_n4888# 1.30614f
C202 plus.t1 a_n2044_n4888# 1.30614f
C203 plus.n19 a_n2044_n4888# 0.495203f
C204 plus.t0 a_n2044_n4888# 1.31582f
C205 plus.n20 a_n2044_n4888# 0.481327f
C206 plus.n21 a_n2044_n4888# 0.151662f
C207 plus.n22 a_n2044_n4888# 0.010466f
C208 plus.n23 a_n2044_n4888# 0.495488f
C209 plus.n24 a_n2044_n4888# 0.50112f
C210 plus.n25 a_n2044_n4888# 0.0614f
C211 plus.n26 a_n2044_n4888# 0.061545f
C212 plus.n27 a_n2044_n4888# 0.046122f
C213 plus.n28 a_n2044_n4888# 0.010466f
C214 plus.n29 a_n2044_n4888# 0.495203f
C215 plus.n30 a_n2044_n4888# 0.490654f
C216 plus.n31 a_n2044_n4888# 1.68231f
.ends

