* NGSPICE file created from diffpair117.ext - technology: sky130A

.subckt diffpair117 minus drain_right drain_left source plus
X0 a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X1 source.t31 minus.t0 drain_right.t13 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X2 source.t0 plus.t0 drain_left.t15 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X3 drain_left.t14 plus.t1 source.t14 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X4 source.t30 minus.t1 drain_right.t3 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 drain_right.t14 minus.t2 source.t29 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X6 a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X7 drain_right.t0 minus.t3 source.t28 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X8 drain_left.t13 plus.t2 source.t2 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X9 source.t9 plus.t3 drain_left.t12 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X10 drain_right.t4 minus.t4 source.t27 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X11 source.t26 minus.t5 drain_right.t6 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X12 drain_right.t10 minus.t6 source.t25 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X13 drain_left.t11 plus.t4 source.t11 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X14 source.t6 plus.t5 drain_left.t10 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 drain_left.t9 plus.t6 source.t15 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X16 source.t24 minus.t7 drain_right.t11 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 source.t7 plus.t7 drain_left.t8 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X18 source.t23 minus.t8 drain_right.t1 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X19 source.t10 plus.t8 drain_left.t7 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X20 drain_right.t7 minus.t9 source.t22 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X21 drain_left.t6 plus.t9 source.t12 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X22 a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X23 drain_right.t15 minus.t10 source.t21 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X24 drain_right.t2 minus.t11 source.t20 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X25 drain_left.t5 plus.t10 source.t4 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X26 source.t1 plus.t11 drain_left.t4 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X27 source.t19 minus.t12 drain_right.t12 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X28 source.t3 plus.t12 drain_left.t3 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X29 drain_right.t9 minus.t13 source.t18 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X30 a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X31 source.t17 minus.t14 drain_right.t5 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X32 source.t16 minus.t15 drain_right.t8 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X33 drain_left.t2 plus.t13 source.t5 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X34 source.t13 plus.t14 drain_left.t1 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X35 drain_left.t0 plus.t15 source.t8 a_n1850_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n21 minus.t15 295.043
R1 minus.n5 minus.t9 295.043
R2 minus.n44 minus.t4 295.043
R3 minus.n28 minus.t0 295.043
R4 minus.n20 minus.t6 265.101
R5 minus.n1 minus.t1 265.101
R6 minus.n14 minus.t13 265.101
R7 minus.n12 minus.t8 265.101
R8 minus.n3 minus.t2 265.101
R9 minus.n6 minus.t14 265.101
R10 minus.n43 minus.t5 265.101
R11 minus.n24 minus.t10 265.101
R12 minus.n37 minus.t12 265.101
R13 minus.n35 minus.t3 265.101
R14 minus.n26 minus.t7 265.101
R15 minus.n29 minus.t11 265.101
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 64.9975
R39 minus.n11 minus.n3 64.9975
R40 minus.n34 minus.n26 64.9975
R41 minus.n38 minus.n24 64.9975
R42 minus.n21 minus.n20 62.0763
R43 minus.n6 minus.n5 62.0763
R44 minus.n29 minus.n28 62.0763
R45 minus.n44 minus.n43 62.0763
R46 minus.n14 minus.n13 46.0096
R47 minus.n13 minus.n12 46.0096
R48 minus.n36 minus.n35 46.0096
R49 minus.n37 minus.n36 46.0096
R50 minus.n46 minus.n22 28.5194
R51 minus.n15 minus.n14 27.0217
R52 minus.n12 minus.n11 27.0217
R53 minus.n35 minus.n34 27.0217
R54 minus.n38 minus.n37 27.0217
R55 minus.n20 minus.n19 10.955
R56 minus.n7 minus.n6 10.955
R57 minus.n30 minus.n29 10.955
R58 minus.n43 minus.n42 10.955
R59 minus.n18 minus.n1 8.03383
R60 minus.n8 minus.n3 8.03383
R61 minus.n31 minus.n26 8.03383
R62 minus.n41 minus.n24 8.03383
R63 minus.n46 minus.n45 6.46641
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 drain_right.n9 drain_right.n7 101.338
R80 drain_right.n5 drain_right.n3 101.338
R81 drain_right.n2 drain_right.n0 101.338
R82 drain_right.n9 drain_right.n8 100.796
R83 drain_right.n11 drain_right.n10 100.796
R84 drain_right.n13 drain_right.n12 100.796
R85 drain_right.n5 drain_right.n4 100.796
R86 drain_right.n2 drain_right.n1 100.796
R87 drain_right drain_right.n6 22.7683
R88 drain_right.n3 drain_right.t6 9.9005
R89 drain_right.n3 drain_right.t4 9.9005
R90 drain_right.n4 drain_right.t12 9.9005
R91 drain_right.n4 drain_right.t15 9.9005
R92 drain_right.n1 drain_right.t11 9.9005
R93 drain_right.n1 drain_right.t0 9.9005
R94 drain_right.n0 drain_right.t13 9.9005
R95 drain_right.n0 drain_right.t2 9.9005
R96 drain_right.n7 drain_right.t5 9.9005
R97 drain_right.n7 drain_right.t7 9.9005
R98 drain_right.n8 drain_right.t1 9.9005
R99 drain_right.n8 drain_right.t14 9.9005
R100 drain_right.n10 drain_right.t3 9.9005
R101 drain_right.n10 drain_right.t9 9.9005
R102 drain_right.n12 drain_right.t8 9.9005
R103 drain_right.n12 drain_right.t10 9.9005
R104 drain_right drain_right.n13 6.19632
R105 drain_right.n13 drain_right.n11 0.543603
R106 drain_right.n11 drain_right.n9 0.543603
R107 drain_right.n6 drain_right.n5 0.216706
R108 drain_right.n6 drain_right.n2 0.216706
R109 source.n82 source.n80 289.615
R110 source.n68 source.n66 289.615
R111 source.n60 source.n58 289.615
R112 source.n46 source.n44 289.615
R113 source.n2 source.n0 289.615
R114 source.n16 source.n14 289.615
R115 source.n24 source.n22 289.615
R116 source.n38 source.n36 289.615
R117 source.n83 source.n82 185
R118 source.n69 source.n68 185
R119 source.n61 source.n60 185
R120 source.n47 source.n46 185
R121 source.n3 source.n2 185
R122 source.n17 source.n16 185
R123 source.n25 source.n24 185
R124 source.n39 source.n38 185
R125 source.t27 source.n81 167.117
R126 source.t31 source.n67 167.117
R127 source.t5 source.n59 167.117
R128 source.t3 source.n45 167.117
R129 source.t14 source.n1 167.117
R130 source.t9 source.n15 167.117
R131 source.t22 source.n23 167.117
R132 source.t16 source.n37 167.117
R133 source.n9 source.n8 84.1169
R134 source.n11 source.n10 84.1169
R135 source.n13 source.n12 84.1169
R136 source.n31 source.n30 84.1169
R137 source.n33 source.n32 84.1169
R138 source.n35 source.n34 84.1169
R139 source.n79 source.n78 84.1168
R140 source.n77 source.n76 84.1168
R141 source.n75 source.n74 84.1168
R142 source.n57 source.n56 84.1168
R143 source.n55 source.n54 84.1168
R144 source.n53 source.n52 84.1168
R145 source.n82 source.t27 52.3082
R146 source.n68 source.t31 52.3082
R147 source.n60 source.t5 52.3082
R148 source.n46 source.t3 52.3082
R149 source.n2 source.t14 52.3082
R150 source.n16 source.t9 52.3082
R151 source.n24 source.t22 52.3082
R152 source.n38 source.t16 52.3082
R153 source.n87 source.n86 31.4096
R154 source.n73 source.n72 31.4096
R155 source.n65 source.n64 31.4096
R156 source.n51 source.n50 31.4096
R157 source.n7 source.n6 31.4096
R158 source.n21 source.n20 31.4096
R159 source.n29 source.n28 31.4096
R160 source.n43 source.n42 31.4096
R161 source.n51 source.n43 14.2551
R162 source.n78 source.t21 9.9005
R163 source.n78 source.t26 9.9005
R164 source.n76 source.t28 9.9005
R165 source.n76 source.t19 9.9005
R166 source.n74 source.t20 9.9005
R167 source.n74 source.t24 9.9005
R168 source.n56 source.t11 9.9005
R169 source.n56 source.t7 9.9005
R170 source.n54 source.t4 9.9005
R171 source.n54 source.t0 9.9005
R172 source.n52 source.t2 9.9005
R173 source.n52 source.t10 9.9005
R174 source.n8 source.t12 9.9005
R175 source.n8 source.t13 9.9005
R176 source.n10 source.t8 9.9005
R177 source.n10 source.t6 9.9005
R178 source.n12 source.t15 9.9005
R179 source.n12 source.t1 9.9005
R180 source.n30 source.t29 9.9005
R181 source.n30 source.t17 9.9005
R182 source.n32 source.t18 9.9005
R183 source.n32 source.t23 9.9005
R184 source.n34 source.t25 9.9005
R185 source.n34 source.t30 9.9005
R186 source.n83 source.n81 9.71174
R187 source.n69 source.n67 9.71174
R188 source.n61 source.n59 9.71174
R189 source.n47 source.n45 9.71174
R190 source.n3 source.n1 9.71174
R191 source.n17 source.n15 9.71174
R192 source.n25 source.n23 9.71174
R193 source.n39 source.n37 9.71174
R194 source.n86 source.n85 9.45567
R195 source.n72 source.n71 9.45567
R196 source.n64 source.n63 9.45567
R197 source.n50 source.n49 9.45567
R198 source.n6 source.n5 9.45567
R199 source.n20 source.n19 9.45567
R200 source.n28 source.n27 9.45567
R201 source.n42 source.n41 9.45567
R202 source.n85 source.n84 9.3005
R203 source.n71 source.n70 9.3005
R204 source.n63 source.n62 9.3005
R205 source.n49 source.n48 9.3005
R206 source.n5 source.n4 9.3005
R207 source.n19 source.n18 9.3005
R208 source.n27 source.n26 9.3005
R209 source.n41 source.n40 9.3005
R210 source.n88 source.n7 8.72059
R211 source.n86 source.n80 8.14595
R212 source.n72 source.n66 8.14595
R213 source.n64 source.n58 8.14595
R214 source.n50 source.n44 8.14595
R215 source.n6 source.n0 8.14595
R216 source.n20 source.n14 8.14595
R217 source.n28 source.n22 8.14595
R218 source.n42 source.n36 8.14595
R219 source.n84 source.n83 7.3702
R220 source.n70 source.n69 7.3702
R221 source.n62 source.n61 7.3702
R222 source.n48 source.n47 7.3702
R223 source.n4 source.n3 7.3702
R224 source.n18 source.n17 7.3702
R225 source.n26 source.n25 7.3702
R226 source.n40 source.n39 7.3702
R227 source.n84 source.n80 5.81868
R228 source.n70 source.n66 5.81868
R229 source.n62 source.n58 5.81868
R230 source.n48 source.n44 5.81868
R231 source.n4 source.n0 5.81868
R232 source.n18 source.n14 5.81868
R233 source.n26 source.n22 5.81868
R234 source.n40 source.n36 5.81868
R235 source.n88 source.n87 5.53498
R236 source.n85 source.n81 3.44771
R237 source.n71 source.n67 3.44771
R238 source.n63 source.n59 3.44771
R239 source.n49 source.n45 3.44771
R240 source.n5 source.n1 3.44771
R241 source.n19 source.n15 3.44771
R242 source.n27 source.n23 3.44771
R243 source.n41 source.n37 3.44771
R244 source.n43 source.n35 0.543603
R245 source.n35 source.n33 0.543603
R246 source.n33 source.n31 0.543603
R247 source.n31 source.n29 0.543603
R248 source.n21 source.n13 0.543603
R249 source.n13 source.n11 0.543603
R250 source.n11 source.n9 0.543603
R251 source.n9 source.n7 0.543603
R252 source.n53 source.n51 0.543603
R253 source.n55 source.n53 0.543603
R254 source.n57 source.n55 0.543603
R255 source.n65 source.n57 0.543603
R256 source.n75 source.n73 0.543603
R257 source.n77 source.n75 0.543603
R258 source.n79 source.n77 0.543603
R259 source.n87 source.n79 0.543603
R260 source.n29 source.n21 0.470328
R261 source.n73 source.n65 0.470328
R262 source source.n88 0.188
R263 plus.n5 plus.t3 295.043
R264 plus.n21 plus.t1 295.043
R265 plus.n28 plus.t13 295.043
R266 plus.n44 plus.t12 295.043
R267 plus.n6 plus.t6 265.101
R268 plus.n3 plus.t11 265.101
R269 plus.n12 plus.t15 265.101
R270 plus.n14 plus.t5 265.101
R271 plus.n1 plus.t9 265.101
R272 plus.n20 plus.t14 265.101
R273 plus.n29 plus.t7 265.101
R274 plus.n26 plus.t4 265.101
R275 plus.n35 plus.t0 265.101
R276 plus.n37 plus.t10 265.101
R277 plus.n24 plus.t8 265.101
R278 plus.n43 plus.t2 265.101
R279 plus.n5 plus.n4 161.489
R280 plus.n28 plus.n27 161.489
R281 plus.n7 plus.n4 161.3
R282 plus.n9 plus.n8 161.3
R283 plus.n11 plus.n10 161.3
R284 plus.n13 plus.n2 161.3
R285 plus.n16 plus.n15 161.3
R286 plus.n18 plus.n17 161.3
R287 plus.n19 plus.n0 161.3
R288 plus.n22 plus.n21 161.3
R289 plus.n30 plus.n27 161.3
R290 plus.n32 plus.n31 161.3
R291 plus.n34 plus.n33 161.3
R292 plus.n36 plus.n25 161.3
R293 plus.n39 plus.n38 161.3
R294 plus.n41 plus.n40 161.3
R295 plus.n42 plus.n23 161.3
R296 plus.n45 plus.n44 161.3
R297 plus.n8 plus.n7 73.0308
R298 plus.n19 plus.n18 73.0308
R299 plus.n42 plus.n41 73.0308
R300 plus.n31 plus.n30 73.0308
R301 plus.n11 plus.n3 64.9975
R302 plus.n15 plus.n1 64.9975
R303 plus.n38 plus.n24 64.9975
R304 plus.n34 plus.n26 64.9975
R305 plus.n6 plus.n5 62.0763
R306 plus.n21 plus.n20 62.0763
R307 plus.n44 plus.n43 62.0763
R308 plus.n29 plus.n28 62.0763
R309 plus.n13 plus.n12 46.0096
R310 plus.n14 plus.n13 46.0096
R311 plus.n37 plus.n36 46.0096
R312 plus.n36 plus.n35 46.0096
R313 plus.n12 plus.n11 27.0217
R314 plus.n15 plus.n14 27.0217
R315 plus.n38 plus.n37 27.0217
R316 plus.n35 plus.n34 27.0217
R317 plus plus.n45 26.1884
R318 plus.n7 plus.n6 10.955
R319 plus.n20 plus.n19 10.955
R320 plus.n43 plus.n42 10.955
R321 plus.n30 plus.n29 10.955
R322 plus plus.n22 8.32247
R323 plus.n8 plus.n3 8.03383
R324 plus.n18 plus.n1 8.03383
R325 plus.n41 plus.n24 8.03383
R326 plus.n31 plus.n26 8.03383
R327 plus.n9 plus.n4 0.189894
R328 plus.n10 plus.n9 0.189894
R329 plus.n10 plus.n2 0.189894
R330 plus.n16 plus.n2 0.189894
R331 plus.n17 plus.n16 0.189894
R332 plus.n17 plus.n0 0.189894
R333 plus.n22 plus.n0 0.189894
R334 plus.n45 plus.n23 0.189894
R335 plus.n40 plus.n23 0.189894
R336 plus.n40 plus.n39 0.189894
R337 plus.n39 plus.n25 0.189894
R338 plus.n33 plus.n25 0.189894
R339 plus.n33 plus.n32 0.189894
R340 plus.n32 plus.n27 0.189894
R341 drain_left.n9 drain_left.n7 101.338
R342 drain_left.n5 drain_left.n3 101.338
R343 drain_left.n2 drain_left.n0 101.338
R344 drain_left.n13 drain_left.n12 100.796
R345 drain_left.n11 drain_left.n10 100.796
R346 drain_left.n9 drain_left.n8 100.796
R347 drain_left.n5 drain_left.n4 100.796
R348 drain_left.n2 drain_left.n1 100.796
R349 drain_left drain_left.n6 23.3215
R350 drain_left.n3 drain_left.t8 9.9005
R351 drain_left.n3 drain_left.t2 9.9005
R352 drain_left.n4 drain_left.t15 9.9005
R353 drain_left.n4 drain_left.t11 9.9005
R354 drain_left.n1 drain_left.t7 9.9005
R355 drain_left.n1 drain_left.t5 9.9005
R356 drain_left.n0 drain_left.t3 9.9005
R357 drain_left.n0 drain_left.t13 9.9005
R358 drain_left.n12 drain_left.t1 9.9005
R359 drain_left.n12 drain_left.t14 9.9005
R360 drain_left.n10 drain_left.t10 9.9005
R361 drain_left.n10 drain_left.t6 9.9005
R362 drain_left.n8 drain_left.t4 9.9005
R363 drain_left.n8 drain_left.t0 9.9005
R364 drain_left.n7 drain_left.t12 9.9005
R365 drain_left.n7 drain_left.t9 9.9005
R366 drain_left drain_left.n13 6.19632
R367 drain_left.n11 drain_left.n9 0.543603
R368 drain_left.n13 drain_left.n11 0.543603
R369 drain_left.n6 drain_left.n5 0.216706
R370 drain_left.n6 drain_left.n2 0.216706
C0 drain_left drain_right 0.948737f
C1 plus source 1.64278f
C2 minus source 1.62881f
C3 plus minus 3.61913f
C4 drain_left source 7.431149f
C5 plus drain_left 1.59168f
C6 drain_left minus 0.177567f
C7 drain_right source 7.43139f
C8 plus drain_right 0.341004f
C9 drain_right minus 1.41201f
C10 drain_right a_n1850_n1288# 3.92919f
C11 drain_left a_n1850_n1288# 4.18098f
C12 source a_n1850_n1288# 3.113032f
C13 minus a_n1850_n1288# 6.426728f
C14 plus a_n1850_n1288# 7.02674f
C15 drain_left.t3 a_n1850_n1288# 0.040891f
C16 drain_left.t13 a_n1850_n1288# 0.040891f
C17 drain_left.n0 a_n1850_n1288# 0.258495f
C18 drain_left.t7 a_n1850_n1288# 0.040891f
C19 drain_left.t5 a_n1850_n1288# 0.040891f
C20 drain_left.n1 a_n1850_n1288# 0.256892f
C21 drain_left.n2 a_n1850_n1288# 0.561512f
C22 drain_left.t8 a_n1850_n1288# 0.040891f
C23 drain_left.t2 a_n1850_n1288# 0.040891f
C24 drain_left.n3 a_n1850_n1288# 0.258495f
C25 drain_left.t15 a_n1850_n1288# 0.040891f
C26 drain_left.t11 a_n1850_n1288# 0.040891f
C27 drain_left.n4 a_n1850_n1288# 0.256892f
C28 drain_left.n5 a_n1850_n1288# 0.561512f
C29 drain_left.n6 a_n1850_n1288# 0.739219f
C30 drain_left.t12 a_n1850_n1288# 0.040891f
C31 drain_left.t9 a_n1850_n1288# 0.040891f
C32 drain_left.n7 a_n1850_n1288# 0.258496f
C33 drain_left.t4 a_n1850_n1288# 0.040891f
C34 drain_left.t0 a_n1850_n1288# 0.040891f
C35 drain_left.n8 a_n1850_n1288# 0.256893f
C36 drain_left.n9 a_n1850_n1288# 0.585989f
C37 drain_left.t10 a_n1850_n1288# 0.040891f
C38 drain_left.t6 a_n1850_n1288# 0.040891f
C39 drain_left.n10 a_n1850_n1288# 0.256893f
C40 drain_left.n11 a_n1850_n1288# 0.288585f
C41 drain_left.t1 a_n1850_n1288# 0.040891f
C42 drain_left.t14 a_n1850_n1288# 0.040891f
C43 drain_left.n12 a_n1850_n1288# 0.256893f
C44 drain_left.n13 a_n1850_n1288# 0.503943f
C45 plus.n0 a_n1850_n1288# 0.027758f
C46 plus.t14 a_n1850_n1288# 0.049008f
C47 plus.t9 a_n1850_n1288# 0.049008f
C48 plus.n1 a_n1850_n1288# 0.034228f
C49 plus.n2 a_n1850_n1288# 0.027758f
C50 plus.t5 a_n1850_n1288# 0.049008f
C51 plus.t15 a_n1850_n1288# 0.049008f
C52 plus.t11 a_n1850_n1288# 0.049008f
C53 plus.n3 a_n1850_n1288# 0.034228f
C54 plus.n4 a_n1850_n1288# 0.059073f
C55 plus.t6 a_n1850_n1288# 0.049008f
C56 plus.t3 a_n1850_n1288# 0.05249f
C57 plus.n5 a_n1850_n1288# 0.042301f
C58 plus.n6 a_n1850_n1288# 0.034228f
C59 plus.n7 a_n1850_n1288# 0.010492f
C60 plus.n8 a_n1850_n1288# 0.010149f
C61 plus.n9 a_n1850_n1288# 0.027758f
C62 plus.n10 a_n1850_n1288# 0.027758f
C63 plus.n11 a_n1850_n1288# 0.011433f
C64 plus.n12 a_n1850_n1288# 0.034228f
C65 plus.n13 a_n1850_n1288# 0.011433f
C66 plus.n14 a_n1850_n1288# 0.034228f
C67 plus.n15 a_n1850_n1288# 0.011433f
C68 plus.n16 a_n1850_n1288# 0.027758f
C69 plus.n17 a_n1850_n1288# 0.027758f
C70 plus.n18 a_n1850_n1288# 0.010149f
C71 plus.n19 a_n1850_n1288# 0.010492f
C72 plus.n20 a_n1850_n1288# 0.034228f
C73 plus.t1 a_n1850_n1288# 0.05249f
C74 plus.n21 a_n1850_n1288# 0.042264f
C75 plus.n22 a_n1850_n1288# 0.19612f
C76 plus.n23 a_n1850_n1288# 0.027758f
C77 plus.t12 a_n1850_n1288# 0.05249f
C78 plus.t2 a_n1850_n1288# 0.049008f
C79 plus.t8 a_n1850_n1288# 0.049008f
C80 plus.n24 a_n1850_n1288# 0.034228f
C81 plus.n25 a_n1850_n1288# 0.027758f
C82 plus.t10 a_n1850_n1288# 0.049008f
C83 plus.t0 a_n1850_n1288# 0.049008f
C84 plus.t4 a_n1850_n1288# 0.049008f
C85 plus.n26 a_n1850_n1288# 0.034228f
C86 plus.n27 a_n1850_n1288# 0.059073f
C87 plus.t7 a_n1850_n1288# 0.049008f
C88 plus.t13 a_n1850_n1288# 0.05249f
C89 plus.n28 a_n1850_n1288# 0.042301f
C90 plus.n29 a_n1850_n1288# 0.034228f
C91 plus.n30 a_n1850_n1288# 0.010492f
C92 plus.n31 a_n1850_n1288# 0.010149f
C93 plus.n32 a_n1850_n1288# 0.027758f
C94 plus.n33 a_n1850_n1288# 0.027758f
C95 plus.n34 a_n1850_n1288# 0.011433f
C96 plus.n35 a_n1850_n1288# 0.034228f
C97 plus.n36 a_n1850_n1288# 0.011433f
C98 plus.n37 a_n1850_n1288# 0.034228f
C99 plus.n38 a_n1850_n1288# 0.011433f
C100 plus.n39 a_n1850_n1288# 0.027758f
C101 plus.n40 a_n1850_n1288# 0.027758f
C102 plus.n41 a_n1850_n1288# 0.010149f
C103 plus.n42 a_n1850_n1288# 0.010492f
C104 plus.n43 a_n1850_n1288# 0.034228f
C105 plus.n44 a_n1850_n1288# 0.042264f
C106 plus.n45 a_n1850_n1288# 0.630642f
C107 source.n0 a_n1850_n1288# 0.039366f
C108 source.n1 a_n1850_n1288# 0.087103f
C109 source.t14 a_n1850_n1288# 0.065366f
C110 source.n2 a_n1850_n1288# 0.06817f
C111 source.n3 a_n1850_n1288# 0.021976f
C112 source.n4 a_n1850_n1288# 0.014493f
C113 source.n5 a_n1850_n1288# 0.191996f
C114 source.n6 a_n1850_n1288# 0.043155f
C115 source.n7 a_n1850_n1288# 0.407224f
C116 source.t12 a_n1850_n1288# 0.042627f
C117 source.t13 a_n1850_n1288# 0.042627f
C118 source.n8 a_n1850_n1288# 0.227884f
C119 source.n9 a_n1850_n1288# 0.30409f
C120 source.t8 a_n1850_n1288# 0.042627f
C121 source.t6 a_n1850_n1288# 0.042627f
C122 source.n10 a_n1850_n1288# 0.227884f
C123 source.n11 a_n1850_n1288# 0.30409f
C124 source.t15 a_n1850_n1288# 0.042627f
C125 source.t1 a_n1850_n1288# 0.042627f
C126 source.n12 a_n1850_n1288# 0.227884f
C127 source.n13 a_n1850_n1288# 0.30409f
C128 source.n14 a_n1850_n1288# 0.039366f
C129 source.n15 a_n1850_n1288# 0.087103f
C130 source.t9 a_n1850_n1288# 0.065366f
C131 source.n16 a_n1850_n1288# 0.06817f
C132 source.n17 a_n1850_n1288# 0.021976f
C133 source.n18 a_n1850_n1288# 0.014493f
C134 source.n19 a_n1850_n1288# 0.191996f
C135 source.n20 a_n1850_n1288# 0.043155f
C136 source.n21 a_n1850_n1288# 0.110236f
C137 source.n22 a_n1850_n1288# 0.039366f
C138 source.n23 a_n1850_n1288# 0.087103f
C139 source.t22 a_n1850_n1288# 0.065366f
C140 source.n24 a_n1850_n1288# 0.06817f
C141 source.n25 a_n1850_n1288# 0.021976f
C142 source.n26 a_n1850_n1288# 0.014493f
C143 source.n27 a_n1850_n1288# 0.191996f
C144 source.n28 a_n1850_n1288# 0.043155f
C145 source.n29 a_n1850_n1288# 0.110236f
C146 source.t29 a_n1850_n1288# 0.042627f
C147 source.t17 a_n1850_n1288# 0.042627f
C148 source.n30 a_n1850_n1288# 0.227884f
C149 source.n31 a_n1850_n1288# 0.30409f
C150 source.t18 a_n1850_n1288# 0.042627f
C151 source.t23 a_n1850_n1288# 0.042627f
C152 source.n32 a_n1850_n1288# 0.227884f
C153 source.n33 a_n1850_n1288# 0.30409f
C154 source.t25 a_n1850_n1288# 0.042627f
C155 source.t30 a_n1850_n1288# 0.042627f
C156 source.n34 a_n1850_n1288# 0.227884f
C157 source.n35 a_n1850_n1288# 0.30409f
C158 source.n36 a_n1850_n1288# 0.039366f
C159 source.n37 a_n1850_n1288# 0.087103f
C160 source.t16 a_n1850_n1288# 0.065366f
C161 source.n38 a_n1850_n1288# 0.06817f
C162 source.n39 a_n1850_n1288# 0.021976f
C163 source.n40 a_n1850_n1288# 0.014493f
C164 source.n41 a_n1850_n1288# 0.191996f
C165 source.n42 a_n1850_n1288# 0.043155f
C166 source.n43 a_n1850_n1288# 0.658679f
C167 source.n44 a_n1850_n1288# 0.039366f
C168 source.n45 a_n1850_n1288# 0.087103f
C169 source.t3 a_n1850_n1288# 0.065366f
C170 source.n46 a_n1850_n1288# 0.06817f
C171 source.n47 a_n1850_n1288# 0.021976f
C172 source.n48 a_n1850_n1288# 0.014493f
C173 source.n49 a_n1850_n1288# 0.191996f
C174 source.n50 a_n1850_n1288# 0.043155f
C175 source.n51 a_n1850_n1288# 0.658679f
C176 source.t2 a_n1850_n1288# 0.042627f
C177 source.t10 a_n1850_n1288# 0.042627f
C178 source.n52 a_n1850_n1288# 0.227883f
C179 source.n53 a_n1850_n1288# 0.304092f
C180 source.t4 a_n1850_n1288# 0.042627f
C181 source.t0 a_n1850_n1288# 0.042627f
C182 source.n54 a_n1850_n1288# 0.227883f
C183 source.n55 a_n1850_n1288# 0.304092f
C184 source.t11 a_n1850_n1288# 0.042627f
C185 source.t7 a_n1850_n1288# 0.042627f
C186 source.n56 a_n1850_n1288# 0.227883f
C187 source.n57 a_n1850_n1288# 0.304092f
C188 source.n58 a_n1850_n1288# 0.039366f
C189 source.n59 a_n1850_n1288# 0.087103f
C190 source.t5 a_n1850_n1288# 0.065366f
C191 source.n60 a_n1850_n1288# 0.06817f
C192 source.n61 a_n1850_n1288# 0.021976f
C193 source.n62 a_n1850_n1288# 0.014493f
C194 source.n63 a_n1850_n1288# 0.191996f
C195 source.n64 a_n1850_n1288# 0.043155f
C196 source.n65 a_n1850_n1288# 0.110236f
C197 source.n66 a_n1850_n1288# 0.039366f
C198 source.n67 a_n1850_n1288# 0.087103f
C199 source.t31 a_n1850_n1288# 0.065366f
C200 source.n68 a_n1850_n1288# 0.06817f
C201 source.n69 a_n1850_n1288# 0.021976f
C202 source.n70 a_n1850_n1288# 0.014493f
C203 source.n71 a_n1850_n1288# 0.191996f
C204 source.n72 a_n1850_n1288# 0.043155f
C205 source.n73 a_n1850_n1288# 0.110236f
C206 source.t20 a_n1850_n1288# 0.042627f
C207 source.t24 a_n1850_n1288# 0.042627f
C208 source.n74 a_n1850_n1288# 0.227883f
C209 source.n75 a_n1850_n1288# 0.304092f
C210 source.t28 a_n1850_n1288# 0.042627f
C211 source.t19 a_n1850_n1288# 0.042627f
C212 source.n76 a_n1850_n1288# 0.227883f
C213 source.n77 a_n1850_n1288# 0.304092f
C214 source.t21 a_n1850_n1288# 0.042627f
C215 source.t26 a_n1850_n1288# 0.042627f
C216 source.n78 a_n1850_n1288# 0.227883f
C217 source.n79 a_n1850_n1288# 0.304092f
C218 source.n80 a_n1850_n1288# 0.039366f
C219 source.n81 a_n1850_n1288# 0.087103f
C220 source.t27 a_n1850_n1288# 0.065366f
C221 source.n82 a_n1850_n1288# 0.06817f
C222 source.n83 a_n1850_n1288# 0.021976f
C223 source.n84 a_n1850_n1288# 0.014493f
C224 source.n85 a_n1850_n1288# 0.191996f
C225 source.n86 a_n1850_n1288# 0.043155f
C226 source.n87 a_n1850_n1288# 0.262489f
C227 source.n88 a_n1850_n1288# 0.66683f
C228 drain_right.t13 a_n1850_n1288# 0.041458f
C229 drain_right.t2 a_n1850_n1288# 0.041458f
C230 drain_right.n0 a_n1850_n1288# 0.262079f
C231 drain_right.t11 a_n1850_n1288# 0.041458f
C232 drain_right.t0 a_n1850_n1288# 0.041458f
C233 drain_right.n1 a_n1850_n1288# 0.260455f
C234 drain_right.n2 a_n1850_n1288# 0.569299f
C235 drain_right.t6 a_n1850_n1288# 0.041458f
C236 drain_right.t4 a_n1850_n1288# 0.041458f
C237 drain_right.n3 a_n1850_n1288# 0.262079f
C238 drain_right.t12 a_n1850_n1288# 0.041458f
C239 drain_right.t15 a_n1850_n1288# 0.041458f
C240 drain_right.n4 a_n1850_n1288# 0.260455f
C241 drain_right.n5 a_n1850_n1288# 0.569299f
C242 drain_right.n6 a_n1850_n1288# 0.698085f
C243 drain_right.t5 a_n1850_n1288# 0.041458f
C244 drain_right.t7 a_n1850_n1288# 0.041458f
C245 drain_right.n7 a_n1850_n1288# 0.26208f
C246 drain_right.t1 a_n1850_n1288# 0.041458f
C247 drain_right.t14 a_n1850_n1288# 0.041458f
C248 drain_right.n8 a_n1850_n1288# 0.260456f
C249 drain_right.n9 a_n1850_n1288# 0.594115f
C250 drain_right.t3 a_n1850_n1288# 0.041458f
C251 drain_right.t9 a_n1850_n1288# 0.041458f
C252 drain_right.n10 a_n1850_n1288# 0.260456f
C253 drain_right.n11 a_n1850_n1288# 0.292587f
C254 drain_right.t8 a_n1850_n1288# 0.041458f
C255 drain_right.t10 a_n1850_n1288# 0.041458f
C256 drain_right.n12 a_n1850_n1288# 0.260456f
C257 drain_right.n13 a_n1850_n1288# 0.510931f
C258 minus.n0 a_n1850_n1288# 0.027332f
C259 minus.t15 a_n1850_n1288# 0.051684f
C260 minus.t6 a_n1850_n1288# 0.048255f
C261 minus.t1 a_n1850_n1288# 0.048255f
C262 minus.n1 a_n1850_n1288# 0.033702f
C263 minus.n2 a_n1850_n1288# 0.027332f
C264 minus.t13 a_n1850_n1288# 0.048255f
C265 minus.t8 a_n1850_n1288# 0.048255f
C266 minus.t2 a_n1850_n1288# 0.048255f
C267 minus.n3 a_n1850_n1288# 0.033702f
C268 minus.n4 a_n1850_n1288# 0.058166f
C269 minus.t14 a_n1850_n1288# 0.048255f
C270 minus.t9 a_n1850_n1288# 0.051684f
C271 minus.n5 a_n1850_n1288# 0.041651f
C272 minus.n6 a_n1850_n1288# 0.033702f
C273 minus.n7 a_n1850_n1288# 0.010331f
C274 minus.n8 a_n1850_n1288# 0.009994f
C275 minus.n9 a_n1850_n1288# 0.027332f
C276 minus.n10 a_n1850_n1288# 0.027332f
C277 minus.n11 a_n1850_n1288# 0.011257f
C278 minus.n12 a_n1850_n1288# 0.033702f
C279 minus.n13 a_n1850_n1288# 0.011257f
C280 minus.n14 a_n1850_n1288# 0.033702f
C281 minus.n15 a_n1850_n1288# 0.011257f
C282 minus.n16 a_n1850_n1288# 0.027332f
C283 minus.n17 a_n1850_n1288# 0.027332f
C284 minus.n18 a_n1850_n1288# 0.009994f
C285 minus.n19 a_n1850_n1288# 0.010331f
C286 minus.n20 a_n1850_n1288# 0.033702f
C287 minus.n21 a_n1850_n1288# 0.041615f
C288 minus.n22 a_n1850_n1288# 0.650503f
C289 minus.n23 a_n1850_n1288# 0.027332f
C290 minus.t5 a_n1850_n1288# 0.048255f
C291 minus.t10 a_n1850_n1288# 0.048255f
C292 minus.n24 a_n1850_n1288# 0.033702f
C293 minus.n25 a_n1850_n1288# 0.027332f
C294 minus.t12 a_n1850_n1288# 0.048255f
C295 minus.t3 a_n1850_n1288# 0.048255f
C296 minus.t7 a_n1850_n1288# 0.048255f
C297 minus.n26 a_n1850_n1288# 0.033702f
C298 minus.n27 a_n1850_n1288# 0.058166f
C299 minus.t11 a_n1850_n1288# 0.048255f
C300 minus.t0 a_n1850_n1288# 0.051684f
C301 minus.n28 a_n1850_n1288# 0.041651f
C302 minus.n29 a_n1850_n1288# 0.033702f
C303 minus.n30 a_n1850_n1288# 0.010331f
C304 minus.n31 a_n1850_n1288# 0.009994f
C305 minus.n32 a_n1850_n1288# 0.027332f
C306 minus.n33 a_n1850_n1288# 0.027332f
C307 minus.n34 a_n1850_n1288# 0.011257f
C308 minus.n35 a_n1850_n1288# 0.033702f
C309 minus.n36 a_n1850_n1288# 0.011257f
C310 minus.n37 a_n1850_n1288# 0.033702f
C311 minus.n38 a_n1850_n1288# 0.011257f
C312 minus.n39 a_n1850_n1288# 0.027332f
C313 minus.n40 a_n1850_n1288# 0.027332f
C314 minus.n41 a_n1850_n1288# 0.009994f
C315 minus.n42 a_n1850_n1288# 0.010331f
C316 minus.n43 a_n1850_n1288# 0.033702f
C317 minus.t4 a_n1850_n1288# 0.051684f
C318 minus.n44 a_n1850_n1288# 0.041615f
C319 minus.n45 a_n1850_n1288# 0.176521f
C320 minus.n46 a_n1850_n1288# 0.805114f
.ends

