* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t26 plus.t0 drain_left.t6 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 source.t6 minus.t0 drain_right.t13 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 source.t25 plus.t1 drain_left.t11 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X3 drain_right.t12 minus.t1 source.t8 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X4 a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X5 drain_left.t12 plus.t2 source.t24 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X6 a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X7 source.t2 minus.t2 drain_right.t11 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X8 a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X9 drain_left.t7 plus.t3 source.t23 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 drain_right.t10 minus.t3 source.t0 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X11 drain_right.t9 minus.t4 source.t1 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X12 a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X13 source.t3 minus.t5 drain_right.t8 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X14 source.t22 plus.t4 drain_left.t4 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X15 drain_right.t7 minus.t6 source.t10 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X16 drain_right.t6 minus.t7 source.t5 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 source.t12 minus.t8 drain_right.t5 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 drain_left.t8 plus.t5 source.t21 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X19 drain_left.t1 plus.t6 source.t20 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X20 drain_right.t4 minus.t9 source.t27 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X21 drain_right.t3 minus.t10 source.t4 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X22 source.t19 plus.t7 drain_left.t9 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 source.t9 minus.t11 drain_right.t2 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X24 source.t11 minus.t12 drain_right.t1 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X25 drain_left.t2 plus.t8 source.t18 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X26 drain_left.t3 plus.t9 source.t17 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X27 drain_left.t0 plus.t10 source.t16 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X28 source.t15 plus.t11 drain_left.t5 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X29 source.t14 plus.t12 drain_left.t10 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X30 drain_right.t0 minus.t13 source.t7 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X31 drain_left.t13 plus.t13 source.t13 a_n1756_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
R0 plus.n3 plus.t6 756.595
R1 plus.n15 plus.t8 756.595
R2 plus.n20 plus.t2 756.595
R3 plus.n32 plus.t10 756.595
R4 plus.n1 plus.t7 690.867
R5 plus.n4 plus.t12 690.867
R6 plus.n6 plus.t9 690.867
R7 plus.n12 plus.t13 690.867
R8 plus.n14 plus.t11 690.867
R9 plus.n18 plus.t4 690.867
R10 plus.n21 plus.t1 690.867
R11 plus.n23 plus.t5 690.867
R12 plus.n29 plus.t3 690.867
R13 plus.n31 plus.t0 690.867
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 51.1217
R33 plus.n13 plus.n12 51.1217
R34 plus.n30 plus.n29 51.1217
R35 plus.n23 plus.n22 51.1217
R36 plus.n5 plus.n4 43.8187
R37 plus.n14 plus.n13 43.8187
R38 plus.n31 plus.n30 43.8187
R39 plus.n22 plus.n21 43.8187
R40 plus.n4 plus.n3 29.2126
R41 plus.n15 plus.n14 29.2126
R42 plus.n32 plus.n31 29.2126
R43 plus.n21 plus.n20 29.2126
R44 plus plus.n33 26.3153
R45 plus.n7 plus.n6 21.9096
R46 plus.n12 plus.n11 21.9096
R47 plus.n29 plus.n28 21.9096
R48 plus.n24 plus.n23 21.9096
R49 plus plus.n16 8.80542
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t1 90.3335
R61 drain_left.n1 drain_left.t0 90.3333
R62 drain_left.n4 drain_left.n2 80.3334
R63 drain_left.n11 drain_left.n10 79.7731
R64 drain_left.n9 drain_left.n8 79.7731
R65 drain_left.n7 drain_left.n6 79.7731
R66 drain_left.n4 drain_left.n3 79.773
R67 drain_left.n1 drain_left.n0 79.773
R68 drain_left drain_left.n5 23.7709
R69 drain_left.n2 drain_left.t11 10.0005
R70 drain_left.n2 drain_left.t12 10.0005
R71 drain_left.n3 drain_left.t4 10.0005
R72 drain_left.n3 drain_left.t8 10.0005
R73 drain_left.n0 drain_left.t6 10.0005
R74 drain_left.n0 drain_left.t7 10.0005
R75 drain_left.n10 drain_left.t5 10.0005
R76 drain_left.n10 drain_left.t2 10.0005
R77 drain_left.n8 drain_left.t9 10.0005
R78 drain_left.n8 drain_left.t13 10.0005
R79 drain_left.n6 drain_left.t10 10.0005
R80 drain_left.n6 drain_left.t3 10.0005
R81 drain_left drain_left.n11 6.21356
R82 drain_left.n9 drain_left.n7 0.560845
R83 drain_left.n11 drain_left.n9 0.560845
R84 drain_left.n5 drain_left.n1 0.365413
R85 drain_left.n5 drain_left.n4 0.0852402
R86 source.n0 source.t18 73.0943
R87 source.n7 source.t10 73.0943
R88 source.n27 source.t8 73.0942
R89 source.n20 source.t24 73.0942
R90 source.n2 source.n1 63.0943
R91 source.n4 source.n3 63.0943
R92 source.n6 source.n5 63.0943
R93 source.n9 source.n8 63.0943
R94 source.n11 source.n10 63.0943
R95 source.n13 source.n12 63.0943
R96 source.n26 source.n25 63.0942
R97 source.n24 source.n23 63.0942
R98 source.n22 source.n21 63.0942
R99 source.n19 source.n18 63.0942
R100 source.n17 source.n16 63.0942
R101 source.n15 source.n14 63.0942
R102 source.n15 source.n13 15.5902
R103 source.n25 source.t0 10.0005
R104 source.n25 source.t2 10.0005
R105 source.n23 source.t7 10.0005
R106 source.n23 source.t11 10.0005
R107 source.n21 source.t1 10.0005
R108 source.n21 source.t6 10.0005
R109 source.n18 source.t21 10.0005
R110 source.n18 source.t25 10.0005
R111 source.n16 source.t23 10.0005
R112 source.n16 source.t22 10.0005
R113 source.n14 source.t16 10.0005
R114 source.n14 source.t26 10.0005
R115 source.n1 source.t13 10.0005
R116 source.n1 source.t15 10.0005
R117 source.n3 source.t17 10.0005
R118 source.n3 source.t19 10.0005
R119 source.n5 source.t20 10.0005
R120 source.n5 source.t14 10.0005
R121 source.n8 source.t27 10.0005
R122 source.n8 source.t3 10.0005
R123 source.n10 source.t5 10.0005
R124 source.n10 source.t12 10.0005
R125 source.n12 source.t4 10.0005
R126 source.n12 source.t9 10.0005
R127 source.n28 source.n0 9.48679
R128 source.n28 source.n27 5.5436
R129 source.n7 source.n6 0.7505
R130 source.n22 source.n20 0.7505
R131 source.n13 source.n11 0.560845
R132 source.n11 source.n9 0.560845
R133 source.n9 source.n7 0.560845
R134 source.n6 source.n4 0.560845
R135 source.n4 source.n2 0.560845
R136 source.n2 source.n0 0.560845
R137 source.n17 source.n15 0.560845
R138 source.n19 source.n17 0.560845
R139 source.n20 source.n19 0.560845
R140 source.n24 source.n22 0.560845
R141 source.n26 source.n24 0.560845
R142 source.n27 source.n26 0.560845
R143 source source.n28 0.188
R144 minus.n15 minus.t10 756.595
R145 minus.n3 minus.t6 756.595
R146 minus.n32 minus.t1 756.595
R147 minus.n20 minus.t4 756.595
R148 minus.n1 minus.t8 690.867
R149 minus.n14 minus.t11 690.867
R150 minus.n12 minus.t7 690.867
R151 minus.n6 minus.t9 690.867
R152 minus.n4 minus.t5 690.867
R153 minus.n18 minus.t12 690.867
R154 minus.n31 minus.t2 690.867
R155 minus.n29 minus.t3 690.867
R156 minus.n23 minus.t13 690.867
R157 minus.n21 minus.t0 690.867
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 51.1217
R177 minus.n6 minus.n5 51.1217
R178 minus.n23 minus.n22 51.1217
R179 minus.n30 minus.n29 51.1217
R180 minus.n14 minus.n13 43.8187
R181 minus.n5 minus.n4 43.8187
R182 minus.n22 minus.n21 43.8187
R183 minus.n31 minus.n30 43.8187
R184 minus.n15 minus.n14 29.2126
R185 minus.n4 minus.n3 29.2126
R186 minus.n21 minus.n20 29.2126
R187 minus.n32 minus.n31 29.2126
R188 minus.n34 minus.n16 29.0251
R189 minus.n12 minus.n11 21.9096
R190 minus.n7 minus.n6 21.9096
R191 minus.n24 minus.n23 21.9096
R192 minus.n29 minus.n28 21.9096
R193 minus.n34 minus.n33 6.57058
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t9 90.3333
R206 drain_right.n11 drain_right.t3 89.7731
R207 drain_right.n8 drain_right.n6 80.3335
R208 drain_right.n4 drain_right.n2 80.3334
R209 drain_right.n8 drain_right.n7 79.7731
R210 drain_right.n10 drain_right.n9 79.7731
R211 drain_right.n4 drain_right.n3 79.773
R212 drain_right.n1 drain_right.n0 79.773
R213 drain_right drain_right.n5 23.2176
R214 drain_right.n2 drain_right.t11 10.0005
R215 drain_right.n2 drain_right.t12 10.0005
R216 drain_right.n3 drain_right.t1 10.0005
R217 drain_right.n3 drain_right.t10 10.0005
R218 drain_right.n0 drain_right.t13 10.0005
R219 drain_right.n0 drain_right.t0 10.0005
R220 drain_right.n6 drain_right.t8 10.0005
R221 drain_right.n6 drain_right.t7 10.0005
R222 drain_right.n7 drain_right.t5 10.0005
R223 drain_right.n7 drain_right.t4 10.0005
R224 drain_right.n9 drain_right.t2 10.0005
R225 drain_right.n9 drain_right.t6 10.0005
R226 drain_right drain_right.n11 5.93339
R227 drain_right.n11 drain_right.n10 0.560845
R228 drain_right.n10 drain_right.n8 0.560845
R229 drain_right.n5 drain_right.n1 0.365413
R230 drain_right.n5 drain_right.n4 0.0852402
C0 drain_right drain_left 0.897783f
C1 drain_right source 9.169371f
C2 minus drain_left 0.176362f
C3 plus drain_left 1.3173f
C4 minus source 1.17314f
C5 plus source 1.1873f
C6 source drain_left 9.17242f
C7 drain_right minus 1.14795f
C8 drain_right plus 0.330156f
C9 plus minus 3.66412f
C10 drain_right a_n1756_n1488# 4.20341f
C11 drain_left a_n1756_n1488# 4.45387f
C12 source a_n1756_n1488# 3.00053f
C13 minus a_n1756_n1488# 5.740038f
C14 plus a_n1756_n1488# 6.547703f
C15 drain_right.t9 a_n1756_n1488# 0.550479f
C16 drain_right.t13 a_n1756_n1488# 0.083829f
C17 drain_right.t0 a_n1756_n1488# 0.083829f
C18 drain_right.n0 a_n1756_n1488# 0.456015f
C19 drain_right.n1 a_n1756_n1488# 0.552658f
C20 drain_right.t11 a_n1756_n1488# 0.083829f
C21 drain_right.t12 a_n1756_n1488# 0.083829f
C22 drain_right.n2 a_n1756_n1488# 0.457971f
C23 drain_right.t1 a_n1756_n1488# 0.083829f
C24 drain_right.t10 a_n1756_n1488# 0.083829f
C25 drain_right.n3 a_n1756_n1488# 0.456015f
C26 drain_right.n4 a_n1756_n1488# 0.520246f
C27 drain_right.n5 a_n1756_n1488# 0.637152f
C28 drain_right.t8 a_n1756_n1488# 0.083829f
C29 drain_right.t7 a_n1756_n1488# 0.083829f
C30 drain_right.n6 a_n1756_n1488# 0.457973f
C31 drain_right.t5 a_n1756_n1488# 0.083829f
C32 drain_right.t4 a_n1756_n1488# 0.083829f
C33 drain_right.n7 a_n1756_n1488# 0.456017f
C34 drain_right.n8 a_n1756_n1488# 0.549623f
C35 drain_right.t2 a_n1756_n1488# 0.083829f
C36 drain_right.t6 a_n1756_n1488# 0.083829f
C37 drain_right.n9 a_n1756_n1488# 0.456017f
C38 drain_right.n10 a_n1756_n1488# 0.27109f
C39 drain_right.t3 a_n1756_n1488# 0.548641f
C40 drain_right.n11 a_n1756_n1488# 0.492313f
C41 minus.n0 a_n1756_n1488# 0.033026f
C42 minus.t10 a_n1756_n1488# 0.045828f
C43 minus.t11 a_n1756_n1488# 0.043038f
C44 minus.t7 a_n1756_n1488# 0.043038f
C45 minus.t8 a_n1756_n1488# 0.043038f
C46 minus.n1 a_n1756_n1488# 0.041036f
C47 minus.n2 a_n1756_n1488# 0.0772f
C48 minus.t9 a_n1756_n1488# 0.043038f
C49 minus.t5 a_n1756_n1488# 0.043038f
C50 minus.t6 a_n1756_n1488# 0.045828f
C51 minus.n3 a_n1756_n1488# 0.043389f
C52 minus.n4 a_n1756_n1488# 0.03008f
C53 minus.n5 a_n1756_n1488# 0.01401f
C54 minus.n6 a_n1756_n1488# 0.03008f
C55 minus.n7 a_n1756_n1488# 0.01401f
C56 minus.n8 a_n1756_n1488# 0.033026f
C57 minus.n9 a_n1756_n1488# 0.033026f
C58 minus.n10 a_n1756_n1488# 0.033026f
C59 minus.n11 a_n1756_n1488# 0.01401f
C60 minus.n12 a_n1756_n1488# 0.03008f
C61 minus.n13 a_n1756_n1488# 0.01401f
C62 minus.n14 a_n1756_n1488# 0.03008f
C63 minus.n15 a_n1756_n1488# 0.043337f
C64 minus.n16 a_n1756_n1488# 0.813879f
C65 minus.n17 a_n1756_n1488# 0.033026f
C66 minus.t2 a_n1756_n1488# 0.043038f
C67 minus.t3 a_n1756_n1488# 0.043038f
C68 minus.t12 a_n1756_n1488# 0.043038f
C69 minus.n18 a_n1756_n1488# 0.041036f
C70 minus.n19 a_n1756_n1488# 0.0772f
C71 minus.t13 a_n1756_n1488# 0.043038f
C72 minus.t0 a_n1756_n1488# 0.043038f
C73 minus.t4 a_n1756_n1488# 0.045828f
C74 minus.n20 a_n1756_n1488# 0.043389f
C75 minus.n21 a_n1756_n1488# 0.03008f
C76 minus.n22 a_n1756_n1488# 0.01401f
C77 minus.n23 a_n1756_n1488# 0.03008f
C78 minus.n24 a_n1756_n1488# 0.01401f
C79 minus.n25 a_n1756_n1488# 0.033026f
C80 minus.n26 a_n1756_n1488# 0.033026f
C81 minus.n27 a_n1756_n1488# 0.033026f
C82 minus.n28 a_n1756_n1488# 0.01401f
C83 minus.n29 a_n1756_n1488# 0.03008f
C84 minus.n30 a_n1756_n1488# 0.01401f
C85 minus.n31 a_n1756_n1488# 0.03008f
C86 minus.t1 a_n1756_n1488# 0.045828f
C87 minus.n32 a_n1756_n1488# 0.043337f
C88 minus.n33 a_n1756_n1488# 0.22139f
C89 minus.n34 a_n1756_n1488# 1.00249f
C90 source.t18 a_n1756_n1488# 0.563911f
C91 source.n0 a_n1756_n1488# 0.744433f
C92 source.t13 a_n1756_n1488# 0.095744f
C93 source.t15 a_n1756_n1488# 0.095744f
C94 source.n1 a_n1756_n1488# 0.465773f
C95 source.n2 a_n1756_n1488# 0.328455f
C96 source.t17 a_n1756_n1488# 0.095744f
C97 source.t19 a_n1756_n1488# 0.095744f
C98 source.n3 a_n1756_n1488# 0.465773f
C99 source.n4 a_n1756_n1488# 0.328455f
C100 source.t20 a_n1756_n1488# 0.095744f
C101 source.t14 a_n1756_n1488# 0.095744f
C102 source.n5 a_n1756_n1488# 0.465773f
C103 source.n6 a_n1756_n1488# 0.344744f
C104 source.t10 a_n1756_n1488# 0.563911f
C105 source.n7 a_n1756_n1488# 0.418946f
C106 source.t27 a_n1756_n1488# 0.095744f
C107 source.t3 a_n1756_n1488# 0.095744f
C108 source.n8 a_n1756_n1488# 0.465773f
C109 source.n9 a_n1756_n1488# 0.328455f
C110 source.t5 a_n1756_n1488# 0.095744f
C111 source.t12 a_n1756_n1488# 0.095744f
C112 source.n10 a_n1756_n1488# 0.465773f
C113 source.n11 a_n1756_n1488# 0.328455f
C114 source.t4 a_n1756_n1488# 0.095744f
C115 source.t9 a_n1756_n1488# 0.095744f
C116 source.n12 a_n1756_n1488# 0.465773f
C117 source.n13 a_n1756_n1488# 0.996556f
C118 source.t16 a_n1756_n1488# 0.095744f
C119 source.t26 a_n1756_n1488# 0.095744f
C120 source.n14 a_n1756_n1488# 0.46577f
C121 source.n15 a_n1756_n1488# 0.996559f
C122 source.t23 a_n1756_n1488# 0.095744f
C123 source.t22 a_n1756_n1488# 0.095744f
C124 source.n16 a_n1756_n1488# 0.46577f
C125 source.n17 a_n1756_n1488# 0.328458f
C126 source.t21 a_n1756_n1488# 0.095744f
C127 source.t25 a_n1756_n1488# 0.095744f
C128 source.n18 a_n1756_n1488# 0.46577f
C129 source.n19 a_n1756_n1488# 0.328458f
C130 source.t24 a_n1756_n1488# 0.563908f
C131 source.n20 a_n1756_n1488# 0.418948f
C132 source.t1 a_n1756_n1488# 0.095744f
C133 source.t6 a_n1756_n1488# 0.095744f
C134 source.n21 a_n1756_n1488# 0.46577f
C135 source.n22 a_n1756_n1488# 0.344747f
C136 source.t7 a_n1756_n1488# 0.095744f
C137 source.t11 a_n1756_n1488# 0.095744f
C138 source.n23 a_n1756_n1488# 0.46577f
C139 source.n24 a_n1756_n1488# 0.328458f
C140 source.t0 a_n1756_n1488# 0.095744f
C141 source.t2 a_n1756_n1488# 0.095744f
C142 source.n25 a_n1756_n1488# 0.46577f
C143 source.n26 a_n1756_n1488# 0.328458f
C144 source.t8 a_n1756_n1488# 0.563908f
C145 source.n27 a_n1756_n1488# 0.546536f
C146 source.n28 a_n1756_n1488# 0.773255f
C147 drain_left.t0 a_n1756_n1488# 0.54507f
C148 drain_left.t6 a_n1756_n1488# 0.083005f
C149 drain_left.t7 a_n1756_n1488# 0.083005f
C150 drain_left.n0 a_n1756_n1488# 0.451534f
C151 drain_left.n1 a_n1756_n1488# 0.547228f
C152 drain_left.t11 a_n1756_n1488# 0.083005f
C153 drain_left.t12 a_n1756_n1488# 0.083005f
C154 drain_left.n2 a_n1756_n1488# 0.453471f
C155 drain_left.t4 a_n1756_n1488# 0.083005f
C156 drain_left.t8 a_n1756_n1488# 0.083005f
C157 drain_left.n3 a_n1756_n1488# 0.451534f
C158 drain_left.n4 a_n1756_n1488# 0.515134f
C159 drain_left.n5 a_n1756_n1488# 0.676727f
C160 drain_left.t1 a_n1756_n1488# 0.545072f
C161 drain_left.t10 a_n1756_n1488# 0.083005f
C162 drain_left.t3 a_n1756_n1488# 0.083005f
C163 drain_left.n6 a_n1756_n1488# 0.451536f
C164 drain_left.n7 a_n1756_n1488# 0.560308f
C165 drain_left.t9 a_n1756_n1488# 0.083005f
C166 drain_left.t13 a_n1756_n1488# 0.083005f
C167 drain_left.n8 a_n1756_n1488# 0.451536f
C168 drain_left.n9 a_n1756_n1488# 0.268426f
C169 drain_left.t5 a_n1756_n1488# 0.083005f
C170 drain_left.t2 a_n1756_n1488# 0.083005f
C171 drain_left.n10 a_n1756_n1488# 0.451536f
C172 drain_left.n11 a_n1756_n1488# 0.461407f
C173 plus.n0 a_n1756_n1488# 0.033633f
C174 plus.t11 a_n1756_n1488# 0.043829f
C175 plus.t13 a_n1756_n1488# 0.043829f
C176 plus.t7 a_n1756_n1488# 0.043829f
C177 plus.n1 a_n1756_n1488# 0.041791f
C178 plus.n2 a_n1756_n1488# 0.078619f
C179 plus.t9 a_n1756_n1488# 0.043829f
C180 plus.t12 a_n1756_n1488# 0.043829f
C181 plus.t6 a_n1756_n1488# 0.046671f
C182 plus.n3 a_n1756_n1488# 0.044186f
C183 plus.n4 a_n1756_n1488# 0.030633f
C184 plus.n5 a_n1756_n1488# 0.014268f
C185 plus.n6 a_n1756_n1488# 0.030633f
C186 plus.n7 a_n1756_n1488# 0.014268f
C187 plus.n8 a_n1756_n1488# 0.033633f
C188 plus.n9 a_n1756_n1488# 0.033633f
C189 plus.n10 a_n1756_n1488# 0.033633f
C190 plus.n11 a_n1756_n1488# 0.014268f
C191 plus.n12 a_n1756_n1488# 0.030633f
C192 plus.n13 a_n1756_n1488# 0.014268f
C193 plus.n14 a_n1756_n1488# 0.030633f
C194 plus.t8 a_n1756_n1488# 0.046671f
C195 plus.n15 a_n1756_n1488# 0.044133f
C196 plus.n16 a_n1756_n1488# 0.257106f
C197 plus.n17 a_n1756_n1488# 0.033633f
C198 plus.t10 a_n1756_n1488# 0.046671f
C199 plus.t0 a_n1756_n1488# 0.043829f
C200 plus.t3 a_n1756_n1488# 0.043829f
C201 plus.t4 a_n1756_n1488# 0.043829f
C202 plus.n18 a_n1756_n1488# 0.041791f
C203 plus.n19 a_n1756_n1488# 0.078619f
C204 plus.t5 a_n1756_n1488# 0.043829f
C205 plus.t1 a_n1756_n1488# 0.043829f
C206 plus.t2 a_n1756_n1488# 0.046671f
C207 plus.n20 a_n1756_n1488# 0.044186f
C208 plus.n21 a_n1756_n1488# 0.030633f
C209 plus.n22 a_n1756_n1488# 0.014268f
C210 plus.n23 a_n1756_n1488# 0.030633f
C211 plus.n24 a_n1756_n1488# 0.014268f
C212 plus.n25 a_n1756_n1488# 0.033633f
C213 plus.n26 a_n1756_n1488# 0.033633f
C214 plus.n27 a_n1756_n1488# 0.033633f
C215 plus.n28 a_n1756_n1488# 0.014268f
C216 plus.n29 a_n1756_n1488# 0.030633f
C217 plus.n30 a_n1756_n1488# 0.014268f
C218 plus.n31 a_n1756_n1488# 0.030633f
C219 plus.n32 a_n1756_n1488# 0.044133f
C220 plus.n33 a_n1756_n1488# 0.780365f
.ends

