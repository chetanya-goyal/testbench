* NGSPICE file created from diffpair516.ext - technology: sky130A

.subckt diffpair516 minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t10 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X1 drain_left.t13 plus.t0 source.t3 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X2 drain_left.t12 plus.t1 source.t8 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X3 drain_right.t8 minus.t1 source.t26 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X4 a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X5 drain_left.t11 plus.t2 source.t12 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X6 drain_right.t6 minus.t2 source.t25 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X7 drain_right.t4 minus.t3 source.t24 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X8 drain_right.t13 minus.t4 source.t23 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X9 a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X10 drain_left.t10 plus.t3 source.t2 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X11 drain_left.t9 plus.t4 source.t11 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X12 drain_left.t8 plus.t5 source.t4 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X13 source.t13 plus.t6 drain_left.t7 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X14 source.t22 minus.t5 drain_right.t1 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X15 drain_right.t3 minus.t6 source.t21 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X16 drain_right.t0 minus.t7 source.t20 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 drain_right.t11 minus.t8 source.t19 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X18 source.t1 plus.t7 drain_left.t6 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X19 source.t7 plus.t8 drain_left.t5 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X20 drain_left.t4 plus.t9 source.t10 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X21 source.t5 plus.t10 drain_left.t3 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X22 source.t6 plus.t11 drain_left.t2 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 drain_right.t9 minus.t9 source.t18 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X24 source.t17 minus.t10 drain_right.t7 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X25 source.t16 minus.t11 drain_right.t5 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X26 a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X27 source.t15 minus.t12 drain_right.t12 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X28 a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X29 drain_left.t1 plus.t12 source.t9 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X30 source.t14 minus.t13 drain_right.t2 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X31 source.t0 plus.t13 drain_left.t0 a_n1724_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 minus.n15 minus.t4 1366.4
R1 minus.n3 minus.t8 1366.4
R2 minus.n32 minus.t6 1366.4
R3 minus.n20 minus.t3 1366.4
R4 minus.n1 minus.t5 1309.43
R5 minus.n14 minus.t0 1309.43
R6 minus.n12 minus.t9 1309.43
R7 minus.n6 minus.t1 1309.43
R8 minus.n4 minus.t12 1309.43
R9 minus.n18 minus.t10 1309.43
R10 minus.n31 minus.t13 1309.43
R11 minus.n29 minus.t7 1309.43
R12 minus.n23 minus.t2 1309.43
R13 minus.n21 minus.t11 1309.43
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n34 minus.n16 37.9607
R41 minus.n15 minus.n14 35.055
R42 minus.n4 minus.n3 35.055
R43 minus.n21 minus.n20 35.055
R44 minus.n32 minus.n31 35.055
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n1 drain_right.t4 62.7427
R62 drain_right.n11 drain_right.t13 62.1998
R63 drain_right.n8 drain_right.n6 61.4227
R64 drain_right.n4 drain_right.n2 61.4227
R65 drain_right.n8 drain_right.n7 60.8798
R66 drain_right.n10 drain_right.n9 60.8798
R67 drain_right.n4 drain_right.n3 60.8796
R68 drain_right.n1 drain_right.n0 60.8796
R69 drain_right drain_right.n5 32.2094
R70 drain_right drain_right.n11 5.92477
R71 drain_right.n2 drain_right.t2 1.3205
R72 drain_right.n2 drain_right.t3 1.3205
R73 drain_right.n3 drain_right.t7 1.3205
R74 drain_right.n3 drain_right.t0 1.3205
R75 drain_right.n0 drain_right.t5 1.3205
R76 drain_right.n0 drain_right.t6 1.3205
R77 drain_right.n6 drain_right.t12 1.3205
R78 drain_right.n6 drain_right.t11 1.3205
R79 drain_right.n7 drain_right.t1 1.3205
R80 drain_right.n7 drain_right.t8 1.3205
R81 drain_right.n9 drain_right.t10 1.3205
R82 drain_right.n9 drain_right.t9 1.3205
R83 drain_right.n11 drain_right.n10 0.543603
R84 drain_right.n10 drain_right.n8 0.543603
R85 drain_right.n5 drain_right.n1 0.352482
R86 drain_right.n5 drain_right.n4 0.0809298
R87 source.n7 source.t19 45.521
R88 source.n27 source.t21 45.5208
R89 source.n20 source.t3 45.5208
R90 source.n0 source.t9 45.5208
R91 source.n2 source.n1 44.201
R92 source.n4 source.n3 44.201
R93 source.n6 source.n5 44.201
R94 source.n9 source.n8 44.201
R95 source.n11 source.n10 44.201
R96 source.n13 source.n12 44.201
R97 source.n26 source.n25 44.2008
R98 source.n24 source.n23 44.2008
R99 source.n22 source.n21 44.2008
R100 source.n19 source.n18 44.2008
R101 source.n17 source.n16 44.2008
R102 source.n15 source.n14 44.2008
R103 source.n15 source.n13 24.6467
R104 source.n28 source.n0 18.5691
R105 source.n28 source.n27 5.53498
R106 source.n25 source.t20 1.3205
R107 source.n25 source.t14 1.3205
R108 source.n23 source.t25 1.3205
R109 source.n23 source.t17 1.3205
R110 source.n21 source.t24 1.3205
R111 source.n21 source.t16 1.3205
R112 source.n18 source.t8 1.3205
R113 source.n18 source.t7 1.3205
R114 source.n16 source.t2 1.3205
R115 source.n16 source.t5 1.3205
R116 source.n14 source.t11 1.3205
R117 source.n14 source.t6 1.3205
R118 source.n1 source.t4 1.3205
R119 source.n1 source.t1 1.3205
R120 source.n3 source.t10 1.3205
R121 source.n3 source.t0 1.3205
R122 source.n5 source.t12 1.3205
R123 source.n5 source.t13 1.3205
R124 source.n8 source.t26 1.3205
R125 source.n8 source.t15 1.3205
R126 source.n10 source.t18 1.3205
R127 source.n10 source.t22 1.3205
R128 source.n12 source.t23 1.3205
R129 source.n12 source.t27 1.3205
R130 source.n7 source.n6 0.741879
R131 source.n22 source.n20 0.741879
R132 source.n13 source.n11 0.543603
R133 source.n11 source.n9 0.543603
R134 source.n9 source.n7 0.543603
R135 source.n6 source.n4 0.543603
R136 source.n4 source.n2 0.543603
R137 source.n2 source.n0 0.543603
R138 source.n17 source.n15 0.543603
R139 source.n19 source.n17 0.543603
R140 source.n20 source.n19 0.543603
R141 source.n24 source.n22 0.543603
R142 source.n26 source.n24 0.543603
R143 source.n27 source.n26 0.543603
R144 source source.n28 0.188
R145 plus.n3 plus.t2 1366.4
R146 plus.n15 plus.t12 1366.4
R147 plus.n20 plus.t0 1366.4
R148 plus.n32 plus.t4 1366.4
R149 plus.n1 plus.t13 1309.43
R150 plus.n4 plus.t6 1309.43
R151 plus.n6 plus.t9 1309.43
R152 plus.n12 plus.t5 1309.43
R153 plus.n14 plus.t7 1309.43
R154 plus.n18 plus.t10 1309.43
R155 plus.n21 plus.t8 1309.43
R156 plus.n23 plus.t1 1309.43
R157 plus.n29 plus.t3 1309.43
R158 plus.n31 plus.t11 1309.43
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 54.0429
R178 plus.n13 plus.n12 54.0429
R179 plus.n30 plus.n29 54.0429
R180 plus.n23 plus.n22 54.0429
R181 plus.n5 plus.n4 37.9763
R182 plus.n14 plus.n13 37.9763
R183 plus.n31 plus.n30 37.9763
R184 plus.n22 plus.n21 37.9763
R185 plus.n4 plus.n3 35.055
R186 plus.n15 plus.n14 35.055
R187 plus.n32 plus.n31 35.055
R188 plus.n21 plus.n20 35.055
R189 plus plus.n33 30.7055
R190 plus.n7 plus.n6 18.9884
R191 plus.n12 plus.n11 18.9884
R192 plus.n29 plus.n28 18.9884
R193 plus.n24 plus.n23 18.9884
R194 plus plus.n16 13.3168
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t11 62.7429
R206 drain_left.n1 drain_left.t9 62.7427
R207 drain_left.n4 drain_left.n2 61.4227
R208 drain_left.n9 drain_left.n8 60.8798
R209 drain_left.n7 drain_left.n6 60.8798
R210 drain_left.n11 drain_left.n10 60.8796
R211 drain_left.n4 drain_left.n3 60.8796
R212 drain_left.n1 drain_left.n0 60.8796
R213 drain_left drain_left.n5 32.7626
R214 drain_left drain_left.n11 6.19632
R215 drain_left.n2 drain_left.t5 1.3205
R216 drain_left.n2 drain_left.t13 1.3205
R217 drain_left.n3 drain_left.t3 1.3205
R218 drain_left.n3 drain_left.t12 1.3205
R219 drain_left.n0 drain_left.t2 1.3205
R220 drain_left.n0 drain_left.t10 1.3205
R221 drain_left.n10 drain_left.t6 1.3205
R222 drain_left.n10 drain_left.t1 1.3205
R223 drain_left.n8 drain_left.t0 1.3205
R224 drain_left.n8 drain_left.t8 1.3205
R225 drain_left.n6 drain_left.t7 1.3205
R226 drain_left.n6 drain_left.t4 1.3205
R227 drain_left.n9 drain_left.n7 0.543603
R228 drain_left.n11 drain_left.n9 0.543603
R229 drain_left.n5 drain_left.n1 0.352482
R230 drain_left.n5 drain_left.n4 0.0809298
C0 drain_right minus 6.46882f
C1 drain_right plus 0.323927f
C2 plus minus 5.85473f
C3 drain_right drain_left 0.884945f
C4 drain_right source 34.3437f
C5 minus drain_left 0.171678f
C6 plus drain_left 6.63194f
C7 minus source 6.00372f
C8 plus source 6.01858f
C9 source drain_left 34.3566f
C10 drain_right a_n1724_n3888# 8.275411f
C11 drain_left a_n1724_n3888# 8.556219f
C12 source a_n1724_n3888# 7.228034f
C13 minus a_n1724_n3888# 6.906449f
C14 plus a_n1724_n3888# 9.09209f
C15 drain_left.t9 a_n1724_n3888# 4.23319f
C16 drain_left.t2 a_n1724_n3888# 0.3666f
C17 drain_left.t10 a_n1724_n3888# 0.3666f
C18 drain_left.n0 a_n1724_n3888# 3.31364f
C19 drain_left.n1 a_n1724_n3888# 0.744718f
C20 drain_left.t5 a_n1724_n3888# 0.3666f
C21 drain_left.t13 a_n1724_n3888# 0.3666f
C22 drain_left.n2 a_n1724_n3888# 3.31694f
C23 drain_left.t3 a_n1724_n3888# 0.3666f
C24 drain_left.t12 a_n1724_n3888# 0.3666f
C25 drain_left.n3 a_n1724_n3888# 3.31364f
C26 drain_left.n4 a_n1724_n3888# 0.695083f
C27 drain_left.n5 a_n1724_n3888# 1.69151f
C28 drain_left.t11 a_n1724_n3888# 4.23319f
C29 drain_left.t7 a_n1724_n3888# 0.3666f
C30 drain_left.t4 a_n1724_n3888# 0.3666f
C31 drain_left.n6 a_n1724_n3888# 3.31364f
C32 drain_left.n7 a_n1724_n3888# 0.761722f
C33 drain_left.t0 a_n1724_n3888# 0.3666f
C34 drain_left.t8 a_n1724_n3888# 0.3666f
C35 drain_left.n8 a_n1724_n3888# 3.31364f
C36 drain_left.n9 a_n1724_n3888# 0.361561f
C37 drain_left.t6 a_n1724_n3888# 0.3666f
C38 drain_left.t1 a_n1724_n3888# 0.3666f
C39 drain_left.n10 a_n1724_n3888# 3.31363f
C40 drain_left.n11 a_n1724_n3888# 0.619003f
C41 plus.n0 a_n1724_n3888# 0.052244f
C42 plus.t7 a_n1724_n3888# 0.663254f
C43 plus.t5 a_n1724_n3888# 0.663254f
C44 plus.t13 a_n1724_n3888# 0.663254f
C45 plus.n1 a_n1724_n3888# 0.272091f
C46 plus.n2 a_n1724_n3888# 0.123088f
C47 plus.t9 a_n1724_n3888# 0.663254f
C48 plus.t6 a_n1724_n3888# 0.663254f
C49 plus.t2 a_n1724_n3888# 0.67413f
C50 plus.n3 a_n1724_n3888# 0.271606f
C51 plus.n4 a_n1724_n3888# 0.25476f
C52 plus.n5 a_n1724_n3888# 0.021519f
C53 plus.n6 a_n1724_n3888# 0.25476f
C54 plus.n7 a_n1724_n3888# 0.021519f
C55 plus.n8 a_n1724_n3888# 0.052244f
C56 plus.n9 a_n1724_n3888# 0.052244f
C57 plus.n10 a_n1724_n3888# 0.052244f
C58 plus.n11 a_n1724_n3888# 0.021519f
C59 plus.n12 a_n1724_n3888# 0.25476f
C60 plus.n13 a_n1724_n3888# 0.021519f
C61 plus.n14 a_n1724_n3888# 0.25476f
C62 plus.t12 a_n1724_n3888# 0.67413f
C63 plus.n15 a_n1724_n3888# 0.271523f
C64 plus.n16 a_n1724_n3888# 0.664693f
C65 plus.n17 a_n1724_n3888# 0.052244f
C66 plus.t4 a_n1724_n3888# 0.67413f
C67 plus.t11 a_n1724_n3888# 0.663254f
C68 plus.t3 a_n1724_n3888# 0.663254f
C69 plus.t10 a_n1724_n3888# 0.663254f
C70 plus.n18 a_n1724_n3888# 0.272091f
C71 plus.n19 a_n1724_n3888# 0.123088f
C72 plus.t1 a_n1724_n3888# 0.663254f
C73 plus.t8 a_n1724_n3888# 0.663254f
C74 plus.t0 a_n1724_n3888# 0.67413f
C75 plus.n20 a_n1724_n3888# 0.271606f
C76 plus.n21 a_n1724_n3888# 0.25476f
C77 plus.n22 a_n1724_n3888# 0.021519f
C78 plus.n23 a_n1724_n3888# 0.25476f
C79 plus.n24 a_n1724_n3888# 0.021519f
C80 plus.n25 a_n1724_n3888# 0.052244f
C81 plus.n26 a_n1724_n3888# 0.052244f
C82 plus.n27 a_n1724_n3888# 0.052244f
C83 plus.n28 a_n1724_n3888# 0.021519f
C84 plus.n29 a_n1724_n3888# 0.25476f
C85 plus.n30 a_n1724_n3888# 0.021519f
C86 plus.n31 a_n1724_n3888# 0.25476f
C87 plus.n32 a_n1724_n3888# 0.271523f
C88 plus.n33 a_n1724_n3888# 1.63511f
C89 source.t9 a_n1724_n3888# 4.20957f
C90 source.n0 a_n1724_n3888# 1.94979f
C91 source.t4 a_n1724_n3888# 0.375632f
C92 source.t1 a_n1724_n3888# 0.375632f
C93 source.n1 a_n1724_n3888# 3.29962f
C94 source.n2 a_n1724_n3888# 0.423061f
C95 source.t10 a_n1724_n3888# 0.375632f
C96 source.t0 a_n1724_n3888# 0.375632f
C97 source.n3 a_n1724_n3888# 3.29962f
C98 source.n4 a_n1724_n3888# 0.423061f
C99 source.t12 a_n1724_n3888# 0.375632f
C100 source.t13 a_n1724_n3888# 0.375632f
C101 source.n5 a_n1724_n3888# 3.29962f
C102 source.n6 a_n1724_n3888# 0.443308f
C103 source.t19 a_n1724_n3888# 4.20957f
C104 source.n7 a_n1724_n3888# 0.557804f
C105 source.t26 a_n1724_n3888# 0.375632f
C106 source.t15 a_n1724_n3888# 0.375632f
C107 source.n8 a_n1724_n3888# 3.29962f
C108 source.n9 a_n1724_n3888# 0.423061f
C109 source.t18 a_n1724_n3888# 0.375632f
C110 source.t22 a_n1724_n3888# 0.375632f
C111 source.n10 a_n1724_n3888# 3.29962f
C112 source.n11 a_n1724_n3888# 0.423061f
C113 source.t23 a_n1724_n3888# 0.375632f
C114 source.t27 a_n1724_n3888# 0.375632f
C115 source.n12 a_n1724_n3888# 3.29962f
C116 source.n13 a_n1724_n3888# 2.41762f
C117 source.t11 a_n1724_n3888# 0.375632f
C118 source.t6 a_n1724_n3888# 0.375632f
C119 source.n14 a_n1724_n3888# 3.29961f
C120 source.n15 a_n1724_n3888# 2.41762f
C121 source.t2 a_n1724_n3888# 0.375632f
C122 source.t5 a_n1724_n3888# 0.375632f
C123 source.n16 a_n1724_n3888# 3.29961f
C124 source.n17 a_n1724_n3888# 0.423066f
C125 source.t8 a_n1724_n3888# 0.375632f
C126 source.t7 a_n1724_n3888# 0.375632f
C127 source.n18 a_n1724_n3888# 3.29961f
C128 source.n19 a_n1724_n3888# 0.423066f
C129 source.t3 a_n1724_n3888# 4.20957f
C130 source.n20 a_n1724_n3888# 0.557809f
C131 source.t24 a_n1724_n3888# 0.375632f
C132 source.t16 a_n1724_n3888# 0.375632f
C133 source.n21 a_n1724_n3888# 3.29961f
C134 source.n22 a_n1724_n3888# 0.443312f
C135 source.t25 a_n1724_n3888# 0.375632f
C136 source.t17 a_n1724_n3888# 0.375632f
C137 source.n23 a_n1724_n3888# 3.29961f
C138 source.n24 a_n1724_n3888# 0.423066f
C139 source.t20 a_n1724_n3888# 0.375632f
C140 source.t14 a_n1724_n3888# 0.375632f
C141 source.n25 a_n1724_n3888# 3.29961f
C142 source.n26 a_n1724_n3888# 0.423066f
C143 source.t21 a_n1724_n3888# 4.20957f
C144 source.n27 a_n1724_n3888# 0.708969f
C145 source.n28 a_n1724_n3888# 2.3171f
C146 drain_right.t4 a_n1724_n3888# 4.225f
C147 drain_right.t5 a_n1724_n3888# 0.365891f
C148 drain_right.t6 a_n1724_n3888# 0.365891f
C149 drain_right.n0 a_n1724_n3888# 3.30723f
C150 drain_right.n1 a_n1724_n3888# 0.743279f
C151 drain_right.t2 a_n1724_n3888# 0.365891f
C152 drain_right.t3 a_n1724_n3888# 0.365891f
C153 drain_right.n2 a_n1724_n3888# 3.31053f
C154 drain_right.t7 a_n1724_n3888# 0.365891f
C155 drain_right.t0 a_n1724_n3888# 0.365891f
C156 drain_right.n3 a_n1724_n3888# 3.30723f
C157 drain_right.n4 a_n1724_n3888# 0.69374f
C158 drain_right.n5 a_n1724_n3888# 1.62387f
C159 drain_right.t12 a_n1724_n3888# 0.365891f
C160 drain_right.t11 a_n1724_n3888# 0.365891f
C161 drain_right.n6 a_n1724_n3888# 3.31052f
C162 drain_right.t1 a_n1724_n3888# 0.365891f
C163 drain_right.t8 a_n1724_n3888# 0.365891f
C164 drain_right.n7 a_n1724_n3888# 3.30723f
C165 drain_right.n8 a_n1724_n3888# 0.730868f
C166 drain_right.t10 a_n1724_n3888# 0.365891f
C167 drain_right.t9 a_n1724_n3888# 0.365891f
C168 drain_right.n9 a_n1724_n3888# 3.30723f
C169 drain_right.n10 a_n1724_n3888# 0.360862f
C170 drain_right.t13 a_n1724_n3888# 4.22152f
C171 drain_right.n11 a_n1724_n3888# 0.660389f
C172 minus.n0 a_n1724_n3888# 0.051667f
C173 minus.t4 a_n1724_n3888# 0.666679f
C174 minus.t0 a_n1724_n3888# 0.655923f
C175 minus.t9 a_n1724_n3888# 0.655923f
C176 minus.t5 a_n1724_n3888# 0.655923f
C177 minus.n1 a_n1724_n3888# 0.269084f
C178 minus.n2 a_n1724_n3888# 0.121728f
C179 minus.t1 a_n1724_n3888# 0.655923f
C180 minus.t12 a_n1724_n3888# 0.655923f
C181 minus.t8 a_n1724_n3888# 0.666679f
C182 minus.n3 a_n1724_n3888# 0.268604f
C183 minus.n4 a_n1724_n3888# 0.251944f
C184 minus.n5 a_n1724_n3888# 0.021281f
C185 minus.n6 a_n1724_n3888# 0.251944f
C186 minus.n7 a_n1724_n3888# 0.021281f
C187 minus.n8 a_n1724_n3888# 0.051667f
C188 minus.n9 a_n1724_n3888# 0.051667f
C189 minus.n10 a_n1724_n3888# 0.051667f
C190 minus.n11 a_n1724_n3888# 0.021281f
C191 minus.n12 a_n1724_n3888# 0.251944f
C192 minus.n13 a_n1724_n3888# 0.021281f
C193 minus.n14 a_n1724_n3888# 0.251944f
C194 minus.n15 a_n1724_n3888# 0.268522f
C195 minus.n16 a_n1724_n3888# 1.96716f
C196 minus.n17 a_n1724_n3888# 0.051667f
C197 minus.t13 a_n1724_n3888# 0.655923f
C198 minus.t7 a_n1724_n3888# 0.655923f
C199 minus.t10 a_n1724_n3888# 0.655923f
C200 minus.n18 a_n1724_n3888# 0.269084f
C201 minus.n19 a_n1724_n3888# 0.121728f
C202 minus.t2 a_n1724_n3888# 0.655923f
C203 minus.t11 a_n1724_n3888# 0.655923f
C204 minus.t3 a_n1724_n3888# 0.666679f
C205 minus.n20 a_n1724_n3888# 0.268604f
C206 minus.n21 a_n1724_n3888# 0.251944f
C207 minus.n22 a_n1724_n3888# 0.021281f
C208 minus.n23 a_n1724_n3888# 0.251944f
C209 minus.n24 a_n1724_n3888# 0.021281f
C210 minus.n25 a_n1724_n3888# 0.051667f
C211 minus.n26 a_n1724_n3888# 0.051667f
C212 minus.n27 a_n1724_n3888# 0.051667f
C213 minus.n28 a_n1724_n3888# 0.021281f
C214 minus.n29 a_n1724_n3888# 0.251944f
C215 minus.n30 a_n1724_n3888# 0.021281f
C216 minus.n31 a_n1724_n3888# 0.251944f
C217 minus.t6 a_n1724_n3888# 0.666679f
C218 minus.n32 a_n1724_n3888# 0.268522f
C219 minus.n33 a_n1724_n3888# 0.34222f
C220 minus.n34 a_n1724_n3888# 2.37573f
.ends

