* NGSPICE file created from diffpair187.ext - technology: sky130A

.subckt diffpair187 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t25 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 drain_left.t14 plus.t1 source.t26 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 drain_right.t15 minus.t0 source.t8 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X3 source.t2 minus.t1 drain_right.t14 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X4 source.t1 minus.t2 drain_right.t13 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X5 drain_right.t12 minus.t3 source.t3 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X6 drain_left.t13 plus.t2 source.t27 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X7 source.t6 minus.t4 drain_right.t11 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X8 a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X9 source.t28 plus.t3 drain_left.t12 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X10 source.t31 plus.t4 drain_left.t11 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X11 drain_left.t10 plus.t5 source.t23 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X12 drain_left.t9 plus.t6 source.t17 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X13 source.t9 minus.t5 drain_right.t10 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X14 source.t11 minus.t6 drain_right.t9 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X15 a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X16 drain_left.t8 plus.t7 source.t19 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X17 drain_left.t7 plus.t8 source.t29 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 source.t30 plus.t9 drain_left.t6 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X19 source.t20 plus.t10 drain_left.t5 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X20 source.t21 plus.t11 drain_left.t4 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X21 source.t16 plus.t12 drain_left.t3 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X22 a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X23 source.t22 plus.t13 drain_left.t2 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X24 source.t24 plus.t14 drain_left.t1 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X25 drain_right.t8 minus.t7 source.t0 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X26 drain_right.t7 minus.t8 source.t13 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X27 drain_right.t6 minus.t9 source.t4 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X28 drain_right.t5 minus.t10 source.t12 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X29 source.t15 minus.t11 drain_right.t4 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X30 drain_right.t3 minus.t12 source.t5 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X31 drain_right.t2 minus.t13 source.t14 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X32 a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X33 source.t7 minus.t14 drain_right.t1 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X34 drain_left.t0 plus.t15 source.t18 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X35 source.t10 minus.t15 drain_right.t0 a_n1760_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n4 plus.t3 455.418
R1 plus.n19 plus.t2 455.418
R2 plus.n25 plus.t6 455.418
R3 plus.n40 plus.t13 455.418
R4 plus.n5 plus.t1 414.521
R5 plus.n3 plus.t12 414.521
R6 plus.n10 plus.t0 414.521
R7 plus.n1 plus.t11 414.521
R8 plus.n16 plus.t15 414.521
R9 plus.n18 plus.t10 414.521
R10 plus.n26 plus.t4 414.521
R11 plus.n24 plus.t8 414.521
R12 plus.n31 plus.t14 414.521
R13 plus.n22 plus.t5 414.521
R14 plus.n37 plus.t9 414.521
R15 plus.n39 plus.t7 414.521
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus.n6 plus.n5 29.2126
R47 plus.n18 plus.n17 29.2126
R48 plus.n39 plus.n38 29.2126
R49 plus.n27 plus.n26 29.2126
R50 plus plus.n41 26.2263
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 8.70126
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n0 source.t27 69.6943
R73 source.n7 source.t28 69.6943
R74 source.n8 source.t13 69.6943
R75 source.n15 source.t9 69.6943
R76 source.n31 source.t8 69.6942
R77 source.n24 source.t10 69.6942
R78 source.n23 source.t17 69.6942
R79 source.n16 source.t22 69.6942
R80 source.n2 source.n1 63.0943
R81 source.n4 source.n3 63.0943
R82 source.n6 source.n5 63.0943
R83 source.n10 source.n9 63.0943
R84 source.n12 source.n11 63.0943
R85 source.n14 source.n13 63.0943
R86 source.n30 source.n29 63.0942
R87 source.n28 source.n27 63.0942
R88 source.n26 source.n25 63.0942
R89 source.n22 source.n21 63.0942
R90 source.n20 source.n19 63.0942
R91 source.n18 source.n17 63.0942
R92 source.n16 source.n15 14.9695
R93 source.n32 source.n0 9.45661
R94 source.n29 source.t3 6.6005
R95 source.n29 source.t2 6.6005
R96 source.n27 source.t12 6.6005
R97 source.n27 source.t7 6.6005
R98 source.n25 source.t4 6.6005
R99 source.n25 source.t15 6.6005
R100 source.n21 source.t29 6.6005
R101 source.n21 source.t31 6.6005
R102 source.n19 source.t23 6.6005
R103 source.n19 source.t24 6.6005
R104 source.n17 source.t19 6.6005
R105 source.n17 source.t30 6.6005
R106 source.n1 source.t18 6.6005
R107 source.n1 source.t20 6.6005
R108 source.n3 source.t25 6.6005
R109 source.n3 source.t21 6.6005
R110 source.n5 source.t26 6.6005
R111 source.n5 source.t16 6.6005
R112 source.n9 source.t0 6.6005
R113 source.n9 source.t6 6.6005
R114 source.n11 source.t5 6.6005
R115 source.n11 source.t1 6.6005
R116 source.n13 source.t14 6.6005
R117 source.n13 source.t11 6.6005
R118 source.n32 source.n31 5.51343
R119 source.n15 source.n14 0.5005
R120 source.n14 source.n12 0.5005
R121 source.n12 source.n10 0.5005
R122 source.n10 source.n8 0.5005
R123 source.n7 source.n6 0.5005
R124 source.n6 source.n4 0.5005
R125 source.n4 source.n2 0.5005
R126 source.n2 source.n0 0.5005
R127 source.n18 source.n16 0.5005
R128 source.n20 source.n18 0.5005
R129 source.n22 source.n20 0.5005
R130 source.n23 source.n22 0.5005
R131 source.n26 source.n24 0.5005
R132 source.n28 source.n26 0.5005
R133 source.n30 source.n28 0.5005
R134 source.n31 source.n30 0.5005
R135 source.n8 source.n7 0.470328
R136 source.n24 source.n23 0.470328
R137 source source.n32 0.188
R138 drain_left.n9 drain_left.n7 80.2731
R139 drain_left.n5 drain_left.n3 80.273
R140 drain_left.n2 drain_left.n0 80.273
R141 drain_left.n13 drain_left.n12 79.7731
R142 drain_left.n11 drain_left.n10 79.7731
R143 drain_left.n9 drain_left.n8 79.7731
R144 drain_left.n5 drain_left.n4 79.773
R145 drain_left.n2 drain_left.n1 79.773
R146 drain_left drain_left.n6 23.7989
R147 drain_left.n3 drain_left.t11 6.6005
R148 drain_left.n3 drain_left.t9 6.6005
R149 drain_left.n4 drain_left.t1 6.6005
R150 drain_left.n4 drain_left.t7 6.6005
R151 drain_left.n1 drain_left.t6 6.6005
R152 drain_left.n1 drain_left.t10 6.6005
R153 drain_left.n0 drain_left.t2 6.6005
R154 drain_left.n0 drain_left.t8 6.6005
R155 drain_left.n12 drain_left.t5 6.6005
R156 drain_left.n12 drain_left.t13 6.6005
R157 drain_left.n10 drain_left.t4 6.6005
R158 drain_left.n10 drain_left.t0 6.6005
R159 drain_left.n8 drain_left.t3 6.6005
R160 drain_left.n8 drain_left.t15 6.6005
R161 drain_left.n7 drain_left.t12 6.6005
R162 drain_left.n7 drain_left.t14 6.6005
R163 drain_left drain_left.n13 6.15322
R164 drain_left.n11 drain_left.n9 0.5005
R165 drain_left.n13 drain_left.n11 0.5005
R166 drain_left.n6 drain_left.n5 0.195154
R167 drain_left.n6 drain_left.n2 0.195154
R168 minus.n19 minus.t5 455.418
R169 minus.n4 minus.t8 455.418
R170 minus.n40 minus.t0 455.418
R171 minus.n25 minus.t15 455.418
R172 minus.n18 minus.t13 414.521
R173 minus.n16 minus.t6 414.521
R174 minus.n1 minus.t12 414.521
R175 minus.n10 minus.t2 414.521
R176 minus.n3 minus.t7 414.521
R177 minus.n5 minus.t4 414.521
R178 minus.n39 minus.t1 414.521
R179 minus.n37 minus.t3 414.521
R180 minus.n22 minus.t14 414.521
R181 minus.n31 minus.t10 414.521
R182 minus.n24 minus.t11 414.521
R183 minus.n26 minus.t9 414.521
R184 minus.n7 minus.n4 161.489
R185 minus.n28 minus.n25 161.489
R186 minus.n20 minus.n19 161.3
R187 minus.n17 minus.n0 161.3
R188 minus.n15 minus.n14 161.3
R189 minus.n13 minus.n12 161.3
R190 minus.n11 minus.n2 161.3
R191 minus.n9 minus.n8 161.3
R192 minus.n7 minus.n6 161.3
R193 minus.n41 minus.n40 161.3
R194 minus.n38 minus.n21 161.3
R195 minus.n36 minus.n35 161.3
R196 minus.n34 minus.n33 161.3
R197 minus.n32 minus.n23 161.3
R198 minus.n30 minus.n29 161.3
R199 minus.n28 minus.n27 161.3
R200 minus.n12 minus.n11 73.0308
R201 minus.n33 minus.n32 73.0308
R202 minus.n15 minus.n1 67.1884
R203 minus.n10 minus.n9 67.1884
R204 minus.n31 minus.n30 67.1884
R205 minus.n36 minus.n22 67.1884
R206 minus.n17 minus.n16 55.5035
R207 minus.n6 minus.n3 55.5035
R208 minus.n27 minus.n24 55.5035
R209 minus.n38 minus.n37 55.5035
R210 minus.n19 minus.n18 43.8187
R211 minus.n5 minus.n4 43.8187
R212 minus.n26 minus.n25 43.8187
R213 minus.n40 minus.n39 43.8187
R214 minus.n18 minus.n17 29.2126
R215 minus.n6 minus.n5 29.2126
R216 minus.n27 minus.n26 29.2126
R217 minus.n39 minus.n38 29.2126
R218 minus.n42 minus.n20 28.9361
R219 minus.n16 minus.n15 17.5278
R220 minus.n9 minus.n3 17.5278
R221 minus.n30 minus.n24 17.5278
R222 minus.n37 minus.n36 17.5278
R223 minus.n42 minus.n41 6.46641
R224 minus.n12 minus.n1 5.84292
R225 minus.n11 minus.n10 5.84292
R226 minus.n32 minus.n31 5.84292
R227 minus.n33 minus.n22 5.84292
R228 minus.n20 minus.n0 0.189894
R229 minus.n14 minus.n0 0.189894
R230 minus.n14 minus.n13 0.189894
R231 minus.n13 minus.n2 0.189894
R232 minus.n8 minus.n2 0.189894
R233 minus.n8 minus.n7 0.189894
R234 minus.n29 minus.n28 0.189894
R235 minus.n29 minus.n23 0.189894
R236 minus.n34 minus.n23 0.189894
R237 minus.n35 minus.n34 0.189894
R238 minus.n35 minus.n21 0.189894
R239 minus.n41 minus.n21 0.189894
R240 minus minus.n42 0.188
R241 drain_right.n9 drain_right.n7 80.2731
R242 drain_right.n5 drain_right.n3 80.273
R243 drain_right.n2 drain_right.n0 80.273
R244 drain_right.n9 drain_right.n8 79.7731
R245 drain_right.n11 drain_right.n10 79.7731
R246 drain_right.n13 drain_right.n12 79.7731
R247 drain_right.n5 drain_right.n4 79.773
R248 drain_right.n2 drain_right.n1 79.773
R249 drain_right drain_right.n6 23.2457
R250 drain_right.n3 drain_right.t14 6.6005
R251 drain_right.n3 drain_right.t15 6.6005
R252 drain_right.n4 drain_right.t1 6.6005
R253 drain_right.n4 drain_right.t12 6.6005
R254 drain_right.n1 drain_right.t4 6.6005
R255 drain_right.n1 drain_right.t5 6.6005
R256 drain_right.n0 drain_right.t0 6.6005
R257 drain_right.n0 drain_right.t6 6.6005
R258 drain_right.n7 drain_right.t11 6.6005
R259 drain_right.n7 drain_right.t7 6.6005
R260 drain_right.n8 drain_right.t13 6.6005
R261 drain_right.n8 drain_right.t8 6.6005
R262 drain_right.n10 drain_right.t9 6.6005
R263 drain_right.n10 drain_right.t3 6.6005
R264 drain_right.n12 drain_right.t10 6.6005
R265 drain_right.n12 drain_right.t2 6.6005
R266 drain_right drain_right.n13 6.15322
R267 drain_right.n13 drain_right.n11 0.5005
R268 drain_right.n11 drain_right.n9 0.5005
R269 drain_right.n6 drain_right.n5 0.195154
R270 drain_right.n6 drain_right.n2 0.195154
C0 source plus 1.79065f
C1 drain_right drain_left 0.897273f
C2 drain_left minus 0.176274f
C3 drain_right plus 0.330041f
C4 minus plus 3.6902f
C5 drain_left plus 1.84693f
C6 drain_right source 10.38f
C7 source minus 1.77665f
C8 source drain_left 10.38f
C9 drain_right minus 1.67661f
C10 drain_right a_n1760_n1488# 4.18283f
C11 drain_left a_n1760_n1488# 4.43058f
C12 source a_n1760_n1488# 3.645067f
C13 minus a_n1760_n1488# 6.128285f
C14 plus a_n1760_n1488# 6.747104f
C15 drain_right.t0 a_n1760_n1488# 0.069052f
C16 drain_right.t6 a_n1760_n1488# 0.069052f
C17 drain_right.n0 a_n1760_n1488# 0.500107f
C18 drain_right.t4 a_n1760_n1488# 0.069052f
C19 drain_right.t5 a_n1760_n1488# 0.069052f
C20 drain_right.n1 a_n1760_n1488# 0.497997f
C21 drain_right.n2 a_n1760_n1488# 0.638464f
C22 drain_right.t14 a_n1760_n1488# 0.069052f
C23 drain_right.t15 a_n1760_n1488# 0.069052f
C24 drain_right.n3 a_n1760_n1488# 0.500107f
C25 drain_right.t1 a_n1760_n1488# 0.069052f
C26 drain_right.t12 a_n1760_n1488# 0.069052f
C27 drain_right.n4 a_n1760_n1488# 0.497997f
C28 drain_right.n5 a_n1760_n1488# 0.638464f
C29 drain_right.n6 a_n1760_n1488# 0.794946f
C30 drain_right.t11 a_n1760_n1488# 0.069052f
C31 drain_right.t7 a_n1760_n1488# 0.069052f
C32 drain_right.n7 a_n1760_n1488# 0.500109f
C33 drain_right.t13 a_n1760_n1488# 0.069052f
C34 drain_right.t8 a_n1760_n1488# 0.069052f
C35 drain_right.n8 a_n1760_n1488# 0.497999f
C36 drain_right.n9 a_n1760_n1488# 0.663648f
C37 drain_right.t9 a_n1760_n1488# 0.069052f
C38 drain_right.t3 a_n1760_n1488# 0.069052f
C39 drain_right.n10 a_n1760_n1488# 0.497999f
C40 drain_right.n11 a_n1760_n1488# 0.327013f
C41 drain_right.t10 a_n1760_n1488# 0.069052f
C42 drain_right.t2 a_n1760_n1488# 0.069052f
C43 drain_right.n12 a_n1760_n1488# 0.497999f
C44 drain_right.n13 a_n1760_n1488# 0.56744f
C45 minus.n0 a_n1760_n1488# 0.026824f
C46 minus.t5 a_n1760_n1488# 0.061466f
C47 minus.t13 a_n1760_n1488# 0.05826f
C48 minus.t6 a_n1760_n1488# 0.05826f
C49 minus.t12 a_n1760_n1488# 0.05826f
C50 minus.n1 a_n1760_n1488# 0.035207f
C51 minus.n2 a_n1760_n1488# 0.026824f
C52 minus.t2 a_n1760_n1488# 0.05826f
C53 minus.t7 a_n1760_n1488# 0.05826f
C54 minus.n3 a_n1760_n1488# 0.035207f
C55 minus.t8 a_n1760_n1488# 0.061466f
C56 minus.n4 a_n1760_n1488# 0.042756f
C57 minus.t4 a_n1760_n1488# 0.05826f
C58 minus.n5 a_n1760_n1488# 0.035207f
C59 minus.n6 a_n1760_n1488# 0.010222f
C60 minus.n7 a_n1760_n1488# 0.058738f
C61 minus.n8 a_n1760_n1488# 0.026824f
C62 minus.n9 a_n1760_n1488# 0.010222f
C63 minus.n10 a_n1760_n1488# 0.035207f
C64 minus.n11 a_n1760_n1488# 0.00956f
C65 minus.n12 a_n1760_n1488# 0.00956f
C66 minus.n13 a_n1760_n1488# 0.026824f
C67 minus.n14 a_n1760_n1488# 0.026824f
C68 minus.n15 a_n1760_n1488# 0.010222f
C69 minus.n16 a_n1760_n1488# 0.035207f
C70 minus.n17 a_n1760_n1488# 0.010222f
C71 minus.n18 a_n1760_n1488# 0.035207f
C72 minus.n19 a_n1760_n1488# 0.042718f
C73 minus.n20 a_n1760_n1488# 0.654844f
C74 minus.n21 a_n1760_n1488# 0.026824f
C75 minus.t1 a_n1760_n1488# 0.05826f
C76 minus.t3 a_n1760_n1488# 0.05826f
C77 minus.t14 a_n1760_n1488# 0.05826f
C78 minus.n22 a_n1760_n1488# 0.035207f
C79 minus.n23 a_n1760_n1488# 0.026824f
C80 minus.t10 a_n1760_n1488# 0.05826f
C81 minus.t11 a_n1760_n1488# 0.05826f
C82 minus.n24 a_n1760_n1488# 0.035207f
C83 minus.t15 a_n1760_n1488# 0.061466f
C84 minus.n25 a_n1760_n1488# 0.042756f
C85 minus.t9 a_n1760_n1488# 0.05826f
C86 minus.n26 a_n1760_n1488# 0.035207f
C87 minus.n27 a_n1760_n1488# 0.010222f
C88 minus.n28 a_n1760_n1488# 0.058738f
C89 minus.n29 a_n1760_n1488# 0.026824f
C90 minus.n30 a_n1760_n1488# 0.010222f
C91 minus.n31 a_n1760_n1488# 0.035207f
C92 minus.n32 a_n1760_n1488# 0.00956f
C93 minus.n33 a_n1760_n1488# 0.00956f
C94 minus.n34 a_n1760_n1488# 0.026824f
C95 minus.n35 a_n1760_n1488# 0.026824f
C96 minus.n36 a_n1760_n1488# 0.010222f
C97 minus.n37 a_n1760_n1488# 0.035207f
C98 minus.n38 a_n1760_n1488# 0.010222f
C99 minus.n39 a_n1760_n1488# 0.035207f
C100 minus.t0 a_n1760_n1488# 0.061466f
C101 minus.n40 a_n1760_n1488# 0.042718f
C102 minus.n41 a_n1760_n1488# 0.173245f
C103 minus.n42 a_n1760_n1488# 0.810144f
C104 drain_left.t2 a_n1760_n1488# 0.068304f
C105 drain_left.t8 a_n1760_n1488# 0.068304f
C106 drain_left.n0 a_n1760_n1488# 0.494687f
C107 drain_left.t6 a_n1760_n1488# 0.068304f
C108 drain_left.t10 a_n1760_n1488# 0.068304f
C109 drain_left.n1 a_n1760_n1488# 0.4926f
C110 drain_left.n2 a_n1760_n1488# 0.631545f
C111 drain_left.t11 a_n1760_n1488# 0.068304f
C112 drain_left.t9 a_n1760_n1488# 0.068304f
C113 drain_left.n3 a_n1760_n1488# 0.494687f
C114 drain_left.t1 a_n1760_n1488# 0.068304f
C115 drain_left.t7 a_n1760_n1488# 0.068304f
C116 drain_left.n4 a_n1760_n1488# 0.4926f
C117 drain_left.n5 a_n1760_n1488# 0.631545f
C118 drain_left.n6 a_n1760_n1488# 0.843472f
C119 drain_left.t12 a_n1760_n1488# 0.068304f
C120 drain_left.t14 a_n1760_n1488# 0.068304f
C121 drain_left.n7 a_n1760_n1488# 0.494689f
C122 drain_left.t3 a_n1760_n1488# 0.068304f
C123 drain_left.t15 a_n1760_n1488# 0.068304f
C124 drain_left.n8 a_n1760_n1488# 0.492602f
C125 drain_left.n9 a_n1760_n1488# 0.656456f
C126 drain_left.t4 a_n1760_n1488# 0.068304f
C127 drain_left.t0 a_n1760_n1488# 0.068304f
C128 drain_left.n10 a_n1760_n1488# 0.492602f
C129 drain_left.n11 a_n1760_n1488# 0.323469f
C130 drain_left.t5 a_n1760_n1488# 0.068304f
C131 drain_left.t13 a_n1760_n1488# 0.068304f
C132 drain_left.n12 a_n1760_n1488# 0.492602f
C133 drain_left.n13 a_n1760_n1488# 0.561291f
C134 source.t27 a_n1760_n1488# 0.551123f
C135 source.n0 a_n1760_n1488# 0.745066f
C136 source.t18 a_n1760_n1488# 0.06637f
C137 source.t20 a_n1760_n1488# 0.06637f
C138 source.n1 a_n1760_n1488# 0.420823f
C139 source.n2 a_n1760_n1488# 0.33409f
C140 source.t25 a_n1760_n1488# 0.06637f
C141 source.t21 a_n1760_n1488# 0.06637f
C142 source.n3 a_n1760_n1488# 0.420823f
C143 source.n4 a_n1760_n1488# 0.33409f
C144 source.t26 a_n1760_n1488# 0.06637f
C145 source.t16 a_n1760_n1488# 0.06637f
C146 source.n5 a_n1760_n1488# 0.420823f
C147 source.n6 a_n1760_n1488# 0.33409f
C148 source.t28 a_n1760_n1488# 0.551123f
C149 source.n7 a_n1760_n1488# 0.382077f
C150 source.t13 a_n1760_n1488# 0.551123f
C151 source.n8 a_n1760_n1488# 0.382077f
C152 source.t0 a_n1760_n1488# 0.06637f
C153 source.t6 a_n1760_n1488# 0.06637f
C154 source.n9 a_n1760_n1488# 0.420823f
C155 source.n10 a_n1760_n1488# 0.33409f
C156 source.t5 a_n1760_n1488# 0.06637f
C157 source.t1 a_n1760_n1488# 0.06637f
C158 source.n11 a_n1760_n1488# 0.420823f
C159 source.n12 a_n1760_n1488# 0.33409f
C160 source.t14 a_n1760_n1488# 0.06637f
C161 source.t11 a_n1760_n1488# 0.06637f
C162 source.n13 a_n1760_n1488# 0.420823f
C163 source.n14 a_n1760_n1488# 0.33409f
C164 source.t9 a_n1760_n1488# 0.551123f
C165 source.n15 a_n1760_n1488# 1.03596f
C166 source.t22 a_n1760_n1488# 0.55112f
C167 source.n16 a_n1760_n1488# 1.03596f
C168 source.t19 a_n1760_n1488# 0.06637f
C169 source.t30 a_n1760_n1488# 0.06637f
C170 source.n17 a_n1760_n1488# 0.42082f
C171 source.n18 a_n1760_n1488# 0.334093f
C172 source.t23 a_n1760_n1488# 0.06637f
C173 source.t24 a_n1760_n1488# 0.06637f
C174 source.n19 a_n1760_n1488# 0.42082f
C175 source.n20 a_n1760_n1488# 0.334093f
C176 source.t29 a_n1760_n1488# 0.06637f
C177 source.t31 a_n1760_n1488# 0.06637f
C178 source.n21 a_n1760_n1488# 0.42082f
C179 source.n22 a_n1760_n1488# 0.334093f
C180 source.t17 a_n1760_n1488# 0.55112f
C181 source.n23 a_n1760_n1488# 0.382079f
C182 source.t10 a_n1760_n1488# 0.55112f
C183 source.n24 a_n1760_n1488# 0.382079f
C184 source.t4 a_n1760_n1488# 0.06637f
C185 source.t15 a_n1760_n1488# 0.06637f
C186 source.n25 a_n1760_n1488# 0.42082f
C187 source.n26 a_n1760_n1488# 0.334093f
C188 source.t12 a_n1760_n1488# 0.06637f
C189 source.t7 a_n1760_n1488# 0.06637f
C190 source.n27 a_n1760_n1488# 0.42082f
C191 source.n28 a_n1760_n1488# 0.334093f
C192 source.t3 a_n1760_n1488# 0.06637f
C193 source.t2 a_n1760_n1488# 0.06637f
C194 source.n29 a_n1760_n1488# 0.42082f
C195 source.n30 a_n1760_n1488# 0.334093f
C196 source.t8 a_n1760_n1488# 0.55112f
C197 source.n31 a_n1760_n1488# 0.537004f
C198 source.n32 a_n1760_n1488# 0.809766f
C199 plus.n0 a_n1760_n1488# 0.027223f
C200 plus.t10 a_n1760_n1488# 0.059127f
C201 plus.t15 a_n1760_n1488# 0.059127f
C202 plus.t11 a_n1760_n1488# 0.059127f
C203 plus.n1 a_n1760_n1488# 0.035731f
C204 plus.n2 a_n1760_n1488# 0.027223f
C205 plus.t0 a_n1760_n1488# 0.059127f
C206 plus.t12 a_n1760_n1488# 0.059127f
C207 plus.n3 a_n1760_n1488# 0.035731f
C208 plus.t3 a_n1760_n1488# 0.062381f
C209 plus.n4 a_n1760_n1488# 0.043392f
C210 plus.t1 a_n1760_n1488# 0.059127f
C211 plus.n5 a_n1760_n1488# 0.035731f
C212 plus.n6 a_n1760_n1488# 0.010374f
C213 plus.n7 a_n1760_n1488# 0.059612f
C214 plus.n8 a_n1760_n1488# 0.027223f
C215 plus.n9 a_n1760_n1488# 0.010374f
C216 plus.n10 a_n1760_n1488# 0.035731f
C217 plus.n11 a_n1760_n1488# 0.009702f
C218 plus.n12 a_n1760_n1488# 0.009702f
C219 plus.n13 a_n1760_n1488# 0.027223f
C220 plus.n14 a_n1760_n1488# 0.027223f
C221 plus.n15 a_n1760_n1488# 0.010374f
C222 plus.n16 a_n1760_n1488# 0.035731f
C223 plus.n17 a_n1760_n1488# 0.010374f
C224 plus.n18 a_n1760_n1488# 0.035731f
C225 plus.t2 a_n1760_n1488# 0.062381f
C226 plus.n19 a_n1760_n1488# 0.043354f
C227 plus.n20 a_n1760_n1488# 0.201086f
C228 plus.n21 a_n1760_n1488# 0.027223f
C229 plus.t13 a_n1760_n1488# 0.062381f
C230 plus.t7 a_n1760_n1488# 0.059127f
C231 plus.t9 a_n1760_n1488# 0.059127f
C232 plus.t5 a_n1760_n1488# 0.059127f
C233 plus.n22 a_n1760_n1488# 0.035731f
C234 plus.n23 a_n1760_n1488# 0.027223f
C235 plus.t14 a_n1760_n1488# 0.059127f
C236 plus.t8 a_n1760_n1488# 0.059127f
C237 plus.n24 a_n1760_n1488# 0.035731f
C238 plus.t6 a_n1760_n1488# 0.062381f
C239 plus.n25 a_n1760_n1488# 0.043392f
C240 plus.t4 a_n1760_n1488# 0.059127f
C241 plus.n26 a_n1760_n1488# 0.035731f
C242 plus.n27 a_n1760_n1488# 0.010374f
C243 plus.n28 a_n1760_n1488# 0.059612f
C244 plus.n29 a_n1760_n1488# 0.027223f
C245 plus.n30 a_n1760_n1488# 0.010374f
C246 plus.n31 a_n1760_n1488# 0.035731f
C247 plus.n32 a_n1760_n1488# 0.009702f
C248 plus.n33 a_n1760_n1488# 0.009702f
C249 plus.n34 a_n1760_n1488# 0.027223f
C250 plus.n35 a_n1760_n1488# 0.027223f
C251 plus.n36 a_n1760_n1488# 0.010374f
C252 plus.n37 a_n1760_n1488# 0.035731f
C253 plus.n38 a_n1760_n1488# 0.010374f
C254 plus.n39 a_n1760_n1488# 0.035731f
C255 plus.n40 a_n1760_n1488# 0.043354f
C256 plus.n41 a_n1760_n1488# 0.625383f
.ends

