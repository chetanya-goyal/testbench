* NGSPICE file created from diffpair394.ext - technology: sky130A

.subckt diffpair394 minus drain_right drain_left source plus
X0 source.t18 minus.t0 drain_right.t7 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X1 source.t19 plus.t0 drain_left.t9 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X2 a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X3 a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X4 source.t0 plus.t1 drain_left.t8 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X5 source.t17 minus.t1 drain_right.t6 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X7 drain_right.t8 minus.t2 source.t16 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 drain_left.t7 plus.t2 source.t3 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X9 drain_left.t6 plus.t3 source.t7 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 source.t15 minus.t3 drain_right.t0 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 drain_right.t2 minus.t4 source.t14 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X12 drain_right.t4 minus.t5 source.t13 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X13 source.t12 minus.t6 drain_right.t5 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X14 drain_left.t5 plus.t4 source.t4 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X15 drain_right.t3 minus.t7 source.t11 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X16 a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X17 drain_right.t9 minus.t8 source.t10 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X18 source.t6 plus.t5 drain_left.t4 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 drain_right.t1 minus.t9 source.t9 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X20 drain_left.t3 plus.t6 source.t1 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X21 drain_left.t2 plus.t7 source.t2 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X22 source.t5 plus.t8 drain_left.t1 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X23 drain_left.t0 plus.t9 source.t8 a_n2072_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n3 minus.t5 343.425
R1 minus.n13 minus.t9 343.425
R2 minus.n2 minus.t3 320.229
R3 minus.n1 minus.t2 320.229
R4 minus.n6 minus.t6 320.229
R5 minus.n8 minus.t7 320.229
R6 minus.n12 minus.t1 320.229
R7 minus.n11 minus.t4 320.229
R8 minus.n16 minus.t0 320.229
R9 minus.n18 minus.t8 320.229
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n19 minus.n18 161.3
R13 minus.n17 minus.n10 161.3
R14 minus.n6 minus.n5 80.6037
R15 minus.n4 minus.n1 80.6037
R16 minus.n16 minus.n15 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n20 minus.n9 34.8736
R23 minus.n7 minus.n6 32.1338
R24 minus.n17 minus.n16 32.1338
R25 minus.n4 minus.n3 31.8629
R26 minus.n14 minus.n13 31.8629
R27 minus.n3 minus.n2 16.2333
R28 minus.n13 minus.n12 16.2333
R29 minus.n8 minus.n7 16.0672
R30 minus.n18 minus.n17 16.0672
R31 minus.n20 minus.n19 6.67664
R32 minus.n5 minus.n4 0.380177
R33 minus.n15 minus.n14 0.380177
R34 minus.n5 minus.n0 0.285035
R35 minus.n15 minus.n10 0.285035
R36 minus.n9 minus.n0 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 drain_right.n1 drain_right.t1 68.7115
R40 drain_right.n7 drain_right.t3 67.7376
R41 drain_right.n6 drain_right.n4 66.5116
R42 drain_right.n3 drain_right.n2 66.2126
R43 drain_right.n6 drain_right.n5 65.5376
R44 drain_right.n1 drain_right.n0 65.5373
R45 drain_right drain_right.n3 28.6812
R46 drain_right drain_right.n7 6.14028
R47 drain_right.n2 drain_right.t7 2.2005
R48 drain_right.n2 drain_right.t9 2.2005
R49 drain_right.n0 drain_right.t6 2.2005
R50 drain_right.n0 drain_right.t2 2.2005
R51 drain_right.n4 drain_right.t0 2.2005
R52 drain_right.n4 drain_right.t4 2.2005
R53 drain_right.n5 drain_right.t5 2.2005
R54 drain_right.n5 drain_right.t8 2.2005
R55 drain_right.n7 drain_right.n6 0.974638
R56 drain_right.n3 drain_right.n1 0.188688
R57 source.n5 source.t13 51.0588
R58 source.n19 source.t10 51.0586
R59 source.n14 source.t4 51.0586
R60 source.n0 source.t2 51.0586
R61 source.n2 source.n1 48.8588
R62 source.n4 source.n3 48.8588
R63 source.n7 source.n6 48.8588
R64 source.n9 source.n8 48.8588
R65 source.n18 source.n17 48.8586
R66 source.n16 source.n15 48.8586
R67 source.n13 source.n12 48.8586
R68 source.n11 source.n10 48.8586
R69 source.n11 source.n9 20.9633
R70 source.n20 source.n0 14.2391
R71 source.n20 source.n19 5.7505
R72 source.n17 source.t14 2.2005
R73 source.n17 source.t18 2.2005
R74 source.n15 source.t9 2.2005
R75 source.n15 source.t17 2.2005
R76 source.n12 source.t7 2.2005
R77 source.n12 source.t0 2.2005
R78 source.n10 source.t3 2.2005
R79 source.n10 source.t19 2.2005
R80 source.n1 source.t1 2.2005
R81 source.n1 source.t6 2.2005
R82 source.n3 source.t8 2.2005
R83 source.n3 source.t5 2.2005
R84 source.n6 source.t16 2.2005
R85 source.n6 source.t15 2.2005
R86 source.n8 source.t11 2.2005
R87 source.n8 source.t12 2.2005
R88 source.n9 source.n7 0.974638
R89 source.n7 source.n5 0.974638
R90 source.n4 source.n2 0.974638
R91 source.n2 source.n0 0.974638
R92 source.n13 source.n11 0.974638
R93 source.n14 source.n13 0.974638
R94 source.n18 source.n16 0.974638
R95 source.n19 source.n18 0.974638
R96 source.n5 source.n4 0.957397
R97 source.n16 source.n14 0.957397
R98 source source.n20 0.188
R99 plus.n3 plus.t9 343.425
R100 plus.n13 plus.t4 343.425
R101 plus.n8 plus.t7 320.229
R102 plus.n6 plus.t5 320.229
R103 plus.n5 plus.t6 320.229
R104 plus.n4 plus.t8 320.229
R105 plus.n18 plus.t2 320.229
R106 plus.n16 plus.t0 320.229
R107 plus.n15 plus.t3 320.229
R108 plus.n14 plus.t1 320.229
R109 plus.n7 plus.n0 161.3
R110 plus.n9 plus.n8 161.3
R111 plus.n17 plus.n10 161.3
R112 plus.n19 plus.n18 161.3
R113 plus.n5 plus.n2 80.6037
R114 plus.n6 plus.n1 80.6037
R115 plus.n15 plus.n12 80.6037
R116 plus.n16 plus.n11 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n7 plus.n6 32.1338
R122 plus.n17 plus.n16 32.1338
R123 plus.n3 plus.n2 31.8629
R124 plus.n13 plus.n12 31.8629
R125 plus plus.n19 29.8911
R126 plus.n4 plus.n3 16.2333
R127 plus.n14 plus.n13 16.2333
R128 plus.n8 plus.n7 16.0672
R129 plus.n18 plus.n17 16.0672
R130 plus plus.n9 11.1842
R131 plus.n2 plus.n1 0.380177
R132 plus.n12 plus.n11 0.380177
R133 plus.n1 plus.n0 0.285035
R134 plus.n11 plus.n10 0.285035
R135 plus.n9 plus.n0 0.189894
R136 plus.n19 plus.n10 0.189894
R137 drain_left.n5 drain_left.t0 68.7117
R138 drain_left.n1 drain_left.t7 68.7115
R139 drain_left.n3 drain_left.n2 66.2126
R140 drain_left.n5 drain_left.n4 65.5376
R141 drain_left.n7 drain_left.n6 65.5374
R142 drain_left.n1 drain_left.n0 65.5373
R143 drain_left drain_left.n3 29.2344
R144 drain_left drain_left.n7 6.62735
R145 drain_left.n2 drain_left.t8 2.2005
R146 drain_left.n2 drain_left.t5 2.2005
R147 drain_left.n0 drain_left.t9 2.2005
R148 drain_left.n0 drain_left.t6 2.2005
R149 drain_left.n6 drain_left.t4 2.2005
R150 drain_left.n6 drain_left.t2 2.2005
R151 drain_left.n4 drain_left.t1 2.2005
R152 drain_left.n4 drain_left.t3 2.2005
R153 drain_left.n7 drain_left.n5 0.974638
R154 drain_left.n3 drain_left.n1 0.188688
C0 plus minus 5.16886f
C1 plus source 5.50677f
C2 drain_left minus 0.172418f
C3 drain_right minus 5.49392f
C4 drain_left source 10.8584f
C5 drain_right source 10.854599f
C6 drain_left plus 5.69501f
C7 drain_right plus 0.359732f
C8 drain_left drain_right 1.03301f
C9 minus source 5.49237f
C10 drain_right a_n2072_n2688# 6.22573f
C11 drain_left a_n2072_n2688# 6.54087f
C12 source a_n2072_n2688# 5.528064f
C13 minus a_n2072_n2688# 7.914271f
C14 plus a_n2072_n2688# 9.40828f
C15 drain_left.t7 a_n2072_n2688# 1.90973f
C16 drain_left.t9 a_n2072_n2688# 0.171098f
C17 drain_left.t6 a_n2072_n2688# 0.171098f
C18 drain_left.n0 a_n2072_n2688# 1.49654f
C19 drain_left.n1 a_n2072_n2688# 0.617114f
C20 drain_left.t8 a_n2072_n2688# 0.171098f
C21 drain_left.t5 a_n2072_n2688# 0.171098f
C22 drain_left.n2 a_n2072_n2688# 1.49992f
C23 drain_left.n3 a_n2072_n2688# 1.42606f
C24 drain_left.t0 a_n2072_n2688# 1.90974f
C25 drain_left.t1 a_n2072_n2688# 0.171098f
C26 drain_left.t3 a_n2072_n2688# 0.171098f
C27 drain_left.n4 a_n2072_n2688# 1.49654f
C28 drain_left.n5 a_n2072_n2688# 0.67507f
C29 drain_left.t4 a_n2072_n2688# 0.171098f
C30 drain_left.t2 a_n2072_n2688# 0.171098f
C31 drain_left.n6 a_n2072_n2688# 1.49654f
C32 drain_left.n7 a_n2072_n2688# 0.559456f
C33 plus.n0 a_n2072_n2688# 0.055727f
C34 plus.t7 a_n2072_n2688# 0.862334f
C35 plus.t5 a_n2072_n2688# 0.862334f
C36 plus.n1 a_n2072_n2688# 0.069561f
C37 plus.t6 a_n2072_n2688# 0.862334f
C38 plus.n2 a_n2072_n2688# 0.256282f
C39 plus.t8 a_n2072_n2688# 0.862334f
C40 plus.t9 a_n2072_n2688# 0.886759f
C41 plus.n3 a_n2072_n2688# 0.341935f
C42 plus.n4 a_n2072_n2688# 0.370305f
C43 plus.n5 a_n2072_n2688# 0.371315f
C44 plus.n6 a_n2072_n2688# 0.368483f
C45 plus.n7 a_n2072_n2688# 0.009477f
C46 plus.n8 a_n2072_n2688# 0.356174f
C47 plus.n9 a_n2072_n2688# 0.428032f
C48 plus.n10 a_n2072_n2688# 0.055727f
C49 plus.t2 a_n2072_n2688# 0.862334f
C50 plus.n11 a_n2072_n2688# 0.069561f
C51 plus.t0 a_n2072_n2688# 0.862334f
C52 plus.n12 a_n2072_n2688# 0.256282f
C53 plus.t3 a_n2072_n2688# 0.862334f
C54 plus.t4 a_n2072_n2688# 0.886759f
C55 plus.n13 a_n2072_n2688# 0.341935f
C56 plus.t1 a_n2072_n2688# 0.862334f
C57 plus.n14 a_n2072_n2688# 0.370305f
C58 plus.n15 a_n2072_n2688# 0.371315f
C59 plus.n16 a_n2072_n2688# 0.368483f
C60 plus.n17 a_n2072_n2688# 0.009477f
C61 plus.n18 a_n2072_n2688# 0.356174f
C62 plus.n19 a_n2072_n2688# 1.22256f
C63 source.t2 a_n2072_n2688# 1.95814f
C64 source.n0 a_n2072_n2688# 1.18592f
C65 source.t1 a_n2072_n2688# 0.183631f
C66 source.t6 a_n2072_n2688# 0.183631f
C67 source.n1 a_n2072_n2688# 1.53723f
C68 source.n2 a_n2072_n2688# 0.402732f
C69 source.t8 a_n2072_n2688# 0.183631f
C70 source.t5 a_n2072_n2688# 0.183631f
C71 source.n3 a_n2072_n2688# 1.53723f
C72 source.n4 a_n2072_n2688# 0.401298f
C73 source.t13 a_n2072_n2688# 1.95814f
C74 source.n5 a_n2072_n2688# 0.481201f
C75 source.t16 a_n2072_n2688# 0.183631f
C76 source.t15 a_n2072_n2688# 0.183631f
C77 source.n6 a_n2072_n2688# 1.53723f
C78 source.n7 a_n2072_n2688# 0.402732f
C79 source.t11 a_n2072_n2688# 0.183631f
C80 source.t12 a_n2072_n2688# 0.183631f
C81 source.n8 a_n2072_n2688# 1.53723f
C82 source.n9 a_n2072_n2688# 1.574f
C83 source.t3 a_n2072_n2688# 0.183631f
C84 source.t19 a_n2072_n2688# 0.183631f
C85 source.n10 a_n2072_n2688# 1.53723f
C86 source.n11 a_n2072_n2688# 1.574f
C87 source.t7 a_n2072_n2688# 0.183631f
C88 source.t0 a_n2072_n2688# 0.183631f
C89 source.n12 a_n2072_n2688# 1.53723f
C90 source.n13 a_n2072_n2688# 0.402737f
C91 source.t4 a_n2072_n2688# 1.95814f
C92 source.n14 a_n2072_n2688# 0.481205f
C93 source.t9 a_n2072_n2688# 0.183631f
C94 source.t17 a_n2072_n2688# 0.183631f
C95 source.n15 a_n2072_n2688# 1.53723f
C96 source.n16 a_n2072_n2688# 0.401302f
C97 source.t14 a_n2072_n2688# 0.183631f
C98 source.t18 a_n2072_n2688# 0.183631f
C99 source.n17 a_n2072_n2688# 1.53723f
C100 source.n18 a_n2072_n2688# 0.402737f
C101 source.t10 a_n2072_n2688# 1.95814f
C102 source.n19 a_n2072_n2688# 0.614695f
C103 source.n20 a_n2072_n2688# 1.36347f
C104 drain_right.t1 a_n2072_n2688# 1.89748f
C105 drain_right.t6 a_n2072_n2688# 0.170001f
C106 drain_right.t2 a_n2072_n2688# 0.170001f
C107 drain_right.n0 a_n2072_n2688# 1.48694f
C108 drain_right.n1 a_n2072_n2688# 0.613155f
C109 drain_right.t7 a_n2072_n2688# 0.170001f
C110 drain_right.t9 a_n2072_n2688# 0.170001f
C111 drain_right.n2 a_n2072_n2688# 1.49029f
C112 drain_right.n3 a_n2072_n2688# 1.36788f
C113 drain_right.t0 a_n2072_n2688# 0.170001f
C114 drain_right.t4 a_n2072_n2688# 0.170001f
C115 drain_right.n4 a_n2072_n2688# 1.49208f
C116 drain_right.t5 a_n2072_n2688# 0.170001f
C117 drain_right.t8 a_n2072_n2688# 0.170001f
C118 drain_right.n5 a_n2072_n2688# 1.48694f
C119 drain_right.n6 a_n2072_n2688# 0.687536f
C120 drain_right.t3 a_n2072_n2688# 1.89275f
C121 drain_right.n7 a_n2072_n2688# 0.558641f
C122 minus.n0 a_n2072_n2688# 0.054765f
C123 minus.t2 a_n2072_n2688# 0.847454f
C124 minus.n1 a_n2072_n2688# 0.364908f
C125 minus.t6 a_n2072_n2688# 0.847454f
C126 minus.t5 a_n2072_n2688# 0.871457f
C127 minus.t3 a_n2072_n2688# 0.847454f
C128 minus.n2 a_n2072_n2688# 0.363915f
C129 minus.n3 a_n2072_n2688# 0.336035f
C130 minus.n4 a_n2072_n2688# 0.25186f
C131 minus.n5 a_n2072_n2688# 0.06836f
C132 minus.n6 a_n2072_n2688# 0.362124f
C133 minus.n7 a_n2072_n2688# 0.009313f
C134 minus.t7 a_n2072_n2688# 0.847454f
C135 minus.n8 a_n2072_n2688# 0.350028f
C136 minus.n9 a_n2072_n2688# 1.37375f
C137 minus.n10 a_n2072_n2688# 0.054765f
C138 minus.t4 a_n2072_n2688# 0.847454f
C139 minus.n11 a_n2072_n2688# 0.364908f
C140 minus.t9 a_n2072_n2688# 0.871457f
C141 minus.t1 a_n2072_n2688# 0.847454f
C142 minus.n12 a_n2072_n2688# 0.363915f
C143 minus.n13 a_n2072_n2688# 0.336035f
C144 minus.n14 a_n2072_n2688# 0.25186f
C145 minus.n15 a_n2072_n2688# 0.06836f
C146 minus.t0 a_n2072_n2688# 0.847454f
C147 minus.n16 a_n2072_n2688# 0.362124f
C148 minus.n17 a_n2072_n2688# 0.009313f
C149 minus.t8 a_n2072_n2688# 0.847454f
C150 minus.n18 a_n2072_n2688# 0.350028f
C151 minus.n19 a_n2072_n2688# 0.28526f
C152 minus.n20 a_n2072_n2688# 1.66888f
.ends

