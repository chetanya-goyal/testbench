* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t34 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 drain_left.t18 plus.t1 source.t37 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 drain_right.t19 minus.t0 source.t10 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X3 source.t12 minus.t1 drain_right.t18 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X4 drain_left.t17 plus.t2 source.t29 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X5 source.t13 minus.t2 drain_right.t17 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X6 drain_right.t16 minus.t3 source.t16 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X7 drain_left.t16 plus.t3 source.t33 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X8 source.t2 minus.t4 drain_right.t15 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X9 drain_right.t14 minus.t5 source.t7 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X10 a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X11 source.t21 plus.t4 drain_left.t15 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X12 source.t22 plus.t5 drain_left.t14 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X13 drain_left.t13 plus.t6 source.t23 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X14 drain_left.t12 plus.t7 source.t36 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X15 source.t1 minus.t6 drain_right.t13 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X16 source.t5 minus.t7 drain_right.t12 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X17 drain_left.t11 plus.t8 source.t35 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 source.t11 minus.t8 drain_right.t11 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X19 drain_left.t10 plus.t9 source.t28 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X20 source.t32 plus.t10 drain_left.t9 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X21 source.t25 plus.t11 drain_left.t8 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X22 source.t24 plus.t12 drain_left.t7 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X23 source.t26 plus.t13 drain_left.t6 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X24 a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X25 source.t18 plus.t14 drain_left.t5 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X26 source.t27 plus.t15 drain_left.t4 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X27 drain_right.t10 minus.t9 source.t15 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X28 source.t31 plus.t16 drain_left.t3 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X29 drain_right.t9 minus.t10 source.t9 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X30 drain_right.t8 minus.t11 source.t8 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X31 source.t20 plus.t17 drain_left.t2 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X32 a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X33 drain_left.t1 plus.t18 source.t19 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X34 drain_right.t7 minus.t12 source.t38 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X35 source.t39 minus.t13 drain_right.t6 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X36 drain_right.t5 minus.t14 source.t4 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X37 drain_right.t4 minus.t15 source.t0 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X38 drain_right.t3 minus.t16 source.t3 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X39 source.t17 minus.t17 drain_right.t2 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X40 drain_left.t0 plus.t19 source.t30 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X41 source.t14 minus.t18 drain_right.t1 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X42 source.t6 minus.t19 drain_right.t0 a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X43 a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# a_n1992_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
R0 plus.n6 plus.t4 467.103
R1 plus.n25 plus.t2 467.103
R2 plus.n33 plus.t7 467.103
R3 plus.n52 plus.t17 467.103
R4 plus.n5 plus.t1 414.521
R5 plus.n9 plus.t13 414.521
R6 plus.n11 plus.t0 414.521
R7 plus.n3 plus.t12 414.521
R8 plus.n17 plus.t19 414.521
R9 plus.n1 plus.t11 414.521
R10 plus.n22 plus.t3 414.521
R11 plus.n24 plus.t16 414.521
R12 plus.n32 plus.t5 414.521
R13 plus.n36 plus.t9 414.521
R14 plus.n38 plus.t15 414.521
R15 plus.n30 plus.t6 414.521
R16 plus.n44 plus.t10 414.521
R17 plus.n28 plus.t8 414.521
R18 plus.n49 plus.t14 414.521
R19 plus.n51 plus.t18 414.521
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus.n10 plus.n9 29.2126
R63 plus.n22 plus.n21 29.2126
R64 plus.n49 plus.n48 29.2126
R65 plus.n37 plus.n36 29.2126
R66 plus plus.n53 27.1354
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 8.73156
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n0 source.t29 69.6943
R93 source.n9 source.t21 69.6943
R94 source.n10 source.t9 69.6943
R95 source.n19 source.t11 69.6943
R96 source.n39 source.t7 69.6942
R97 source.n30 source.t6 69.6942
R98 source.n29 source.t36 69.6942
R99 source.n20 source.t20 69.6942
R100 source.n2 source.n1 63.0943
R101 source.n4 source.n3 63.0943
R102 source.n6 source.n5 63.0943
R103 source.n8 source.n7 63.0943
R104 source.n12 source.n11 63.0943
R105 source.n14 source.n13 63.0943
R106 source.n16 source.n15 63.0943
R107 source.n18 source.n17 63.0943
R108 source.n38 source.n37 63.0942
R109 source.n36 source.n35 63.0942
R110 source.n34 source.n33 63.0942
R111 source.n32 source.n31 63.0942
R112 source.n28 source.n27 63.0942
R113 source.n26 source.n25 63.0942
R114 source.n24 source.n23 63.0942
R115 source.n22 source.n21 63.0942
R116 source.n20 source.n19 14.9695
R117 source.n40 source.n0 9.45661
R118 source.n37 source.t10 6.6005
R119 source.n37 source.t14 6.6005
R120 source.n35 source.t16 6.6005
R121 source.n35 source.t12 6.6005
R122 source.n33 source.t38 6.6005
R123 source.n33 source.t17 6.6005
R124 source.n31 source.t8 6.6005
R125 source.n31 source.t39 6.6005
R126 source.n27 source.t28 6.6005
R127 source.n27 source.t22 6.6005
R128 source.n25 source.t23 6.6005
R129 source.n25 source.t27 6.6005
R130 source.n23 source.t35 6.6005
R131 source.n23 source.t32 6.6005
R132 source.n21 source.t19 6.6005
R133 source.n21 source.t18 6.6005
R134 source.n1 source.t33 6.6005
R135 source.n1 source.t31 6.6005
R136 source.n3 source.t30 6.6005
R137 source.n3 source.t25 6.6005
R138 source.n5 source.t34 6.6005
R139 source.n5 source.t24 6.6005
R140 source.n7 source.t37 6.6005
R141 source.n7 source.t26 6.6005
R142 source.n11 source.t15 6.6005
R143 source.n11 source.t2 6.6005
R144 source.n13 source.t4 6.6005
R145 source.n13 source.t13 6.6005
R146 source.n15 source.t0 6.6005
R147 source.n15 source.t5 6.6005
R148 source.n17 source.t3 6.6005
R149 source.n17 source.t1 6.6005
R150 source.n40 source.n39 5.51343
R151 source.n19 source.n18 0.5005
R152 source.n18 source.n16 0.5005
R153 source.n16 source.n14 0.5005
R154 source.n14 source.n12 0.5005
R155 source.n12 source.n10 0.5005
R156 source.n9 source.n8 0.5005
R157 source.n8 source.n6 0.5005
R158 source.n6 source.n4 0.5005
R159 source.n4 source.n2 0.5005
R160 source.n2 source.n0 0.5005
R161 source.n22 source.n20 0.5005
R162 source.n24 source.n22 0.5005
R163 source.n26 source.n24 0.5005
R164 source.n28 source.n26 0.5005
R165 source.n29 source.n28 0.5005
R166 source.n32 source.n30 0.5005
R167 source.n34 source.n32 0.5005
R168 source.n36 source.n34 0.5005
R169 source.n38 source.n36 0.5005
R170 source.n39 source.n38 0.5005
R171 source.n10 source.n9 0.470328
R172 source.n30 source.n29 0.470328
R173 source source.n40 0.188
R174 drain_left.n10 drain_left.n8 80.2731
R175 drain_left.n6 drain_left.n4 80.273
R176 drain_left.n2 drain_left.n0 80.273
R177 drain_left.n16 drain_left.n15 79.7731
R178 drain_left.n14 drain_left.n13 79.7731
R179 drain_left.n12 drain_left.n11 79.7731
R180 drain_left.n10 drain_left.n9 79.7731
R181 drain_left.n7 drain_left.n3 79.773
R182 drain_left.n6 drain_left.n5 79.773
R183 drain_left.n2 drain_left.n1 79.773
R184 drain_left drain_left.n7 24.5489
R185 drain_left.n3 drain_left.t9 6.6005
R186 drain_left.n3 drain_left.t13 6.6005
R187 drain_left.n4 drain_left.t14 6.6005
R188 drain_left.n4 drain_left.t12 6.6005
R189 drain_left.n5 drain_left.t4 6.6005
R190 drain_left.n5 drain_left.t10 6.6005
R191 drain_left.n1 drain_left.t5 6.6005
R192 drain_left.n1 drain_left.t11 6.6005
R193 drain_left.n0 drain_left.t2 6.6005
R194 drain_left.n0 drain_left.t1 6.6005
R195 drain_left.n15 drain_left.t3 6.6005
R196 drain_left.n15 drain_left.t17 6.6005
R197 drain_left.n13 drain_left.t8 6.6005
R198 drain_left.n13 drain_left.t16 6.6005
R199 drain_left.n11 drain_left.t7 6.6005
R200 drain_left.n11 drain_left.t0 6.6005
R201 drain_left.n9 drain_left.t6 6.6005
R202 drain_left.n9 drain_left.t19 6.6005
R203 drain_left.n8 drain_left.t15 6.6005
R204 drain_left.n8 drain_left.t18 6.6005
R205 drain_left drain_left.n16 6.15322
R206 drain_left.n12 drain_left.n10 0.5005
R207 drain_left.n14 drain_left.n12 0.5005
R208 drain_left.n16 drain_left.n14 0.5005
R209 drain_left.n7 drain_left.n6 0.445154
R210 drain_left.n7 drain_left.n2 0.445154
R211 minus.n25 minus.t8 467.103
R212 minus.n6 minus.t10 467.103
R213 minus.n52 minus.t5 467.103
R214 minus.n33 minus.t19 467.103
R215 minus.n24 minus.t16 414.521
R216 minus.n22 minus.t6 414.521
R217 minus.n1 minus.t15 414.521
R218 minus.n17 minus.t7 414.521
R219 minus.n3 minus.t14 414.521
R220 minus.n11 minus.t2 414.521
R221 minus.n9 minus.t9 414.521
R222 minus.n5 minus.t4 414.521
R223 minus.n51 minus.t18 414.521
R224 minus.n49 minus.t0 414.521
R225 minus.n28 minus.t1 414.521
R226 minus.n44 minus.t3 414.521
R227 minus.n30 minus.t17 414.521
R228 minus.n38 minus.t12 414.521
R229 minus.n36 minus.t13 414.521
R230 minus.n32 minus.t11 414.521
R231 minus.n7 minus.n6 161.489
R232 minus.n34 minus.n33 161.489
R233 minus.n26 minus.n25 161.3
R234 minus.n23 minus.n0 161.3
R235 minus.n21 minus.n20 161.3
R236 minus.n19 minus.n18 161.3
R237 minus.n16 minus.n2 161.3
R238 minus.n15 minus.n14 161.3
R239 minus.n13 minus.n12 161.3
R240 minus.n10 minus.n4 161.3
R241 minus.n8 minus.n7 161.3
R242 minus.n53 minus.n52 161.3
R243 minus.n50 minus.n27 161.3
R244 minus.n48 minus.n47 161.3
R245 minus.n46 minus.n45 161.3
R246 minus.n43 minus.n29 161.3
R247 minus.n42 minus.n41 161.3
R248 minus.n40 minus.n39 161.3
R249 minus.n37 minus.n31 161.3
R250 minus.n35 minus.n34 161.3
R251 minus.n16 minus.n15 73.0308
R252 minus.n43 minus.n42 73.0308
R253 minus.n18 minus.n17 67.1884
R254 minus.n12 minus.n3 67.1884
R255 minus.n39 minus.n30 67.1884
R256 minus.n45 minus.n44 67.1884
R257 minus.n21 minus.n1 55.5035
R258 minus.n11 minus.n10 55.5035
R259 minus.n38 minus.n37 55.5035
R260 minus.n48 minus.n28 55.5035
R261 minus.n23 minus.n22 43.8187
R262 minus.n9 minus.n8 43.8187
R263 minus.n36 minus.n35 43.8187
R264 minus.n50 minus.n49 43.8187
R265 minus.n24 minus.n23 40.8975
R266 minus.n8 minus.n5 40.8975
R267 minus.n35 minus.n32 40.8975
R268 minus.n51 minus.n50 40.8975
R269 minus.n25 minus.n24 32.1338
R270 minus.n6 minus.n5 32.1338
R271 minus.n33 minus.n32 32.1338
R272 minus.n52 minus.n51 32.1338
R273 minus.n54 minus.n26 29.8452
R274 minus.n22 minus.n21 29.2126
R275 minus.n10 minus.n9 29.2126
R276 minus.n37 minus.n36 29.2126
R277 minus.n49 minus.n48 29.2126
R278 minus.n18 minus.n1 17.5278
R279 minus.n12 minus.n11 17.5278
R280 minus.n39 minus.n38 17.5278
R281 minus.n45 minus.n28 17.5278
R282 minus.n54 minus.n53 6.49671
R283 minus.n17 minus.n16 5.84292
R284 minus.n15 minus.n3 5.84292
R285 minus.n42 minus.n30 5.84292
R286 minus.n44 minus.n43 5.84292
R287 minus.n26 minus.n0 0.189894
R288 minus.n20 minus.n0 0.189894
R289 minus.n20 minus.n19 0.189894
R290 minus.n19 minus.n2 0.189894
R291 minus.n14 minus.n2 0.189894
R292 minus.n14 minus.n13 0.189894
R293 minus.n13 minus.n4 0.189894
R294 minus.n7 minus.n4 0.189894
R295 minus.n34 minus.n31 0.189894
R296 minus.n40 minus.n31 0.189894
R297 minus.n41 minus.n40 0.189894
R298 minus.n41 minus.n29 0.189894
R299 minus.n46 minus.n29 0.189894
R300 minus.n47 minus.n46 0.189894
R301 minus.n47 minus.n27 0.189894
R302 minus.n53 minus.n27 0.189894
R303 minus minus.n54 0.188
R304 drain_right.n10 drain_right.n8 80.2731
R305 drain_right.n6 drain_right.n4 80.273
R306 drain_right.n2 drain_right.n0 80.273
R307 drain_right.n10 drain_right.n9 79.7731
R308 drain_right.n12 drain_right.n11 79.7731
R309 drain_right.n14 drain_right.n13 79.7731
R310 drain_right.n16 drain_right.n15 79.7731
R311 drain_right.n7 drain_right.n3 79.773
R312 drain_right.n6 drain_right.n5 79.773
R313 drain_right.n2 drain_right.n1 79.773
R314 drain_right drain_right.n7 23.9957
R315 drain_right.n3 drain_right.t2 6.6005
R316 drain_right.n3 drain_right.t16 6.6005
R317 drain_right.n4 drain_right.t1 6.6005
R318 drain_right.n4 drain_right.t14 6.6005
R319 drain_right.n5 drain_right.t18 6.6005
R320 drain_right.n5 drain_right.t19 6.6005
R321 drain_right.n1 drain_right.t6 6.6005
R322 drain_right.n1 drain_right.t7 6.6005
R323 drain_right.n0 drain_right.t0 6.6005
R324 drain_right.n0 drain_right.t8 6.6005
R325 drain_right.n8 drain_right.t15 6.6005
R326 drain_right.n8 drain_right.t9 6.6005
R327 drain_right.n9 drain_right.t17 6.6005
R328 drain_right.n9 drain_right.t10 6.6005
R329 drain_right.n11 drain_right.t12 6.6005
R330 drain_right.n11 drain_right.t5 6.6005
R331 drain_right.n13 drain_right.t13 6.6005
R332 drain_right.n13 drain_right.t4 6.6005
R333 drain_right.n15 drain_right.t11 6.6005
R334 drain_right.n15 drain_right.t3 6.6005
R335 drain_right drain_right.n16 6.15322
R336 drain_right.n16 drain_right.n14 0.5005
R337 drain_right.n14 drain_right.n12 0.5005
R338 drain_right.n12 drain_right.n10 0.5005
R339 drain_right.n7 drain_right.n6 0.445154
R340 drain_right.n7 drain_right.n2 0.445154
C0 drain_right source 12.6508f
C1 source plus 2.18429f
C2 source drain_left 12.650499f
C3 drain_right plus 0.354786f
C4 drain_right drain_left 1.04655f
C5 drain_left plus 2.20113f
C6 source minus 2.17029f
C7 drain_right minus 2.00664f
C8 minus plus 3.9782f
C9 drain_left minus 0.176785f
C10 drain_right a_n1992_n1488# 4.82941f
C11 drain_left a_n1992_n1488# 5.1444f
C12 source a_n1992_n1488# 3.749464f
C13 minus a_n1992_n1488# 7.064308f
C14 plus a_n1992_n1488# 8.5042f
C15 drain_right.t0 a_n1992_n1488# 0.08142f
C16 drain_right.t8 a_n1992_n1488# 0.08142f
C17 drain_right.n0 a_n1992_n1488# 0.589681f
C18 drain_right.t6 a_n1992_n1488# 0.08142f
C19 drain_right.t7 a_n1992_n1488# 0.08142f
C20 drain_right.n1 a_n1992_n1488# 0.587193f
C21 drain_right.n2 a_n1992_n1488# 0.778186f
C22 drain_right.t2 a_n1992_n1488# 0.08142f
C23 drain_right.t16 a_n1992_n1488# 0.08142f
C24 drain_right.n3 a_n1992_n1488# 0.587193f
C25 drain_right.t1 a_n1992_n1488# 0.08142f
C26 drain_right.t14 a_n1992_n1488# 0.08142f
C27 drain_right.n4 a_n1992_n1488# 0.589681f
C28 drain_right.t18 a_n1992_n1488# 0.08142f
C29 drain_right.t19 a_n1992_n1488# 0.08142f
C30 drain_right.n5 a_n1992_n1488# 0.587193f
C31 drain_right.n6 a_n1992_n1488# 0.778186f
C32 drain_right.n7 a_n1992_n1488# 1.35165f
C33 drain_right.t15 a_n1992_n1488# 0.08142f
C34 drain_right.t9 a_n1992_n1488# 0.08142f
C35 drain_right.n8 a_n1992_n1488# 0.589684f
C36 drain_right.t17 a_n1992_n1488# 0.08142f
C37 drain_right.t10 a_n1992_n1488# 0.08142f
C38 drain_right.n9 a_n1992_n1488# 0.587196f
C39 drain_right.n10 a_n1992_n1488# 0.782515f
C40 drain_right.t12 a_n1992_n1488# 0.08142f
C41 drain_right.t5 a_n1992_n1488# 0.08142f
C42 drain_right.n11 a_n1992_n1488# 0.587196f
C43 drain_right.n12 a_n1992_n1488# 0.385585f
C44 drain_right.t13 a_n1992_n1488# 0.08142f
C45 drain_right.t4 a_n1992_n1488# 0.08142f
C46 drain_right.n13 a_n1992_n1488# 0.587196f
C47 drain_right.n14 a_n1992_n1488# 0.385585f
C48 drain_right.t11 a_n1992_n1488# 0.08142f
C49 drain_right.t3 a_n1992_n1488# 0.08142f
C50 drain_right.n15 a_n1992_n1488# 0.587196f
C51 drain_right.n16 a_n1992_n1488# 0.669075f
C52 minus.n0 a_n1992_n1488# 0.05098f
C53 minus.t8 a_n1992_n1488# 0.118645f
C54 minus.t16 a_n1992_n1488# 0.110723f
C55 minus.t6 a_n1992_n1488# 0.110723f
C56 minus.t15 a_n1992_n1488# 0.110723f
C57 minus.n1 a_n1992_n1488# 0.06691f
C58 minus.n2 a_n1992_n1488# 0.05098f
C59 minus.t7 a_n1992_n1488# 0.110723f
C60 minus.t14 a_n1992_n1488# 0.110723f
C61 minus.n3 a_n1992_n1488# 0.06691f
C62 minus.n4 a_n1992_n1488# 0.05098f
C63 minus.t2 a_n1992_n1488# 0.110723f
C64 minus.t9 a_n1992_n1488# 0.110723f
C65 minus.t4 a_n1992_n1488# 0.110723f
C66 minus.n5 a_n1992_n1488# 0.06691f
C67 minus.t10 a_n1992_n1488# 0.118645f
C68 minus.n6 a_n1992_n1488# 0.081949f
C69 minus.n7 a_n1992_n1488# 0.116655f
C70 minus.n8 a_n1992_n1488# 0.019426f
C71 minus.n9 a_n1992_n1488# 0.06691f
C72 minus.n10 a_n1992_n1488# 0.019426f
C73 minus.n11 a_n1992_n1488# 0.06691f
C74 minus.n12 a_n1992_n1488# 0.019426f
C75 minus.n13 a_n1992_n1488# 0.05098f
C76 minus.n14 a_n1992_n1488# 0.05098f
C77 minus.n15 a_n1992_n1488# 0.018169f
C78 minus.n16 a_n1992_n1488# 0.018169f
C79 minus.n17 a_n1992_n1488# 0.06691f
C80 minus.n18 a_n1992_n1488# 0.019426f
C81 minus.n19 a_n1992_n1488# 0.05098f
C82 minus.n20 a_n1992_n1488# 0.05098f
C83 minus.n21 a_n1992_n1488# 0.019426f
C84 minus.n22 a_n1992_n1488# 0.06691f
C85 minus.n23 a_n1992_n1488# 0.019426f
C86 minus.n24 a_n1992_n1488# 0.06691f
C87 minus.n25 a_n1992_n1488# 0.081872f
C88 minus.n26 a_n1992_n1488# 1.31436f
C89 minus.n27 a_n1992_n1488# 0.05098f
C90 minus.t18 a_n1992_n1488# 0.110723f
C91 minus.t0 a_n1992_n1488# 0.110723f
C92 minus.t1 a_n1992_n1488# 0.110723f
C93 minus.n28 a_n1992_n1488# 0.06691f
C94 minus.n29 a_n1992_n1488# 0.05098f
C95 minus.t3 a_n1992_n1488# 0.110723f
C96 minus.t17 a_n1992_n1488# 0.110723f
C97 minus.n30 a_n1992_n1488# 0.06691f
C98 minus.n31 a_n1992_n1488# 0.05098f
C99 minus.t12 a_n1992_n1488# 0.110723f
C100 minus.t13 a_n1992_n1488# 0.110723f
C101 minus.t11 a_n1992_n1488# 0.110723f
C102 minus.n32 a_n1992_n1488# 0.06691f
C103 minus.t19 a_n1992_n1488# 0.118645f
C104 minus.n33 a_n1992_n1488# 0.081949f
C105 minus.n34 a_n1992_n1488# 0.116655f
C106 minus.n35 a_n1992_n1488# 0.019426f
C107 minus.n36 a_n1992_n1488# 0.06691f
C108 minus.n37 a_n1992_n1488# 0.019426f
C109 minus.n38 a_n1992_n1488# 0.06691f
C110 minus.n39 a_n1992_n1488# 0.019426f
C111 minus.n40 a_n1992_n1488# 0.05098f
C112 minus.n41 a_n1992_n1488# 0.05098f
C113 minus.n42 a_n1992_n1488# 0.018169f
C114 minus.n43 a_n1992_n1488# 0.018169f
C115 minus.n44 a_n1992_n1488# 0.06691f
C116 minus.n45 a_n1992_n1488# 0.019426f
C117 minus.n46 a_n1992_n1488# 0.05098f
C118 minus.n47 a_n1992_n1488# 0.05098f
C119 minus.n48 a_n1992_n1488# 0.019426f
C120 minus.n49 a_n1992_n1488# 0.06691f
C121 minus.n50 a_n1992_n1488# 0.019426f
C122 minus.n51 a_n1992_n1488# 0.06691f
C123 minus.t5 a_n1992_n1488# 0.118645f
C124 minus.n52 a_n1992_n1488# 0.081872f
C125 minus.n53 a_n1992_n1488# 0.332897f
C126 minus.n54 a_n1992_n1488# 1.6221f
C127 drain_left.t2 a_n1992_n1488# 0.08178f
C128 drain_left.t1 a_n1992_n1488# 0.08178f
C129 drain_left.n0 a_n1992_n1488# 0.592291f
C130 drain_left.t5 a_n1992_n1488# 0.08178f
C131 drain_left.t11 a_n1992_n1488# 0.08178f
C132 drain_left.n1 a_n1992_n1488# 0.589792f
C133 drain_left.n2 a_n1992_n1488# 0.78163f
C134 drain_left.t9 a_n1992_n1488# 0.08178f
C135 drain_left.t13 a_n1992_n1488# 0.08178f
C136 drain_left.n3 a_n1992_n1488# 0.589792f
C137 drain_left.t14 a_n1992_n1488# 0.08178f
C138 drain_left.t12 a_n1992_n1488# 0.08178f
C139 drain_left.n4 a_n1992_n1488# 0.592291f
C140 drain_left.t4 a_n1992_n1488# 0.08178f
C141 drain_left.t10 a_n1992_n1488# 0.08178f
C142 drain_left.n5 a_n1992_n1488# 0.589792f
C143 drain_left.n6 a_n1992_n1488# 0.78163f
C144 drain_left.n7 a_n1992_n1488# 1.42585f
C145 drain_left.t15 a_n1992_n1488# 0.08178f
C146 drain_left.t18 a_n1992_n1488# 0.08178f
C147 drain_left.n8 a_n1992_n1488# 0.592294f
C148 drain_left.t6 a_n1992_n1488# 0.08178f
C149 drain_left.t19 a_n1992_n1488# 0.08178f
C150 drain_left.n9 a_n1992_n1488# 0.589795f
C151 drain_left.n10 a_n1992_n1488# 0.785978f
C152 drain_left.t7 a_n1992_n1488# 0.08178f
C153 drain_left.t0 a_n1992_n1488# 0.08178f
C154 drain_left.n11 a_n1992_n1488# 0.589795f
C155 drain_left.n12 a_n1992_n1488# 0.387291f
C156 drain_left.t8 a_n1992_n1488# 0.08178f
C157 drain_left.t16 a_n1992_n1488# 0.08178f
C158 drain_left.n13 a_n1992_n1488# 0.589795f
C159 drain_left.n14 a_n1992_n1488# 0.387291f
C160 drain_left.t3 a_n1992_n1488# 0.08178f
C161 drain_left.t17 a_n1992_n1488# 0.08178f
C162 drain_left.n15 a_n1992_n1488# 0.589795f
C163 drain_left.n16 a_n1992_n1488# 0.672036f
C164 source.t29 a_n1992_n1488# 0.674458f
C165 source.n0 a_n1992_n1488# 0.911803f
C166 source.t33 a_n1992_n1488# 0.081223f
C167 source.t31 a_n1992_n1488# 0.081223f
C168 source.n1 a_n1992_n1488# 0.514998f
C169 source.n2 a_n1992_n1488# 0.408856f
C170 source.t30 a_n1992_n1488# 0.081223f
C171 source.t25 a_n1992_n1488# 0.081223f
C172 source.n3 a_n1992_n1488# 0.514998f
C173 source.n4 a_n1992_n1488# 0.408856f
C174 source.t34 a_n1992_n1488# 0.081223f
C175 source.t24 a_n1992_n1488# 0.081223f
C176 source.n5 a_n1992_n1488# 0.514998f
C177 source.n6 a_n1992_n1488# 0.408856f
C178 source.t37 a_n1992_n1488# 0.081223f
C179 source.t26 a_n1992_n1488# 0.081223f
C180 source.n7 a_n1992_n1488# 0.514998f
C181 source.n8 a_n1992_n1488# 0.408856f
C182 source.t21 a_n1992_n1488# 0.674458f
C183 source.n9 a_n1992_n1488# 0.467581f
C184 source.t9 a_n1992_n1488# 0.674458f
C185 source.n10 a_n1992_n1488# 0.467581f
C186 source.t15 a_n1992_n1488# 0.081223f
C187 source.t2 a_n1992_n1488# 0.081223f
C188 source.n11 a_n1992_n1488# 0.514998f
C189 source.n12 a_n1992_n1488# 0.408856f
C190 source.t4 a_n1992_n1488# 0.081223f
C191 source.t13 a_n1992_n1488# 0.081223f
C192 source.n13 a_n1992_n1488# 0.514998f
C193 source.n14 a_n1992_n1488# 0.408856f
C194 source.t0 a_n1992_n1488# 0.081223f
C195 source.t5 a_n1992_n1488# 0.081223f
C196 source.n15 a_n1992_n1488# 0.514998f
C197 source.n16 a_n1992_n1488# 0.408856f
C198 source.t3 a_n1992_n1488# 0.081223f
C199 source.t1 a_n1992_n1488# 0.081223f
C200 source.n17 a_n1992_n1488# 0.514998f
C201 source.n18 a_n1992_n1488# 0.408856f
C202 source.t11 a_n1992_n1488# 0.674458f
C203 source.n19 a_n1992_n1488# 1.2678f
C204 source.t20 a_n1992_n1488# 0.674455f
C205 source.n20 a_n1992_n1488# 1.2678f
C206 source.t19 a_n1992_n1488# 0.081223f
C207 source.t18 a_n1992_n1488# 0.081223f
C208 source.n21 a_n1992_n1488# 0.514994f
C209 source.n22 a_n1992_n1488# 0.40886f
C210 source.t35 a_n1992_n1488# 0.081223f
C211 source.t32 a_n1992_n1488# 0.081223f
C212 source.n23 a_n1992_n1488# 0.514994f
C213 source.n24 a_n1992_n1488# 0.40886f
C214 source.t23 a_n1992_n1488# 0.081223f
C215 source.t27 a_n1992_n1488# 0.081223f
C216 source.n25 a_n1992_n1488# 0.514994f
C217 source.n26 a_n1992_n1488# 0.40886f
C218 source.t28 a_n1992_n1488# 0.081223f
C219 source.t22 a_n1992_n1488# 0.081223f
C220 source.n27 a_n1992_n1488# 0.514994f
C221 source.n28 a_n1992_n1488# 0.40886f
C222 source.t36 a_n1992_n1488# 0.674455f
C223 source.n29 a_n1992_n1488# 0.467584f
C224 source.t6 a_n1992_n1488# 0.674455f
C225 source.n30 a_n1992_n1488# 0.467584f
C226 source.t8 a_n1992_n1488# 0.081223f
C227 source.t39 a_n1992_n1488# 0.081223f
C228 source.n31 a_n1992_n1488# 0.514994f
C229 source.n32 a_n1992_n1488# 0.40886f
C230 source.t38 a_n1992_n1488# 0.081223f
C231 source.t17 a_n1992_n1488# 0.081223f
C232 source.n33 a_n1992_n1488# 0.514994f
C233 source.n34 a_n1992_n1488# 0.40886f
C234 source.t16 a_n1992_n1488# 0.081223f
C235 source.t12 a_n1992_n1488# 0.081223f
C236 source.n35 a_n1992_n1488# 0.514994f
C237 source.n36 a_n1992_n1488# 0.40886f
C238 source.t10 a_n1992_n1488# 0.081223f
C239 source.t14 a_n1992_n1488# 0.081223f
C240 source.n37 a_n1992_n1488# 0.514994f
C241 source.n38 a_n1992_n1488# 0.40886f
C242 source.t7 a_n1992_n1488# 0.674455f
C243 source.n39 a_n1992_n1488# 0.657179f
C244 source.n40 a_n1992_n1488# 0.990982f
C245 plus.n0 a_n1992_n1488# 0.052888f
C246 plus.t16 a_n1992_n1488# 0.114868f
C247 plus.t3 a_n1992_n1488# 0.114868f
C248 plus.t11 a_n1992_n1488# 0.114868f
C249 plus.n1 a_n1992_n1488# 0.069415f
C250 plus.n2 a_n1992_n1488# 0.052888f
C251 plus.t19 a_n1992_n1488# 0.114868f
C252 plus.t12 a_n1992_n1488# 0.114868f
C253 plus.n3 a_n1992_n1488# 0.069415f
C254 plus.n4 a_n1992_n1488# 0.052888f
C255 plus.t0 a_n1992_n1488# 0.114868f
C256 plus.t13 a_n1992_n1488# 0.114868f
C257 plus.t1 a_n1992_n1488# 0.114868f
C258 plus.n5 a_n1992_n1488# 0.069415f
C259 plus.t4 a_n1992_n1488# 0.123086f
C260 plus.n6 a_n1992_n1488# 0.085017f
C261 plus.n7 a_n1992_n1488# 0.121022f
C262 plus.n8 a_n1992_n1488# 0.020153f
C263 plus.n9 a_n1992_n1488# 0.069415f
C264 plus.n10 a_n1992_n1488# 0.020153f
C265 plus.n11 a_n1992_n1488# 0.069415f
C266 plus.n12 a_n1992_n1488# 0.020153f
C267 plus.n13 a_n1992_n1488# 0.052888f
C268 plus.n14 a_n1992_n1488# 0.052888f
C269 plus.n15 a_n1992_n1488# 0.018849f
C270 plus.n16 a_n1992_n1488# 0.018849f
C271 plus.n17 a_n1992_n1488# 0.069415f
C272 plus.n18 a_n1992_n1488# 0.020153f
C273 plus.n19 a_n1992_n1488# 0.052888f
C274 plus.n20 a_n1992_n1488# 0.052888f
C275 plus.n21 a_n1992_n1488# 0.020153f
C276 plus.n22 a_n1992_n1488# 0.069415f
C277 plus.n23 a_n1992_n1488# 0.020153f
C278 plus.n24 a_n1992_n1488# 0.069415f
C279 plus.t2 a_n1992_n1488# 0.123086f
C280 plus.n25 a_n1992_n1488# 0.084937f
C281 plus.n26 a_n1992_n1488# 0.394636f
C282 plus.n27 a_n1992_n1488# 0.052888f
C283 plus.t17 a_n1992_n1488# 0.123086f
C284 plus.t18 a_n1992_n1488# 0.114868f
C285 plus.t14 a_n1992_n1488# 0.114868f
C286 plus.t8 a_n1992_n1488# 0.114868f
C287 plus.n28 a_n1992_n1488# 0.069415f
C288 plus.n29 a_n1992_n1488# 0.052888f
C289 plus.t10 a_n1992_n1488# 0.114868f
C290 plus.t6 a_n1992_n1488# 0.114868f
C291 plus.n30 a_n1992_n1488# 0.069415f
C292 plus.n31 a_n1992_n1488# 0.052888f
C293 plus.t15 a_n1992_n1488# 0.114868f
C294 plus.t9 a_n1992_n1488# 0.114868f
C295 plus.t5 a_n1992_n1488# 0.114868f
C296 plus.n32 a_n1992_n1488# 0.069415f
C297 plus.t7 a_n1992_n1488# 0.123086f
C298 plus.n33 a_n1992_n1488# 0.085017f
C299 plus.n34 a_n1992_n1488# 0.121022f
C300 plus.n35 a_n1992_n1488# 0.020153f
C301 plus.n36 a_n1992_n1488# 0.069415f
C302 plus.n37 a_n1992_n1488# 0.020153f
C303 plus.n38 a_n1992_n1488# 0.069415f
C304 plus.n39 a_n1992_n1488# 0.020153f
C305 plus.n40 a_n1992_n1488# 0.052888f
C306 plus.n41 a_n1992_n1488# 0.052888f
C307 plus.n42 a_n1992_n1488# 0.018849f
C308 plus.n43 a_n1992_n1488# 0.018849f
C309 plus.n44 a_n1992_n1488# 0.069415f
C310 plus.n45 a_n1992_n1488# 0.020153f
C311 plus.n46 a_n1992_n1488# 0.052888f
C312 plus.n47 a_n1992_n1488# 0.052888f
C313 plus.n48 a_n1992_n1488# 0.020153f
C314 plus.n49 a_n1992_n1488# 0.069415f
C315 plus.n50 a_n1992_n1488# 0.020153f
C316 plus.n51 a_n1992_n1488# 0.069415f
C317 plus.n52 a_n1992_n1488# 0.084937f
C318 plus.n53 a_n1992_n1488# 1.28155f
.ends

