* NGSPICE file created from diffpair157.ext - technology: sky130A

.subckt diffpair157 minus drain_right drain_left source plus
X0 a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X1 source.t17 plus.t0 drain_left.t10 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X2 drain_right.t15 minus.t0 source.t19 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X4 a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X5 drain_right.t14 minus.t1 source.t1 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X6 a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X7 drain_right.t13 minus.t2 source.t20 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X8 drain_right.t12 minus.t3 source.t18 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X9 source.t16 plus.t1 drain_left.t11 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X10 source.t15 plus.t2 drain_left.t1 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X11 source.t14 plus.t3 drain_left.t5 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X12 drain_right.t11 minus.t4 source.t0 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X13 source.t30 minus.t5 drain_right.t10 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X14 drain_right.t9 minus.t6 source.t28 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X15 drain_right.t8 minus.t7 source.t25 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X16 source.t26 minus.t8 drain_right.t7 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X17 source.t27 minus.t9 drain_right.t6 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X18 source.t31 minus.t10 drain_right.t5 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X19 drain_left.t15 plus.t4 source.t13 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X20 drain_left.t2 plus.t5 source.t12 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X21 source.t29 minus.t11 drain_right.t4 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X22 drain_left.t12 plus.t6 source.t11 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X23 drain_right.t3 minus.t12 source.t24 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X24 source.t10 plus.t7 drain_left.t8 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X25 drain_left.t3 plus.t8 source.t9 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X26 drain_left.t6 plus.t9 source.t8 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X27 source.t22 minus.t13 drain_right.t2 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X28 source.t21 minus.t14 drain_right.t1 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X29 source.t7 plus.t10 drain_left.t13 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X30 source.t23 minus.t15 drain_right.t0 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X31 source.t6 plus.t11 drain_left.t4 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X32 drain_left.t9 plus.t12 source.t5 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X33 drain_left.t7 plus.t13 source.t4 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X34 source.t3 plus.t14 drain_left.t0 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X35 drain_left.t14 plus.t15 source.t2 a_n2750_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 plus.n10 plus.n9 161.3
R1 plus.n11 plus.n4 161.3
R2 plus.n13 plus.n12 161.3
R3 plus.n14 plus.n3 161.3
R4 plus.n16 plus.n15 161.3
R5 plus.n19 plus.n0 161.3
R6 plus.n21 plus.n20 161.3
R7 plus.n32 plus.n31 161.3
R8 plus.n33 plus.n26 161.3
R9 plus.n35 plus.n34 161.3
R10 plus.n36 plus.n25 161.3
R11 plus.n38 plus.n37 161.3
R12 plus.n41 plus.n22 161.3
R13 plus.n43 plus.n42 161.3
R14 plus.n7 plus.t14 130.377
R15 plus.n29 plus.t13 130.377
R16 plus.n20 plus.t5 109.355
R17 plus.n18 plus.t7 109.355
R18 plus.n17 plus.t8 109.355
R19 plus.n3 plus.t11 109.355
R20 plus.n11 plus.t9 109.355
R21 plus.n5 plus.t10 109.355
R22 plus.n6 plus.t12 109.355
R23 plus.n42 plus.t0 109.355
R24 plus.n40 plus.t6 109.355
R25 plus.n39 plus.t3 109.355
R26 plus.n25 plus.t4 109.355
R27 plus.n33 plus.t2 109.355
R28 plus.n27 plus.t15 109.355
R29 plus.n28 plus.t1 109.355
R30 plus.n8 plus.n5 80.6037
R31 plus.n17 plus.n2 80.6037
R32 plus.n18 plus.n1 80.6037
R33 plus.n30 plus.n27 80.6037
R34 plus.n39 plus.n24 80.6037
R35 plus.n40 plus.n23 80.6037
R36 plus.n18 plus.n17 48.2005
R37 plus.n6 plus.n5 48.2005
R38 plus.n40 plus.n39 48.2005
R39 plus.n28 plus.n27 48.2005
R40 plus.n17 plus.n16 43.0884
R41 plus.n10 plus.n5 43.0884
R42 plus.n39 plus.n38 43.0884
R43 plus.n32 plus.n27 43.0884
R44 plus.n19 plus.n18 40.1672
R45 plus.n41 plus.n40 40.1672
R46 plus.n8 plus.n7 31.6481
R47 plus.n30 plus.n29 31.6481
R48 plus plus.n43 29.7869
R49 plus.n12 plus.n11 24.1005
R50 plus.n12 plus.n3 24.1005
R51 plus.n34 plus.n25 24.1005
R52 plus.n34 plus.n33 24.1005
R53 plus.n7 plus.n6 17.444
R54 plus.n29 plus.n28 17.444
R55 plus plus.n21 8.51186
R56 plus.n20 plus.n19 8.03383
R57 plus.n42 plus.n41 8.03383
R58 plus.n16 plus.n3 5.11262
R59 plus.n11 plus.n10 5.11262
R60 plus.n38 plus.n25 5.11262
R61 plus.n33 plus.n32 5.11262
R62 plus.n2 plus.n1 0.380177
R63 plus.n24 plus.n23 0.380177
R64 plus.n9 plus.n8 0.285035
R65 plus.n15 plus.n2 0.285035
R66 plus.n1 plus.n0 0.285035
R67 plus.n23 plus.n22 0.285035
R68 plus.n37 plus.n24 0.285035
R69 plus.n31 plus.n30 0.285035
R70 plus.n9 plus.n4 0.189894
R71 plus.n13 plus.n4 0.189894
R72 plus.n14 plus.n13 0.189894
R73 plus.n15 plus.n14 0.189894
R74 plus.n21 plus.n0 0.189894
R75 plus.n43 plus.n22 0.189894
R76 plus.n37 plus.n36 0.189894
R77 plus.n36 plus.n35 0.189894
R78 plus.n35 plus.n26 0.189894
R79 plus.n31 plus.n26 0.189894
R80 drain_left.n9 drain_left.n7 101.769
R81 drain_left.n5 drain_left.n3 101.769
R82 drain_left.n2 drain_left.n0 101.769
R83 drain_left.n13 drain_left.n12 100.796
R84 drain_left.n11 drain_left.n10 100.796
R85 drain_left.n9 drain_left.n8 100.796
R86 drain_left.n5 drain_left.n4 100.796
R87 drain_left.n2 drain_left.n1 100.796
R88 drain_left drain_left.n6 26.1232
R89 drain_left.n3 drain_left.t11 9.9005
R90 drain_left.n3 drain_left.t7 9.9005
R91 drain_left.n4 drain_left.t1 9.9005
R92 drain_left.n4 drain_left.t14 9.9005
R93 drain_left.n1 drain_left.t5 9.9005
R94 drain_left.n1 drain_left.t15 9.9005
R95 drain_left.n0 drain_left.t10 9.9005
R96 drain_left.n0 drain_left.t12 9.9005
R97 drain_left.n12 drain_left.t8 9.9005
R98 drain_left.n12 drain_left.t2 9.9005
R99 drain_left.n10 drain_left.t4 9.9005
R100 drain_left.n10 drain_left.t3 9.9005
R101 drain_left.n8 drain_left.t13 9.9005
R102 drain_left.n8 drain_left.t6 9.9005
R103 drain_left.n7 drain_left.t0 9.9005
R104 drain_left.n7 drain_left.t9 9.9005
R105 drain_left drain_left.n13 6.62735
R106 drain_left.n11 drain_left.n9 0.974638
R107 drain_left.n13 drain_left.n11 0.974638
R108 drain_left.n6 drain_left.n5 0.432223
R109 drain_left.n6 drain_left.n2 0.432223
R110 source.n82 source.n80 289.615
R111 source.n68 source.n66 289.615
R112 source.n60 source.n58 289.615
R113 source.n46 source.n44 289.615
R114 source.n2 source.n0 289.615
R115 source.n16 source.n14 289.615
R116 source.n24 source.n22 289.615
R117 source.n38 source.n36 289.615
R118 source.n83 source.n82 185
R119 source.n69 source.n68 185
R120 source.n61 source.n60 185
R121 source.n47 source.n46 185
R122 source.n3 source.n2 185
R123 source.n17 source.n16 185
R124 source.n25 source.n24 185
R125 source.n39 source.n38 185
R126 source.t18 source.n81 167.117
R127 source.t21 source.n67 167.117
R128 source.t4 source.n59 167.117
R129 source.t17 source.n45 167.117
R130 source.t12 source.n1 167.117
R131 source.t3 source.n15 167.117
R132 source.t25 source.n23 167.117
R133 source.t22 source.n37 167.117
R134 source.n9 source.n8 84.1169
R135 source.n11 source.n10 84.1169
R136 source.n13 source.n12 84.1169
R137 source.n31 source.n30 84.1169
R138 source.n33 source.n32 84.1169
R139 source.n35 source.n34 84.1169
R140 source.n79 source.n78 84.1168
R141 source.n77 source.n76 84.1168
R142 source.n75 source.n74 84.1168
R143 source.n57 source.n56 84.1168
R144 source.n55 source.n54 84.1168
R145 source.n53 source.n52 84.1168
R146 source.n82 source.t18 52.3082
R147 source.n68 source.t21 52.3082
R148 source.n60 source.t4 52.3082
R149 source.n46 source.t17 52.3082
R150 source.n2 source.t12 52.3082
R151 source.n16 source.t3 52.3082
R152 source.n24 source.t25 52.3082
R153 source.n38 source.t22 52.3082
R154 source.n87 source.n86 31.4096
R155 source.n73 source.n72 31.4096
R156 source.n65 source.n64 31.4096
R157 source.n51 source.n50 31.4096
R158 source.n7 source.n6 31.4096
R159 source.n21 source.n20 31.4096
R160 source.n29 source.n28 31.4096
R161 source.n43 source.n42 31.4096
R162 source.n51 source.n43 14.6861
R163 source.n78 source.t20 9.9005
R164 source.n78 source.t31 9.9005
R165 source.n76 source.t1 9.9005
R166 source.n76 source.t26 9.9005
R167 source.n74 source.t19 9.9005
R168 source.n74 source.t23 9.9005
R169 source.n56 source.t2 9.9005
R170 source.n56 source.t16 9.9005
R171 source.n54 source.t13 9.9005
R172 source.n54 source.t15 9.9005
R173 source.n52 source.t11 9.9005
R174 source.n52 source.t14 9.9005
R175 source.n8 source.t9 9.9005
R176 source.n8 source.t10 9.9005
R177 source.n10 source.t8 9.9005
R178 source.n10 source.t6 9.9005
R179 source.n12 source.t5 9.9005
R180 source.n12 source.t7 9.9005
R181 source.n30 source.t0 9.9005
R182 source.n30 source.t30 9.9005
R183 source.n32 source.t24 9.9005
R184 source.n32 source.t29 9.9005
R185 source.n34 source.t28 9.9005
R186 source.n34 source.t27 9.9005
R187 source.n83 source.n81 9.71174
R188 source.n69 source.n67 9.71174
R189 source.n61 source.n59 9.71174
R190 source.n47 source.n45 9.71174
R191 source.n3 source.n1 9.71174
R192 source.n17 source.n15 9.71174
R193 source.n25 source.n23 9.71174
R194 source.n39 source.n37 9.71174
R195 source.n86 source.n85 9.45567
R196 source.n72 source.n71 9.45567
R197 source.n64 source.n63 9.45567
R198 source.n50 source.n49 9.45567
R199 source.n6 source.n5 9.45567
R200 source.n20 source.n19 9.45567
R201 source.n28 source.n27 9.45567
R202 source.n42 source.n41 9.45567
R203 source.n85 source.n84 9.3005
R204 source.n71 source.n70 9.3005
R205 source.n63 source.n62 9.3005
R206 source.n49 source.n48 9.3005
R207 source.n5 source.n4 9.3005
R208 source.n19 source.n18 9.3005
R209 source.n27 source.n26 9.3005
R210 source.n41 source.n40 9.3005
R211 source.n88 source.n7 8.93611
R212 source.n86 source.n80 8.14595
R213 source.n72 source.n66 8.14595
R214 source.n64 source.n58 8.14595
R215 source.n50 source.n44 8.14595
R216 source.n6 source.n0 8.14595
R217 source.n20 source.n14 8.14595
R218 source.n28 source.n22 8.14595
R219 source.n42 source.n36 8.14595
R220 source.n84 source.n83 7.3702
R221 source.n70 source.n69 7.3702
R222 source.n62 source.n61 7.3702
R223 source.n48 source.n47 7.3702
R224 source.n4 source.n3 7.3702
R225 source.n18 source.n17 7.3702
R226 source.n26 source.n25 7.3702
R227 source.n40 source.n39 7.3702
R228 source.n84 source.n80 5.81868
R229 source.n70 source.n66 5.81868
R230 source.n62 source.n58 5.81868
R231 source.n48 source.n44 5.81868
R232 source.n4 source.n0 5.81868
R233 source.n18 source.n14 5.81868
R234 source.n26 source.n22 5.81868
R235 source.n40 source.n36 5.81868
R236 source.n88 source.n87 5.7505
R237 source.n85 source.n81 3.44771
R238 source.n71 source.n67 3.44771
R239 source.n63 source.n59 3.44771
R240 source.n49 source.n45 3.44771
R241 source.n5 source.n1 3.44771
R242 source.n19 source.n15 3.44771
R243 source.n27 source.n23 3.44771
R244 source.n41 source.n37 3.44771
R245 source.n43 source.n35 0.974638
R246 source.n35 source.n33 0.974638
R247 source.n33 source.n31 0.974638
R248 source.n31 source.n29 0.974638
R249 source.n21 source.n13 0.974638
R250 source.n13 source.n11 0.974638
R251 source.n11 source.n9 0.974638
R252 source.n9 source.n7 0.974638
R253 source.n53 source.n51 0.974638
R254 source.n55 source.n53 0.974638
R255 source.n57 source.n55 0.974638
R256 source.n65 source.n57 0.974638
R257 source.n75 source.n73 0.974638
R258 source.n77 source.n75 0.974638
R259 source.n79 source.n77 0.974638
R260 source.n87 source.n79 0.974638
R261 source.n29 source.n21 0.470328
R262 source.n73 source.n65 0.470328
R263 source source.n88 0.188
R264 minus.n21 minus.n20 161.3
R265 minus.n19 minus.n0 161.3
R266 minus.n15 minus.n14 161.3
R267 minus.n13 minus.n2 161.3
R268 minus.n12 minus.n11 161.3
R269 minus.n10 minus.n3 161.3
R270 minus.n9 minus.n8 161.3
R271 minus.n43 minus.n42 161.3
R272 minus.n41 minus.n22 161.3
R273 minus.n37 minus.n36 161.3
R274 minus.n35 minus.n24 161.3
R275 minus.n34 minus.n33 161.3
R276 minus.n32 minus.n25 161.3
R277 minus.n31 minus.n30 161.3
R278 minus.n5 minus.t7 130.377
R279 minus.n27 minus.t14 130.377
R280 minus.n6 minus.t5 109.355
R281 minus.n7 minus.t4 109.355
R282 minus.n3 minus.t11 109.355
R283 minus.n13 minus.t12 109.355
R284 minus.n1 minus.t9 109.355
R285 minus.n18 minus.t6 109.355
R286 minus.n20 minus.t13 109.355
R287 minus.n28 minus.t0 109.355
R288 minus.n29 minus.t15 109.355
R289 minus.n25 minus.t1 109.355
R290 minus.n35 minus.t8 109.355
R291 minus.n23 minus.t2 109.355
R292 minus.n40 minus.t10 109.355
R293 minus.n42 minus.t3 109.355
R294 minus.n18 minus.n17 80.6037
R295 minus.n16 minus.n1 80.6037
R296 minus.n7 minus.n4 80.6037
R297 minus.n40 minus.n39 80.6037
R298 minus.n38 minus.n23 80.6037
R299 minus.n29 minus.n26 80.6037
R300 minus.n7 minus.n6 48.2005
R301 minus.n18 minus.n1 48.2005
R302 minus.n29 minus.n28 48.2005
R303 minus.n40 minus.n23 48.2005
R304 minus.n8 minus.n7 43.0884
R305 minus.n14 minus.n1 43.0884
R306 minus.n30 minus.n29 43.0884
R307 minus.n36 minus.n23 43.0884
R308 minus.n19 minus.n18 40.1672
R309 minus.n41 minus.n40 40.1672
R310 minus.n44 minus.n21 32.1179
R311 minus.n5 minus.n4 31.6481
R312 minus.n27 minus.n26 31.6481
R313 minus.n13 minus.n12 24.1005
R314 minus.n12 minus.n3 24.1005
R315 minus.n34 minus.n25 24.1005
R316 minus.n35 minus.n34 24.1005
R317 minus.n6 minus.n5 17.444
R318 minus.n28 minus.n27 17.444
R319 minus.n20 minus.n19 8.03383
R320 minus.n42 minus.n41 8.03383
R321 minus.n44 minus.n43 6.6558
R322 minus.n8 minus.n3 5.11262
R323 minus.n14 minus.n13 5.11262
R324 minus.n30 minus.n25 5.11262
R325 minus.n36 minus.n35 5.11262
R326 minus.n17 minus.n16 0.380177
R327 minus.n39 minus.n38 0.380177
R328 minus.n17 minus.n0 0.285035
R329 minus.n16 minus.n15 0.285035
R330 minus.n9 minus.n4 0.285035
R331 minus.n31 minus.n26 0.285035
R332 minus.n38 minus.n37 0.285035
R333 minus.n39 minus.n22 0.285035
R334 minus.n21 minus.n0 0.189894
R335 minus.n15 minus.n2 0.189894
R336 minus.n11 minus.n2 0.189894
R337 minus.n11 minus.n10 0.189894
R338 minus.n10 minus.n9 0.189894
R339 minus.n32 minus.n31 0.189894
R340 minus.n33 minus.n32 0.189894
R341 minus.n33 minus.n24 0.189894
R342 minus.n37 minus.n24 0.189894
R343 minus.n43 minus.n22 0.189894
R344 minus minus.n44 0.188
R345 drain_right.n9 drain_right.n7 101.769
R346 drain_right.n5 drain_right.n3 101.769
R347 drain_right.n2 drain_right.n0 101.769
R348 drain_right.n9 drain_right.n8 100.796
R349 drain_right.n11 drain_right.n10 100.796
R350 drain_right.n13 drain_right.n12 100.796
R351 drain_right.n5 drain_right.n4 100.796
R352 drain_right.n2 drain_right.n1 100.796
R353 drain_right drain_right.n6 25.57
R354 drain_right.n3 drain_right.t5 9.9005
R355 drain_right.n3 drain_right.t12 9.9005
R356 drain_right.n4 drain_right.t7 9.9005
R357 drain_right.n4 drain_right.t13 9.9005
R358 drain_right.n1 drain_right.t0 9.9005
R359 drain_right.n1 drain_right.t14 9.9005
R360 drain_right.n0 drain_right.t1 9.9005
R361 drain_right.n0 drain_right.t15 9.9005
R362 drain_right.n7 drain_right.t10 9.9005
R363 drain_right.n7 drain_right.t8 9.9005
R364 drain_right.n8 drain_right.t4 9.9005
R365 drain_right.n8 drain_right.t11 9.9005
R366 drain_right.n10 drain_right.t6 9.9005
R367 drain_right.n10 drain_right.t3 9.9005
R368 drain_right.n12 drain_right.t2 9.9005
R369 drain_right.n12 drain_right.t9 9.9005
R370 drain_right drain_right.n13 6.62735
R371 drain_right.n13 drain_right.n11 0.974638
R372 drain_right.n11 drain_right.n9 0.974638
R373 drain_right.n6 drain_right.n5 0.432223
R374 drain_right.n6 drain_right.n2 0.432223
C0 minus drain_left 0.179408f
C1 plus source 3.01388f
C2 source drain_right 6.12752f
C3 plus drain_right 0.437249f
C4 drain_left source 6.12476f
C5 plus drain_left 2.60295f
C6 drain_left drain_right 1.44945f
C7 minus source 2.99992f
C8 plus minus 4.73206f
C9 minus drain_right 2.32972f
C10 drain_right a_n2750_n1288# 4.99156f
C11 drain_left a_n2750_n1288# 5.40373f
C12 source a_n2750_n1288# 3.4367f
C13 minus a_n2750_n1288# 10.180932f
C14 plus a_n2750_n1288# 11.46417f
C15 drain_right.t1 a_n2750_n1288# 0.041005f
C16 drain_right.t15 a_n2750_n1288# 0.041005f
C17 drain_right.n0 a_n2750_n1288# 0.261163f
C18 drain_right.t0 a_n2750_n1288# 0.041005f
C19 drain_right.t14 a_n2750_n1288# 0.041005f
C20 drain_right.n1 a_n2750_n1288# 0.257603f
C21 drain_right.n2 a_n2750_n1288# 0.685843f
C22 drain_right.t5 a_n2750_n1288# 0.041005f
C23 drain_right.t12 a_n2750_n1288# 0.041005f
C24 drain_right.n3 a_n2750_n1288# 0.261163f
C25 drain_right.t7 a_n2750_n1288# 0.041005f
C26 drain_right.t13 a_n2750_n1288# 0.041005f
C27 drain_right.n4 a_n2750_n1288# 0.257603f
C28 drain_right.n5 a_n2750_n1288# 0.685843f
C29 drain_right.n6 a_n2750_n1288# 0.952138f
C30 drain_right.t10 a_n2750_n1288# 0.041005f
C31 drain_right.t8 a_n2750_n1288# 0.041005f
C32 drain_right.n7 a_n2750_n1288# 0.261164f
C33 drain_right.t4 a_n2750_n1288# 0.041005f
C34 drain_right.t11 a_n2750_n1288# 0.041005f
C35 drain_right.n8 a_n2750_n1288# 0.257604f
C36 drain_right.n9 a_n2750_n1288# 0.729793f
C37 drain_right.t6 a_n2750_n1288# 0.041005f
C38 drain_right.t3 a_n2750_n1288# 0.041005f
C39 drain_right.n10 a_n2750_n1288# 0.257604f
C40 drain_right.n11 a_n2750_n1288# 0.361452f
C41 drain_right.t2 a_n2750_n1288# 0.041005f
C42 drain_right.t9 a_n2750_n1288# 0.041005f
C43 drain_right.n12 a_n2750_n1288# 0.257604f
C44 drain_right.n13 a_n2750_n1288# 0.594096f
C45 minus.n0 a_n2750_n1288# 0.055133f
C46 minus.t9 a_n2750_n1288# 0.204717f
C47 minus.n1 a_n2750_n1288# 0.150324f
C48 minus.t6 a_n2750_n1288# 0.204717f
C49 minus.n2 a_n2750_n1288# 0.041317f
C50 minus.t11 a_n2750_n1288# 0.204717f
C51 minus.n3 a_n2750_n1288# 0.138528f
C52 minus.n4 a_n2750_n1288# 0.236975f
C53 minus.t7 a_n2750_n1288# 0.227637f
C54 minus.n5 a_n2750_n1288# 0.12292f
C55 minus.t5 a_n2750_n1288# 0.204717f
C56 minus.n6 a_n2750_n1288# 0.150648f
C57 minus.t4 a_n2750_n1288# 0.204717f
C58 minus.n7 a_n2750_n1288# 0.150324f
C59 minus.n8 a_n2750_n1288# 0.009376f
C60 minus.n9 a_n2750_n1288# 0.055133f
C61 minus.n10 a_n2750_n1288# 0.041317f
C62 minus.n11 a_n2750_n1288# 0.041317f
C63 minus.n12 a_n2750_n1288# 0.009376f
C64 minus.t12 a_n2750_n1288# 0.204717f
C65 minus.n13 a_n2750_n1288# 0.138528f
C66 minus.n14 a_n2750_n1288# 0.009376f
C67 minus.n15 a_n2750_n1288# 0.055133f
C68 minus.n16 a_n2750_n1288# 0.068819f
C69 minus.n17 a_n2750_n1288# 0.068819f
C70 minus.n18 a_n2750_n1288# 0.149814f
C71 minus.n19 a_n2750_n1288# 0.009376f
C72 minus.t13 a_n2750_n1288# 0.204717f
C73 minus.n20 a_n2750_n1288# 0.134834f
C74 minus.n21 a_n2750_n1288# 1.21085f
C75 minus.n22 a_n2750_n1288# 0.055133f
C76 minus.t2 a_n2750_n1288# 0.204717f
C77 minus.n23 a_n2750_n1288# 0.150324f
C78 minus.n24 a_n2750_n1288# 0.041317f
C79 minus.t1 a_n2750_n1288# 0.204717f
C80 minus.n25 a_n2750_n1288# 0.138528f
C81 minus.n26 a_n2750_n1288# 0.236975f
C82 minus.t14 a_n2750_n1288# 0.227637f
C83 minus.n27 a_n2750_n1288# 0.12292f
C84 minus.t0 a_n2750_n1288# 0.204717f
C85 minus.n28 a_n2750_n1288# 0.150648f
C86 minus.t15 a_n2750_n1288# 0.204717f
C87 minus.n29 a_n2750_n1288# 0.150324f
C88 minus.n30 a_n2750_n1288# 0.009376f
C89 minus.n31 a_n2750_n1288# 0.055133f
C90 minus.n32 a_n2750_n1288# 0.041317f
C91 minus.n33 a_n2750_n1288# 0.041317f
C92 minus.n34 a_n2750_n1288# 0.009376f
C93 minus.t8 a_n2750_n1288# 0.204717f
C94 minus.n35 a_n2750_n1288# 0.138528f
C95 minus.n36 a_n2750_n1288# 0.009376f
C96 minus.n37 a_n2750_n1288# 0.055133f
C97 minus.n38 a_n2750_n1288# 0.068819f
C98 minus.n39 a_n2750_n1288# 0.068819f
C99 minus.t10 a_n2750_n1288# 0.204717f
C100 minus.n40 a_n2750_n1288# 0.149814f
C101 minus.n41 a_n2750_n1288# 0.009376f
C102 minus.t3 a_n2750_n1288# 0.204717f
C103 minus.n42 a_n2750_n1288# 0.134834f
C104 minus.n43 a_n2750_n1288# 0.285177f
C105 minus.n44 a_n2750_n1288# 1.48076f
C106 source.n0 a_n2750_n1288# 0.044367f
C107 source.n1 a_n2750_n1288# 0.098168f
C108 source.t12 a_n2750_n1288# 0.07367f
C109 source.n2 a_n2750_n1288# 0.07683f
C110 source.n3 a_n2750_n1288# 0.024767f
C111 source.n4 a_n2750_n1288# 0.016334f
C112 source.n5 a_n2750_n1288# 0.216387f
C113 source.n6 a_n2750_n1288# 0.048637f
C114 source.n7 a_n2750_n1288# 0.533702f
C115 source.t9 a_n2750_n1288# 0.048042f
C116 source.t10 a_n2750_n1288# 0.048042f
C117 source.n8 a_n2750_n1288# 0.256833f
C118 source.n9 a_n2750_n1288# 0.427158f
C119 source.t8 a_n2750_n1288# 0.048042f
C120 source.t6 a_n2750_n1288# 0.048042f
C121 source.n10 a_n2750_n1288# 0.256833f
C122 source.n11 a_n2750_n1288# 0.427158f
C123 source.t5 a_n2750_n1288# 0.048042f
C124 source.t7 a_n2750_n1288# 0.048042f
C125 source.n12 a_n2750_n1288# 0.256833f
C126 source.n13 a_n2750_n1288# 0.427158f
C127 source.n14 a_n2750_n1288# 0.044367f
C128 source.n15 a_n2750_n1288# 0.098168f
C129 source.t3 a_n2750_n1288# 0.07367f
C130 source.n16 a_n2750_n1288# 0.07683f
C131 source.n17 a_n2750_n1288# 0.024767f
C132 source.n18 a_n2750_n1288# 0.016334f
C133 source.n19 a_n2750_n1288# 0.216387f
C134 source.n20 a_n2750_n1288# 0.048637f
C135 source.n21 a_n2750_n1288# 0.166458f
C136 source.n22 a_n2750_n1288# 0.044367f
C137 source.n23 a_n2750_n1288# 0.098168f
C138 source.t25 a_n2750_n1288# 0.07367f
C139 source.n24 a_n2750_n1288# 0.07683f
C140 source.n25 a_n2750_n1288# 0.024767f
C141 source.n26 a_n2750_n1288# 0.016334f
C142 source.n27 a_n2750_n1288# 0.216387f
C143 source.n28 a_n2750_n1288# 0.048637f
C144 source.n29 a_n2750_n1288# 0.166458f
C145 source.t0 a_n2750_n1288# 0.048042f
C146 source.t30 a_n2750_n1288# 0.048042f
C147 source.n30 a_n2750_n1288# 0.256833f
C148 source.n31 a_n2750_n1288# 0.427158f
C149 source.t24 a_n2750_n1288# 0.048042f
C150 source.t29 a_n2750_n1288# 0.048042f
C151 source.n32 a_n2750_n1288# 0.256833f
C152 source.n33 a_n2750_n1288# 0.427158f
C153 source.t28 a_n2750_n1288# 0.048042f
C154 source.t27 a_n2750_n1288# 0.048042f
C155 source.n34 a_n2750_n1288# 0.256833f
C156 source.n35 a_n2750_n1288# 0.427158f
C157 source.n36 a_n2750_n1288# 0.044367f
C158 source.n37 a_n2750_n1288# 0.098168f
C159 source.t22 a_n2750_n1288# 0.07367f
C160 source.n38 a_n2750_n1288# 0.07683f
C161 source.n39 a_n2750_n1288# 0.024767f
C162 source.n40 a_n2750_n1288# 0.016334f
C163 source.n41 a_n2750_n1288# 0.216387f
C164 source.n42 a_n2750_n1288# 0.048637f
C165 source.n43 a_n2750_n1288# 0.826793f
C166 source.n44 a_n2750_n1288# 0.044367f
C167 source.n45 a_n2750_n1288# 0.098168f
C168 source.t17 a_n2750_n1288# 0.07367f
C169 source.n46 a_n2750_n1288# 0.07683f
C170 source.n47 a_n2750_n1288# 0.024767f
C171 source.n48 a_n2750_n1288# 0.016334f
C172 source.n49 a_n2750_n1288# 0.216387f
C173 source.n50 a_n2750_n1288# 0.048637f
C174 source.n51 a_n2750_n1288# 0.826793f
C175 source.t11 a_n2750_n1288# 0.048042f
C176 source.t14 a_n2750_n1288# 0.048042f
C177 source.n52 a_n2750_n1288# 0.256832f
C178 source.n53 a_n2750_n1288# 0.42716f
C179 source.t13 a_n2750_n1288# 0.048042f
C180 source.t15 a_n2750_n1288# 0.048042f
C181 source.n54 a_n2750_n1288# 0.256832f
C182 source.n55 a_n2750_n1288# 0.42716f
C183 source.t2 a_n2750_n1288# 0.048042f
C184 source.t16 a_n2750_n1288# 0.048042f
C185 source.n56 a_n2750_n1288# 0.256832f
C186 source.n57 a_n2750_n1288# 0.42716f
C187 source.n58 a_n2750_n1288# 0.044367f
C188 source.n59 a_n2750_n1288# 0.098168f
C189 source.t4 a_n2750_n1288# 0.07367f
C190 source.n60 a_n2750_n1288# 0.07683f
C191 source.n61 a_n2750_n1288# 0.024767f
C192 source.n62 a_n2750_n1288# 0.016334f
C193 source.n63 a_n2750_n1288# 0.216387f
C194 source.n64 a_n2750_n1288# 0.048637f
C195 source.n65 a_n2750_n1288# 0.166458f
C196 source.n66 a_n2750_n1288# 0.044367f
C197 source.n67 a_n2750_n1288# 0.098168f
C198 source.t21 a_n2750_n1288# 0.07367f
C199 source.n68 a_n2750_n1288# 0.07683f
C200 source.n69 a_n2750_n1288# 0.024767f
C201 source.n70 a_n2750_n1288# 0.016334f
C202 source.n71 a_n2750_n1288# 0.216387f
C203 source.n72 a_n2750_n1288# 0.048637f
C204 source.n73 a_n2750_n1288# 0.166458f
C205 source.t19 a_n2750_n1288# 0.048042f
C206 source.t23 a_n2750_n1288# 0.048042f
C207 source.n74 a_n2750_n1288# 0.256832f
C208 source.n75 a_n2750_n1288# 0.42716f
C209 source.t1 a_n2750_n1288# 0.048042f
C210 source.t26 a_n2750_n1288# 0.048042f
C211 source.n76 a_n2750_n1288# 0.256832f
C212 source.n77 a_n2750_n1288# 0.42716f
C213 source.t20 a_n2750_n1288# 0.048042f
C214 source.t31 a_n2750_n1288# 0.048042f
C215 source.n78 a_n2750_n1288# 0.256832f
C216 source.n79 a_n2750_n1288# 0.42716f
C217 source.n80 a_n2750_n1288# 0.044367f
C218 source.n81 a_n2750_n1288# 0.098168f
C219 source.t18 a_n2750_n1288# 0.07367f
C220 source.n82 a_n2750_n1288# 0.07683f
C221 source.n83 a_n2750_n1288# 0.024767f
C222 source.n84 a_n2750_n1288# 0.016334f
C223 source.n85 a_n2750_n1288# 0.216387f
C224 source.n86 a_n2750_n1288# 0.048637f
C225 source.n87 a_n2750_n1288# 0.371324f
C226 source.n88 a_n2750_n1288# 0.77018f
C227 drain_left.t10 a_n2750_n1288# 0.041962f
C228 drain_left.t12 a_n2750_n1288# 0.041962f
C229 drain_left.n0 a_n2750_n1288# 0.267261f
C230 drain_left.t5 a_n2750_n1288# 0.041962f
C231 drain_left.t15 a_n2750_n1288# 0.041962f
C232 drain_left.n1 a_n2750_n1288# 0.263618f
C233 drain_left.n2 a_n2750_n1288# 0.701858f
C234 drain_left.t11 a_n2750_n1288# 0.041962f
C235 drain_left.t7 a_n2750_n1288# 0.041962f
C236 drain_left.n3 a_n2750_n1288# 0.267261f
C237 drain_left.t1 a_n2750_n1288# 0.041962f
C238 drain_left.t14 a_n2750_n1288# 0.041962f
C239 drain_left.n4 a_n2750_n1288# 0.263618f
C240 drain_left.n5 a_n2750_n1288# 0.701858f
C241 drain_left.n6 a_n2750_n1288# 1.02594f
C242 drain_left.t0 a_n2750_n1288# 0.041962f
C243 drain_left.t9 a_n2750_n1288# 0.041962f
C244 drain_left.n7 a_n2750_n1288# 0.267262f
C245 drain_left.t13 a_n2750_n1288# 0.041962f
C246 drain_left.t6 a_n2750_n1288# 0.041962f
C247 drain_left.n8 a_n2750_n1288# 0.263619f
C248 drain_left.n9 a_n2750_n1288# 0.746834f
C249 drain_left.t4 a_n2750_n1288# 0.041962f
C250 drain_left.t3 a_n2750_n1288# 0.041962f
C251 drain_left.n10 a_n2750_n1288# 0.263619f
C252 drain_left.n11 a_n2750_n1288# 0.369891f
C253 drain_left.t8 a_n2750_n1288# 0.041962f
C254 drain_left.t2 a_n2750_n1288# 0.041962f
C255 drain_left.n12 a_n2750_n1288# 0.263619f
C256 drain_left.n13 a_n2750_n1288# 0.607968f
C257 plus.n0 a_n2750_n1288# 0.057265f
C258 plus.t5 a_n2750_n1288# 0.212635f
C259 plus.t7 a_n2750_n1288# 0.212635f
C260 plus.n1 a_n2750_n1288# 0.071481f
C261 plus.t8 a_n2750_n1288# 0.212635f
C262 plus.n2 a_n2750_n1288# 0.071481f
C263 plus.t11 a_n2750_n1288# 0.212635f
C264 plus.n3 a_n2750_n1288# 0.143886f
C265 plus.n4 a_n2750_n1288# 0.042915f
C266 plus.t9 a_n2750_n1288# 0.212635f
C267 plus.t10 a_n2750_n1288# 0.212635f
C268 plus.n5 a_n2750_n1288# 0.156138f
C269 plus.t12 a_n2750_n1288# 0.212635f
C270 plus.n6 a_n2750_n1288# 0.156474f
C271 plus.t14 a_n2750_n1288# 0.236441f
C272 plus.n7 a_n2750_n1288# 0.127675f
C273 plus.n8 a_n2750_n1288# 0.24614f
C274 plus.n9 a_n2750_n1288# 0.057265f
C275 plus.n10 a_n2750_n1288# 0.009738f
C276 plus.n11 a_n2750_n1288# 0.143886f
C277 plus.n12 a_n2750_n1288# 0.009738f
C278 plus.n13 a_n2750_n1288# 0.042915f
C279 plus.n14 a_n2750_n1288# 0.042915f
C280 plus.n15 a_n2750_n1288# 0.057265f
C281 plus.n16 a_n2750_n1288# 0.009738f
C282 plus.n17 a_n2750_n1288# 0.156138f
C283 plus.n18 a_n2750_n1288# 0.155609f
C284 plus.n19 a_n2750_n1288# 0.009738f
C285 plus.n20 a_n2750_n1288# 0.14005f
C286 plus.n21 a_n2750_n1288# 0.323292f
C287 plus.n22 a_n2750_n1288# 0.057265f
C288 plus.t0 a_n2750_n1288# 0.212635f
C289 plus.n23 a_n2750_n1288# 0.071481f
C290 plus.t6 a_n2750_n1288# 0.212635f
C291 plus.n24 a_n2750_n1288# 0.071481f
C292 plus.t3 a_n2750_n1288# 0.212635f
C293 plus.t4 a_n2750_n1288# 0.212635f
C294 plus.n25 a_n2750_n1288# 0.143886f
C295 plus.n26 a_n2750_n1288# 0.042915f
C296 plus.t2 a_n2750_n1288# 0.212635f
C297 plus.t15 a_n2750_n1288# 0.212635f
C298 plus.n27 a_n2750_n1288# 0.156138f
C299 plus.t1 a_n2750_n1288# 0.212635f
C300 plus.n28 a_n2750_n1288# 0.156474f
C301 plus.t13 a_n2750_n1288# 0.236441f
C302 plus.n29 a_n2750_n1288# 0.127675f
C303 plus.n30 a_n2750_n1288# 0.24614f
C304 plus.n31 a_n2750_n1288# 0.057265f
C305 plus.n32 a_n2750_n1288# 0.009738f
C306 plus.n33 a_n2750_n1288# 0.143886f
C307 plus.n34 a_n2750_n1288# 0.009738f
C308 plus.n35 a_n2750_n1288# 0.042915f
C309 plus.n36 a_n2750_n1288# 0.042915f
C310 plus.n37 a_n2750_n1288# 0.057265f
C311 plus.n38 a_n2750_n1288# 0.009738f
C312 plus.n39 a_n2750_n1288# 0.156138f
C313 plus.n40 a_n2750_n1288# 0.155609f
C314 plus.n41 a_n2750_n1288# 0.009738f
C315 plus.n42 a_n2750_n1288# 0.14005f
C316 plus.n43 a_n2750_n1288# 1.19605f
.ends

