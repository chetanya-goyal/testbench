* NGSPICE file created from diffpair366.ext - technology: sky130A

.subckt diffpair366 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t24 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X1 a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X2 drain_right.t12 minus.t1 source.t25 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 drain_left.t13 plus.t0 source.t11 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X5 drain_left.t12 plus.t1 source.t4 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 source.t21 minus.t2 drain_right.t11 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X7 drain_left.t11 plus.t2 source.t9 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X8 drain_right.t10 minus.t3 source.t20 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 source.t0 plus.t3 drain_left.t10 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 source.t27 minus.t4 drain_right.t9 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 drain_right.t8 minus.t5 source.t26 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 drain_right.t7 minus.t6 source.t19 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 source.t12 plus.t4 drain_left.t9 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 drain_right.t6 minus.t7 source.t18 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X15 a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X16 source.t23 minus.t8 drain_right.t5 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 drain_left.t8 plus.t5 source.t1 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X18 source.t16 minus.t9 drain_right.t4 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 drain_right.t3 minus.t10 source.t14 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X20 source.t5 plus.t6 drain_left.t7 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X21 drain_left.t6 plus.t7 source.t8 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X22 source.t3 plus.t8 drain_left.t5 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X24 source.t17 minus.t11 drain_right.t2 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 drain_left.t4 plus.t9 source.t6 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 source.t13 plus.t10 drain_left.t3 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X27 drain_left.t2 plus.t11 source.t2 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X28 drain_left.t1 plus.t12 source.t7 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 source.t15 minus.t12 drain_right.t1 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X30 drain_right.t0 minus.t13 source.t22 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X31 source.t10 plus.t13 drain_left.t0 a_n2044_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n4 minus.t10 533.348
R1 minus.n20 minus.t13 533.348
R2 minus.n3 minus.t2 512.366
R3 minus.n7 minus.t5 512.366
R4 minus.n8 minus.t11 512.366
R5 minus.n1 minus.t3 512.366
R6 minus.n13 minus.t9 512.366
R7 minus.n14 minus.t0 512.366
R8 minus.n19 minus.t12 512.366
R9 minus.n23 minus.t6 512.366
R10 minus.n24 minus.t4 512.366
R11 minus.n17 minus.t1 512.366
R12 minus.n29 minus.t8 512.366
R13 minus.n30 minus.t7 512.366
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n0 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n1 161.3
R18 minus.n7 minus.n2 161.3
R19 minus.n6 minus.n5 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n16 161.3
R22 minus.n28 minus.n27 161.3
R23 minus.n26 minus.n17 161.3
R24 minus.n23 minus.n18 161.3
R25 minus.n22 minus.n21 161.3
R26 minus.n9 minus.n8 80.6037
R27 minus.n25 minus.n24 80.6037
R28 minus.n5 minus.n4 70.4033
R29 minus.n21 minus.n20 70.4033
R30 minus.n8 minus.n7 48.2005
R31 minus.n8 minus.n1 48.2005
R32 minus.n14 minus.n13 48.2005
R33 minus.n24 minus.n23 48.2005
R34 minus.n24 minus.n17 48.2005
R35 minus.n30 minus.n29 48.2005
R36 minus.n32 minus.n15 34.6842
R37 minus.n7 minus.n6 24.8308
R38 minus.n12 minus.n1 24.8308
R39 minus.n23 minus.n22 24.8308
R40 minus.n28 minus.n17 24.8308
R41 minus.n6 minus.n3 23.3702
R42 minus.n13 minus.n12 23.3702
R43 minus.n22 minus.n19 23.3702
R44 minus.n29 minus.n28 23.3702
R45 minus.n4 minus.n3 20.9576
R46 minus.n20 minus.n19 20.9576
R47 minus.n32 minus.n31 6.5933
R48 minus.n10 minus.n9 0.285035
R49 minus.n9 minus.n2 0.285035
R50 minus.n25 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n5 minus.n2 0.189894
R56 minus.n21 minus.n18 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n16 0.189894
R59 minus.n31 minus.n16 0.189894
R60 minus minus.n32 0.188
R61 source.n7 source.t14 51.0588
R62 source.n27 source.t18 51.0586
R63 source.n20 source.t8 51.0586
R64 source.n0 source.t1 51.0586
R65 source.n2 source.n1 48.8588
R66 source.n4 source.n3 48.8588
R67 source.n6 source.n5 48.8588
R68 source.n9 source.n8 48.8588
R69 source.n11 source.n10 48.8588
R70 source.n13 source.n12 48.8588
R71 source.n26 source.n25 48.8586
R72 source.n24 source.n23 48.8586
R73 source.n22 source.n21 48.8586
R74 source.n19 source.n18 48.8586
R75 source.n17 source.n16 48.8586
R76 source.n15 source.n14 48.8586
R77 source.n15 source.n13 20.446
R78 source.n28 source.n0 14.1098
R79 source.n28 source.n27 5.62119
R80 source.n25 source.t25 2.2005
R81 source.n25 source.t23 2.2005
R82 source.n23 source.t19 2.2005
R83 source.n23 source.t27 2.2005
R84 source.n21 source.t22 2.2005
R85 source.n21 source.t15 2.2005
R86 source.n18 source.t4 2.2005
R87 source.n18 source.t3 2.2005
R88 source.n16 source.t2 2.2005
R89 source.n16 source.t13 2.2005
R90 source.n14 source.t11 2.2005
R91 source.n14 source.t0 2.2005
R92 source.n1 source.t6 2.2005
R93 source.n1 source.t10 2.2005
R94 source.n3 source.t7 2.2005
R95 source.n3 source.t12 2.2005
R96 source.n5 source.t9 2.2005
R97 source.n5 source.t5 2.2005
R98 source.n8 source.t26 2.2005
R99 source.n8 source.t21 2.2005
R100 source.n10 source.t20 2.2005
R101 source.n10 source.t17 2.2005
R102 source.n12 source.t24 2.2005
R103 source.n12 source.t16 2.2005
R104 source.n7 source.n6 0.828086
R105 source.n22 source.n20 0.828086
R106 source.n13 source.n11 0.716017
R107 source.n11 source.n9 0.716017
R108 source.n9 source.n7 0.716017
R109 source.n6 source.n4 0.716017
R110 source.n4 source.n2 0.716017
R111 source.n2 source.n0 0.716017
R112 source.n17 source.n15 0.716017
R113 source.n19 source.n17 0.716017
R114 source.n20 source.n19 0.716017
R115 source.n24 source.n22 0.716017
R116 source.n26 source.n24 0.716017
R117 source.n27 source.n26 0.716017
R118 source source.n28 0.188
R119 drain_right.n1 drain_right.t0 68.4529
R120 drain_right.n11 drain_right.t13 67.7376
R121 drain_right.n8 drain_right.n6 66.2529
R122 drain_right.n4 drain_right.n2 66.2529
R123 drain_right.n8 drain_right.n7 65.5376
R124 drain_right.n10 drain_right.n9 65.5376
R125 drain_right.n4 drain_right.n3 65.5373
R126 drain_right.n1 drain_right.n0 65.5373
R127 drain_right drain_right.n5 28.6553
R128 drain_right drain_right.n11 6.01097
R129 drain_right.n2 drain_right.t5 2.2005
R130 drain_right.n2 drain_right.t6 2.2005
R131 drain_right.n3 drain_right.t9 2.2005
R132 drain_right.n3 drain_right.t12 2.2005
R133 drain_right.n0 drain_right.t1 2.2005
R134 drain_right.n0 drain_right.t7 2.2005
R135 drain_right.n6 drain_right.t11 2.2005
R136 drain_right.n6 drain_right.t3 2.2005
R137 drain_right.n7 drain_right.t2 2.2005
R138 drain_right.n7 drain_right.t8 2.2005
R139 drain_right.n9 drain_right.t4 2.2005
R140 drain_right.n9 drain_right.t10 2.2005
R141 drain_right.n11 drain_right.n10 0.716017
R142 drain_right.n10 drain_right.n8 0.716017
R143 drain_right.n5 drain_right.n1 0.481792
R144 drain_right.n5 drain_right.n4 0.124033
R145 plus.n4 plus.t2 533.348
R146 plus.n20 plus.t7 533.348
R147 plus.n14 plus.t5 512.366
R148 plus.n13 plus.t13 512.366
R149 plus.n1 plus.t9 512.366
R150 plus.n8 plus.t4 512.366
R151 plus.n7 plus.t12 512.366
R152 plus.n3 plus.t6 512.366
R153 plus.n30 plus.t0 512.366
R154 plus.n29 plus.t3 512.366
R155 plus.n17 plus.t11 512.366
R156 plus.n24 plus.t10 512.366
R157 plus.n23 plus.t1 512.366
R158 plus.n19 plus.t8 512.366
R159 plus.n6 plus.n5 161.3
R160 plus.n7 plus.n2 161.3
R161 plus.n10 plus.n1 161.3
R162 plus.n12 plus.n11 161.3
R163 plus.n13 plus.n0 161.3
R164 plus.n15 plus.n14 161.3
R165 plus.n22 plus.n21 161.3
R166 plus.n23 plus.n18 161.3
R167 plus.n26 plus.n17 161.3
R168 plus.n28 plus.n27 161.3
R169 plus.n29 plus.n16 161.3
R170 plus.n31 plus.n30 161.3
R171 plus.n9 plus.n8 80.6037
R172 plus.n25 plus.n24 80.6037
R173 plus.n5 plus.n4 70.4033
R174 plus.n21 plus.n20 70.4033
R175 plus.n14 plus.n13 48.2005
R176 plus.n8 plus.n1 48.2005
R177 plus.n8 plus.n7 48.2005
R178 plus.n30 plus.n29 48.2005
R179 plus.n24 plus.n17 48.2005
R180 plus.n24 plus.n23 48.2005
R181 plus plus.n31 29.7017
R182 plus.n12 plus.n1 24.8308
R183 plus.n7 plus.n6 24.8308
R184 plus.n28 plus.n17 24.8308
R185 plus.n23 plus.n22 24.8308
R186 plus.n13 plus.n12 23.3702
R187 plus.n6 plus.n3 23.3702
R188 plus.n29 plus.n28 23.3702
R189 plus.n22 plus.n19 23.3702
R190 plus.n4 plus.n3 20.9576
R191 plus.n20 plus.n19 20.9576
R192 plus plus.n15 11.1009
R193 plus.n9 plus.n2 0.285035
R194 plus.n10 plus.n9 0.285035
R195 plus.n26 plus.n25 0.285035
R196 plus.n25 plus.n18 0.285035
R197 plus.n5 plus.n2 0.189894
R198 plus.n11 plus.n10 0.189894
R199 plus.n11 plus.n0 0.189894
R200 plus.n15 plus.n0 0.189894
R201 plus.n31 plus.n16 0.189894
R202 plus.n27 plus.n16 0.189894
R203 plus.n27 plus.n26 0.189894
R204 plus.n21 plus.n18 0.189894
R205 drain_left.n7 drain_left.t11 68.4531
R206 drain_left.n1 drain_left.t13 68.4529
R207 drain_left.n4 drain_left.n2 66.2529
R208 drain_left.n9 drain_left.n8 65.5376
R209 drain_left.n7 drain_left.n6 65.5376
R210 drain_left.n11 drain_left.n10 65.5374
R211 drain_left.n4 drain_left.n3 65.5373
R212 drain_left.n1 drain_left.n0 65.5373
R213 drain_left drain_left.n5 29.2086
R214 drain_left drain_left.n11 6.36873
R215 drain_left.n2 drain_left.t5 2.2005
R216 drain_left.n2 drain_left.t6 2.2005
R217 drain_left.n3 drain_left.t3 2.2005
R218 drain_left.n3 drain_left.t12 2.2005
R219 drain_left.n0 drain_left.t10 2.2005
R220 drain_left.n0 drain_left.t2 2.2005
R221 drain_left.n10 drain_left.t0 2.2005
R222 drain_left.n10 drain_left.t8 2.2005
R223 drain_left.n8 drain_left.t9 2.2005
R224 drain_left.n8 drain_left.t4 2.2005
R225 drain_left.n6 drain_left.t7 2.2005
R226 drain_left.n6 drain_left.t1 2.2005
R227 drain_left.n9 drain_left.n7 0.716017
R228 drain_left.n11 drain_left.n9 0.716017
R229 drain_left.n5 drain_left.n1 0.481792
R230 drain_left.n5 drain_left.n4 0.124033
C0 drain_right drain_left 1.05823f
C1 drain_right minus 5.69379f
C2 drain_left minus 0.172393f
C3 drain_right source 17.1593f
C4 drain_left source 17.1654f
C5 source minus 5.64252f
C6 drain_right plus 0.356914f
C7 drain_left plus 5.89174f
C8 plus minus 5.14027f
C9 plus source 5.65698f
C10 drain_right a_n2044_n2688# 6.51003f
C11 drain_left a_n2044_n2688# 6.82534f
C12 source a_n2044_n2688# 5.376417f
C13 minus a_n2044_n2688# 7.837464f
C14 plus a_n2044_n2688# 9.51304f
C15 drain_left.t13 a_n2044_n2688# 2.13362f
C16 drain_left.t10 a_n2044_n2688# 0.191304f
C17 drain_left.t2 a_n2044_n2688# 0.191304f
C18 drain_left.n0 a_n2044_n2688# 1.67327f
C19 drain_left.n1 a_n2044_n2688# 0.670179f
C20 drain_left.t5 a_n2044_n2688# 0.191304f
C21 drain_left.t6 a_n2044_n2688# 0.191304f
C22 drain_left.n2 a_n2044_n2688# 1.67705f
C23 drain_left.t3 a_n2044_n2688# 0.191304f
C24 drain_left.t12 a_n2044_n2688# 0.191304f
C25 drain_left.n3 a_n2044_n2688# 1.67327f
C26 drain_left.n4 a_n2044_n2688# 0.639773f
C27 drain_left.n5 a_n2044_n2688# 1.20132f
C28 drain_left.t11 a_n2044_n2688# 2.13363f
C29 drain_left.t7 a_n2044_n2688# 0.191304f
C30 drain_left.t1 a_n2044_n2688# 0.191304f
C31 drain_left.n6 a_n2044_n2688# 1.67327f
C32 drain_left.n7 a_n2044_n2688# 0.689178f
C33 drain_left.t9 a_n2044_n2688# 0.191304f
C34 drain_left.t4 a_n2044_n2688# 0.191304f
C35 drain_left.n8 a_n2044_n2688# 1.67327f
C36 drain_left.n9 a_n2044_n2688# 0.339488f
C37 drain_left.t0 a_n2044_n2688# 0.191304f
C38 drain_left.t8 a_n2044_n2688# 0.191304f
C39 drain_left.n10 a_n2044_n2688# 1.67327f
C40 drain_left.n11 a_n2044_n2688# 0.57059f
C41 plus.n0 a_n2044_n2688# 0.046742f
C42 plus.t5 a_n2044_n2688# 0.603227f
C43 plus.t13 a_n2044_n2688# 0.603227f
C44 plus.t9 a_n2044_n2688# 0.603227f
C45 plus.n1 a_n2044_n2688# 0.261993f
C46 plus.n2 a_n2044_n2688# 0.062372f
C47 plus.t4 a_n2044_n2688# 0.603227f
C48 plus.t12 a_n2044_n2688# 0.603227f
C49 plus.t6 a_n2044_n2688# 0.603227f
C50 plus.n3 a_n2044_n2688# 0.261705f
C51 plus.t2 a_n2044_n2688# 0.613344f
C52 plus.n4 a_n2044_n2688# 0.247337f
C53 plus.n5 a_n2044_n2688# 0.1537f
C54 plus.n6 a_n2044_n2688# 0.010607f
C55 plus.n7 a_n2044_n2688# 0.261993f
C56 plus.n8 a_n2044_n2688# 0.267701f
C57 plus.n9 a_n2044_n2688# 0.062226f
C58 plus.n10 a_n2044_n2688# 0.062372f
C59 plus.n11 a_n2044_n2688# 0.046742f
C60 plus.n12 a_n2044_n2688# 0.010607f
C61 plus.n13 a_n2044_n2688# 0.261705f
C62 plus.n14 a_n2044_n2688# 0.257094f
C63 plus.n15 a_n2044_n2688# 0.469699f
C64 plus.n16 a_n2044_n2688# 0.046742f
C65 plus.t0 a_n2044_n2688# 0.603227f
C66 plus.t3 a_n2044_n2688# 0.603227f
C67 plus.t11 a_n2044_n2688# 0.603227f
C68 plus.n17 a_n2044_n2688# 0.261993f
C69 plus.n18 a_n2044_n2688# 0.062372f
C70 plus.t10 a_n2044_n2688# 0.603227f
C71 plus.t1 a_n2044_n2688# 0.603227f
C72 plus.t8 a_n2044_n2688# 0.603227f
C73 plus.n19 a_n2044_n2688# 0.261705f
C74 plus.t7 a_n2044_n2688# 0.613344f
C75 plus.n20 a_n2044_n2688# 0.247337f
C76 plus.n21 a_n2044_n2688# 0.1537f
C77 plus.n22 a_n2044_n2688# 0.010607f
C78 plus.n23 a_n2044_n2688# 0.261993f
C79 plus.n24 a_n2044_n2688# 0.267701f
C80 plus.n25 a_n2044_n2688# 0.062226f
C81 plus.n26 a_n2044_n2688# 0.062372f
C82 plus.n27 a_n2044_n2688# 0.046742f
C83 plus.n28 a_n2044_n2688# 0.010607f
C84 plus.n29 a_n2044_n2688# 0.261705f
C85 plus.n30 a_n2044_n2688# 0.257094f
C86 plus.n31 a_n2044_n2688# 1.35261f
C87 drain_right.t0 a_n2044_n2688# 2.12483f
C88 drain_right.t1 a_n2044_n2688# 0.190515f
C89 drain_right.t7 a_n2044_n2688# 0.190515f
C90 drain_right.n0 a_n2044_n2688# 1.66637f
C91 drain_right.n1 a_n2044_n2688# 0.667417f
C92 drain_right.t5 a_n2044_n2688# 0.190515f
C93 drain_right.t6 a_n2044_n2688# 0.190515f
C94 drain_right.n2 a_n2044_n2688# 1.67014f
C95 drain_right.t9 a_n2044_n2688# 0.190515f
C96 drain_right.t12 a_n2044_n2688# 0.190515f
C97 drain_right.n3 a_n2044_n2688# 1.66637f
C98 drain_right.n4 a_n2044_n2688# 0.637136f
C99 drain_right.n5 a_n2044_n2688# 1.14142f
C100 drain_right.t11 a_n2044_n2688# 0.190515f
C101 drain_right.t3 a_n2044_n2688# 0.190515f
C102 drain_right.n6 a_n2044_n2688# 1.67014f
C103 drain_right.t2 a_n2044_n2688# 0.190515f
C104 drain_right.t8 a_n2044_n2688# 0.190515f
C105 drain_right.n7 a_n2044_n2688# 1.66638f
C106 drain_right.n8 a_n2044_n2688# 0.683206f
C107 drain_right.t4 a_n2044_n2688# 0.190515f
C108 drain_right.t10 a_n2044_n2688# 0.190515f
C109 drain_right.n9 a_n2044_n2688# 1.66638f
C110 drain_right.n10 a_n2044_n2688# 0.338089f
C111 drain_right.t13 a_n2044_n2688# 2.12115f
C112 drain_right.n11 a_n2044_n2688# 0.586817f
C113 source.t1 a_n2044_n2688# 2.16464f
C114 source.n0 a_n2044_n2688# 1.27125f
C115 source.t6 a_n2044_n2688# 0.202996f
C116 source.t10 a_n2044_n2688# 0.202996f
C117 source.n1 a_n2044_n2688# 1.69935f
C118 source.n2 a_n2044_n2688# 0.397632f
C119 source.t7 a_n2044_n2688# 0.202996f
C120 source.t12 a_n2044_n2688# 0.202996f
C121 source.n3 a_n2044_n2688# 1.69935f
C122 source.n4 a_n2044_n2688# 0.397632f
C123 source.t9 a_n2044_n2688# 0.202996f
C124 source.t5 a_n2044_n2688# 0.202996f
C125 source.n5 a_n2044_n2688# 1.69935f
C126 source.n6 a_n2044_n2688# 0.407939f
C127 source.t14 a_n2044_n2688# 2.16464f
C128 source.n7 a_n2044_n2688# 0.496268f
C129 source.t26 a_n2044_n2688# 0.202996f
C130 source.t21 a_n2044_n2688# 0.202996f
C131 source.n8 a_n2044_n2688# 1.69935f
C132 source.n9 a_n2044_n2688# 0.397632f
C133 source.t20 a_n2044_n2688# 0.202996f
C134 source.t17 a_n2044_n2688# 0.202996f
C135 source.n10 a_n2044_n2688# 1.69935f
C136 source.n11 a_n2044_n2688# 0.397632f
C137 source.t24 a_n2044_n2688# 0.202996f
C138 source.t16 a_n2044_n2688# 0.202996f
C139 source.n12 a_n2044_n2688# 1.69935f
C140 source.n13 a_n2044_n2688# 1.66863f
C141 source.t11 a_n2044_n2688# 0.202996f
C142 source.t0 a_n2044_n2688# 0.202996f
C143 source.n14 a_n2044_n2688# 1.69934f
C144 source.n15 a_n2044_n2688# 1.66864f
C145 source.t2 a_n2044_n2688# 0.202996f
C146 source.t13 a_n2044_n2688# 0.202996f
C147 source.n16 a_n2044_n2688# 1.69934f
C148 source.n17 a_n2044_n2688# 0.397637f
C149 source.t4 a_n2044_n2688# 0.202996f
C150 source.t3 a_n2044_n2688# 0.202996f
C151 source.n18 a_n2044_n2688# 1.69934f
C152 source.n19 a_n2044_n2688# 0.397637f
C153 source.t8 a_n2044_n2688# 2.16464f
C154 source.n20 a_n2044_n2688# 0.496274f
C155 source.t22 a_n2044_n2688# 0.202996f
C156 source.t15 a_n2044_n2688# 0.202996f
C157 source.n21 a_n2044_n2688# 1.69934f
C158 source.n22 a_n2044_n2688# 0.407944f
C159 source.t19 a_n2044_n2688# 0.202996f
C160 source.t27 a_n2044_n2688# 0.202996f
C161 source.n23 a_n2044_n2688# 1.69934f
C162 source.n24 a_n2044_n2688# 0.397637f
C163 source.t25 a_n2044_n2688# 0.202996f
C164 source.t23 a_n2044_n2688# 0.202996f
C165 source.n25 a_n2044_n2688# 1.69934f
C166 source.n26 a_n2044_n2688# 0.397637f
C167 source.t18 a_n2044_n2688# 2.16464f
C168 source.n27 a_n2044_n2688# 0.637094f
C169 source.n28 a_n2044_n2688# 1.49427f
C170 minus.n0 a_n2044_n2688# 0.045644f
C171 minus.t3 a_n2044_n2688# 0.589056f
C172 minus.n1 a_n2044_n2688# 0.255838f
C173 minus.n2 a_n2044_n2688# 0.060907f
C174 minus.t2 a_n2044_n2688# 0.589056f
C175 minus.n3 a_n2044_n2688# 0.255557f
C176 minus.t10 a_n2044_n2688# 0.598936f
C177 minus.n4 a_n2044_n2688# 0.241526f
C178 minus.n5 a_n2044_n2688# 0.15009f
C179 minus.n6 a_n2044_n2688# 0.010358f
C180 minus.t5 a_n2044_n2688# 0.589056f
C181 minus.n7 a_n2044_n2688# 0.255838f
C182 minus.t11 a_n2044_n2688# 0.589056f
C183 minus.n8 a_n2044_n2688# 0.261412f
C184 minus.n9 a_n2044_n2688# 0.060764f
C185 minus.n10 a_n2044_n2688# 0.060907f
C186 minus.n11 a_n2044_n2688# 0.045644f
C187 minus.n12 a_n2044_n2688# 0.010358f
C188 minus.t9 a_n2044_n2688# 0.589056f
C189 minus.n13 a_n2044_n2688# 0.255557f
C190 minus.t0 a_n2044_n2688# 0.589056f
C191 minus.n14 a_n2044_n2688# 0.251054f
C192 minus.n15 a_n2044_n2688# 1.51166f
C193 minus.n16 a_n2044_n2688# 0.045644f
C194 minus.t1 a_n2044_n2688# 0.589056f
C195 minus.n17 a_n2044_n2688# 0.255838f
C196 minus.n18 a_n2044_n2688# 0.060907f
C197 minus.t12 a_n2044_n2688# 0.589056f
C198 minus.n19 a_n2044_n2688# 0.255557f
C199 minus.t13 a_n2044_n2688# 0.598936f
C200 minus.n20 a_n2044_n2688# 0.241526f
C201 minus.n21 a_n2044_n2688# 0.15009f
C202 minus.n22 a_n2044_n2688# 0.010358f
C203 minus.t6 a_n2044_n2688# 0.589056f
C204 minus.n23 a_n2044_n2688# 0.255838f
C205 minus.t4 a_n2044_n2688# 0.589056f
C206 minus.n24 a_n2044_n2688# 0.261412f
C207 minus.n25 a_n2044_n2688# 0.060764f
C208 minus.n26 a_n2044_n2688# 0.060907f
C209 minus.n27 a_n2044_n2688# 0.045644f
C210 minus.n28 a_n2044_n2688# 0.010358f
C211 minus.t8 a_n2044_n2688# 0.589056f
C212 minus.n29 a_n2044_n2688# 0.255557f
C213 minus.t7 a_n2044_n2688# 0.589056f
C214 minus.n30 a_n2044_n2688# 0.251054f
C215 minus.n31 a_n2044_n2688# 0.3084f
C216 minus.n32 a_n2044_n2688# 1.84051f
.ends

