* NGSPICE file created from diffpair261.ext - technology: sky130A

.subckt diffpair261 minus drain_right drain_left source plus
X0 source minus drain_right a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_right minus source a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X2 drain_right minus source a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X3 a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X4 a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X5 drain_left plus source a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X6 source minus drain_right a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X7 a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X8 source plus drain_left a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X9 a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X10 source plus drain_left a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X11 drain_left plus source a_n1064_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
.ends

