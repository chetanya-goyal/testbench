* NGSPICE file created from diffpair503.ext - technology: sky130A

.subckt diffpair503 minus drain_right drain_left source plus
X0 a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X1 drain_left.t7 plus.t0 source.t4 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X2 drain_left.t6 plus.t1 source.t11 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X3 drain_left.t5 plus.t2 source.t8 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X4 source.t1 minus.t0 drain_right.t7 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X5 source.t12 minus.t1 drain_right.t6 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X6 source.t13 minus.t2 drain_right.t5 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X7 source.t7 plus.t3 drain_left.t4 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 source.t9 plus.t4 drain_left.t3 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X9 a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X10 drain_right.t4 minus.t3 source.t14 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X11 a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X12 a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X13 source.t10 plus.t5 drain_left.t2 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X14 drain_left.t1 plus.t6 source.t5 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X15 drain_right.t3 minus.t4 source.t15 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X16 drain_right.t2 minus.t5 source.t0 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X17 drain_right.t1 minus.t6 source.t3 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X18 source.t6 plus.t7 drain_left.t0 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X19 source.t2 minus.t7 drain_right.t0 a_n1296_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
R0 plus.n1 plus.t4 1625.36
R1 plus.n5 plus.t0 1625.36
R2 plus.n8 plus.t2 1625.36
R3 plus.n12 plus.t3 1625.36
R4 plus.n2 plus.t1 1571.32
R5 plus.n4 plus.t5 1571.32
R6 plus.n9 plus.t7 1571.32
R7 plus.n11 plus.t6 1571.32
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 29.0483
R23 plus plus.n6 13.2808
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n3 source.t9 45.521
R27 source.n4 source.t0 45.521
R28 source.n7 source.t1 45.521
R29 source.n15 source.t3 45.5208
R30 source.n12 source.t13 45.5208
R31 source.n11 source.t8 45.5208
R32 source.n8 source.t7 45.5208
R33 source.n0 source.t4 45.5208
R34 source.n2 source.n1 44.201
R35 source.n6 source.n5 44.201
R36 source.n14 source.n13 44.2008
R37 source.n10 source.n9 44.2008
R38 source.n8 source.n7 24.0605
R39 source.n16 source.n0 18.5475
R40 source.n16 source.n15 5.51343
R41 source.n13 source.t14 1.3205
R42 source.n13 source.t2 1.3205
R43 source.n9 source.t5 1.3205
R44 source.n9 source.t6 1.3205
R45 source.n1 source.t11 1.3205
R46 source.n1 source.t10 1.3205
R47 source.n5 source.t15 1.3205
R48 source.n5 source.t12 1.3205
R49 source.n7 source.n6 0.5005
R50 source.n6 source.n4 0.5005
R51 source.n3 source.n2 0.5005
R52 source.n2 source.n0 0.5005
R53 source.n10 source.n8 0.5005
R54 source.n11 source.n10 0.5005
R55 source.n14 source.n12 0.5005
R56 source.n15 source.n14 0.5005
R57 source.n4 source.n3 0.470328
R58 source.n12 source.n11 0.470328
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 61.3798
R61 drain_left.n2 drain_left.n1 61.0742
R62 drain_left.n2 drain_left.n0 61.0742
R63 drain_left.n5 drain_left.n4 60.8796
R64 drain_left drain_left.n2 31.3898
R65 drain_left drain_left.n5 6.15322
R66 drain_left.n1 drain_left.t0 1.3205
R67 drain_left.n1 drain_left.t5 1.3205
R68 drain_left.n0 drain_left.t4 1.3205
R69 drain_left.n0 drain_left.t1 1.3205
R70 drain_left.n4 drain_left.t2 1.3205
R71 drain_left.n4 drain_left.t7 1.3205
R72 drain_left.n3 drain_left.t3 1.3205
R73 drain_left.n3 drain_left.t6 1.3205
R74 minus.n5 minus.t0 1625.36
R75 minus.n1 minus.t5 1625.36
R76 minus.n12 minus.t6 1625.36
R77 minus.n8 minus.t2 1625.36
R78 minus.n4 minus.t4 1571.32
R79 minus.n2 minus.t1 1571.32
R80 minus.n11 minus.t7 1571.32
R81 minus.n9 minus.t3 1571.32
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 42.3581
R89 minus.n3 minus.n2 42.3581
R90 minus.n10 minus.n9 42.3581
R91 minus.n11 minus.n10 42.3581
R92 minus.n14 minus.n6 36.3035
R93 minus.n5 minus.n4 30.6732
R94 minus.n2 minus.n1 30.6732
R95 minus.n9 minus.n8 30.6732
R96 minus.n12 minus.n11 30.6732
R97 minus.n14 minus.n13 6.5005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 61.3796
R102 drain_right.n2 drain_right.n1 61.0742
R103 drain_right.n2 drain_right.n0 61.0742
R104 drain_right.n5 drain_right.n4 60.8798
R105 drain_right drain_right.n2 30.8366
R106 drain_right drain_right.n5 6.15322
R107 drain_right.n1 drain_right.t0 1.3205
R108 drain_right.n1 drain_right.t1 1.3205
R109 drain_right.n0 drain_right.t5 1.3205
R110 drain_right.n0 drain_right.t4 1.3205
R111 drain_right.n3 drain_right.t6 1.3205
R112 drain_right.n3 drain_right.t2 1.3205
R113 drain_right.n4 drain_right.t7 1.3205
R114 drain_right.n4 drain_right.t3 1.3205
C0 source minus 3.07681f
C1 minus plus 5.32169f
C2 drain_right drain_left 0.605638f
C3 drain_right source 21.9694f
C4 drain_right plus 0.275273f
C5 drain_right minus 3.6673f
C6 source drain_left 21.970499f
C7 drain_left plus 3.78929f
C8 drain_left minus 0.170438f
C9 source plus 3.09085f
C10 drain_right a_n1296_n3888# 6.55053f
C11 drain_left a_n1296_n3888# 6.74519f
C12 source a_n1296_n3888# 10.080214f
C13 minus a_n1296_n3888# 5.181356f
C14 plus a_n1296_n3888# 7.474121f
C15 drain_right.t5 a_n1296_n3888# 0.418587f
C16 drain_right.t4 a_n1296_n3888# 0.418587f
C17 drain_right.n0 a_n1296_n3888# 3.78477f
C18 drain_right.t0 a_n1296_n3888# 0.418587f
C19 drain_right.t1 a_n1296_n3888# 0.418587f
C20 drain_right.n1 a_n1296_n3888# 3.78477f
C21 drain_right.n2 a_n1296_n3888# 2.4712f
C22 drain_right.t6 a_n1296_n3888# 0.418587f
C23 drain_right.t2 a_n1296_n3888# 0.418587f
C24 drain_right.n3 a_n1296_n3888# 3.78693f
C25 drain_right.t7 a_n1296_n3888# 0.418587f
C26 drain_right.t3 a_n1296_n3888# 0.418587f
C27 drain_right.n4 a_n1296_n3888# 3.78354f
C28 drain_right.n5 a_n1296_n3888# 1.10838f
C29 minus.n0 a_n1296_n3888# 0.132202f
C30 minus.t0 a_n1296_n3888# 0.61594f
C31 minus.t4 a_n1296_n3888# 0.607936f
C32 minus.t1 a_n1296_n3888# 0.607936f
C33 minus.t5 a_n1296_n3888# 0.61594f
C34 minus.n1 a_n1296_n3888# 0.254697f
C35 minus.n2 a_n1296_n3888# 0.236464f
C36 minus.n3 a_n1296_n3888# 0.021897f
C37 minus.n4 a_n1296_n3888# 0.236464f
C38 minus.n5 a_n1296_n3888# 0.25461f
C39 minus.n6 a_n1296_n3888# 2.04051f
C40 minus.n7 a_n1296_n3888# 0.132202f
C41 minus.t7 a_n1296_n3888# 0.607936f
C42 minus.t3 a_n1296_n3888# 0.607936f
C43 minus.t2 a_n1296_n3888# 0.61594f
C44 minus.n8 a_n1296_n3888# 0.254697f
C45 minus.n9 a_n1296_n3888# 0.236464f
C46 minus.n10 a_n1296_n3888# 0.021897f
C47 minus.n11 a_n1296_n3888# 0.236464f
C48 minus.t6 a_n1296_n3888# 0.61594f
C49 minus.n12 a_n1296_n3888# 0.25461f
C50 minus.n13 a_n1296_n3888# 0.375757f
C51 minus.n14 a_n1296_n3888# 2.47782f
C52 drain_left.t4 a_n1296_n3888# 0.417969f
C53 drain_left.t1 a_n1296_n3888# 0.417969f
C54 drain_left.n0 a_n1296_n3888# 3.77918f
C55 drain_left.t0 a_n1296_n3888# 0.417969f
C56 drain_left.t5 a_n1296_n3888# 0.417969f
C57 drain_left.n1 a_n1296_n3888# 3.77918f
C58 drain_left.n2 a_n1296_n3888# 2.54166f
C59 drain_left.t3 a_n1296_n3888# 0.417969f
C60 drain_left.t6 a_n1296_n3888# 0.417969f
C61 drain_left.n3 a_n1296_n3888# 3.78135f
C62 drain_left.t2 a_n1296_n3888# 0.417969f
C63 drain_left.t7 a_n1296_n3888# 0.417969f
C64 drain_left.n4 a_n1296_n3888# 3.77794f
C65 drain_left.n5 a_n1296_n3888# 1.10674f
C66 source.t4 a_n1296_n3888# 3.32332f
C67 source.n0 a_n1296_n3888# 1.53369f
C68 source.t11 a_n1296_n3888# 0.29655f
C69 source.t10 a_n1296_n3888# 0.29655f
C70 source.n1 a_n1296_n3888# 2.60494f
C71 source.n2 a_n1296_n3888# 0.327044f
C72 source.t9 a_n1296_n3888# 3.32332f
C73 source.n3 a_n1296_n3888# 0.415003f
C74 source.t0 a_n1296_n3888# 3.32332f
C75 source.n4 a_n1296_n3888# 0.415003f
C76 source.t15 a_n1296_n3888# 0.29655f
C77 source.t12 a_n1296_n3888# 0.29655f
C78 source.n5 a_n1296_n3888# 2.60494f
C79 source.n6 a_n1296_n3888# 0.327044f
C80 source.t1 a_n1296_n3888# 3.32332f
C81 source.n7 a_n1296_n3888# 1.94829f
C82 source.t7 a_n1296_n3888# 3.32332f
C83 source.n8 a_n1296_n3888# 1.9483f
C84 source.t5 a_n1296_n3888# 0.29655f
C85 source.t6 a_n1296_n3888# 0.29655f
C86 source.n9 a_n1296_n3888# 2.60494f
C87 source.n10 a_n1296_n3888# 0.327047f
C88 source.t8 a_n1296_n3888# 3.32332f
C89 source.n11 a_n1296_n3888# 0.415007f
C90 source.t13 a_n1296_n3888# 3.32332f
C91 source.n12 a_n1296_n3888# 0.415007f
C92 source.t14 a_n1296_n3888# 0.29655f
C93 source.t2 a_n1296_n3888# 0.29655f
C94 source.n13 a_n1296_n3888# 2.60494f
C95 source.n14 a_n1296_n3888# 0.327047f
C96 source.t3 a_n1296_n3888# 3.32332f
C97 source.n15 a_n1296_n3888# 0.553452f
C98 source.n16 a_n1296_n3888# 1.82724f
C99 plus.n0 a_n1296_n3888# 0.134587f
C100 plus.t5 a_n1296_n3888# 0.618905f
C101 plus.t1 a_n1296_n3888# 0.618905f
C102 plus.t4 a_n1296_n3888# 0.627053f
C103 plus.n1 a_n1296_n3888# 0.259293f
C104 plus.n2 a_n1296_n3888# 0.240731f
C105 plus.n3 a_n1296_n3888# 0.022292f
C106 plus.n4 a_n1296_n3888# 0.240731f
C107 plus.t0 a_n1296_n3888# 0.627053f
C108 plus.n5 a_n1296_n3888# 0.259203f
C109 plus.n6 a_n1296_n3888# 0.739341f
C110 plus.n7 a_n1296_n3888# 0.134587f
C111 plus.t3 a_n1296_n3888# 0.627053f
C112 plus.t6 a_n1296_n3888# 0.618905f
C113 plus.t7 a_n1296_n3888# 0.618905f
C114 plus.t2 a_n1296_n3888# 0.627053f
C115 plus.n8 a_n1296_n3888# 0.259293f
C116 plus.n9 a_n1296_n3888# 0.240731f
C117 plus.n10 a_n1296_n3888# 0.022292f
C118 plus.n11 a_n1296_n3888# 0.240731f
C119 plus.n12 a_n1296_n3888# 0.259203f
C120 plus.n13 a_n1296_n3888# 1.69963f
.ends

