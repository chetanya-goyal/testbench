* NGSPICE file created from diffpair163.ext - technology: sky130A

.subckt diffpair163 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t6 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 source.t14 plus.t0 drain_left.t7 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X3 drain_left.t6 plus.t1 source.t3 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X4 source.t10 minus.t1 drain_right.t6 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X5 a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X6 source.t9 minus.t2 drain_right.t5 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X7 source.t0 plus.t2 drain_left.t5 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X8 drain_right.t4 minus.t3 source.t8 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X9 source.t13 minus.t4 drain_right.t3 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X10 drain_left.t4 plus.t3 source.t15 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X11 source.t1 plus.t4 drain_left.t3 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X12 drain_right.t2 minus.t5 source.t11 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X13 drain_left.t2 plus.t5 source.t2 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X14 drain_right.t1 minus.t6 source.t12 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X15 a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X16 a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X17 source.t5 plus.t6 drain_left.t1 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 drain_left.t0 plus.t7 source.t4 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X19 source.t7 minus.t7 drain_right.t0 a_n1366_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
R0 minus.n5 minus.t4 760.245
R1 minus.n1 minus.t3 760.245
R2 minus.n12 minus.t6 760.245
R3 minus.n8 minus.t1 760.245
R4 minus.n4 minus.t5 690.867
R5 minus.n2 minus.t2 690.867
R6 minus.n11 minus.t7 690.867
R7 minus.n9 minus.t0 690.867
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 27.5573
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n0 source.t2 73.0943
R28 source.n3 source.t1 73.0943
R29 source.n4 source.t8 73.0943
R30 source.n7 source.t13 73.0943
R31 source.n15 source.t12 73.0942
R32 source.n12 source.t10 73.0942
R33 source.n11 source.t3 73.0942
R34 source.n8 source.t0 73.0942
R35 source.n2 source.n1 63.0943
R36 source.n6 source.n5 63.0943
R37 source.n14 source.n13 63.0942
R38 source.n10 source.n9 63.0942
R39 source.n8 source.n7 15.0299
R40 source.n13 source.t6 10.0005
R41 source.n13 source.t7 10.0005
R42 source.n9 source.t15 10.0005
R43 source.n9 source.t14 10.0005
R44 source.n1 source.t4 10.0005
R45 source.n1 source.t5 10.0005
R46 source.n5 source.t11 10.0005
R47 source.n5 source.t9 10.0005
R48 source.n16 source.n0 9.48679
R49 source.n16 source.n15 5.5436
R50 source.n7 source.n6 0.560845
R51 source.n6 source.n4 0.560845
R52 source.n3 source.n2 0.560845
R53 source.n2 source.n0 0.560845
R54 source.n10 source.n8 0.560845
R55 source.n11 source.n10 0.560845
R56 source.n14 source.n12 0.560845
R57 source.n15 source.n14 0.560845
R58 source.n4 source.n3 0.470328
R59 source.n12 source.n11 0.470328
R60 source source.n16 0.188
R61 drain_right.n5 drain_right.n3 80.3335
R62 drain_right.n2 drain_right.n1 79.9978
R63 drain_right.n2 drain_right.n0 79.9978
R64 drain_right.n5 drain_right.n4 79.7731
R65 drain_right drain_right.n2 21.9569
R66 drain_right.n1 drain_right.t0 10.0005
R67 drain_right.n1 drain_right.t1 10.0005
R68 drain_right.n0 drain_right.t6 10.0005
R69 drain_right.n0 drain_right.t7 10.0005
R70 drain_right.n3 drain_right.t5 10.0005
R71 drain_right.n3 drain_right.t4 10.0005
R72 drain_right.n4 drain_right.t3 10.0005
R73 drain_right.n4 drain_right.t2 10.0005
R74 drain_right drain_right.n5 6.21356
R75 plus.n1 plus.t4 760.245
R76 plus.n5 plus.t5 760.245
R77 plus.n8 plus.t1 760.245
R78 plus.n12 plus.t2 760.245
R79 plus.n2 plus.t7 690.867
R80 plus.n4 plus.t6 690.867
R81 plus.n9 plus.t0 690.867
R82 plus.n11 plus.t3 690.867
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus.n2 plus.n1 25.5611
R94 plus.n5 plus.n4 25.5611
R95 plus.n12 plus.n11 25.5611
R96 plus.n9 plus.n8 25.5611
R97 plus plus.n13 24.8475
R98 plus plus.n6 8.81489
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 80.3335
R102 drain_left.n2 drain_left.n1 79.9978
R103 drain_left.n2 drain_left.n0 79.9978
R104 drain_left.n5 drain_left.n4 79.7731
R105 drain_left drain_left.n2 22.5101
R106 drain_left.n1 drain_left.t7 10.0005
R107 drain_left.n1 drain_left.t6 10.0005
R108 drain_left.n0 drain_left.t5 10.0005
R109 drain_left.n0 drain_left.t4 10.0005
R110 drain_left.n4 drain_left.t1 10.0005
R111 drain_left.n4 drain_left.t2 10.0005
R112 drain_left.n3 drain_left.t3 10.0005
R113 drain_left.n3 drain_left.t0 10.0005
R114 drain_left drain_left.n5 6.21356
C0 source drain_left 5.6175f
C1 drain_left plus 0.934686f
C2 drain_left minus 0.175459f
C3 source plus 0.765875f
C4 source minus 0.751877f
C5 minus plus 3.17498f
C6 drain_right drain_left 0.640281f
C7 drain_right source 5.61683f
C8 drain_right plus 0.28799f
C9 drain_right minus 0.805282f
C10 drain_right a_n1366_n1488# 3.29483f
C11 drain_left a_n1366_n1488# 3.46306f
C12 source a_n1366_n1488# 3.49915f
C13 minus a_n1366_n1488# 4.283154f
C14 plus a_n1366_n1488# 5.16203f
C15 drain_left.t5 a_n1366_n1488# 0.083228f
C16 drain_left.t4 a_n1366_n1488# 0.083228f
C17 drain_left.n0 a_n1366_n1488# 0.453465f
C18 drain_left.t7 a_n1366_n1488# 0.083228f
C19 drain_left.t6 a_n1366_n1488# 0.083228f
C20 drain_left.n1 a_n1366_n1488# 0.453465f
C21 drain_left.n2 a_n1366_n1488# 1.10227f
C22 drain_left.t3 a_n1366_n1488# 0.083228f
C23 drain_left.t0 a_n1366_n1488# 0.083228f
C24 drain_left.n3 a_n1366_n1488# 0.45469f
C25 drain_left.t1 a_n1366_n1488# 0.083228f
C26 drain_left.t2 a_n1366_n1488# 0.083228f
C27 drain_left.n4 a_n1366_n1488# 0.452748f
C28 drain_left.n5 a_n1366_n1488# 0.739182f
C29 plus.n0 a_n1366_n1488# 0.093687f
C30 plus.t6 a_n1366_n1488# 0.05155f
C31 plus.t7 a_n1366_n1488# 0.05155f
C32 plus.t4 a_n1366_n1488# 0.055116f
C33 plus.n1 a_n1366_n1488# 0.052357f
C34 plus.n2 a_n1366_n1488# 0.03603f
C35 plus.n3 a_n1366_n1488# 0.016781f
C36 plus.n4 a_n1366_n1488# 0.03603f
C37 plus.t5 a_n1366_n1488# 0.055116f
C38 plus.n5 a_n1366_n1488# 0.052293f
C39 plus.n6 a_n1366_n1488# 0.303322f
C40 plus.n7 a_n1366_n1488# 0.093687f
C41 plus.t2 a_n1366_n1488# 0.055116f
C42 plus.t3 a_n1366_n1488# 0.05155f
C43 plus.t0 a_n1366_n1488# 0.05155f
C44 plus.t1 a_n1366_n1488# 0.055116f
C45 plus.n8 a_n1366_n1488# 0.052357f
C46 plus.n9 a_n1366_n1488# 0.03603f
C47 plus.n10 a_n1366_n1488# 0.016781f
C48 plus.n11 a_n1366_n1488# 0.03603f
C49 plus.n12 a_n1366_n1488# 0.052293f
C50 plus.n13 a_n1366_n1488# 0.841495f
C51 drain_right.t6 a_n1366_n1488# 0.084597f
C52 drain_right.t7 a_n1366_n1488# 0.084597f
C53 drain_right.n0 a_n1366_n1488# 0.460925f
C54 drain_right.t0 a_n1366_n1488# 0.084597f
C55 drain_right.t1 a_n1366_n1488# 0.084597f
C56 drain_right.n1 a_n1366_n1488# 0.460925f
C57 drain_right.n2 a_n1366_n1488# 1.07345f
C58 drain_right.t5 a_n1366_n1488# 0.084597f
C59 drain_right.t4 a_n1366_n1488# 0.084597f
C60 drain_right.n3 a_n1366_n1488# 0.462171f
C61 drain_right.t3 a_n1366_n1488# 0.084597f
C62 drain_right.t2 a_n1366_n1488# 0.084597f
C63 drain_right.n4 a_n1366_n1488# 0.460197f
C64 drain_right.n5 a_n1366_n1488# 0.751343f
C65 source.t2 a_n1366_n1488# 0.44515f
C66 source.n0 a_n1366_n1488# 0.587654f
C67 source.t4 a_n1366_n1488# 0.07558f
C68 source.t5 a_n1366_n1488# 0.07558f
C69 source.n1 a_n1366_n1488# 0.36768f
C70 source.n2 a_n1366_n1488# 0.259282f
C71 source.t1 a_n1366_n1488# 0.44515f
C72 source.n3 a_n1366_n1488# 0.311719f
C73 source.t8 a_n1366_n1488# 0.44515f
C74 source.n4 a_n1366_n1488# 0.311719f
C75 source.t11 a_n1366_n1488# 0.07558f
C76 source.t9 a_n1366_n1488# 0.07558f
C77 source.n5 a_n1366_n1488# 0.36768f
C78 source.n6 a_n1366_n1488# 0.259282f
C79 source.t13 a_n1366_n1488# 0.44515f
C80 source.n7 a_n1366_n1488# 0.807262f
C81 source.t0 a_n1366_n1488# 0.445148f
C82 source.n8 a_n1366_n1488# 0.807265f
C83 source.t15 a_n1366_n1488# 0.07558f
C84 source.t14 a_n1366_n1488# 0.07558f
C85 source.n9 a_n1366_n1488# 0.367678f
C86 source.n10 a_n1366_n1488# 0.259284f
C87 source.t3 a_n1366_n1488# 0.445148f
C88 source.n11 a_n1366_n1488# 0.311721f
C89 source.t10 a_n1366_n1488# 0.445148f
C90 source.n12 a_n1366_n1488# 0.311721f
C91 source.t6 a_n1366_n1488# 0.07558f
C92 source.t7 a_n1366_n1488# 0.07558f
C93 source.n13 a_n1366_n1488# 0.367678f
C94 source.n14 a_n1366_n1488# 0.259284f
C95 source.t12 a_n1366_n1488# 0.445148f
C96 source.n15 a_n1366_n1488# 0.431434f
C97 source.n16 a_n1366_n1488# 0.610405f
C98 minus.n0 a_n1366_n1488# 0.091402f
C99 minus.t4 a_n1366_n1488# 0.053772f
C100 minus.t5 a_n1366_n1488# 0.050293f
C101 minus.t2 a_n1366_n1488# 0.050293f
C102 minus.t3 a_n1366_n1488# 0.053772f
C103 minus.n1 a_n1366_n1488# 0.05108f
C104 minus.n2 a_n1366_n1488# 0.035151f
C105 minus.n3 a_n1366_n1488# 0.016372f
C106 minus.n4 a_n1366_n1488# 0.035151f
C107 minus.n5 a_n1366_n1488# 0.051018f
C108 minus.n6 a_n1366_n1488# 0.868748f
C109 minus.n7 a_n1366_n1488# 0.091402f
C110 minus.t7 a_n1366_n1488# 0.050293f
C111 minus.t0 a_n1366_n1488# 0.050293f
C112 minus.t1 a_n1366_n1488# 0.053772f
C113 minus.n8 a_n1366_n1488# 0.05108f
C114 minus.n9 a_n1366_n1488# 0.035151f
C115 minus.n10 a_n1366_n1488# 0.016372f
C116 minus.n11 a_n1366_n1488# 0.035151f
C117 minus.t6 a_n1366_n1488# 0.053772f
C118 minus.n12 a_n1366_n1488# 0.051018f
C119 minus.n13 a_n1366_n1488# 0.259564f
C120 minus.n14 a_n1366_n1488# 1.06974f
.ends

