* NGSPICE file created from diffpair53.ext - technology: sky130A

.subckt diffpair53 minus drain_right drain_left source plus
X0 a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X1 a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X2 source.t15 plus.t0 drain_left.t4 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X3 a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X4 source.t0 minus.t0 drain_right.t7 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 drain_right.t6 minus.t1 source.t7 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X6 source.t1 minus.t2 drain_right.t5 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X7 drain_right.t4 minus.t3 source.t4 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 drain_left.t2 plus.t1 source.t14 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X9 drain_left.t6 plus.t2 source.t13 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X10 source.t6 minus.t4 drain_right.t3 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 source.t12 plus.t3 drain_left.t5 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X12 drain_right.t2 minus.t5 source.t2 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X13 drain_left.t3 plus.t4 source.t11 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 source.t10 plus.t5 drain_left.t1 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X15 a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X16 source.t9 plus.t6 drain_left.t0 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X17 drain_right.t1 minus.t6 source.t3 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X18 source.t5 minus.t7 drain_right.t0 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X19 drain_left.t7 plus.t7 source.t8 a_n1646_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n5 plus.n4 161.3
R1 plus.n11 plus.n10 161.3
R2 plus.n1 plus.t5 132.459
R3 plus.n7 plus.t1 132.459
R4 plus.n4 plus.t2 105.638
R5 plus.n3 plus.t3 105.638
R6 plus.n2 plus.t4 105.638
R7 plus.n10 plus.t6 105.638
R8 plus.n9 plus.t7 105.638
R9 plus.n8 plus.t0 105.638
R10 plus.n3 plus.n0 80.6037
R11 plus.n9 plus.n6 80.6037
R12 plus.n4 plus.n3 48.2005
R13 plus.n3 plus.n2 48.2005
R14 plus.n10 plus.n9 48.2005
R15 plus.n9 plus.n8 48.2005
R16 plus.n1 plus.n0 45.2318
R17 plus.n7 plus.n6 45.2318
R18 plus plus.n11 25.1846
R19 plus.n2 plus.n1 13.3799
R20 plus.n8 plus.n7 13.3799
R21 plus plus.n5 8.09141
R22 plus.n5 plus.n0 0.285035
R23 plus.n11 plus.n6 0.285035
R24 drain_left.n5 drain_left.n3 240.935
R25 drain_left.n2 drain_left.n1 240.477
R26 drain_left.n2 drain_left.n0 240.477
R27 drain_left.n5 drain_left.n4 240.132
R28 drain_left drain_left.n2 21.8398
R29 drain_left.n1 drain_left.t4 19.8005
R30 drain_left.n1 drain_left.t2 19.8005
R31 drain_left.n0 drain_left.t0 19.8005
R32 drain_left.n0 drain_left.t7 19.8005
R33 drain_left.n4 drain_left.t5 19.8005
R34 drain_left.n4 drain_left.t6 19.8005
R35 drain_left.n3 drain_left.t1 19.8005
R36 drain_left.n3 drain_left.t3 19.8005
R37 drain_left drain_left.n5 6.45494
R38 source.n0 source.t13 243.255
R39 source.n3 source.t10 243.255
R40 source.n4 source.t2 243.255
R41 source.n7 source.t1 243.255
R42 source.n15 source.t3 243.254
R43 source.n12 source.t5 243.254
R44 source.n11 source.t14 243.254
R45 source.n8 source.t9 243.254
R46 source.n2 source.n1 223.454
R47 source.n6 source.n5 223.454
R48 source.n14 source.n13 223.453
R49 source.n10 source.n9 223.453
R50 source.n13 source.t7 19.8005
R51 source.n13 source.t0 19.8005
R52 source.n9 source.t8 19.8005
R53 source.n9 source.t15 19.8005
R54 source.n1 source.t11 19.8005
R55 source.n1 source.t12 19.8005
R56 source.n5 source.t4 19.8005
R57 source.n5 source.t6 19.8005
R58 source.n8 source.n7 13.7561
R59 source.n16 source.n0 8.09232
R60 source.n16 source.n15 5.66429
R61 source.n7 source.n6 0.802224
R62 source.n6 source.n4 0.802224
R63 source.n3 source.n2 0.802224
R64 source.n2 source.n0 0.802224
R65 source.n10 source.n8 0.802224
R66 source.n11 source.n10 0.802224
R67 source.n14 source.n12 0.802224
R68 source.n15 source.n14 0.802224
R69 source.n4 source.n3 0.470328
R70 source.n12 source.n11 0.470328
R71 source source.n16 0.188
R72 minus.n5 minus.n4 161.3
R73 minus.n11 minus.n10 161.3
R74 minus.n1 minus.t5 132.459
R75 minus.n7 minus.t7 132.459
R76 minus.n2 minus.t4 105.638
R77 minus.n3 minus.t3 105.638
R78 minus.n4 minus.t2 105.638
R79 minus.n8 minus.t1 105.638
R80 minus.n9 minus.t0 105.638
R81 minus.n10 minus.t6 105.638
R82 minus.n3 minus.n0 80.6037
R83 minus.n9 minus.n6 80.6037
R84 minus.n3 minus.n2 48.2005
R85 minus.n4 minus.n3 48.2005
R86 minus.n9 minus.n8 48.2005
R87 minus.n10 minus.n9 48.2005
R88 minus.n1 minus.n0 45.2318
R89 minus.n7 minus.n6 45.2318
R90 minus.n12 minus.n5 27.1369
R91 minus.n2 minus.n1 13.3799
R92 minus.n8 minus.n7 13.3799
R93 minus.n12 minus.n11 6.61414
R94 minus.n5 minus.n0 0.285035
R95 minus.n11 minus.n6 0.285035
R96 minus minus.n12 0.188
R97 drain_right.n5 drain_right.n3 240.935
R98 drain_right.n2 drain_right.n1 240.477
R99 drain_right.n2 drain_right.n0 240.477
R100 drain_right.n5 drain_right.n4 240.132
R101 drain_right drain_right.n2 21.2865
R102 drain_right.n1 drain_right.t7 19.8005
R103 drain_right.n1 drain_right.t1 19.8005
R104 drain_right.n0 drain_right.t0 19.8005
R105 drain_right.n0 drain_right.t6 19.8005
R106 drain_right.n3 drain_right.t3 19.8005
R107 drain_right.n3 drain_right.t2 19.8005
R108 drain_right.n4 drain_right.t5 19.8005
R109 drain_right.n4 drain_right.t4 19.8005
R110 drain_right drain_right.n5 6.45494
C0 drain_right source 2.90573f
C1 source plus 1.09889f
C2 minus drain_left 0.178437f
C3 drain_right minus 0.772271f
C4 minus plus 3.16769f
C5 drain_right drain_left 0.776011f
C6 plus drain_left 0.930596f
C7 source minus 1.08502f
C8 drain_right plus 0.321038f
C9 source drain_left 2.9046f
C10 drain_right a_n1646_n1088# 3.055085f
C11 drain_left a_n1646_n1088# 3.257414f
C12 source a_n1646_n1088# 2.404576f
C13 minus a_n1646_n1088# 5.453362f
C14 plus a_n1646_n1088# 6.107221f
C15 drain_right.t0 a_n1646_n1088# 0.015779f
C16 drain_right.t6 a_n1646_n1088# 0.015779f
C17 drain_right.n0 a_n1646_n1088# 0.061632f
C18 drain_right.t7 a_n1646_n1088# 0.015779f
C19 drain_right.t1 a_n1646_n1088# 0.015779f
C20 drain_right.n1 a_n1646_n1088# 0.061632f
C21 drain_right.n2 a_n1646_n1088# 0.919248f
C22 drain_right.t3 a_n1646_n1088# 0.015779f
C23 drain_right.t2 a_n1646_n1088# 0.015779f
C24 drain_right.n3 a_n1646_n1088# 0.062146f
C25 drain_right.t5 a_n1646_n1088# 0.015779f
C26 drain_right.t4 a_n1646_n1088# 0.015779f
C27 drain_right.n4 a_n1646_n1088# 0.061312f
C28 drain_right.n5 a_n1646_n1088# 0.666916f
C29 minus.n0 a_n1646_n1088# 0.155127f
C30 minus.t4 a_n1646_n1088# 0.064728f
C31 minus.t5 a_n1646_n1088# 0.078086f
C32 minus.n1 a_n1646_n1088# 0.053479f
C33 minus.n2 a_n1646_n1088# 0.073103f
C34 minus.t3 a_n1646_n1088# 0.064728f
C35 minus.n3 a_n1646_n1088# 0.073103f
C36 minus.t2 a_n1646_n1088# 0.064728f
C37 minus.n4 a_n1646_n1088# 0.065884f
C38 minus.n5 a_n1646_n1088# 0.708521f
C39 minus.n6 a_n1646_n1088# 0.155127f
C40 minus.t7 a_n1646_n1088# 0.078086f
C41 minus.n7 a_n1646_n1088# 0.053479f
C42 minus.t1 a_n1646_n1088# 0.064728f
C43 minus.n8 a_n1646_n1088# 0.073103f
C44 minus.t0 a_n1646_n1088# 0.064728f
C45 minus.n9 a_n1646_n1088# 0.073103f
C46 minus.t6 a_n1646_n1088# 0.064728f
C47 minus.n10 a_n1646_n1088# 0.065884f
C48 minus.n11 a_n1646_n1088# 0.227136f
C49 minus.n12 a_n1646_n1088# 0.857518f
C50 source.t13 a_n1646_n1088# 0.099695f
C51 source.n0 a_n1646_n1088# 0.461833f
C52 source.t11 a_n1646_n1088# 0.017912f
C53 source.t12 a_n1646_n1088# 0.017912f
C54 source.n1 a_n1646_n1088# 0.058091f
C55 source.n2 a_n1646_n1088# 0.256321f
C56 source.t10 a_n1646_n1088# 0.099695f
C57 source.n3 a_n1646_n1088# 0.239327f
C58 source.t2 a_n1646_n1088# 0.099695f
C59 source.n4 a_n1646_n1088# 0.239327f
C60 source.t4 a_n1646_n1088# 0.017912f
C61 source.t6 a_n1646_n1088# 0.017912f
C62 source.n5 a_n1646_n1088# 0.058091f
C63 source.n6 a_n1646_n1088# 0.256321f
C64 source.t1 a_n1646_n1088# 0.099695f
C65 source.n7 a_n1646_n1088# 0.647478f
C66 source.t9 a_n1646_n1088# 0.099694f
C67 source.n8 a_n1646_n1088# 0.647478f
C68 source.t8 a_n1646_n1088# 0.017912f
C69 source.t15 a_n1646_n1088# 0.017912f
C70 source.n9 a_n1646_n1088# 0.058091f
C71 source.n10 a_n1646_n1088# 0.256321f
C72 source.t14 a_n1646_n1088# 0.099694f
C73 source.n11 a_n1646_n1088# 0.239327f
C74 source.t5 a_n1646_n1088# 0.099694f
C75 source.n12 a_n1646_n1088# 0.239327f
C76 source.t7 a_n1646_n1088# 0.017912f
C77 source.t0 a_n1646_n1088# 0.017912f
C78 source.n13 a_n1646_n1088# 0.058091f
C79 source.n14 a_n1646_n1088# 0.256321f
C80 source.t3 a_n1646_n1088# 0.099694f
C81 source.n15 a_n1646_n1088# 0.382249f
C82 source.n16 a_n1646_n1088# 0.466997f
C83 drain_left.t0 a_n1646_n1088# 0.015365f
C84 drain_left.t7 a_n1646_n1088# 0.015365f
C85 drain_left.n0 a_n1646_n1088# 0.060015f
C86 drain_left.t4 a_n1646_n1088# 0.015365f
C87 drain_left.t2 a_n1646_n1088# 0.015365f
C88 drain_left.n1 a_n1646_n1088# 0.060015f
C89 drain_left.n2 a_n1646_n1088# 0.932773f
C90 drain_left.t1 a_n1646_n1088# 0.015365f
C91 drain_left.t3 a_n1646_n1088# 0.015365f
C92 drain_left.n3 a_n1646_n1088# 0.060516f
C93 drain_left.t5 a_n1646_n1088# 0.015365f
C94 drain_left.t6 a_n1646_n1088# 0.015365f
C95 drain_left.n4 a_n1646_n1088# 0.059704f
C96 drain_left.n5 a_n1646_n1088# 0.649424f
C97 plus.n0 a_n1646_n1088# 0.15831f
C98 plus.t2 a_n1646_n1088# 0.066056f
C99 plus.t3 a_n1646_n1088# 0.066056f
C100 plus.t4 a_n1646_n1088# 0.066056f
C101 plus.t5 a_n1646_n1088# 0.079688f
C102 plus.n1 a_n1646_n1088# 0.054576f
C103 plus.n2 a_n1646_n1088# 0.074603f
C104 plus.n3 a_n1646_n1088# 0.074603f
C105 plus.n4 a_n1646_n1088# 0.067236f
C106 plus.n5 a_n1646_n1088# 0.2426f
C107 plus.n6 a_n1646_n1088# 0.15831f
C108 plus.t6 a_n1646_n1088# 0.066056f
C109 plus.t7 a_n1646_n1088# 0.066056f
C110 plus.t1 a_n1646_n1088# 0.079688f
C111 plus.n7 a_n1646_n1088# 0.054576f
C112 plus.t0 a_n1646_n1088# 0.066056f
C113 plus.n8 a_n1646_n1088# 0.074603f
C114 plus.n9 a_n1646_n1088# 0.074603f
C115 plus.n10 a_n1646_n1088# 0.067236f
C116 plus.n11 a_n1646_n1088# 0.7034f
.ends

