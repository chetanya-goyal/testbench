* NGSPICE file created from diffpair705.ext - technology: sky130A

.subckt diffpair705 minus drain_right drain_left source plus
X0 source.t20 minus.t0 drain_right.t6 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X1 source.t21 plus.t0 drain_left.t11 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X2 drain_right.t3 minus.t1 source.t19 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X3 source.t22 plus.t1 drain_left.t10 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X4 source.t18 minus.t2 drain_right.t2 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X5 a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.7
X6 source.t17 minus.t3 drain_right.t1 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X7 source.t2 plus.t2 drain_left.t9 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X8 source.t1 plus.t3 drain_left.t8 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X9 source.t7 plus.t4 drain_left.t7 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X10 drain_right.t0 minus.t4 source.t16 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X11 source.t15 minus.t5 drain_right.t8 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X12 drain_right.t7 minus.t6 source.t14 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X13 drain_right.t10 minus.t7 source.t13 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X14 source.t3 plus.t5 drain_left.t6 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X15 drain_left.t5 plus.t6 source.t5 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X16 drain_left.t4 plus.t7 source.t8 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X17 drain_left.t3 plus.t8 source.t0 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X18 a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X19 drain_right.t9 minus.t8 source.t12 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X20 drain_left.t2 plus.t9 source.t23 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X21 drain_left.t1 plus.t10 source.t4 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X22 a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X23 drain_right.t5 minus.t9 source.t11 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X24 source.t10 minus.t10 drain_right.t4 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X25 source.t9 minus.t11 drain_right.t11 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X26 a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X27 drain_left.t0 plus.t11 source.t6 a_n2158_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
R0 minus.n5 minus.t8 940.138
R1 minus.n23 minus.t5 940.138
R2 minus.n4 minus.t2 916.833
R3 minus.n8 minus.t7 916.833
R4 minus.n10 minus.t10 916.833
R5 minus.n14 minus.t6 916.833
R6 minus.n16 minus.t11 916.833
R7 minus.n22 minus.t4 916.833
R8 minus.n26 minus.t0 916.833
R9 minus.n28 minus.t1 916.833
R10 minus.n32 minus.t3 916.833
R11 minus.n34 minus.t9 916.833
R12 minus.n17 minus.n16 161.3
R13 minus.n15 minus.n0 161.3
R14 minus.n14 minus.n13 161.3
R15 minus.n12 minus.n1 161.3
R16 minus.n11 minus.n10 161.3
R17 minus.n9 minus.n2 161.3
R18 minus.n8 minus.n7 161.3
R19 minus.n6 minus.n3 161.3
R20 minus.n35 minus.n34 161.3
R21 minus.n33 minus.n18 161.3
R22 minus.n32 minus.n31 161.3
R23 minus.n30 minus.n19 161.3
R24 minus.n29 minus.n28 161.3
R25 minus.n27 minus.n20 161.3
R26 minus.n26 minus.n25 161.3
R27 minus.n24 minus.n21 161.3
R28 minus.n36 minus.n17 47.2884
R29 minus.n6 minus.n5 44.8907
R30 minus.n24 minus.n23 44.8907
R31 minus.n16 minus.n15 32.8641
R32 minus.n34 minus.n33 32.8641
R33 minus.n4 minus.n3 28.4823
R34 minus.n14 minus.n1 28.4823
R35 minus.n22 minus.n21 28.4823
R36 minus.n32 minus.n19 28.4823
R37 minus.n10 minus.n9 24.1005
R38 minus.n9 minus.n8 24.1005
R39 minus.n27 minus.n26 24.1005
R40 minus.n28 minus.n27 24.1005
R41 minus.n8 minus.n3 19.7187
R42 minus.n10 minus.n1 19.7187
R43 minus.n26 minus.n21 19.7187
R44 minus.n28 minus.n19 19.7187
R45 minus.n5 minus.n4 18.4104
R46 minus.n23 minus.n22 18.4104
R47 minus.n15 minus.n14 15.3369
R48 minus.n33 minus.n32 15.3369
R49 minus.n36 minus.n35 6.64444
R50 minus.n17 minus.n0 0.189894
R51 minus.n13 minus.n0 0.189894
R52 minus.n13 minus.n12 0.189894
R53 minus.n12 minus.n11 0.189894
R54 minus.n11 minus.n2 0.189894
R55 minus.n7 minus.n2 0.189894
R56 minus.n7 minus.n6 0.189894
R57 minus.n25 minus.n24 0.189894
R58 minus.n25 minus.n20 0.189894
R59 minus.n29 minus.n20 0.189894
R60 minus.n30 minus.n29 0.189894
R61 minus.n31 minus.n30 0.189894
R62 minus.n31 minus.n18 0.189894
R63 minus.n35 minus.n18 0.189894
R64 minus minus.n36 0.188
R65 drain_right.n6 drain_right.n4 59.6032
R66 drain_right.n3 drain_right.n2 59.548
R67 drain_right.n3 drain_right.n0 59.548
R68 drain_right.n3 drain_right.n1 58.7154
R69 drain_right.n6 drain_right.n5 58.7154
R70 drain_right.n8 drain_right.n7 58.7154
R71 drain_right drain_right.n3 41.102
R72 drain_right drain_right.n8 6.54115
R73 drain_right.n8 drain_right.n6 0.888431
R74 drain_right.n1 drain_right.t6 0.7925
R75 drain_right.n1 drain_right.t3 0.7925
R76 drain_right.n2 drain_right.t1 0.7925
R77 drain_right.n2 drain_right.t5 0.7925
R78 drain_right.n0 drain_right.t8 0.7925
R79 drain_right.n0 drain_right.t0 0.7925
R80 drain_right.n4 drain_right.t2 0.7925
R81 drain_right.n4 drain_right.t9 0.7925
R82 drain_right.n5 drain_right.t4 0.7925
R83 drain_right.n5 drain_right.t10 0.7925
R84 drain_right.n7 drain_right.t11 0.7925
R85 drain_right.n7 drain_right.t7 0.7925
R86 source.n1130 source.n996 289.615
R87 source.n986 source.n852 289.615
R88 source.n846 source.n712 289.615
R89 source.n702 source.n568 289.615
R90 source.n134 source.n0 289.615
R91 source.n278 source.n144 289.615
R92 source.n418 source.n284 289.615
R93 source.n562 source.n428 289.615
R94 source.n1040 source.n1039 185
R95 source.n1045 source.n1044 185
R96 source.n1047 source.n1046 185
R97 source.n1036 source.n1035 185
R98 source.n1053 source.n1052 185
R99 source.n1055 source.n1054 185
R100 source.n1032 source.n1031 185
R101 source.n1062 source.n1061 185
R102 source.n1063 source.n1030 185
R103 source.n1065 source.n1064 185
R104 source.n1028 source.n1027 185
R105 source.n1071 source.n1070 185
R106 source.n1073 source.n1072 185
R107 source.n1024 source.n1023 185
R108 source.n1079 source.n1078 185
R109 source.n1081 source.n1080 185
R110 source.n1020 source.n1019 185
R111 source.n1087 source.n1086 185
R112 source.n1089 source.n1088 185
R113 source.n1016 source.n1015 185
R114 source.n1095 source.n1094 185
R115 source.n1097 source.n1096 185
R116 source.n1012 source.n1011 185
R117 source.n1103 source.n1102 185
R118 source.n1106 source.n1105 185
R119 source.n1104 source.n1008 185
R120 source.n1111 source.n1007 185
R121 source.n1113 source.n1112 185
R122 source.n1115 source.n1114 185
R123 source.n1004 source.n1003 185
R124 source.n1121 source.n1120 185
R125 source.n1123 source.n1122 185
R126 source.n1000 source.n999 185
R127 source.n1129 source.n1128 185
R128 source.n1131 source.n1130 185
R129 source.n896 source.n895 185
R130 source.n901 source.n900 185
R131 source.n903 source.n902 185
R132 source.n892 source.n891 185
R133 source.n909 source.n908 185
R134 source.n911 source.n910 185
R135 source.n888 source.n887 185
R136 source.n918 source.n917 185
R137 source.n919 source.n886 185
R138 source.n921 source.n920 185
R139 source.n884 source.n883 185
R140 source.n927 source.n926 185
R141 source.n929 source.n928 185
R142 source.n880 source.n879 185
R143 source.n935 source.n934 185
R144 source.n937 source.n936 185
R145 source.n876 source.n875 185
R146 source.n943 source.n942 185
R147 source.n945 source.n944 185
R148 source.n872 source.n871 185
R149 source.n951 source.n950 185
R150 source.n953 source.n952 185
R151 source.n868 source.n867 185
R152 source.n959 source.n958 185
R153 source.n962 source.n961 185
R154 source.n960 source.n864 185
R155 source.n967 source.n863 185
R156 source.n969 source.n968 185
R157 source.n971 source.n970 185
R158 source.n860 source.n859 185
R159 source.n977 source.n976 185
R160 source.n979 source.n978 185
R161 source.n856 source.n855 185
R162 source.n985 source.n984 185
R163 source.n987 source.n986 185
R164 source.n756 source.n755 185
R165 source.n761 source.n760 185
R166 source.n763 source.n762 185
R167 source.n752 source.n751 185
R168 source.n769 source.n768 185
R169 source.n771 source.n770 185
R170 source.n748 source.n747 185
R171 source.n778 source.n777 185
R172 source.n779 source.n746 185
R173 source.n781 source.n780 185
R174 source.n744 source.n743 185
R175 source.n787 source.n786 185
R176 source.n789 source.n788 185
R177 source.n740 source.n739 185
R178 source.n795 source.n794 185
R179 source.n797 source.n796 185
R180 source.n736 source.n735 185
R181 source.n803 source.n802 185
R182 source.n805 source.n804 185
R183 source.n732 source.n731 185
R184 source.n811 source.n810 185
R185 source.n813 source.n812 185
R186 source.n728 source.n727 185
R187 source.n819 source.n818 185
R188 source.n822 source.n821 185
R189 source.n820 source.n724 185
R190 source.n827 source.n723 185
R191 source.n829 source.n828 185
R192 source.n831 source.n830 185
R193 source.n720 source.n719 185
R194 source.n837 source.n836 185
R195 source.n839 source.n838 185
R196 source.n716 source.n715 185
R197 source.n845 source.n844 185
R198 source.n847 source.n846 185
R199 source.n612 source.n611 185
R200 source.n617 source.n616 185
R201 source.n619 source.n618 185
R202 source.n608 source.n607 185
R203 source.n625 source.n624 185
R204 source.n627 source.n626 185
R205 source.n604 source.n603 185
R206 source.n634 source.n633 185
R207 source.n635 source.n602 185
R208 source.n637 source.n636 185
R209 source.n600 source.n599 185
R210 source.n643 source.n642 185
R211 source.n645 source.n644 185
R212 source.n596 source.n595 185
R213 source.n651 source.n650 185
R214 source.n653 source.n652 185
R215 source.n592 source.n591 185
R216 source.n659 source.n658 185
R217 source.n661 source.n660 185
R218 source.n588 source.n587 185
R219 source.n667 source.n666 185
R220 source.n669 source.n668 185
R221 source.n584 source.n583 185
R222 source.n675 source.n674 185
R223 source.n678 source.n677 185
R224 source.n676 source.n580 185
R225 source.n683 source.n579 185
R226 source.n685 source.n684 185
R227 source.n687 source.n686 185
R228 source.n576 source.n575 185
R229 source.n693 source.n692 185
R230 source.n695 source.n694 185
R231 source.n572 source.n571 185
R232 source.n701 source.n700 185
R233 source.n703 source.n702 185
R234 source.n135 source.n134 185
R235 source.n133 source.n132 185
R236 source.n4 source.n3 185
R237 source.n127 source.n126 185
R238 source.n125 source.n124 185
R239 source.n8 source.n7 185
R240 source.n119 source.n118 185
R241 source.n117 source.n116 185
R242 source.n115 source.n11 185
R243 source.n15 source.n12 185
R244 source.n110 source.n109 185
R245 source.n108 source.n107 185
R246 source.n17 source.n16 185
R247 source.n102 source.n101 185
R248 source.n100 source.n99 185
R249 source.n21 source.n20 185
R250 source.n94 source.n93 185
R251 source.n92 source.n91 185
R252 source.n25 source.n24 185
R253 source.n86 source.n85 185
R254 source.n84 source.n83 185
R255 source.n29 source.n28 185
R256 source.n78 source.n77 185
R257 source.n76 source.n75 185
R258 source.n33 source.n32 185
R259 source.n70 source.n69 185
R260 source.n68 source.n35 185
R261 source.n67 source.n66 185
R262 source.n38 source.n36 185
R263 source.n61 source.n60 185
R264 source.n59 source.n58 185
R265 source.n42 source.n41 185
R266 source.n53 source.n52 185
R267 source.n51 source.n50 185
R268 source.n46 source.n45 185
R269 source.n279 source.n278 185
R270 source.n277 source.n276 185
R271 source.n148 source.n147 185
R272 source.n271 source.n270 185
R273 source.n269 source.n268 185
R274 source.n152 source.n151 185
R275 source.n263 source.n262 185
R276 source.n261 source.n260 185
R277 source.n259 source.n155 185
R278 source.n159 source.n156 185
R279 source.n254 source.n253 185
R280 source.n252 source.n251 185
R281 source.n161 source.n160 185
R282 source.n246 source.n245 185
R283 source.n244 source.n243 185
R284 source.n165 source.n164 185
R285 source.n238 source.n237 185
R286 source.n236 source.n235 185
R287 source.n169 source.n168 185
R288 source.n230 source.n229 185
R289 source.n228 source.n227 185
R290 source.n173 source.n172 185
R291 source.n222 source.n221 185
R292 source.n220 source.n219 185
R293 source.n177 source.n176 185
R294 source.n214 source.n213 185
R295 source.n212 source.n179 185
R296 source.n211 source.n210 185
R297 source.n182 source.n180 185
R298 source.n205 source.n204 185
R299 source.n203 source.n202 185
R300 source.n186 source.n185 185
R301 source.n197 source.n196 185
R302 source.n195 source.n194 185
R303 source.n190 source.n189 185
R304 source.n419 source.n418 185
R305 source.n417 source.n416 185
R306 source.n288 source.n287 185
R307 source.n411 source.n410 185
R308 source.n409 source.n408 185
R309 source.n292 source.n291 185
R310 source.n403 source.n402 185
R311 source.n401 source.n400 185
R312 source.n399 source.n295 185
R313 source.n299 source.n296 185
R314 source.n394 source.n393 185
R315 source.n392 source.n391 185
R316 source.n301 source.n300 185
R317 source.n386 source.n385 185
R318 source.n384 source.n383 185
R319 source.n305 source.n304 185
R320 source.n378 source.n377 185
R321 source.n376 source.n375 185
R322 source.n309 source.n308 185
R323 source.n370 source.n369 185
R324 source.n368 source.n367 185
R325 source.n313 source.n312 185
R326 source.n362 source.n361 185
R327 source.n360 source.n359 185
R328 source.n317 source.n316 185
R329 source.n354 source.n353 185
R330 source.n352 source.n319 185
R331 source.n351 source.n350 185
R332 source.n322 source.n320 185
R333 source.n345 source.n344 185
R334 source.n343 source.n342 185
R335 source.n326 source.n325 185
R336 source.n337 source.n336 185
R337 source.n335 source.n334 185
R338 source.n330 source.n329 185
R339 source.n563 source.n562 185
R340 source.n561 source.n560 185
R341 source.n432 source.n431 185
R342 source.n555 source.n554 185
R343 source.n553 source.n552 185
R344 source.n436 source.n435 185
R345 source.n547 source.n546 185
R346 source.n545 source.n544 185
R347 source.n543 source.n439 185
R348 source.n443 source.n440 185
R349 source.n538 source.n537 185
R350 source.n536 source.n535 185
R351 source.n445 source.n444 185
R352 source.n530 source.n529 185
R353 source.n528 source.n527 185
R354 source.n449 source.n448 185
R355 source.n522 source.n521 185
R356 source.n520 source.n519 185
R357 source.n453 source.n452 185
R358 source.n514 source.n513 185
R359 source.n512 source.n511 185
R360 source.n457 source.n456 185
R361 source.n506 source.n505 185
R362 source.n504 source.n503 185
R363 source.n461 source.n460 185
R364 source.n498 source.n497 185
R365 source.n496 source.n463 185
R366 source.n495 source.n494 185
R367 source.n466 source.n464 185
R368 source.n489 source.n488 185
R369 source.n487 source.n486 185
R370 source.n470 source.n469 185
R371 source.n481 source.n480 185
R372 source.n479 source.n478 185
R373 source.n474 source.n473 185
R374 source.n1041 source.t11 149.524
R375 source.n897 source.t15 149.524
R376 source.n757 source.t6 149.524
R377 source.n613 source.t2 149.524
R378 source.n47 source.t0 149.524
R379 source.n191 source.t7 149.524
R380 source.n331 source.t12 149.524
R381 source.n475 source.t9 149.524
R382 source.n1045 source.n1039 104.615
R383 source.n1046 source.n1045 104.615
R384 source.n1046 source.n1035 104.615
R385 source.n1053 source.n1035 104.615
R386 source.n1054 source.n1053 104.615
R387 source.n1054 source.n1031 104.615
R388 source.n1062 source.n1031 104.615
R389 source.n1063 source.n1062 104.615
R390 source.n1064 source.n1063 104.615
R391 source.n1064 source.n1027 104.615
R392 source.n1071 source.n1027 104.615
R393 source.n1072 source.n1071 104.615
R394 source.n1072 source.n1023 104.615
R395 source.n1079 source.n1023 104.615
R396 source.n1080 source.n1079 104.615
R397 source.n1080 source.n1019 104.615
R398 source.n1087 source.n1019 104.615
R399 source.n1088 source.n1087 104.615
R400 source.n1088 source.n1015 104.615
R401 source.n1095 source.n1015 104.615
R402 source.n1096 source.n1095 104.615
R403 source.n1096 source.n1011 104.615
R404 source.n1103 source.n1011 104.615
R405 source.n1105 source.n1103 104.615
R406 source.n1105 source.n1104 104.615
R407 source.n1104 source.n1007 104.615
R408 source.n1113 source.n1007 104.615
R409 source.n1114 source.n1113 104.615
R410 source.n1114 source.n1003 104.615
R411 source.n1121 source.n1003 104.615
R412 source.n1122 source.n1121 104.615
R413 source.n1122 source.n999 104.615
R414 source.n1129 source.n999 104.615
R415 source.n1130 source.n1129 104.615
R416 source.n901 source.n895 104.615
R417 source.n902 source.n901 104.615
R418 source.n902 source.n891 104.615
R419 source.n909 source.n891 104.615
R420 source.n910 source.n909 104.615
R421 source.n910 source.n887 104.615
R422 source.n918 source.n887 104.615
R423 source.n919 source.n918 104.615
R424 source.n920 source.n919 104.615
R425 source.n920 source.n883 104.615
R426 source.n927 source.n883 104.615
R427 source.n928 source.n927 104.615
R428 source.n928 source.n879 104.615
R429 source.n935 source.n879 104.615
R430 source.n936 source.n935 104.615
R431 source.n936 source.n875 104.615
R432 source.n943 source.n875 104.615
R433 source.n944 source.n943 104.615
R434 source.n944 source.n871 104.615
R435 source.n951 source.n871 104.615
R436 source.n952 source.n951 104.615
R437 source.n952 source.n867 104.615
R438 source.n959 source.n867 104.615
R439 source.n961 source.n959 104.615
R440 source.n961 source.n960 104.615
R441 source.n960 source.n863 104.615
R442 source.n969 source.n863 104.615
R443 source.n970 source.n969 104.615
R444 source.n970 source.n859 104.615
R445 source.n977 source.n859 104.615
R446 source.n978 source.n977 104.615
R447 source.n978 source.n855 104.615
R448 source.n985 source.n855 104.615
R449 source.n986 source.n985 104.615
R450 source.n761 source.n755 104.615
R451 source.n762 source.n761 104.615
R452 source.n762 source.n751 104.615
R453 source.n769 source.n751 104.615
R454 source.n770 source.n769 104.615
R455 source.n770 source.n747 104.615
R456 source.n778 source.n747 104.615
R457 source.n779 source.n778 104.615
R458 source.n780 source.n779 104.615
R459 source.n780 source.n743 104.615
R460 source.n787 source.n743 104.615
R461 source.n788 source.n787 104.615
R462 source.n788 source.n739 104.615
R463 source.n795 source.n739 104.615
R464 source.n796 source.n795 104.615
R465 source.n796 source.n735 104.615
R466 source.n803 source.n735 104.615
R467 source.n804 source.n803 104.615
R468 source.n804 source.n731 104.615
R469 source.n811 source.n731 104.615
R470 source.n812 source.n811 104.615
R471 source.n812 source.n727 104.615
R472 source.n819 source.n727 104.615
R473 source.n821 source.n819 104.615
R474 source.n821 source.n820 104.615
R475 source.n820 source.n723 104.615
R476 source.n829 source.n723 104.615
R477 source.n830 source.n829 104.615
R478 source.n830 source.n719 104.615
R479 source.n837 source.n719 104.615
R480 source.n838 source.n837 104.615
R481 source.n838 source.n715 104.615
R482 source.n845 source.n715 104.615
R483 source.n846 source.n845 104.615
R484 source.n617 source.n611 104.615
R485 source.n618 source.n617 104.615
R486 source.n618 source.n607 104.615
R487 source.n625 source.n607 104.615
R488 source.n626 source.n625 104.615
R489 source.n626 source.n603 104.615
R490 source.n634 source.n603 104.615
R491 source.n635 source.n634 104.615
R492 source.n636 source.n635 104.615
R493 source.n636 source.n599 104.615
R494 source.n643 source.n599 104.615
R495 source.n644 source.n643 104.615
R496 source.n644 source.n595 104.615
R497 source.n651 source.n595 104.615
R498 source.n652 source.n651 104.615
R499 source.n652 source.n591 104.615
R500 source.n659 source.n591 104.615
R501 source.n660 source.n659 104.615
R502 source.n660 source.n587 104.615
R503 source.n667 source.n587 104.615
R504 source.n668 source.n667 104.615
R505 source.n668 source.n583 104.615
R506 source.n675 source.n583 104.615
R507 source.n677 source.n675 104.615
R508 source.n677 source.n676 104.615
R509 source.n676 source.n579 104.615
R510 source.n685 source.n579 104.615
R511 source.n686 source.n685 104.615
R512 source.n686 source.n575 104.615
R513 source.n693 source.n575 104.615
R514 source.n694 source.n693 104.615
R515 source.n694 source.n571 104.615
R516 source.n701 source.n571 104.615
R517 source.n702 source.n701 104.615
R518 source.n134 source.n133 104.615
R519 source.n133 source.n3 104.615
R520 source.n126 source.n3 104.615
R521 source.n126 source.n125 104.615
R522 source.n125 source.n7 104.615
R523 source.n118 source.n7 104.615
R524 source.n118 source.n117 104.615
R525 source.n117 source.n11 104.615
R526 source.n15 source.n11 104.615
R527 source.n109 source.n15 104.615
R528 source.n109 source.n108 104.615
R529 source.n108 source.n16 104.615
R530 source.n101 source.n16 104.615
R531 source.n101 source.n100 104.615
R532 source.n100 source.n20 104.615
R533 source.n93 source.n20 104.615
R534 source.n93 source.n92 104.615
R535 source.n92 source.n24 104.615
R536 source.n85 source.n24 104.615
R537 source.n85 source.n84 104.615
R538 source.n84 source.n28 104.615
R539 source.n77 source.n28 104.615
R540 source.n77 source.n76 104.615
R541 source.n76 source.n32 104.615
R542 source.n69 source.n32 104.615
R543 source.n69 source.n68 104.615
R544 source.n68 source.n67 104.615
R545 source.n67 source.n36 104.615
R546 source.n60 source.n36 104.615
R547 source.n60 source.n59 104.615
R548 source.n59 source.n41 104.615
R549 source.n52 source.n41 104.615
R550 source.n52 source.n51 104.615
R551 source.n51 source.n45 104.615
R552 source.n278 source.n277 104.615
R553 source.n277 source.n147 104.615
R554 source.n270 source.n147 104.615
R555 source.n270 source.n269 104.615
R556 source.n269 source.n151 104.615
R557 source.n262 source.n151 104.615
R558 source.n262 source.n261 104.615
R559 source.n261 source.n155 104.615
R560 source.n159 source.n155 104.615
R561 source.n253 source.n159 104.615
R562 source.n253 source.n252 104.615
R563 source.n252 source.n160 104.615
R564 source.n245 source.n160 104.615
R565 source.n245 source.n244 104.615
R566 source.n244 source.n164 104.615
R567 source.n237 source.n164 104.615
R568 source.n237 source.n236 104.615
R569 source.n236 source.n168 104.615
R570 source.n229 source.n168 104.615
R571 source.n229 source.n228 104.615
R572 source.n228 source.n172 104.615
R573 source.n221 source.n172 104.615
R574 source.n221 source.n220 104.615
R575 source.n220 source.n176 104.615
R576 source.n213 source.n176 104.615
R577 source.n213 source.n212 104.615
R578 source.n212 source.n211 104.615
R579 source.n211 source.n180 104.615
R580 source.n204 source.n180 104.615
R581 source.n204 source.n203 104.615
R582 source.n203 source.n185 104.615
R583 source.n196 source.n185 104.615
R584 source.n196 source.n195 104.615
R585 source.n195 source.n189 104.615
R586 source.n418 source.n417 104.615
R587 source.n417 source.n287 104.615
R588 source.n410 source.n287 104.615
R589 source.n410 source.n409 104.615
R590 source.n409 source.n291 104.615
R591 source.n402 source.n291 104.615
R592 source.n402 source.n401 104.615
R593 source.n401 source.n295 104.615
R594 source.n299 source.n295 104.615
R595 source.n393 source.n299 104.615
R596 source.n393 source.n392 104.615
R597 source.n392 source.n300 104.615
R598 source.n385 source.n300 104.615
R599 source.n385 source.n384 104.615
R600 source.n384 source.n304 104.615
R601 source.n377 source.n304 104.615
R602 source.n377 source.n376 104.615
R603 source.n376 source.n308 104.615
R604 source.n369 source.n308 104.615
R605 source.n369 source.n368 104.615
R606 source.n368 source.n312 104.615
R607 source.n361 source.n312 104.615
R608 source.n361 source.n360 104.615
R609 source.n360 source.n316 104.615
R610 source.n353 source.n316 104.615
R611 source.n353 source.n352 104.615
R612 source.n352 source.n351 104.615
R613 source.n351 source.n320 104.615
R614 source.n344 source.n320 104.615
R615 source.n344 source.n343 104.615
R616 source.n343 source.n325 104.615
R617 source.n336 source.n325 104.615
R618 source.n336 source.n335 104.615
R619 source.n335 source.n329 104.615
R620 source.n562 source.n561 104.615
R621 source.n561 source.n431 104.615
R622 source.n554 source.n431 104.615
R623 source.n554 source.n553 104.615
R624 source.n553 source.n435 104.615
R625 source.n546 source.n435 104.615
R626 source.n546 source.n545 104.615
R627 source.n545 source.n439 104.615
R628 source.n443 source.n439 104.615
R629 source.n537 source.n443 104.615
R630 source.n537 source.n536 104.615
R631 source.n536 source.n444 104.615
R632 source.n529 source.n444 104.615
R633 source.n529 source.n528 104.615
R634 source.n528 source.n448 104.615
R635 source.n521 source.n448 104.615
R636 source.n521 source.n520 104.615
R637 source.n520 source.n452 104.615
R638 source.n513 source.n452 104.615
R639 source.n513 source.n512 104.615
R640 source.n512 source.n456 104.615
R641 source.n505 source.n456 104.615
R642 source.n505 source.n504 104.615
R643 source.n504 source.n460 104.615
R644 source.n497 source.n460 104.615
R645 source.n497 source.n496 104.615
R646 source.n496 source.n495 104.615
R647 source.n495 source.n464 104.615
R648 source.n488 source.n464 104.615
R649 source.n488 source.n487 104.615
R650 source.n487 source.n469 104.615
R651 source.n480 source.n469 104.615
R652 source.n480 source.n479 104.615
R653 source.n479 source.n473 104.615
R654 source.t11 source.n1039 52.3082
R655 source.t15 source.n895 52.3082
R656 source.t6 source.n755 52.3082
R657 source.t2 source.n611 52.3082
R658 source.t0 source.n45 52.3082
R659 source.t7 source.n189 52.3082
R660 source.t12 source.n329 52.3082
R661 source.t9 source.n473 52.3082
R662 source.n995 source.n994 42.0366
R663 source.n993 source.n992 42.0366
R664 source.n711 source.n710 42.0366
R665 source.n709 source.n708 42.0366
R666 source.n141 source.n140 42.0366
R667 source.n143 source.n142 42.0366
R668 source.n425 source.n424 42.0366
R669 source.n427 source.n426 42.0366
R670 source.n707 source.n567 32.0241
R671 source.n1135 source.n1134 30.6338
R672 source.n991 source.n990 30.6338
R673 source.n851 source.n850 30.6338
R674 source.n707 source.n706 30.6338
R675 source.n139 source.n138 30.6338
R676 source.n283 source.n282 30.6338
R677 source.n423 source.n422 30.6338
R678 source.n567 source.n566 30.6338
R679 source.n1136 source.n139 26.3172
R680 source.n1065 source.n1030 13.1884
R681 source.n1112 source.n1111 13.1884
R682 source.n921 source.n886 13.1884
R683 source.n968 source.n967 13.1884
R684 source.n781 source.n746 13.1884
R685 source.n828 source.n827 13.1884
R686 source.n637 source.n602 13.1884
R687 source.n684 source.n683 13.1884
R688 source.n116 source.n115 13.1884
R689 source.n70 source.n35 13.1884
R690 source.n260 source.n259 13.1884
R691 source.n214 source.n179 13.1884
R692 source.n400 source.n399 13.1884
R693 source.n354 source.n319 13.1884
R694 source.n544 source.n543 13.1884
R695 source.n498 source.n463 13.1884
R696 source.n1061 source.n1060 12.8005
R697 source.n1066 source.n1028 12.8005
R698 source.n1110 source.n1008 12.8005
R699 source.n1115 source.n1006 12.8005
R700 source.n917 source.n916 12.8005
R701 source.n922 source.n884 12.8005
R702 source.n966 source.n864 12.8005
R703 source.n971 source.n862 12.8005
R704 source.n777 source.n776 12.8005
R705 source.n782 source.n744 12.8005
R706 source.n826 source.n724 12.8005
R707 source.n831 source.n722 12.8005
R708 source.n633 source.n632 12.8005
R709 source.n638 source.n600 12.8005
R710 source.n682 source.n580 12.8005
R711 source.n687 source.n578 12.8005
R712 source.n119 source.n10 12.8005
R713 source.n114 source.n12 12.8005
R714 source.n71 source.n33 12.8005
R715 source.n66 source.n37 12.8005
R716 source.n263 source.n154 12.8005
R717 source.n258 source.n156 12.8005
R718 source.n215 source.n177 12.8005
R719 source.n210 source.n181 12.8005
R720 source.n403 source.n294 12.8005
R721 source.n398 source.n296 12.8005
R722 source.n355 source.n317 12.8005
R723 source.n350 source.n321 12.8005
R724 source.n547 source.n438 12.8005
R725 source.n542 source.n440 12.8005
R726 source.n499 source.n461 12.8005
R727 source.n494 source.n465 12.8005
R728 source.n1059 source.n1032 12.0247
R729 source.n1070 source.n1069 12.0247
R730 source.n1107 source.n1106 12.0247
R731 source.n1116 source.n1004 12.0247
R732 source.n915 source.n888 12.0247
R733 source.n926 source.n925 12.0247
R734 source.n963 source.n962 12.0247
R735 source.n972 source.n860 12.0247
R736 source.n775 source.n748 12.0247
R737 source.n786 source.n785 12.0247
R738 source.n823 source.n822 12.0247
R739 source.n832 source.n720 12.0247
R740 source.n631 source.n604 12.0247
R741 source.n642 source.n641 12.0247
R742 source.n679 source.n678 12.0247
R743 source.n688 source.n576 12.0247
R744 source.n120 source.n8 12.0247
R745 source.n111 source.n110 12.0247
R746 source.n75 source.n74 12.0247
R747 source.n65 source.n38 12.0247
R748 source.n264 source.n152 12.0247
R749 source.n255 source.n254 12.0247
R750 source.n219 source.n218 12.0247
R751 source.n209 source.n182 12.0247
R752 source.n404 source.n292 12.0247
R753 source.n395 source.n394 12.0247
R754 source.n359 source.n358 12.0247
R755 source.n349 source.n322 12.0247
R756 source.n548 source.n436 12.0247
R757 source.n539 source.n538 12.0247
R758 source.n503 source.n502 12.0247
R759 source.n493 source.n466 12.0247
R760 source.n1056 source.n1055 11.249
R761 source.n1073 source.n1026 11.249
R762 source.n1102 source.n1010 11.249
R763 source.n1120 source.n1119 11.249
R764 source.n912 source.n911 11.249
R765 source.n929 source.n882 11.249
R766 source.n958 source.n866 11.249
R767 source.n976 source.n975 11.249
R768 source.n772 source.n771 11.249
R769 source.n789 source.n742 11.249
R770 source.n818 source.n726 11.249
R771 source.n836 source.n835 11.249
R772 source.n628 source.n627 11.249
R773 source.n645 source.n598 11.249
R774 source.n674 source.n582 11.249
R775 source.n692 source.n691 11.249
R776 source.n124 source.n123 11.249
R777 source.n107 source.n14 11.249
R778 source.n78 source.n31 11.249
R779 source.n62 source.n61 11.249
R780 source.n268 source.n267 11.249
R781 source.n251 source.n158 11.249
R782 source.n222 source.n175 11.249
R783 source.n206 source.n205 11.249
R784 source.n408 source.n407 11.249
R785 source.n391 source.n298 11.249
R786 source.n362 source.n315 11.249
R787 source.n346 source.n345 11.249
R788 source.n552 source.n551 11.249
R789 source.n535 source.n442 11.249
R790 source.n506 source.n459 11.249
R791 source.n490 source.n489 11.249
R792 source.n1052 source.n1034 10.4732
R793 source.n1074 source.n1024 10.4732
R794 source.n1101 source.n1012 10.4732
R795 source.n1123 source.n1002 10.4732
R796 source.n908 source.n890 10.4732
R797 source.n930 source.n880 10.4732
R798 source.n957 source.n868 10.4732
R799 source.n979 source.n858 10.4732
R800 source.n768 source.n750 10.4732
R801 source.n790 source.n740 10.4732
R802 source.n817 source.n728 10.4732
R803 source.n839 source.n718 10.4732
R804 source.n624 source.n606 10.4732
R805 source.n646 source.n596 10.4732
R806 source.n673 source.n584 10.4732
R807 source.n695 source.n574 10.4732
R808 source.n127 source.n6 10.4732
R809 source.n106 source.n17 10.4732
R810 source.n79 source.n29 10.4732
R811 source.n58 source.n40 10.4732
R812 source.n271 source.n150 10.4732
R813 source.n250 source.n161 10.4732
R814 source.n223 source.n173 10.4732
R815 source.n202 source.n184 10.4732
R816 source.n411 source.n290 10.4732
R817 source.n390 source.n301 10.4732
R818 source.n363 source.n313 10.4732
R819 source.n342 source.n324 10.4732
R820 source.n555 source.n434 10.4732
R821 source.n534 source.n445 10.4732
R822 source.n507 source.n457 10.4732
R823 source.n486 source.n468 10.4732
R824 source.n1041 source.n1040 10.2747
R825 source.n897 source.n896 10.2747
R826 source.n757 source.n756 10.2747
R827 source.n613 source.n612 10.2747
R828 source.n47 source.n46 10.2747
R829 source.n191 source.n190 10.2747
R830 source.n331 source.n330 10.2747
R831 source.n475 source.n474 10.2747
R832 source.n1051 source.n1036 9.69747
R833 source.n1078 source.n1077 9.69747
R834 source.n1098 source.n1097 9.69747
R835 source.n1124 source.n1000 9.69747
R836 source.n907 source.n892 9.69747
R837 source.n934 source.n933 9.69747
R838 source.n954 source.n953 9.69747
R839 source.n980 source.n856 9.69747
R840 source.n767 source.n752 9.69747
R841 source.n794 source.n793 9.69747
R842 source.n814 source.n813 9.69747
R843 source.n840 source.n716 9.69747
R844 source.n623 source.n608 9.69747
R845 source.n650 source.n649 9.69747
R846 source.n670 source.n669 9.69747
R847 source.n696 source.n572 9.69747
R848 source.n128 source.n4 9.69747
R849 source.n103 source.n102 9.69747
R850 source.n83 source.n82 9.69747
R851 source.n57 source.n42 9.69747
R852 source.n272 source.n148 9.69747
R853 source.n247 source.n246 9.69747
R854 source.n227 source.n226 9.69747
R855 source.n201 source.n186 9.69747
R856 source.n412 source.n288 9.69747
R857 source.n387 source.n386 9.69747
R858 source.n367 source.n366 9.69747
R859 source.n341 source.n326 9.69747
R860 source.n556 source.n432 9.69747
R861 source.n531 source.n530 9.69747
R862 source.n511 source.n510 9.69747
R863 source.n485 source.n470 9.69747
R864 source.n1134 source.n1133 9.45567
R865 source.n990 source.n989 9.45567
R866 source.n850 source.n849 9.45567
R867 source.n706 source.n705 9.45567
R868 source.n138 source.n137 9.45567
R869 source.n282 source.n281 9.45567
R870 source.n422 source.n421 9.45567
R871 source.n566 source.n565 9.45567
R872 source.n998 source.n997 9.3005
R873 source.n1127 source.n1126 9.3005
R874 source.n1125 source.n1124 9.3005
R875 source.n1002 source.n1001 9.3005
R876 source.n1119 source.n1118 9.3005
R877 source.n1117 source.n1116 9.3005
R878 source.n1006 source.n1005 9.3005
R879 source.n1085 source.n1084 9.3005
R880 source.n1083 source.n1082 9.3005
R881 source.n1022 source.n1021 9.3005
R882 source.n1077 source.n1076 9.3005
R883 source.n1075 source.n1074 9.3005
R884 source.n1026 source.n1025 9.3005
R885 source.n1069 source.n1068 9.3005
R886 source.n1067 source.n1066 9.3005
R887 source.n1043 source.n1042 9.3005
R888 source.n1038 source.n1037 9.3005
R889 source.n1049 source.n1048 9.3005
R890 source.n1051 source.n1050 9.3005
R891 source.n1034 source.n1033 9.3005
R892 source.n1057 source.n1056 9.3005
R893 source.n1059 source.n1058 9.3005
R894 source.n1060 source.n1029 9.3005
R895 source.n1018 source.n1017 9.3005
R896 source.n1091 source.n1090 9.3005
R897 source.n1093 source.n1092 9.3005
R898 source.n1014 source.n1013 9.3005
R899 source.n1099 source.n1098 9.3005
R900 source.n1101 source.n1100 9.3005
R901 source.n1010 source.n1009 9.3005
R902 source.n1108 source.n1107 9.3005
R903 source.n1110 source.n1109 9.3005
R904 source.n1133 source.n1132 9.3005
R905 source.n854 source.n853 9.3005
R906 source.n983 source.n982 9.3005
R907 source.n981 source.n980 9.3005
R908 source.n858 source.n857 9.3005
R909 source.n975 source.n974 9.3005
R910 source.n973 source.n972 9.3005
R911 source.n862 source.n861 9.3005
R912 source.n941 source.n940 9.3005
R913 source.n939 source.n938 9.3005
R914 source.n878 source.n877 9.3005
R915 source.n933 source.n932 9.3005
R916 source.n931 source.n930 9.3005
R917 source.n882 source.n881 9.3005
R918 source.n925 source.n924 9.3005
R919 source.n923 source.n922 9.3005
R920 source.n899 source.n898 9.3005
R921 source.n894 source.n893 9.3005
R922 source.n905 source.n904 9.3005
R923 source.n907 source.n906 9.3005
R924 source.n890 source.n889 9.3005
R925 source.n913 source.n912 9.3005
R926 source.n915 source.n914 9.3005
R927 source.n916 source.n885 9.3005
R928 source.n874 source.n873 9.3005
R929 source.n947 source.n946 9.3005
R930 source.n949 source.n948 9.3005
R931 source.n870 source.n869 9.3005
R932 source.n955 source.n954 9.3005
R933 source.n957 source.n956 9.3005
R934 source.n866 source.n865 9.3005
R935 source.n964 source.n963 9.3005
R936 source.n966 source.n965 9.3005
R937 source.n989 source.n988 9.3005
R938 source.n714 source.n713 9.3005
R939 source.n843 source.n842 9.3005
R940 source.n841 source.n840 9.3005
R941 source.n718 source.n717 9.3005
R942 source.n835 source.n834 9.3005
R943 source.n833 source.n832 9.3005
R944 source.n722 source.n721 9.3005
R945 source.n801 source.n800 9.3005
R946 source.n799 source.n798 9.3005
R947 source.n738 source.n737 9.3005
R948 source.n793 source.n792 9.3005
R949 source.n791 source.n790 9.3005
R950 source.n742 source.n741 9.3005
R951 source.n785 source.n784 9.3005
R952 source.n783 source.n782 9.3005
R953 source.n759 source.n758 9.3005
R954 source.n754 source.n753 9.3005
R955 source.n765 source.n764 9.3005
R956 source.n767 source.n766 9.3005
R957 source.n750 source.n749 9.3005
R958 source.n773 source.n772 9.3005
R959 source.n775 source.n774 9.3005
R960 source.n776 source.n745 9.3005
R961 source.n734 source.n733 9.3005
R962 source.n807 source.n806 9.3005
R963 source.n809 source.n808 9.3005
R964 source.n730 source.n729 9.3005
R965 source.n815 source.n814 9.3005
R966 source.n817 source.n816 9.3005
R967 source.n726 source.n725 9.3005
R968 source.n824 source.n823 9.3005
R969 source.n826 source.n825 9.3005
R970 source.n849 source.n848 9.3005
R971 source.n570 source.n569 9.3005
R972 source.n699 source.n698 9.3005
R973 source.n697 source.n696 9.3005
R974 source.n574 source.n573 9.3005
R975 source.n691 source.n690 9.3005
R976 source.n689 source.n688 9.3005
R977 source.n578 source.n577 9.3005
R978 source.n657 source.n656 9.3005
R979 source.n655 source.n654 9.3005
R980 source.n594 source.n593 9.3005
R981 source.n649 source.n648 9.3005
R982 source.n647 source.n646 9.3005
R983 source.n598 source.n597 9.3005
R984 source.n641 source.n640 9.3005
R985 source.n639 source.n638 9.3005
R986 source.n615 source.n614 9.3005
R987 source.n610 source.n609 9.3005
R988 source.n621 source.n620 9.3005
R989 source.n623 source.n622 9.3005
R990 source.n606 source.n605 9.3005
R991 source.n629 source.n628 9.3005
R992 source.n631 source.n630 9.3005
R993 source.n632 source.n601 9.3005
R994 source.n590 source.n589 9.3005
R995 source.n663 source.n662 9.3005
R996 source.n665 source.n664 9.3005
R997 source.n586 source.n585 9.3005
R998 source.n671 source.n670 9.3005
R999 source.n673 source.n672 9.3005
R1000 source.n582 source.n581 9.3005
R1001 source.n680 source.n679 9.3005
R1002 source.n682 source.n681 9.3005
R1003 source.n705 source.n704 9.3005
R1004 source.n49 source.n48 9.3005
R1005 source.n44 source.n43 9.3005
R1006 source.n55 source.n54 9.3005
R1007 source.n57 source.n56 9.3005
R1008 source.n40 source.n39 9.3005
R1009 source.n63 source.n62 9.3005
R1010 source.n65 source.n64 9.3005
R1011 source.n37 source.n34 9.3005
R1012 source.n96 source.n95 9.3005
R1013 source.n98 source.n97 9.3005
R1014 source.n19 source.n18 9.3005
R1015 source.n104 source.n103 9.3005
R1016 source.n106 source.n105 9.3005
R1017 source.n14 source.n13 9.3005
R1018 source.n112 source.n111 9.3005
R1019 source.n114 source.n113 9.3005
R1020 source.n137 source.n136 9.3005
R1021 source.n2 source.n1 9.3005
R1022 source.n131 source.n130 9.3005
R1023 source.n129 source.n128 9.3005
R1024 source.n6 source.n5 9.3005
R1025 source.n123 source.n122 9.3005
R1026 source.n121 source.n120 9.3005
R1027 source.n10 source.n9 9.3005
R1028 source.n23 source.n22 9.3005
R1029 source.n90 source.n89 9.3005
R1030 source.n88 source.n87 9.3005
R1031 source.n27 source.n26 9.3005
R1032 source.n82 source.n81 9.3005
R1033 source.n80 source.n79 9.3005
R1034 source.n31 source.n30 9.3005
R1035 source.n74 source.n73 9.3005
R1036 source.n72 source.n71 9.3005
R1037 source.n193 source.n192 9.3005
R1038 source.n188 source.n187 9.3005
R1039 source.n199 source.n198 9.3005
R1040 source.n201 source.n200 9.3005
R1041 source.n184 source.n183 9.3005
R1042 source.n207 source.n206 9.3005
R1043 source.n209 source.n208 9.3005
R1044 source.n181 source.n178 9.3005
R1045 source.n240 source.n239 9.3005
R1046 source.n242 source.n241 9.3005
R1047 source.n163 source.n162 9.3005
R1048 source.n248 source.n247 9.3005
R1049 source.n250 source.n249 9.3005
R1050 source.n158 source.n157 9.3005
R1051 source.n256 source.n255 9.3005
R1052 source.n258 source.n257 9.3005
R1053 source.n281 source.n280 9.3005
R1054 source.n146 source.n145 9.3005
R1055 source.n275 source.n274 9.3005
R1056 source.n273 source.n272 9.3005
R1057 source.n150 source.n149 9.3005
R1058 source.n267 source.n266 9.3005
R1059 source.n265 source.n264 9.3005
R1060 source.n154 source.n153 9.3005
R1061 source.n167 source.n166 9.3005
R1062 source.n234 source.n233 9.3005
R1063 source.n232 source.n231 9.3005
R1064 source.n171 source.n170 9.3005
R1065 source.n226 source.n225 9.3005
R1066 source.n224 source.n223 9.3005
R1067 source.n175 source.n174 9.3005
R1068 source.n218 source.n217 9.3005
R1069 source.n216 source.n215 9.3005
R1070 source.n333 source.n332 9.3005
R1071 source.n328 source.n327 9.3005
R1072 source.n339 source.n338 9.3005
R1073 source.n341 source.n340 9.3005
R1074 source.n324 source.n323 9.3005
R1075 source.n347 source.n346 9.3005
R1076 source.n349 source.n348 9.3005
R1077 source.n321 source.n318 9.3005
R1078 source.n380 source.n379 9.3005
R1079 source.n382 source.n381 9.3005
R1080 source.n303 source.n302 9.3005
R1081 source.n388 source.n387 9.3005
R1082 source.n390 source.n389 9.3005
R1083 source.n298 source.n297 9.3005
R1084 source.n396 source.n395 9.3005
R1085 source.n398 source.n397 9.3005
R1086 source.n421 source.n420 9.3005
R1087 source.n286 source.n285 9.3005
R1088 source.n415 source.n414 9.3005
R1089 source.n413 source.n412 9.3005
R1090 source.n290 source.n289 9.3005
R1091 source.n407 source.n406 9.3005
R1092 source.n405 source.n404 9.3005
R1093 source.n294 source.n293 9.3005
R1094 source.n307 source.n306 9.3005
R1095 source.n374 source.n373 9.3005
R1096 source.n372 source.n371 9.3005
R1097 source.n311 source.n310 9.3005
R1098 source.n366 source.n365 9.3005
R1099 source.n364 source.n363 9.3005
R1100 source.n315 source.n314 9.3005
R1101 source.n358 source.n357 9.3005
R1102 source.n356 source.n355 9.3005
R1103 source.n477 source.n476 9.3005
R1104 source.n472 source.n471 9.3005
R1105 source.n483 source.n482 9.3005
R1106 source.n485 source.n484 9.3005
R1107 source.n468 source.n467 9.3005
R1108 source.n491 source.n490 9.3005
R1109 source.n493 source.n492 9.3005
R1110 source.n465 source.n462 9.3005
R1111 source.n524 source.n523 9.3005
R1112 source.n526 source.n525 9.3005
R1113 source.n447 source.n446 9.3005
R1114 source.n532 source.n531 9.3005
R1115 source.n534 source.n533 9.3005
R1116 source.n442 source.n441 9.3005
R1117 source.n540 source.n539 9.3005
R1118 source.n542 source.n541 9.3005
R1119 source.n565 source.n564 9.3005
R1120 source.n430 source.n429 9.3005
R1121 source.n559 source.n558 9.3005
R1122 source.n557 source.n556 9.3005
R1123 source.n434 source.n433 9.3005
R1124 source.n551 source.n550 9.3005
R1125 source.n549 source.n548 9.3005
R1126 source.n438 source.n437 9.3005
R1127 source.n451 source.n450 9.3005
R1128 source.n518 source.n517 9.3005
R1129 source.n516 source.n515 9.3005
R1130 source.n455 source.n454 9.3005
R1131 source.n510 source.n509 9.3005
R1132 source.n508 source.n507 9.3005
R1133 source.n459 source.n458 9.3005
R1134 source.n502 source.n501 9.3005
R1135 source.n500 source.n499 9.3005
R1136 source.n1048 source.n1047 8.92171
R1137 source.n1081 source.n1022 8.92171
R1138 source.n1094 source.n1014 8.92171
R1139 source.n1128 source.n1127 8.92171
R1140 source.n904 source.n903 8.92171
R1141 source.n937 source.n878 8.92171
R1142 source.n950 source.n870 8.92171
R1143 source.n984 source.n983 8.92171
R1144 source.n764 source.n763 8.92171
R1145 source.n797 source.n738 8.92171
R1146 source.n810 source.n730 8.92171
R1147 source.n844 source.n843 8.92171
R1148 source.n620 source.n619 8.92171
R1149 source.n653 source.n594 8.92171
R1150 source.n666 source.n586 8.92171
R1151 source.n700 source.n699 8.92171
R1152 source.n132 source.n131 8.92171
R1153 source.n99 source.n19 8.92171
R1154 source.n86 source.n27 8.92171
R1155 source.n54 source.n53 8.92171
R1156 source.n276 source.n275 8.92171
R1157 source.n243 source.n163 8.92171
R1158 source.n230 source.n171 8.92171
R1159 source.n198 source.n197 8.92171
R1160 source.n416 source.n415 8.92171
R1161 source.n383 source.n303 8.92171
R1162 source.n370 source.n311 8.92171
R1163 source.n338 source.n337 8.92171
R1164 source.n560 source.n559 8.92171
R1165 source.n527 source.n447 8.92171
R1166 source.n514 source.n455 8.92171
R1167 source.n482 source.n481 8.92171
R1168 source.n1044 source.n1038 8.14595
R1169 source.n1082 source.n1020 8.14595
R1170 source.n1093 source.n1016 8.14595
R1171 source.n1131 source.n998 8.14595
R1172 source.n900 source.n894 8.14595
R1173 source.n938 source.n876 8.14595
R1174 source.n949 source.n872 8.14595
R1175 source.n987 source.n854 8.14595
R1176 source.n760 source.n754 8.14595
R1177 source.n798 source.n736 8.14595
R1178 source.n809 source.n732 8.14595
R1179 source.n847 source.n714 8.14595
R1180 source.n616 source.n610 8.14595
R1181 source.n654 source.n592 8.14595
R1182 source.n665 source.n588 8.14595
R1183 source.n703 source.n570 8.14595
R1184 source.n135 source.n2 8.14595
R1185 source.n98 source.n21 8.14595
R1186 source.n87 source.n25 8.14595
R1187 source.n50 source.n44 8.14595
R1188 source.n279 source.n146 8.14595
R1189 source.n242 source.n165 8.14595
R1190 source.n231 source.n169 8.14595
R1191 source.n194 source.n188 8.14595
R1192 source.n419 source.n286 8.14595
R1193 source.n382 source.n305 8.14595
R1194 source.n371 source.n309 8.14595
R1195 source.n334 source.n328 8.14595
R1196 source.n563 source.n430 8.14595
R1197 source.n526 source.n449 8.14595
R1198 source.n515 source.n453 8.14595
R1199 source.n478 source.n472 8.14595
R1200 source.n1043 source.n1040 7.3702
R1201 source.n1086 source.n1085 7.3702
R1202 source.n1090 source.n1089 7.3702
R1203 source.n1132 source.n996 7.3702
R1204 source.n899 source.n896 7.3702
R1205 source.n942 source.n941 7.3702
R1206 source.n946 source.n945 7.3702
R1207 source.n988 source.n852 7.3702
R1208 source.n759 source.n756 7.3702
R1209 source.n802 source.n801 7.3702
R1210 source.n806 source.n805 7.3702
R1211 source.n848 source.n712 7.3702
R1212 source.n615 source.n612 7.3702
R1213 source.n658 source.n657 7.3702
R1214 source.n662 source.n661 7.3702
R1215 source.n704 source.n568 7.3702
R1216 source.n136 source.n0 7.3702
R1217 source.n95 source.n94 7.3702
R1218 source.n91 source.n90 7.3702
R1219 source.n49 source.n46 7.3702
R1220 source.n280 source.n144 7.3702
R1221 source.n239 source.n238 7.3702
R1222 source.n235 source.n234 7.3702
R1223 source.n193 source.n190 7.3702
R1224 source.n420 source.n284 7.3702
R1225 source.n379 source.n378 7.3702
R1226 source.n375 source.n374 7.3702
R1227 source.n333 source.n330 7.3702
R1228 source.n564 source.n428 7.3702
R1229 source.n523 source.n522 7.3702
R1230 source.n519 source.n518 7.3702
R1231 source.n477 source.n474 7.3702
R1232 source.n1086 source.n1018 6.59444
R1233 source.n1089 source.n1018 6.59444
R1234 source.n1134 source.n996 6.59444
R1235 source.n942 source.n874 6.59444
R1236 source.n945 source.n874 6.59444
R1237 source.n990 source.n852 6.59444
R1238 source.n802 source.n734 6.59444
R1239 source.n805 source.n734 6.59444
R1240 source.n850 source.n712 6.59444
R1241 source.n658 source.n590 6.59444
R1242 source.n661 source.n590 6.59444
R1243 source.n706 source.n568 6.59444
R1244 source.n138 source.n0 6.59444
R1245 source.n94 source.n23 6.59444
R1246 source.n91 source.n23 6.59444
R1247 source.n282 source.n144 6.59444
R1248 source.n238 source.n167 6.59444
R1249 source.n235 source.n167 6.59444
R1250 source.n422 source.n284 6.59444
R1251 source.n378 source.n307 6.59444
R1252 source.n375 source.n307 6.59444
R1253 source.n566 source.n428 6.59444
R1254 source.n522 source.n451 6.59444
R1255 source.n519 source.n451 6.59444
R1256 source.n1044 source.n1043 5.81868
R1257 source.n1085 source.n1020 5.81868
R1258 source.n1090 source.n1016 5.81868
R1259 source.n1132 source.n1131 5.81868
R1260 source.n900 source.n899 5.81868
R1261 source.n941 source.n876 5.81868
R1262 source.n946 source.n872 5.81868
R1263 source.n988 source.n987 5.81868
R1264 source.n760 source.n759 5.81868
R1265 source.n801 source.n736 5.81868
R1266 source.n806 source.n732 5.81868
R1267 source.n848 source.n847 5.81868
R1268 source.n616 source.n615 5.81868
R1269 source.n657 source.n592 5.81868
R1270 source.n662 source.n588 5.81868
R1271 source.n704 source.n703 5.81868
R1272 source.n136 source.n135 5.81868
R1273 source.n95 source.n21 5.81868
R1274 source.n90 source.n25 5.81868
R1275 source.n50 source.n49 5.81868
R1276 source.n280 source.n279 5.81868
R1277 source.n239 source.n165 5.81868
R1278 source.n234 source.n169 5.81868
R1279 source.n194 source.n193 5.81868
R1280 source.n420 source.n419 5.81868
R1281 source.n379 source.n305 5.81868
R1282 source.n374 source.n309 5.81868
R1283 source.n334 source.n333 5.81868
R1284 source.n564 source.n563 5.81868
R1285 source.n523 source.n449 5.81868
R1286 source.n518 source.n453 5.81868
R1287 source.n478 source.n477 5.81868
R1288 source.n1136 source.n1135 5.7074
R1289 source.n1047 source.n1038 5.04292
R1290 source.n1082 source.n1081 5.04292
R1291 source.n1094 source.n1093 5.04292
R1292 source.n1128 source.n998 5.04292
R1293 source.n903 source.n894 5.04292
R1294 source.n938 source.n937 5.04292
R1295 source.n950 source.n949 5.04292
R1296 source.n984 source.n854 5.04292
R1297 source.n763 source.n754 5.04292
R1298 source.n798 source.n797 5.04292
R1299 source.n810 source.n809 5.04292
R1300 source.n844 source.n714 5.04292
R1301 source.n619 source.n610 5.04292
R1302 source.n654 source.n653 5.04292
R1303 source.n666 source.n665 5.04292
R1304 source.n700 source.n570 5.04292
R1305 source.n132 source.n2 5.04292
R1306 source.n99 source.n98 5.04292
R1307 source.n87 source.n86 5.04292
R1308 source.n53 source.n44 5.04292
R1309 source.n276 source.n146 5.04292
R1310 source.n243 source.n242 5.04292
R1311 source.n231 source.n230 5.04292
R1312 source.n197 source.n188 5.04292
R1313 source.n416 source.n286 5.04292
R1314 source.n383 source.n382 5.04292
R1315 source.n371 source.n370 5.04292
R1316 source.n337 source.n328 5.04292
R1317 source.n560 source.n430 5.04292
R1318 source.n527 source.n526 5.04292
R1319 source.n515 source.n514 5.04292
R1320 source.n481 source.n472 5.04292
R1321 source.n1048 source.n1036 4.26717
R1322 source.n1078 source.n1022 4.26717
R1323 source.n1097 source.n1014 4.26717
R1324 source.n1127 source.n1000 4.26717
R1325 source.n904 source.n892 4.26717
R1326 source.n934 source.n878 4.26717
R1327 source.n953 source.n870 4.26717
R1328 source.n983 source.n856 4.26717
R1329 source.n764 source.n752 4.26717
R1330 source.n794 source.n738 4.26717
R1331 source.n813 source.n730 4.26717
R1332 source.n843 source.n716 4.26717
R1333 source.n620 source.n608 4.26717
R1334 source.n650 source.n594 4.26717
R1335 source.n669 source.n586 4.26717
R1336 source.n699 source.n572 4.26717
R1337 source.n131 source.n4 4.26717
R1338 source.n102 source.n19 4.26717
R1339 source.n83 source.n27 4.26717
R1340 source.n54 source.n42 4.26717
R1341 source.n275 source.n148 4.26717
R1342 source.n246 source.n163 4.26717
R1343 source.n227 source.n171 4.26717
R1344 source.n198 source.n186 4.26717
R1345 source.n415 source.n288 4.26717
R1346 source.n386 source.n303 4.26717
R1347 source.n367 source.n311 4.26717
R1348 source.n338 source.n326 4.26717
R1349 source.n559 source.n432 4.26717
R1350 source.n530 source.n447 4.26717
R1351 source.n511 source.n455 4.26717
R1352 source.n482 source.n470 4.26717
R1353 source.n1052 source.n1051 3.49141
R1354 source.n1077 source.n1024 3.49141
R1355 source.n1098 source.n1012 3.49141
R1356 source.n1124 source.n1123 3.49141
R1357 source.n908 source.n907 3.49141
R1358 source.n933 source.n880 3.49141
R1359 source.n954 source.n868 3.49141
R1360 source.n980 source.n979 3.49141
R1361 source.n768 source.n767 3.49141
R1362 source.n793 source.n740 3.49141
R1363 source.n814 source.n728 3.49141
R1364 source.n840 source.n839 3.49141
R1365 source.n624 source.n623 3.49141
R1366 source.n649 source.n596 3.49141
R1367 source.n670 source.n584 3.49141
R1368 source.n696 source.n695 3.49141
R1369 source.n128 source.n127 3.49141
R1370 source.n103 source.n17 3.49141
R1371 source.n82 source.n29 3.49141
R1372 source.n58 source.n57 3.49141
R1373 source.n272 source.n271 3.49141
R1374 source.n247 source.n161 3.49141
R1375 source.n226 source.n173 3.49141
R1376 source.n202 source.n201 3.49141
R1377 source.n412 source.n411 3.49141
R1378 source.n387 source.n301 3.49141
R1379 source.n366 source.n313 3.49141
R1380 source.n342 source.n341 3.49141
R1381 source.n556 source.n555 3.49141
R1382 source.n531 source.n445 3.49141
R1383 source.n510 source.n457 3.49141
R1384 source.n486 source.n485 3.49141
R1385 source.n48 source.n47 2.84303
R1386 source.n192 source.n191 2.84303
R1387 source.n332 source.n331 2.84303
R1388 source.n476 source.n475 2.84303
R1389 source.n1042 source.n1041 2.84303
R1390 source.n898 source.n897 2.84303
R1391 source.n758 source.n757 2.84303
R1392 source.n614 source.n613 2.84303
R1393 source.n1055 source.n1034 2.71565
R1394 source.n1074 source.n1073 2.71565
R1395 source.n1102 source.n1101 2.71565
R1396 source.n1120 source.n1002 2.71565
R1397 source.n911 source.n890 2.71565
R1398 source.n930 source.n929 2.71565
R1399 source.n958 source.n957 2.71565
R1400 source.n976 source.n858 2.71565
R1401 source.n771 source.n750 2.71565
R1402 source.n790 source.n789 2.71565
R1403 source.n818 source.n817 2.71565
R1404 source.n836 source.n718 2.71565
R1405 source.n627 source.n606 2.71565
R1406 source.n646 source.n645 2.71565
R1407 source.n674 source.n673 2.71565
R1408 source.n692 source.n574 2.71565
R1409 source.n124 source.n6 2.71565
R1410 source.n107 source.n106 2.71565
R1411 source.n79 source.n78 2.71565
R1412 source.n61 source.n40 2.71565
R1413 source.n268 source.n150 2.71565
R1414 source.n251 source.n250 2.71565
R1415 source.n223 source.n222 2.71565
R1416 source.n205 source.n184 2.71565
R1417 source.n408 source.n290 2.71565
R1418 source.n391 source.n390 2.71565
R1419 source.n363 source.n362 2.71565
R1420 source.n345 source.n324 2.71565
R1421 source.n552 source.n434 2.71565
R1422 source.n535 source.n534 2.71565
R1423 source.n507 source.n506 2.71565
R1424 source.n489 source.n468 2.71565
R1425 source.n1056 source.n1032 1.93989
R1426 source.n1070 source.n1026 1.93989
R1427 source.n1106 source.n1010 1.93989
R1428 source.n1119 source.n1004 1.93989
R1429 source.n912 source.n888 1.93989
R1430 source.n926 source.n882 1.93989
R1431 source.n962 source.n866 1.93989
R1432 source.n975 source.n860 1.93989
R1433 source.n772 source.n748 1.93989
R1434 source.n786 source.n742 1.93989
R1435 source.n822 source.n726 1.93989
R1436 source.n835 source.n720 1.93989
R1437 source.n628 source.n604 1.93989
R1438 source.n642 source.n598 1.93989
R1439 source.n678 source.n582 1.93989
R1440 source.n691 source.n576 1.93989
R1441 source.n123 source.n8 1.93989
R1442 source.n110 source.n14 1.93989
R1443 source.n75 source.n31 1.93989
R1444 source.n62 source.n38 1.93989
R1445 source.n267 source.n152 1.93989
R1446 source.n254 source.n158 1.93989
R1447 source.n219 source.n175 1.93989
R1448 source.n206 source.n182 1.93989
R1449 source.n407 source.n292 1.93989
R1450 source.n394 source.n298 1.93989
R1451 source.n359 source.n315 1.93989
R1452 source.n346 source.n322 1.93989
R1453 source.n551 source.n436 1.93989
R1454 source.n538 source.n442 1.93989
R1455 source.n503 source.n459 1.93989
R1456 source.n490 source.n466 1.93989
R1457 source.n1061 source.n1059 1.16414
R1458 source.n1069 source.n1028 1.16414
R1459 source.n1107 source.n1008 1.16414
R1460 source.n1116 source.n1115 1.16414
R1461 source.n917 source.n915 1.16414
R1462 source.n925 source.n884 1.16414
R1463 source.n963 source.n864 1.16414
R1464 source.n972 source.n971 1.16414
R1465 source.n777 source.n775 1.16414
R1466 source.n785 source.n744 1.16414
R1467 source.n823 source.n724 1.16414
R1468 source.n832 source.n831 1.16414
R1469 source.n633 source.n631 1.16414
R1470 source.n641 source.n600 1.16414
R1471 source.n679 source.n580 1.16414
R1472 source.n688 source.n687 1.16414
R1473 source.n120 source.n119 1.16414
R1474 source.n111 source.n12 1.16414
R1475 source.n74 source.n33 1.16414
R1476 source.n66 source.n65 1.16414
R1477 source.n264 source.n263 1.16414
R1478 source.n255 source.n156 1.16414
R1479 source.n218 source.n177 1.16414
R1480 source.n210 source.n209 1.16414
R1481 source.n404 source.n403 1.16414
R1482 source.n395 source.n296 1.16414
R1483 source.n358 source.n317 1.16414
R1484 source.n350 source.n349 1.16414
R1485 source.n548 source.n547 1.16414
R1486 source.n539 source.n440 1.16414
R1487 source.n502 source.n461 1.16414
R1488 source.n494 source.n493 1.16414
R1489 source.n567 source.n427 0.888431
R1490 source.n427 source.n425 0.888431
R1491 source.n425 source.n423 0.888431
R1492 source.n283 source.n143 0.888431
R1493 source.n143 source.n141 0.888431
R1494 source.n141 source.n139 0.888431
R1495 source.n709 source.n707 0.888431
R1496 source.n711 source.n709 0.888431
R1497 source.n851 source.n711 0.888431
R1498 source.n993 source.n991 0.888431
R1499 source.n995 source.n993 0.888431
R1500 source.n1135 source.n995 0.888431
R1501 source.n994 source.t19 0.7925
R1502 source.n994 source.t17 0.7925
R1503 source.n992 source.t16 0.7925
R1504 source.n992 source.t20 0.7925
R1505 source.n710 source.t4 0.7925
R1506 source.n710 source.t21 0.7925
R1507 source.n708 source.t8 0.7925
R1508 source.n708 source.t3 0.7925
R1509 source.n140 source.t5 0.7925
R1510 source.n140 source.t1 0.7925
R1511 source.n142 source.t23 0.7925
R1512 source.n142 source.t22 0.7925
R1513 source.n424 source.t13 0.7925
R1514 source.n424 source.t18 0.7925
R1515 source.n426 source.t14 0.7925
R1516 source.n426 source.t10 0.7925
R1517 source.n423 source.n283 0.470328
R1518 source.n991 source.n851 0.470328
R1519 source.n1060 source.n1030 0.388379
R1520 source.n1066 source.n1065 0.388379
R1521 source.n1111 source.n1110 0.388379
R1522 source.n1112 source.n1006 0.388379
R1523 source.n916 source.n886 0.388379
R1524 source.n922 source.n921 0.388379
R1525 source.n967 source.n966 0.388379
R1526 source.n968 source.n862 0.388379
R1527 source.n776 source.n746 0.388379
R1528 source.n782 source.n781 0.388379
R1529 source.n827 source.n826 0.388379
R1530 source.n828 source.n722 0.388379
R1531 source.n632 source.n602 0.388379
R1532 source.n638 source.n637 0.388379
R1533 source.n683 source.n682 0.388379
R1534 source.n684 source.n578 0.388379
R1535 source.n116 source.n10 0.388379
R1536 source.n115 source.n114 0.388379
R1537 source.n71 source.n70 0.388379
R1538 source.n37 source.n35 0.388379
R1539 source.n260 source.n154 0.388379
R1540 source.n259 source.n258 0.388379
R1541 source.n215 source.n214 0.388379
R1542 source.n181 source.n179 0.388379
R1543 source.n400 source.n294 0.388379
R1544 source.n399 source.n398 0.388379
R1545 source.n355 source.n354 0.388379
R1546 source.n321 source.n319 0.388379
R1547 source.n544 source.n438 0.388379
R1548 source.n543 source.n542 0.388379
R1549 source.n499 source.n498 0.388379
R1550 source.n465 source.n463 0.388379
R1551 source source.n1136 0.188
R1552 source.n1042 source.n1037 0.155672
R1553 source.n1049 source.n1037 0.155672
R1554 source.n1050 source.n1049 0.155672
R1555 source.n1050 source.n1033 0.155672
R1556 source.n1057 source.n1033 0.155672
R1557 source.n1058 source.n1057 0.155672
R1558 source.n1058 source.n1029 0.155672
R1559 source.n1067 source.n1029 0.155672
R1560 source.n1068 source.n1067 0.155672
R1561 source.n1068 source.n1025 0.155672
R1562 source.n1075 source.n1025 0.155672
R1563 source.n1076 source.n1075 0.155672
R1564 source.n1076 source.n1021 0.155672
R1565 source.n1083 source.n1021 0.155672
R1566 source.n1084 source.n1083 0.155672
R1567 source.n1084 source.n1017 0.155672
R1568 source.n1091 source.n1017 0.155672
R1569 source.n1092 source.n1091 0.155672
R1570 source.n1092 source.n1013 0.155672
R1571 source.n1099 source.n1013 0.155672
R1572 source.n1100 source.n1099 0.155672
R1573 source.n1100 source.n1009 0.155672
R1574 source.n1108 source.n1009 0.155672
R1575 source.n1109 source.n1108 0.155672
R1576 source.n1109 source.n1005 0.155672
R1577 source.n1117 source.n1005 0.155672
R1578 source.n1118 source.n1117 0.155672
R1579 source.n1118 source.n1001 0.155672
R1580 source.n1125 source.n1001 0.155672
R1581 source.n1126 source.n1125 0.155672
R1582 source.n1126 source.n997 0.155672
R1583 source.n1133 source.n997 0.155672
R1584 source.n898 source.n893 0.155672
R1585 source.n905 source.n893 0.155672
R1586 source.n906 source.n905 0.155672
R1587 source.n906 source.n889 0.155672
R1588 source.n913 source.n889 0.155672
R1589 source.n914 source.n913 0.155672
R1590 source.n914 source.n885 0.155672
R1591 source.n923 source.n885 0.155672
R1592 source.n924 source.n923 0.155672
R1593 source.n924 source.n881 0.155672
R1594 source.n931 source.n881 0.155672
R1595 source.n932 source.n931 0.155672
R1596 source.n932 source.n877 0.155672
R1597 source.n939 source.n877 0.155672
R1598 source.n940 source.n939 0.155672
R1599 source.n940 source.n873 0.155672
R1600 source.n947 source.n873 0.155672
R1601 source.n948 source.n947 0.155672
R1602 source.n948 source.n869 0.155672
R1603 source.n955 source.n869 0.155672
R1604 source.n956 source.n955 0.155672
R1605 source.n956 source.n865 0.155672
R1606 source.n964 source.n865 0.155672
R1607 source.n965 source.n964 0.155672
R1608 source.n965 source.n861 0.155672
R1609 source.n973 source.n861 0.155672
R1610 source.n974 source.n973 0.155672
R1611 source.n974 source.n857 0.155672
R1612 source.n981 source.n857 0.155672
R1613 source.n982 source.n981 0.155672
R1614 source.n982 source.n853 0.155672
R1615 source.n989 source.n853 0.155672
R1616 source.n758 source.n753 0.155672
R1617 source.n765 source.n753 0.155672
R1618 source.n766 source.n765 0.155672
R1619 source.n766 source.n749 0.155672
R1620 source.n773 source.n749 0.155672
R1621 source.n774 source.n773 0.155672
R1622 source.n774 source.n745 0.155672
R1623 source.n783 source.n745 0.155672
R1624 source.n784 source.n783 0.155672
R1625 source.n784 source.n741 0.155672
R1626 source.n791 source.n741 0.155672
R1627 source.n792 source.n791 0.155672
R1628 source.n792 source.n737 0.155672
R1629 source.n799 source.n737 0.155672
R1630 source.n800 source.n799 0.155672
R1631 source.n800 source.n733 0.155672
R1632 source.n807 source.n733 0.155672
R1633 source.n808 source.n807 0.155672
R1634 source.n808 source.n729 0.155672
R1635 source.n815 source.n729 0.155672
R1636 source.n816 source.n815 0.155672
R1637 source.n816 source.n725 0.155672
R1638 source.n824 source.n725 0.155672
R1639 source.n825 source.n824 0.155672
R1640 source.n825 source.n721 0.155672
R1641 source.n833 source.n721 0.155672
R1642 source.n834 source.n833 0.155672
R1643 source.n834 source.n717 0.155672
R1644 source.n841 source.n717 0.155672
R1645 source.n842 source.n841 0.155672
R1646 source.n842 source.n713 0.155672
R1647 source.n849 source.n713 0.155672
R1648 source.n614 source.n609 0.155672
R1649 source.n621 source.n609 0.155672
R1650 source.n622 source.n621 0.155672
R1651 source.n622 source.n605 0.155672
R1652 source.n629 source.n605 0.155672
R1653 source.n630 source.n629 0.155672
R1654 source.n630 source.n601 0.155672
R1655 source.n639 source.n601 0.155672
R1656 source.n640 source.n639 0.155672
R1657 source.n640 source.n597 0.155672
R1658 source.n647 source.n597 0.155672
R1659 source.n648 source.n647 0.155672
R1660 source.n648 source.n593 0.155672
R1661 source.n655 source.n593 0.155672
R1662 source.n656 source.n655 0.155672
R1663 source.n656 source.n589 0.155672
R1664 source.n663 source.n589 0.155672
R1665 source.n664 source.n663 0.155672
R1666 source.n664 source.n585 0.155672
R1667 source.n671 source.n585 0.155672
R1668 source.n672 source.n671 0.155672
R1669 source.n672 source.n581 0.155672
R1670 source.n680 source.n581 0.155672
R1671 source.n681 source.n680 0.155672
R1672 source.n681 source.n577 0.155672
R1673 source.n689 source.n577 0.155672
R1674 source.n690 source.n689 0.155672
R1675 source.n690 source.n573 0.155672
R1676 source.n697 source.n573 0.155672
R1677 source.n698 source.n697 0.155672
R1678 source.n698 source.n569 0.155672
R1679 source.n705 source.n569 0.155672
R1680 source.n137 source.n1 0.155672
R1681 source.n130 source.n1 0.155672
R1682 source.n130 source.n129 0.155672
R1683 source.n129 source.n5 0.155672
R1684 source.n122 source.n5 0.155672
R1685 source.n122 source.n121 0.155672
R1686 source.n121 source.n9 0.155672
R1687 source.n113 source.n9 0.155672
R1688 source.n113 source.n112 0.155672
R1689 source.n112 source.n13 0.155672
R1690 source.n105 source.n13 0.155672
R1691 source.n105 source.n104 0.155672
R1692 source.n104 source.n18 0.155672
R1693 source.n97 source.n18 0.155672
R1694 source.n97 source.n96 0.155672
R1695 source.n96 source.n22 0.155672
R1696 source.n89 source.n22 0.155672
R1697 source.n89 source.n88 0.155672
R1698 source.n88 source.n26 0.155672
R1699 source.n81 source.n26 0.155672
R1700 source.n81 source.n80 0.155672
R1701 source.n80 source.n30 0.155672
R1702 source.n73 source.n30 0.155672
R1703 source.n73 source.n72 0.155672
R1704 source.n72 source.n34 0.155672
R1705 source.n64 source.n34 0.155672
R1706 source.n64 source.n63 0.155672
R1707 source.n63 source.n39 0.155672
R1708 source.n56 source.n39 0.155672
R1709 source.n56 source.n55 0.155672
R1710 source.n55 source.n43 0.155672
R1711 source.n48 source.n43 0.155672
R1712 source.n281 source.n145 0.155672
R1713 source.n274 source.n145 0.155672
R1714 source.n274 source.n273 0.155672
R1715 source.n273 source.n149 0.155672
R1716 source.n266 source.n149 0.155672
R1717 source.n266 source.n265 0.155672
R1718 source.n265 source.n153 0.155672
R1719 source.n257 source.n153 0.155672
R1720 source.n257 source.n256 0.155672
R1721 source.n256 source.n157 0.155672
R1722 source.n249 source.n157 0.155672
R1723 source.n249 source.n248 0.155672
R1724 source.n248 source.n162 0.155672
R1725 source.n241 source.n162 0.155672
R1726 source.n241 source.n240 0.155672
R1727 source.n240 source.n166 0.155672
R1728 source.n233 source.n166 0.155672
R1729 source.n233 source.n232 0.155672
R1730 source.n232 source.n170 0.155672
R1731 source.n225 source.n170 0.155672
R1732 source.n225 source.n224 0.155672
R1733 source.n224 source.n174 0.155672
R1734 source.n217 source.n174 0.155672
R1735 source.n217 source.n216 0.155672
R1736 source.n216 source.n178 0.155672
R1737 source.n208 source.n178 0.155672
R1738 source.n208 source.n207 0.155672
R1739 source.n207 source.n183 0.155672
R1740 source.n200 source.n183 0.155672
R1741 source.n200 source.n199 0.155672
R1742 source.n199 source.n187 0.155672
R1743 source.n192 source.n187 0.155672
R1744 source.n421 source.n285 0.155672
R1745 source.n414 source.n285 0.155672
R1746 source.n414 source.n413 0.155672
R1747 source.n413 source.n289 0.155672
R1748 source.n406 source.n289 0.155672
R1749 source.n406 source.n405 0.155672
R1750 source.n405 source.n293 0.155672
R1751 source.n397 source.n293 0.155672
R1752 source.n397 source.n396 0.155672
R1753 source.n396 source.n297 0.155672
R1754 source.n389 source.n297 0.155672
R1755 source.n389 source.n388 0.155672
R1756 source.n388 source.n302 0.155672
R1757 source.n381 source.n302 0.155672
R1758 source.n381 source.n380 0.155672
R1759 source.n380 source.n306 0.155672
R1760 source.n373 source.n306 0.155672
R1761 source.n373 source.n372 0.155672
R1762 source.n372 source.n310 0.155672
R1763 source.n365 source.n310 0.155672
R1764 source.n365 source.n364 0.155672
R1765 source.n364 source.n314 0.155672
R1766 source.n357 source.n314 0.155672
R1767 source.n357 source.n356 0.155672
R1768 source.n356 source.n318 0.155672
R1769 source.n348 source.n318 0.155672
R1770 source.n348 source.n347 0.155672
R1771 source.n347 source.n323 0.155672
R1772 source.n340 source.n323 0.155672
R1773 source.n340 source.n339 0.155672
R1774 source.n339 source.n327 0.155672
R1775 source.n332 source.n327 0.155672
R1776 source.n565 source.n429 0.155672
R1777 source.n558 source.n429 0.155672
R1778 source.n558 source.n557 0.155672
R1779 source.n557 source.n433 0.155672
R1780 source.n550 source.n433 0.155672
R1781 source.n550 source.n549 0.155672
R1782 source.n549 source.n437 0.155672
R1783 source.n541 source.n437 0.155672
R1784 source.n541 source.n540 0.155672
R1785 source.n540 source.n441 0.155672
R1786 source.n533 source.n441 0.155672
R1787 source.n533 source.n532 0.155672
R1788 source.n532 source.n446 0.155672
R1789 source.n525 source.n446 0.155672
R1790 source.n525 source.n524 0.155672
R1791 source.n524 source.n450 0.155672
R1792 source.n517 source.n450 0.155672
R1793 source.n517 source.n516 0.155672
R1794 source.n516 source.n454 0.155672
R1795 source.n509 source.n454 0.155672
R1796 source.n509 source.n508 0.155672
R1797 source.n508 source.n458 0.155672
R1798 source.n501 source.n458 0.155672
R1799 source.n501 source.n500 0.155672
R1800 source.n500 source.n462 0.155672
R1801 source.n492 source.n462 0.155672
R1802 source.n492 source.n491 0.155672
R1803 source.n491 source.n467 0.155672
R1804 source.n484 source.n467 0.155672
R1805 source.n484 source.n483 0.155672
R1806 source.n483 source.n471 0.155672
R1807 source.n476 source.n471 0.155672
R1808 plus.n5 plus.t4 940.138
R1809 plus.n23 plus.t11 940.138
R1810 plus.n16 plus.t8 916.833
R1811 plus.n14 plus.t3 916.833
R1812 plus.n2 plus.t6 916.833
R1813 plus.n8 plus.t1 916.833
R1814 plus.n4 plus.t9 916.833
R1815 plus.n34 plus.t2 916.833
R1816 plus.n32 plus.t7 916.833
R1817 plus.n20 plus.t5 916.833
R1818 plus.n26 plus.t10 916.833
R1819 plus.n22 plus.t0 916.833
R1820 plus.n7 plus.n6 161.3
R1821 plus.n8 plus.n3 161.3
R1822 plus.n10 plus.n9 161.3
R1823 plus.n11 plus.n2 161.3
R1824 plus.n13 plus.n12 161.3
R1825 plus.n14 plus.n1 161.3
R1826 plus.n15 plus.n0 161.3
R1827 plus.n17 plus.n16 161.3
R1828 plus.n25 plus.n24 161.3
R1829 plus.n26 plus.n21 161.3
R1830 plus.n28 plus.n27 161.3
R1831 plus.n29 plus.n20 161.3
R1832 plus.n31 plus.n30 161.3
R1833 plus.n32 plus.n19 161.3
R1834 plus.n33 plus.n18 161.3
R1835 plus.n35 plus.n34 161.3
R1836 plus.n6 plus.n5 44.8907
R1837 plus.n24 plus.n23 44.8907
R1838 plus plus.n35 36.2452
R1839 plus.n16 plus.n15 32.8641
R1840 plus.n34 plus.n33 32.8641
R1841 plus.n14 plus.n13 28.4823
R1842 plus.n7 plus.n4 28.4823
R1843 plus.n32 plus.n31 28.4823
R1844 plus.n25 plus.n22 28.4823
R1845 plus.n9 plus.n8 24.1005
R1846 plus.n9 plus.n2 24.1005
R1847 plus.n27 plus.n20 24.1005
R1848 plus.n27 plus.n26 24.1005
R1849 plus.n13 plus.n2 19.7187
R1850 plus.n8 plus.n7 19.7187
R1851 plus.n31 plus.n20 19.7187
R1852 plus.n26 plus.n25 19.7187
R1853 plus.n5 plus.n4 18.4104
R1854 plus.n23 plus.n22 18.4104
R1855 plus plus.n17 17.2126
R1856 plus.n15 plus.n14 15.3369
R1857 plus.n33 plus.n32 15.3369
R1858 plus.n6 plus.n3 0.189894
R1859 plus.n10 plus.n3 0.189894
R1860 plus.n11 plus.n10 0.189894
R1861 plus.n12 plus.n11 0.189894
R1862 plus.n12 plus.n1 0.189894
R1863 plus.n1 plus.n0 0.189894
R1864 plus.n17 plus.n0 0.189894
R1865 plus.n35 plus.n18 0.189894
R1866 plus.n19 plus.n18 0.189894
R1867 plus.n30 plus.n19 0.189894
R1868 plus.n30 plus.n29 0.189894
R1869 plus.n29 plus.n28 0.189894
R1870 plus.n28 plus.n21 0.189894
R1871 plus.n24 plus.n21 0.189894
R1872 drain_left.n6 drain_left.n4 59.6034
R1873 drain_left.n3 drain_left.n2 59.548
R1874 drain_left.n3 drain_left.n0 59.548
R1875 drain_left.n3 drain_left.n1 58.7154
R1876 drain_left.n6 drain_left.n5 58.7154
R1877 drain_left.n8 drain_left.n7 58.7153
R1878 drain_left drain_left.n3 41.6552
R1879 drain_left drain_left.n8 6.54115
R1880 drain_left.n8 drain_left.n6 0.888431
R1881 drain_left.n1 drain_left.t6 0.7925
R1882 drain_left.n1 drain_left.t1 0.7925
R1883 drain_left.n2 drain_left.t11 0.7925
R1884 drain_left.n2 drain_left.t0 0.7925
R1885 drain_left.n0 drain_left.t9 0.7925
R1886 drain_left.n0 drain_left.t4 0.7925
R1887 drain_left.n7 drain_left.t8 0.7925
R1888 drain_left.n7 drain_left.t3 0.7925
R1889 drain_left.n5 drain_left.t10 0.7925
R1890 drain_left.n5 drain_left.t5 0.7925
R1891 drain_left.n4 drain_left.t7 0.7925
R1892 drain_left.n4 drain_left.t2 0.7925
C0 source plus 15.301901f
C1 drain_left plus 16.1126f
C2 source drain_left 29.2552f
C3 minus plus 8.2422f
C4 minus source 15.287901f
C5 minus drain_left 0.17184f
C6 drain_right plus 0.366822f
C7 source drain_right 29.257198f
C8 drain_left drain_right 1.08491f
C9 minus drain_right 15.900801f
C10 drain_right a_n2158_n5888# 8.587501f
C11 drain_left a_n2158_n5888# 8.89558f
C12 source a_n2158_n5888# 16.423769f
C13 minus a_n2158_n5888# 9.385561f
C14 plus a_n2158_n5888# 11.746301f
C15 drain_left.t9 a_n2158_n5888# 0.54064f
C16 drain_left.t4 a_n2158_n5888# 0.54064f
C17 drain_left.n0 a_n2158_n5888# 4.98811f
C18 drain_left.t6 a_n2158_n5888# 0.54064f
C19 drain_left.t1 a_n2158_n5888# 0.54064f
C20 drain_left.n1 a_n2158_n5888# 4.98259f
C21 drain_left.t11 a_n2158_n5888# 0.54064f
C22 drain_left.t0 a_n2158_n5888# 0.54064f
C23 drain_left.n2 a_n2158_n5888# 4.98811f
C24 drain_left.n3 a_n2158_n5888# 3.44097f
C25 drain_left.t7 a_n2158_n5888# 0.54064f
C26 drain_left.t2 a_n2158_n5888# 0.54064f
C27 drain_left.n4 a_n2158_n5888# 4.98853f
C28 drain_left.t10 a_n2158_n5888# 0.54064f
C29 drain_left.t5 a_n2158_n5888# 0.54064f
C30 drain_left.n5 a_n2158_n5888# 4.98259f
C31 drain_left.n6 a_n2158_n5888# 0.780916f
C32 drain_left.t8 a_n2158_n5888# 0.54064f
C33 drain_left.t3 a_n2158_n5888# 0.54064f
C34 drain_left.n7 a_n2158_n5888# 4.98257f
C35 drain_left.n8 a_n2158_n5888# 0.629987f
C36 plus.n0 a_n2158_n5888# 0.041568f
C37 plus.t8 a_n2158_n5888# 2.05576f
C38 plus.t3 a_n2158_n5888# 2.05576f
C39 plus.n1 a_n2158_n5888# 0.041568f
C40 plus.t6 a_n2158_n5888# 2.05576f
C41 plus.n2 a_n2158_n5888# 0.750457f
C42 plus.n3 a_n2158_n5888# 0.041568f
C43 plus.t1 a_n2158_n5888# 2.05576f
C44 plus.t9 a_n2158_n5888# 2.05576f
C45 plus.n4 a_n2158_n5888# 0.755106f
C46 plus.t4 a_n2158_n5888# 2.07436f
C47 plus.n5 a_n2158_n5888# 0.735577f
C48 plus.n6 a_n2158_n5888# 0.174384f
C49 plus.n7 a_n2158_n5888# 0.009433f
C50 plus.n8 a_n2158_n5888# 0.750457f
C51 plus.n9 a_n2158_n5888# 0.009433f
C52 plus.n10 a_n2158_n5888# 0.041568f
C53 plus.n11 a_n2158_n5888# 0.041568f
C54 plus.n12 a_n2158_n5888# 0.041568f
C55 plus.n13 a_n2158_n5888# 0.009433f
C56 plus.n14 a_n2158_n5888# 0.750457f
C57 plus.n15 a_n2158_n5888# 0.009433f
C58 plus.n16 a_n2158_n5888# 0.748535f
C59 plus.n17 a_n2158_n5888# 0.755496f
C60 plus.n18 a_n2158_n5888# 0.041568f
C61 plus.t2 a_n2158_n5888# 2.05576f
C62 plus.n19 a_n2158_n5888# 0.041568f
C63 plus.t7 a_n2158_n5888# 2.05576f
C64 plus.t5 a_n2158_n5888# 2.05576f
C65 plus.n20 a_n2158_n5888# 0.750457f
C66 plus.n21 a_n2158_n5888# 0.041568f
C67 plus.t10 a_n2158_n5888# 2.05576f
C68 plus.t0 a_n2158_n5888# 2.05576f
C69 plus.n22 a_n2158_n5888# 0.755106f
C70 plus.t11 a_n2158_n5888# 2.07436f
C71 plus.n23 a_n2158_n5888# 0.735577f
C72 plus.n24 a_n2158_n5888# 0.174384f
C73 plus.n25 a_n2158_n5888# 0.009433f
C74 plus.n26 a_n2158_n5888# 0.750457f
C75 plus.n27 a_n2158_n5888# 0.009433f
C76 plus.n28 a_n2158_n5888# 0.041568f
C77 plus.n29 a_n2158_n5888# 0.041568f
C78 plus.n30 a_n2158_n5888# 0.041568f
C79 plus.n31 a_n2158_n5888# 0.009433f
C80 plus.n32 a_n2158_n5888# 0.750457f
C81 plus.n33 a_n2158_n5888# 0.009433f
C82 plus.n34 a_n2158_n5888# 0.748535f
C83 plus.n35 a_n2158_n5888# 1.6856f
C84 source.n0 a_n2158_n5888# 0.029047f
C85 source.n1 a_n2158_n5888# 0.02107f
C86 source.n2 a_n2158_n5888# 0.011322f
C87 source.n3 a_n2158_n5888# 0.026761f
C88 source.n4 a_n2158_n5888# 0.011988f
C89 source.n5 a_n2158_n5888# 0.02107f
C90 source.n6 a_n2158_n5888# 0.011322f
C91 source.n7 a_n2158_n5888# 0.026761f
C92 source.n8 a_n2158_n5888# 0.011988f
C93 source.n9 a_n2158_n5888# 0.02107f
C94 source.n10 a_n2158_n5888# 0.011322f
C95 source.n11 a_n2158_n5888# 0.026761f
C96 source.n12 a_n2158_n5888# 0.011988f
C97 source.n13 a_n2158_n5888# 0.02107f
C98 source.n14 a_n2158_n5888# 0.011322f
C99 source.n15 a_n2158_n5888# 0.026761f
C100 source.n16 a_n2158_n5888# 0.026761f
C101 source.n17 a_n2158_n5888# 0.011988f
C102 source.n18 a_n2158_n5888# 0.02107f
C103 source.n19 a_n2158_n5888# 0.011322f
C104 source.n20 a_n2158_n5888# 0.026761f
C105 source.n21 a_n2158_n5888# 0.011988f
C106 source.n22 a_n2158_n5888# 0.02107f
C107 source.n23 a_n2158_n5888# 0.011322f
C108 source.n24 a_n2158_n5888# 0.026761f
C109 source.n25 a_n2158_n5888# 0.011988f
C110 source.n26 a_n2158_n5888# 0.02107f
C111 source.n27 a_n2158_n5888# 0.011322f
C112 source.n28 a_n2158_n5888# 0.026761f
C113 source.n29 a_n2158_n5888# 0.011988f
C114 source.n30 a_n2158_n5888# 0.02107f
C115 source.n31 a_n2158_n5888# 0.011322f
C116 source.n32 a_n2158_n5888# 0.026761f
C117 source.n33 a_n2158_n5888# 0.011988f
C118 source.n34 a_n2158_n5888# 0.02107f
C119 source.n35 a_n2158_n5888# 0.011655f
C120 source.n36 a_n2158_n5888# 0.026761f
C121 source.n37 a_n2158_n5888# 0.011322f
C122 source.n38 a_n2158_n5888# 0.011988f
C123 source.n39 a_n2158_n5888# 0.02107f
C124 source.n40 a_n2158_n5888# 0.011322f
C125 source.n41 a_n2158_n5888# 0.026761f
C126 source.n42 a_n2158_n5888# 0.011988f
C127 source.n43 a_n2158_n5888# 0.02107f
C128 source.n44 a_n2158_n5888# 0.011322f
C129 source.n45 a_n2158_n5888# 0.020071f
C130 source.n46 a_n2158_n5888# 0.018918f
C131 source.t0 a_n2158_n5888# 0.046673f
C132 source.n47 a_n2158_n5888# 0.257071f
C133 source.n48 a_n2158_n5888# 2.28126f
C134 source.n49 a_n2158_n5888# 0.011322f
C135 source.n50 a_n2158_n5888# 0.011988f
C136 source.n51 a_n2158_n5888# 0.026761f
C137 source.n52 a_n2158_n5888# 0.026761f
C138 source.n53 a_n2158_n5888# 0.011988f
C139 source.n54 a_n2158_n5888# 0.011322f
C140 source.n55 a_n2158_n5888# 0.02107f
C141 source.n56 a_n2158_n5888# 0.02107f
C142 source.n57 a_n2158_n5888# 0.011322f
C143 source.n58 a_n2158_n5888# 0.011988f
C144 source.n59 a_n2158_n5888# 0.026761f
C145 source.n60 a_n2158_n5888# 0.026761f
C146 source.n61 a_n2158_n5888# 0.011988f
C147 source.n62 a_n2158_n5888# 0.011322f
C148 source.n63 a_n2158_n5888# 0.02107f
C149 source.n64 a_n2158_n5888# 0.02107f
C150 source.n65 a_n2158_n5888# 0.011322f
C151 source.n66 a_n2158_n5888# 0.011988f
C152 source.n67 a_n2158_n5888# 0.026761f
C153 source.n68 a_n2158_n5888# 0.026761f
C154 source.n69 a_n2158_n5888# 0.026761f
C155 source.n70 a_n2158_n5888# 0.011655f
C156 source.n71 a_n2158_n5888# 0.011322f
C157 source.n72 a_n2158_n5888# 0.02107f
C158 source.n73 a_n2158_n5888# 0.02107f
C159 source.n74 a_n2158_n5888# 0.011322f
C160 source.n75 a_n2158_n5888# 0.011988f
C161 source.n76 a_n2158_n5888# 0.026761f
C162 source.n77 a_n2158_n5888# 0.026761f
C163 source.n78 a_n2158_n5888# 0.011988f
C164 source.n79 a_n2158_n5888# 0.011322f
C165 source.n80 a_n2158_n5888# 0.02107f
C166 source.n81 a_n2158_n5888# 0.02107f
C167 source.n82 a_n2158_n5888# 0.011322f
C168 source.n83 a_n2158_n5888# 0.011988f
C169 source.n84 a_n2158_n5888# 0.026761f
C170 source.n85 a_n2158_n5888# 0.026761f
C171 source.n86 a_n2158_n5888# 0.011988f
C172 source.n87 a_n2158_n5888# 0.011322f
C173 source.n88 a_n2158_n5888# 0.02107f
C174 source.n89 a_n2158_n5888# 0.02107f
C175 source.n90 a_n2158_n5888# 0.011322f
C176 source.n91 a_n2158_n5888# 0.011988f
C177 source.n92 a_n2158_n5888# 0.026761f
C178 source.n93 a_n2158_n5888# 0.026761f
C179 source.n94 a_n2158_n5888# 0.011988f
C180 source.n95 a_n2158_n5888# 0.011322f
C181 source.n96 a_n2158_n5888# 0.02107f
C182 source.n97 a_n2158_n5888# 0.02107f
C183 source.n98 a_n2158_n5888# 0.011322f
C184 source.n99 a_n2158_n5888# 0.011988f
C185 source.n100 a_n2158_n5888# 0.026761f
C186 source.n101 a_n2158_n5888# 0.026761f
C187 source.n102 a_n2158_n5888# 0.011988f
C188 source.n103 a_n2158_n5888# 0.011322f
C189 source.n104 a_n2158_n5888# 0.02107f
C190 source.n105 a_n2158_n5888# 0.02107f
C191 source.n106 a_n2158_n5888# 0.011322f
C192 source.n107 a_n2158_n5888# 0.011988f
C193 source.n108 a_n2158_n5888# 0.026761f
C194 source.n109 a_n2158_n5888# 0.026761f
C195 source.n110 a_n2158_n5888# 0.011988f
C196 source.n111 a_n2158_n5888# 0.011322f
C197 source.n112 a_n2158_n5888# 0.02107f
C198 source.n113 a_n2158_n5888# 0.02107f
C199 source.n114 a_n2158_n5888# 0.011322f
C200 source.n115 a_n2158_n5888# 0.011655f
C201 source.n116 a_n2158_n5888# 0.011655f
C202 source.n117 a_n2158_n5888# 0.026761f
C203 source.n118 a_n2158_n5888# 0.026761f
C204 source.n119 a_n2158_n5888# 0.011988f
C205 source.n120 a_n2158_n5888# 0.011322f
C206 source.n121 a_n2158_n5888# 0.02107f
C207 source.n122 a_n2158_n5888# 0.02107f
C208 source.n123 a_n2158_n5888# 0.011322f
C209 source.n124 a_n2158_n5888# 0.011988f
C210 source.n125 a_n2158_n5888# 0.026761f
C211 source.n126 a_n2158_n5888# 0.026761f
C212 source.n127 a_n2158_n5888# 0.011988f
C213 source.n128 a_n2158_n5888# 0.011322f
C214 source.n129 a_n2158_n5888# 0.02107f
C215 source.n130 a_n2158_n5888# 0.02107f
C216 source.n131 a_n2158_n5888# 0.011322f
C217 source.n132 a_n2158_n5888# 0.011988f
C218 source.n133 a_n2158_n5888# 0.026761f
C219 source.n134 a_n2158_n5888# 0.056928f
C220 source.n135 a_n2158_n5888# 0.011988f
C221 source.n136 a_n2158_n5888# 0.011322f
C222 source.n137 a_n2158_n5888# 0.0464f
C223 source.n138 a_n2158_n5888# 0.031678f
C224 source.n139 a_n2158_n5888# 1.69218f
C225 source.t5 a_n2158_n5888# 0.416253f
C226 source.t1 a_n2158_n5888# 0.416253f
C227 source.n140 a_n2158_n5888# 3.76715f
C228 source.n141 a_n2158_n5888# 0.339104f
C229 source.t23 a_n2158_n5888# 0.416253f
C230 source.t22 a_n2158_n5888# 0.416253f
C231 source.n142 a_n2158_n5888# 3.76715f
C232 source.n143 a_n2158_n5888# 0.339104f
C233 source.n144 a_n2158_n5888# 0.029047f
C234 source.n145 a_n2158_n5888# 0.02107f
C235 source.n146 a_n2158_n5888# 0.011322f
C236 source.n147 a_n2158_n5888# 0.026761f
C237 source.n148 a_n2158_n5888# 0.011988f
C238 source.n149 a_n2158_n5888# 0.02107f
C239 source.n150 a_n2158_n5888# 0.011322f
C240 source.n151 a_n2158_n5888# 0.026761f
C241 source.n152 a_n2158_n5888# 0.011988f
C242 source.n153 a_n2158_n5888# 0.02107f
C243 source.n154 a_n2158_n5888# 0.011322f
C244 source.n155 a_n2158_n5888# 0.026761f
C245 source.n156 a_n2158_n5888# 0.011988f
C246 source.n157 a_n2158_n5888# 0.02107f
C247 source.n158 a_n2158_n5888# 0.011322f
C248 source.n159 a_n2158_n5888# 0.026761f
C249 source.n160 a_n2158_n5888# 0.026761f
C250 source.n161 a_n2158_n5888# 0.011988f
C251 source.n162 a_n2158_n5888# 0.02107f
C252 source.n163 a_n2158_n5888# 0.011322f
C253 source.n164 a_n2158_n5888# 0.026761f
C254 source.n165 a_n2158_n5888# 0.011988f
C255 source.n166 a_n2158_n5888# 0.02107f
C256 source.n167 a_n2158_n5888# 0.011322f
C257 source.n168 a_n2158_n5888# 0.026761f
C258 source.n169 a_n2158_n5888# 0.011988f
C259 source.n170 a_n2158_n5888# 0.02107f
C260 source.n171 a_n2158_n5888# 0.011322f
C261 source.n172 a_n2158_n5888# 0.026761f
C262 source.n173 a_n2158_n5888# 0.011988f
C263 source.n174 a_n2158_n5888# 0.02107f
C264 source.n175 a_n2158_n5888# 0.011322f
C265 source.n176 a_n2158_n5888# 0.026761f
C266 source.n177 a_n2158_n5888# 0.011988f
C267 source.n178 a_n2158_n5888# 0.02107f
C268 source.n179 a_n2158_n5888# 0.011655f
C269 source.n180 a_n2158_n5888# 0.026761f
C270 source.n181 a_n2158_n5888# 0.011322f
C271 source.n182 a_n2158_n5888# 0.011988f
C272 source.n183 a_n2158_n5888# 0.02107f
C273 source.n184 a_n2158_n5888# 0.011322f
C274 source.n185 a_n2158_n5888# 0.026761f
C275 source.n186 a_n2158_n5888# 0.011988f
C276 source.n187 a_n2158_n5888# 0.02107f
C277 source.n188 a_n2158_n5888# 0.011322f
C278 source.n189 a_n2158_n5888# 0.020071f
C279 source.n190 a_n2158_n5888# 0.018918f
C280 source.t7 a_n2158_n5888# 0.046673f
C281 source.n191 a_n2158_n5888# 0.257071f
C282 source.n192 a_n2158_n5888# 2.28126f
C283 source.n193 a_n2158_n5888# 0.011322f
C284 source.n194 a_n2158_n5888# 0.011988f
C285 source.n195 a_n2158_n5888# 0.026761f
C286 source.n196 a_n2158_n5888# 0.026761f
C287 source.n197 a_n2158_n5888# 0.011988f
C288 source.n198 a_n2158_n5888# 0.011322f
C289 source.n199 a_n2158_n5888# 0.02107f
C290 source.n200 a_n2158_n5888# 0.02107f
C291 source.n201 a_n2158_n5888# 0.011322f
C292 source.n202 a_n2158_n5888# 0.011988f
C293 source.n203 a_n2158_n5888# 0.026761f
C294 source.n204 a_n2158_n5888# 0.026761f
C295 source.n205 a_n2158_n5888# 0.011988f
C296 source.n206 a_n2158_n5888# 0.011322f
C297 source.n207 a_n2158_n5888# 0.02107f
C298 source.n208 a_n2158_n5888# 0.02107f
C299 source.n209 a_n2158_n5888# 0.011322f
C300 source.n210 a_n2158_n5888# 0.011988f
C301 source.n211 a_n2158_n5888# 0.026761f
C302 source.n212 a_n2158_n5888# 0.026761f
C303 source.n213 a_n2158_n5888# 0.026761f
C304 source.n214 a_n2158_n5888# 0.011655f
C305 source.n215 a_n2158_n5888# 0.011322f
C306 source.n216 a_n2158_n5888# 0.02107f
C307 source.n217 a_n2158_n5888# 0.02107f
C308 source.n218 a_n2158_n5888# 0.011322f
C309 source.n219 a_n2158_n5888# 0.011988f
C310 source.n220 a_n2158_n5888# 0.026761f
C311 source.n221 a_n2158_n5888# 0.026761f
C312 source.n222 a_n2158_n5888# 0.011988f
C313 source.n223 a_n2158_n5888# 0.011322f
C314 source.n224 a_n2158_n5888# 0.02107f
C315 source.n225 a_n2158_n5888# 0.02107f
C316 source.n226 a_n2158_n5888# 0.011322f
C317 source.n227 a_n2158_n5888# 0.011988f
C318 source.n228 a_n2158_n5888# 0.026761f
C319 source.n229 a_n2158_n5888# 0.026761f
C320 source.n230 a_n2158_n5888# 0.011988f
C321 source.n231 a_n2158_n5888# 0.011322f
C322 source.n232 a_n2158_n5888# 0.02107f
C323 source.n233 a_n2158_n5888# 0.02107f
C324 source.n234 a_n2158_n5888# 0.011322f
C325 source.n235 a_n2158_n5888# 0.011988f
C326 source.n236 a_n2158_n5888# 0.026761f
C327 source.n237 a_n2158_n5888# 0.026761f
C328 source.n238 a_n2158_n5888# 0.011988f
C329 source.n239 a_n2158_n5888# 0.011322f
C330 source.n240 a_n2158_n5888# 0.02107f
C331 source.n241 a_n2158_n5888# 0.02107f
C332 source.n242 a_n2158_n5888# 0.011322f
C333 source.n243 a_n2158_n5888# 0.011988f
C334 source.n244 a_n2158_n5888# 0.026761f
C335 source.n245 a_n2158_n5888# 0.026761f
C336 source.n246 a_n2158_n5888# 0.011988f
C337 source.n247 a_n2158_n5888# 0.011322f
C338 source.n248 a_n2158_n5888# 0.02107f
C339 source.n249 a_n2158_n5888# 0.02107f
C340 source.n250 a_n2158_n5888# 0.011322f
C341 source.n251 a_n2158_n5888# 0.011988f
C342 source.n252 a_n2158_n5888# 0.026761f
C343 source.n253 a_n2158_n5888# 0.026761f
C344 source.n254 a_n2158_n5888# 0.011988f
C345 source.n255 a_n2158_n5888# 0.011322f
C346 source.n256 a_n2158_n5888# 0.02107f
C347 source.n257 a_n2158_n5888# 0.02107f
C348 source.n258 a_n2158_n5888# 0.011322f
C349 source.n259 a_n2158_n5888# 0.011655f
C350 source.n260 a_n2158_n5888# 0.011655f
C351 source.n261 a_n2158_n5888# 0.026761f
C352 source.n262 a_n2158_n5888# 0.026761f
C353 source.n263 a_n2158_n5888# 0.011988f
C354 source.n264 a_n2158_n5888# 0.011322f
C355 source.n265 a_n2158_n5888# 0.02107f
C356 source.n266 a_n2158_n5888# 0.02107f
C357 source.n267 a_n2158_n5888# 0.011322f
C358 source.n268 a_n2158_n5888# 0.011988f
C359 source.n269 a_n2158_n5888# 0.026761f
C360 source.n270 a_n2158_n5888# 0.026761f
C361 source.n271 a_n2158_n5888# 0.011988f
C362 source.n272 a_n2158_n5888# 0.011322f
C363 source.n273 a_n2158_n5888# 0.02107f
C364 source.n274 a_n2158_n5888# 0.02107f
C365 source.n275 a_n2158_n5888# 0.011322f
C366 source.n276 a_n2158_n5888# 0.011988f
C367 source.n277 a_n2158_n5888# 0.026761f
C368 source.n278 a_n2158_n5888# 0.056928f
C369 source.n279 a_n2158_n5888# 0.011988f
C370 source.n280 a_n2158_n5888# 0.011322f
C371 source.n281 a_n2158_n5888# 0.0464f
C372 source.n282 a_n2158_n5888# 0.031678f
C373 source.n283 a_n2158_n5888# 0.108878f
C374 source.n284 a_n2158_n5888# 0.029047f
C375 source.n285 a_n2158_n5888# 0.02107f
C376 source.n286 a_n2158_n5888# 0.011322f
C377 source.n287 a_n2158_n5888# 0.026761f
C378 source.n288 a_n2158_n5888# 0.011988f
C379 source.n289 a_n2158_n5888# 0.02107f
C380 source.n290 a_n2158_n5888# 0.011322f
C381 source.n291 a_n2158_n5888# 0.026761f
C382 source.n292 a_n2158_n5888# 0.011988f
C383 source.n293 a_n2158_n5888# 0.02107f
C384 source.n294 a_n2158_n5888# 0.011322f
C385 source.n295 a_n2158_n5888# 0.026761f
C386 source.n296 a_n2158_n5888# 0.011988f
C387 source.n297 a_n2158_n5888# 0.02107f
C388 source.n298 a_n2158_n5888# 0.011322f
C389 source.n299 a_n2158_n5888# 0.026761f
C390 source.n300 a_n2158_n5888# 0.026761f
C391 source.n301 a_n2158_n5888# 0.011988f
C392 source.n302 a_n2158_n5888# 0.02107f
C393 source.n303 a_n2158_n5888# 0.011322f
C394 source.n304 a_n2158_n5888# 0.026761f
C395 source.n305 a_n2158_n5888# 0.011988f
C396 source.n306 a_n2158_n5888# 0.02107f
C397 source.n307 a_n2158_n5888# 0.011322f
C398 source.n308 a_n2158_n5888# 0.026761f
C399 source.n309 a_n2158_n5888# 0.011988f
C400 source.n310 a_n2158_n5888# 0.02107f
C401 source.n311 a_n2158_n5888# 0.011322f
C402 source.n312 a_n2158_n5888# 0.026761f
C403 source.n313 a_n2158_n5888# 0.011988f
C404 source.n314 a_n2158_n5888# 0.02107f
C405 source.n315 a_n2158_n5888# 0.011322f
C406 source.n316 a_n2158_n5888# 0.026761f
C407 source.n317 a_n2158_n5888# 0.011988f
C408 source.n318 a_n2158_n5888# 0.02107f
C409 source.n319 a_n2158_n5888# 0.011655f
C410 source.n320 a_n2158_n5888# 0.026761f
C411 source.n321 a_n2158_n5888# 0.011322f
C412 source.n322 a_n2158_n5888# 0.011988f
C413 source.n323 a_n2158_n5888# 0.02107f
C414 source.n324 a_n2158_n5888# 0.011322f
C415 source.n325 a_n2158_n5888# 0.026761f
C416 source.n326 a_n2158_n5888# 0.011988f
C417 source.n327 a_n2158_n5888# 0.02107f
C418 source.n328 a_n2158_n5888# 0.011322f
C419 source.n329 a_n2158_n5888# 0.020071f
C420 source.n330 a_n2158_n5888# 0.018918f
C421 source.t12 a_n2158_n5888# 0.046673f
C422 source.n331 a_n2158_n5888# 0.257071f
C423 source.n332 a_n2158_n5888# 2.28126f
C424 source.n333 a_n2158_n5888# 0.011322f
C425 source.n334 a_n2158_n5888# 0.011988f
C426 source.n335 a_n2158_n5888# 0.026761f
C427 source.n336 a_n2158_n5888# 0.026761f
C428 source.n337 a_n2158_n5888# 0.011988f
C429 source.n338 a_n2158_n5888# 0.011322f
C430 source.n339 a_n2158_n5888# 0.02107f
C431 source.n340 a_n2158_n5888# 0.02107f
C432 source.n341 a_n2158_n5888# 0.011322f
C433 source.n342 a_n2158_n5888# 0.011988f
C434 source.n343 a_n2158_n5888# 0.026761f
C435 source.n344 a_n2158_n5888# 0.026761f
C436 source.n345 a_n2158_n5888# 0.011988f
C437 source.n346 a_n2158_n5888# 0.011322f
C438 source.n347 a_n2158_n5888# 0.02107f
C439 source.n348 a_n2158_n5888# 0.02107f
C440 source.n349 a_n2158_n5888# 0.011322f
C441 source.n350 a_n2158_n5888# 0.011988f
C442 source.n351 a_n2158_n5888# 0.026761f
C443 source.n352 a_n2158_n5888# 0.026761f
C444 source.n353 a_n2158_n5888# 0.026761f
C445 source.n354 a_n2158_n5888# 0.011655f
C446 source.n355 a_n2158_n5888# 0.011322f
C447 source.n356 a_n2158_n5888# 0.02107f
C448 source.n357 a_n2158_n5888# 0.02107f
C449 source.n358 a_n2158_n5888# 0.011322f
C450 source.n359 a_n2158_n5888# 0.011988f
C451 source.n360 a_n2158_n5888# 0.026761f
C452 source.n361 a_n2158_n5888# 0.026761f
C453 source.n362 a_n2158_n5888# 0.011988f
C454 source.n363 a_n2158_n5888# 0.011322f
C455 source.n364 a_n2158_n5888# 0.02107f
C456 source.n365 a_n2158_n5888# 0.02107f
C457 source.n366 a_n2158_n5888# 0.011322f
C458 source.n367 a_n2158_n5888# 0.011988f
C459 source.n368 a_n2158_n5888# 0.026761f
C460 source.n369 a_n2158_n5888# 0.026761f
C461 source.n370 a_n2158_n5888# 0.011988f
C462 source.n371 a_n2158_n5888# 0.011322f
C463 source.n372 a_n2158_n5888# 0.02107f
C464 source.n373 a_n2158_n5888# 0.02107f
C465 source.n374 a_n2158_n5888# 0.011322f
C466 source.n375 a_n2158_n5888# 0.011988f
C467 source.n376 a_n2158_n5888# 0.026761f
C468 source.n377 a_n2158_n5888# 0.026761f
C469 source.n378 a_n2158_n5888# 0.011988f
C470 source.n379 a_n2158_n5888# 0.011322f
C471 source.n380 a_n2158_n5888# 0.02107f
C472 source.n381 a_n2158_n5888# 0.02107f
C473 source.n382 a_n2158_n5888# 0.011322f
C474 source.n383 a_n2158_n5888# 0.011988f
C475 source.n384 a_n2158_n5888# 0.026761f
C476 source.n385 a_n2158_n5888# 0.026761f
C477 source.n386 a_n2158_n5888# 0.011988f
C478 source.n387 a_n2158_n5888# 0.011322f
C479 source.n388 a_n2158_n5888# 0.02107f
C480 source.n389 a_n2158_n5888# 0.02107f
C481 source.n390 a_n2158_n5888# 0.011322f
C482 source.n391 a_n2158_n5888# 0.011988f
C483 source.n392 a_n2158_n5888# 0.026761f
C484 source.n393 a_n2158_n5888# 0.026761f
C485 source.n394 a_n2158_n5888# 0.011988f
C486 source.n395 a_n2158_n5888# 0.011322f
C487 source.n396 a_n2158_n5888# 0.02107f
C488 source.n397 a_n2158_n5888# 0.02107f
C489 source.n398 a_n2158_n5888# 0.011322f
C490 source.n399 a_n2158_n5888# 0.011655f
C491 source.n400 a_n2158_n5888# 0.011655f
C492 source.n401 a_n2158_n5888# 0.026761f
C493 source.n402 a_n2158_n5888# 0.026761f
C494 source.n403 a_n2158_n5888# 0.011988f
C495 source.n404 a_n2158_n5888# 0.011322f
C496 source.n405 a_n2158_n5888# 0.02107f
C497 source.n406 a_n2158_n5888# 0.02107f
C498 source.n407 a_n2158_n5888# 0.011322f
C499 source.n408 a_n2158_n5888# 0.011988f
C500 source.n409 a_n2158_n5888# 0.026761f
C501 source.n410 a_n2158_n5888# 0.026761f
C502 source.n411 a_n2158_n5888# 0.011988f
C503 source.n412 a_n2158_n5888# 0.011322f
C504 source.n413 a_n2158_n5888# 0.02107f
C505 source.n414 a_n2158_n5888# 0.02107f
C506 source.n415 a_n2158_n5888# 0.011322f
C507 source.n416 a_n2158_n5888# 0.011988f
C508 source.n417 a_n2158_n5888# 0.026761f
C509 source.n418 a_n2158_n5888# 0.056928f
C510 source.n419 a_n2158_n5888# 0.011988f
C511 source.n420 a_n2158_n5888# 0.011322f
C512 source.n421 a_n2158_n5888# 0.0464f
C513 source.n422 a_n2158_n5888# 0.031678f
C514 source.n423 a_n2158_n5888# 0.108878f
C515 source.t13 a_n2158_n5888# 0.416253f
C516 source.t18 a_n2158_n5888# 0.416253f
C517 source.n424 a_n2158_n5888# 3.76715f
C518 source.n425 a_n2158_n5888# 0.339104f
C519 source.t14 a_n2158_n5888# 0.416253f
C520 source.t10 a_n2158_n5888# 0.416253f
C521 source.n426 a_n2158_n5888# 3.76715f
C522 source.n427 a_n2158_n5888# 0.339104f
C523 source.n428 a_n2158_n5888# 0.029047f
C524 source.n429 a_n2158_n5888# 0.02107f
C525 source.n430 a_n2158_n5888# 0.011322f
C526 source.n431 a_n2158_n5888# 0.026761f
C527 source.n432 a_n2158_n5888# 0.011988f
C528 source.n433 a_n2158_n5888# 0.02107f
C529 source.n434 a_n2158_n5888# 0.011322f
C530 source.n435 a_n2158_n5888# 0.026761f
C531 source.n436 a_n2158_n5888# 0.011988f
C532 source.n437 a_n2158_n5888# 0.02107f
C533 source.n438 a_n2158_n5888# 0.011322f
C534 source.n439 a_n2158_n5888# 0.026761f
C535 source.n440 a_n2158_n5888# 0.011988f
C536 source.n441 a_n2158_n5888# 0.02107f
C537 source.n442 a_n2158_n5888# 0.011322f
C538 source.n443 a_n2158_n5888# 0.026761f
C539 source.n444 a_n2158_n5888# 0.026761f
C540 source.n445 a_n2158_n5888# 0.011988f
C541 source.n446 a_n2158_n5888# 0.02107f
C542 source.n447 a_n2158_n5888# 0.011322f
C543 source.n448 a_n2158_n5888# 0.026761f
C544 source.n449 a_n2158_n5888# 0.011988f
C545 source.n450 a_n2158_n5888# 0.02107f
C546 source.n451 a_n2158_n5888# 0.011322f
C547 source.n452 a_n2158_n5888# 0.026761f
C548 source.n453 a_n2158_n5888# 0.011988f
C549 source.n454 a_n2158_n5888# 0.02107f
C550 source.n455 a_n2158_n5888# 0.011322f
C551 source.n456 a_n2158_n5888# 0.026761f
C552 source.n457 a_n2158_n5888# 0.011988f
C553 source.n458 a_n2158_n5888# 0.02107f
C554 source.n459 a_n2158_n5888# 0.011322f
C555 source.n460 a_n2158_n5888# 0.026761f
C556 source.n461 a_n2158_n5888# 0.011988f
C557 source.n462 a_n2158_n5888# 0.02107f
C558 source.n463 a_n2158_n5888# 0.011655f
C559 source.n464 a_n2158_n5888# 0.026761f
C560 source.n465 a_n2158_n5888# 0.011322f
C561 source.n466 a_n2158_n5888# 0.011988f
C562 source.n467 a_n2158_n5888# 0.02107f
C563 source.n468 a_n2158_n5888# 0.011322f
C564 source.n469 a_n2158_n5888# 0.026761f
C565 source.n470 a_n2158_n5888# 0.011988f
C566 source.n471 a_n2158_n5888# 0.02107f
C567 source.n472 a_n2158_n5888# 0.011322f
C568 source.n473 a_n2158_n5888# 0.020071f
C569 source.n474 a_n2158_n5888# 0.018918f
C570 source.t9 a_n2158_n5888# 0.046673f
C571 source.n475 a_n2158_n5888# 0.257071f
C572 source.n476 a_n2158_n5888# 2.28126f
C573 source.n477 a_n2158_n5888# 0.011322f
C574 source.n478 a_n2158_n5888# 0.011988f
C575 source.n479 a_n2158_n5888# 0.026761f
C576 source.n480 a_n2158_n5888# 0.026761f
C577 source.n481 a_n2158_n5888# 0.011988f
C578 source.n482 a_n2158_n5888# 0.011322f
C579 source.n483 a_n2158_n5888# 0.02107f
C580 source.n484 a_n2158_n5888# 0.02107f
C581 source.n485 a_n2158_n5888# 0.011322f
C582 source.n486 a_n2158_n5888# 0.011988f
C583 source.n487 a_n2158_n5888# 0.026761f
C584 source.n488 a_n2158_n5888# 0.026761f
C585 source.n489 a_n2158_n5888# 0.011988f
C586 source.n490 a_n2158_n5888# 0.011322f
C587 source.n491 a_n2158_n5888# 0.02107f
C588 source.n492 a_n2158_n5888# 0.02107f
C589 source.n493 a_n2158_n5888# 0.011322f
C590 source.n494 a_n2158_n5888# 0.011988f
C591 source.n495 a_n2158_n5888# 0.026761f
C592 source.n496 a_n2158_n5888# 0.026761f
C593 source.n497 a_n2158_n5888# 0.026761f
C594 source.n498 a_n2158_n5888# 0.011655f
C595 source.n499 a_n2158_n5888# 0.011322f
C596 source.n500 a_n2158_n5888# 0.02107f
C597 source.n501 a_n2158_n5888# 0.02107f
C598 source.n502 a_n2158_n5888# 0.011322f
C599 source.n503 a_n2158_n5888# 0.011988f
C600 source.n504 a_n2158_n5888# 0.026761f
C601 source.n505 a_n2158_n5888# 0.026761f
C602 source.n506 a_n2158_n5888# 0.011988f
C603 source.n507 a_n2158_n5888# 0.011322f
C604 source.n508 a_n2158_n5888# 0.02107f
C605 source.n509 a_n2158_n5888# 0.02107f
C606 source.n510 a_n2158_n5888# 0.011322f
C607 source.n511 a_n2158_n5888# 0.011988f
C608 source.n512 a_n2158_n5888# 0.026761f
C609 source.n513 a_n2158_n5888# 0.026761f
C610 source.n514 a_n2158_n5888# 0.011988f
C611 source.n515 a_n2158_n5888# 0.011322f
C612 source.n516 a_n2158_n5888# 0.02107f
C613 source.n517 a_n2158_n5888# 0.02107f
C614 source.n518 a_n2158_n5888# 0.011322f
C615 source.n519 a_n2158_n5888# 0.011988f
C616 source.n520 a_n2158_n5888# 0.026761f
C617 source.n521 a_n2158_n5888# 0.026761f
C618 source.n522 a_n2158_n5888# 0.011988f
C619 source.n523 a_n2158_n5888# 0.011322f
C620 source.n524 a_n2158_n5888# 0.02107f
C621 source.n525 a_n2158_n5888# 0.02107f
C622 source.n526 a_n2158_n5888# 0.011322f
C623 source.n527 a_n2158_n5888# 0.011988f
C624 source.n528 a_n2158_n5888# 0.026761f
C625 source.n529 a_n2158_n5888# 0.026761f
C626 source.n530 a_n2158_n5888# 0.011988f
C627 source.n531 a_n2158_n5888# 0.011322f
C628 source.n532 a_n2158_n5888# 0.02107f
C629 source.n533 a_n2158_n5888# 0.02107f
C630 source.n534 a_n2158_n5888# 0.011322f
C631 source.n535 a_n2158_n5888# 0.011988f
C632 source.n536 a_n2158_n5888# 0.026761f
C633 source.n537 a_n2158_n5888# 0.026761f
C634 source.n538 a_n2158_n5888# 0.011988f
C635 source.n539 a_n2158_n5888# 0.011322f
C636 source.n540 a_n2158_n5888# 0.02107f
C637 source.n541 a_n2158_n5888# 0.02107f
C638 source.n542 a_n2158_n5888# 0.011322f
C639 source.n543 a_n2158_n5888# 0.011655f
C640 source.n544 a_n2158_n5888# 0.011655f
C641 source.n545 a_n2158_n5888# 0.026761f
C642 source.n546 a_n2158_n5888# 0.026761f
C643 source.n547 a_n2158_n5888# 0.011988f
C644 source.n548 a_n2158_n5888# 0.011322f
C645 source.n549 a_n2158_n5888# 0.02107f
C646 source.n550 a_n2158_n5888# 0.02107f
C647 source.n551 a_n2158_n5888# 0.011322f
C648 source.n552 a_n2158_n5888# 0.011988f
C649 source.n553 a_n2158_n5888# 0.026761f
C650 source.n554 a_n2158_n5888# 0.026761f
C651 source.n555 a_n2158_n5888# 0.011988f
C652 source.n556 a_n2158_n5888# 0.011322f
C653 source.n557 a_n2158_n5888# 0.02107f
C654 source.n558 a_n2158_n5888# 0.02107f
C655 source.n559 a_n2158_n5888# 0.011322f
C656 source.n560 a_n2158_n5888# 0.011988f
C657 source.n561 a_n2158_n5888# 0.026761f
C658 source.n562 a_n2158_n5888# 0.056928f
C659 source.n563 a_n2158_n5888# 0.011988f
C660 source.n564 a_n2158_n5888# 0.011322f
C661 source.n565 a_n2158_n5888# 0.0464f
C662 source.n566 a_n2158_n5888# 0.031678f
C663 source.n567 a_n2158_n5888# 2.09254f
C664 source.n568 a_n2158_n5888# 0.029047f
C665 source.n569 a_n2158_n5888# 0.02107f
C666 source.n570 a_n2158_n5888# 0.011322f
C667 source.n571 a_n2158_n5888# 0.026761f
C668 source.n572 a_n2158_n5888# 0.011988f
C669 source.n573 a_n2158_n5888# 0.02107f
C670 source.n574 a_n2158_n5888# 0.011322f
C671 source.n575 a_n2158_n5888# 0.026761f
C672 source.n576 a_n2158_n5888# 0.011988f
C673 source.n577 a_n2158_n5888# 0.02107f
C674 source.n578 a_n2158_n5888# 0.011322f
C675 source.n579 a_n2158_n5888# 0.026761f
C676 source.n580 a_n2158_n5888# 0.011988f
C677 source.n581 a_n2158_n5888# 0.02107f
C678 source.n582 a_n2158_n5888# 0.011322f
C679 source.n583 a_n2158_n5888# 0.026761f
C680 source.n584 a_n2158_n5888# 0.011988f
C681 source.n585 a_n2158_n5888# 0.02107f
C682 source.n586 a_n2158_n5888# 0.011322f
C683 source.n587 a_n2158_n5888# 0.026761f
C684 source.n588 a_n2158_n5888# 0.011988f
C685 source.n589 a_n2158_n5888# 0.02107f
C686 source.n590 a_n2158_n5888# 0.011322f
C687 source.n591 a_n2158_n5888# 0.026761f
C688 source.n592 a_n2158_n5888# 0.011988f
C689 source.n593 a_n2158_n5888# 0.02107f
C690 source.n594 a_n2158_n5888# 0.011322f
C691 source.n595 a_n2158_n5888# 0.026761f
C692 source.n596 a_n2158_n5888# 0.011988f
C693 source.n597 a_n2158_n5888# 0.02107f
C694 source.n598 a_n2158_n5888# 0.011322f
C695 source.n599 a_n2158_n5888# 0.026761f
C696 source.n600 a_n2158_n5888# 0.011988f
C697 source.n601 a_n2158_n5888# 0.02107f
C698 source.n602 a_n2158_n5888# 0.011655f
C699 source.n603 a_n2158_n5888# 0.026761f
C700 source.n604 a_n2158_n5888# 0.011988f
C701 source.n605 a_n2158_n5888# 0.02107f
C702 source.n606 a_n2158_n5888# 0.011322f
C703 source.n607 a_n2158_n5888# 0.026761f
C704 source.n608 a_n2158_n5888# 0.011988f
C705 source.n609 a_n2158_n5888# 0.02107f
C706 source.n610 a_n2158_n5888# 0.011322f
C707 source.n611 a_n2158_n5888# 0.020071f
C708 source.n612 a_n2158_n5888# 0.018918f
C709 source.t2 a_n2158_n5888# 0.046673f
C710 source.n613 a_n2158_n5888# 0.257071f
C711 source.n614 a_n2158_n5888# 2.28126f
C712 source.n615 a_n2158_n5888# 0.011322f
C713 source.n616 a_n2158_n5888# 0.011988f
C714 source.n617 a_n2158_n5888# 0.026761f
C715 source.n618 a_n2158_n5888# 0.026761f
C716 source.n619 a_n2158_n5888# 0.011988f
C717 source.n620 a_n2158_n5888# 0.011322f
C718 source.n621 a_n2158_n5888# 0.02107f
C719 source.n622 a_n2158_n5888# 0.02107f
C720 source.n623 a_n2158_n5888# 0.011322f
C721 source.n624 a_n2158_n5888# 0.011988f
C722 source.n625 a_n2158_n5888# 0.026761f
C723 source.n626 a_n2158_n5888# 0.026761f
C724 source.n627 a_n2158_n5888# 0.011988f
C725 source.n628 a_n2158_n5888# 0.011322f
C726 source.n629 a_n2158_n5888# 0.02107f
C727 source.n630 a_n2158_n5888# 0.02107f
C728 source.n631 a_n2158_n5888# 0.011322f
C729 source.n632 a_n2158_n5888# 0.011322f
C730 source.n633 a_n2158_n5888# 0.011988f
C731 source.n634 a_n2158_n5888# 0.026761f
C732 source.n635 a_n2158_n5888# 0.026761f
C733 source.n636 a_n2158_n5888# 0.026761f
C734 source.n637 a_n2158_n5888# 0.011655f
C735 source.n638 a_n2158_n5888# 0.011322f
C736 source.n639 a_n2158_n5888# 0.02107f
C737 source.n640 a_n2158_n5888# 0.02107f
C738 source.n641 a_n2158_n5888# 0.011322f
C739 source.n642 a_n2158_n5888# 0.011988f
C740 source.n643 a_n2158_n5888# 0.026761f
C741 source.n644 a_n2158_n5888# 0.026761f
C742 source.n645 a_n2158_n5888# 0.011988f
C743 source.n646 a_n2158_n5888# 0.011322f
C744 source.n647 a_n2158_n5888# 0.02107f
C745 source.n648 a_n2158_n5888# 0.02107f
C746 source.n649 a_n2158_n5888# 0.011322f
C747 source.n650 a_n2158_n5888# 0.011988f
C748 source.n651 a_n2158_n5888# 0.026761f
C749 source.n652 a_n2158_n5888# 0.026761f
C750 source.n653 a_n2158_n5888# 0.011988f
C751 source.n654 a_n2158_n5888# 0.011322f
C752 source.n655 a_n2158_n5888# 0.02107f
C753 source.n656 a_n2158_n5888# 0.02107f
C754 source.n657 a_n2158_n5888# 0.011322f
C755 source.n658 a_n2158_n5888# 0.011988f
C756 source.n659 a_n2158_n5888# 0.026761f
C757 source.n660 a_n2158_n5888# 0.026761f
C758 source.n661 a_n2158_n5888# 0.011988f
C759 source.n662 a_n2158_n5888# 0.011322f
C760 source.n663 a_n2158_n5888# 0.02107f
C761 source.n664 a_n2158_n5888# 0.02107f
C762 source.n665 a_n2158_n5888# 0.011322f
C763 source.n666 a_n2158_n5888# 0.011988f
C764 source.n667 a_n2158_n5888# 0.026761f
C765 source.n668 a_n2158_n5888# 0.026761f
C766 source.n669 a_n2158_n5888# 0.011988f
C767 source.n670 a_n2158_n5888# 0.011322f
C768 source.n671 a_n2158_n5888# 0.02107f
C769 source.n672 a_n2158_n5888# 0.02107f
C770 source.n673 a_n2158_n5888# 0.011322f
C771 source.n674 a_n2158_n5888# 0.011988f
C772 source.n675 a_n2158_n5888# 0.026761f
C773 source.n676 a_n2158_n5888# 0.026761f
C774 source.n677 a_n2158_n5888# 0.026761f
C775 source.n678 a_n2158_n5888# 0.011988f
C776 source.n679 a_n2158_n5888# 0.011322f
C777 source.n680 a_n2158_n5888# 0.02107f
C778 source.n681 a_n2158_n5888# 0.02107f
C779 source.n682 a_n2158_n5888# 0.011322f
C780 source.n683 a_n2158_n5888# 0.011655f
C781 source.n684 a_n2158_n5888# 0.011655f
C782 source.n685 a_n2158_n5888# 0.026761f
C783 source.n686 a_n2158_n5888# 0.026761f
C784 source.n687 a_n2158_n5888# 0.011988f
C785 source.n688 a_n2158_n5888# 0.011322f
C786 source.n689 a_n2158_n5888# 0.02107f
C787 source.n690 a_n2158_n5888# 0.02107f
C788 source.n691 a_n2158_n5888# 0.011322f
C789 source.n692 a_n2158_n5888# 0.011988f
C790 source.n693 a_n2158_n5888# 0.026761f
C791 source.n694 a_n2158_n5888# 0.026761f
C792 source.n695 a_n2158_n5888# 0.011988f
C793 source.n696 a_n2158_n5888# 0.011322f
C794 source.n697 a_n2158_n5888# 0.02107f
C795 source.n698 a_n2158_n5888# 0.02107f
C796 source.n699 a_n2158_n5888# 0.011322f
C797 source.n700 a_n2158_n5888# 0.011988f
C798 source.n701 a_n2158_n5888# 0.026761f
C799 source.n702 a_n2158_n5888# 0.056928f
C800 source.n703 a_n2158_n5888# 0.011988f
C801 source.n704 a_n2158_n5888# 0.011322f
C802 source.n705 a_n2158_n5888# 0.0464f
C803 source.n706 a_n2158_n5888# 0.031678f
C804 source.n707 a_n2158_n5888# 2.09254f
C805 source.t8 a_n2158_n5888# 0.416253f
C806 source.t3 a_n2158_n5888# 0.416253f
C807 source.n708 a_n2158_n5888# 3.76715f
C808 source.n709 a_n2158_n5888# 0.339106f
C809 source.t4 a_n2158_n5888# 0.416253f
C810 source.t21 a_n2158_n5888# 0.416253f
C811 source.n710 a_n2158_n5888# 3.76715f
C812 source.n711 a_n2158_n5888# 0.339106f
C813 source.n712 a_n2158_n5888# 0.029047f
C814 source.n713 a_n2158_n5888# 0.02107f
C815 source.n714 a_n2158_n5888# 0.011322f
C816 source.n715 a_n2158_n5888# 0.026761f
C817 source.n716 a_n2158_n5888# 0.011988f
C818 source.n717 a_n2158_n5888# 0.02107f
C819 source.n718 a_n2158_n5888# 0.011322f
C820 source.n719 a_n2158_n5888# 0.026761f
C821 source.n720 a_n2158_n5888# 0.011988f
C822 source.n721 a_n2158_n5888# 0.02107f
C823 source.n722 a_n2158_n5888# 0.011322f
C824 source.n723 a_n2158_n5888# 0.026761f
C825 source.n724 a_n2158_n5888# 0.011988f
C826 source.n725 a_n2158_n5888# 0.02107f
C827 source.n726 a_n2158_n5888# 0.011322f
C828 source.n727 a_n2158_n5888# 0.026761f
C829 source.n728 a_n2158_n5888# 0.011988f
C830 source.n729 a_n2158_n5888# 0.02107f
C831 source.n730 a_n2158_n5888# 0.011322f
C832 source.n731 a_n2158_n5888# 0.026761f
C833 source.n732 a_n2158_n5888# 0.011988f
C834 source.n733 a_n2158_n5888# 0.02107f
C835 source.n734 a_n2158_n5888# 0.011322f
C836 source.n735 a_n2158_n5888# 0.026761f
C837 source.n736 a_n2158_n5888# 0.011988f
C838 source.n737 a_n2158_n5888# 0.02107f
C839 source.n738 a_n2158_n5888# 0.011322f
C840 source.n739 a_n2158_n5888# 0.026761f
C841 source.n740 a_n2158_n5888# 0.011988f
C842 source.n741 a_n2158_n5888# 0.02107f
C843 source.n742 a_n2158_n5888# 0.011322f
C844 source.n743 a_n2158_n5888# 0.026761f
C845 source.n744 a_n2158_n5888# 0.011988f
C846 source.n745 a_n2158_n5888# 0.02107f
C847 source.n746 a_n2158_n5888# 0.011655f
C848 source.n747 a_n2158_n5888# 0.026761f
C849 source.n748 a_n2158_n5888# 0.011988f
C850 source.n749 a_n2158_n5888# 0.02107f
C851 source.n750 a_n2158_n5888# 0.011322f
C852 source.n751 a_n2158_n5888# 0.026761f
C853 source.n752 a_n2158_n5888# 0.011988f
C854 source.n753 a_n2158_n5888# 0.02107f
C855 source.n754 a_n2158_n5888# 0.011322f
C856 source.n755 a_n2158_n5888# 0.020071f
C857 source.n756 a_n2158_n5888# 0.018918f
C858 source.t6 a_n2158_n5888# 0.046673f
C859 source.n757 a_n2158_n5888# 0.257071f
C860 source.n758 a_n2158_n5888# 2.28126f
C861 source.n759 a_n2158_n5888# 0.011322f
C862 source.n760 a_n2158_n5888# 0.011988f
C863 source.n761 a_n2158_n5888# 0.026761f
C864 source.n762 a_n2158_n5888# 0.026761f
C865 source.n763 a_n2158_n5888# 0.011988f
C866 source.n764 a_n2158_n5888# 0.011322f
C867 source.n765 a_n2158_n5888# 0.02107f
C868 source.n766 a_n2158_n5888# 0.02107f
C869 source.n767 a_n2158_n5888# 0.011322f
C870 source.n768 a_n2158_n5888# 0.011988f
C871 source.n769 a_n2158_n5888# 0.026761f
C872 source.n770 a_n2158_n5888# 0.026761f
C873 source.n771 a_n2158_n5888# 0.011988f
C874 source.n772 a_n2158_n5888# 0.011322f
C875 source.n773 a_n2158_n5888# 0.02107f
C876 source.n774 a_n2158_n5888# 0.02107f
C877 source.n775 a_n2158_n5888# 0.011322f
C878 source.n776 a_n2158_n5888# 0.011322f
C879 source.n777 a_n2158_n5888# 0.011988f
C880 source.n778 a_n2158_n5888# 0.026761f
C881 source.n779 a_n2158_n5888# 0.026761f
C882 source.n780 a_n2158_n5888# 0.026761f
C883 source.n781 a_n2158_n5888# 0.011655f
C884 source.n782 a_n2158_n5888# 0.011322f
C885 source.n783 a_n2158_n5888# 0.02107f
C886 source.n784 a_n2158_n5888# 0.02107f
C887 source.n785 a_n2158_n5888# 0.011322f
C888 source.n786 a_n2158_n5888# 0.011988f
C889 source.n787 a_n2158_n5888# 0.026761f
C890 source.n788 a_n2158_n5888# 0.026761f
C891 source.n789 a_n2158_n5888# 0.011988f
C892 source.n790 a_n2158_n5888# 0.011322f
C893 source.n791 a_n2158_n5888# 0.02107f
C894 source.n792 a_n2158_n5888# 0.02107f
C895 source.n793 a_n2158_n5888# 0.011322f
C896 source.n794 a_n2158_n5888# 0.011988f
C897 source.n795 a_n2158_n5888# 0.026761f
C898 source.n796 a_n2158_n5888# 0.026761f
C899 source.n797 a_n2158_n5888# 0.011988f
C900 source.n798 a_n2158_n5888# 0.011322f
C901 source.n799 a_n2158_n5888# 0.02107f
C902 source.n800 a_n2158_n5888# 0.02107f
C903 source.n801 a_n2158_n5888# 0.011322f
C904 source.n802 a_n2158_n5888# 0.011988f
C905 source.n803 a_n2158_n5888# 0.026761f
C906 source.n804 a_n2158_n5888# 0.026761f
C907 source.n805 a_n2158_n5888# 0.011988f
C908 source.n806 a_n2158_n5888# 0.011322f
C909 source.n807 a_n2158_n5888# 0.02107f
C910 source.n808 a_n2158_n5888# 0.02107f
C911 source.n809 a_n2158_n5888# 0.011322f
C912 source.n810 a_n2158_n5888# 0.011988f
C913 source.n811 a_n2158_n5888# 0.026761f
C914 source.n812 a_n2158_n5888# 0.026761f
C915 source.n813 a_n2158_n5888# 0.011988f
C916 source.n814 a_n2158_n5888# 0.011322f
C917 source.n815 a_n2158_n5888# 0.02107f
C918 source.n816 a_n2158_n5888# 0.02107f
C919 source.n817 a_n2158_n5888# 0.011322f
C920 source.n818 a_n2158_n5888# 0.011988f
C921 source.n819 a_n2158_n5888# 0.026761f
C922 source.n820 a_n2158_n5888# 0.026761f
C923 source.n821 a_n2158_n5888# 0.026761f
C924 source.n822 a_n2158_n5888# 0.011988f
C925 source.n823 a_n2158_n5888# 0.011322f
C926 source.n824 a_n2158_n5888# 0.02107f
C927 source.n825 a_n2158_n5888# 0.02107f
C928 source.n826 a_n2158_n5888# 0.011322f
C929 source.n827 a_n2158_n5888# 0.011655f
C930 source.n828 a_n2158_n5888# 0.011655f
C931 source.n829 a_n2158_n5888# 0.026761f
C932 source.n830 a_n2158_n5888# 0.026761f
C933 source.n831 a_n2158_n5888# 0.011988f
C934 source.n832 a_n2158_n5888# 0.011322f
C935 source.n833 a_n2158_n5888# 0.02107f
C936 source.n834 a_n2158_n5888# 0.02107f
C937 source.n835 a_n2158_n5888# 0.011322f
C938 source.n836 a_n2158_n5888# 0.011988f
C939 source.n837 a_n2158_n5888# 0.026761f
C940 source.n838 a_n2158_n5888# 0.026761f
C941 source.n839 a_n2158_n5888# 0.011988f
C942 source.n840 a_n2158_n5888# 0.011322f
C943 source.n841 a_n2158_n5888# 0.02107f
C944 source.n842 a_n2158_n5888# 0.02107f
C945 source.n843 a_n2158_n5888# 0.011322f
C946 source.n844 a_n2158_n5888# 0.011988f
C947 source.n845 a_n2158_n5888# 0.026761f
C948 source.n846 a_n2158_n5888# 0.056928f
C949 source.n847 a_n2158_n5888# 0.011988f
C950 source.n848 a_n2158_n5888# 0.011322f
C951 source.n849 a_n2158_n5888# 0.0464f
C952 source.n850 a_n2158_n5888# 0.031678f
C953 source.n851 a_n2158_n5888# 0.108878f
C954 source.n852 a_n2158_n5888# 0.029047f
C955 source.n853 a_n2158_n5888# 0.02107f
C956 source.n854 a_n2158_n5888# 0.011322f
C957 source.n855 a_n2158_n5888# 0.026761f
C958 source.n856 a_n2158_n5888# 0.011988f
C959 source.n857 a_n2158_n5888# 0.02107f
C960 source.n858 a_n2158_n5888# 0.011322f
C961 source.n859 a_n2158_n5888# 0.026761f
C962 source.n860 a_n2158_n5888# 0.011988f
C963 source.n861 a_n2158_n5888# 0.02107f
C964 source.n862 a_n2158_n5888# 0.011322f
C965 source.n863 a_n2158_n5888# 0.026761f
C966 source.n864 a_n2158_n5888# 0.011988f
C967 source.n865 a_n2158_n5888# 0.02107f
C968 source.n866 a_n2158_n5888# 0.011322f
C969 source.n867 a_n2158_n5888# 0.026761f
C970 source.n868 a_n2158_n5888# 0.011988f
C971 source.n869 a_n2158_n5888# 0.02107f
C972 source.n870 a_n2158_n5888# 0.011322f
C973 source.n871 a_n2158_n5888# 0.026761f
C974 source.n872 a_n2158_n5888# 0.011988f
C975 source.n873 a_n2158_n5888# 0.02107f
C976 source.n874 a_n2158_n5888# 0.011322f
C977 source.n875 a_n2158_n5888# 0.026761f
C978 source.n876 a_n2158_n5888# 0.011988f
C979 source.n877 a_n2158_n5888# 0.02107f
C980 source.n878 a_n2158_n5888# 0.011322f
C981 source.n879 a_n2158_n5888# 0.026761f
C982 source.n880 a_n2158_n5888# 0.011988f
C983 source.n881 a_n2158_n5888# 0.02107f
C984 source.n882 a_n2158_n5888# 0.011322f
C985 source.n883 a_n2158_n5888# 0.026761f
C986 source.n884 a_n2158_n5888# 0.011988f
C987 source.n885 a_n2158_n5888# 0.02107f
C988 source.n886 a_n2158_n5888# 0.011655f
C989 source.n887 a_n2158_n5888# 0.026761f
C990 source.n888 a_n2158_n5888# 0.011988f
C991 source.n889 a_n2158_n5888# 0.02107f
C992 source.n890 a_n2158_n5888# 0.011322f
C993 source.n891 a_n2158_n5888# 0.026761f
C994 source.n892 a_n2158_n5888# 0.011988f
C995 source.n893 a_n2158_n5888# 0.02107f
C996 source.n894 a_n2158_n5888# 0.011322f
C997 source.n895 a_n2158_n5888# 0.020071f
C998 source.n896 a_n2158_n5888# 0.018918f
C999 source.t15 a_n2158_n5888# 0.046673f
C1000 source.n897 a_n2158_n5888# 0.257071f
C1001 source.n898 a_n2158_n5888# 2.28126f
C1002 source.n899 a_n2158_n5888# 0.011322f
C1003 source.n900 a_n2158_n5888# 0.011988f
C1004 source.n901 a_n2158_n5888# 0.026761f
C1005 source.n902 a_n2158_n5888# 0.026761f
C1006 source.n903 a_n2158_n5888# 0.011988f
C1007 source.n904 a_n2158_n5888# 0.011322f
C1008 source.n905 a_n2158_n5888# 0.02107f
C1009 source.n906 a_n2158_n5888# 0.02107f
C1010 source.n907 a_n2158_n5888# 0.011322f
C1011 source.n908 a_n2158_n5888# 0.011988f
C1012 source.n909 a_n2158_n5888# 0.026761f
C1013 source.n910 a_n2158_n5888# 0.026761f
C1014 source.n911 a_n2158_n5888# 0.011988f
C1015 source.n912 a_n2158_n5888# 0.011322f
C1016 source.n913 a_n2158_n5888# 0.02107f
C1017 source.n914 a_n2158_n5888# 0.02107f
C1018 source.n915 a_n2158_n5888# 0.011322f
C1019 source.n916 a_n2158_n5888# 0.011322f
C1020 source.n917 a_n2158_n5888# 0.011988f
C1021 source.n918 a_n2158_n5888# 0.026761f
C1022 source.n919 a_n2158_n5888# 0.026761f
C1023 source.n920 a_n2158_n5888# 0.026761f
C1024 source.n921 a_n2158_n5888# 0.011655f
C1025 source.n922 a_n2158_n5888# 0.011322f
C1026 source.n923 a_n2158_n5888# 0.02107f
C1027 source.n924 a_n2158_n5888# 0.02107f
C1028 source.n925 a_n2158_n5888# 0.011322f
C1029 source.n926 a_n2158_n5888# 0.011988f
C1030 source.n927 a_n2158_n5888# 0.026761f
C1031 source.n928 a_n2158_n5888# 0.026761f
C1032 source.n929 a_n2158_n5888# 0.011988f
C1033 source.n930 a_n2158_n5888# 0.011322f
C1034 source.n931 a_n2158_n5888# 0.02107f
C1035 source.n932 a_n2158_n5888# 0.02107f
C1036 source.n933 a_n2158_n5888# 0.011322f
C1037 source.n934 a_n2158_n5888# 0.011988f
C1038 source.n935 a_n2158_n5888# 0.026761f
C1039 source.n936 a_n2158_n5888# 0.026761f
C1040 source.n937 a_n2158_n5888# 0.011988f
C1041 source.n938 a_n2158_n5888# 0.011322f
C1042 source.n939 a_n2158_n5888# 0.02107f
C1043 source.n940 a_n2158_n5888# 0.02107f
C1044 source.n941 a_n2158_n5888# 0.011322f
C1045 source.n942 a_n2158_n5888# 0.011988f
C1046 source.n943 a_n2158_n5888# 0.026761f
C1047 source.n944 a_n2158_n5888# 0.026761f
C1048 source.n945 a_n2158_n5888# 0.011988f
C1049 source.n946 a_n2158_n5888# 0.011322f
C1050 source.n947 a_n2158_n5888# 0.02107f
C1051 source.n948 a_n2158_n5888# 0.02107f
C1052 source.n949 a_n2158_n5888# 0.011322f
C1053 source.n950 a_n2158_n5888# 0.011988f
C1054 source.n951 a_n2158_n5888# 0.026761f
C1055 source.n952 a_n2158_n5888# 0.026761f
C1056 source.n953 a_n2158_n5888# 0.011988f
C1057 source.n954 a_n2158_n5888# 0.011322f
C1058 source.n955 a_n2158_n5888# 0.02107f
C1059 source.n956 a_n2158_n5888# 0.02107f
C1060 source.n957 a_n2158_n5888# 0.011322f
C1061 source.n958 a_n2158_n5888# 0.011988f
C1062 source.n959 a_n2158_n5888# 0.026761f
C1063 source.n960 a_n2158_n5888# 0.026761f
C1064 source.n961 a_n2158_n5888# 0.026761f
C1065 source.n962 a_n2158_n5888# 0.011988f
C1066 source.n963 a_n2158_n5888# 0.011322f
C1067 source.n964 a_n2158_n5888# 0.02107f
C1068 source.n965 a_n2158_n5888# 0.02107f
C1069 source.n966 a_n2158_n5888# 0.011322f
C1070 source.n967 a_n2158_n5888# 0.011655f
C1071 source.n968 a_n2158_n5888# 0.011655f
C1072 source.n969 a_n2158_n5888# 0.026761f
C1073 source.n970 a_n2158_n5888# 0.026761f
C1074 source.n971 a_n2158_n5888# 0.011988f
C1075 source.n972 a_n2158_n5888# 0.011322f
C1076 source.n973 a_n2158_n5888# 0.02107f
C1077 source.n974 a_n2158_n5888# 0.02107f
C1078 source.n975 a_n2158_n5888# 0.011322f
C1079 source.n976 a_n2158_n5888# 0.011988f
C1080 source.n977 a_n2158_n5888# 0.026761f
C1081 source.n978 a_n2158_n5888# 0.026761f
C1082 source.n979 a_n2158_n5888# 0.011988f
C1083 source.n980 a_n2158_n5888# 0.011322f
C1084 source.n981 a_n2158_n5888# 0.02107f
C1085 source.n982 a_n2158_n5888# 0.02107f
C1086 source.n983 a_n2158_n5888# 0.011322f
C1087 source.n984 a_n2158_n5888# 0.011988f
C1088 source.n985 a_n2158_n5888# 0.026761f
C1089 source.n986 a_n2158_n5888# 0.056928f
C1090 source.n987 a_n2158_n5888# 0.011988f
C1091 source.n988 a_n2158_n5888# 0.011322f
C1092 source.n989 a_n2158_n5888# 0.0464f
C1093 source.n990 a_n2158_n5888# 0.031678f
C1094 source.n991 a_n2158_n5888# 0.108878f
C1095 source.t16 a_n2158_n5888# 0.416253f
C1096 source.t20 a_n2158_n5888# 0.416253f
C1097 source.n992 a_n2158_n5888# 3.76715f
C1098 source.n993 a_n2158_n5888# 0.339106f
C1099 source.t19 a_n2158_n5888# 0.416253f
C1100 source.t17 a_n2158_n5888# 0.416253f
C1101 source.n994 a_n2158_n5888# 3.76715f
C1102 source.n995 a_n2158_n5888# 0.339106f
C1103 source.n996 a_n2158_n5888# 0.029047f
C1104 source.n997 a_n2158_n5888# 0.02107f
C1105 source.n998 a_n2158_n5888# 0.011322f
C1106 source.n999 a_n2158_n5888# 0.026761f
C1107 source.n1000 a_n2158_n5888# 0.011988f
C1108 source.n1001 a_n2158_n5888# 0.02107f
C1109 source.n1002 a_n2158_n5888# 0.011322f
C1110 source.n1003 a_n2158_n5888# 0.026761f
C1111 source.n1004 a_n2158_n5888# 0.011988f
C1112 source.n1005 a_n2158_n5888# 0.02107f
C1113 source.n1006 a_n2158_n5888# 0.011322f
C1114 source.n1007 a_n2158_n5888# 0.026761f
C1115 source.n1008 a_n2158_n5888# 0.011988f
C1116 source.n1009 a_n2158_n5888# 0.02107f
C1117 source.n1010 a_n2158_n5888# 0.011322f
C1118 source.n1011 a_n2158_n5888# 0.026761f
C1119 source.n1012 a_n2158_n5888# 0.011988f
C1120 source.n1013 a_n2158_n5888# 0.02107f
C1121 source.n1014 a_n2158_n5888# 0.011322f
C1122 source.n1015 a_n2158_n5888# 0.026761f
C1123 source.n1016 a_n2158_n5888# 0.011988f
C1124 source.n1017 a_n2158_n5888# 0.02107f
C1125 source.n1018 a_n2158_n5888# 0.011322f
C1126 source.n1019 a_n2158_n5888# 0.026761f
C1127 source.n1020 a_n2158_n5888# 0.011988f
C1128 source.n1021 a_n2158_n5888# 0.02107f
C1129 source.n1022 a_n2158_n5888# 0.011322f
C1130 source.n1023 a_n2158_n5888# 0.026761f
C1131 source.n1024 a_n2158_n5888# 0.011988f
C1132 source.n1025 a_n2158_n5888# 0.02107f
C1133 source.n1026 a_n2158_n5888# 0.011322f
C1134 source.n1027 a_n2158_n5888# 0.026761f
C1135 source.n1028 a_n2158_n5888# 0.011988f
C1136 source.n1029 a_n2158_n5888# 0.02107f
C1137 source.n1030 a_n2158_n5888# 0.011655f
C1138 source.n1031 a_n2158_n5888# 0.026761f
C1139 source.n1032 a_n2158_n5888# 0.011988f
C1140 source.n1033 a_n2158_n5888# 0.02107f
C1141 source.n1034 a_n2158_n5888# 0.011322f
C1142 source.n1035 a_n2158_n5888# 0.026761f
C1143 source.n1036 a_n2158_n5888# 0.011988f
C1144 source.n1037 a_n2158_n5888# 0.02107f
C1145 source.n1038 a_n2158_n5888# 0.011322f
C1146 source.n1039 a_n2158_n5888# 0.020071f
C1147 source.n1040 a_n2158_n5888# 0.018918f
C1148 source.t11 a_n2158_n5888# 0.046673f
C1149 source.n1041 a_n2158_n5888# 0.257071f
C1150 source.n1042 a_n2158_n5888# 2.28126f
C1151 source.n1043 a_n2158_n5888# 0.011322f
C1152 source.n1044 a_n2158_n5888# 0.011988f
C1153 source.n1045 a_n2158_n5888# 0.026761f
C1154 source.n1046 a_n2158_n5888# 0.026761f
C1155 source.n1047 a_n2158_n5888# 0.011988f
C1156 source.n1048 a_n2158_n5888# 0.011322f
C1157 source.n1049 a_n2158_n5888# 0.02107f
C1158 source.n1050 a_n2158_n5888# 0.02107f
C1159 source.n1051 a_n2158_n5888# 0.011322f
C1160 source.n1052 a_n2158_n5888# 0.011988f
C1161 source.n1053 a_n2158_n5888# 0.026761f
C1162 source.n1054 a_n2158_n5888# 0.026761f
C1163 source.n1055 a_n2158_n5888# 0.011988f
C1164 source.n1056 a_n2158_n5888# 0.011322f
C1165 source.n1057 a_n2158_n5888# 0.02107f
C1166 source.n1058 a_n2158_n5888# 0.02107f
C1167 source.n1059 a_n2158_n5888# 0.011322f
C1168 source.n1060 a_n2158_n5888# 0.011322f
C1169 source.n1061 a_n2158_n5888# 0.011988f
C1170 source.n1062 a_n2158_n5888# 0.026761f
C1171 source.n1063 a_n2158_n5888# 0.026761f
C1172 source.n1064 a_n2158_n5888# 0.026761f
C1173 source.n1065 a_n2158_n5888# 0.011655f
C1174 source.n1066 a_n2158_n5888# 0.011322f
C1175 source.n1067 a_n2158_n5888# 0.02107f
C1176 source.n1068 a_n2158_n5888# 0.02107f
C1177 source.n1069 a_n2158_n5888# 0.011322f
C1178 source.n1070 a_n2158_n5888# 0.011988f
C1179 source.n1071 a_n2158_n5888# 0.026761f
C1180 source.n1072 a_n2158_n5888# 0.026761f
C1181 source.n1073 a_n2158_n5888# 0.011988f
C1182 source.n1074 a_n2158_n5888# 0.011322f
C1183 source.n1075 a_n2158_n5888# 0.02107f
C1184 source.n1076 a_n2158_n5888# 0.02107f
C1185 source.n1077 a_n2158_n5888# 0.011322f
C1186 source.n1078 a_n2158_n5888# 0.011988f
C1187 source.n1079 a_n2158_n5888# 0.026761f
C1188 source.n1080 a_n2158_n5888# 0.026761f
C1189 source.n1081 a_n2158_n5888# 0.011988f
C1190 source.n1082 a_n2158_n5888# 0.011322f
C1191 source.n1083 a_n2158_n5888# 0.02107f
C1192 source.n1084 a_n2158_n5888# 0.02107f
C1193 source.n1085 a_n2158_n5888# 0.011322f
C1194 source.n1086 a_n2158_n5888# 0.011988f
C1195 source.n1087 a_n2158_n5888# 0.026761f
C1196 source.n1088 a_n2158_n5888# 0.026761f
C1197 source.n1089 a_n2158_n5888# 0.011988f
C1198 source.n1090 a_n2158_n5888# 0.011322f
C1199 source.n1091 a_n2158_n5888# 0.02107f
C1200 source.n1092 a_n2158_n5888# 0.02107f
C1201 source.n1093 a_n2158_n5888# 0.011322f
C1202 source.n1094 a_n2158_n5888# 0.011988f
C1203 source.n1095 a_n2158_n5888# 0.026761f
C1204 source.n1096 a_n2158_n5888# 0.026761f
C1205 source.n1097 a_n2158_n5888# 0.011988f
C1206 source.n1098 a_n2158_n5888# 0.011322f
C1207 source.n1099 a_n2158_n5888# 0.02107f
C1208 source.n1100 a_n2158_n5888# 0.02107f
C1209 source.n1101 a_n2158_n5888# 0.011322f
C1210 source.n1102 a_n2158_n5888# 0.011988f
C1211 source.n1103 a_n2158_n5888# 0.026761f
C1212 source.n1104 a_n2158_n5888# 0.026761f
C1213 source.n1105 a_n2158_n5888# 0.026761f
C1214 source.n1106 a_n2158_n5888# 0.011988f
C1215 source.n1107 a_n2158_n5888# 0.011322f
C1216 source.n1108 a_n2158_n5888# 0.02107f
C1217 source.n1109 a_n2158_n5888# 0.02107f
C1218 source.n1110 a_n2158_n5888# 0.011322f
C1219 source.n1111 a_n2158_n5888# 0.011655f
C1220 source.n1112 a_n2158_n5888# 0.011655f
C1221 source.n1113 a_n2158_n5888# 0.026761f
C1222 source.n1114 a_n2158_n5888# 0.026761f
C1223 source.n1115 a_n2158_n5888# 0.011988f
C1224 source.n1116 a_n2158_n5888# 0.011322f
C1225 source.n1117 a_n2158_n5888# 0.02107f
C1226 source.n1118 a_n2158_n5888# 0.02107f
C1227 source.n1119 a_n2158_n5888# 0.011322f
C1228 source.n1120 a_n2158_n5888# 0.011988f
C1229 source.n1121 a_n2158_n5888# 0.026761f
C1230 source.n1122 a_n2158_n5888# 0.026761f
C1231 source.n1123 a_n2158_n5888# 0.011988f
C1232 source.n1124 a_n2158_n5888# 0.011322f
C1233 source.n1125 a_n2158_n5888# 0.02107f
C1234 source.n1126 a_n2158_n5888# 0.02107f
C1235 source.n1127 a_n2158_n5888# 0.011322f
C1236 source.n1128 a_n2158_n5888# 0.011988f
C1237 source.n1129 a_n2158_n5888# 0.026761f
C1238 source.n1130 a_n2158_n5888# 0.056928f
C1239 source.n1131 a_n2158_n5888# 0.011988f
C1240 source.n1132 a_n2158_n5888# 0.011322f
C1241 source.n1133 a_n2158_n5888# 0.0464f
C1242 source.n1134 a_n2158_n5888# 0.031678f
C1243 source.n1135 a_n2158_n5888# 0.246319f
C1244 source.n1136 a_n2158_n5888# 2.26157f
C1245 drain_right.t8 a_n2158_n5888# 0.539531f
C1246 drain_right.t0 a_n2158_n5888# 0.539531f
C1247 drain_right.n0 a_n2158_n5888# 4.97787f
C1248 drain_right.t6 a_n2158_n5888# 0.539531f
C1249 drain_right.t3 a_n2158_n5888# 0.539531f
C1250 drain_right.n1 a_n2158_n5888# 4.97236f
C1251 drain_right.t1 a_n2158_n5888# 0.539531f
C1252 drain_right.t5 a_n2158_n5888# 0.539531f
C1253 drain_right.n2 a_n2158_n5888# 4.97787f
C1254 drain_right.n3 a_n2158_n5888# 3.3775f
C1255 drain_right.t2 a_n2158_n5888# 0.539531f
C1256 drain_right.t9 a_n2158_n5888# 0.539531f
C1257 drain_right.n4 a_n2158_n5888# 4.97828f
C1258 drain_right.t4 a_n2158_n5888# 0.539531f
C1259 drain_right.t10 a_n2158_n5888# 0.539531f
C1260 drain_right.n5 a_n2158_n5888# 4.97236f
C1261 drain_right.n6 a_n2158_n5888# 0.779326f
C1262 drain_right.t11 a_n2158_n5888# 0.539531f
C1263 drain_right.t7 a_n2158_n5888# 0.539531f
C1264 drain_right.n7 a_n2158_n5888# 4.97236f
C1265 drain_right.n8 a_n2158_n5888# 0.628681f
C1266 minus.n0 a_n2158_n5888# 0.041271f
C1267 minus.n1 a_n2158_n5888# 0.009365f
C1268 minus.t6 a_n2158_n5888# 2.04105f
C1269 minus.n2 a_n2158_n5888# 0.041271f
C1270 minus.n3 a_n2158_n5888# 0.009365f
C1271 minus.t7 a_n2158_n5888# 2.04105f
C1272 minus.t8 a_n2158_n5888# 2.05952f
C1273 minus.t2 a_n2158_n5888# 2.04105f
C1274 minus.n4 a_n2158_n5888# 0.749701f
C1275 minus.n5 a_n2158_n5888# 0.730311f
C1276 minus.n6 a_n2158_n5888# 0.173135f
C1277 minus.n7 a_n2158_n5888# 0.041271f
C1278 minus.n8 a_n2158_n5888# 0.745085f
C1279 minus.n9 a_n2158_n5888# 0.009365f
C1280 minus.t10 a_n2158_n5888# 2.04105f
C1281 minus.n10 a_n2158_n5888# 0.745085f
C1282 minus.n11 a_n2158_n5888# 0.041271f
C1283 minus.n12 a_n2158_n5888# 0.041271f
C1284 minus.n13 a_n2158_n5888# 0.041271f
C1285 minus.n14 a_n2158_n5888# 0.745085f
C1286 minus.n15 a_n2158_n5888# 0.009365f
C1287 minus.t11 a_n2158_n5888# 2.04105f
C1288 minus.n16 a_n2158_n5888# 0.743176f
C1289 minus.n17 a_n2158_n5888# 2.17196f
C1290 minus.n18 a_n2158_n5888# 0.041271f
C1291 minus.n19 a_n2158_n5888# 0.009365f
C1292 minus.n20 a_n2158_n5888# 0.041271f
C1293 minus.n21 a_n2158_n5888# 0.009365f
C1294 minus.t5 a_n2158_n5888# 2.05952f
C1295 minus.t4 a_n2158_n5888# 2.04105f
C1296 minus.n22 a_n2158_n5888# 0.749701f
C1297 minus.n23 a_n2158_n5888# 0.730311f
C1298 minus.n24 a_n2158_n5888# 0.173135f
C1299 minus.n25 a_n2158_n5888# 0.041271f
C1300 minus.t0 a_n2158_n5888# 2.04105f
C1301 minus.n26 a_n2158_n5888# 0.745085f
C1302 minus.n27 a_n2158_n5888# 0.009365f
C1303 minus.t1 a_n2158_n5888# 2.04105f
C1304 minus.n28 a_n2158_n5888# 0.745085f
C1305 minus.n29 a_n2158_n5888# 0.041271f
C1306 minus.n30 a_n2158_n5888# 0.041271f
C1307 minus.n31 a_n2158_n5888# 0.041271f
C1308 minus.t3 a_n2158_n5888# 2.04105f
C1309 minus.n32 a_n2158_n5888# 0.745085f
C1310 minus.n33 a_n2158_n5888# 0.009365f
C1311 minus.t9 a_n2158_n5888# 2.04105f
C1312 minus.n34 a_n2158_n5888# 0.743176f
C1313 minus.n35 a_n2158_n5888# 0.283767f
C1314 minus.n36 a_n2158_n5888# 2.55433f
.ends

