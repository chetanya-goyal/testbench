* NGSPICE file created from diffpair97.ext - technology: sky130A

.subckt diffpair97 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t18 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X1 source.t9 minus.t0 drain_right.t15 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X2 drain_right.t14 minus.t1 source.t5 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t17 plus.t1 drain_left.t14 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 drain_right.t13 minus.t2 source.t6 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 drain_right.t12 minus.t3 source.t15 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X6 source.t26 plus.t2 drain_left.t13 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X7 a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X8 drain_right.t11 minus.t4 source.t14 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X9 source.t19 plus.t3 drain_left.t12 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X10 drain_left.t11 plus.t4 source.t20 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X11 drain_left.t10 plus.t5 source.t29 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 source.t10 minus.t5 drain_right.t10 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X13 source.t4 minus.t6 drain_right.t9 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X14 drain_left.t9 plus.t6 source.t25 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X15 source.t24 plus.t7 drain_left.t8 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X16 a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X17 drain_right.t8 minus.t7 source.t8 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X18 source.t22 plus.t8 drain_left.t7 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X19 source.t11 minus.t8 drain_right.t7 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X20 drain_left.t6 plus.t9 source.t31 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X21 drain_right.t6 minus.t9 source.t0 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X22 drain_right.t5 minus.t10 source.t12 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X23 source.t1 minus.t11 drain_right.t4 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X24 source.t21 plus.t10 drain_left.t5 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X25 drain_left.t4 plus.t11 source.t28 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X26 drain_right.t3 minus.t12 source.t7 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X27 source.t30 plus.t12 drain_left.t3 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X28 source.t2 minus.t13 drain_right.t2 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X29 source.t3 minus.t14 drain_right.t1 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X30 source.t13 minus.t15 drain_right.t0 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X31 a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X32 a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X33 drain_left.t2 plus.t13 source.t23 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X34 drain_left.t1 plus.t14 source.t27 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X35 source.t16 plus.t15 drain_left.t0 a_n1670_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 plus.n4 plus.t7 449.502
R1 plus.n17 plus.t14 449.502
R2 plus.n23 plus.t13 449.502
R3 plus.n36 plus.t8 449.502
R4 plus.n3 plus.t4 397.651
R5 plus.n7 plus.t15 397.651
R6 plus.n9 plus.t11 397.651
R7 plus.n1 plus.t10 397.651
R8 plus.n14 plus.t6 397.651
R9 plus.n16 plus.t3 397.651
R10 plus.n22 plus.t2 397.651
R11 plus.n26 plus.t9 397.651
R12 plus.n28 plus.t1 397.651
R13 plus.n20 plus.t5 397.651
R14 plus.n33 plus.t12 397.651
R15 plus.n35 plus.t0 397.651
R16 plus.n5 plus.n4 161.489
R17 plus.n24 plus.n23 161.489
R18 plus.n6 plus.n5 161.3
R19 plus.n8 plus.n2 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n0 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n25 plus.n24 161.3
R25 plus.n27 plus.n21 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n19 161.3
R29 plus.n37 plus.n36 161.3
R30 plus.n6 plus.n3 47.4702
R31 plus.n16 plus.n15 47.4702
R32 plus.n35 plus.n34 47.4702
R33 plus.n25 plus.n22 47.4702
R34 plus.n8 plus.n7 43.0884
R35 plus.n14 plus.n13 43.0884
R36 plus.n33 plus.n32 43.0884
R37 plus.n27 plus.n26 43.0884
R38 plus.n10 plus.n9 38.7066
R39 plus.n10 plus.n1 38.7066
R40 plus.n29 plus.n20 38.7066
R41 plus.n29 plus.n28 38.7066
R42 plus.n9 plus.n8 34.3247
R43 plus.n13 plus.n1 34.3247
R44 plus.n32 plus.n20 34.3247
R45 plus.n28 plus.n27 34.3247
R46 plus.n7 plus.n6 29.9429
R47 plus.n15 plus.n14 29.9429
R48 plus.n34 plus.n33 29.9429
R49 plus.n26 plus.n25 29.9429
R50 plus.n4 plus.n3 25.5611
R51 plus.n17 plus.n16 25.5611
R52 plus.n36 plus.n35 25.5611
R53 plus.n23 plus.n22 25.5611
R54 plus plus.n37 25.5066
R55 plus plus.n18 8.32247
R56 plus.n5 plus.n2 0.189894
R57 plus.n11 plus.n2 0.189894
R58 plus.n12 plus.n11 0.189894
R59 plus.n12 plus.n0 0.189894
R60 plus.n18 plus.n0 0.189894
R61 plus.n37 plus.n19 0.189894
R62 plus.n31 plus.n19 0.189894
R63 plus.n31 plus.n30 0.189894
R64 plus.n30 plus.n21 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n82 source.n80 289.615
R67 source.n68 source.n66 289.615
R68 source.n60 source.n58 289.615
R69 source.n46 source.n44 289.615
R70 source.n2 source.n0 289.615
R71 source.n16 source.n14 289.615
R72 source.n24 source.n22 289.615
R73 source.n38 source.n36 289.615
R74 source.n83 source.n82 185
R75 source.n69 source.n68 185
R76 source.n61 source.n60 185
R77 source.n47 source.n46 185
R78 source.n3 source.n2 185
R79 source.n17 source.n16 185
R80 source.n25 source.n24 185
R81 source.n39 source.n38 185
R82 source.t14 source.n81 167.117
R83 source.t13 source.n67 167.117
R84 source.t23 source.n59 167.117
R85 source.t22 source.n45 167.117
R86 source.t27 source.n1 167.117
R87 source.t24 source.n15 167.117
R88 source.t0 source.n23 167.117
R89 source.t3 source.n37 167.117
R90 source.n9 source.n8 84.1169
R91 source.n11 source.n10 84.1169
R92 source.n13 source.n12 84.1169
R93 source.n31 source.n30 84.1169
R94 source.n33 source.n32 84.1169
R95 source.n35 source.n34 84.1169
R96 source.n79 source.n78 84.1168
R97 source.n77 source.n76 84.1168
R98 source.n75 source.n74 84.1168
R99 source.n57 source.n56 84.1168
R100 source.n55 source.n54 84.1168
R101 source.n53 source.n52 84.1168
R102 source.n82 source.t14 52.3082
R103 source.n68 source.t13 52.3082
R104 source.n60 source.t23 52.3082
R105 source.n46 source.t22 52.3082
R106 source.n2 source.t27 52.3082
R107 source.n16 source.t24 52.3082
R108 source.n24 source.t0 52.3082
R109 source.n38 source.t3 52.3082
R110 source.n87 source.n86 31.4096
R111 source.n73 source.n72 31.4096
R112 source.n65 source.n64 31.4096
R113 source.n51 source.n50 31.4096
R114 source.n7 source.n6 31.4096
R115 source.n21 source.n20 31.4096
R116 source.n29 source.n28 31.4096
R117 source.n43 source.n42 31.4096
R118 source.n51 source.n43 14.1689
R119 source.n78 source.t8 9.9005
R120 source.n78 source.t1 9.9005
R121 source.n76 source.t7 9.9005
R122 source.n76 source.t9 9.9005
R123 source.n74 source.t5 9.9005
R124 source.n74 source.t11 9.9005
R125 source.n56 source.t31 9.9005
R126 source.n56 source.t26 9.9005
R127 source.n54 source.t29 9.9005
R128 source.n54 source.t17 9.9005
R129 source.n52 source.t18 9.9005
R130 source.n52 source.t30 9.9005
R131 source.n8 source.t25 9.9005
R132 source.n8 source.t19 9.9005
R133 source.n10 source.t28 9.9005
R134 source.n10 source.t21 9.9005
R135 source.n12 source.t20 9.9005
R136 source.n12 source.t16 9.9005
R137 source.n30 source.t6 9.9005
R138 source.n30 source.t4 9.9005
R139 source.n32 source.t12 9.9005
R140 source.n32 source.t2 9.9005
R141 source.n34 source.t15 9.9005
R142 source.n34 source.t10 9.9005
R143 source.n83 source.n81 9.71174
R144 source.n69 source.n67 9.71174
R145 source.n61 source.n59 9.71174
R146 source.n47 source.n45 9.71174
R147 source.n3 source.n1 9.71174
R148 source.n17 source.n15 9.71174
R149 source.n25 source.n23 9.71174
R150 source.n39 source.n37 9.71174
R151 source.n86 source.n85 9.45567
R152 source.n72 source.n71 9.45567
R153 source.n64 source.n63 9.45567
R154 source.n50 source.n49 9.45567
R155 source.n6 source.n5 9.45567
R156 source.n20 source.n19 9.45567
R157 source.n28 source.n27 9.45567
R158 source.n42 source.n41 9.45567
R159 source.n85 source.n84 9.3005
R160 source.n71 source.n70 9.3005
R161 source.n63 source.n62 9.3005
R162 source.n49 source.n48 9.3005
R163 source.n5 source.n4 9.3005
R164 source.n19 source.n18 9.3005
R165 source.n27 source.n26 9.3005
R166 source.n41 source.n40 9.3005
R167 source.n88 source.n7 8.67749
R168 source.n86 source.n80 8.14595
R169 source.n72 source.n66 8.14595
R170 source.n64 source.n58 8.14595
R171 source.n50 source.n44 8.14595
R172 source.n6 source.n0 8.14595
R173 source.n20 source.n14 8.14595
R174 source.n28 source.n22 8.14595
R175 source.n42 source.n36 8.14595
R176 source.n84 source.n83 7.3702
R177 source.n70 source.n69 7.3702
R178 source.n62 source.n61 7.3702
R179 source.n48 source.n47 7.3702
R180 source.n4 source.n3 7.3702
R181 source.n18 source.n17 7.3702
R182 source.n26 source.n25 7.3702
R183 source.n40 source.n39 7.3702
R184 source.n84 source.n80 5.81868
R185 source.n70 source.n66 5.81868
R186 source.n62 source.n58 5.81868
R187 source.n48 source.n44 5.81868
R188 source.n4 source.n0 5.81868
R189 source.n18 source.n14 5.81868
R190 source.n26 source.n22 5.81868
R191 source.n40 source.n36 5.81868
R192 source.n88 source.n87 5.49188
R193 source.n85 source.n81 3.44771
R194 source.n71 source.n67 3.44771
R195 source.n63 source.n59 3.44771
R196 source.n49 source.n45 3.44771
R197 source.n5 source.n1 3.44771
R198 source.n19 source.n15 3.44771
R199 source.n27 source.n23 3.44771
R200 source.n41 source.n37 3.44771
R201 source.n29 source.n21 0.470328
R202 source.n73 source.n65 0.470328
R203 source.n43 source.n35 0.457397
R204 source.n35 source.n33 0.457397
R205 source.n33 source.n31 0.457397
R206 source.n31 source.n29 0.457397
R207 source.n21 source.n13 0.457397
R208 source.n13 source.n11 0.457397
R209 source.n11 source.n9 0.457397
R210 source.n9 source.n7 0.457397
R211 source.n53 source.n51 0.457397
R212 source.n55 source.n53 0.457397
R213 source.n57 source.n55 0.457397
R214 source.n65 source.n57 0.457397
R215 source.n75 source.n73 0.457397
R216 source.n77 source.n75 0.457397
R217 source.n79 source.n77 0.457397
R218 source.n87 source.n79 0.457397
R219 source source.n88 0.188
R220 drain_left.n9 drain_left.n7 101.252
R221 drain_left.n5 drain_left.n3 101.252
R222 drain_left.n2 drain_left.n0 101.252
R223 drain_left.n13 drain_left.n12 100.796
R224 drain_left.n11 drain_left.n10 100.796
R225 drain_left.n9 drain_left.n8 100.796
R226 drain_left.n5 drain_left.n4 100.796
R227 drain_left.n2 drain_left.n1 100.796
R228 drain_left drain_left.n6 22.7611
R229 drain_left.n3 drain_left.t13 9.9005
R230 drain_left.n3 drain_left.t2 9.9005
R231 drain_left.n4 drain_left.t14 9.9005
R232 drain_left.n4 drain_left.t6 9.9005
R233 drain_left.n1 drain_left.t3 9.9005
R234 drain_left.n1 drain_left.t10 9.9005
R235 drain_left.n0 drain_left.t7 9.9005
R236 drain_left.n0 drain_left.t15 9.9005
R237 drain_left.n12 drain_left.t12 9.9005
R238 drain_left.n12 drain_left.t1 9.9005
R239 drain_left.n10 drain_left.t5 9.9005
R240 drain_left.n10 drain_left.t9 9.9005
R241 drain_left.n8 drain_left.t0 9.9005
R242 drain_left.n8 drain_left.t4 9.9005
R243 drain_left.n7 drain_left.t8 9.9005
R244 drain_left.n7 drain_left.t11 9.9005
R245 drain_left drain_left.n13 6.11011
R246 drain_left.n11 drain_left.n9 0.457397
R247 drain_left.n13 drain_left.n11 0.457397
R248 drain_left.n6 drain_left.n5 0.173602
R249 drain_left.n6 drain_left.n2 0.173602
R250 minus.n17 minus.t14 449.502
R251 minus.n4 minus.t9 449.502
R252 minus.n36 minus.t4 449.502
R253 minus.n23 minus.t15 449.502
R254 minus.n16 minus.t3 397.651
R255 minus.n14 minus.t5 397.651
R256 minus.n1 minus.t10 397.651
R257 minus.n9 minus.t13 397.651
R258 minus.n7 minus.t2 397.651
R259 minus.n3 minus.t6 397.651
R260 minus.n35 minus.t11 397.651
R261 minus.n33 minus.t7 397.651
R262 minus.n20 minus.t0 397.651
R263 minus.n28 minus.t12 397.651
R264 minus.n26 minus.t8 397.651
R265 minus.n22 minus.t1 397.651
R266 minus.n5 minus.n4 161.489
R267 minus.n24 minus.n23 161.489
R268 minus.n18 minus.n17 161.3
R269 minus.n15 minus.n0 161.3
R270 minus.n13 minus.n12 161.3
R271 minus.n11 minus.n10 161.3
R272 minus.n8 minus.n2 161.3
R273 minus.n6 minus.n5 161.3
R274 minus.n37 minus.n36 161.3
R275 minus.n34 minus.n19 161.3
R276 minus.n32 minus.n31 161.3
R277 minus.n30 minus.n29 161.3
R278 minus.n27 minus.n21 161.3
R279 minus.n25 minus.n24 161.3
R280 minus.n16 minus.n15 47.4702
R281 minus.n6 minus.n3 47.4702
R282 minus.n25 minus.n22 47.4702
R283 minus.n35 minus.n34 47.4702
R284 minus.n14 minus.n13 43.0884
R285 minus.n8 minus.n7 43.0884
R286 minus.n27 minus.n26 43.0884
R287 minus.n33 minus.n32 43.0884
R288 minus.n10 minus.n1 38.7066
R289 minus.n10 minus.n9 38.7066
R290 minus.n29 minus.n28 38.7066
R291 minus.n29 minus.n20 38.7066
R292 minus.n13 minus.n1 34.3247
R293 minus.n9 minus.n8 34.3247
R294 minus.n28 minus.n27 34.3247
R295 minus.n32 minus.n20 34.3247
R296 minus.n15 minus.n14 29.9429
R297 minus.n7 minus.n6 29.9429
R298 minus.n26 minus.n25 29.9429
R299 minus.n34 minus.n33 29.9429
R300 minus.n38 minus.n18 27.8376
R301 minus.n17 minus.n16 25.5611
R302 minus.n4 minus.n3 25.5611
R303 minus.n23 minus.n22 25.5611
R304 minus.n36 minus.n35 25.5611
R305 minus.n38 minus.n37 6.46641
R306 minus.n18 minus.n0 0.189894
R307 minus.n12 minus.n0 0.189894
R308 minus.n12 minus.n11 0.189894
R309 minus.n11 minus.n2 0.189894
R310 minus.n5 minus.n2 0.189894
R311 minus.n24 minus.n21 0.189894
R312 minus.n30 minus.n21 0.189894
R313 minus.n31 minus.n30 0.189894
R314 minus.n31 minus.n19 0.189894
R315 minus.n37 minus.n19 0.189894
R316 minus minus.n38 0.188
R317 drain_right.n9 drain_right.n7 101.252
R318 drain_right.n5 drain_right.n3 101.252
R319 drain_right.n2 drain_right.n0 101.252
R320 drain_right.n9 drain_right.n8 100.796
R321 drain_right.n11 drain_right.n10 100.796
R322 drain_right.n13 drain_right.n12 100.796
R323 drain_right.n5 drain_right.n4 100.796
R324 drain_right.n2 drain_right.n1 100.796
R325 drain_right drain_right.n6 22.2079
R326 drain_right.n3 drain_right.t4 9.9005
R327 drain_right.n3 drain_right.t11 9.9005
R328 drain_right.n4 drain_right.t15 9.9005
R329 drain_right.n4 drain_right.t8 9.9005
R330 drain_right.n1 drain_right.t7 9.9005
R331 drain_right.n1 drain_right.t3 9.9005
R332 drain_right.n0 drain_right.t0 9.9005
R333 drain_right.n0 drain_right.t14 9.9005
R334 drain_right.n7 drain_right.t9 9.9005
R335 drain_right.n7 drain_right.t6 9.9005
R336 drain_right.n8 drain_right.t2 9.9005
R337 drain_right.n8 drain_right.t13 9.9005
R338 drain_right.n10 drain_right.t10 9.9005
R339 drain_right.n10 drain_right.t5 9.9005
R340 drain_right.n12 drain_right.t1 9.9005
R341 drain_right.n12 drain_right.t12 9.9005
R342 drain_right drain_right.n13 6.11011
R343 drain_right.n13 drain_right.n11 0.457397
R344 drain_right.n11 drain_right.n9 0.457397
R345 drain_right.n6 drain_right.n5 0.173602
R346 drain_right.n6 drain_right.n2 0.173602
C0 drain_right drain_left 0.846053f
C1 source drain_left 8.37424f
C2 drain_right plus 0.321281f
C3 source plus 1.28815f
C4 drain_left minus 0.176775f
C5 plus minus 3.39327f
C6 drain_right source 8.37391f
C7 drain_right minus 1.15454f
C8 source minus 1.27418f
C9 drain_left plus 1.31552f
C10 drain_right a_n1670_n1288# 3.93185f
C11 drain_left a_n1670_n1288# 4.16878f
C12 source a_n1670_n1288# 3.039674f
C13 minus a_n1670_n1288# 5.671903f
C14 plus a_n1670_n1288# 6.346002f
C15 drain_right.t0 a_n1670_n1288# 0.048493f
C16 drain_right.t14 a_n1670_n1288# 0.048493f
C17 drain_right.n0 a_n1670_n1288# 0.306174f
C18 drain_right.t7 a_n1670_n1288# 0.048493f
C19 drain_right.t3 a_n1670_n1288# 0.048493f
C20 drain_right.n1 a_n1670_n1288# 0.304651f
C21 drain_right.n2 a_n1670_n1288# 0.637268f
C22 drain_right.t4 a_n1670_n1288# 0.048493f
C23 drain_right.t11 a_n1670_n1288# 0.048493f
C24 drain_right.n3 a_n1670_n1288# 0.306174f
C25 drain_right.t15 a_n1670_n1288# 0.048493f
C26 drain_right.t8 a_n1670_n1288# 0.048493f
C27 drain_right.n4 a_n1670_n1288# 0.304651f
C28 drain_right.n5 a_n1670_n1288# 0.637268f
C29 drain_right.n6 a_n1670_n1288# 0.754067f
C30 drain_right.t9 a_n1670_n1288# 0.048493f
C31 drain_right.t6 a_n1670_n1288# 0.048493f
C32 drain_right.n7 a_n1670_n1288# 0.306175f
C33 drain_right.t2 a_n1670_n1288# 0.048493f
C34 drain_right.t13 a_n1670_n1288# 0.048493f
C35 drain_right.n8 a_n1670_n1288# 0.304652f
C36 drain_right.n9 a_n1670_n1288# 0.661214f
C37 drain_right.t10 a_n1670_n1288# 0.048493f
C38 drain_right.t5 a_n1670_n1288# 0.048493f
C39 drain_right.n10 a_n1670_n1288# 0.304652f
C40 drain_right.n11 a_n1670_n1288# 0.325189f
C41 drain_right.t1 a_n1670_n1288# 0.048493f
C42 drain_right.t12 a_n1670_n1288# 0.048493f
C43 drain_right.n12 a_n1670_n1288# 0.304652f
C44 drain_right.n13 a_n1670_n1288# 0.576301f
C45 minus.n0 a_n1670_n1288# 0.031099f
C46 minus.t14 a_n1670_n1288# 0.040044f
C47 minus.t3 a_n1670_n1288# 0.036605f
C48 minus.t5 a_n1670_n1288# 0.036605f
C49 minus.t10 a_n1670_n1288# 0.036605f
C50 minus.n1 a_n1670_n1288# 0.028761f
C51 minus.n2 a_n1670_n1288# 0.031099f
C52 minus.t13 a_n1670_n1288# 0.036605f
C53 minus.t2 a_n1670_n1288# 0.036605f
C54 minus.t6 a_n1670_n1288# 0.036605f
C55 minus.n3 a_n1670_n1288# 0.028761f
C56 minus.t9 a_n1670_n1288# 0.040044f
C57 minus.n4 a_n1670_n1288# 0.037314f
C58 minus.n5 a_n1670_n1288# 0.070014f
C59 minus.n6 a_n1670_n1288# 0.010892f
C60 minus.n7 a_n1670_n1288# 0.028761f
C61 minus.n8 a_n1670_n1288# 0.010892f
C62 minus.n9 a_n1670_n1288# 0.028761f
C63 minus.n10 a_n1670_n1288# 0.010892f
C64 minus.n11 a_n1670_n1288# 0.031099f
C65 minus.n12 a_n1670_n1288# 0.031099f
C66 minus.n13 a_n1670_n1288# 0.010892f
C67 minus.n14 a_n1670_n1288# 0.028761f
C68 minus.n15 a_n1670_n1288# 0.010892f
C69 minus.n16 a_n1670_n1288# 0.028761f
C70 minus.n17 a_n1670_n1288# 0.037268f
C71 minus.n18 a_n1670_n1288# 0.70917f
C72 minus.n19 a_n1670_n1288# 0.031099f
C73 minus.t11 a_n1670_n1288# 0.036605f
C74 minus.t7 a_n1670_n1288# 0.036605f
C75 minus.t0 a_n1670_n1288# 0.036605f
C76 minus.n20 a_n1670_n1288# 0.028761f
C77 minus.n21 a_n1670_n1288# 0.031099f
C78 minus.t12 a_n1670_n1288# 0.036605f
C79 minus.t8 a_n1670_n1288# 0.036605f
C80 minus.t1 a_n1670_n1288# 0.036605f
C81 minus.n22 a_n1670_n1288# 0.028761f
C82 minus.t15 a_n1670_n1288# 0.040044f
C83 minus.n23 a_n1670_n1288# 0.037314f
C84 minus.n24 a_n1670_n1288# 0.070014f
C85 minus.n25 a_n1670_n1288# 0.010892f
C86 minus.n26 a_n1670_n1288# 0.028761f
C87 minus.n27 a_n1670_n1288# 0.010892f
C88 minus.n28 a_n1670_n1288# 0.028761f
C89 minus.n29 a_n1670_n1288# 0.010892f
C90 minus.n30 a_n1670_n1288# 0.031099f
C91 minus.n31 a_n1670_n1288# 0.031099f
C92 minus.n32 a_n1670_n1288# 0.010892f
C93 minus.n33 a_n1670_n1288# 0.028761f
C94 minus.n34 a_n1670_n1288# 0.010892f
C95 minus.n35 a_n1670_n1288# 0.028761f
C96 minus.t4 a_n1670_n1288# 0.040044f
C97 minus.n36 a_n1670_n1288# 0.037268f
C98 minus.n37 a_n1670_n1288# 0.200854f
C99 minus.n38 a_n1670_n1288# 0.878078f
C100 drain_left.t7 a_n1670_n1288# 0.04781f
C101 drain_left.t15 a_n1670_n1288# 0.04781f
C102 drain_left.n0 a_n1670_n1288# 0.301861f
C103 drain_left.t3 a_n1670_n1288# 0.04781f
C104 drain_left.t10 a_n1670_n1288# 0.04781f
C105 drain_left.n1 a_n1670_n1288# 0.300359f
C106 drain_left.n2 a_n1670_n1288# 0.62829f
C107 drain_left.t13 a_n1670_n1288# 0.04781f
C108 drain_left.t2 a_n1670_n1288# 0.04781f
C109 drain_left.n3 a_n1670_n1288# 0.301861f
C110 drain_left.t14 a_n1670_n1288# 0.04781f
C111 drain_left.t6 a_n1670_n1288# 0.04781f
C112 drain_left.n4 a_n1670_n1288# 0.300359f
C113 drain_left.n5 a_n1670_n1288# 0.62829f
C114 drain_left.n6 a_n1670_n1288# 0.802806f
C115 drain_left.t8 a_n1670_n1288# 0.04781f
C116 drain_left.t11 a_n1670_n1288# 0.04781f
C117 drain_left.n7 a_n1670_n1288# 0.301862f
C118 drain_left.t0 a_n1670_n1288# 0.04781f
C119 drain_left.t4 a_n1670_n1288# 0.04781f
C120 drain_left.n8 a_n1670_n1288# 0.30036f
C121 drain_left.n9 a_n1670_n1288# 0.651899f
C122 drain_left.t5 a_n1670_n1288# 0.04781f
C123 drain_left.t9 a_n1670_n1288# 0.04781f
C124 drain_left.n10 a_n1670_n1288# 0.30036f
C125 drain_left.n11 a_n1670_n1288# 0.320608f
C126 drain_left.t12 a_n1670_n1288# 0.04781f
C127 drain_left.t1 a_n1670_n1288# 0.04781f
C128 drain_left.n12 a_n1670_n1288# 0.30036f
C129 drain_left.n13 a_n1670_n1288# 0.568182f
C130 source.n0 a_n1670_n1288# 0.045516f
C131 source.n1 a_n1670_n1288# 0.100709f
C132 source.t27 a_n1670_n1288# 0.075577f
C133 source.n2 a_n1670_n1288# 0.078819f
C134 source.n3 a_n1670_n1288# 0.025408f
C135 source.n4 a_n1670_n1288# 0.016757f
C136 source.n5 a_n1670_n1288# 0.221987f
C137 source.n6 a_n1670_n1288# 0.049896f
C138 source.n7 a_n1670_n1288# 0.455429f
C139 source.t25 a_n1670_n1288# 0.049286f
C140 source.t19 a_n1670_n1288# 0.049286f
C141 source.n8 a_n1670_n1288# 0.263481f
C142 source.n9 a_n1670_n1288# 0.334266f
C143 source.t28 a_n1670_n1288# 0.049286f
C144 source.t21 a_n1670_n1288# 0.049286f
C145 source.n10 a_n1670_n1288# 0.263481f
C146 source.n11 a_n1670_n1288# 0.334266f
C147 source.t20 a_n1670_n1288# 0.049286f
C148 source.t16 a_n1670_n1288# 0.049286f
C149 source.n12 a_n1670_n1288# 0.263481f
C150 source.n13 a_n1670_n1288# 0.334266f
C151 source.n14 a_n1670_n1288# 0.045516f
C152 source.n15 a_n1670_n1288# 0.100709f
C153 source.t24 a_n1670_n1288# 0.075577f
C154 source.n16 a_n1670_n1288# 0.078819f
C155 source.n17 a_n1670_n1288# 0.025408f
C156 source.n18 a_n1670_n1288# 0.016757f
C157 source.n19 a_n1670_n1288# 0.221987f
C158 source.n20 a_n1670_n1288# 0.049896f
C159 source.n21 a_n1670_n1288# 0.118793f
C160 source.n22 a_n1670_n1288# 0.045516f
C161 source.n23 a_n1670_n1288# 0.100709f
C162 source.t0 a_n1670_n1288# 0.075577f
C163 source.n24 a_n1670_n1288# 0.078819f
C164 source.n25 a_n1670_n1288# 0.025408f
C165 source.n26 a_n1670_n1288# 0.016757f
C166 source.n27 a_n1670_n1288# 0.221987f
C167 source.n28 a_n1670_n1288# 0.049896f
C168 source.n29 a_n1670_n1288# 0.118793f
C169 source.t6 a_n1670_n1288# 0.049286f
C170 source.t4 a_n1670_n1288# 0.049286f
C171 source.n30 a_n1670_n1288# 0.263481f
C172 source.n31 a_n1670_n1288# 0.334266f
C173 source.t12 a_n1670_n1288# 0.049286f
C174 source.t2 a_n1670_n1288# 0.049286f
C175 source.n32 a_n1670_n1288# 0.263481f
C176 source.n33 a_n1670_n1288# 0.334266f
C177 source.t15 a_n1670_n1288# 0.049286f
C178 source.t10 a_n1670_n1288# 0.049286f
C179 source.n34 a_n1670_n1288# 0.263481f
C180 source.n35 a_n1670_n1288# 0.334266f
C181 source.n36 a_n1670_n1288# 0.045516f
C182 source.n37 a_n1670_n1288# 0.100709f
C183 source.t3 a_n1670_n1288# 0.075577f
C184 source.n38 a_n1670_n1288# 0.078819f
C185 source.n39 a_n1670_n1288# 0.025408f
C186 source.n40 a_n1670_n1288# 0.016757f
C187 source.n41 a_n1670_n1288# 0.221987f
C188 source.n42 a_n1670_n1288# 0.049896f
C189 source.n43 a_n1670_n1288# 0.744244f
C190 source.n44 a_n1670_n1288# 0.045516f
C191 source.n45 a_n1670_n1288# 0.100709f
C192 source.t22 a_n1670_n1288# 0.075577f
C193 source.n46 a_n1670_n1288# 0.078819f
C194 source.n47 a_n1670_n1288# 0.025408f
C195 source.n48 a_n1670_n1288# 0.016757f
C196 source.n49 a_n1670_n1288# 0.221987f
C197 source.n50 a_n1670_n1288# 0.049896f
C198 source.n51 a_n1670_n1288# 0.744244f
C199 source.t18 a_n1670_n1288# 0.049286f
C200 source.t30 a_n1670_n1288# 0.049286f
C201 source.n52 a_n1670_n1288# 0.263479f
C202 source.n53 a_n1670_n1288# 0.334268f
C203 source.t29 a_n1670_n1288# 0.049286f
C204 source.t17 a_n1670_n1288# 0.049286f
C205 source.n54 a_n1670_n1288# 0.263479f
C206 source.n55 a_n1670_n1288# 0.334268f
C207 source.t31 a_n1670_n1288# 0.049286f
C208 source.t26 a_n1670_n1288# 0.049286f
C209 source.n56 a_n1670_n1288# 0.263479f
C210 source.n57 a_n1670_n1288# 0.334268f
C211 source.n58 a_n1670_n1288# 0.045516f
C212 source.n59 a_n1670_n1288# 0.100709f
C213 source.t23 a_n1670_n1288# 0.075577f
C214 source.n60 a_n1670_n1288# 0.078819f
C215 source.n61 a_n1670_n1288# 0.025408f
C216 source.n62 a_n1670_n1288# 0.016757f
C217 source.n63 a_n1670_n1288# 0.221987f
C218 source.n64 a_n1670_n1288# 0.049896f
C219 source.n65 a_n1670_n1288# 0.118793f
C220 source.n66 a_n1670_n1288# 0.045516f
C221 source.n67 a_n1670_n1288# 0.100709f
C222 source.t13 a_n1670_n1288# 0.075577f
C223 source.n68 a_n1670_n1288# 0.078819f
C224 source.n69 a_n1670_n1288# 0.025408f
C225 source.n70 a_n1670_n1288# 0.016757f
C226 source.n71 a_n1670_n1288# 0.221987f
C227 source.n72 a_n1670_n1288# 0.049896f
C228 source.n73 a_n1670_n1288# 0.118793f
C229 source.t5 a_n1670_n1288# 0.049286f
C230 source.t11 a_n1670_n1288# 0.049286f
C231 source.n74 a_n1670_n1288# 0.263479f
C232 source.n75 a_n1670_n1288# 0.334268f
C233 source.t7 a_n1670_n1288# 0.049286f
C234 source.t9 a_n1670_n1288# 0.049286f
C235 source.n76 a_n1670_n1288# 0.263479f
C236 source.n77 a_n1670_n1288# 0.334268f
C237 source.t8 a_n1670_n1288# 0.049286f
C238 source.t1 a_n1670_n1288# 0.049286f
C239 source.n78 a_n1670_n1288# 0.263479f
C240 source.n79 a_n1670_n1288# 0.334268f
C241 source.n80 a_n1670_n1288# 0.045516f
C242 source.n81 a_n1670_n1288# 0.100709f
C243 source.t14 a_n1670_n1288# 0.075577f
C244 source.n82 a_n1670_n1288# 0.078819f
C245 source.n83 a_n1670_n1288# 0.025408f
C246 source.n84 a_n1670_n1288# 0.016757f
C247 source.n85 a_n1670_n1288# 0.221987f
C248 source.n86 a_n1670_n1288# 0.049896f
C249 source.n87 a_n1670_n1288# 0.287885f
C250 source.n88 a_n1670_n1288# 0.767356f
C251 plus.n0 a_n1670_n1288# 0.031685f
C252 plus.t3 a_n1670_n1288# 0.037295f
C253 plus.t6 a_n1670_n1288# 0.037295f
C254 plus.t10 a_n1670_n1288# 0.037295f
C255 plus.n1 a_n1670_n1288# 0.029303f
C256 plus.n2 a_n1670_n1288# 0.031685f
C257 plus.t11 a_n1670_n1288# 0.037295f
C258 plus.t15 a_n1670_n1288# 0.037295f
C259 plus.t4 a_n1670_n1288# 0.037295f
C260 plus.n3 a_n1670_n1288# 0.029303f
C261 plus.t7 a_n1670_n1288# 0.040799f
C262 plus.n4 a_n1670_n1288# 0.038017f
C263 plus.n5 a_n1670_n1288# 0.071334f
C264 plus.n6 a_n1670_n1288# 0.011097f
C265 plus.n7 a_n1670_n1288# 0.029303f
C266 plus.n8 a_n1670_n1288# 0.011097f
C267 plus.n9 a_n1670_n1288# 0.029303f
C268 plus.n10 a_n1670_n1288# 0.011097f
C269 plus.n11 a_n1670_n1288# 0.031685f
C270 plus.n12 a_n1670_n1288# 0.031685f
C271 plus.n13 a_n1670_n1288# 0.011097f
C272 plus.n14 a_n1670_n1288# 0.029303f
C273 plus.n15 a_n1670_n1288# 0.011097f
C274 plus.n16 a_n1670_n1288# 0.029303f
C275 plus.t14 a_n1670_n1288# 0.040799f
C276 plus.n17 a_n1670_n1288# 0.037971f
C277 plus.n18 a_n1670_n1288# 0.22387f
C278 plus.n19 a_n1670_n1288# 0.031685f
C279 plus.t8 a_n1670_n1288# 0.040799f
C280 plus.t0 a_n1670_n1288# 0.037295f
C281 plus.t12 a_n1670_n1288# 0.037295f
C282 plus.t5 a_n1670_n1288# 0.037295f
C283 plus.n20 a_n1670_n1288# 0.029303f
C284 plus.n21 a_n1670_n1288# 0.031685f
C285 plus.t1 a_n1670_n1288# 0.037295f
C286 plus.t9 a_n1670_n1288# 0.037295f
C287 plus.t2 a_n1670_n1288# 0.037295f
C288 plus.n22 a_n1670_n1288# 0.029303f
C289 plus.t13 a_n1670_n1288# 0.040799f
C290 plus.n23 a_n1670_n1288# 0.038017f
C291 plus.n24 a_n1670_n1288# 0.071334f
C292 plus.n25 a_n1670_n1288# 0.011097f
C293 plus.n26 a_n1670_n1288# 0.029303f
C294 plus.n27 a_n1670_n1288# 0.011097f
C295 plus.n28 a_n1670_n1288# 0.029303f
C296 plus.n29 a_n1670_n1288# 0.011097f
C297 plus.n30 a_n1670_n1288# 0.031685f
C298 plus.n31 a_n1670_n1288# 0.031685f
C299 plus.n32 a_n1670_n1288# 0.011097f
C300 plus.n33 a_n1670_n1288# 0.029303f
C301 plus.n34 a_n1670_n1288# 0.011097f
C302 plus.n35 a_n1670_n1288# 0.029303f
C303 plus.n36 a_n1670_n1288# 0.037971f
C304 plus.n37 a_n1670_n1288# 0.69091f
.ends

