* NGSPICE file created from diffpair319.ext - technology: sky130A

.subckt diffpair319 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t16 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X1 source.t8 plus.t0 drain_left.t23 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 drain_left.t22 plus.t1 source.t7 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X3 drain_left.t21 plus.t2 source.t17 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X4 drain_right.t5 minus.t1 source.t46 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X5 drain_left.t20 plus.t3 source.t19 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X6 drain_left.t19 plus.t4 source.t3 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X7 drain_left.t18 plus.t5 source.t0 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X8 source.t45 minus.t2 drain_right.t1 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X9 source.t44 minus.t3 drain_right.t0 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X10 source.t43 minus.t4 drain_right.t2 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X11 source.t42 minus.t5 drain_right.t3 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X12 drain_left.t17 plus.t6 source.t5 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X13 source.t11 plus.t7 drain_left.t16 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X14 source.t23 plus.t8 drain_left.t15 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X15 drain_right.t14 minus.t6 source.t41 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X16 drain_left.t14 plus.t9 source.t12 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X17 drain_right.t22 minus.t7 source.t40 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X18 source.t39 minus.t8 drain_right.t20 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X19 drain_left.t13 plus.t10 source.t10 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X20 source.t38 minus.t9 drain_right.t19 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X21 source.t37 minus.t10 drain_right.t12 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X22 drain_right.t13 minus.t11 source.t36 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X23 drain_right.t23 minus.t12 source.t35 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X24 source.t34 minus.t13 drain_right.t6 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X25 source.t18 plus.t11 drain_left.t12 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X26 drain_right.t8 minus.t14 source.t33 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X27 source.t1 plus.t12 drain_left.t11 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X28 source.t20 plus.t13 drain_left.t10 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X29 source.t32 minus.t15 drain_right.t10 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X30 drain_right.t17 minus.t16 source.t31 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X31 drain_left.t9 plus.t14 source.t21 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X32 source.t30 minus.t17 drain_right.t7 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X33 drain_right.t9 minus.t18 source.t29 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X34 drain_right.t4 minus.t19 source.t28 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X35 drain_right.t15 minus.t20 source.t27 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X36 a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X37 source.t13 plus.t15 drain_left.t8 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X38 a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X39 source.t4 plus.t16 drain_left.t7 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X40 drain_left.t6 plus.t17 source.t6 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X41 drain_left.t5 plus.t18 source.t2 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X42 source.t26 minus.t21 drain_right.t11 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X43 source.t14 plus.t19 drain_left.t4 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X44 drain_right.t21 minus.t22 source.t25 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X45 source.t16 plus.t20 drain_left.t3 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X46 drain_left.t2 plus.t21 source.t9 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X47 a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X48 source.t15 plus.t22 drain_left.t1 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X49 drain_right.t18 minus.t23 source.t24 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X50 source.t22 plus.t23 drain_left.t0 a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X51 a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# a_n3654_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
R0 minus.n8 minus.t14 251.291
R1 minus.n44 minus.t13 251.291
R2 minus.n9 minus.t9 229.855
R3 minus.n10 minus.t6 229.855
R4 minus.n14 minus.t17 229.855
R5 minus.n16 minus.t19 229.855
R6 minus.n20 minus.t15 229.855
R7 minus.n21 minus.t11 229.855
R8 minus.n3 minus.t21 229.855
R9 minus.n27 minus.t18 229.855
R10 minus.n1 minus.t3 229.855
R11 minus.n32 minus.t12 229.855
R12 minus.n34 minus.t10 229.855
R13 minus.n45 minus.t1 229.855
R14 minus.n46 minus.t5 229.855
R15 minus.n50 minus.t23 229.855
R16 minus.n52 minus.t8 229.855
R17 minus.n56 minus.t22 229.855
R18 minus.n57 minus.t2 229.855
R19 minus.n39 minus.t16 229.855
R20 minus.n63 minus.t4 229.855
R21 minus.n37 minus.t20 229.855
R22 minus.n68 minus.t0 229.855
R23 minus.n70 minus.t7 229.855
R24 minus.n35 minus.n34 161.3
R25 minus.n33 minus.n0 161.3
R26 minus.n29 minus.n28 161.3
R27 minus.n27 minus.n2 161.3
R28 minus.n26 minus.n25 161.3
R29 minus.n24 minus.n3 161.3
R30 minus.n23 minus.n22 161.3
R31 minus.n18 minus.n5 161.3
R32 minus.n17 minus.n16 161.3
R33 minus.n15 minus.n6 161.3
R34 minus.n14 minus.n13 161.3
R35 minus.n12 minus.n7 161.3
R36 minus.n71 minus.n70 161.3
R37 minus.n69 minus.n36 161.3
R38 minus.n65 minus.n64 161.3
R39 minus.n63 minus.n38 161.3
R40 minus.n62 minus.n61 161.3
R41 minus.n60 minus.n39 161.3
R42 minus.n59 minus.n58 161.3
R43 minus.n54 minus.n41 161.3
R44 minus.n53 minus.n52 161.3
R45 minus.n51 minus.n42 161.3
R46 minus.n50 minus.n49 161.3
R47 minus.n48 minus.n43 161.3
R48 minus.n32 minus.n31 80.6037
R49 minus.n30 minus.n1 80.6037
R50 minus.n21 minus.n4 80.6037
R51 minus.n20 minus.n19 80.6037
R52 minus.n11 minus.n10 80.6037
R53 minus.n68 minus.n67 80.6037
R54 minus.n66 minus.n37 80.6037
R55 minus.n57 minus.n40 80.6037
R56 minus.n56 minus.n55 80.6037
R57 minus.n47 minus.n46 80.6037
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n20 minus.n5 41.6278
R69 minus.n22 minus.n21 41.6278
R70 minus.n56 minus.n41 41.6278
R71 minus.n58 minus.n57 41.6278
R72 minus.n33 minus.n32 38.7066
R73 minus.n69 minus.n68 38.7066
R74 minus.n72 minus.n35 38.5763
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 drain_right.n7 drain_right.n5 68.1648
R132 drain_right.n2 drain_right.n0 68.1648
R133 drain_right.n13 drain_right.n11 68.1648
R134 drain_right.n13 drain_right.n12 67.1908
R135 drain_right.n15 drain_right.n14 67.1908
R136 drain_right.n17 drain_right.n16 67.1908
R137 drain_right.n19 drain_right.n18 67.1908
R138 drain_right.n21 drain_right.n20 67.1908
R139 drain_right.n7 drain_right.n6 67.1907
R140 drain_right.n9 drain_right.n8 67.1907
R141 drain_right.n4 drain_right.n3 67.1907
R142 drain_right.n2 drain_right.n1 67.1907
R143 drain_right drain_right.n10 31.5227
R144 drain_right drain_right.n21 6.62735
R145 drain_right.n5 drain_right.t16 3.3005
R146 drain_right.n5 drain_right.t22 3.3005
R147 drain_right.n6 drain_right.t2 3.3005
R148 drain_right.n6 drain_right.t15 3.3005
R149 drain_right.n8 drain_right.t1 3.3005
R150 drain_right.n8 drain_right.t17 3.3005
R151 drain_right.n3 drain_right.t20 3.3005
R152 drain_right.n3 drain_right.t21 3.3005
R153 drain_right.n1 drain_right.t3 3.3005
R154 drain_right.n1 drain_right.t18 3.3005
R155 drain_right.n0 drain_right.t6 3.3005
R156 drain_right.n0 drain_right.t5 3.3005
R157 drain_right.n11 drain_right.t19 3.3005
R158 drain_right.n11 drain_right.t8 3.3005
R159 drain_right.n12 drain_right.t7 3.3005
R160 drain_right.n12 drain_right.t14 3.3005
R161 drain_right.n14 drain_right.t10 3.3005
R162 drain_right.n14 drain_right.t4 3.3005
R163 drain_right.n16 drain_right.t11 3.3005
R164 drain_right.n16 drain_right.t13 3.3005
R165 drain_right.n18 drain_right.t0 3.3005
R166 drain_right.n18 drain_right.t9 3.3005
R167 drain_right.n20 drain_right.t12 3.3005
R168 drain_right.n20 drain_right.t23 3.3005
R169 drain_right.n9 drain_right.n7 0.974638
R170 drain_right.n4 drain_right.n2 0.974638
R171 drain_right.n21 drain_right.n19 0.974638
R172 drain_right.n19 drain_right.n17 0.974638
R173 drain_right.n17 drain_right.n15 0.974638
R174 drain_right.n15 drain_right.n13 0.974638
R175 drain_right.n10 drain_right.n9 0.432223
R176 drain_right.n10 drain_right.n4 0.432223
R177 source.n290 source.n264 289.615
R178 source.n248 source.n222 289.615
R179 source.n216 source.n190 289.615
R180 source.n174 source.n148 289.615
R181 source.n26 source.n0 289.615
R182 source.n68 source.n42 289.615
R183 source.n100 source.n74 289.615
R184 source.n142 source.n116 289.615
R185 source.n275 source.n274 185
R186 source.n272 source.n271 185
R187 source.n281 source.n280 185
R188 source.n283 source.n282 185
R189 source.n268 source.n267 185
R190 source.n289 source.n288 185
R191 source.n291 source.n290 185
R192 source.n233 source.n232 185
R193 source.n230 source.n229 185
R194 source.n239 source.n238 185
R195 source.n241 source.n240 185
R196 source.n226 source.n225 185
R197 source.n247 source.n246 185
R198 source.n249 source.n248 185
R199 source.n201 source.n200 185
R200 source.n198 source.n197 185
R201 source.n207 source.n206 185
R202 source.n209 source.n208 185
R203 source.n194 source.n193 185
R204 source.n215 source.n214 185
R205 source.n217 source.n216 185
R206 source.n159 source.n158 185
R207 source.n156 source.n155 185
R208 source.n165 source.n164 185
R209 source.n167 source.n166 185
R210 source.n152 source.n151 185
R211 source.n173 source.n172 185
R212 source.n175 source.n174 185
R213 source.n27 source.n26 185
R214 source.n25 source.n24 185
R215 source.n4 source.n3 185
R216 source.n19 source.n18 185
R217 source.n17 source.n16 185
R218 source.n8 source.n7 185
R219 source.n11 source.n10 185
R220 source.n69 source.n68 185
R221 source.n67 source.n66 185
R222 source.n46 source.n45 185
R223 source.n61 source.n60 185
R224 source.n59 source.n58 185
R225 source.n50 source.n49 185
R226 source.n53 source.n52 185
R227 source.n101 source.n100 185
R228 source.n99 source.n98 185
R229 source.n78 source.n77 185
R230 source.n93 source.n92 185
R231 source.n91 source.n90 185
R232 source.n82 source.n81 185
R233 source.n85 source.n84 185
R234 source.n143 source.n142 185
R235 source.n141 source.n140 185
R236 source.n120 source.n119 185
R237 source.n135 source.n134 185
R238 source.n133 source.n132 185
R239 source.n124 source.n123 185
R240 source.n127 source.n126 185
R241 source.t40 source.n273 147.661
R242 source.t34 source.n231 147.661
R243 source.t12 source.n199 147.661
R244 source.t1 source.n157 147.661
R245 source.t5 source.n9 147.661
R246 source.t15 source.n51 147.661
R247 source.t33 source.n83 147.661
R248 source.t37 source.n125 147.661
R249 source.n274 source.n271 104.615
R250 source.n281 source.n271 104.615
R251 source.n282 source.n281 104.615
R252 source.n282 source.n267 104.615
R253 source.n289 source.n267 104.615
R254 source.n290 source.n289 104.615
R255 source.n232 source.n229 104.615
R256 source.n239 source.n229 104.615
R257 source.n240 source.n239 104.615
R258 source.n240 source.n225 104.615
R259 source.n247 source.n225 104.615
R260 source.n248 source.n247 104.615
R261 source.n200 source.n197 104.615
R262 source.n207 source.n197 104.615
R263 source.n208 source.n207 104.615
R264 source.n208 source.n193 104.615
R265 source.n215 source.n193 104.615
R266 source.n216 source.n215 104.615
R267 source.n158 source.n155 104.615
R268 source.n165 source.n155 104.615
R269 source.n166 source.n165 104.615
R270 source.n166 source.n151 104.615
R271 source.n173 source.n151 104.615
R272 source.n174 source.n173 104.615
R273 source.n26 source.n25 104.615
R274 source.n25 source.n3 104.615
R275 source.n18 source.n3 104.615
R276 source.n18 source.n17 104.615
R277 source.n17 source.n7 104.615
R278 source.n10 source.n7 104.615
R279 source.n68 source.n67 104.615
R280 source.n67 source.n45 104.615
R281 source.n60 source.n45 104.615
R282 source.n60 source.n59 104.615
R283 source.n59 source.n49 104.615
R284 source.n52 source.n49 104.615
R285 source.n100 source.n99 104.615
R286 source.n99 source.n77 104.615
R287 source.n92 source.n77 104.615
R288 source.n92 source.n91 104.615
R289 source.n91 source.n81 104.615
R290 source.n84 source.n81 104.615
R291 source.n142 source.n141 104.615
R292 source.n141 source.n119 104.615
R293 source.n134 source.n119 104.615
R294 source.n134 source.n133 104.615
R295 source.n133 source.n123 104.615
R296 source.n126 source.n123 104.615
R297 source.n274 source.t40 52.3082
R298 source.n232 source.t34 52.3082
R299 source.n200 source.t12 52.3082
R300 source.n158 source.t1 52.3082
R301 source.n10 source.t5 52.3082
R302 source.n52 source.t15 52.3082
R303 source.n84 source.t33 52.3082
R304 source.n126 source.t37 52.3082
R305 source.n33 source.n32 50.512
R306 source.n35 source.n34 50.512
R307 source.n37 source.n36 50.512
R308 source.n39 source.n38 50.512
R309 source.n41 source.n40 50.512
R310 source.n107 source.n106 50.512
R311 source.n109 source.n108 50.512
R312 source.n111 source.n110 50.512
R313 source.n113 source.n112 50.512
R314 source.n115 source.n114 50.512
R315 source.n263 source.n262 50.5119
R316 source.n261 source.n260 50.5119
R317 source.n259 source.n258 50.5119
R318 source.n257 source.n256 50.5119
R319 source.n255 source.n254 50.5119
R320 source.n189 source.n188 50.5119
R321 source.n187 source.n186 50.5119
R322 source.n185 source.n184 50.5119
R323 source.n183 source.n182 50.5119
R324 source.n181 source.n180 50.5119
R325 source.n295 source.n294 32.1853
R326 source.n253 source.n252 32.1853
R327 source.n221 source.n220 32.1853
R328 source.n179 source.n178 32.1853
R329 source.n31 source.n30 32.1853
R330 source.n73 source.n72 32.1853
R331 source.n105 source.n104 32.1853
R332 source.n147 source.n146 32.1853
R333 source.n179 source.n147 17.7164
R334 source.n275 source.n273 15.6674
R335 source.n233 source.n231 15.6674
R336 source.n201 source.n199 15.6674
R337 source.n159 source.n157 15.6674
R338 source.n11 source.n9 15.6674
R339 source.n53 source.n51 15.6674
R340 source.n85 source.n83 15.6674
R341 source.n127 source.n125 15.6674
R342 source.n276 source.n272 12.8005
R343 source.n234 source.n230 12.8005
R344 source.n202 source.n198 12.8005
R345 source.n160 source.n156 12.8005
R346 source.n12 source.n8 12.8005
R347 source.n54 source.n50 12.8005
R348 source.n86 source.n82 12.8005
R349 source.n128 source.n124 12.8005
R350 source.n280 source.n279 12.0247
R351 source.n238 source.n237 12.0247
R352 source.n206 source.n205 12.0247
R353 source.n164 source.n163 12.0247
R354 source.n16 source.n15 12.0247
R355 source.n58 source.n57 12.0247
R356 source.n90 source.n89 12.0247
R357 source.n132 source.n131 12.0247
R358 source.n296 source.n31 11.9664
R359 source.n283 source.n270 11.249
R360 source.n241 source.n228 11.249
R361 source.n209 source.n196 11.249
R362 source.n167 source.n154 11.249
R363 source.n19 source.n6 11.249
R364 source.n61 source.n48 11.249
R365 source.n93 source.n80 11.249
R366 source.n135 source.n122 11.249
R367 source.n284 source.n268 10.4732
R368 source.n242 source.n226 10.4732
R369 source.n210 source.n194 10.4732
R370 source.n168 source.n152 10.4732
R371 source.n20 source.n4 10.4732
R372 source.n62 source.n46 10.4732
R373 source.n94 source.n78 10.4732
R374 source.n136 source.n120 10.4732
R375 source.n288 source.n287 9.69747
R376 source.n246 source.n245 9.69747
R377 source.n214 source.n213 9.69747
R378 source.n172 source.n171 9.69747
R379 source.n24 source.n23 9.69747
R380 source.n66 source.n65 9.69747
R381 source.n98 source.n97 9.69747
R382 source.n140 source.n139 9.69747
R383 source.n294 source.n293 9.45567
R384 source.n252 source.n251 9.45567
R385 source.n220 source.n219 9.45567
R386 source.n178 source.n177 9.45567
R387 source.n30 source.n29 9.45567
R388 source.n72 source.n71 9.45567
R389 source.n104 source.n103 9.45567
R390 source.n146 source.n145 9.45567
R391 source.n293 source.n292 9.3005
R392 source.n266 source.n265 9.3005
R393 source.n287 source.n286 9.3005
R394 source.n285 source.n284 9.3005
R395 source.n270 source.n269 9.3005
R396 source.n279 source.n278 9.3005
R397 source.n277 source.n276 9.3005
R398 source.n251 source.n250 9.3005
R399 source.n224 source.n223 9.3005
R400 source.n245 source.n244 9.3005
R401 source.n243 source.n242 9.3005
R402 source.n228 source.n227 9.3005
R403 source.n237 source.n236 9.3005
R404 source.n235 source.n234 9.3005
R405 source.n219 source.n218 9.3005
R406 source.n192 source.n191 9.3005
R407 source.n213 source.n212 9.3005
R408 source.n211 source.n210 9.3005
R409 source.n196 source.n195 9.3005
R410 source.n205 source.n204 9.3005
R411 source.n203 source.n202 9.3005
R412 source.n177 source.n176 9.3005
R413 source.n150 source.n149 9.3005
R414 source.n171 source.n170 9.3005
R415 source.n169 source.n168 9.3005
R416 source.n154 source.n153 9.3005
R417 source.n163 source.n162 9.3005
R418 source.n161 source.n160 9.3005
R419 source.n29 source.n28 9.3005
R420 source.n2 source.n1 9.3005
R421 source.n23 source.n22 9.3005
R422 source.n21 source.n20 9.3005
R423 source.n6 source.n5 9.3005
R424 source.n15 source.n14 9.3005
R425 source.n13 source.n12 9.3005
R426 source.n71 source.n70 9.3005
R427 source.n44 source.n43 9.3005
R428 source.n65 source.n64 9.3005
R429 source.n63 source.n62 9.3005
R430 source.n48 source.n47 9.3005
R431 source.n57 source.n56 9.3005
R432 source.n55 source.n54 9.3005
R433 source.n103 source.n102 9.3005
R434 source.n76 source.n75 9.3005
R435 source.n97 source.n96 9.3005
R436 source.n95 source.n94 9.3005
R437 source.n80 source.n79 9.3005
R438 source.n89 source.n88 9.3005
R439 source.n87 source.n86 9.3005
R440 source.n145 source.n144 9.3005
R441 source.n118 source.n117 9.3005
R442 source.n139 source.n138 9.3005
R443 source.n137 source.n136 9.3005
R444 source.n122 source.n121 9.3005
R445 source.n131 source.n130 9.3005
R446 source.n129 source.n128 9.3005
R447 source.n291 source.n266 8.92171
R448 source.n249 source.n224 8.92171
R449 source.n217 source.n192 8.92171
R450 source.n175 source.n150 8.92171
R451 source.n27 source.n2 8.92171
R452 source.n69 source.n44 8.92171
R453 source.n101 source.n76 8.92171
R454 source.n143 source.n118 8.92171
R455 source.n292 source.n264 8.14595
R456 source.n250 source.n222 8.14595
R457 source.n218 source.n190 8.14595
R458 source.n176 source.n148 8.14595
R459 source.n28 source.n0 8.14595
R460 source.n70 source.n42 8.14595
R461 source.n102 source.n74 8.14595
R462 source.n144 source.n116 8.14595
R463 source.n294 source.n264 5.81868
R464 source.n252 source.n222 5.81868
R465 source.n220 source.n190 5.81868
R466 source.n178 source.n148 5.81868
R467 source.n30 source.n0 5.81868
R468 source.n72 source.n42 5.81868
R469 source.n104 source.n74 5.81868
R470 source.n146 source.n116 5.81868
R471 source.n296 source.n295 5.7505
R472 source.n292 source.n291 5.04292
R473 source.n250 source.n249 5.04292
R474 source.n218 source.n217 5.04292
R475 source.n176 source.n175 5.04292
R476 source.n28 source.n27 5.04292
R477 source.n70 source.n69 5.04292
R478 source.n102 source.n101 5.04292
R479 source.n144 source.n143 5.04292
R480 source.n277 source.n273 4.38594
R481 source.n235 source.n231 4.38594
R482 source.n203 source.n199 4.38594
R483 source.n161 source.n157 4.38594
R484 source.n13 source.n9 4.38594
R485 source.n55 source.n51 4.38594
R486 source.n87 source.n83 4.38594
R487 source.n129 source.n125 4.38594
R488 source.n288 source.n266 4.26717
R489 source.n246 source.n224 4.26717
R490 source.n214 source.n192 4.26717
R491 source.n172 source.n150 4.26717
R492 source.n24 source.n2 4.26717
R493 source.n66 source.n44 4.26717
R494 source.n98 source.n76 4.26717
R495 source.n140 source.n118 4.26717
R496 source.n287 source.n268 3.49141
R497 source.n245 source.n226 3.49141
R498 source.n213 source.n194 3.49141
R499 source.n171 source.n152 3.49141
R500 source.n23 source.n4 3.49141
R501 source.n65 source.n46 3.49141
R502 source.n97 source.n78 3.49141
R503 source.n139 source.n120 3.49141
R504 source.n262 source.t27 3.3005
R505 source.n262 source.t47 3.3005
R506 source.n260 source.t31 3.3005
R507 source.n260 source.t43 3.3005
R508 source.n258 source.t25 3.3005
R509 source.n258 source.t45 3.3005
R510 source.n256 source.t24 3.3005
R511 source.n256 source.t39 3.3005
R512 source.n254 source.t46 3.3005
R513 source.n254 source.t42 3.3005
R514 source.n188 source.t3 3.3005
R515 source.n188 source.t8 3.3005
R516 source.n186 source.t0 3.3005
R517 source.n186 source.t22 3.3005
R518 source.n184 source.t19 3.3005
R519 source.n184 source.t18 3.3005
R520 source.n182 source.t7 3.3005
R521 source.n182 source.t4 3.3005
R522 source.n180 source.t17 3.3005
R523 source.n180 source.t11 3.3005
R524 source.n32 source.t10 3.3005
R525 source.n32 source.t23 3.3005
R526 source.n34 source.t21 3.3005
R527 source.n34 source.t20 3.3005
R528 source.n36 source.t6 3.3005
R529 source.n36 source.t13 3.3005
R530 source.n38 source.t2 3.3005
R531 source.n38 source.t16 3.3005
R532 source.n40 source.t9 3.3005
R533 source.n40 source.t14 3.3005
R534 source.n106 source.t41 3.3005
R535 source.n106 source.t38 3.3005
R536 source.n108 source.t28 3.3005
R537 source.n108 source.t30 3.3005
R538 source.n110 source.t36 3.3005
R539 source.n110 source.t32 3.3005
R540 source.n112 source.t29 3.3005
R541 source.n112 source.t26 3.3005
R542 source.n114 source.t35 3.3005
R543 source.n114 source.t44 3.3005
R544 source.n284 source.n283 2.71565
R545 source.n242 source.n241 2.71565
R546 source.n210 source.n209 2.71565
R547 source.n168 source.n167 2.71565
R548 source.n20 source.n19 2.71565
R549 source.n62 source.n61 2.71565
R550 source.n94 source.n93 2.71565
R551 source.n136 source.n135 2.71565
R552 source.n280 source.n270 1.93989
R553 source.n238 source.n228 1.93989
R554 source.n206 source.n196 1.93989
R555 source.n164 source.n154 1.93989
R556 source.n16 source.n6 1.93989
R557 source.n58 source.n48 1.93989
R558 source.n90 source.n80 1.93989
R559 source.n132 source.n122 1.93989
R560 source.n279 source.n272 1.16414
R561 source.n237 source.n230 1.16414
R562 source.n205 source.n198 1.16414
R563 source.n163 source.n156 1.16414
R564 source.n15 source.n8 1.16414
R565 source.n57 source.n50 1.16414
R566 source.n89 source.n82 1.16414
R567 source.n131 source.n124 1.16414
R568 source.n147 source.n115 0.974638
R569 source.n115 source.n113 0.974638
R570 source.n113 source.n111 0.974638
R571 source.n111 source.n109 0.974638
R572 source.n109 source.n107 0.974638
R573 source.n107 source.n105 0.974638
R574 source.n73 source.n41 0.974638
R575 source.n41 source.n39 0.974638
R576 source.n39 source.n37 0.974638
R577 source.n37 source.n35 0.974638
R578 source.n35 source.n33 0.974638
R579 source.n33 source.n31 0.974638
R580 source.n181 source.n179 0.974638
R581 source.n183 source.n181 0.974638
R582 source.n185 source.n183 0.974638
R583 source.n187 source.n185 0.974638
R584 source.n189 source.n187 0.974638
R585 source.n221 source.n189 0.974638
R586 source.n255 source.n253 0.974638
R587 source.n257 source.n255 0.974638
R588 source.n259 source.n257 0.974638
R589 source.n261 source.n259 0.974638
R590 source.n263 source.n261 0.974638
R591 source.n295 source.n263 0.974638
R592 source.n105 source.n73 0.470328
R593 source.n253 source.n221 0.470328
R594 source.n276 source.n275 0.388379
R595 source.n234 source.n233 0.388379
R596 source.n202 source.n201 0.388379
R597 source.n160 source.n159 0.388379
R598 source.n12 source.n11 0.388379
R599 source.n54 source.n53 0.388379
R600 source.n86 source.n85 0.388379
R601 source.n128 source.n127 0.388379
R602 source source.n296 0.188
R603 source.n278 source.n277 0.155672
R604 source.n278 source.n269 0.155672
R605 source.n285 source.n269 0.155672
R606 source.n286 source.n285 0.155672
R607 source.n286 source.n265 0.155672
R608 source.n293 source.n265 0.155672
R609 source.n236 source.n235 0.155672
R610 source.n236 source.n227 0.155672
R611 source.n243 source.n227 0.155672
R612 source.n244 source.n243 0.155672
R613 source.n244 source.n223 0.155672
R614 source.n251 source.n223 0.155672
R615 source.n204 source.n203 0.155672
R616 source.n204 source.n195 0.155672
R617 source.n211 source.n195 0.155672
R618 source.n212 source.n211 0.155672
R619 source.n212 source.n191 0.155672
R620 source.n219 source.n191 0.155672
R621 source.n162 source.n161 0.155672
R622 source.n162 source.n153 0.155672
R623 source.n169 source.n153 0.155672
R624 source.n170 source.n169 0.155672
R625 source.n170 source.n149 0.155672
R626 source.n177 source.n149 0.155672
R627 source.n29 source.n1 0.155672
R628 source.n22 source.n1 0.155672
R629 source.n22 source.n21 0.155672
R630 source.n21 source.n5 0.155672
R631 source.n14 source.n5 0.155672
R632 source.n14 source.n13 0.155672
R633 source.n71 source.n43 0.155672
R634 source.n64 source.n43 0.155672
R635 source.n64 source.n63 0.155672
R636 source.n63 source.n47 0.155672
R637 source.n56 source.n47 0.155672
R638 source.n56 source.n55 0.155672
R639 source.n103 source.n75 0.155672
R640 source.n96 source.n75 0.155672
R641 source.n96 source.n95 0.155672
R642 source.n95 source.n79 0.155672
R643 source.n88 source.n79 0.155672
R644 source.n88 source.n87 0.155672
R645 source.n145 source.n117 0.155672
R646 source.n138 source.n117 0.155672
R647 source.n138 source.n137 0.155672
R648 source.n137 source.n121 0.155672
R649 source.n130 source.n121 0.155672
R650 source.n130 source.n129 0.155672
R651 plus.n10 plus.t22 251.291
R652 plus.n46 plus.t9 251.291
R653 plus.n34 plus.t6 229.855
R654 plus.n32 plus.t8 229.855
R655 plus.n31 plus.t10 229.855
R656 plus.n3 plus.t13 229.855
R657 plus.n25 plus.t14 229.855
R658 plus.n5 plus.t15 229.855
R659 plus.n20 plus.t17 229.855
R660 plus.n18 plus.t20 229.855
R661 plus.n8 plus.t18 229.855
R662 plus.n12 plus.t19 229.855
R663 plus.n11 plus.t21 229.855
R664 plus.n70 plus.t12 229.855
R665 plus.n68 plus.t2 229.855
R666 plus.n67 plus.t7 229.855
R667 plus.n39 plus.t1 229.855
R668 plus.n61 plus.t16 229.855
R669 plus.n41 plus.t3 229.855
R670 plus.n56 plus.t11 229.855
R671 plus.n54 plus.t5 229.855
R672 plus.n44 plus.t23 229.855
R673 plus.n48 plus.t4 229.855
R674 plus.n47 plus.t0 229.855
R675 plus.n14 plus.n13 161.3
R676 plus.n15 plus.n8 161.3
R677 plus.n17 plus.n16 161.3
R678 plus.n18 plus.n7 161.3
R679 plus.n19 plus.n6 161.3
R680 plus.n24 plus.n23 161.3
R681 plus.n25 plus.n4 161.3
R682 plus.n27 plus.n26 161.3
R683 plus.n28 plus.n3 161.3
R684 plus.n30 plus.n29 161.3
R685 plus.n33 plus.n0 161.3
R686 plus.n35 plus.n34 161.3
R687 plus.n50 plus.n49 161.3
R688 plus.n51 plus.n44 161.3
R689 plus.n53 plus.n52 161.3
R690 plus.n54 plus.n43 161.3
R691 plus.n55 plus.n42 161.3
R692 plus.n60 plus.n59 161.3
R693 plus.n61 plus.n40 161.3
R694 plus.n63 plus.n62 161.3
R695 plus.n64 plus.n39 161.3
R696 plus.n66 plus.n65 161.3
R697 plus.n69 plus.n36 161.3
R698 plus.n71 plus.n70 161.3
R699 plus.n12 plus.n9 80.6037
R700 plus.n21 plus.n20 80.6037
R701 plus.n22 plus.n5 80.6037
R702 plus.n31 plus.n2 80.6037
R703 plus.n32 plus.n1 80.6037
R704 plus.n48 plus.n45 80.6037
R705 plus.n57 plus.n56 80.6037
R706 plus.n58 plus.n41 80.6037
R707 plus.n67 plus.n38 80.6037
R708 plus.n68 plus.n37 80.6037
R709 plus.n32 plus.n31 48.2005
R710 plus.n20 plus.n5 48.2005
R711 plus.n12 plus.n11 48.2005
R712 plus.n68 plus.n67 48.2005
R713 plus.n56 plus.n41 48.2005
R714 plus.n48 plus.n47 48.2005
R715 plus.n31 plus.n30 44.549
R716 plus.n13 plus.n12 44.549
R717 plus.n67 plus.n66 44.549
R718 plus.n49 plus.n48 44.549
R719 plus.n24 plus.n5 41.6278
R720 plus.n20 plus.n19 41.6278
R721 plus.n60 plus.n41 41.6278
R722 plus.n56 plus.n55 41.6278
R723 plus.n33 plus.n32 38.7066
R724 plus.n69 plus.n68 38.7066
R725 plus plus.n71 34.7301
R726 plus.n10 plus.n9 31.6825
R727 plus.n46 plus.n45 31.6825
R728 plus.n26 plus.n3 25.5611
R729 plus.n17 plus.n8 25.5611
R730 plus.n62 plus.n39 25.5611
R731 plus.n53 plus.n44 25.5611
R732 plus.n26 plus.n25 22.6399
R733 plus.n18 plus.n17 22.6399
R734 plus.n62 plus.n61 22.6399
R735 plus.n54 plus.n53 22.6399
R736 plus.n11 plus.n10 17.2341
R737 plus.n47 plus.n46 17.2341
R738 plus plus.n35 10.0308
R739 plus.n34 plus.n33 9.49444
R740 plus.n70 plus.n69 9.49444
R741 plus.n25 plus.n24 6.57323
R742 plus.n19 plus.n18 6.57323
R743 plus.n61 plus.n60 6.57323
R744 plus.n55 plus.n54 6.57323
R745 plus.n30 plus.n3 3.65202
R746 plus.n13 plus.n8 3.65202
R747 plus.n66 plus.n39 3.65202
R748 plus.n49 plus.n44 3.65202
R749 plus.n22 plus.n21 0.380177
R750 plus.n2 plus.n1 0.380177
R751 plus.n38 plus.n37 0.380177
R752 plus.n58 plus.n57 0.380177
R753 plus.n14 plus.n9 0.285035
R754 plus.n21 plus.n6 0.285035
R755 plus.n23 plus.n22 0.285035
R756 plus.n29 plus.n2 0.285035
R757 plus.n1 plus.n0 0.285035
R758 plus.n37 plus.n36 0.285035
R759 plus.n65 plus.n38 0.285035
R760 plus.n59 plus.n58 0.285035
R761 plus.n57 plus.n42 0.285035
R762 plus.n50 plus.n45 0.285035
R763 plus.n15 plus.n14 0.189894
R764 plus.n16 plus.n15 0.189894
R765 plus.n16 plus.n7 0.189894
R766 plus.n7 plus.n6 0.189894
R767 plus.n23 plus.n4 0.189894
R768 plus.n27 plus.n4 0.189894
R769 plus.n28 plus.n27 0.189894
R770 plus.n29 plus.n28 0.189894
R771 plus.n35 plus.n0 0.189894
R772 plus.n71 plus.n36 0.189894
R773 plus.n65 plus.n64 0.189894
R774 plus.n64 plus.n63 0.189894
R775 plus.n63 plus.n40 0.189894
R776 plus.n59 plus.n40 0.189894
R777 plus.n43 plus.n42 0.189894
R778 plus.n52 plus.n43 0.189894
R779 plus.n52 plus.n51 0.189894
R780 plus.n51 plus.n50 0.189894
R781 drain_left.n13 drain_left.n11 68.165
R782 drain_left.n7 drain_left.n5 68.1648
R783 drain_left.n2 drain_left.n0 68.1648
R784 drain_left.n19 drain_left.n18 67.1908
R785 drain_left.n17 drain_left.n16 67.1908
R786 drain_left.n15 drain_left.n14 67.1908
R787 drain_left.n13 drain_left.n12 67.1908
R788 drain_left.n21 drain_left.n20 67.1907
R789 drain_left.n7 drain_left.n6 67.1907
R790 drain_left.n9 drain_left.n8 67.1907
R791 drain_left.n4 drain_left.n3 67.1907
R792 drain_left.n2 drain_left.n1 67.1907
R793 drain_left drain_left.n10 32.0759
R794 drain_left drain_left.n21 6.62735
R795 drain_left.n5 drain_left.t23 3.3005
R796 drain_left.n5 drain_left.t14 3.3005
R797 drain_left.n6 drain_left.t0 3.3005
R798 drain_left.n6 drain_left.t19 3.3005
R799 drain_left.n8 drain_left.t12 3.3005
R800 drain_left.n8 drain_left.t18 3.3005
R801 drain_left.n3 drain_left.t7 3.3005
R802 drain_left.n3 drain_left.t20 3.3005
R803 drain_left.n1 drain_left.t16 3.3005
R804 drain_left.n1 drain_left.t22 3.3005
R805 drain_left.n0 drain_left.t11 3.3005
R806 drain_left.n0 drain_left.t21 3.3005
R807 drain_left.n20 drain_left.t15 3.3005
R808 drain_left.n20 drain_left.t17 3.3005
R809 drain_left.n18 drain_left.t10 3.3005
R810 drain_left.n18 drain_left.t13 3.3005
R811 drain_left.n16 drain_left.t8 3.3005
R812 drain_left.n16 drain_left.t9 3.3005
R813 drain_left.n14 drain_left.t3 3.3005
R814 drain_left.n14 drain_left.t6 3.3005
R815 drain_left.n12 drain_left.t4 3.3005
R816 drain_left.n12 drain_left.t5 3.3005
R817 drain_left.n11 drain_left.t1 3.3005
R818 drain_left.n11 drain_left.t2 3.3005
R819 drain_left.n9 drain_left.n7 0.974638
R820 drain_left.n4 drain_left.n2 0.974638
R821 drain_left.n15 drain_left.n13 0.974638
R822 drain_left.n17 drain_left.n15 0.974638
R823 drain_left.n19 drain_left.n17 0.974638
R824 drain_left.n21 drain_left.n19 0.974638
R825 drain_left.n10 drain_left.n9 0.432223
R826 drain_left.n10 drain_left.n4 0.432223
C0 drain_left source 15.7426f
C1 drain_right minus 8.43596f
C2 plus minus 6.59768f
C3 drain_right plus 0.526806f
C4 drain_left minus 0.175388f
C5 drain_right drain_left 2.02887f
C6 drain_left plus 8.803451f
C7 source minus 9.218071f
C8 drain_right source 15.745701f
C9 source plus 9.23209f
C10 drain_right a_n3654_n2088# 7.20867f
C11 drain_left a_n3654_n2088# 7.72614f
C12 source a_n3654_n2088# 6.050945f
C13 minus a_n3654_n2088# 14.308546f
C14 plus a_n3654_n2088# 15.90264f
C15 drain_left.t11 a_n3654_n2088# 0.137069f
C16 drain_left.t21 a_n3654_n2088# 0.137069f
C17 drain_left.n0 a_n3654_n2088# 1.14927f
C18 drain_left.t16 a_n3654_n2088# 0.137069f
C19 drain_left.t22 a_n3654_n2088# 0.137069f
C20 drain_left.n1 a_n3654_n2088# 1.14316f
C21 drain_left.n2 a_n3654_n2088# 0.837773f
C22 drain_left.t7 a_n3654_n2088# 0.137069f
C23 drain_left.t20 a_n3654_n2088# 0.137069f
C24 drain_left.n3 a_n3654_n2088# 1.14316f
C25 drain_left.n4 a_n3654_n2088# 0.367147f
C26 drain_left.t23 a_n3654_n2088# 0.137069f
C27 drain_left.t14 a_n3654_n2088# 0.137069f
C28 drain_left.n5 a_n3654_n2088# 1.14927f
C29 drain_left.t0 a_n3654_n2088# 0.137069f
C30 drain_left.t19 a_n3654_n2088# 0.137069f
C31 drain_left.n6 a_n3654_n2088# 1.14316f
C32 drain_left.n7 a_n3654_n2088# 0.837773f
C33 drain_left.t12 a_n3654_n2088# 0.137069f
C34 drain_left.t18 a_n3654_n2088# 0.137069f
C35 drain_left.n8 a_n3654_n2088# 1.14316f
C36 drain_left.n9 a_n3654_n2088# 0.367147f
C37 drain_left.n10 a_n3654_n2088# 1.60691f
C38 drain_left.t1 a_n3654_n2088# 0.137069f
C39 drain_left.t2 a_n3654_n2088# 0.137069f
C40 drain_left.n11 a_n3654_n2088# 1.14927f
C41 drain_left.t4 a_n3654_n2088# 0.137069f
C42 drain_left.t5 a_n3654_n2088# 0.137069f
C43 drain_left.n12 a_n3654_n2088# 1.14316f
C44 drain_left.n13 a_n3654_n2088# 0.837762f
C45 drain_left.t3 a_n3654_n2088# 0.137069f
C46 drain_left.t6 a_n3654_n2088# 0.137069f
C47 drain_left.n14 a_n3654_n2088# 1.14316f
C48 drain_left.n15 a_n3654_n2088# 0.416116f
C49 drain_left.t8 a_n3654_n2088# 0.137069f
C50 drain_left.t9 a_n3654_n2088# 0.137069f
C51 drain_left.n16 a_n3654_n2088# 1.14316f
C52 drain_left.n17 a_n3654_n2088# 0.416116f
C53 drain_left.t10 a_n3654_n2088# 0.137069f
C54 drain_left.t13 a_n3654_n2088# 0.137069f
C55 drain_left.n18 a_n3654_n2088# 1.14316f
C56 drain_left.n19 a_n3654_n2088# 0.416116f
C57 drain_left.t15 a_n3654_n2088# 0.137069f
C58 drain_left.t17 a_n3654_n2088# 0.137069f
C59 drain_left.n20 a_n3654_n2088# 1.14316f
C60 drain_left.n21 a_n3654_n2088# 0.675347f
C61 plus.n0 a_n3654_n2088# 0.051693f
C62 plus.t6 a_n3654_n2088# 0.539361f
C63 plus.t8 a_n3654_n2088# 0.539361f
C64 plus.n1 a_n3654_n2088# 0.064526f
C65 plus.t10 a_n3654_n2088# 0.539361f
C66 plus.n2 a_n3654_n2088# 0.064526f
C67 plus.t13 a_n3654_n2088# 0.539361f
C68 plus.n3 a_n3654_n2088# 0.245692f
C69 plus.n4 a_n3654_n2088# 0.03874f
C70 plus.t14 a_n3654_n2088# 0.539361f
C71 plus.t15 a_n3654_n2088# 0.539361f
C72 plus.n5 a_n3654_n2088# 0.256513f
C73 plus.n6 a_n3654_n2088# 0.051693f
C74 plus.t17 a_n3654_n2088# 0.539361f
C75 plus.t20 a_n3654_n2088# 0.539361f
C76 plus.n7 a_n3654_n2088# 0.03874f
C77 plus.t18 a_n3654_n2088# 0.539361f
C78 plus.n8 a_n3654_n2088# 0.245692f
C79 plus.n9 a_n3654_n2088# 0.222662f
C80 plus.t19 a_n3654_n2088# 0.539361f
C81 plus.t21 a_n3654_n2088# 0.539361f
C82 plus.t22 a_n3654_n2088# 0.560599f
C83 plus.n10 a_n3654_n2088# 0.231402f
C84 plus.n11 a_n3654_n2088# 0.25697f
C85 plus.n12 a_n3654_n2088# 0.25699f
C86 plus.n13 a_n3654_n2088# 0.008791f
C87 plus.n14 a_n3654_n2088# 0.051693f
C88 plus.n15 a_n3654_n2088# 0.03874f
C89 plus.n16 a_n3654_n2088# 0.03874f
C90 plus.n17 a_n3654_n2088# 0.008791f
C91 plus.n18 a_n3654_n2088# 0.245692f
C92 plus.n19 a_n3654_n2088# 0.008791f
C93 plus.n20 a_n3654_n2088# 0.256513f
C94 plus.n21 a_n3654_n2088# 0.064526f
C95 plus.n22 a_n3654_n2088# 0.064526f
C96 plus.n23 a_n3654_n2088# 0.051693f
C97 plus.n24 a_n3654_n2088# 0.008791f
C98 plus.n25 a_n3654_n2088# 0.245692f
C99 plus.n26 a_n3654_n2088# 0.008791f
C100 plus.n27 a_n3654_n2088# 0.03874f
C101 plus.n28 a_n3654_n2088# 0.03874f
C102 plus.n29 a_n3654_n2088# 0.051693f
C103 plus.n30 a_n3654_n2088# 0.008791f
C104 plus.n31 a_n3654_n2088# 0.25699f
C105 plus.n32 a_n3654_n2088# 0.256035f
C106 plus.n33 a_n3654_n2088# 0.008791f
C107 plus.n34 a_n3654_n2088# 0.242467f
C108 plus.n35 a_n3654_n2088# 0.34707f
C109 plus.n36 a_n3654_n2088# 0.051693f
C110 plus.t12 a_n3654_n2088# 0.539361f
C111 plus.n37 a_n3654_n2088# 0.064526f
C112 plus.t2 a_n3654_n2088# 0.539361f
C113 plus.n38 a_n3654_n2088# 0.064526f
C114 plus.t7 a_n3654_n2088# 0.539361f
C115 plus.t1 a_n3654_n2088# 0.539361f
C116 plus.n39 a_n3654_n2088# 0.245692f
C117 plus.n40 a_n3654_n2088# 0.03874f
C118 plus.t16 a_n3654_n2088# 0.539361f
C119 plus.t3 a_n3654_n2088# 0.539361f
C120 plus.n41 a_n3654_n2088# 0.256513f
C121 plus.n42 a_n3654_n2088# 0.051693f
C122 plus.t11 a_n3654_n2088# 0.539361f
C123 plus.n43 a_n3654_n2088# 0.03874f
C124 plus.t5 a_n3654_n2088# 0.539361f
C125 plus.t23 a_n3654_n2088# 0.539361f
C126 plus.n44 a_n3654_n2088# 0.245692f
C127 plus.n45 a_n3654_n2088# 0.222662f
C128 plus.t4 a_n3654_n2088# 0.539361f
C129 plus.t9 a_n3654_n2088# 0.560599f
C130 plus.n46 a_n3654_n2088# 0.231402f
C131 plus.t0 a_n3654_n2088# 0.539361f
C132 plus.n47 a_n3654_n2088# 0.25697f
C133 plus.n48 a_n3654_n2088# 0.25699f
C134 plus.n49 a_n3654_n2088# 0.008791f
C135 plus.n50 a_n3654_n2088# 0.051693f
C136 plus.n51 a_n3654_n2088# 0.03874f
C137 plus.n52 a_n3654_n2088# 0.03874f
C138 plus.n53 a_n3654_n2088# 0.008791f
C139 plus.n54 a_n3654_n2088# 0.245692f
C140 plus.n55 a_n3654_n2088# 0.008791f
C141 plus.n56 a_n3654_n2088# 0.256513f
C142 plus.n57 a_n3654_n2088# 0.064526f
C143 plus.n58 a_n3654_n2088# 0.064526f
C144 plus.n59 a_n3654_n2088# 0.051693f
C145 plus.n60 a_n3654_n2088# 0.008791f
C146 plus.n61 a_n3654_n2088# 0.245692f
C147 plus.n62 a_n3654_n2088# 0.008791f
C148 plus.n63 a_n3654_n2088# 0.03874f
C149 plus.n64 a_n3654_n2088# 0.03874f
C150 plus.n65 a_n3654_n2088# 0.051693f
C151 plus.n66 a_n3654_n2088# 0.008791f
C152 plus.n67 a_n3654_n2088# 0.25699f
C153 plus.n68 a_n3654_n2088# 0.256035f
C154 plus.n69 a_n3654_n2088# 0.008791f
C155 plus.n70 a_n3654_n2088# 0.242467f
C156 plus.n71 a_n3654_n2088# 1.37862f
C157 source.n0 a_n3654_n2088# 0.036994f
C158 source.n1 a_n3654_n2088# 0.026319f
C159 source.n2 a_n3654_n2088# 0.014143f
C160 source.n3 a_n3654_n2088# 0.033429f
C161 source.n4 a_n3654_n2088# 0.014975f
C162 source.n5 a_n3654_n2088# 0.026319f
C163 source.n6 a_n3654_n2088# 0.014143f
C164 source.n7 a_n3654_n2088# 0.033429f
C165 source.n8 a_n3654_n2088# 0.014975f
C166 source.n9 a_n3654_n2088# 0.112628f
C167 source.t5 a_n3654_n2088# 0.054484f
C168 source.n10 a_n3654_n2088# 0.025071f
C169 source.n11 a_n3654_n2088# 0.019746f
C170 source.n12 a_n3654_n2088# 0.014143f
C171 source.n13 a_n3654_n2088# 0.626241f
C172 source.n14 a_n3654_n2088# 0.026319f
C173 source.n15 a_n3654_n2088# 0.014143f
C174 source.n16 a_n3654_n2088# 0.014975f
C175 source.n17 a_n3654_n2088# 0.033429f
C176 source.n18 a_n3654_n2088# 0.033429f
C177 source.n19 a_n3654_n2088# 0.014975f
C178 source.n20 a_n3654_n2088# 0.014143f
C179 source.n21 a_n3654_n2088# 0.026319f
C180 source.n22 a_n3654_n2088# 0.026319f
C181 source.n23 a_n3654_n2088# 0.014143f
C182 source.n24 a_n3654_n2088# 0.014975f
C183 source.n25 a_n3654_n2088# 0.033429f
C184 source.n26 a_n3654_n2088# 0.072367f
C185 source.n27 a_n3654_n2088# 0.014975f
C186 source.n28 a_n3654_n2088# 0.014143f
C187 source.n29 a_n3654_n2088# 0.060836f
C188 source.n30 a_n3654_n2088# 0.040492f
C189 source.n31 a_n3654_n2088# 0.700036f
C190 source.t10 a_n3654_n2088# 0.12479f
C191 source.t23 a_n3654_n2088# 0.12479f
C192 source.n32 a_n3654_n2088# 0.971871f
C193 source.n33 a_n3654_n2088# 0.411944f
C194 source.t21 a_n3654_n2088# 0.12479f
C195 source.t20 a_n3654_n2088# 0.12479f
C196 source.n34 a_n3654_n2088# 0.971871f
C197 source.n35 a_n3654_n2088# 0.411944f
C198 source.t6 a_n3654_n2088# 0.12479f
C199 source.t13 a_n3654_n2088# 0.12479f
C200 source.n36 a_n3654_n2088# 0.971871f
C201 source.n37 a_n3654_n2088# 0.411944f
C202 source.t2 a_n3654_n2088# 0.12479f
C203 source.t16 a_n3654_n2088# 0.12479f
C204 source.n38 a_n3654_n2088# 0.971871f
C205 source.n39 a_n3654_n2088# 0.411944f
C206 source.t9 a_n3654_n2088# 0.12479f
C207 source.t14 a_n3654_n2088# 0.12479f
C208 source.n40 a_n3654_n2088# 0.971871f
C209 source.n41 a_n3654_n2088# 0.411944f
C210 source.n42 a_n3654_n2088# 0.036994f
C211 source.n43 a_n3654_n2088# 0.026319f
C212 source.n44 a_n3654_n2088# 0.014143f
C213 source.n45 a_n3654_n2088# 0.033429f
C214 source.n46 a_n3654_n2088# 0.014975f
C215 source.n47 a_n3654_n2088# 0.026319f
C216 source.n48 a_n3654_n2088# 0.014143f
C217 source.n49 a_n3654_n2088# 0.033429f
C218 source.n50 a_n3654_n2088# 0.014975f
C219 source.n51 a_n3654_n2088# 0.112628f
C220 source.t15 a_n3654_n2088# 0.054484f
C221 source.n52 a_n3654_n2088# 0.025071f
C222 source.n53 a_n3654_n2088# 0.019746f
C223 source.n54 a_n3654_n2088# 0.014143f
C224 source.n55 a_n3654_n2088# 0.626241f
C225 source.n56 a_n3654_n2088# 0.026319f
C226 source.n57 a_n3654_n2088# 0.014143f
C227 source.n58 a_n3654_n2088# 0.014975f
C228 source.n59 a_n3654_n2088# 0.033429f
C229 source.n60 a_n3654_n2088# 0.033429f
C230 source.n61 a_n3654_n2088# 0.014975f
C231 source.n62 a_n3654_n2088# 0.014143f
C232 source.n63 a_n3654_n2088# 0.026319f
C233 source.n64 a_n3654_n2088# 0.026319f
C234 source.n65 a_n3654_n2088# 0.014143f
C235 source.n66 a_n3654_n2088# 0.014975f
C236 source.n67 a_n3654_n2088# 0.033429f
C237 source.n68 a_n3654_n2088# 0.072367f
C238 source.n69 a_n3654_n2088# 0.014975f
C239 source.n70 a_n3654_n2088# 0.014143f
C240 source.n71 a_n3654_n2088# 0.060836f
C241 source.n72 a_n3654_n2088# 0.040492f
C242 source.n73 a_n3654_n2088# 0.144936f
C243 source.n74 a_n3654_n2088# 0.036994f
C244 source.n75 a_n3654_n2088# 0.026319f
C245 source.n76 a_n3654_n2088# 0.014143f
C246 source.n77 a_n3654_n2088# 0.033429f
C247 source.n78 a_n3654_n2088# 0.014975f
C248 source.n79 a_n3654_n2088# 0.026319f
C249 source.n80 a_n3654_n2088# 0.014143f
C250 source.n81 a_n3654_n2088# 0.033429f
C251 source.n82 a_n3654_n2088# 0.014975f
C252 source.n83 a_n3654_n2088# 0.112628f
C253 source.t33 a_n3654_n2088# 0.054484f
C254 source.n84 a_n3654_n2088# 0.025071f
C255 source.n85 a_n3654_n2088# 0.019746f
C256 source.n86 a_n3654_n2088# 0.014143f
C257 source.n87 a_n3654_n2088# 0.626241f
C258 source.n88 a_n3654_n2088# 0.026319f
C259 source.n89 a_n3654_n2088# 0.014143f
C260 source.n90 a_n3654_n2088# 0.014975f
C261 source.n91 a_n3654_n2088# 0.033429f
C262 source.n92 a_n3654_n2088# 0.033429f
C263 source.n93 a_n3654_n2088# 0.014975f
C264 source.n94 a_n3654_n2088# 0.014143f
C265 source.n95 a_n3654_n2088# 0.026319f
C266 source.n96 a_n3654_n2088# 0.026319f
C267 source.n97 a_n3654_n2088# 0.014143f
C268 source.n98 a_n3654_n2088# 0.014975f
C269 source.n99 a_n3654_n2088# 0.033429f
C270 source.n100 a_n3654_n2088# 0.072367f
C271 source.n101 a_n3654_n2088# 0.014975f
C272 source.n102 a_n3654_n2088# 0.014143f
C273 source.n103 a_n3654_n2088# 0.060836f
C274 source.n104 a_n3654_n2088# 0.040492f
C275 source.n105 a_n3654_n2088# 0.144936f
C276 source.t41 a_n3654_n2088# 0.12479f
C277 source.t38 a_n3654_n2088# 0.12479f
C278 source.n106 a_n3654_n2088# 0.971871f
C279 source.n107 a_n3654_n2088# 0.411944f
C280 source.t28 a_n3654_n2088# 0.12479f
C281 source.t30 a_n3654_n2088# 0.12479f
C282 source.n108 a_n3654_n2088# 0.971871f
C283 source.n109 a_n3654_n2088# 0.411944f
C284 source.t36 a_n3654_n2088# 0.12479f
C285 source.t32 a_n3654_n2088# 0.12479f
C286 source.n110 a_n3654_n2088# 0.971871f
C287 source.n111 a_n3654_n2088# 0.411944f
C288 source.t29 a_n3654_n2088# 0.12479f
C289 source.t26 a_n3654_n2088# 0.12479f
C290 source.n112 a_n3654_n2088# 0.971871f
C291 source.n113 a_n3654_n2088# 0.411944f
C292 source.t35 a_n3654_n2088# 0.12479f
C293 source.t44 a_n3654_n2088# 0.12479f
C294 source.n114 a_n3654_n2088# 0.971871f
C295 source.n115 a_n3654_n2088# 0.411944f
C296 source.n116 a_n3654_n2088# 0.036994f
C297 source.n117 a_n3654_n2088# 0.026319f
C298 source.n118 a_n3654_n2088# 0.014143f
C299 source.n119 a_n3654_n2088# 0.033429f
C300 source.n120 a_n3654_n2088# 0.014975f
C301 source.n121 a_n3654_n2088# 0.026319f
C302 source.n122 a_n3654_n2088# 0.014143f
C303 source.n123 a_n3654_n2088# 0.033429f
C304 source.n124 a_n3654_n2088# 0.014975f
C305 source.n125 a_n3654_n2088# 0.112628f
C306 source.t37 a_n3654_n2088# 0.054484f
C307 source.n126 a_n3654_n2088# 0.025071f
C308 source.n127 a_n3654_n2088# 0.019746f
C309 source.n128 a_n3654_n2088# 0.014143f
C310 source.n129 a_n3654_n2088# 0.626241f
C311 source.n130 a_n3654_n2088# 0.026319f
C312 source.n131 a_n3654_n2088# 0.014143f
C313 source.n132 a_n3654_n2088# 0.014975f
C314 source.n133 a_n3654_n2088# 0.033429f
C315 source.n134 a_n3654_n2088# 0.033429f
C316 source.n135 a_n3654_n2088# 0.014975f
C317 source.n136 a_n3654_n2088# 0.014143f
C318 source.n137 a_n3654_n2088# 0.026319f
C319 source.n138 a_n3654_n2088# 0.026319f
C320 source.n139 a_n3654_n2088# 0.014143f
C321 source.n140 a_n3654_n2088# 0.014975f
C322 source.n141 a_n3654_n2088# 0.033429f
C323 source.n142 a_n3654_n2088# 0.072367f
C324 source.n143 a_n3654_n2088# 0.014975f
C325 source.n144 a_n3654_n2088# 0.014143f
C326 source.n145 a_n3654_n2088# 0.060836f
C327 source.n146 a_n3654_n2088# 0.040492f
C328 source.n147 a_n3654_n2088# 1.04945f
C329 source.n148 a_n3654_n2088# 0.036994f
C330 source.n149 a_n3654_n2088# 0.026319f
C331 source.n150 a_n3654_n2088# 0.014143f
C332 source.n151 a_n3654_n2088# 0.033429f
C333 source.n152 a_n3654_n2088# 0.014975f
C334 source.n153 a_n3654_n2088# 0.026319f
C335 source.n154 a_n3654_n2088# 0.014143f
C336 source.n155 a_n3654_n2088# 0.033429f
C337 source.n156 a_n3654_n2088# 0.014975f
C338 source.n157 a_n3654_n2088# 0.112628f
C339 source.t1 a_n3654_n2088# 0.054484f
C340 source.n158 a_n3654_n2088# 0.025071f
C341 source.n159 a_n3654_n2088# 0.019746f
C342 source.n160 a_n3654_n2088# 0.014143f
C343 source.n161 a_n3654_n2088# 0.626241f
C344 source.n162 a_n3654_n2088# 0.026319f
C345 source.n163 a_n3654_n2088# 0.014143f
C346 source.n164 a_n3654_n2088# 0.014975f
C347 source.n165 a_n3654_n2088# 0.033429f
C348 source.n166 a_n3654_n2088# 0.033429f
C349 source.n167 a_n3654_n2088# 0.014975f
C350 source.n168 a_n3654_n2088# 0.014143f
C351 source.n169 a_n3654_n2088# 0.026319f
C352 source.n170 a_n3654_n2088# 0.026319f
C353 source.n171 a_n3654_n2088# 0.014143f
C354 source.n172 a_n3654_n2088# 0.014975f
C355 source.n173 a_n3654_n2088# 0.033429f
C356 source.n174 a_n3654_n2088# 0.072367f
C357 source.n175 a_n3654_n2088# 0.014975f
C358 source.n176 a_n3654_n2088# 0.014143f
C359 source.n177 a_n3654_n2088# 0.060836f
C360 source.n178 a_n3654_n2088# 0.040492f
C361 source.n179 a_n3654_n2088# 1.04945f
C362 source.t17 a_n3654_n2088# 0.12479f
C363 source.t11 a_n3654_n2088# 0.12479f
C364 source.n180 a_n3654_n2088# 0.971864f
C365 source.n181 a_n3654_n2088# 0.411951f
C366 source.t7 a_n3654_n2088# 0.12479f
C367 source.t4 a_n3654_n2088# 0.12479f
C368 source.n182 a_n3654_n2088# 0.971864f
C369 source.n183 a_n3654_n2088# 0.411951f
C370 source.t19 a_n3654_n2088# 0.12479f
C371 source.t18 a_n3654_n2088# 0.12479f
C372 source.n184 a_n3654_n2088# 0.971864f
C373 source.n185 a_n3654_n2088# 0.411951f
C374 source.t0 a_n3654_n2088# 0.12479f
C375 source.t22 a_n3654_n2088# 0.12479f
C376 source.n186 a_n3654_n2088# 0.971864f
C377 source.n187 a_n3654_n2088# 0.411951f
C378 source.t3 a_n3654_n2088# 0.12479f
C379 source.t8 a_n3654_n2088# 0.12479f
C380 source.n188 a_n3654_n2088# 0.971864f
C381 source.n189 a_n3654_n2088# 0.411951f
C382 source.n190 a_n3654_n2088# 0.036994f
C383 source.n191 a_n3654_n2088# 0.026319f
C384 source.n192 a_n3654_n2088# 0.014143f
C385 source.n193 a_n3654_n2088# 0.033429f
C386 source.n194 a_n3654_n2088# 0.014975f
C387 source.n195 a_n3654_n2088# 0.026319f
C388 source.n196 a_n3654_n2088# 0.014143f
C389 source.n197 a_n3654_n2088# 0.033429f
C390 source.n198 a_n3654_n2088# 0.014975f
C391 source.n199 a_n3654_n2088# 0.112628f
C392 source.t12 a_n3654_n2088# 0.054484f
C393 source.n200 a_n3654_n2088# 0.025071f
C394 source.n201 a_n3654_n2088# 0.019746f
C395 source.n202 a_n3654_n2088# 0.014143f
C396 source.n203 a_n3654_n2088# 0.626241f
C397 source.n204 a_n3654_n2088# 0.026319f
C398 source.n205 a_n3654_n2088# 0.014143f
C399 source.n206 a_n3654_n2088# 0.014975f
C400 source.n207 a_n3654_n2088# 0.033429f
C401 source.n208 a_n3654_n2088# 0.033429f
C402 source.n209 a_n3654_n2088# 0.014975f
C403 source.n210 a_n3654_n2088# 0.014143f
C404 source.n211 a_n3654_n2088# 0.026319f
C405 source.n212 a_n3654_n2088# 0.026319f
C406 source.n213 a_n3654_n2088# 0.014143f
C407 source.n214 a_n3654_n2088# 0.014975f
C408 source.n215 a_n3654_n2088# 0.033429f
C409 source.n216 a_n3654_n2088# 0.072367f
C410 source.n217 a_n3654_n2088# 0.014975f
C411 source.n218 a_n3654_n2088# 0.014143f
C412 source.n219 a_n3654_n2088# 0.060836f
C413 source.n220 a_n3654_n2088# 0.040492f
C414 source.n221 a_n3654_n2088# 0.144936f
C415 source.n222 a_n3654_n2088# 0.036994f
C416 source.n223 a_n3654_n2088# 0.026319f
C417 source.n224 a_n3654_n2088# 0.014143f
C418 source.n225 a_n3654_n2088# 0.033429f
C419 source.n226 a_n3654_n2088# 0.014975f
C420 source.n227 a_n3654_n2088# 0.026319f
C421 source.n228 a_n3654_n2088# 0.014143f
C422 source.n229 a_n3654_n2088# 0.033429f
C423 source.n230 a_n3654_n2088# 0.014975f
C424 source.n231 a_n3654_n2088# 0.112628f
C425 source.t34 a_n3654_n2088# 0.054484f
C426 source.n232 a_n3654_n2088# 0.025071f
C427 source.n233 a_n3654_n2088# 0.019746f
C428 source.n234 a_n3654_n2088# 0.014143f
C429 source.n235 a_n3654_n2088# 0.626241f
C430 source.n236 a_n3654_n2088# 0.026319f
C431 source.n237 a_n3654_n2088# 0.014143f
C432 source.n238 a_n3654_n2088# 0.014975f
C433 source.n239 a_n3654_n2088# 0.033429f
C434 source.n240 a_n3654_n2088# 0.033429f
C435 source.n241 a_n3654_n2088# 0.014975f
C436 source.n242 a_n3654_n2088# 0.014143f
C437 source.n243 a_n3654_n2088# 0.026319f
C438 source.n244 a_n3654_n2088# 0.026319f
C439 source.n245 a_n3654_n2088# 0.014143f
C440 source.n246 a_n3654_n2088# 0.014975f
C441 source.n247 a_n3654_n2088# 0.033429f
C442 source.n248 a_n3654_n2088# 0.072367f
C443 source.n249 a_n3654_n2088# 0.014975f
C444 source.n250 a_n3654_n2088# 0.014143f
C445 source.n251 a_n3654_n2088# 0.060836f
C446 source.n252 a_n3654_n2088# 0.040492f
C447 source.n253 a_n3654_n2088# 0.144936f
C448 source.t46 a_n3654_n2088# 0.12479f
C449 source.t42 a_n3654_n2088# 0.12479f
C450 source.n254 a_n3654_n2088# 0.971864f
C451 source.n255 a_n3654_n2088# 0.411951f
C452 source.t24 a_n3654_n2088# 0.12479f
C453 source.t39 a_n3654_n2088# 0.12479f
C454 source.n256 a_n3654_n2088# 0.971864f
C455 source.n257 a_n3654_n2088# 0.411951f
C456 source.t25 a_n3654_n2088# 0.12479f
C457 source.t45 a_n3654_n2088# 0.12479f
C458 source.n258 a_n3654_n2088# 0.971864f
C459 source.n259 a_n3654_n2088# 0.411951f
C460 source.t31 a_n3654_n2088# 0.12479f
C461 source.t43 a_n3654_n2088# 0.12479f
C462 source.n260 a_n3654_n2088# 0.971864f
C463 source.n261 a_n3654_n2088# 0.411951f
C464 source.t27 a_n3654_n2088# 0.12479f
C465 source.t47 a_n3654_n2088# 0.12479f
C466 source.n262 a_n3654_n2088# 0.971864f
C467 source.n263 a_n3654_n2088# 0.411951f
C468 source.n264 a_n3654_n2088# 0.036994f
C469 source.n265 a_n3654_n2088# 0.026319f
C470 source.n266 a_n3654_n2088# 0.014143f
C471 source.n267 a_n3654_n2088# 0.033429f
C472 source.n268 a_n3654_n2088# 0.014975f
C473 source.n269 a_n3654_n2088# 0.026319f
C474 source.n270 a_n3654_n2088# 0.014143f
C475 source.n271 a_n3654_n2088# 0.033429f
C476 source.n272 a_n3654_n2088# 0.014975f
C477 source.n273 a_n3654_n2088# 0.112628f
C478 source.t40 a_n3654_n2088# 0.054484f
C479 source.n274 a_n3654_n2088# 0.025071f
C480 source.n275 a_n3654_n2088# 0.019746f
C481 source.n276 a_n3654_n2088# 0.014143f
C482 source.n277 a_n3654_n2088# 0.626241f
C483 source.n278 a_n3654_n2088# 0.026319f
C484 source.n279 a_n3654_n2088# 0.014143f
C485 source.n280 a_n3654_n2088# 0.014975f
C486 source.n281 a_n3654_n2088# 0.033429f
C487 source.n282 a_n3654_n2088# 0.033429f
C488 source.n283 a_n3654_n2088# 0.014975f
C489 source.n284 a_n3654_n2088# 0.014143f
C490 source.n285 a_n3654_n2088# 0.026319f
C491 source.n286 a_n3654_n2088# 0.026319f
C492 source.n287 a_n3654_n2088# 0.014143f
C493 source.n288 a_n3654_n2088# 0.014975f
C494 source.n289 a_n3654_n2088# 0.033429f
C495 source.n290 a_n3654_n2088# 0.072367f
C496 source.n291 a_n3654_n2088# 0.014975f
C497 source.n292 a_n3654_n2088# 0.014143f
C498 source.n293 a_n3654_n2088# 0.060836f
C499 source.n294 a_n3654_n2088# 0.040492f
C500 source.n295 a_n3654_n2088# 0.322315f
C501 source.n296 a_n3654_n2088# 1.09526f
C502 drain_right.t6 a_n3654_n2088# 0.135579f
C503 drain_right.t5 a_n3654_n2088# 0.135579f
C504 drain_right.n0 a_n3654_n2088# 1.13677f
C505 drain_right.t3 a_n3654_n2088# 0.135579f
C506 drain_right.t18 a_n3654_n2088# 0.135579f
C507 drain_right.n1 a_n3654_n2088# 1.13073f
C508 drain_right.n2 a_n3654_n2088# 0.828664f
C509 drain_right.t20 a_n3654_n2088# 0.135579f
C510 drain_right.t21 a_n3654_n2088# 0.135579f
C511 drain_right.n3 a_n3654_n2088# 1.13073f
C512 drain_right.n4 a_n3654_n2088# 0.363155f
C513 drain_right.t16 a_n3654_n2088# 0.135579f
C514 drain_right.t22 a_n3654_n2088# 0.135579f
C515 drain_right.n5 a_n3654_n2088# 1.13677f
C516 drain_right.t2 a_n3654_n2088# 0.135579f
C517 drain_right.t15 a_n3654_n2088# 0.135579f
C518 drain_right.n6 a_n3654_n2088# 1.13073f
C519 drain_right.n7 a_n3654_n2088# 0.828663f
C520 drain_right.t1 a_n3654_n2088# 0.135579f
C521 drain_right.t17 a_n3654_n2088# 0.135579f
C522 drain_right.n8 a_n3654_n2088# 1.13073f
C523 drain_right.n9 a_n3654_n2088# 0.363155f
C524 drain_right.n10 a_n3654_n2088# 1.53285f
C525 drain_right.t19 a_n3654_n2088# 0.135579f
C526 drain_right.t8 a_n3654_n2088# 0.135579f
C527 drain_right.n11 a_n3654_n2088# 1.13677f
C528 drain_right.t7 a_n3654_n2088# 0.135579f
C529 drain_right.t14 a_n3654_n2088# 0.135579f
C530 drain_right.n12 a_n3654_n2088# 1.13073f
C531 drain_right.n13 a_n3654_n2088# 0.828658f
C532 drain_right.t10 a_n3654_n2088# 0.135579f
C533 drain_right.t4 a_n3654_n2088# 0.135579f
C534 drain_right.n14 a_n3654_n2088# 1.13073f
C535 drain_right.n15 a_n3654_n2088# 0.411591f
C536 drain_right.t11 a_n3654_n2088# 0.135579f
C537 drain_right.t13 a_n3654_n2088# 0.135579f
C538 drain_right.n16 a_n3654_n2088# 1.13073f
C539 drain_right.n17 a_n3654_n2088# 0.411591f
C540 drain_right.t0 a_n3654_n2088# 0.135579f
C541 drain_right.t9 a_n3654_n2088# 0.135579f
C542 drain_right.n18 a_n3654_n2088# 1.13073f
C543 drain_right.n19 a_n3654_n2088# 0.411591f
C544 drain_right.t12 a_n3654_n2088# 0.135579f
C545 drain_right.t23 a_n3654_n2088# 0.135579f
C546 drain_right.n20 a_n3654_n2088# 1.13073f
C547 drain_right.n21 a_n3654_n2088# 0.667998f
C548 minus.n0 a_n3654_n2088# 0.050692f
C549 minus.t3 a_n3654_n2088# 0.528907f
C550 minus.n1 a_n3654_n2088# 0.252009f
C551 minus.t12 a_n3654_n2088# 0.528907f
C552 minus.n2 a_n3654_n2088# 0.037989f
C553 minus.t21 a_n3654_n2088# 0.528907f
C554 minus.n3 a_n3654_n2088# 0.240929f
C555 minus.n4 a_n3654_n2088# 0.063275f
C556 minus.n5 a_n3654_n2088# 0.00862f
C557 minus.t15 a_n3654_n2088# 0.528907f
C558 minus.n6 a_n3654_n2088# 0.037989f
C559 minus.n7 a_n3654_n2088# 0.00862f
C560 minus.t17 a_n3654_n2088# 0.528907f
C561 minus.t14 a_n3654_n2088# 0.549733f
C562 minus.n8 a_n3654_n2088# 0.226917f
C563 minus.t9 a_n3654_n2088# 0.528907f
C564 minus.n9 a_n3654_n2088# 0.251989f
C565 minus.t6 a_n3654_n2088# 0.528907f
C566 minus.n10 a_n3654_n2088# 0.252009f
C567 minus.n11 a_n3654_n2088# 0.218346f
C568 minus.n12 a_n3654_n2088# 0.050692f
C569 minus.n13 a_n3654_n2088# 0.037989f
C570 minus.n14 a_n3654_n2088# 0.240929f
C571 minus.n15 a_n3654_n2088# 0.00862f
C572 minus.t19 a_n3654_n2088# 0.528907f
C573 minus.n16 a_n3654_n2088# 0.240929f
C574 minus.n17 a_n3654_n2088# 0.037989f
C575 minus.n18 a_n3654_n2088# 0.050692f
C576 minus.n19 a_n3654_n2088# 0.063275f
C577 minus.n20 a_n3654_n2088# 0.251541f
C578 minus.t11 a_n3654_n2088# 0.528907f
C579 minus.n21 a_n3654_n2088# 0.251541f
C580 minus.n22 a_n3654_n2088# 0.00862f
C581 minus.n23 a_n3654_n2088# 0.050692f
C582 minus.n24 a_n3654_n2088# 0.037989f
C583 minus.n25 a_n3654_n2088# 0.037989f
C584 minus.n26 a_n3654_n2088# 0.00862f
C585 minus.t18 a_n3654_n2088# 0.528907f
C586 minus.n27 a_n3654_n2088# 0.240929f
C587 minus.n28 a_n3654_n2088# 0.00862f
C588 minus.n29 a_n3654_n2088# 0.050692f
C589 minus.n30 a_n3654_n2088# 0.063275f
C590 minus.n31 a_n3654_n2088# 0.063275f
C591 minus.n32 a_n3654_n2088# 0.251072f
C592 minus.n33 a_n3654_n2088# 0.00862f
C593 minus.t10 a_n3654_n2088# 0.528907f
C594 minus.n34 a_n3654_n2088# 0.237767f
C595 minus.n35 a_n3654_n2088# 1.4857f
C596 minus.n36 a_n3654_n2088# 0.050692f
C597 minus.t20 a_n3654_n2088# 0.528907f
C598 minus.n37 a_n3654_n2088# 0.252009f
C599 minus.n38 a_n3654_n2088# 0.037989f
C600 minus.t16 a_n3654_n2088# 0.528907f
C601 minus.n39 a_n3654_n2088# 0.240929f
C602 minus.n40 a_n3654_n2088# 0.063275f
C603 minus.n41 a_n3654_n2088# 0.00862f
C604 minus.n42 a_n3654_n2088# 0.037989f
C605 minus.n43 a_n3654_n2088# 0.00862f
C606 minus.t13 a_n3654_n2088# 0.549733f
C607 minus.n44 a_n3654_n2088# 0.226917f
C608 minus.t1 a_n3654_n2088# 0.528907f
C609 minus.n45 a_n3654_n2088# 0.251989f
C610 minus.t5 a_n3654_n2088# 0.528907f
C611 minus.n46 a_n3654_n2088# 0.252009f
C612 minus.n47 a_n3654_n2088# 0.218346f
C613 minus.n48 a_n3654_n2088# 0.050692f
C614 minus.n49 a_n3654_n2088# 0.037989f
C615 minus.t23 a_n3654_n2088# 0.528907f
C616 minus.n50 a_n3654_n2088# 0.240929f
C617 minus.n51 a_n3654_n2088# 0.00862f
C618 minus.t8 a_n3654_n2088# 0.528907f
C619 minus.n52 a_n3654_n2088# 0.240929f
C620 minus.n53 a_n3654_n2088# 0.037989f
C621 minus.n54 a_n3654_n2088# 0.050692f
C622 minus.n55 a_n3654_n2088# 0.063275f
C623 minus.t22 a_n3654_n2088# 0.528907f
C624 minus.n56 a_n3654_n2088# 0.251541f
C625 minus.t2 a_n3654_n2088# 0.528907f
C626 minus.n57 a_n3654_n2088# 0.251541f
C627 minus.n58 a_n3654_n2088# 0.00862f
C628 minus.n59 a_n3654_n2088# 0.050692f
C629 minus.n60 a_n3654_n2088# 0.037989f
C630 minus.n61 a_n3654_n2088# 0.037989f
C631 minus.n62 a_n3654_n2088# 0.00862f
C632 minus.t4 a_n3654_n2088# 0.528907f
C633 minus.n63 a_n3654_n2088# 0.240929f
C634 minus.n64 a_n3654_n2088# 0.00862f
C635 minus.n65 a_n3654_n2088# 0.050692f
C636 minus.n66 a_n3654_n2088# 0.063275f
C637 minus.n67 a_n3654_n2088# 0.063275f
C638 minus.t0 a_n3654_n2088# 0.528907f
C639 minus.n68 a_n3654_n2088# 0.251072f
C640 minus.n69 a_n3654_n2088# 0.00862f
C641 minus.t7 a_n3654_n2088# 0.528907f
C642 minus.n70 a_n3654_n2088# 0.237767f
C643 minus.n71 a_n3654_n2088# 0.262539f
C644 minus.n72 a_n3654_n2088# 1.7879f
.ends

