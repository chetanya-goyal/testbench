* NGSPICE file created from diffpair474.ext - technology: sky130A

.subckt diffpair474 minus drain_right drain_left source plus
X0 a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X1 source.t19 minus.t0 drain_right.t3 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X2 source.t0 plus.t0 drain_left.t9 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X3 a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X4 a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X5 source.t6 plus.t1 drain_left.t8 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X6 source.t18 minus.t1 drain_right.t2 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X7 drain_right.t7 minus.t2 source.t17 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X8 source.t16 minus.t3 drain_right.t8 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X9 drain_right.t0 minus.t4 source.t15 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X10 drain_left.t7 plus.t2 source.t9 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X11 source.t14 minus.t5 drain_right.t9 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X12 drain_left.t6 plus.t3 source.t4 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X13 drain_right.t1 minus.t6 source.t13 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X14 drain_right.t5 minus.t7 source.t12 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X15 source.t8 plus.t4 drain_left.t5 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X16 drain_left.t4 plus.t5 source.t5 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X17 drain_left.t3 plus.t6 source.t7 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X18 drain_left.t2 plus.t7 source.t1 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X19 source.t3 plus.t8 drain_left.t1 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X20 a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X21 drain_right.t6 minus.t8 source.t11 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X22 drain_left.t0 plus.t9 source.t2 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X23 drain_right.t4 minus.t9 source.t10 a_n2072_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
R0 minus.n3 minus.t4 433.8
R1 minus.n13 minus.t9 433.8
R2 minus.n2 minus.t3 410.604
R3 minus.n1 minus.t2 410.604
R4 minus.n6 minus.t5 410.604
R5 minus.n8 minus.t6 410.604
R6 minus.n12 minus.t1 410.604
R7 minus.n11 minus.t7 410.604
R8 minus.n16 minus.t0 410.604
R9 minus.n18 minus.t8 410.604
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n19 minus.n18 161.3
R13 minus.n17 minus.n10 161.3
R14 minus.n6 minus.n5 80.6037
R15 minus.n4 minus.n1 80.6037
R16 minus.n16 minus.n15 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n20 minus.n9 37.1463
R23 minus.n7 minus.n6 32.1338
R24 minus.n17 minus.n16 32.1338
R25 minus.n4 minus.n3 31.8629
R26 minus.n14 minus.n13 31.8629
R27 minus.n3 minus.n2 16.2333
R28 minus.n13 minus.n12 16.2333
R29 minus.n8 minus.n7 16.0672
R30 minus.n18 minus.n17 16.0672
R31 minus.n20 minus.n19 6.67664
R32 minus.n5 minus.n4 0.380177
R33 minus.n15 minus.n14 0.380177
R34 minus.n5 minus.n0 0.285035
R35 minus.n15 minus.n10 0.285035
R36 minus.n9 minus.n0 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 drain_right.n60 drain_right.n0 289.615
R40 drain_right.n132 drain_right.n72 289.615
R41 drain_right.n20 drain_right.n19 185
R42 drain_right.n25 drain_right.n24 185
R43 drain_right.n27 drain_right.n26 185
R44 drain_right.n16 drain_right.n15 185
R45 drain_right.n33 drain_right.n32 185
R46 drain_right.n35 drain_right.n34 185
R47 drain_right.n12 drain_right.n11 185
R48 drain_right.n42 drain_right.n41 185
R49 drain_right.n43 drain_right.n10 185
R50 drain_right.n45 drain_right.n44 185
R51 drain_right.n8 drain_right.n7 185
R52 drain_right.n51 drain_right.n50 185
R53 drain_right.n53 drain_right.n52 185
R54 drain_right.n4 drain_right.n3 185
R55 drain_right.n59 drain_right.n58 185
R56 drain_right.n61 drain_right.n60 185
R57 drain_right.n133 drain_right.n132 185
R58 drain_right.n131 drain_right.n130 185
R59 drain_right.n76 drain_right.n75 185
R60 drain_right.n125 drain_right.n124 185
R61 drain_right.n123 drain_right.n122 185
R62 drain_right.n80 drain_right.n79 185
R63 drain_right.n117 drain_right.n116 185
R64 drain_right.n115 drain_right.n82 185
R65 drain_right.n114 drain_right.n113 185
R66 drain_right.n85 drain_right.n83 185
R67 drain_right.n108 drain_right.n107 185
R68 drain_right.n106 drain_right.n105 185
R69 drain_right.n89 drain_right.n88 185
R70 drain_right.n100 drain_right.n99 185
R71 drain_right.n98 drain_right.n97 185
R72 drain_right.n93 drain_right.n92 185
R73 drain_right.n21 drain_right.t4 149.524
R74 drain_right.n94 drain_right.t1 149.524
R75 drain_right.n25 drain_right.n19 104.615
R76 drain_right.n26 drain_right.n25 104.615
R77 drain_right.n26 drain_right.n15 104.615
R78 drain_right.n33 drain_right.n15 104.615
R79 drain_right.n34 drain_right.n33 104.615
R80 drain_right.n34 drain_right.n11 104.615
R81 drain_right.n42 drain_right.n11 104.615
R82 drain_right.n43 drain_right.n42 104.615
R83 drain_right.n44 drain_right.n43 104.615
R84 drain_right.n44 drain_right.n7 104.615
R85 drain_right.n51 drain_right.n7 104.615
R86 drain_right.n52 drain_right.n51 104.615
R87 drain_right.n52 drain_right.n3 104.615
R88 drain_right.n59 drain_right.n3 104.615
R89 drain_right.n60 drain_right.n59 104.615
R90 drain_right.n132 drain_right.n131 104.615
R91 drain_right.n131 drain_right.n75 104.615
R92 drain_right.n124 drain_right.n75 104.615
R93 drain_right.n124 drain_right.n123 104.615
R94 drain_right.n123 drain_right.n79 104.615
R95 drain_right.n116 drain_right.n79 104.615
R96 drain_right.n116 drain_right.n115 104.615
R97 drain_right.n115 drain_right.n114 104.615
R98 drain_right.n114 drain_right.n83 104.615
R99 drain_right.n107 drain_right.n83 104.615
R100 drain_right.n107 drain_right.n106 104.615
R101 drain_right.n106 drain_right.n88 104.615
R102 drain_right.n99 drain_right.n88 104.615
R103 drain_right.n99 drain_right.n98 104.615
R104 drain_right.n98 drain_right.n92 104.615
R105 drain_right.n71 drain_right.n69 60.5266
R106 drain_right.n68 drain_right.n67 60.2278
R107 drain_right.n71 drain_right.n70 59.5527
R108 drain_right.n66 drain_right.n65 59.5525
R109 drain_right.t4 drain_right.n19 52.3082
R110 drain_right.t1 drain_right.n92 52.3082
R111 drain_right.n66 drain_right.n64 47.511
R112 drain_right.n137 drain_right.n136 46.5369
R113 drain_right drain_right.n68 30.9539
R114 drain_right.n45 drain_right.n10 13.1884
R115 drain_right.n117 drain_right.n82 13.1884
R116 drain_right.n41 drain_right.n40 12.8005
R117 drain_right.n46 drain_right.n8 12.8005
R118 drain_right.n118 drain_right.n80 12.8005
R119 drain_right.n113 drain_right.n84 12.8005
R120 drain_right.n39 drain_right.n12 12.0247
R121 drain_right.n50 drain_right.n49 12.0247
R122 drain_right.n122 drain_right.n121 12.0247
R123 drain_right.n112 drain_right.n85 12.0247
R124 drain_right.n36 drain_right.n35 11.249
R125 drain_right.n53 drain_right.n6 11.249
R126 drain_right.n125 drain_right.n78 11.249
R127 drain_right.n109 drain_right.n108 11.249
R128 drain_right.n32 drain_right.n14 10.4732
R129 drain_right.n54 drain_right.n4 10.4732
R130 drain_right.n126 drain_right.n76 10.4732
R131 drain_right.n105 drain_right.n87 10.4732
R132 drain_right.n21 drain_right.n20 10.2747
R133 drain_right.n94 drain_right.n93 10.2747
R134 drain_right.n31 drain_right.n16 9.69747
R135 drain_right.n58 drain_right.n57 9.69747
R136 drain_right.n130 drain_right.n129 9.69747
R137 drain_right.n104 drain_right.n89 9.69747
R138 drain_right.n64 drain_right.n63 9.45567
R139 drain_right.n136 drain_right.n135 9.45567
R140 drain_right.n63 drain_right.n62 9.3005
R141 drain_right.n2 drain_right.n1 9.3005
R142 drain_right.n57 drain_right.n56 9.3005
R143 drain_right.n55 drain_right.n54 9.3005
R144 drain_right.n6 drain_right.n5 9.3005
R145 drain_right.n49 drain_right.n48 9.3005
R146 drain_right.n47 drain_right.n46 9.3005
R147 drain_right.n23 drain_right.n22 9.3005
R148 drain_right.n18 drain_right.n17 9.3005
R149 drain_right.n29 drain_right.n28 9.3005
R150 drain_right.n31 drain_right.n30 9.3005
R151 drain_right.n14 drain_right.n13 9.3005
R152 drain_right.n37 drain_right.n36 9.3005
R153 drain_right.n39 drain_right.n38 9.3005
R154 drain_right.n40 drain_right.n9 9.3005
R155 drain_right.n96 drain_right.n95 9.3005
R156 drain_right.n91 drain_right.n90 9.3005
R157 drain_right.n102 drain_right.n101 9.3005
R158 drain_right.n104 drain_right.n103 9.3005
R159 drain_right.n87 drain_right.n86 9.3005
R160 drain_right.n110 drain_right.n109 9.3005
R161 drain_right.n112 drain_right.n111 9.3005
R162 drain_right.n84 drain_right.n81 9.3005
R163 drain_right.n135 drain_right.n134 9.3005
R164 drain_right.n74 drain_right.n73 9.3005
R165 drain_right.n129 drain_right.n128 9.3005
R166 drain_right.n127 drain_right.n126 9.3005
R167 drain_right.n78 drain_right.n77 9.3005
R168 drain_right.n121 drain_right.n120 9.3005
R169 drain_right.n119 drain_right.n118 9.3005
R170 drain_right.n28 drain_right.n27 8.92171
R171 drain_right.n61 drain_right.n2 8.92171
R172 drain_right.n133 drain_right.n74 8.92171
R173 drain_right.n101 drain_right.n100 8.92171
R174 drain_right.n24 drain_right.n18 8.14595
R175 drain_right.n62 drain_right.n0 8.14595
R176 drain_right.n134 drain_right.n72 8.14595
R177 drain_right.n97 drain_right.n91 8.14595
R178 drain_right.n23 drain_right.n20 7.3702
R179 drain_right.n96 drain_right.n93 7.3702
R180 drain_right drain_right.n137 6.14028
R181 drain_right.n24 drain_right.n23 5.81868
R182 drain_right.n64 drain_right.n0 5.81868
R183 drain_right.n136 drain_right.n72 5.81868
R184 drain_right.n97 drain_right.n96 5.81868
R185 drain_right.n27 drain_right.n18 5.04292
R186 drain_right.n62 drain_right.n61 5.04292
R187 drain_right.n134 drain_right.n133 5.04292
R188 drain_right.n100 drain_right.n91 5.04292
R189 drain_right.n28 drain_right.n16 4.26717
R190 drain_right.n58 drain_right.n2 4.26717
R191 drain_right.n130 drain_right.n74 4.26717
R192 drain_right.n101 drain_right.n89 4.26717
R193 drain_right.n32 drain_right.n31 3.49141
R194 drain_right.n57 drain_right.n4 3.49141
R195 drain_right.n129 drain_right.n76 3.49141
R196 drain_right.n105 drain_right.n104 3.49141
R197 drain_right.n22 drain_right.n21 2.84303
R198 drain_right.n95 drain_right.n94 2.84303
R199 drain_right.n35 drain_right.n14 2.71565
R200 drain_right.n54 drain_right.n53 2.71565
R201 drain_right.n126 drain_right.n125 2.71565
R202 drain_right.n108 drain_right.n87 2.71565
R203 drain_right.n36 drain_right.n12 1.93989
R204 drain_right.n50 drain_right.n6 1.93989
R205 drain_right.n122 drain_right.n78 1.93989
R206 drain_right.n109 drain_right.n85 1.93989
R207 drain_right.n67 drain_right.t3 1.6505
R208 drain_right.n67 drain_right.t6 1.6505
R209 drain_right.n65 drain_right.t2 1.6505
R210 drain_right.n65 drain_right.t5 1.6505
R211 drain_right.n69 drain_right.t8 1.6505
R212 drain_right.n69 drain_right.t0 1.6505
R213 drain_right.n70 drain_right.t9 1.6505
R214 drain_right.n70 drain_right.t7 1.6505
R215 drain_right.n41 drain_right.n39 1.16414
R216 drain_right.n49 drain_right.n8 1.16414
R217 drain_right.n121 drain_right.n80 1.16414
R218 drain_right.n113 drain_right.n112 1.16414
R219 drain_right.n137 drain_right.n71 0.974638
R220 drain_right.n40 drain_right.n10 0.388379
R221 drain_right.n46 drain_right.n45 0.388379
R222 drain_right.n118 drain_right.n117 0.388379
R223 drain_right.n84 drain_right.n82 0.388379
R224 drain_right.n68 drain_right.n66 0.188688
R225 drain_right.n22 drain_right.n17 0.155672
R226 drain_right.n29 drain_right.n17 0.155672
R227 drain_right.n30 drain_right.n29 0.155672
R228 drain_right.n30 drain_right.n13 0.155672
R229 drain_right.n37 drain_right.n13 0.155672
R230 drain_right.n38 drain_right.n37 0.155672
R231 drain_right.n38 drain_right.n9 0.155672
R232 drain_right.n47 drain_right.n9 0.155672
R233 drain_right.n48 drain_right.n47 0.155672
R234 drain_right.n48 drain_right.n5 0.155672
R235 drain_right.n55 drain_right.n5 0.155672
R236 drain_right.n56 drain_right.n55 0.155672
R237 drain_right.n56 drain_right.n1 0.155672
R238 drain_right.n63 drain_right.n1 0.155672
R239 drain_right.n135 drain_right.n73 0.155672
R240 drain_right.n128 drain_right.n73 0.155672
R241 drain_right.n128 drain_right.n127 0.155672
R242 drain_right.n127 drain_right.n77 0.155672
R243 drain_right.n120 drain_right.n77 0.155672
R244 drain_right.n120 drain_right.n119 0.155672
R245 drain_right.n119 drain_right.n81 0.155672
R246 drain_right.n111 drain_right.n81 0.155672
R247 drain_right.n111 drain_right.n110 0.155672
R248 drain_right.n110 drain_right.n86 0.155672
R249 drain_right.n103 drain_right.n86 0.155672
R250 drain_right.n103 drain_right.n102 0.155672
R251 drain_right.n102 drain_right.n90 0.155672
R252 drain_right.n95 drain_right.n90 0.155672
R253 source.n274 source.n214 289.615
R254 source.n204 source.n144 289.615
R255 source.n60 source.n0 289.615
R256 source.n130 source.n70 289.615
R257 source.n234 source.n233 185
R258 source.n239 source.n238 185
R259 source.n241 source.n240 185
R260 source.n230 source.n229 185
R261 source.n247 source.n246 185
R262 source.n249 source.n248 185
R263 source.n226 source.n225 185
R264 source.n256 source.n255 185
R265 source.n257 source.n224 185
R266 source.n259 source.n258 185
R267 source.n222 source.n221 185
R268 source.n265 source.n264 185
R269 source.n267 source.n266 185
R270 source.n218 source.n217 185
R271 source.n273 source.n272 185
R272 source.n275 source.n274 185
R273 source.n164 source.n163 185
R274 source.n169 source.n168 185
R275 source.n171 source.n170 185
R276 source.n160 source.n159 185
R277 source.n177 source.n176 185
R278 source.n179 source.n178 185
R279 source.n156 source.n155 185
R280 source.n186 source.n185 185
R281 source.n187 source.n154 185
R282 source.n189 source.n188 185
R283 source.n152 source.n151 185
R284 source.n195 source.n194 185
R285 source.n197 source.n196 185
R286 source.n148 source.n147 185
R287 source.n203 source.n202 185
R288 source.n205 source.n204 185
R289 source.n61 source.n60 185
R290 source.n59 source.n58 185
R291 source.n4 source.n3 185
R292 source.n53 source.n52 185
R293 source.n51 source.n50 185
R294 source.n8 source.n7 185
R295 source.n45 source.n44 185
R296 source.n43 source.n10 185
R297 source.n42 source.n41 185
R298 source.n13 source.n11 185
R299 source.n36 source.n35 185
R300 source.n34 source.n33 185
R301 source.n17 source.n16 185
R302 source.n28 source.n27 185
R303 source.n26 source.n25 185
R304 source.n21 source.n20 185
R305 source.n131 source.n130 185
R306 source.n129 source.n128 185
R307 source.n74 source.n73 185
R308 source.n123 source.n122 185
R309 source.n121 source.n120 185
R310 source.n78 source.n77 185
R311 source.n115 source.n114 185
R312 source.n113 source.n80 185
R313 source.n112 source.n111 185
R314 source.n83 source.n81 185
R315 source.n106 source.n105 185
R316 source.n104 source.n103 185
R317 source.n87 source.n86 185
R318 source.n98 source.n97 185
R319 source.n96 source.n95 185
R320 source.n91 source.n90 185
R321 source.n235 source.t11 149.524
R322 source.n165 source.t7 149.524
R323 source.n22 source.t1 149.524
R324 source.n92 source.t15 149.524
R325 source.n239 source.n233 104.615
R326 source.n240 source.n239 104.615
R327 source.n240 source.n229 104.615
R328 source.n247 source.n229 104.615
R329 source.n248 source.n247 104.615
R330 source.n248 source.n225 104.615
R331 source.n256 source.n225 104.615
R332 source.n257 source.n256 104.615
R333 source.n258 source.n257 104.615
R334 source.n258 source.n221 104.615
R335 source.n265 source.n221 104.615
R336 source.n266 source.n265 104.615
R337 source.n266 source.n217 104.615
R338 source.n273 source.n217 104.615
R339 source.n274 source.n273 104.615
R340 source.n169 source.n163 104.615
R341 source.n170 source.n169 104.615
R342 source.n170 source.n159 104.615
R343 source.n177 source.n159 104.615
R344 source.n178 source.n177 104.615
R345 source.n178 source.n155 104.615
R346 source.n186 source.n155 104.615
R347 source.n187 source.n186 104.615
R348 source.n188 source.n187 104.615
R349 source.n188 source.n151 104.615
R350 source.n195 source.n151 104.615
R351 source.n196 source.n195 104.615
R352 source.n196 source.n147 104.615
R353 source.n203 source.n147 104.615
R354 source.n204 source.n203 104.615
R355 source.n60 source.n59 104.615
R356 source.n59 source.n3 104.615
R357 source.n52 source.n3 104.615
R358 source.n52 source.n51 104.615
R359 source.n51 source.n7 104.615
R360 source.n44 source.n7 104.615
R361 source.n44 source.n43 104.615
R362 source.n43 source.n42 104.615
R363 source.n42 source.n11 104.615
R364 source.n35 source.n11 104.615
R365 source.n35 source.n34 104.615
R366 source.n34 source.n16 104.615
R367 source.n27 source.n16 104.615
R368 source.n27 source.n26 104.615
R369 source.n26 source.n20 104.615
R370 source.n130 source.n129 104.615
R371 source.n129 source.n73 104.615
R372 source.n122 source.n73 104.615
R373 source.n122 source.n121 104.615
R374 source.n121 source.n77 104.615
R375 source.n114 source.n77 104.615
R376 source.n114 source.n113 104.615
R377 source.n113 source.n112 104.615
R378 source.n112 source.n81 104.615
R379 source.n105 source.n81 104.615
R380 source.n105 source.n104 104.615
R381 source.n104 source.n86 104.615
R382 source.n97 source.n86 104.615
R383 source.n97 source.n96 104.615
R384 source.n96 source.n90 104.615
R385 source.t11 source.n233 52.3082
R386 source.t7 source.n163 52.3082
R387 source.t1 source.n20 52.3082
R388 source.t15 source.n90 52.3082
R389 source.n67 source.n66 42.8739
R390 source.n69 source.n68 42.8739
R391 source.n137 source.n136 42.8739
R392 source.n139 source.n138 42.8739
R393 source.n213 source.n212 42.8737
R394 source.n211 source.n210 42.8737
R395 source.n143 source.n142 42.8737
R396 source.n141 source.n140 42.8737
R397 source.n279 source.n278 29.8581
R398 source.n209 source.n208 29.8581
R399 source.n65 source.n64 29.8581
R400 source.n135 source.n134 29.8581
R401 source.n141 source.n139 23.236
R402 source.n280 source.n65 16.5119
R403 source.n259 source.n224 13.1884
R404 source.n189 source.n154 13.1884
R405 source.n45 source.n10 13.1884
R406 source.n115 source.n80 13.1884
R407 source.n255 source.n254 12.8005
R408 source.n260 source.n222 12.8005
R409 source.n185 source.n184 12.8005
R410 source.n190 source.n152 12.8005
R411 source.n46 source.n8 12.8005
R412 source.n41 source.n12 12.8005
R413 source.n116 source.n78 12.8005
R414 source.n111 source.n82 12.8005
R415 source.n253 source.n226 12.0247
R416 source.n264 source.n263 12.0247
R417 source.n183 source.n156 12.0247
R418 source.n194 source.n193 12.0247
R419 source.n50 source.n49 12.0247
R420 source.n40 source.n13 12.0247
R421 source.n120 source.n119 12.0247
R422 source.n110 source.n83 12.0247
R423 source.n250 source.n249 11.249
R424 source.n267 source.n220 11.249
R425 source.n180 source.n179 11.249
R426 source.n197 source.n150 11.249
R427 source.n53 source.n6 11.249
R428 source.n37 source.n36 11.249
R429 source.n123 source.n76 11.249
R430 source.n107 source.n106 11.249
R431 source.n246 source.n228 10.4732
R432 source.n268 source.n218 10.4732
R433 source.n176 source.n158 10.4732
R434 source.n198 source.n148 10.4732
R435 source.n54 source.n4 10.4732
R436 source.n33 source.n15 10.4732
R437 source.n124 source.n74 10.4732
R438 source.n103 source.n85 10.4732
R439 source.n235 source.n234 10.2747
R440 source.n165 source.n164 10.2747
R441 source.n22 source.n21 10.2747
R442 source.n92 source.n91 10.2747
R443 source.n245 source.n230 9.69747
R444 source.n272 source.n271 9.69747
R445 source.n175 source.n160 9.69747
R446 source.n202 source.n201 9.69747
R447 source.n58 source.n57 9.69747
R448 source.n32 source.n17 9.69747
R449 source.n128 source.n127 9.69747
R450 source.n102 source.n87 9.69747
R451 source.n278 source.n277 9.45567
R452 source.n208 source.n207 9.45567
R453 source.n64 source.n63 9.45567
R454 source.n134 source.n133 9.45567
R455 source.n277 source.n276 9.3005
R456 source.n216 source.n215 9.3005
R457 source.n271 source.n270 9.3005
R458 source.n269 source.n268 9.3005
R459 source.n220 source.n219 9.3005
R460 source.n263 source.n262 9.3005
R461 source.n261 source.n260 9.3005
R462 source.n237 source.n236 9.3005
R463 source.n232 source.n231 9.3005
R464 source.n243 source.n242 9.3005
R465 source.n245 source.n244 9.3005
R466 source.n228 source.n227 9.3005
R467 source.n251 source.n250 9.3005
R468 source.n253 source.n252 9.3005
R469 source.n254 source.n223 9.3005
R470 source.n207 source.n206 9.3005
R471 source.n146 source.n145 9.3005
R472 source.n201 source.n200 9.3005
R473 source.n199 source.n198 9.3005
R474 source.n150 source.n149 9.3005
R475 source.n193 source.n192 9.3005
R476 source.n191 source.n190 9.3005
R477 source.n167 source.n166 9.3005
R478 source.n162 source.n161 9.3005
R479 source.n173 source.n172 9.3005
R480 source.n175 source.n174 9.3005
R481 source.n158 source.n157 9.3005
R482 source.n181 source.n180 9.3005
R483 source.n183 source.n182 9.3005
R484 source.n184 source.n153 9.3005
R485 source.n24 source.n23 9.3005
R486 source.n19 source.n18 9.3005
R487 source.n30 source.n29 9.3005
R488 source.n32 source.n31 9.3005
R489 source.n15 source.n14 9.3005
R490 source.n38 source.n37 9.3005
R491 source.n40 source.n39 9.3005
R492 source.n12 source.n9 9.3005
R493 source.n63 source.n62 9.3005
R494 source.n2 source.n1 9.3005
R495 source.n57 source.n56 9.3005
R496 source.n55 source.n54 9.3005
R497 source.n6 source.n5 9.3005
R498 source.n49 source.n48 9.3005
R499 source.n47 source.n46 9.3005
R500 source.n94 source.n93 9.3005
R501 source.n89 source.n88 9.3005
R502 source.n100 source.n99 9.3005
R503 source.n102 source.n101 9.3005
R504 source.n85 source.n84 9.3005
R505 source.n108 source.n107 9.3005
R506 source.n110 source.n109 9.3005
R507 source.n82 source.n79 9.3005
R508 source.n133 source.n132 9.3005
R509 source.n72 source.n71 9.3005
R510 source.n127 source.n126 9.3005
R511 source.n125 source.n124 9.3005
R512 source.n76 source.n75 9.3005
R513 source.n119 source.n118 9.3005
R514 source.n117 source.n116 9.3005
R515 source.n242 source.n241 8.92171
R516 source.n275 source.n216 8.92171
R517 source.n172 source.n171 8.92171
R518 source.n205 source.n146 8.92171
R519 source.n61 source.n2 8.92171
R520 source.n29 source.n28 8.92171
R521 source.n131 source.n72 8.92171
R522 source.n99 source.n98 8.92171
R523 source.n238 source.n232 8.14595
R524 source.n276 source.n214 8.14595
R525 source.n168 source.n162 8.14595
R526 source.n206 source.n144 8.14595
R527 source.n62 source.n0 8.14595
R528 source.n25 source.n19 8.14595
R529 source.n132 source.n70 8.14595
R530 source.n95 source.n89 8.14595
R531 source.n237 source.n234 7.3702
R532 source.n167 source.n164 7.3702
R533 source.n24 source.n21 7.3702
R534 source.n94 source.n91 7.3702
R535 source.n238 source.n237 5.81868
R536 source.n278 source.n214 5.81868
R537 source.n168 source.n167 5.81868
R538 source.n208 source.n144 5.81868
R539 source.n64 source.n0 5.81868
R540 source.n25 source.n24 5.81868
R541 source.n134 source.n70 5.81868
R542 source.n95 source.n94 5.81868
R543 source.n280 source.n279 5.7505
R544 source.n241 source.n232 5.04292
R545 source.n276 source.n275 5.04292
R546 source.n171 source.n162 5.04292
R547 source.n206 source.n205 5.04292
R548 source.n62 source.n61 5.04292
R549 source.n28 source.n19 5.04292
R550 source.n132 source.n131 5.04292
R551 source.n98 source.n89 5.04292
R552 source.n242 source.n230 4.26717
R553 source.n272 source.n216 4.26717
R554 source.n172 source.n160 4.26717
R555 source.n202 source.n146 4.26717
R556 source.n58 source.n2 4.26717
R557 source.n29 source.n17 4.26717
R558 source.n128 source.n72 4.26717
R559 source.n99 source.n87 4.26717
R560 source.n246 source.n245 3.49141
R561 source.n271 source.n218 3.49141
R562 source.n176 source.n175 3.49141
R563 source.n201 source.n148 3.49141
R564 source.n57 source.n4 3.49141
R565 source.n33 source.n32 3.49141
R566 source.n127 source.n74 3.49141
R567 source.n103 source.n102 3.49141
R568 source.n236 source.n235 2.84303
R569 source.n166 source.n165 2.84303
R570 source.n23 source.n22 2.84303
R571 source.n93 source.n92 2.84303
R572 source.n249 source.n228 2.71565
R573 source.n268 source.n267 2.71565
R574 source.n179 source.n158 2.71565
R575 source.n198 source.n197 2.71565
R576 source.n54 source.n53 2.71565
R577 source.n36 source.n15 2.71565
R578 source.n124 source.n123 2.71565
R579 source.n106 source.n85 2.71565
R580 source.n250 source.n226 1.93989
R581 source.n264 source.n220 1.93989
R582 source.n180 source.n156 1.93989
R583 source.n194 source.n150 1.93989
R584 source.n50 source.n6 1.93989
R585 source.n37 source.n13 1.93989
R586 source.n120 source.n76 1.93989
R587 source.n107 source.n83 1.93989
R588 source.n212 source.t12 1.6505
R589 source.n212 source.t19 1.6505
R590 source.n210 source.t10 1.6505
R591 source.n210 source.t18 1.6505
R592 source.n142 source.t4 1.6505
R593 source.n142 source.t6 1.6505
R594 source.n140 source.t9 1.6505
R595 source.n140 source.t0 1.6505
R596 source.n66 source.t5 1.6505
R597 source.n66 source.t8 1.6505
R598 source.n68 source.t2 1.6505
R599 source.n68 source.t3 1.6505
R600 source.n136 source.t17 1.6505
R601 source.n136 source.t16 1.6505
R602 source.n138 source.t13 1.6505
R603 source.n138 source.t14 1.6505
R604 source.n255 source.n253 1.16414
R605 source.n263 source.n222 1.16414
R606 source.n185 source.n183 1.16414
R607 source.n193 source.n152 1.16414
R608 source.n49 source.n8 1.16414
R609 source.n41 source.n40 1.16414
R610 source.n119 source.n78 1.16414
R611 source.n111 source.n110 1.16414
R612 source.n139 source.n137 0.974638
R613 source.n137 source.n135 0.974638
R614 source.n69 source.n67 0.974638
R615 source.n67 source.n65 0.974638
R616 source.n143 source.n141 0.974638
R617 source.n209 source.n143 0.974638
R618 source.n213 source.n211 0.974638
R619 source.n279 source.n213 0.974638
R620 source.n135 source.n69 0.957397
R621 source.n211 source.n209 0.957397
R622 source.n254 source.n224 0.388379
R623 source.n260 source.n259 0.388379
R624 source.n184 source.n154 0.388379
R625 source.n190 source.n189 0.388379
R626 source.n46 source.n45 0.388379
R627 source.n12 source.n10 0.388379
R628 source.n116 source.n115 0.388379
R629 source.n82 source.n80 0.388379
R630 source source.n280 0.188
R631 source.n236 source.n231 0.155672
R632 source.n243 source.n231 0.155672
R633 source.n244 source.n243 0.155672
R634 source.n244 source.n227 0.155672
R635 source.n251 source.n227 0.155672
R636 source.n252 source.n251 0.155672
R637 source.n252 source.n223 0.155672
R638 source.n261 source.n223 0.155672
R639 source.n262 source.n261 0.155672
R640 source.n262 source.n219 0.155672
R641 source.n269 source.n219 0.155672
R642 source.n270 source.n269 0.155672
R643 source.n270 source.n215 0.155672
R644 source.n277 source.n215 0.155672
R645 source.n166 source.n161 0.155672
R646 source.n173 source.n161 0.155672
R647 source.n174 source.n173 0.155672
R648 source.n174 source.n157 0.155672
R649 source.n181 source.n157 0.155672
R650 source.n182 source.n181 0.155672
R651 source.n182 source.n153 0.155672
R652 source.n191 source.n153 0.155672
R653 source.n192 source.n191 0.155672
R654 source.n192 source.n149 0.155672
R655 source.n199 source.n149 0.155672
R656 source.n200 source.n199 0.155672
R657 source.n200 source.n145 0.155672
R658 source.n207 source.n145 0.155672
R659 source.n63 source.n1 0.155672
R660 source.n56 source.n1 0.155672
R661 source.n56 source.n55 0.155672
R662 source.n55 source.n5 0.155672
R663 source.n48 source.n5 0.155672
R664 source.n48 source.n47 0.155672
R665 source.n47 source.n9 0.155672
R666 source.n39 source.n9 0.155672
R667 source.n39 source.n38 0.155672
R668 source.n38 source.n14 0.155672
R669 source.n31 source.n14 0.155672
R670 source.n31 source.n30 0.155672
R671 source.n30 source.n18 0.155672
R672 source.n23 source.n18 0.155672
R673 source.n133 source.n71 0.155672
R674 source.n126 source.n71 0.155672
R675 source.n126 source.n125 0.155672
R676 source.n125 source.n75 0.155672
R677 source.n118 source.n75 0.155672
R678 source.n118 source.n117 0.155672
R679 source.n117 source.n79 0.155672
R680 source.n109 source.n79 0.155672
R681 source.n109 source.n108 0.155672
R682 source.n108 source.n84 0.155672
R683 source.n101 source.n84 0.155672
R684 source.n101 source.n100 0.155672
R685 source.n100 source.n88 0.155672
R686 source.n93 source.n88 0.155672
R687 plus.n3 plus.t9 433.8
R688 plus.n13 plus.t6 433.8
R689 plus.n8 plus.t7 410.604
R690 plus.n6 plus.t4 410.604
R691 plus.n5 plus.t5 410.604
R692 plus.n4 plus.t8 410.604
R693 plus.n18 plus.t2 410.604
R694 plus.n16 plus.t0 410.604
R695 plus.n15 plus.t3 410.604
R696 plus.n14 plus.t1 410.604
R697 plus.n7 plus.n0 161.3
R698 plus.n9 plus.n8 161.3
R699 plus.n17 plus.n10 161.3
R700 plus.n19 plus.n18 161.3
R701 plus.n5 plus.n2 80.6037
R702 plus.n6 plus.n1 80.6037
R703 plus.n15 plus.n12 80.6037
R704 plus.n16 plus.n11 80.6037
R705 plus.n6 plus.n5 48.2005
R706 plus.n5 plus.n4 48.2005
R707 plus.n16 plus.n15 48.2005
R708 plus.n15 plus.n14 48.2005
R709 plus.n7 plus.n6 32.1338
R710 plus.n17 plus.n16 32.1338
R711 plus.n3 plus.n2 31.8629
R712 plus.n13 plus.n12 31.8629
R713 plus plus.n19 31.0274
R714 plus.n4 plus.n3 16.2333
R715 plus.n14 plus.n13 16.2333
R716 plus.n8 plus.n7 16.0672
R717 plus.n18 plus.n17 16.0672
R718 plus plus.n9 12.3206
R719 plus.n2 plus.n1 0.380177
R720 plus.n12 plus.n11 0.380177
R721 plus.n1 plus.n0 0.285035
R722 plus.n11 plus.n10 0.285035
R723 plus.n9 plus.n0 0.189894
R724 plus.n19 plus.n10 0.189894
R725 drain_left.n60 drain_left.n0 289.615
R726 drain_left.n129 drain_left.n69 289.615
R727 drain_left.n20 drain_left.n19 185
R728 drain_left.n25 drain_left.n24 185
R729 drain_left.n27 drain_left.n26 185
R730 drain_left.n16 drain_left.n15 185
R731 drain_left.n33 drain_left.n32 185
R732 drain_left.n35 drain_left.n34 185
R733 drain_left.n12 drain_left.n11 185
R734 drain_left.n42 drain_left.n41 185
R735 drain_left.n43 drain_left.n10 185
R736 drain_left.n45 drain_left.n44 185
R737 drain_left.n8 drain_left.n7 185
R738 drain_left.n51 drain_left.n50 185
R739 drain_left.n53 drain_left.n52 185
R740 drain_left.n4 drain_left.n3 185
R741 drain_left.n59 drain_left.n58 185
R742 drain_left.n61 drain_left.n60 185
R743 drain_left.n130 drain_left.n129 185
R744 drain_left.n128 drain_left.n127 185
R745 drain_left.n73 drain_left.n72 185
R746 drain_left.n122 drain_left.n121 185
R747 drain_left.n120 drain_left.n119 185
R748 drain_left.n77 drain_left.n76 185
R749 drain_left.n114 drain_left.n113 185
R750 drain_left.n112 drain_left.n79 185
R751 drain_left.n111 drain_left.n110 185
R752 drain_left.n82 drain_left.n80 185
R753 drain_left.n105 drain_left.n104 185
R754 drain_left.n103 drain_left.n102 185
R755 drain_left.n86 drain_left.n85 185
R756 drain_left.n97 drain_left.n96 185
R757 drain_left.n95 drain_left.n94 185
R758 drain_left.n90 drain_left.n89 185
R759 drain_left.n21 drain_left.t7 149.524
R760 drain_left.n91 drain_left.t0 149.524
R761 drain_left.n25 drain_left.n19 104.615
R762 drain_left.n26 drain_left.n25 104.615
R763 drain_left.n26 drain_left.n15 104.615
R764 drain_left.n33 drain_left.n15 104.615
R765 drain_left.n34 drain_left.n33 104.615
R766 drain_left.n34 drain_left.n11 104.615
R767 drain_left.n42 drain_left.n11 104.615
R768 drain_left.n43 drain_left.n42 104.615
R769 drain_left.n44 drain_left.n43 104.615
R770 drain_left.n44 drain_left.n7 104.615
R771 drain_left.n51 drain_left.n7 104.615
R772 drain_left.n52 drain_left.n51 104.615
R773 drain_left.n52 drain_left.n3 104.615
R774 drain_left.n59 drain_left.n3 104.615
R775 drain_left.n60 drain_left.n59 104.615
R776 drain_left.n129 drain_left.n128 104.615
R777 drain_left.n128 drain_left.n72 104.615
R778 drain_left.n121 drain_left.n72 104.615
R779 drain_left.n121 drain_left.n120 104.615
R780 drain_left.n120 drain_left.n76 104.615
R781 drain_left.n113 drain_left.n76 104.615
R782 drain_left.n113 drain_left.n112 104.615
R783 drain_left.n112 drain_left.n111 104.615
R784 drain_left.n111 drain_left.n80 104.615
R785 drain_left.n104 drain_left.n80 104.615
R786 drain_left.n104 drain_left.n103 104.615
R787 drain_left.n103 drain_left.n85 104.615
R788 drain_left.n96 drain_left.n85 104.615
R789 drain_left.n96 drain_left.n95 104.615
R790 drain_left.n95 drain_left.n89 104.615
R791 drain_left.n68 drain_left.n67 60.2278
R792 drain_left.n135 drain_left.n134 59.5527
R793 drain_left.n66 drain_left.n65 59.5525
R794 drain_left.n137 drain_left.n136 59.5525
R795 drain_left.t7 drain_left.n19 52.3082
R796 drain_left.t0 drain_left.n89 52.3082
R797 drain_left.n66 drain_left.n64 47.511
R798 drain_left.n135 drain_left.n133 47.511
R799 drain_left drain_left.n68 31.5072
R800 drain_left.n45 drain_left.n10 13.1884
R801 drain_left.n114 drain_left.n79 13.1884
R802 drain_left.n41 drain_left.n40 12.8005
R803 drain_left.n46 drain_left.n8 12.8005
R804 drain_left.n115 drain_left.n77 12.8005
R805 drain_left.n110 drain_left.n81 12.8005
R806 drain_left.n39 drain_left.n12 12.0247
R807 drain_left.n50 drain_left.n49 12.0247
R808 drain_left.n119 drain_left.n118 12.0247
R809 drain_left.n109 drain_left.n82 12.0247
R810 drain_left.n36 drain_left.n35 11.249
R811 drain_left.n53 drain_left.n6 11.249
R812 drain_left.n122 drain_left.n75 11.249
R813 drain_left.n106 drain_left.n105 11.249
R814 drain_left.n32 drain_left.n14 10.4732
R815 drain_left.n54 drain_left.n4 10.4732
R816 drain_left.n123 drain_left.n73 10.4732
R817 drain_left.n102 drain_left.n84 10.4732
R818 drain_left.n21 drain_left.n20 10.2747
R819 drain_left.n91 drain_left.n90 10.2747
R820 drain_left.n31 drain_left.n16 9.69747
R821 drain_left.n58 drain_left.n57 9.69747
R822 drain_left.n127 drain_left.n126 9.69747
R823 drain_left.n101 drain_left.n86 9.69747
R824 drain_left.n64 drain_left.n63 9.45567
R825 drain_left.n133 drain_left.n132 9.45567
R826 drain_left.n63 drain_left.n62 9.3005
R827 drain_left.n2 drain_left.n1 9.3005
R828 drain_left.n57 drain_left.n56 9.3005
R829 drain_left.n55 drain_left.n54 9.3005
R830 drain_left.n6 drain_left.n5 9.3005
R831 drain_left.n49 drain_left.n48 9.3005
R832 drain_left.n47 drain_left.n46 9.3005
R833 drain_left.n23 drain_left.n22 9.3005
R834 drain_left.n18 drain_left.n17 9.3005
R835 drain_left.n29 drain_left.n28 9.3005
R836 drain_left.n31 drain_left.n30 9.3005
R837 drain_left.n14 drain_left.n13 9.3005
R838 drain_left.n37 drain_left.n36 9.3005
R839 drain_left.n39 drain_left.n38 9.3005
R840 drain_left.n40 drain_left.n9 9.3005
R841 drain_left.n93 drain_left.n92 9.3005
R842 drain_left.n88 drain_left.n87 9.3005
R843 drain_left.n99 drain_left.n98 9.3005
R844 drain_left.n101 drain_left.n100 9.3005
R845 drain_left.n84 drain_left.n83 9.3005
R846 drain_left.n107 drain_left.n106 9.3005
R847 drain_left.n109 drain_left.n108 9.3005
R848 drain_left.n81 drain_left.n78 9.3005
R849 drain_left.n132 drain_left.n131 9.3005
R850 drain_left.n71 drain_left.n70 9.3005
R851 drain_left.n126 drain_left.n125 9.3005
R852 drain_left.n124 drain_left.n123 9.3005
R853 drain_left.n75 drain_left.n74 9.3005
R854 drain_left.n118 drain_left.n117 9.3005
R855 drain_left.n116 drain_left.n115 9.3005
R856 drain_left.n28 drain_left.n27 8.92171
R857 drain_left.n61 drain_left.n2 8.92171
R858 drain_left.n130 drain_left.n71 8.92171
R859 drain_left.n98 drain_left.n97 8.92171
R860 drain_left.n24 drain_left.n18 8.14595
R861 drain_left.n62 drain_left.n0 8.14595
R862 drain_left.n131 drain_left.n69 8.14595
R863 drain_left.n94 drain_left.n88 8.14595
R864 drain_left.n23 drain_left.n20 7.3702
R865 drain_left.n93 drain_left.n90 7.3702
R866 drain_left drain_left.n137 6.62735
R867 drain_left.n24 drain_left.n23 5.81868
R868 drain_left.n64 drain_left.n0 5.81868
R869 drain_left.n133 drain_left.n69 5.81868
R870 drain_left.n94 drain_left.n93 5.81868
R871 drain_left.n27 drain_left.n18 5.04292
R872 drain_left.n62 drain_left.n61 5.04292
R873 drain_left.n131 drain_left.n130 5.04292
R874 drain_left.n97 drain_left.n88 5.04292
R875 drain_left.n28 drain_left.n16 4.26717
R876 drain_left.n58 drain_left.n2 4.26717
R877 drain_left.n127 drain_left.n71 4.26717
R878 drain_left.n98 drain_left.n86 4.26717
R879 drain_left.n32 drain_left.n31 3.49141
R880 drain_left.n57 drain_left.n4 3.49141
R881 drain_left.n126 drain_left.n73 3.49141
R882 drain_left.n102 drain_left.n101 3.49141
R883 drain_left.n22 drain_left.n21 2.84303
R884 drain_left.n92 drain_left.n91 2.84303
R885 drain_left.n35 drain_left.n14 2.71565
R886 drain_left.n54 drain_left.n53 2.71565
R887 drain_left.n123 drain_left.n122 2.71565
R888 drain_left.n105 drain_left.n84 2.71565
R889 drain_left.n36 drain_left.n12 1.93989
R890 drain_left.n50 drain_left.n6 1.93989
R891 drain_left.n119 drain_left.n75 1.93989
R892 drain_left.n106 drain_left.n82 1.93989
R893 drain_left.n67 drain_left.t8 1.6505
R894 drain_left.n67 drain_left.t3 1.6505
R895 drain_left.n65 drain_left.t9 1.6505
R896 drain_left.n65 drain_left.t6 1.6505
R897 drain_left.n136 drain_left.t5 1.6505
R898 drain_left.n136 drain_left.t2 1.6505
R899 drain_left.n134 drain_left.t1 1.6505
R900 drain_left.n134 drain_left.t4 1.6505
R901 drain_left.n41 drain_left.n39 1.16414
R902 drain_left.n49 drain_left.n8 1.16414
R903 drain_left.n118 drain_left.n77 1.16414
R904 drain_left.n110 drain_left.n109 1.16414
R905 drain_left.n137 drain_left.n135 0.974638
R906 drain_left.n40 drain_left.n10 0.388379
R907 drain_left.n46 drain_left.n45 0.388379
R908 drain_left.n115 drain_left.n114 0.388379
R909 drain_left.n81 drain_left.n79 0.388379
R910 drain_left.n68 drain_left.n66 0.188688
R911 drain_left.n22 drain_left.n17 0.155672
R912 drain_left.n29 drain_left.n17 0.155672
R913 drain_left.n30 drain_left.n29 0.155672
R914 drain_left.n30 drain_left.n13 0.155672
R915 drain_left.n37 drain_left.n13 0.155672
R916 drain_left.n38 drain_left.n37 0.155672
R917 drain_left.n38 drain_left.n9 0.155672
R918 drain_left.n47 drain_left.n9 0.155672
R919 drain_left.n48 drain_left.n47 0.155672
R920 drain_left.n48 drain_left.n5 0.155672
R921 drain_left.n55 drain_left.n5 0.155672
R922 drain_left.n56 drain_left.n55 0.155672
R923 drain_left.n56 drain_left.n1 0.155672
R924 drain_left.n63 drain_left.n1 0.155672
R925 drain_left.n132 drain_left.n70 0.155672
R926 drain_left.n125 drain_left.n70 0.155672
R927 drain_left.n125 drain_left.n124 0.155672
R928 drain_left.n124 drain_left.n74 0.155672
R929 drain_left.n117 drain_left.n74 0.155672
R930 drain_left.n117 drain_left.n116 0.155672
R931 drain_left.n116 drain_left.n78 0.155672
R932 drain_left.n108 drain_left.n78 0.155672
R933 drain_left.n108 drain_left.n107 0.155672
R934 drain_left.n107 drain_left.n83 0.155672
R935 drain_left.n100 drain_left.n83 0.155672
R936 drain_left.n100 drain_left.n99 0.155672
R937 drain_left.n99 drain_left.n87 0.155672
R938 drain_left.n92 drain_left.n87 0.155672
C0 minus source 7.05966f
C1 minus plus 5.72441f
C2 minus drain_left 0.172418f
C3 source plus 7.07417f
C4 drain_left source 13.5812f
C5 minus drain_right 7.17872f
C6 source drain_right 13.575701f
C7 drain_left plus 7.37925f
C8 drain_right plus 0.360171f
C9 drain_left drain_right 1.03391f
C10 drain_right a_n2072_n3288# 7.05052f
C11 drain_left a_n2072_n3288# 7.36373f
C12 source a_n2072_n3288# 6.635383f
C13 minus a_n2072_n3288# 8.116245f
C14 plus a_n2072_n3288# 9.75319f
C15 drain_left.n0 a_n2072_n3288# 0.031747f
C16 drain_left.n1 a_n2072_n3288# 0.023967f
C17 drain_left.n2 a_n2072_n3288# 0.012879f
C18 drain_left.n3 a_n2072_n3288# 0.03044f
C19 drain_left.n4 a_n2072_n3288# 0.013636f
C20 drain_left.n5 a_n2072_n3288# 0.023967f
C21 drain_left.n6 a_n2072_n3288# 0.012879f
C22 drain_left.n7 a_n2072_n3288# 0.03044f
C23 drain_left.n8 a_n2072_n3288# 0.013636f
C24 drain_left.n9 a_n2072_n3288# 0.023967f
C25 drain_left.n10 a_n2072_n3288# 0.013257f
C26 drain_left.n11 a_n2072_n3288# 0.03044f
C27 drain_left.n12 a_n2072_n3288# 0.013636f
C28 drain_left.n13 a_n2072_n3288# 0.023967f
C29 drain_left.n14 a_n2072_n3288# 0.012879f
C30 drain_left.n15 a_n2072_n3288# 0.03044f
C31 drain_left.n16 a_n2072_n3288# 0.013636f
C32 drain_left.n17 a_n2072_n3288# 0.023967f
C33 drain_left.n18 a_n2072_n3288# 0.012879f
C34 drain_left.n19 a_n2072_n3288# 0.02283f
C35 drain_left.n20 a_n2072_n3288# 0.021519f
C36 drain_left.t7 a_n2072_n3288# 0.051412f
C37 drain_left.n21 a_n2072_n3288# 0.172796f
C38 drain_left.n22 a_n2072_n3288# 1.20907f
C39 drain_left.n23 a_n2072_n3288# 0.012879f
C40 drain_left.n24 a_n2072_n3288# 0.013636f
C41 drain_left.n25 a_n2072_n3288# 0.03044f
C42 drain_left.n26 a_n2072_n3288# 0.03044f
C43 drain_left.n27 a_n2072_n3288# 0.013636f
C44 drain_left.n28 a_n2072_n3288# 0.012879f
C45 drain_left.n29 a_n2072_n3288# 0.023967f
C46 drain_left.n30 a_n2072_n3288# 0.023967f
C47 drain_left.n31 a_n2072_n3288# 0.012879f
C48 drain_left.n32 a_n2072_n3288# 0.013636f
C49 drain_left.n33 a_n2072_n3288# 0.03044f
C50 drain_left.n34 a_n2072_n3288# 0.03044f
C51 drain_left.n35 a_n2072_n3288# 0.013636f
C52 drain_left.n36 a_n2072_n3288# 0.012879f
C53 drain_left.n37 a_n2072_n3288# 0.023967f
C54 drain_left.n38 a_n2072_n3288# 0.023967f
C55 drain_left.n39 a_n2072_n3288# 0.012879f
C56 drain_left.n40 a_n2072_n3288# 0.012879f
C57 drain_left.n41 a_n2072_n3288# 0.013636f
C58 drain_left.n42 a_n2072_n3288# 0.03044f
C59 drain_left.n43 a_n2072_n3288# 0.03044f
C60 drain_left.n44 a_n2072_n3288# 0.03044f
C61 drain_left.n45 a_n2072_n3288# 0.013257f
C62 drain_left.n46 a_n2072_n3288# 0.012879f
C63 drain_left.n47 a_n2072_n3288# 0.023967f
C64 drain_left.n48 a_n2072_n3288# 0.023967f
C65 drain_left.n49 a_n2072_n3288# 0.012879f
C66 drain_left.n50 a_n2072_n3288# 0.013636f
C67 drain_left.n51 a_n2072_n3288# 0.03044f
C68 drain_left.n52 a_n2072_n3288# 0.03044f
C69 drain_left.n53 a_n2072_n3288# 0.013636f
C70 drain_left.n54 a_n2072_n3288# 0.012879f
C71 drain_left.n55 a_n2072_n3288# 0.023967f
C72 drain_left.n56 a_n2072_n3288# 0.023967f
C73 drain_left.n57 a_n2072_n3288# 0.012879f
C74 drain_left.n58 a_n2072_n3288# 0.013636f
C75 drain_left.n59 a_n2072_n3288# 0.03044f
C76 drain_left.n60 a_n2072_n3288# 0.062467f
C77 drain_left.n61 a_n2072_n3288# 0.013636f
C78 drain_left.n62 a_n2072_n3288# 0.012879f
C79 drain_left.n63 a_n2072_n3288# 0.051469f
C80 drain_left.n64 a_n2072_n3288# 0.0535f
C81 drain_left.t9 a_n2072_n3288# 0.227269f
C82 drain_left.t6 a_n2072_n3288# 0.227269f
C83 drain_left.n65 a_n2072_n3288# 2.02234f
C84 drain_left.n66 a_n2072_n3288# 0.410542f
C85 drain_left.t8 a_n2072_n3288# 0.227269f
C86 drain_left.t3 a_n2072_n3288# 0.227269f
C87 drain_left.n67 a_n2072_n3288# 2.02614f
C88 drain_left.n68 a_n2072_n3288# 1.59156f
C89 drain_left.n69 a_n2072_n3288# 0.031747f
C90 drain_left.n70 a_n2072_n3288# 0.023967f
C91 drain_left.n71 a_n2072_n3288# 0.012879f
C92 drain_left.n72 a_n2072_n3288# 0.03044f
C93 drain_left.n73 a_n2072_n3288# 0.013636f
C94 drain_left.n74 a_n2072_n3288# 0.023967f
C95 drain_left.n75 a_n2072_n3288# 0.012879f
C96 drain_left.n76 a_n2072_n3288# 0.03044f
C97 drain_left.n77 a_n2072_n3288# 0.013636f
C98 drain_left.n78 a_n2072_n3288# 0.023967f
C99 drain_left.n79 a_n2072_n3288# 0.013257f
C100 drain_left.n80 a_n2072_n3288# 0.03044f
C101 drain_left.n81 a_n2072_n3288# 0.012879f
C102 drain_left.n82 a_n2072_n3288# 0.013636f
C103 drain_left.n83 a_n2072_n3288# 0.023967f
C104 drain_left.n84 a_n2072_n3288# 0.012879f
C105 drain_left.n85 a_n2072_n3288# 0.03044f
C106 drain_left.n86 a_n2072_n3288# 0.013636f
C107 drain_left.n87 a_n2072_n3288# 0.023967f
C108 drain_left.n88 a_n2072_n3288# 0.012879f
C109 drain_left.n89 a_n2072_n3288# 0.02283f
C110 drain_left.n90 a_n2072_n3288# 0.021519f
C111 drain_left.t0 a_n2072_n3288# 0.051412f
C112 drain_left.n91 a_n2072_n3288# 0.172796f
C113 drain_left.n92 a_n2072_n3288# 1.20907f
C114 drain_left.n93 a_n2072_n3288# 0.012879f
C115 drain_left.n94 a_n2072_n3288# 0.013636f
C116 drain_left.n95 a_n2072_n3288# 0.03044f
C117 drain_left.n96 a_n2072_n3288# 0.03044f
C118 drain_left.n97 a_n2072_n3288# 0.013636f
C119 drain_left.n98 a_n2072_n3288# 0.012879f
C120 drain_left.n99 a_n2072_n3288# 0.023967f
C121 drain_left.n100 a_n2072_n3288# 0.023967f
C122 drain_left.n101 a_n2072_n3288# 0.012879f
C123 drain_left.n102 a_n2072_n3288# 0.013636f
C124 drain_left.n103 a_n2072_n3288# 0.03044f
C125 drain_left.n104 a_n2072_n3288# 0.03044f
C126 drain_left.n105 a_n2072_n3288# 0.013636f
C127 drain_left.n106 a_n2072_n3288# 0.012879f
C128 drain_left.n107 a_n2072_n3288# 0.023967f
C129 drain_left.n108 a_n2072_n3288# 0.023967f
C130 drain_left.n109 a_n2072_n3288# 0.012879f
C131 drain_left.n110 a_n2072_n3288# 0.013636f
C132 drain_left.n111 a_n2072_n3288# 0.03044f
C133 drain_left.n112 a_n2072_n3288# 0.03044f
C134 drain_left.n113 a_n2072_n3288# 0.03044f
C135 drain_left.n114 a_n2072_n3288# 0.013257f
C136 drain_left.n115 a_n2072_n3288# 0.012879f
C137 drain_left.n116 a_n2072_n3288# 0.023967f
C138 drain_left.n117 a_n2072_n3288# 0.023967f
C139 drain_left.n118 a_n2072_n3288# 0.012879f
C140 drain_left.n119 a_n2072_n3288# 0.013636f
C141 drain_left.n120 a_n2072_n3288# 0.03044f
C142 drain_left.n121 a_n2072_n3288# 0.03044f
C143 drain_left.n122 a_n2072_n3288# 0.013636f
C144 drain_left.n123 a_n2072_n3288# 0.012879f
C145 drain_left.n124 a_n2072_n3288# 0.023967f
C146 drain_left.n125 a_n2072_n3288# 0.023967f
C147 drain_left.n126 a_n2072_n3288# 0.012879f
C148 drain_left.n127 a_n2072_n3288# 0.013636f
C149 drain_left.n128 a_n2072_n3288# 0.03044f
C150 drain_left.n129 a_n2072_n3288# 0.062467f
C151 drain_left.n130 a_n2072_n3288# 0.013636f
C152 drain_left.n131 a_n2072_n3288# 0.012879f
C153 drain_left.n132 a_n2072_n3288# 0.051469f
C154 drain_left.n133 a_n2072_n3288# 0.0535f
C155 drain_left.t1 a_n2072_n3288# 0.227269f
C156 drain_left.t4 a_n2072_n3288# 0.227269f
C157 drain_left.n134 a_n2072_n3288# 2.02235f
C158 drain_left.n135 a_n2072_n3288# 0.468277f
C159 drain_left.t5 a_n2072_n3288# 0.227269f
C160 drain_left.t2 a_n2072_n3288# 0.227269f
C161 drain_left.n136 a_n2072_n3288# 2.02234f
C162 drain_left.n137 a_n2072_n3288# 0.566504f
C163 plus.n0 a_n2072_n3288# 0.055034f
C164 plus.t7 a_n2072_n3288# 1.12902f
C165 plus.t4 a_n2072_n3288# 1.12902f
C166 plus.n1 a_n2072_n3288# 0.068696f
C167 plus.t5 a_n2072_n3288# 1.12902f
C168 plus.n2 a_n2072_n3288# 0.253097f
C169 plus.t8 a_n2072_n3288# 1.12902f
C170 plus.t9 a_n2072_n3288# 1.15306f
C171 plus.n3 a_n2072_n3288# 0.430233f
C172 plus.n4 a_n2072_n3288# 0.45817f
C173 plus.n5 a_n2072_n3288# 0.459167f
C174 plus.n6 a_n2072_n3288# 0.45637f
C175 plus.n7 a_n2072_n3288# 0.009359f
C176 plus.n8 a_n2072_n3288# 0.444214f
C177 plus.n9 a_n2072_n3288# 0.478789f
C178 plus.n10 a_n2072_n3288# 0.055034f
C179 plus.t2 a_n2072_n3288# 1.12902f
C180 plus.n11 a_n2072_n3288# 0.068696f
C181 plus.t0 a_n2072_n3288# 1.12902f
C182 plus.n12 a_n2072_n3288# 0.253097f
C183 plus.t3 a_n2072_n3288# 1.12902f
C184 plus.t6 a_n2072_n3288# 1.15306f
C185 plus.n13 a_n2072_n3288# 0.430233f
C186 plus.t1 a_n2072_n3288# 1.12902f
C187 plus.n14 a_n2072_n3288# 0.45817f
C188 plus.n15 a_n2072_n3288# 0.459167f
C189 plus.n16 a_n2072_n3288# 0.45637f
C190 plus.n17 a_n2072_n3288# 0.009359f
C191 plus.n18 a_n2072_n3288# 0.444214f
C192 plus.n19 a_n2072_n3288# 1.29288f
C193 source.n0 a_n2072_n3288# 0.033382f
C194 source.n1 a_n2072_n3288# 0.025201f
C195 source.n2 a_n2072_n3288# 0.013542f
C196 source.n3 a_n2072_n3288# 0.032009f
C197 source.n4 a_n2072_n3288# 0.014339f
C198 source.n5 a_n2072_n3288# 0.025201f
C199 source.n6 a_n2072_n3288# 0.013542f
C200 source.n7 a_n2072_n3288# 0.032009f
C201 source.n8 a_n2072_n3288# 0.014339f
C202 source.n9 a_n2072_n3288# 0.025201f
C203 source.n10 a_n2072_n3288# 0.01394f
C204 source.n11 a_n2072_n3288# 0.032009f
C205 source.n12 a_n2072_n3288# 0.013542f
C206 source.n13 a_n2072_n3288# 0.014339f
C207 source.n14 a_n2072_n3288# 0.025201f
C208 source.n15 a_n2072_n3288# 0.013542f
C209 source.n16 a_n2072_n3288# 0.032009f
C210 source.n17 a_n2072_n3288# 0.014339f
C211 source.n18 a_n2072_n3288# 0.025201f
C212 source.n19 a_n2072_n3288# 0.013542f
C213 source.n20 a_n2072_n3288# 0.024007f
C214 source.n21 a_n2072_n3288# 0.022628f
C215 source.t1 a_n2072_n3288# 0.05406f
C216 source.n22 a_n2072_n3288# 0.181699f
C217 source.n23 a_n2072_n3288# 1.27136f
C218 source.n24 a_n2072_n3288# 0.013542f
C219 source.n25 a_n2072_n3288# 0.014339f
C220 source.n26 a_n2072_n3288# 0.032009f
C221 source.n27 a_n2072_n3288# 0.032009f
C222 source.n28 a_n2072_n3288# 0.014339f
C223 source.n29 a_n2072_n3288# 0.013542f
C224 source.n30 a_n2072_n3288# 0.025201f
C225 source.n31 a_n2072_n3288# 0.025201f
C226 source.n32 a_n2072_n3288# 0.013542f
C227 source.n33 a_n2072_n3288# 0.014339f
C228 source.n34 a_n2072_n3288# 0.032009f
C229 source.n35 a_n2072_n3288# 0.032009f
C230 source.n36 a_n2072_n3288# 0.014339f
C231 source.n37 a_n2072_n3288# 0.013542f
C232 source.n38 a_n2072_n3288# 0.025201f
C233 source.n39 a_n2072_n3288# 0.025201f
C234 source.n40 a_n2072_n3288# 0.013542f
C235 source.n41 a_n2072_n3288# 0.014339f
C236 source.n42 a_n2072_n3288# 0.032009f
C237 source.n43 a_n2072_n3288# 0.032009f
C238 source.n44 a_n2072_n3288# 0.032009f
C239 source.n45 a_n2072_n3288# 0.01394f
C240 source.n46 a_n2072_n3288# 0.013542f
C241 source.n47 a_n2072_n3288# 0.025201f
C242 source.n48 a_n2072_n3288# 0.025201f
C243 source.n49 a_n2072_n3288# 0.013542f
C244 source.n50 a_n2072_n3288# 0.014339f
C245 source.n51 a_n2072_n3288# 0.032009f
C246 source.n52 a_n2072_n3288# 0.032009f
C247 source.n53 a_n2072_n3288# 0.014339f
C248 source.n54 a_n2072_n3288# 0.013542f
C249 source.n55 a_n2072_n3288# 0.025201f
C250 source.n56 a_n2072_n3288# 0.025201f
C251 source.n57 a_n2072_n3288# 0.013542f
C252 source.n58 a_n2072_n3288# 0.014339f
C253 source.n59 a_n2072_n3288# 0.032009f
C254 source.n60 a_n2072_n3288# 0.065685f
C255 source.n61 a_n2072_n3288# 0.014339f
C256 source.n62 a_n2072_n3288# 0.013542f
C257 source.n63 a_n2072_n3288# 0.05412f
C258 source.n64 a_n2072_n3288# 0.036251f
C259 source.n65 a_n2072_n3288# 1.07159f
C260 source.t5 a_n2072_n3288# 0.238978f
C261 source.t8 a_n2072_n3288# 0.238978f
C262 source.n66 a_n2072_n3288# 2.04614f
C263 source.n67 a_n2072_n3288# 0.41586f
C264 source.t2 a_n2072_n3288# 0.238978f
C265 source.t3 a_n2072_n3288# 0.238978f
C266 source.n68 a_n2072_n3288# 2.04614f
C267 source.n69 a_n2072_n3288# 0.41446f
C268 source.n70 a_n2072_n3288# 0.033382f
C269 source.n71 a_n2072_n3288# 0.025201f
C270 source.n72 a_n2072_n3288# 0.013542f
C271 source.n73 a_n2072_n3288# 0.032009f
C272 source.n74 a_n2072_n3288# 0.014339f
C273 source.n75 a_n2072_n3288# 0.025201f
C274 source.n76 a_n2072_n3288# 0.013542f
C275 source.n77 a_n2072_n3288# 0.032009f
C276 source.n78 a_n2072_n3288# 0.014339f
C277 source.n79 a_n2072_n3288# 0.025201f
C278 source.n80 a_n2072_n3288# 0.01394f
C279 source.n81 a_n2072_n3288# 0.032009f
C280 source.n82 a_n2072_n3288# 0.013542f
C281 source.n83 a_n2072_n3288# 0.014339f
C282 source.n84 a_n2072_n3288# 0.025201f
C283 source.n85 a_n2072_n3288# 0.013542f
C284 source.n86 a_n2072_n3288# 0.032009f
C285 source.n87 a_n2072_n3288# 0.014339f
C286 source.n88 a_n2072_n3288# 0.025201f
C287 source.n89 a_n2072_n3288# 0.013542f
C288 source.n90 a_n2072_n3288# 0.024007f
C289 source.n91 a_n2072_n3288# 0.022628f
C290 source.t15 a_n2072_n3288# 0.05406f
C291 source.n92 a_n2072_n3288# 0.181699f
C292 source.n93 a_n2072_n3288# 1.27136f
C293 source.n94 a_n2072_n3288# 0.013542f
C294 source.n95 a_n2072_n3288# 0.014339f
C295 source.n96 a_n2072_n3288# 0.032009f
C296 source.n97 a_n2072_n3288# 0.032009f
C297 source.n98 a_n2072_n3288# 0.014339f
C298 source.n99 a_n2072_n3288# 0.013542f
C299 source.n100 a_n2072_n3288# 0.025201f
C300 source.n101 a_n2072_n3288# 0.025201f
C301 source.n102 a_n2072_n3288# 0.013542f
C302 source.n103 a_n2072_n3288# 0.014339f
C303 source.n104 a_n2072_n3288# 0.032009f
C304 source.n105 a_n2072_n3288# 0.032009f
C305 source.n106 a_n2072_n3288# 0.014339f
C306 source.n107 a_n2072_n3288# 0.013542f
C307 source.n108 a_n2072_n3288# 0.025201f
C308 source.n109 a_n2072_n3288# 0.025201f
C309 source.n110 a_n2072_n3288# 0.013542f
C310 source.n111 a_n2072_n3288# 0.014339f
C311 source.n112 a_n2072_n3288# 0.032009f
C312 source.n113 a_n2072_n3288# 0.032009f
C313 source.n114 a_n2072_n3288# 0.032009f
C314 source.n115 a_n2072_n3288# 0.01394f
C315 source.n116 a_n2072_n3288# 0.013542f
C316 source.n117 a_n2072_n3288# 0.025201f
C317 source.n118 a_n2072_n3288# 0.025201f
C318 source.n119 a_n2072_n3288# 0.013542f
C319 source.n120 a_n2072_n3288# 0.014339f
C320 source.n121 a_n2072_n3288# 0.032009f
C321 source.n122 a_n2072_n3288# 0.032009f
C322 source.n123 a_n2072_n3288# 0.014339f
C323 source.n124 a_n2072_n3288# 0.013542f
C324 source.n125 a_n2072_n3288# 0.025201f
C325 source.n126 a_n2072_n3288# 0.025201f
C326 source.n127 a_n2072_n3288# 0.013542f
C327 source.n128 a_n2072_n3288# 0.014339f
C328 source.n129 a_n2072_n3288# 0.032009f
C329 source.n130 a_n2072_n3288# 0.065685f
C330 source.n131 a_n2072_n3288# 0.014339f
C331 source.n132 a_n2072_n3288# 0.013542f
C332 source.n133 a_n2072_n3288# 0.05412f
C333 source.n134 a_n2072_n3288# 0.036251f
C334 source.n135 a_n2072_n3288# 0.176005f
C335 source.t17 a_n2072_n3288# 0.238978f
C336 source.t16 a_n2072_n3288# 0.238978f
C337 source.n136 a_n2072_n3288# 2.04614f
C338 source.n137 a_n2072_n3288# 0.41586f
C339 source.t13 a_n2072_n3288# 0.238978f
C340 source.t14 a_n2072_n3288# 0.238978f
C341 source.n138 a_n2072_n3288# 2.04614f
C342 source.n139 a_n2072_n3288# 1.79806f
C343 source.t9 a_n2072_n3288# 0.238978f
C344 source.t0 a_n2072_n3288# 0.238978f
C345 source.n140 a_n2072_n3288# 2.04612f
C346 source.n141 a_n2072_n3288# 1.79807f
C347 source.t4 a_n2072_n3288# 0.238978f
C348 source.t6 a_n2072_n3288# 0.238978f
C349 source.n142 a_n2072_n3288# 2.04612f
C350 source.n143 a_n2072_n3288# 0.415873f
C351 source.n144 a_n2072_n3288# 0.033382f
C352 source.n145 a_n2072_n3288# 0.025201f
C353 source.n146 a_n2072_n3288# 0.013542f
C354 source.n147 a_n2072_n3288# 0.032009f
C355 source.n148 a_n2072_n3288# 0.014339f
C356 source.n149 a_n2072_n3288# 0.025201f
C357 source.n150 a_n2072_n3288# 0.013542f
C358 source.n151 a_n2072_n3288# 0.032009f
C359 source.n152 a_n2072_n3288# 0.014339f
C360 source.n153 a_n2072_n3288# 0.025201f
C361 source.n154 a_n2072_n3288# 0.01394f
C362 source.n155 a_n2072_n3288# 0.032009f
C363 source.n156 a_n2072_n3288# 0.014339f
C364 source.n157 a_n2072_n3288# 0.025201f
C365 source.n158 a_n2072_n3288# 0.013542f
C366 source.n159 a_n2072_n3288# 0.032009f
C367 source.n160 a_n2072_n3288# 0.014339f
C368 source.n161 a_n2072_n3288# 0.025201f
C369 source.n162 a_n2072_n3288# 0.013542f
C370 source.n163 a_n2072_n3288# 0.024007f
C371 source.n164 a_n2072_n3288# 0.022628f
C372 source.t7 a_n2072_n3288# 0.05406f
C373 source.n165 a_n2072_n3288# 0.181699f
C374 source.n166 a_n2072_n3288# 1.27136f
C375 source.n167 a_n2072_n3288# 0.013542f
C376 source.n168 a_n2072_n3288# 0.014339f
C377 source.n169 a_n2072_n3288# 0.032009f
C378 source.n170 a_n2072_n3288# 0.032009f
C379 source.n171 a_n2072_n3288# 0.014339f
C380 source.n172 a_n2072_n3288# 0.013542f
C381 source.n173 a_n2072_n3288# 0.025201f
C382 source.n174 a_n2072_n3288# 0.025201f
C383 source.n175 a_n2072_n3288# 0.013542f
C384 source.n176 a_n2072_n3288# 0.014339f
C385 source.n177 a_n2072_n3288# 0.032009f
C386 source.n178 a_n2072_n3288# 0.032009f
C387 source.n179 a_n2072_n3288# 0.014339f
C388 source.n180 a_n2072_n3288# 0.013542f
C389 source.n181 a_n2072_n3288# 0.025201f
C390 source.n182 a_n2072_n3288# 0.025201f
C391 source.n183 a_n2072_n3288# 0.013542f
C392 source.n184 a_n2072_n3288# 0.013542f
C393 source.n185 a_n2072_n3288# 0.014339f
C394 source.n186 a_n2072_n3288# 0.032009f
C395 source.n187 a_n2072_n3288# 0.032009f
C396 source.n188 a_n2072_n3288# 0.032009f
C397 source.n189 a_n2072_n3288# 0.01394f
C398 source.n190 a_n2072_n3288# 0.013542f
C399 source.n191 a_n2072_n3288# 0.025201f
C400 source.n192 a_n2072_n3288# 0.025201f
C401 source.n193 a_n2072_n3288# 0.013542f
C402 source.n194 a_n2072_n3288# 0.014339f
C403 source.n195 a_n2072_n3288# 0.032009f
C404 source.n196 a_n2072_n3288# 0.032009f
C405 source.n197 a_n2072_n3288# 0.014339f
C406 source.n198 a_n2072_n3288# 0.013542f
C407 source.n199 a_n2072_n3288# 0.025201f
C408 source.n200 a_n2072_n3288# 0.025201f
C409 source.n201 a_n2072_n3288# 0.013542f
C410 source.n202 a_n2072_n3288# 0.014339f
C411 source.n203 a_n2072_n3288# 0.032009f
C412 source.n204 a_n2072_n3288# 0.065685f
C413 source.n205 a_n2072_n3288# 0.014339f
C414 source.n206 a_n2072_n3288# 0.013542f
C415 source.n207 a_n2072_n3288# 0.05412f
C416 source.n208 a_n2072_n3288# 0.036251f
C417 source.n209 a_n2072_n3288# 0.176005f
C418 source.t10 a_n2072_n3288# 0.238978f
C419 source.t18 a_n2072_n3288# 0.238978f
C420 source.n210 a_n2072_n3288# 2.04612f
C421 source.n211 a_n2072_n3288# 0.414472f
C422 source.t12 a_n2072_n3288# 0.238978f
C423 source.t19 a_n2072_n3288# 0.238978f
C424 source.n212 a_n2072_n3288# 2.04612f
C425 source.n213 a_n2072_n3288# 0.415873f
C426 source.n214 a_n2072_n3288# 0.033382f
C427 source.n215 a_n2072_n3288# 0.025201f
C428 source.n216 a_n2072_n3288# 0.013542f
C429 source.n217 a_n2072_n3288# 0.032009f
C430 source.n218 a_n2072_n3288# 0.014339f
C431 source.n219 a_n2072_n3288# 0.025201f
C432 source.n220 a_n2072_n3288# 0.013542f
C433 source.n221 a_n2072_n3288# 0.032009f
C434 source.n222 a_n2072_n3288# 0.014339f
C435 source.n223 a_n2072_n3288# 0.025201f
C436 source.n224 a_n2072_n3288# 0.01394f
C437 source.n225 a_n2072_n3288# 0.032009f
C438 source.n226 a_n2072_n3288# 0.014339f
C439 source.n227 a_n2072_n3288# 0.025201f
C440 source.n228 a_n2072_n3288# 0.013542f
C441 source.n229 a_n2072_n3288# 0.032009f
C442 source.n230 a_n2072_n3288# 0.014339f
C443 source.n231 a_n2072_n3288# 0.025201f
C444 source.n232 a_n2072_n3288# 0.013542f
C445 source.n233 a_n2072_n3288# 0.024007f
C446 source.n234 a_n2072_n3288# 0.022628f
C447 source.t11 a_n2072_n3288# 0.05406f
C448 source.n235 a_n2072_n3288# 0.181699f
C449 source.n236 a_n2072_n3288# 1.27136f
C450 source.n237 a_n2072_n3288# 0.013542f
C451 source.n238 a_n2072_n3288# 0.014339f
C452 source.n239 a_n2072_n3288# 0.032009f
C453 source.n240 a_n2072_n3288# 0.032009f
C454 source.n241 a_n2072_n3288# 0.014339f
C455 source.n242 a_n2072_n3288# 0.013542f
C456 source.n243 a_n2072_n3288# 0.025201f
C457 source.n244 a_n2072_n3288# 0.025201f
C458 source.n245 a_n2072_n3288# 0.013542f
C459 source.n246 a_n2072_n3288# 0.014339f
C460 source.n247 a_n2072_n3288# 0.032009f
C461 source.n248 a_n2072_n3288# 0.032009f
C462 source.n249 a_n2072_n3288# 0.014339f
C463 source.n250 a_n2072_n3288# 0.013542f
C464 source.n251 a_n2072_n3288# 0.025201f
C465 source.n252 a_n2072_n3288# 0.025201f
C466 source.n253 a_n2072_n3288# 0.013542f
C467 source.n254 a_n2072_n3288# 0.013542f
C468 source.n255 a_n2072_n3288# 0.014339f
C469 source.n256 a_n2072_n3288# 0.032009f
C470 source.n257 a_n2072_n3288# 0.032009f
C471 source.n258 a_n2072_n3288# 0.032009f
C472 source.n259 a_n2072_n3288# 0.01394f
C473 source.n260 a_n2072_n3288# 0.013542f
C474 source.n261 a_n2072_n3288# 0.025201f
C475 source.n262 a_n2072_n3288# 0.025201f
C476 source.n263 a_n2072_n3288# 0.013542f
C477 source.n264 a_n2072_n3288# 0.014339f
C478 source.n265 a_n2072_n3288# 0.032009f
C479 source.n266 a_n2072_n3288# 0.032009f
C480 source.n267 a_n2072_n3288# 0.014339f
C481 source.n268 a_n2072_n3288# 0.013542f
C482 source.n269 a_n2072_n3288# 0.025201f
C483 source.n270 a_n2072_n3288# 0.025201f
C484 source.n271 a_n2072_n3288# 0.013542f
C485 source.n272 a_n2072_n3288# 0.014339f
C486 source.n273 a_n2072_n3288# 0.032009f
C487 source.n274 a_n2072_n3288# 0.065685f
C488 source.n275 a_n2072_n3288# 0.014339f
C489 source.n276 a_n2072_n3288# 0.013542f
C490 source.n277 a_n2072_n3288# 0.05412f
C491 source.n278 a_n2072_n3288# 0.036251f
C492 source.n279 a_n2072_n3288# 0.306298f
C493 source.n280 a_n2072_n3288# 1.60104f
C494 drain_right.n0 a_n2072_n3288# 0.031585f
C495 drain_right.n1 a_n2072_n3288# 0.023845f
C496 drain_right.n2 a_n2072_n3288# 0.012813f
C497 drain_right.n3 a_n2072_n3288# 0.030286f
C498 drain_right.n4 a_n2072_n3288# 0.013567f
C499 drain_right.n5 a_n2072_n3288# 0.023845f
C500 drain_right.n6 a_n2072_n3288# 0.012813f
C501 drain_right.n7 a_n2072_n3288# 0.030286f
C502 drain_right.n8 a_n2072_n3288# 0.013567f
C503 drain_right.n9 a_n2072_n3288# 0.023845f
C504 drain_right.n10 a_n2072_n3288# 0.01319f
C505 drain_right.n11 a_n2072_n3288# 0.030286f
C506 drain_right.n12 a_n2072_n3288# 0.013567f
C507 drain_right.n13 a_n2072_n3288# 0.023845f
C508 drain_right.n14 a_n2072_n3288# 0.012813f
C509 drain_right.n15 a_n2072_n3288# 0.030286f
C510 drain_right.n16 a_n2072_n3288# 0.013567f
C511 drain_right.n17 a_n2072_n3288# 0.023845f
C512 drain_right.n18 a_n2072_n3288# 0.012813f
C513 drain_right.n19 a_n2072_n3288# 0.022714f
C514 drain_right.n20 a_n2072_n3288# 0.02141f
C515 drain_right.t4 a_n2072_n3288# 0.05115f
C516 drain_right.n21 a_n2072_n3288# 0.171918f
C517 drain_right.n22 a_n2072_n3288# 1.20293f
C518 drain_right.n23 a_n2072_n3288# 0.012813f
C519 drain_right.n24 a_n2072_n3288# 0.013567f
C520 drain_right.n25 a_n2072_n3288# 0.030286f
C521 drain_right.n26 a_n2072_n3288# 0.030286f
C522 drain_right.n27 a_n2072_n3288# 0.013567f
C523 drain_right.n28 a_n2072_n3288# 0.012813f
C524 drain_right.n29 a_n2072_n3288# 0.023845f
C525 drain_right.n30 a_n2072_n3288# 0.023845f
C526 drain_right.n31 a_n2072_n3288# 0.012813f
C527 drain_right.n32 a_n2072_n3288# 0.013567f
C528 drain_right.n33 a_n2072_n3288# 0.030286f
C529 drain_right.n34 a_n2072_n3288# 0.030286f
C530 drain_right.n35 a_n2072_n3288# 0.013567f
C531 drain_right.n36 a_n2072_n3288# 0.012813f
C532 drain_right.n37 a_n2072_n3288# 0.023845f
C533 drain_right.n38 a_n2072_n3288# 0.023845f
C534 drain_right.n39 a_n2072_n3288# 0.012813f
C535 drain_right.n40 a_n2072_n3288# 0.012813f
C536 drain_right.n41 a_n2072_n3288# 0.013567f
C537 drain_right.n42 a_n2072_n3288# 0.030286f
C538 drain_right.n43 a_n2072_n3288# 0.030286f
C539 drain_right.n44 a_n2072_n3288# 0.030286f
C540 drain_right.n45 a_n2072_n3288# 0.01319f
C541 drain_right.n46 a_n2072_n3288# 0.012813f
C542 drain_right.n47 a_n2072_n3288# 0.023845f
C543 drain_right.n48 a_n2072_n3288# 0.023845f
C544 drain_right.n49 a_n2072_n3288# 0.012813f
C545 drain_right.n50 a_n2072_n3288# 0.013567f
C546 drain_right.n51 a_n2072_n3288# 0.030286f
C547 drain_right.n52 a_n2072_n3288# 0.030286f
C548 drain_right.n53 a_n2072_n3288# 0.013567f
C549 drain_right.n54 a_n2072_n3288# 0.012813f
C550 drain_right.n55 a_n2072_n3288# 0.023845f
C551 drain_right.n56 a_n2072_n3288# 0.023845f
C552 drain_right.n57 a_n2072_n3288# 0.012813f
C553 drain_right.n58 a_n2072_n3288# 0.013567f
C554 drain_right.n59 a_n2072_n3288# 0.030286f
C555 drain_right.n60 a_n2072_n3288# 0.062149f
C556 drain_right.n61 a_n2072_n3288# 0.013567f
C557 drain_right.n62 a_n2072_n3288# 0.012813f
C558 drain_right.n63 a_n2072_n3288# 0.051207f
C559 drain_right.n64 a_n2072_n3288# 0.053228f
C560 drain_right.t2 a_n2072_n3288# 0.226114f
C561 drain_right.t5 a_n2072_n3288# 0.226114f
C562 drain_right.n65 a_n2072_n3288# 2.01207f
C563 drain_right.n66 a_n2072_n3288# 0.408456f
C564 drain_right.t3 a_n2072_n3288# 0.226114f
C565 drain_right.t6 a_n2072_n3288# 0.226114f
C566 drain_right.n67 a_n2072_n3288# 2.01585f
C567 drain_right.n68 a_n2072_n3288# 1.53419f
C568 drain_right.t8 a_n2072_n3288# 0.226114f
C569 drain_right.t0 a_n2072_n3288# 0.226114f
C570 drain_right.n69 a_n2072_n3288# 2.01785f
C571 drain_right.t9 a_n2072_n3288# 0.226114f
C572 drain_right.t7 a_n2072_n3288# 0.226114f
C573 drain_right.n70 a_n2072_n3288# 2.01207f
C574 drain_right.n71 a_n2072_n3288# 0.703432f
C575 drain_right.n72 a_n2072_n3288# 0.031585f
C576 drain_right.n73 a_n2072_n3288# 0.023845f
C577 drain_right.n74 a_n2072_n3288# 0.012813f
C578 drain_right.n75 a_n2072_n3288# 0.030286f
C579 drain_right.n76 a_n2072_n3288# 0.013567f
C580 drain_right.n77 a_n2072_n3288# 0.023845f
C581 drain_right.n78 a_n2072_n3288# 0.012813f
C582 drain_right.n79 a_n2072_n3288# 0.030286f
C583 drain_right.n80 a_n2072_n3288# 0.013567f
C584 drain_right.n81 a_n2072_n3288# 0.023845f
C585 drain_right.n82 a_n2072_n3288# 0.01319f
C586 drain_right.n83 a_n2072_n3288# 0.030286f
C587 drain_right.n84 a_n2072_n3288# 0.012813f
C588 drain_right.n85 a_n2072_n3288# 0.013567f
C589 drain_right.n86 a_n2072_n3288# 0.023845f
C590 drain_right.n87 a_n2072_n3288# 0.012813f
C591 drain_right.n88 a_n2072_n3288# 0.030286f
C592 drain_right.n89 a_n2072_n3288# 0.013567f
C593 drain_right.n90 a_n2072_n3288# 0.023845f
C594 drain_right.n91 a_n2072_n3288# 0.012813f
C595 drain_right.n92 a_n2072_n3288# 0.022714f
C596 drain_right.n93 a_n2072_n3288# 0.02141f
C597 drain_right.t1 a_n2072_n3288# 0.05115f
C598 drain_right.n94 a_n2072_n3288# 0.171918f
C599 drain_right.n95 a_n2072_n3288# 1.20293f
C600 drain_right.n96 a_n2072_n3288# 0.012813f
C601 drain_right.n97 a_n2072_n3288# 0.013567f
C602 drain_right.n98 a_n2072_n3288# 0.030286f
C603 drain_right.n99 a_n2072_n3288# 0.030286f
C604 drain_right.n100 a_n2072_n3288# 0.013567f
C605 drain_right.n101 a_n2072_n3288# 0.012813f
C606 drain_right.n102 a_n2072_n3288# 0.023845f
C607 drain_right.n103 a_n2072_n3288# 0.023845f
C608 drain_right.n104 a_n2072_n3288# 0.012813f
C609 drain_right.n105 a_n2072_n3288# 0.013567f
C610 drain_right.n106 a_n2072_n3288# 0.030286f
C611 drain_right.n107 a_n2072_n3288# 0.030286f
C612 drain_right.n108 a_n2072_n3288# 0.013567f
C613 drain_right.n109 a_n2072_n3288# 0.012813f
C614 drain_right.n110 a_n2072_n3288# 0.023845f
C615 drain_right.n111 a_n2072_n3288# 0.023845f
C616 drain_right.n112 a_n2072_n3288# 0.012813f
C617 drain_right.n113 a_n2072_n3288# 0.013567f
C618 drain_right.n114 a_n2072_n3288# 0.030286f
C619 drain_right.n115 a_n2072_n3288# 0.030286f
C620 drain_right.n116 a_n2072_n3288# 0.030286f
C621 drain_right.n117 a_n2072_n3288# 0.01319f
C622 drain_right.n118 a_n2072_n3288# 0.012813f
C623 drain_right.n119 a_n2072_n3288# 0.023845f
C624 drain_right.n120 a_n2072_n3288# 0.023845f
C625 drain_right.n121 a_n2072_n3288# 0.012813f
C626 drain_right.n122 a_n2072_n3288# 0.013567f
C627 drain_right.n123 a_n2072_n3288# 0.030286f
C628 drain_right.n124 a_n2072_n3288# 0.030286f
C629 drain_right.n125 a_n2072_n3288# 0.013567f
C630 drain_right.n126 a_n2072_n3288# 0.012813f
C631 drain_right.n127 a_n2072_n3288# 0.023845f
C632 drain_right.n128 a_n2072_n3288# 0.023845f
C633 drain_right.n129 a_n2072_n3288# 0.012813f
C634 drain_right.n130 a_n2072_n3288# 0.013567f
C635 drain_right.n131 a_n2072_n3288# 0.030286f
C636 drain_right.n132 a_n2072_n3288# 0.062149f
C637 drain_right.n133 a_n2072_n3288# 0.013567f
C638 drain_right.n134 a_n2072_n3288# 0.012813f
C639 drain_right.n135 a_n2072_n3288# 0.051207f
C640 drain_right.n136 a_n2072_n3288# 0.050798f
C641 drain_right.n137 a_n2072_n3288# 0.342666f
C642 minus.n0 a_n2072_n3288# 0.054265f
C643 minus.t2 a_n2072_n3288# 1.11324f
C644 minus.n1 a_n2072_n3288# 0.452752f
C645 minus.t5 a_n2072_n3288# 1.11324f
C646 minus.t4 a_n2072_n3288# 1.13695f
C647 minus.t3 a_n2072_n3288# 1.11324f
C648 minus.n2 a_n2072_n3288# 0.451768f
C649 minus.n3 a_n2072_n3288# 0.424222f
C650 minus.n4 a_n2072_n3288# 0.249561f
C651 minus.n5 a_n2072_n3288# 0.067736f
C652 minus.n6 a_n2072_n3288# 0.449994f
C653 minus.n7 a_n2072_n3288# 0.009228f
C654 minus.t6 a_n2072_n3288# 1.11324f
C655 minus.n8 a_n2072_n3288# 0.438008f
C656 minus.n9 a_n2072_n3288# 1.50186f
C657 minus.n10 a_n2072_n3288# 0.054265f
C658 minus.t7 a_n2072_n3288# 1.11324f
C659 minus.n11 a_n2072_n3288# 0.452752f
C660 minus.t9 a_n2072_n3288# 1.13695f
C661 minus.t1 a_n2072_n3288# 1.11324f
C662 minus.n12 a_n2072_n3288# 0.451768f
C663 minus.n13 a_n2072_n3288# 0.424222f
C664 minus.n14 a_n2072_n3288# 0.249561f
C665 minus.n15 a_n2072_n3288# 0.067736f
C666 minus.t0 a_n2072_n3288# 1.11324f
C667 minus.n16 a_n2072_n3288# 0.449994f
C668 minus.n17 a_n2072_n3288# 0.009228f
C669 minus.t8 a_n2072_n3288# 1.11324f
C670 minus.n18 a_n2072_n3288# 0.438008f
C671 minus.n19 a_n2072_n3288# 0.282656f
C672 minus.n20 a_n2072_n3288# 1.81388f
.ends

