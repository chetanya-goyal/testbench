* NGSPICE file created from diffpair647.ext - technology: sky130A

.subckt diffpair647 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t25 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X1 drain_right.t14 minus.t1 source.t23 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X2 source.t16 minus.t2 drain_right.t13 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X3 source.t3 plus.t0 drain_left.t15 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X4 drain_left.t14 plus.t1 source.t7 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X5 source.t9 plus.t2 drain_left.t13 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X6 drain_left.t12 plus.t3 source.t0 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X7 a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X8 a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X9 source.t21 minus.t3 drain_right.t12 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X10 source.t13 plus.t4 drain_left.t11 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X11 a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X12 drain_right.t11 minus.t4 source.t28 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X13 drain_right.t10 minus.t5 source.t30 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X14 source.t18 minus.t6 drain_right.t9 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X15 drain_left.t10 plus.t5 source.t1 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X16 source.t24 minus.t7 drain_right.t8 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 drain_left.t9 plus.t6 source.t11 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X18 drain_left.t8 plus.t7 source.t15 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X19 source.t2 plus.t8 drain_left.t7 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X20 drain_right.t7 minus.t8 source.t31 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X21 drain_right.t6 minus.t9 source.t27 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X22 drain_right.t5 minus.t10 source.t17 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X23 source.t20 minus.t11 drain_right.t4 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X24 drain_left.t6 plus.t9 source.t14 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X25 source.t26 minus.t12 drain_right.t3 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X26 drain_right.t2 minus.t13 source.t29 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X27 source.t4 plus.t10 drain_left.t5 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X28 source.t8 plus.t11 drain_left.t4 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X29 source.t10 plus.t12 drain_left.t3 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X30 a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X31 drain_left.t2 plus.t13 source.t5 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X32 drain_left.t1 plus.t14 source.t12 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X33 source.t19 minus.t14 drain_right.t1 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X34 source.t6 plus.t15 drain_left.t0 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X35 source.t22 minus.t15 drain_right.t0 a_n1886_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
R0 minus.n21 minus.t11 4265.7
R1 minus.n5 minus.t4 4265.7
R2 minus.n44 minus.t1 4265.7
R3 minus.n28 minus.t2 4265.7
R4 minus.n20 minus.t9 4225.53
R5 minus.n1 minus.t12 4225.53
R6 minus.n14 minus.t5 4225.53
R7 minus.n12 minus.t7 4225.53
R8 minus.n3 minus.t8 4225.53
R9 minus.n6 minus.t3 4225.53
R10 minus.n43 minus.t15 4225.53
R11 minus.n24 minus.t13 4225.53
R12 minus.n37 minus.t6 4225.53
R13 minus.n35 minus.t0 4225.53
R14 minus.n26 minus.t14 4225.53
R15 minus.n29 minus.t10 4225.53
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 69.3793
R39 minus.n11 minus.n3 69.3793
R40 minus.n34 minus.n26 69.3793
R41 minus.n38 minus.n24 69.3793
R42 minus.n21 minus.n20 54.7732
R43 minus.n6 minus.n5 54.7732
R44 minus.n29 minus.n28 54.7732
R45 minus.n44 minus.n43 54.7732
R46 minus.n14 minus.n13 47.4702
R47 minus.n13 minus.n12 47.4702
R48 minus.n36 minus.n35 47.4702
R49 minus.n37 minus.n36 47.4702
R50 minus.n46 minus.n22 46.1179
R51 minus.n15 minus.n14 25.5611
R52 minus.n12 minus.n11 25.5611
R53 minus.n35 minus.n34 25.5611
R54 minus.n38 minus.n37 25.5611
R55 minus.n20 minus.n19 18.2581
R56 minus.n7 minus.n6 18.2581
R57 minus.n30 minus.n29 18.2581
R58 minus.n43 minus.n42 18.2581
R59 minus.n46 minus.n45 6.50429
R60 minus.n18 minus.n1 3.65202
R61 minus.n8 minus.n3 3.65202
R62 minus.n31 minus.n26 3.65202
R63 minus.n41 minus.n24 3.65202
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 source.n7 source.t2 43.2366
R80 source.n8 source.t28 43.2366
R81 source.n15 source.t20 43.2366
R82 source.n31 source.t23 43.2365
R83 source.n24 source.t16 43.2365
R84 source.n23 source.t1 43.2365
R85 source.n16 source.t9 43.2365
R86 source.n0 source.t15 43.2365
R87 source.n30 source.n29 42.0366
R88 source.n28 source.n27 42.0366
R89 source.n26 source.n25 42.0366
R90 source.n22 source.n21 42.0366
R91 source.n20 source.n19 42.0366
R92 source.n18 source.n17 42.0366
R93 source.n2 source.n1 42.0366
R94 source.n4 source.n3 42.0366
R95 source.n6 source.n5 42.0366
R96 source.n10 source.n9 42.0366
R97 source.n12 source.n11 42.0366
R98 source.n14 source.n13 42.0366
R99 source.n16 source.n15 31.6966
R100 source.n32 source.n0 26.1535
R101 source.n32 source.n31 5.5436
R102 source.n29 source.t29 1.2005
R103 source.n29 source.t22 1.2005
R104 source.n27 source.t25 1.2005
R105 source.n27 source.t18 1.2005
R106 source.n25 source.t17 1.2005
R107 source.n25 source.t19 1.2005
R108 source.n21 source.t7 1.2005
R109 source.n21 source.t4 1.2005
R110 source.n19 source.t11 1.2005
R111 source.n19 source.t13 1.2005
R112 source.n17 source.t0 1.2005
R113 source.n17 source.t3 1.2005
R114 source.n1 source.t5 1.2005
R115 source.n1 source.t8 1.2005
R116 source.n3 source.t14 1.2005
R117 source.n3 source.t6 1.2005
R118 source.n5 source.t12 1.2005
R119 source.n5 source.t10 1.2005
R120 source.n9 source.t31 1.2005
R121 source.n9 source.t21 1.2005
R122 source.n11 source.t30 1.2005
R123 source.n11 source.t24 1.2005
R124 source.n13 source.t27 1.2005
R125 source.n13 source.t26 1.2005
R126 source.n15 source.n14 0.560845
R127 source.n14 source.n12 0.560845
R128 source.n12 source.n10 0.560845
R129 source.n10 source.n8 0.560845
R130 source.n7 source.n6 0.560845
R131 source.n6 source.n4 0.560845
R132 source.n4 source.n2 0.560845
R133 source.n2 source.n0 0.560845
R134 source.n18 source.n16 0.560845
R135 source.n20 source.n18 0.560845
R136 source.n22 source.n20 0.560845
R137 source.n23 source.n22 0.560845
R138 source.n26 source.n24 0.560845
R139 source.n28 source.n26 0.560845
R140 source.n30 source.n28 0.560845
R141 source.n31 source.n30 0.560845
R142 source.n8 source.n7 0.470328
R143 source.n24 source.n23 0.470328
R144 source source.n32 0.188
R145 drain_right.n5 drain_right.n3 59.2758
R146 drain_right.n2 drain_right.n0 59.2758
R147 drain_right.n9 drain_right.n7 59.2756
R148 drain_right.n5 drain_right.n4 58.7154
R149 drain_right.n2 drain_right.n1 58.7154
R150 drain_right.n9 drain_right.n8 58.7154
R151 drain_right.n11 drain_right.n10 58.7154
R152 drain_right.n13 drain_right.n12 58.7154
R153 drain_right drain_right.n6 40.3046
R154 drain_right drain_right.n13 6.21356
R155 drain_right.n3 drain_right.t0 1.2005
R156 drain_right.n3 drain_right.t14 1.2005
R157 drain_right.n4 drain_right.t9 1.2005
R158 drain_right.n4 drain_right.t2 1.2005
R159 drain_right.n1 drain_right.t1 1.2005
R160 drain_right.n1 drain_right.t15 1.2005
R161 drain_right.n0 drain_right.t13 1.2005
R162 drain_right.n0 drain_right.t5 1.2005
R163 drain_right.n7 drain_right.t12 1.2005
R164 drain_right.n7 drain_right.t11 1.2005
R165 drain_right.n8 drain_right.t8 1.2005
R166 drain_right.n8 drain_right.t7 1.2005
R167 drain_right.n10 drain_right.t3 1.2005
R168 drain_right.n10 drain_right.t10 1.2005
R169 drain_right.n12 drain_right.t4 1.2005
R170 drain_right.n12 drain_right.t6 1.2005
R171 drain_right.n13 drain_right.n11 0.560845
R172 drain_right.n11 drain_right.n9 0.560845
R173 drain_right.n6 drain_right.n5 0.225326
R174 drain_right.n6 drain_right.n2 0.225326
R175 plus.n5 plus.t8 4265.7
R176 plus.n21 plus.t7 4265.7
R177 plus.n28 plus.t5 4265.7
R178 plus.n44 plus.t2 4265.7
R179 plus.n6 plus.t14 4225.53
R180 plus.n3 plus.t12 4225.53
R181 plus.n12 plus.t9 4225.53
R182 plus.n14 plus.t15 4225.53
R183 plus.n1 plus.t13 4225.53
R184 plus.n20 plus.t11 4225.53
R185 plus.n29 plus.t10 4225.53
R186 plus.n26 plus.t1 4225.53
R187 plus.n35 plus.t4 4225.53
R188 plus.n37 plus.t6 4225.53
R189 plus.n24 plus.t0 4225.53
R190 plus.n43 plus.t3 4225.53
R191 plus.n5 plus.n4 161.489
R192 plus.n28 plus.n27 161.489
R193 plus.n7 plus.n4 161.3
R194 plus.n9 plus.n8 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n13 plus.n2 161.3
R197 plus.n16 plus.n15 161.3
R198 plus.n18 plus.n17 161.3
R199 plus.n19 plus.n0 161.3
R200 plus.n22 plus.n21 161.3
R201 plus.n30 plus.n27 161.3
R202 plus.n32 plus.n31 161.3
R203 plus.n34 plus.n33 161.3
R204 plus.n36 plus.n25 161.3
R205 plus.n39 plus.n38 161.3
R206 plus.n41 plus.n40 161.3
R207 plus.n42 plus.n23 161.3
R208 plus.n45 plus.n44 161.3
R209 plus.n8 plus.n7 73.0308
R210 plus.n19 plus.n18 73.0308
R211 plus.n42 plus.n41 73.0308
R212 plus.n31 plus.n30 73.0308
R213 plus.n11 plus.n3 69.3793
R214 plus.n15 plus.n1 69.3793
R215 plus.n38 plus.n24 69.3793
R216 plus.n34 plus.n26 69.3793
R217 plus.n6 plus.n5 54.7732
R218 plus.n21 plus.n20 54.7732
R219 plus.n44 plus.n43 54.7732
R220 plus.n29 plus.n28 54.7732
R221 plus.n13 plus.n12 47.4702
R222 plus.n14 plus.n13 47.4702
R223 plus.n37 plus.n36 47.4702
R224 plus.n36 plus.n35 47.4702
R225 plus plus.n45 35.0748
R226 plus.n12 plus.n11 25.5611
R227 plus.n15 plus.n14 25.5611
R228 plus.n38 plus.n37 25.5611
R229 plus.n35 plus.n34 25.5611
R230 plus.n7 plus.n6 18.2581
R231 plus.n20 plus.n19 18.2581
R232 plus.n43 plus.n42 18.2581
R233 plus.n30 plus.n29 18.2581
R234 plus plus.n22 17.0725
R235 plus.n8 plus.n3 3.65202
R236 plus.n18 plus.n1 3.65202
R237 plus.n41 plus.n24 3.65202
R238 plus.n31 plus.n26 3.65202
R239 plus.n9 plus.n4 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n2 0.189894
R242 plus.n16 plus.n2 0.189894
R243 plus.n17 plus.n16 0.189894
R244 plus.n17 plus.n0 0.189894
R245 plus.n22 plus.n0 0.189894
R246 plus.n45 plus.n23 0.189894
R247 plus.n40 plus.n23 0.189894
R248 plus.n40 plus.n39 0.189894
R249 plus.n39 plus.n25 0.189894
R250 plus.n33 plus.n25 0.189894
R251 plus.n33 plus.n32 0.189894
R252 plus.n32 plus.n27 0.189894
R253 drain_left.n5 drain_left.n3 59.2758
R254 drain_left.n2 drain_left.n0 59.2758
R255 drain_left.n9 drain_left.n7 59.2758
R256 drain_left.n5 drain_left.n4 58.7154
R257 drain_left.n2 drain_left.n1 58.7154
R258 drain_left.n11 drain_left.n10 58.7154
R259 drain_left.n9 drain_left.n8 58.7154
R260 drain_left.n13 drain_left.n12 58.7153
R261 drain_left drain_left.n6 40.8578
R262 drain_left drain_left.n13 6.21356
R263 drain_left.n3 drain_left.t5 1.2005
R264 drain_left.n3 drain_left.t10 1.2005
R265 drain_left.n4 drain_left.t11 1.2005
R266 drain_left.n4 drain_left.t14 1.2005
R267 drain_left.n1 drain_left.t15 1.2005
R268 drain_left.n1 drain_left.t9 1.2005
R269 drain_left.n0 drain_left.t13 1.2005
R270 drain_left.n0 drain_left.t12 1.2005
R271 drain_left.n12 drain_left.t4 1.2005
R272 drain_left.n12 drain_left.t8 1.2005
R273 drain_left.n10 drain_left.t0 1.2005
R274 drain_left.n10 drain_left.t2 1.2005
R275 drain_left.n8 drain_left.t3 1.2005
R276 drain_left.n8 drain_left.t6 1.2005
R277 drain_left.n7 drain_left.t7 1.2005
R278 drain_left.n7 drain_left.t1 1.2005
R279 drain_left.n11 drain_left.n9 0.560845
R280 drain_left.n13 drain_left.n11 0.560845
R281 drain_left.n6 drain_left.n5 0.225326
R282 drain_left.n6 drain_left.n2 0.225326
C0 drain_left source 61.7512f
C1 drain_right drain_left 0.96779f
C2 drain_right source 61.7515f
C3 plus drain_left 6.99884f
C4 plus source 5.718359f
C5 drain_right plus 0.337321f
C6 minus drain_left 0.170952f
C7 minus source 5.704319f
C8 drain_right minus 6.81525f
C9 plus minus 7.89976f
C10 drain_right a_n1886_n5888# 8.48391f
C11 drain_left a_n1886_n5888# 8.76537f
C12 source a_n1886_n5888# 15.797586f
C13 minus a_n1886_n5888# 7.843384f
C14 plus a_n1886_n5888# 10.928731f
C15 drain_left.t13 a_n1886_n5888# 0.846411f
C16 drain_left.t12 a_n1886_n5888# 0.846411f
C17 drain_left.n0 a_n1886_n5888# 5.72729f
C18 drain_left.t15 a_n1886_n5888# 0.846411f
C19 drain_left.t9 a_n1886_n5888# 0.846411f
C20 drain_left.n1 a_n1886_n5888# 5.72395f
C21 drain_left.n2 a_n1886_n5888# 0.662668f
C22 drain_left.t5 a_n1886_n5888# 0.846411f
C23 drain_left.t10 a_n1886_n5888# 0.846411f
C24 drain_left.n3 a_n1886_n5888# 5.72729f
C25 drain_left.t11 a_n1886_n5888# 0.846411f
C26 drain_left.t14 a_n1886_n5888# 0.846411f
C27 drain_left.n4 a_n1886_n5888# 5.72395f
C28 drain_left.n5 a_n1886_n5888# 0.662668f
C29 drain_left.n6 a_n1886_n5888# 2.32498f
C30 drain_left.t7 a_n1886_n5888# 0.846411f
C31 drain_left.t1 a_n1886_n5888# 0.846411f
C32 drain_left.n7 a_n1886_n5888# 5.72729f
C33 drain_left.t3 a_n1886_n5888# 0.846411f
C34 drain_left.t6 a_n1886_n5888# 0.846411f
C35 drain_left.n8 a_n1886_n5888# 5.72395f
C36 drain_left.n9 a_n1886_n5888# 0.69032f
C37 drain_left.t0 a_n1886_n5888# 0.846411f
C38 drain_left.t2 a_n1886_n5888# 0.846411f
C39 drain_left.n10 a_n1886_n5888# 5.72395f
C40 drain_left.n11 a_n1886_n5888# 0.341132f
C41 drain_left.t4 a_n1886_n5888# 0.846411f
C42 drain_left.t8 a_n1886_n5888# 0.846411f
C43 drain_left.n12 a_n1886_n5888# 5.72394f
C44 drain_left.n13 a_n1886_n5888# 0.577286f
C45 plus.n0 a_n1886_n5888# 0.055405f
C46 plus.t11 a_n1886_n5888# 0.584594f
C47 plus.t13 a_n1886_n5888# 0.584594f
C48 plus.n1 a_n1886_n5888# 0.221261f
C49 plus.n2 a_n1886_n5888# 0.055405f
C50 plus.t15 a_n1886_n5888# 0.584594f
C51 plus.t9 a_n1886_n5888# 0.584594f
C52 plus.t12 a_n1886_n5888# 0.584594f
C53 plus.n3 a_n1886_n5888# 0.221261f
C54 plus.n4 a_n1886_n5888# 0.117569f
C55 plus.t14 a_n1886_n5888# 0.584594f
C56 plus.t8 a_n1886_n5888# 0.586654f
C57 plus.n5 a_n1886_n5888# 0.240216f
C58 plus.n6 a_n1886_n5888# 0.221261f
C59 plus.n7 a_n1886_n5888# 0.02265f
C60 plus.n8 a_n1886_n5888# 0.019234f
C61 plus.n9 a_n1886_n5888# 0.055405f
C62 plus.n10 a_n1886_n5888# 0.055405f
C63 plus.n11 a_n1886_n5888# 0.023504f
C64 plus.n12 a_n1886_n5888# 0.221261f
C65 plus.n13 a_n1886_n5888# 0.023504f
C66 plus.n14 a_n1886_n5888# 0.221261f
C67 plus.n15 a_n1886_n5888# 0.023504f
C68 plus.n16 a_n1886_n5888# 0.055405f
C69 plus.n17 a_n1886_n5888# 0.055405f
C70 plus.n18 a_n1886_n5888# 0.019234f
C71 plus.n19 a_n1886_n5888# 0.02265f
C72 plus.n20 a_n1886_n5888# 0.221261f
C73 plus.t7 a_n1886_n5888# 0.586654f
C74 plus.n21 a_n1886_n5888# 0.240143f
C75 plus.n22 a_n1886_n5888# 0.989547f
C76 plus.n23 a_n1886_n5888# 0.055405f
C77 plus.t2 a_n1886_n5888# 0.586654f
C78 plus.t3 a_n1886_n5888# 0.584594f
C79 plus.t0 a_n1886_n5888# 0.584594f
C80 plus.n24 a_n1886_n5888# 0.221261f
C81 plus.n25 a_n1886_n5888# 0.055405f
C82 plus.t6 a_n1886_n5888# 0.584594f
C83 plus.t4 a_n1886_n5888# 0.584594f
C84 plus.t1 a_n1886_n5888# 0.584594f
C85 plus.n26 a_n1886_n5888# 0.221261f
C86 plus.n27 a_n1886_n5888# 0.117569f
C87 plus.t10 a_n1886_n5888# 0.584594f
C88 plus.t5 a_n1886_n5888# 0.586654f
C89 plus.n28 a_n1886_n5888# 0.240216f
C90 plus.n29 a_n1886_n5888# 0.221261f
C91 plus.n30 a_n1886_n5888# 0.02265f
C92 plus.n31 a_n1886_n5888# 0.019234f
C93 plus.n32 a_n1886_n5888# 0.055405f
C94 plus.n33 a_n1886_n5888# 0.055405f
C95 plus.n34 a_n1886_n5888# 0.023504f
C96 plus.n35 a_n1886_n5888# 0.221261f
C97 plus.n36 a_n1886_n5888# 0.023504f
C98 plus.n37 a_n1886_n5888# 0.221261f
C99 plus.n38 a_n1886_n5888# 0.023504f
C100 plus.n39 a_n1886_n5888# 0.055405f
C101 plus.n40 a_n1886_n5888# 0.055405f
C102 plus.n41 a_n1886_n5888# 0.019234f
C103 plus.n42 a_n1886_n5888# 0.02265f
C104 plus.n43 a_n1886_n5888# 0.221261f
C105 plus.n44 a_n1886_n5888# 0.240143f
C106 plus.n45 a_n1886_n5888# 2.15118f
C107 drain_right.t13 a_n1886_n5888# 0.84531f
C108 drain_right.t5 a_n1886_n5888# 0.84531f
C109 drain_right.n0 a_n1886_n5888# 5.71983f
C110 drain_right.t1 a_n1886_n5888# 0.84531f
C111 drain_right.t15 a_n1886_n5888# 0.84531f
C112 drain_right.n1 a_n1886_n5888# 5.7165f
C113 drain_right.n2 a_n1886_n5888# 0.661806f
C114 drain_right.t0 a_n1886_n5888# 0.84531f
C115 drain_right.t14 a_n1886_n5888# 0.84531f
C116 drain_right.n3 a_n1886_n5888# 5.71983f
C117 drain_right.t9 a_n1886_n5888# 0.84531f
C118 drain_right.t2 a_n1886_n5888# 0.84531f
C119 drain_right.n4 a_n1886_n5888# 5.7165f
C120 drain_right.n5 a_n1886_n5888# 0.661806f
C121 drain_right.n6 a_n1886_n5888# 2.26345f
C122 drain_right.t12 a_n1886_n5888# 0.84531f
C123 drain_right.t11 a_n1886_n5888# 0.84531f
C124 drain_right.n7 a_n1886_n5888# 5.71982f
C125 drain_right.t8 a_n1886_n5888# 0.84531f
C126 drain_right.t7 a_n1886_n5888# 0.84531f
C127 drain_right.n8 a_n1886_n5888# 5.7165f
C128 drain_right.n9 a_n1886_n5888# 0.689434f
C129 drain_right.t3 a_n1886_n5888# 0.84531f
C130 drain_right.t10 a_n1886_n5888# 0.84531f
C131 drain_right.n10 a_n1886_n5888# 5.7165f
C132 drain_right.n11 a_n1886_n5888# 0.340688f
C133 drain_right.t4 a_n1886_n5888# 0.84531f
C134 drain_right.t6 a_n1886_n5888# 0.84531f
C135 drain_right.n12 a_n1886_n5888# 5.7165f
C136 drain_right.n13 a_n1886_n5888# 0.576522f
C137 source.t15 a_n1886_n5888# 5.76071f
C138 source.n0 a_n1886_n5888# 2.20432f
C139 source.t5 a_n1886_n5888# 0.698589f
C140 source.t8 a_n1886_n5888# 0.698589f
C141 source.n1 a_n1886_n5888# 4.64777f
C142 source.n2 a_n1886_n5888# 0.326344f
C143 source.t14 a_n1886_n5888# 0.698589f
C144 source.t6 a_n1886_n5888# 0.698589f
C145 source.n3 a_n1886_n5888# 4.64777f
C146 source.n4 a_n1886_n5888# 0.326344f
C147 source.t12 a_n1886_n5888# 0.698589f
C148 source.t10 a_n1886_n5888# 0.698589f
C149 source.n5 a_n1886_n5888# 4.64777f
C150 source.n6 a_n1886_n5888# 0.326344f
C151 source.t2 a_n1886_n5888# 5.76073f
C152 source.n7 a_n1886_n5888# 0.464045f
C153 source.t28 a_n1886_n5888# 5.76073f
C154 source.n8 a_n1886_n5888# 0.464045f
C155 source.t31 a_n1886_n5888# 0.698589f
C156 source.t21 a_n1886_n5888# 0.698589f
C157 source.n9 a_n1886_n5888# 4.64777f
C158 source.n10 a_n1886_n5888# 0.326344f
C159 source.t30 a_n1886_n5888# 0.698589f
C160 source.t24 a_n1886_n5888# 0.698589f
C161 source.n11 a_n1886_n5888# 4.64777f
C162 source.n12 a_n1886_n5888# 0.326344f
C163 source.t27 a_n1886_n5888# 0.698589f
C164 source.t26 a_n1886_n5888# 0.698589f
C165 source.n13 a_n1886_n5888# 4.64777f
C166 source.n14 a_n1886_n5888# 0.326344f
C167 source.t20 a_n1886_n5888# 5.76073f
C168 source.n15 a_n1886_n5888# 2.63664f
C169 source.t9 a_n1886_n5888# 5.76071f
C170 source.n16 a_n1886_n5888# 2.63666f
C171 source.t0 a_n1886_n5888# 0.698589f
C172 source.t3 a_n1886_n5888# 0.698589f
C173 source.n17 a_n1886_n5888# 4.64777f
C174 source.n18 a_n1886_n5888# 0.326345f
C175 source.t11 a_n1886_n5888# 0.698589f
C176 source.t13 a_n1886_n5888# 0.698589f
C177 source.n19 a_n1886_n5888# 4.64777f
C178 source.n20 a_n1886_n5888# 0.326345f
C179 source.t7 a_n1886_n5888# 0.698589f
C180 source.t4 a_n1886_n5888# 0.698589f
C181 source.n21 a_n1886_n5888# 4.64777f
C182 source.n22 a_n1886_n5888# 0.326345f
C183 source.t1 a_n1886_n5888# 5.76071f
C184 source.n23 a_n1886_n5888# 0.46406f
C185 source.t16 a_n1886_n5888# 5.76071f
C186 source.n24 a_n1886_n5888# 0.46406f
C187 source.t17 a_n1886_n5888# 0.698589f
C188 source.t19 a_n1886_n5888# 0.698589f
C189 source.n25 a_n1886_n5888# 4.64777f
C190 source.n26 a_n1886_n5888# 0.326345f
C191 source.t25 a_n1886_n5888# 0.698589f
C192 source.t18 a_n1886_n5888# 0.698589f
C193 source.n27 a_n1886_n5888# 4.64777f
C194 source.n28 a_n1886_n5888# 0.326345f
C195 source.t29 a_n1886_n5888# 0.698589f
C196 source.t22 a_n1886_n5888# 0.698589f
C197 source.n29 a_n1886_n5888# 4.64777f
C198 source.n30 a_n1886_n5888# 0.326345f
C199 source.t23 a_n1886_n5888# 5.76071f
C200 source.n31 a_n1886_n5888# 0.596841f
C201 source.n32 a_n1886_n5888# 2.48876f
C202 minus.n0 a_n1886_n5888# 0.05457f
C203 minus.t11 a_n1886_n5888# 0.577815f
C204 minus.t9 a_n1886_n5888# 0.575787f
C205 minus.t12 a_n1886_n5888# 0.575787f
C206 minus.n1 a_n1886_n5888# 0.217927f
C207 minus.n2 a_n1886_n5888# 0.05457f
C208 minus.t5 a_n1886_n5888# 0.575787f
C209 minus.t7 a_n1886_n5888# 0.575787f
C210 minus.t8 a_n1886_n5888# 0.575787f
C211 minus.n3 a_n1886_n5888# 0.217927f
C212 minus.n4 a_n1886_n5888# 0.115798f
C213 minus.t3 a_n1886_n5888# 0.575787f
C214 minus.t4 a_n1886_n5888# 0.577815f
C215 minus.n5 a_n1886_n5888# 0.236597f
C216 minus.n6 a_n1886_n5888# 0.217927f
C217 minus.n7 a_n1886_n5888# 0.022308f
C218 minus.n8 a_n1886_n5888# 0.018944f
C219 minus.n9 a_n1886_n5888# 0.05457f
C220 minus.n10 a_n1886_n5888# 0.05457f
C221 minus.n11 a_n1886_n5888# 0.023149f
C222 minus.n12 a_n1886_n5888# 0.217927f
C223 minus.n13 a_n1886_n5888# 0.023149f
C224 minus.n14 a_n1886_n5888# 0.217927f
C225 minus.n15 a_n1886_n5888# 0.023149f
C226 minus.n16 a_n1886_n5888# 0.05457f
C227 minus.n17 a_n1886_n5888# 0.05457f
C228 minus.n18 a_n1886_n5888# 0.018944f
C229 minus.n19 a_n1886_n5888# 0.022308f
C230 minus.n20 a_n1886_n5888# 0.217927f
C231 minus.n21 a_n1886_n5888# 0.236525f
C232 minus.n22 a_n1886_n5888# 2.76728f
C233 minus.n23 a_n1886_n5888# 0.05457f
C234 minus.t15 a_n1886_n5888# 0.575787f
C235 minus.t13 a_n1886_n5888# 0.575787f
C236 minus.n24 a_n1886_n5888# 0.217927f
C237 minus.n25 a_n1886_n5888# 0.05457f
C238 minus.t6 a_n1886_n5888# 0.575787f
C239 minus.t0 a_n1886_n5888# 0.575787f
C240 minus.t14 a_n1886_n5888# 0.575787f
C241 minus.n26 a_n1886_n5888# 0.217927f
C242 minus.n27 a_n1886_n5888# 0.115798f
C243 minus.t10 a_n1886_n5888# 0.575787f
C244 minus.t2 a_n1886_n5888# 0.577815f
C245 minus.n28 a_n1886_n5888# 0.236597f
C246 minus.n29 a_n1886_n5888# 0.217927f
C247 minus.n30 a_n1886_n5888# 0.022308f
C248 minus.n31 a_n1886_n5888# 0.018944f
C249 minus.n32 a_n1886_n5888# 0.05457f
C250 minus.n33 a_n1886_n5888# 0.05457f
C251 minus.n34 a_n1886_n5888# 0.023149f
C252 minus.n35 a_n1886_n5888# 0.217927f
C253 minus.n36 a_n1886_n5888# 0.023149f
C254 minus.n37 a_n1886_n5888# 0.217927f
C255 minus.n38 a_n1886_n5888# 0.023149f
C256 minus.n39 a_n1886_n5888# 0.05457f
C257 minus.n40 a_n1886_n5888# 0.05457f
C258 minus.n41 a_n1886_n5888# 0.018944f
C259 minus.n42 a_n1886_n5888# 0.022308f
C260 minus.n43 a_n1886_n5888# 0.217927f
C261 minus.t1 a_n1886_n5888# 0.577815f
C262 minus.n44 a_n1886_n5888# 0.236525f
C263 minus.n45 a_n1886_n5888# 0.357318f
C264 minus.n46 a_n1886_n5888# 3.26714f
.ends

