* NGSPICE file created from diffpair406.ext - technology: sky130A

.subckt diffpair406 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t16 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X1 source.t2 plus.t0 drain_left.t13 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X2 a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X3 drain_left.t12 plus.t1 source.t6 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X4 a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X5 a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X6 drain_left.t11 plus.t2 source.t8 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X7 source.t1 plus.t3 drain_left.t10 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X8 drain_right.t12 minus.t1 source.t15 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X9 a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X10 drain_left.t9 plus.t4 source.t0 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X11 source.t27 minus.t2 drain_right.t11 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X12 drain_left.t8 plus.t5 source.t11 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 drain_right.t10 minus.t3 source.t24 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X14 drain_right.t9 minus.t4 source.t23 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X15 source.t25 minus.t5 drain_right.t8 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X16 source.t26 minus.t6 drain_right.t7 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 source.t18 minus.t7 drain_right.t6 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X18 source.t7 plus.t6 drain_left.t7 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 drain_left.t6 plus.t7 source.t10 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X20 drain_right.t5 minus.t8 source.t17 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X21 drain_right.t4 minus.t9 source.t20 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X22 source.t4 plus.t8 drain_left.t5 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X23 source.t19 minus.t10 drain_right.t3 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X24 drain_right.t2 minus.t11 source.t14 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X25 drain_left.t4 plus.t9 source.t12 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X26 drain_left.t3 plus.t10 source.t13 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X27 drain_right.t1 minus.t12 source.t21 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X28 source.t3 plus.t11 drain_left.t2 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X29 source.t9 plus.t12 drain_left.t1 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X30 drain_left.t0 plus.t13 source.t5 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X31 source.t22 minus.t13 drain_right.t0 a_n1756_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
R0 minus.n15 minus.t9 2202.59
R1 minus.n3 minus.t3 2202.59
R2 minus.n32 minus.t12 2202.59
R3 minus.n20 minus.t0 2202.59
R4 minus.n1 minus.t6 2136.87
R5 minus.n14 minus.t10 2136.87
R6 minus.n12 minus.t4 2136.87
R7 minus.n6 minus.t8 2136.87
R8 minus.n4 minus.t2 2136.87
R9 minus.n18 minus.t13 2136.87
R10 minus.n31 minus.t7 2136.87
R11 minus.n29 minus.t1 2136.87
R12 minus.n23 minus.t11 2136.87
R13 minus.n21 minus.t5 2136.87
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 51.1217
R33 minus.n6 minus.n5 51.1217
R34 minus.n23 minus.n22 51.1217
R35 minus.n30 minus.n29 51.1217
R36 minus.n14 minus.n13 43.8187
R37 minus.n5 minus.n4 43.8187
R38 minus.n22 minus.n21 43.8187
R39 minus.n31 minus.n30 43.8187
R40 minus.n34 minus.n16 35.8433
R41 minus.n15 minus.n14 29.2126
R42 minus.n4 minus.n3 29.2126
R43 minus.n21 minus.n20 29.2126
R44 minus.n32 minus.n31 29.2126
R45 minus.n12 minus.n11 21.9096
R46 minus.n7 minus.n6 21.9096
R47 minus.n24 minus.n23 21.9096
R48 minus.n29 minus.n28 21.9096
R49 minus.n34 minus.n33 6.57058
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 source.n7 source.t24 45.3739
R62 source.n27 source.t21 45.3737
R63 source.n20 source.t0 45.3737
R64 source.n0 source.t12 45.3737
R65 source.n2 source.n1 42.8739
R66 source.n4 source.n3 42.8739
R67 source.n6 source.n5 42.8739
R68 source.n9 source.n8 42.8739
R69 source.n11 source.n10 42.8739
R70 source.n13 source.n12 42.8739
R71 source.n26 source.n25 42.8737
R72 source.n24 source.n23 42.8737
R73 source.n22 source.n21 42.8737
R74 source.n19 source.n18 42.8737
R75 source.n17 source.n16 42.8737
R76 source.n15 source.n14 42.8737
R77 source.n15 source.n13 22.4084
R78 source.n28 source.n0 16.305
R79 source.n28 source.n27 5.5436
R80 source.n25 source.t15 2.5005
R81 source.n25 source.t18 2.5005
R82 source.n23 source.t14 2.5005
R83 source.n23 source.t22 2.5005
R84 source.n21 source.t16 2.5005
R85 source.n21 source.t25 2.5005
R86 source.n18 source.t6 2.5005
R87 source.n18 source.t7 2.5005
R88 source.n16 source.t11 2.5005
R89 source.n16 source.t1 2.5005
R90 source.n14 source.t8 2.5005
R91 source.n14 source.t2 2.5005
R92 source.n1 source.t5 2.5005
R93 source.n1 source.t3 2.5005
R94 source.n3 source.t13 2.5005
R95 source.n3 source.t4 2.5005
R96 source.n5 source.t10 2.5005
R97 source.n5 source.t9 2.5005
R98 source.n8 source.t17 2.5005
R99 source.n8 source.t27 2.5005
R100 source.n10 source.t23 2.5005
R101 source.n10 source.t26 2.5005
R102 source.n12 source.t20 2.5005
R103 source.n12 source.t19 2.5005
R104 source.n7 source.n6 0.7505
R105 source.n22 source.n20 0.7505
R106 source.n13 source.n11 0.560845
R107 source.n11 source.n9 0.560845
R108 source.n9 source.n7 0.560845
R109 source.n6 source.n4 0.560845
R110 source.n4 source.n2 0.560845
R111 source.n2 source.n0 0.560845
R112 source.n17 source.n15 0.560845
R113 source.n19 source.n17 0.560845
R114 source.n20 source.n19 0.560845
R115 source.n24 source.n22 0.560845
R116 source.n26 source.n24 0.560845
R117 source.n27 source.n26 0.560845
R118 source source.n28 0.188
R119 drain_right.n1 drain_right.t13 62.6128
R120 drain_right.n11 drain_right.t4 62.0527
R121 drain_right.n4 drain_right.n2 60.1128
R122 drain_right.n8 drain_right.n6 60.1128
R123 drain_right.n8 drain_right.n7 59.5527
R124 drain_right.n10 drain_right.n9 59.5527
R125 drain_right.n4 drain_right.n3 59.5525
R126 drain_right.n1 drain_right.n0 59.5525
R127 drain_right drain_right.n5 30.0358
R128 drain_right drain_right.n11 5.93339
R129 drain_right.n2 drain_right.t6 2.5005
R130 drain_right.n2 drain_right.t1 2.5005
R131 drain_right.n3 drain_right.t0 2.5005
R132 drain_right.n3 drain_right.t12 2.5005
R133 drain_right.n0 drain_right.t8 2.5005
R134 drain_right.n0 drain_right.t2 2.5005
R135 drain_right.n6 drain_right.t11 2.5005
R136 drain_right.n6 drain_right.t10 2.5005
R137 drain_right.n7 drain_right.t7 2.5005
R138 drain_right.n7 drain_right.t5 2.5005
R139 drain_right.n9 drain_right.t3 2.5005
R140 drain_right.n9 drain_right.t9 2.5005
R141 drain_right.n11 drain_right.n10 0.560845
R142 drain_right.n10 drain_right.n8 0.560845
R143 drain_right.n5 drain_right.n1 0.365413
R144 drain_right.n5 drain_right.n4 0.0852402
R145 plus.n3 plus.t7 2202.59
R146 plus.n15 plus.t9 2202.59
R147 plus.n20 plus.t4 2202.59
R148 plus.n32 plus.t2 2202.59
R149 plus.n1 plus.t8 2136.87
R150 plus.n4 plus.t12 2136.87
R151 plus.n6 plus.t10 2136.87
R152 plus.n12 plus.t13 2136.87
R153 plus.n14 plus.t11 2136.87
R154 plus.n18 plus.t3 2136.87
R155 plus.n21 plus.t6 2136.87
R156 plus.n23 plus.t1 2136.87
R157 plus.n29 plus.t5 2136.87
R158 plus.n31 plus.t0 2136.87
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 51.1217
R178 plus.n13 plus.n12 51.1217
R179 plus.n30 plus.n29 51.1217
R180 plus.n23 plus.n22 51.1217
R181 plus.n5 plus.n4 43.8187
R182 plus.n14 plus.n13 43.8187
R183 plus.n31 plus.n30 43.8187
R184 plus.n22 plus.n21 43.8187
R185 plus plus.n33 29.7244
R186 plus.n4 plus.n3 29.2126
R187 plus.n15 plus.n14 29.2126
R188 plus.n32 plus.n31 29.2126
R189 plus.n21 plus.n20 29.2126
R190 plus.n7 plus.n6 21.9096
R191 plus.n12 plus.n11 21.9096
R192 plus.n29 plus.n28 21.9096
R193 plus.n24 plus.n23 21.9096
R194 plus plus.n16 12.2145
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t6 62.613
R206 drain_left.n1 drain_left.t11 62.6128
R207 drain_left.n4 drain_left.n2 60.1128
R208 drain_left.n9 drain_left.n8 59.5527
R209 drain_left.n7 drain_left.n6 59.5527
R210 drain_left.n4 drain_left.n3 59.5525
R211 drain_left.n1 drain_left.n0 59.5525
R212 drain_left.n11 drain_left.n10 59.5525
R213 drain_left drain_left.n5 30.5891
R214 drain_left drain_left.n11 6.21356
R215 drain_left.n2 drain_left.t7 2.5005
R216 drain_left.n2 drain_left.t9 2.5005
R217 drain_left.n3 drain_left.t10 2.5005
R218 drain_left.n3 drain_left.t12 2.5005
R219 drain_left.n0 drain_left.t13 2.5005
R220 drain_left.n0 drain_left.t8 2.5005
R221 drain_left.n10 drain_left.t2 2.5005
R222 drain_left.n10 drain_left.t4 2.5005
R223 drain_left.n8 drain_left.t5 2.5005
R224 drain_left.n8 drain_left.t0 2.5005
R225 drain_left.n6 drain_left.t1 2.5005
R226 drain_left.n6 drain_left.t3 2.5005
R227 drain_left.n9 drain_left.n7 0.560845
R228 drain_left.n11 drain_left.n9 0.560845
R229 drain_left.n5 drain_left.n1 0.365413
R230 drain_left.n5 drain_left.n4 0.0852402
C0 source drain_left 28.586098f
C1 drain_right minus 3.19515f
C2 drain_right plus 0.326127f
C3 plus minus 5.32397f
C4 drain_right drain_left 0.901368f
C5 drain_right source 28.575802f
C6 minus drain_left 0.171187f
C7 plus drain_left 3.36241f
C8 minus source 2.69676f
C9 plus source 2.71145f
C10 drain_right a_n1756_n3288# 6.9784f
C11 drain_left a_n1756_n3288# 7.25394f
C12 source a_n1756_n3288# 6.268777f
C13 minus a_n1756_n3288# 6.459813f
C14 plus a_n1756_n3288# 8.619491f
C15 drain_left.t11 a_n1756_n3288# 3.032f
C16 drain_left.t13 a_n1756_n3288# 0.375899f
C17 drain_left.t8 a_n1756_n3288# 0.375899f
C18 drain_left.n0 a_n1756_n3288# 2.46326f
C19 drain_left.n1 a_n1756_n3288# 0.684459f
C20 drain_left.t7 a_n1756_n3288# 0.375899f
C21 drain_left.t9 a_n1756_n3288# 0.375899f
C22 drain_left.n2 a_n1756_n3288# 2.46628f
C23 drain_left.t10 a_n1756_n3288# 0.375899f
C24 drain_left.t12 a_n1756_n3288# 0.375899f
C25 drain_left.n3 a_n1756_n3288# 2.46326f
C26 drain_left.n4 a_n1756_n3288# 0.602669f
C27 drain_left.n5 a_n1756_n3288# 1.25471f
C28 drain_left.t6 a_n1756_n3288# 3.03201f
C29 drain_left.t1 a_n1756_n3288# 0.375899f
C30 drain_left.t3 a_n1756_n3288# 0.375899f
C31 drain_left.n6 a_n1756_n3288# 2.46327f
C32 drain_left.n7 a_n1756_n3288# 0.699254f
C33 drain_left.t5 a_n1756_n3288# 0.375899f
C34 drain_left.t0 a_n1756_n3288# 0.375899f
C35 drain_left.n8 a_n1756_n3288# 2.46327f
C36 drain_left.n9 a_n1756_n3288# 0.314038f
C37 drain_left.t2 a_n1756_n3288# 0.375899f
C38 drain_left.t4 a_n1756_n3288# 0.375899f
C39 drain_left.n10 a_n1756_n3288# 2.46326f
C40 drain_left.n11 a_n1756_n3288# 0.532532f
C41 plus.n0 a_n1756_n3288# 0.056205f
C42 plus.t11 a_n1756_n3288# 0.285887f
C43 plus.t13 a_n1756_n3288# 0.285887f
C44 plus.t8 a_n1756_n3288# 0.285887f
C45 plus.n1 a_n1756_n3288# 0.140718f
C46 plus.n2 a_n1756_n3288# 0.131382f
C47 plus.t10 a_n1756_n3288# 0.285887f
C48 plus.t12 a_n1756_n3288# 0.285887f
C49 plus.t7 a_n1756_n3288# 0.289634f
C50 plus.n3 a_n1756_n3288# 0.145724f
C51 plus.n4 a_n1756_n3288# 0.122073f
C52 plus.n5 a_n1756_n3288# 0.023843f
C53 plus.n6 a_n1756_n3288# 0.122073f
C54 plus.n7 a_n1756_n3288# 0.023843f
C55 plus.n8 a_n1756_n3288# 0.056205f
C56 plus.n9 a_n1756_n3288# 0.056205f
C57 plus.n10 a_n1756_n3288# 0.056205f
C58 plus.n11 a_n1756_n3288# 0.023843f
C59 plus.n12 a_n1756_n3288# 0.122073f
C60 plus.n13 a_n1756_n3288# 0.023843f
C61 plus.n14 a_n1756_n3288# 0.122073f
C62 plus.t9 a_n1756_n3288# 0.289634f
C63 plus.n15 a_n1756_n3288# 0.145635f
C64 plus.n16 a_n1756_n3288# 0.638319f
C65 plus.n17 a_n1756_n3288# 0.056205f
C66 plus.t2 a_n1756_n3288# 0.289634f
C67 plus.t0 a_n1756_n3288# 0.285887f
C68 plus.t5 a_n1756_n3288# 0.285887f
C69 plus.t3 a_n1756_n3288# 0.285887f
C70 plus.n18 a_n1756_n3288# 0.140718f
C71 plus.n19 a_n1756_n3288# 0.131382f
C72 plus.t1 a_n1756_n3288# 0.285887f
C73 plus.t6 a_n1756_n3288# 0.285887f
C74 plus.t4 a_n1756_n3288# 0.289634f
C75 plus.n20 a_n1756_n3288# 0.145724f
C76 plus.n21 a_n1756_n3288# 0.122073f
C77 plus.n22 a_n1756_n3288# 0.023843f
C78 plus.n23 a_n1756_n3288# 0.122073f
C79 plus.n24 a_n1756_n3288# 0.023843f
C80 plus.n25 a_n1756_n3288# 0.056205f
C81 plus.n26 a_n1756_n3288# 0.056205f
C82 plus.n27 a_n1756_n3288# 0.056205f
C83 plus.n28 a_n1756_n3288# 0.023843f
C84 plus.n29 a_n1756_n3288# 0.122073f
C85 plus.n30 a_n1756_n3288# 0.023843f
C86 plus.n31 a_n1756_n3288# 0.122073f
C87 plus.n32 a_n1756_n3288# 0.145635f
C88 plus.n33 a_n1756_n3288# 1.65698f
C89 drain_right.t13 a_n1756_n3288# 3.02272f
C90 drain_right.t8 a_n1756_n3288# 0.374748f
C91 drain_right.t2 a_n1756_n3288# 0.374748f
C92 drain_right.n0 a_n1756_n3288# 2.45572f
C93 drain_right.n1 a_n1756_n3288# 0.682363f
C94 drain_right.t6 a_n1756_n3288# 0.374748f
C95 drain_right.t1 a_n1756_n3288# 0.374748f
C96 drain_right.n2 a_n1756_n3288# 2.45873f
C97 drain_right.t0 a_n1756_n3288# 0.374748f
C98 drain_right.t12 a_n1756_n3288# 0.374748f
C99 drain_right.n3 a_n1756_n3288# 2.45572f
C100 drain_right.n4 a_n1756_n3288# 0.600824f
C101 drain_right.n5 a_n1756_n3288# 1.19669f
C102 drain_right.t11 a_n1756_n3288# 0.374748f
C103 drain_right.t10 a_n1756_n3288# 0.374748f
C104 drain_right.n6 a_n1756_n3288# 2.45873f
C105 drain_right.t7 a_n1756_n3288# 0.374748f
C106 drain_right.t5 a_n1756_n3288# 0.374748f
C107 drain_right.n7 a_n1756_n3288# 2.45573f
C108 drain_right.n8 a_n1756_n3288# 0.633651f
C109 drain_right.t3 a_n1756_n3288# 0.374748f
C110 drain_right.t9 a_n1756_n3288# 0.374748f
C111 drain_right.n9 a_n1756_n3288# 2.45573f
C112 drain_right.n10 a_n1756_n3288# 0.313076f
C113 drain_right.t4 a_n1756_n3288# 3.01926f
C114 drain_right.n11 a_n1756_n3288# 0.606214f
C115 source.t12 a_n1756_n3288# 2.97387f
C116 source.n0 a_n1756_n3288# 1.48305f
C117 source.t5 a_n1756_n3288# 0.384321f
C118 source.t3 a_n1756_n3288# 0.384321f
C119 source.n1 a_n1756_n3288# 2.43311f
C120 source.n2 a_n1756_n3288# 0.370064f
C121 source.t13 a_n1756_n3288# 0.384321f
C122 source.t4 a_n1756_n3288# 0.384321f
C123 source.n3 a_n1756_n3288# 2.43311f
C124 source.n4 a_n1756_n3288# 0.370064f
C125 source.t10 a_n1756_n3288# 0.384321f
C126 source.t9 a_n1756_n3288# 0.384321f
C127 source.n5 a_n1756_n3288# 2.43311f
C128 source.n6 a_n1756_n3288# 0.38641f
C129 source.t24 a_n1756_n3288# 2.97388f
C130 source.n7 a_n1756_n3288# 0.537411f
C131 source.t17 a_n1756_n3288# 0.384321f
C132 source.t27 a_n1756_n3288# 0.384321f
C133 source.n8 a_n1756_n3288# 2.43311f
C134 source.n9 a_n1756_n3288# 0.370064f
C135 source.t23 a_n1756_n3288# 0.384321f
C136 source.t26 a_n1756_n3288# 0.384321f
C137 source.n10 a_n1756_n3288# 2.43311f
C138 source.n11 a_n1756_n3288# 0.370064f
C139 source.t20 a_n1756_n3288# 0.384321f
C140 source.t19 a_n1756_n3288# 0.384321f
C141 source.n12 a_n1756_n3288# 2.43311f
C142 source.n13 a_n1756_n3288# 1.80147f
C143 source.t8 a_n1756_n3288# 0.384321f
C144 source.t2 a_n1756_n3288# 0.384321f
C145 source.n14 a_n1756_n3288# 2.43309f
C146 source.n15 a_n1756_n3288# 1.80148f
C147 source.t11 a_n1756_n3288# 0.384321f
C148 source.t1 a_n1756_n3288# 0.384321f
C149 source.n16 a_n1756_n3288# 2.43309f
C150 source.n17 a_n1756_n3288# 0.370077f
C151 source.t6 a_n1756_n3288# 0.384321f
C152 source.t7 a_n1756_n3288# 0.384321f
C153 source.n18 a_n1756_n3288# 2.43309f
C154 source.n19 a_n1756_n3288# 0.370077f
C155 source.t0 a_n1756_n3288# 2.97387f
C156 source.n20 a_n1756_n3288# 0.537424f
C157 source.t16 a_n1756_n3288# 0.384321f
C158 source.t25 a_n1756_n3288# 0.384321f
C159 source.n21 a_n1756_n3288# 2.43309f
C160 source.n22 a_n1756_n3288# 0.386424f
C161 source.t14 a_n1756_n3288# 0.384321f
C162 source.t22 a_n1756_n3288# 0.384321f
C163 source.n23 a_n1756_n3288# 2.43309f
C164 source.n24 a_n1756_n3288# 0.370077f
C165 source.t15 a_n1756_n3288# 0.384321f
C166 source.t18 a_n1756_n3288# 0.384321f
C167 source.n25 a_n1756_n3288# 2.43309f
C168 source.n26 a_n1756_n3288# 0.370077f
C169 source.t21 a_n1756_n3288# 2.97387f
C170 source.n27 a_n1756_n3288# 0.665459f
C171 source.n28 a_n1756_n3288# 1.67889f
C172 minus.n0 a_n1756_n3288# 0.054674f
C173 minus.t9 a_n1756_n3288# 0.281743f
C174 minus.t10 a_n1756_n3288# 0.278099f
C175 minus.t4 a_n1756_n3288# 0.278099f
C176 minus.t6 a_n1756_n3288# 0.278099f
C177 minus.n1 a_n1756_n3288# 0.136885f
C178 minus.n2 a_n1756_n3288# 0.127802f
C179 minus.t8 a_n1756_n3288# 0.278099f
C180 minus.t2 a_n1756_n3288# 0.278099f
C181 minus.t3 a_n1756_n3288# 0.281743f
C182 minus.n3 a_n1756_n3288# 0.141754f
C183 minus.n4 a_n1756_n3288# 0.118748f
C184 minus.n5 a_n1756_n3288# 0.023194f
C185 minus.n6 a_n1756_n3288# 0.118748f
C186 minus.n7 a_n1756_n3288# 0.023194f
C187 minus.n8 a_n1756_n3288# 0.054674f
C188 minus.n9 a_n1756_n3288# 0.054674f
C189 minus.n10 a_n1756_n3288# 0.054674f
C190 minus.n11 a_n1756_n3288# 0.023194f
C191 minus.n12 a_n1756_n3288# 0.118748f
C192 minus.n13 a_n1756_n3288# 0.023194f
C193 minus.n14 a_n1756_n3288# 0.118748f
C194 minus.n15 a_n1756_n3288# 0.141668f
C195 minus.n16 a_n1756_n3288# 1.90601f
C196 minus.n17 a_n1756_n3288# 0.054674f
C197 minus.t7 a_n1756_n3288# 0.278099f
C198 minus.t1 a_n1756_n3288# 0.278099f
C199 minus.t13 a_n1756_n3288# 0.278099f
C200 minus.n18 a_n1756_n3288# 0.136885f
C201 minus.n19 a_n1756_n3288# 0.127802f
C202 minus.t11 a_n1756_n3288# 0.278099f
C203 minus.t5 a_n1756_n3288# 0.278099f
C204 minus.t0 a_n1756_n3288# 0.281743f
C205 minus.n20 a_n1756_n3288# 0.141754f
C206 minus.n21 a_n1756_n3288# 0.118748f
C207 minus.n22 a_n1756_n3288# 0.023194f
C208 minus.n23 a_n1756_n3288# 0.118748f
C209 minus.n24 a_n1756_n3288# 0.023194f
C210 minus.n25 a_n1756_n3288# 0.054674f
C211 minus.n26 a_n1756_n3288# 0.054674f
C212 minus.n27 a_n1756_n3288# 0.054674f
C213 minus.n28 a_n1756_n3288# 0.023194f
C214 minus.n29 a_n1756_n3288# 0.118748f
C215 minus.n30 a_n1756_n3288# 0.023194f
C216 minus.n31 a_n1756_n3288# 0.118748f
C217 minus.t12 a_n1756_n3288# 0.281743f
C218 minus.n32 a_n1756_n3288# 0.141668f
C219 minus.n33 a_n1756_n3288# 0.366506f
C220 minus.n34 a_n1756_n3288# 2.31447f
.ends

