* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t33 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 drain_left.t18 plus.t1 source.t24 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X2 source.t7 minus.t0 drain_right.t19 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 drain_left.t17 plus.t2 source.t32 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X4 source.t6 minus.t1 drain_right.t18 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X5 drain_left.t16 plus.t3 source.t31 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X6 source.t12 minus.t2 drain_right.t17 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X7 a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X8 source.t5 minus.t3 drain_right.t16 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X9 source.t4 minus.t4 drain_right.t15 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X10 source.t3 minus.t5 drain_right.t14 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X11 source.t15 plus.t4 drain_left.t15 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X12 a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X13 drain_right.t13 minus.t6 source.t11 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X14 source.t9 minus.t7 drain_right.t12 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X15 source.t8 minus.t8 drain_right.t11 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X16 source.t10 minus.t9 drain_right.t10 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X17 drain_right.t9 minus.t10 source.t2 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X18 drain_right.t8 minus.t11 source.t1 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X19 source.t0 minus.t12 drain_right.t7 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X20 source.t22 plus.t5 drain_left.t14 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X21 source.t17 plus.t6 drain_left.t13 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X22 source.t16 plus.t7 drain_left.t12 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X23 source.t18 plus.t8 drain_left.t11 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X24 drain_left.t10 plus.t9 source.t23 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X25 drain_left.t9 plus.t10 source.t28 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X26 drain_right.t6 minus.t13 source.t36 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X27 drain_left.t8 plus.t11 source.t19 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X28 source.t26 plus.t12 drain_left.t7 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X29 drain_right.t5 minus.t14 source.t39 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X30 drain_left.t6 plus.t13 source.t27 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X31 a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X32 source.t20 plus.t14 drain_left.t5 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X33 a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X34 source.t25 plus.t15 drain_left.t4 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X35 source.t21 plus.t16 drain_left.t3 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X36 drain_right.t4 minus.t15 source.t37 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X37 drain_right.t3 minus.t16 source.t35 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X38 source.t34 plus.t17 drain_left.t2 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X39 drain_right.t2 minus.t17 source.t14 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X40 drain_right.t1 minus.t18 source.t13 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X41 drain_left.t1 plus.t18 source.t30 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X42 drain_left.t0 plus.t19 source.t29 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X43 drain_right.t0 minus.t19 source.t38 a_n1992_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
R0 plus.n6 plus.t4 274.303
R1 plus.n25 plus.t2 274.303
R2 plus.n33 plus.t10 274.303
R3 plus.n52 plus.t17 274.303
R4 plus.n5 plus.t1 221.72
R5 plus.n9 plus.t8 221.72
R6 plus.n11 plus.t0 221.72
R7 plus.n3 plus.t7 221.72
R8 plus.n17 plus.t18 221.72
R9 plus.n1 plus.t6 221.72
R10 plus.n22 plus.t3 221.72
R11 plus.n24 plus.t12 221.72
R12 plus.n32 plus.t5 221.72
R13 plus.n36 plus.t13 221.72
R14 plus.n38 plus.t16 221.72
R15 plus.n30 plus.t9 221.72
R16 plus.n44 plus.t14 221.72
R17 plus.n28 plus.t11 221.72
R18 plus.n49 plus.t15 221.72
R19 plus.n51 plus.t19 221.72
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus.n10 plus.n9 29.2126
R63 plus.n22 plus.n21 29.2126
R64 plus.n49 plus.n48 29.2126
R65 plus.n37 plus.n36 29.2126
R66 plus plus.n53 26.3778
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 7.97398
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n0 source.t32 243.255
R93 source.n9 source.t15 243.255
R94 source.n10 source.t39 243.255
R95 source.n19 source.t0 243.255
R96 source.n39 source.t2 243.254
R97 source.n30 source.t3 243.254
R98 source.n29 source.t28 243.254
R99 source.n20 source.t34 243.254
R100 source.n2 source.n1 223.454
R101 source.n4 source.n3 223.454
R102 source.n6 source.n5 223.454
R103 source.n8 source.n7 223.454
R104 source.n12 source.n11 223.454
R105 source.n14 source.n13 223.454
R106 source.n16 source.n15 223.454
R107 source.n18 source.n17 223.454
R108 source.n38 source.n37 223.453
R109 source.n36 source.n35 223.453
R110 source.n34 source.n33 223.453
R111 source.n32 source.n31 223.453
R112 source.n28 source.n27 223.453
R113 source.n26 source.n25 223.453
R114 source.n24 source.n23 223.453
R115 source.n22 source.n21 223.453
R116 source.n37 source.t11 19.8005
R117 source.n37 source.t5 19.8005
R118 source.n35 source.t1 19.8005
R119 source.n35 source.t9 19.8005
R120 source.n33 source.t38 19.8005
R121 source.n33 source.t4 19.8005
R122 source.n31 source.t13 19.8005
R123 source.n31 source.t7 19.8005
R124 source.n27 source.t27 19.8005
R125 source.n27 source.t22 19.8005
R126 source.n25 source.t23 19.8005
R127 source.n25 source.t21 19.8005
R128 source.n23 source.t19 19.8005
R129 source.n23 source.t20 19.8005
R130 source.n21 source.t29 19.8005
R131 source.n21 source.t25 19.8005
R132 source.n1 source.t31 19.8005
R133 source.n1 source.t26 19.8005
R134 source.n3 source.t30 19.8005
R135 source.n3 source.t17 19.8005
R136 source.n5 source.t33 19.8005
R137 source.n5 source.t16 19.8005
R138 source.n7 source.t24 19.8005
R139 source.n7 source.t18 19.8005
R140 source.n11 source.t36 19.8005
R141 source.n11 source.t12 19.8005
R142 source.n13 source.t37 19.8005
R143 source.n13 source.t6 19.8005
R144 source.n15 source.t35 19.8005
R145 source.n15 source.t10 19.8005
R146 source.n17 source.t14 19.8005
R147 source.n17 source.t8 19.8005
R148 source.n20 source.n19 13.4544
R149 source.n40 source.n0 7.94146
R150 source.n40 source.n39 5.51343
R151 source.n19 source.n18 0.5005
R152 source.n18 source.n16 0.5005
R153 source.n16 source.n14 0.5005
R154 source.n14 source.n12 0.5005
R155 source.n12 source.n10 0.5005
R156 source.n9 source.n8 0.5005
R157 source.n8 source.n6 0.5005
R158 source.n6 source.n4 0.5005
R159 source.n4 source.n2 0.5005
R160 source.n2 source.n0 0.5005
R161 source.n22 source.n20 0.5005
R162 source.n24 source.n22 0.5005
R163 source.n26 source.n24 0.5005
R164 source.n28 source.n26 0.5005
R165 source.n29 source.n28 0.5005
R166 source.n32 source.n30 0.5005
R167 source.n34 source.n32 0.5005
R168 source.n36 source.n34 0.5005
R169 source.n38 source.n36 0.5005
R170 source.n39 source.n38 0.5005
R171 source.n10 source.n9 0.470328
R172 source.n30 source.n29 0.470328
R173 source source.n40 0.188
R174 drain_left.n10 drain_left.n8 240.632
R175 drain_left.n6 drain_left.n4 240.631
R176 drain_left.n2 drain_left.n0 240.631
R177 drain_left.n16 drain_left.n15 240.132
R178 drain_left.n14 drain_left.n13 240.132
R179 drain_left.n12 drain_left.n11 240.132
R180 drain_left.n10 drain_left.n9 240.132
R181 drain_left.n7 drain_left.n3 240.131
R182 drain_left.n6 drain_left.n5 240.131
R183 drain_left.n2 drain_left.n1 240.131
R184 drain_left drain_left.n7 23.0337
R185 drain_left.n3 drain_left.t5 19.8005
R186 drain_left.n3 drain_left.t10 19.8005
R187 drain_left.n4 drain_left.t14 19.8005
R188 drain_left.n4 drain_left.t9 19.8005
R189 drain_left.n5 drain_left.t3 19.8005
R190 drain_left.n5 drain_left.t6 19.8005
R191 drain_left.n1 drain_left.t4 19.8005
R192 drain_left.n1 drain_left.t8 19.8005
R193 drain_left.n0 drain_left.t2 19.8005
R194 drain_left.n0 drain_left.t0 19.8005
R195 drain_left.n15 drain_left.t7 19.8005
R196 drain_left.n15 drain_left.t17 19.8005
R197 drain_left.n13 drain_left.t13 19.8005
R198 drain_left.n13 drain_left.t16 19.8005
R199 drain_left.n11 drain_left.t12 19.8005
R200 drain_left.n11 drain_left.t1 19.8005
R201 drain_left.n9 drain_left.t11 19.8005
R202 drain_left.n9 drain_left.t19 19.8005
R203 drain_left.n8 drain_left.t15 19.8005
R204 drain_left.n8 drain_left.t18 19.8005
R205 drain_left drain_left.n16 6.15322
R206 drain_left.n12 drain_left.n10 0.5005
R207 drain_left.n14 drain_left.n12 0.5005
R208 drain_left.n16 drain_left.n14 0.5005
R209 drain_left.n7 drain_left.n6 0.445154
R210 drain_left.n7 drain_left.n2 0.445154
R211 minus.n25 minus.t12 274.303
R212 minus.n6 minus.t14 274.303
R213 minus.n52 minus.t10 274.303
R214 minus.n33 minus.t5 274.303
R215 minus.n24 minus.t17 221.72
R216 minus.n22 minus.t8 221.72
R217 minus.n1 minus.t16 221.72
R218 minus.n17 minus.t9 221.72
R219 minus.n3 minus.t15 221.72
R220 minus.n11 minus.t1 221.72
R221 minus.n9 minus.t13 221.72
R222 minus.n5 minus.t2 221.72
R223 minus.n51 minus.t3 221.72
R224 minus.n49 minus.t6 221.72
R225 minus.n28 minus.t7 221.72
R226 minus.n44 minus.t11 221.72
R227 minus.n30 minus.t4 221.72
R228 minus.n38 minus.t19 221.72
R229 minus.n36 minus.t0 221.72
R230 minus.n32 minus.t18 221.72
R231 minus.n7 minus.n6 161.489
R232 minus.n34 minus.n33 161.489
R233 minus.n26 minus.n25 161.3
R234 minus.n23 minus.n0 161.3
R235 minus.n21 minus.n20 161.3
R236 minus.n19 minus.n18 161.3
R237 minus.n16 minus.n2 161.3
R238 minus.n15 minus.n14 161.3
R239 minus.n13 minus.n12 161.3
R240 minus.n10 minus.n4 161.3
R241 minus.n8 minus.n7 161.3
R242 minus.n53 minus.n52 161.3
R243 minus.n50 minus.n27 161.3
R244 minus.n48 minus.n47 161.3
R245 minus.n46 minus.n45 161.3
R246 minus.n43 minus.n29 161.3
R247 minus.n42 minus.n41 161.3
R248 minus.n40 minus.n39 161.3
R249 minus.n37 minus.n31 161.3
R250 minus.n35 minus.n34 161.3
R251 minus.n16 minus.n15 73.0308
R252 minus.n43 minus.n42 73.0308
R253 minus.n18 minus.n17 67.1884
R254 minus.n12 minus.n3 67.1884
R255 minus.n39 minus.n30 67.1884
R256 minus.n45 minus.n44 67.1884
R257 minus.n21 minus.n1 55.5035
R258 minus.n11 minus.n10 55.5035
R259 minus.n38 minus.n37 55.5035
R260 minus.n48 minus.n28 55.5035
R261 minus.n23 minus.n22 43.8187
R262 minus.n9 minus.n8 43.8187
R263 minus.n36 minus.n35 43.8187
R264 minus.n50 minus.n49 43.8187
R265 minus.n24 minus.n23 40.8975
R266 minus.n8 minus.n5 40.8975
R267 minus.n35 minus.n32 40.8975
R268 minus.n51 minus.n50 40.8975
R269 minus.n25 minus.n24 32.1338
R270 minus.n6 minus.n5 32.1338
R271 minus.n33 minus.n32 32.1338
R272 minus.n52 minus.n51 32.1338
R273 minus.n22 minus.n21 29.2126
R274 minus.n10 minus.n9 29.2126
R275 minus.n37 minus.n36 29.2126
R276 minus.n49 minus.n48 29.2126
R277 minus.n54 minus.n26 28.33
R278 minus.n18 minus.n1 17.5278
R279 minus.n12 minus.n11 17.5278
R280 minus.n39 minus.n38 17.5278
R281 minus.n45 minus.n28 17.5278
R282 minus.n54 minus.n53 6.49671
R283 minus.n17 minus.n16 5.84292
R284 minus.n15 minus.n3 5.84292
R285 minus.n42 minus.n30 5.84292
R286 minus.n44 minus.n43 5.84292
R287 minus.n26 minus.n0 0.189894
R288 minus.n20 minus.n0 0.189894
R289 minus.n20 minus.n19 0.189894
R290 minus.n19 minus.n2 0.189894
R291 minus.n14 minus.n2 0.189894
R292 minus.n14 minus.n13 0.189894
R293 minus.n13 minus.n4 0.189894
R294 minus.n7 minus.n4 0.189894
R295 minus.n34 minus.n31 0.189894
R296 minus.n40 minus.n31 0.189894
R297 minus.n41 minus.n40 0.189894
R298 minus.n41 minus.n29 0.189894
R299 minus.n46 minus.n29 0.189894
R300 minus.n47 minus.n46 0.189894
R301 minus.n47 minus.n27 0.189894
R302 minus.n53 minus.n27 0.189894
R303 minus minus.n54 0.188
R304 drain_right.n10 drain_right.n8 240.632
R305 drain_right.n6 drain_right.n4 240.631
R306 drain_right.n2 drain_right.n0 240.631
R307 drain_right.n10 drain_right.n9 240.132
R308 drain_right.n12 drain_right.n11 240.132
R309 drain_right.n14 drain_right.n13 240.132
R310 drain_right.n16 drain_right.n15 240.132
R311 drain_right.n7 drain_right.n3 240.131
R312 drain_right.n6 drain_right.n5 240.131
R313 drain_right.n2 drain_right.n1 240.131
R314 drain_right drain_right.n7 22.4805
R315 drain_right.n3 drain_right.t15 19.8005
R316 drain_right.n3 drain_right.t8 19.8005
R317 drain_right.n4 drain_right.t16 19.8005
R318 drain_right.n4 drain_right.t9 19.8005
R319 drain_right.n5 drain_right.t12 19.8005
R320 drain_right.n5 drain_right.t13 19.8005
R321 drain_right.n1 drain_right.t19 19.8005
R322 drain_right.n1 drain_right.t0 19.8005
R323 drain_right.n0 drain_right.t14 19.8005
R324 drain_right.n0 drain_right.t1 19.8005
R325 drain_right.n8 drain_right.t17 19.8005
R326 drain_right.n8 drain_right.t5 19.8005
R327 drain_right.n9 drain_right.t18 19.8005
R328 drain_right.n9 drain_right.t6 19.8005
R329 drain_right.n11 drain_right.t10 19.8005
R330 drain_right.n11 drain_right.t4 19.8005
R331 drain_right.n13 drain_right.t11 19.8005
R332 drain_right.n13 drain_right.t3 19.8005
R333 drain_right.n15 drain_right.t7 19.8005
R334 drain_right.n15 drain_right.t2 19.8005
R335 drain_right drain_right.n16 6.15322
R336 drain_right.n16 drain_right.n14 0.5005
R337 drain_right.n14 drain_right.n12 0.5005
R338 drain_right.n12 drain_right.n10 0.5005
R339 drain_right.n7 drain_right.n6 0.445154
R340 drain_right.n7 drain_right.n2 0.445154
C0 drain_right source 6.37228f
C1 source plus 1.38523f
C2 source drain_left 6.37207f
C3 drain_right plus 0.357705f
C4 drain_right drain_left 1.04702f
C5 drain_left plus 1.25327f
C6 source minus 1.37137f
C7 drain_right minus 1.05885f
C8 minus plus 3.61084f
C9 drain_left minus 0.179068f
C10 drain_right a_n1992_n1088# 4.00608f
C11 drain_left a_n1992_n1088# 4.27615f
C12 source a_n1992_n1088# 2.607437f
C13 minus a_n1992_n1088# 6.872941f
C14 plus a_n1992_n1088# 7.547469f
C15 drain_right.t14 a_n1992_n1088# 0.02167f
C16 drain_right.t1 a_n1992_n1088# 0.02167f
C17 drain_right.n0 a_n1992_n1088# 0.08481f
C18 drain_right.t19 a_n1992_n1088# 0.02167f
C19 drain_right.t0 a_n1992_n1088# 0.02167f
C20 drain_right.n1 a_n1992_n1088# 0.084205f
C21 drain_right.n2 a_n1992_n1088# 0.56725f
C22 drain_right.t15 a_n1992_n1088# 0.02167f
C23 drain_right.t8 a_n1992_n1088# 0.02167f
C24 drain_right.n3 a_n1992_n1088# 0.084205f
C25 drain_right.t16 a_n1992_n1088# 0.02167f
C26 drain_right.t9 a_n1992_n1088# 0.02167f
C27 drain_right.n4 a_n1992_n1088# 0.08481f
C28 drain_right.t12 a_n1992_n1088# 0.02167f
C29 drain_right.t13 a_n1992_n1088# 0.02167f
C30 drain_right.n5 a_n1992_n1088# 0.084205f
C31 drain_right.n6 a_n1992_n1088# 0.56725f
C32 drain_right.n7 a_n1992_n1088# 0.959662f
C33 drain_right.t17 a_n1992_n1088# 0.02167f
C34 drain_right.t5 a_n1992_n1088# 0.02167f
C35 drain_right.n8 a_n1992_n1088# 0.08481f
C36 drain_right.t18 a_n1992_n1088# 0.02167f
C37 drain_right.t6 a_n1992_n1088# 0.02167f
C38 drain_right.n9 a_n1992_n1088# 0.084205f
C39 drain_right.n10 a_n1992_n1088# 0.570711f
C40 drain_right.t10 a_n1992_n1088# 0.02167f
C41 drain_right.t4 a_n1992_n1088# 0.02167f
C42 drain_right.n11 a_n1992_n1088# 0.084205f
C43 drain_right.n12 a_n1992_n1088# 0.280135f
C44 drain_right.t11 a_n1992_n1088# 0.02167f
C45 drain_right.t3 a_n1992_n1088# 0.02167f
C46 drain_right.n13 a_n1992_n1088# 0.084205f
C47 drain_right.n14 a_n1992_n1088# 0.280135f
C48 drain_right.t7 a_n1992_n1088# 0.02167f
C49 drain_right.t2 a_n1992_n1088# 0.02167f
C50 drain_right.n15 a_n1992_n1088# 0.084205f
C51 drain_right.n16 a_n1992_n1088# 0.506494f
C52 minus.n0 a_n1992_n1088# 0.030367f
C53 minus.t12 a_n1992_n1088# 0.028719f
C54 minus.t17 a_n1992_n1088# 0.023403f
C55 minus.t8 a_n1992_n1088# 0.023403f
C56 minus.t16 a_n1992_n1088# 0.023403f
C57 minus.n1 a_n1992_n1088# 0.025672f
C58 minus.n2 a_n1992_n1088# 0.030367f
C59 minus.t9 a_n1992_n1088# 0.023403f
C60 minus.t15 a_n1992_n1088# 0.023403f
C61 minus.n3 a_n1992_n1088# 0.025672f
C62 minus.n4 a_n1992_n1088# 0.030367f
C63 minus.t1 a_n1992_n1088# 0.023403f
C64 minus.t13 a_n1992_n1088# 0.023403f
C65 minus.t2 a_n1992_n1088# 0.023403f
C66 minus.n5 a_n1992_n1088# 0.025672f
C67 minus.t14 a_n1992_n1088# 0.028719f
C68 minus.n6 a_n1992_n1088# 0.034033f
C69 minus.n7 a_n1992_n1088# 0.069488f
C70 minus.n8 a_n1992_n1088# 0.011571f
C71 minus.n9 a_n1992_n1088# 0.025672f
C72 minus.n10 a_n1992_n1088# 0.011571f
C73 minus.n11 a_n1992_n1088# 0.025672f
C74 minus.n12 a_n1992_n1088# 0.011571f
C75 minus.n13 a_n1992_n1088# 0.030367f
C76 minus.n14 a_n1992_n1088# 0.030367f
C77 minus.n15 a_n1992_n1088# 0.010823f
C78 minus.n16 a_n1992_n1088# 0.010823f
C79 minus.n17 a_n1992_n1088# 0.025672f
C80 minus.n18 a_n1992_n1088# 0.011571f
C81 minus.n19 a_n1992_n1088# 0.030367f
C82 minus.n20 a_n1992_n1088# 0.030367f
C83 minus.n21 a_n1992_n1088# 0.011571f
C84 minus.n22 a_n1992_n1088# 0.025672f
C85 minus.n23 a_n1992_n1088# 0.011571f
C86 minus.n24 a_n1992_n1088# 0.025672f
C87 minus.n25 a_n1992_n1088# 0.033987f
C88 minus.n26 a_n1992_n1088# 0.715225f
C89 minus.n27 a_n1992_n1088# 0.030367f
C90 minus.t3 a_n1992_n1088# 0.023403f
C91 minus.t6 a_n1992_n1088# 0.023403f
C92 minus.t7 a_n1992_n1088# 0.023403f
C93 minus.n28 a_n1992_n1088# 0.025672f
C94 minus.n29 a_n1992_n1088# 0.030367f
C95 minus.t11 a_n1992_n1088# 0.023403f
C96 minus.t4 a_n1992_n1088# 0.023403f
C97 minus.n30 a_n1992_n1088# 0.025672f
C98 minus.n31 a_n1992_n1088# 0.030367f
C99 minus.t19 a_n1992_n1088# 0.023403f
C100 minus.t0 a_n1992_n1088# 0.023403f
C101 minus.t18 a_n1992_n1088# 0.023403f
C102 minus.n32 a_n1992_n1088# 0.025672f
C103 minus.t5 a_n1992_n1088# 0.028719f
C104 minus.n33 a_n1992_n1088# 0.034033f
C105 minus.n34 a_n1992_n1088# 0.069488f
C106 minus.n35 a_n1992_n1088# 0.011571f
C107 minus.n36 a_n1992_n1088# 0.025672f
C108 minus.n37 a_n1992_n1088# 0.011571f
C109 minus.n38 a_n1992_n1088# 0.025672f
C110 minus.n39 a_n1992_n1088# 0.011571f
C111 minus.n40 a_n1992_n1088# 0.030367f
C112 minus.n41 a_n1992_n1088# 0.030367f
C113 minus.n42 a_n1992_n1088# 0.010823f
C114 minus.n43 a_n1992_n1088# 0.010823f
C115 minus.n44 a_n1992_n1088# 0.025672f
C116 minus.n45 a_n1992_n1088# 0.011571f
C117 minus.n46 a_n1992_n1088# 0.030367f
C118 minus.n47 a_n1992_n1088# 0.030367f
C119 minus.n48 a_n1992_n1088# 0.011571f
C120 minus.n49 a_n1992_n1088# 0.025672f
C121 minus.n50 a_n1992_n1088# 0.011571f
C122 minus.n51 a_n1992_n1088# 0.025672f
C123 minus.t10 a_n1992_n1088# 0.028719f
C124 minus.n52 a_n1992_n1088# 0.033987f
C125 minus.n53 a_n1992_n1088# 0.198296f
C126 minus.n54 a_n1992_n1088# 0.884147f
C127 drain_left.t2 a_n1992_n1088# 0.021313f
C128 drain_left.t0 a_n1992_n1088# 0.021313f
C129 drain_left.n0 a_n1992_n1088# 0.083412f
C130 drain_left.t4 a_n1992_n1088# 0.021313f
C131 drain_left.t8 a_n1992_n1088# 0.021313f
C132 drain_left.n1 a_n1992_n1088# 0.082817f
C133 drain_left.n2 a_n1992_n1088# 0.557899f
C134 drain_left.t5 a_n1992_n1088# 0.021313f
C135 drain_left.t10 a_n1992_n1088# 0.021313f
C136 drain_left.n3 a_n1992_n1088# 0.082817f
C137 drain_left.t14 a_n1992_n1088# 0.021313f
C138 drain_left.t9 a_n1992_n1088# 0.021313f
C139 drain_left.n4 a_n1992_n1088# 0.083412f
C140 drain_left.t3 a_n1992_n1088# 0.021313f
C141 drain_left.t6 a_n1992_n1088# 0.021313f
C142 drain_left.n5 a_n1992_n1088# 0.082817f
C143 drain_left.n6 a_n1992_n1088# 0.557899f
C144 drain_left.n7 a_n1992_n1088# 0.995915f
C145 drain_left.t15 a_n1992_n1088# 0.021313f
C146 drain_left.t18 a_n1992_n1088# 0.021313f
C147 drain_left.n8 a_n1992_n1088# 0.083412f
C148 drain_left.t11 a_n1992_n1088# 0.021313f
C149 drain_left.t19 a_n1992_n1088# 0.021313f
C150 drain_left.n9 a_n1992_n1088# 0.082817f
C151 drain_left.n10 a_n1992_n1088# 0.561302f
C152 drain_left.t12 a_n1992_n1088# 0.021313f
C153 drain_left.t1 a_n1992_n1088# 0.021313f
C154 drain_left.n11 a_n1992_n1088# 0.082817f
C155 drain_left.n12 a_n1992_n1088# 0.275517f
C156 drain_left.t13 a_n1992_n1088# 0.021313f
C157 drain_left.t16 a_n1992_n1088# 0.021313f
C158 drain_left.n13 a_n1992_n1088# 0.082817f
C159 drain_left.n14 a_n1992_n1088# 0.275517f
C160 drain_left.t7 a_n1992_n1088# 0.021313f
C161 drain_left.t17 a_n1992_n1088# 0.021313f
C162 drain_left.n15 a_n1992_n1088# 0.082817f
C163 drain_left.n16 a_n1992_n1088# 0.498144f
C164 source.t32 a_n1992_n1088# 0.141267f
C165 source.n0 a_n1992_n1088# 0.59858f
C166 source.t31 a_n1992_n1088# 0.025381f
C167 source.t26 a_n1992_n1088# 0.025381f
C168 source.n1 a_n1992_n1088# 0.082314f
C169 source.n2 a_n1992_n1088# 0.300753f
C170 source.t30 a_n1992_n1088# 0.025381f
C171 source.t17 a_n1992_n1088# 0.025381f
C172 source.n3 a_n1992_n1088# 0.082314f
C173 source.n4 a_n1992_n1088# 0.300753f
C174 source.t33 a_n1992_n1088# 0.025381f
C175 source.t16 a_n1992_n1088# 0.025381f
C176 source.n5 a_n1992_n1088# 0.082314f
C177 source.n6 a_n1992_n1088# 0.300753f
C178 source.t24 a_n1992_n1088# 0.025381f
C179 source.t18 a_n1992_n1088# 0.025381f
C180 source.n7 a_n1992_n1088# 0.082314f
C181 source.n8 a_n1992_n1088# 0.300753f
C182 source.t15 a_n1992_n1088# 0.141267f
C183 source.n9 a_n1992_n1088# 0.307899f
C184 source.t39 a_n1992_n1088# 0.141267f
C185 source.n10 a_n1992_n1088# 0.307899f
C186 source.t36 a_n1992_n1088# 0.025381f
C187 source.t12 a_n1992_n1088# 0.025381f
C188 source.n11 a_n1992_n1088# 0.082314f
C189 source.n12 a_n1992_n1088# 0.300753f
C190 source.t37 a_n1992_n1088# 0.025381f
C191 source.t6 a_n1992_n1088# 0.025381f
C192 source.n13 a_n1992_n1088# 0.082314f
C193 source.n14 a_n1992_n1088# 0.300753f
C194 source.t35 a_n1992_n1088# 0.025381f
C195 source.t10 a_n1992_n1088# 0.025381f
C196 source.n15 a_n1992_n1088# 0.082314f
C197 source.n16 a_n1992_n1088# 0.300753f
C198 source.t14 a_n1992_n1088# 0.025381f
C199 source.t8 a_n1992_n1088# 0.025381f
C200 source.n17 a_n1992_n1088# 0.082314f
C201 source.n18 a_n1992_n1088# 0.300753f
C202 source.t0 a_n1992_n1088# 0.141267f
C203 source.n19 a_n1992_n1088# 0.85502f
C204 source.t34 a_n1992_n1088# 0.141267f
C205 source.n20 a_n1992_n1088# 0.855021f
C206 source.t29 a_n1992_n1088# 0.025381f
C207 source.t25 a_n1992_n1088# 0.025381f
C208 source.n21 a_n1992_n1088# 0.082314f
C209 source.n22 a_n1992_n1088# 0.300753f
C210 source.t19 a_n1992_n1088# 0.025381f
C211 source.t20 a_n1992_n1088# 0.025381f
C212 source.n23 a_n1992_n1088# 0.082314f
C213 source.n24 a_n1992_n1088# 0.300753f
C214 source.t23 a_n1992_n1088# 0.025381f
C215 source.t21 a_n1992_n1088# 0.025381f
C216 source.n25 a_n1992_n1088# 0.082314f
C217 source.n26 a_n1992_n1088# 0.300753f
C218 source.t27 a_n1992_n1088# 0.025381f
C219 source.t22 a_n1992_n1088# 0.025381f
C220 source.n27 a_n1992_n1088# 0.082314f
C221 source.n28 a_n1992_n1088# 0.300753f
C222 source.t28 a_n1992_n1088# 0.141267f
C223 source.n29 a_n1992_n1088# 0.307899f
C224 source.t3 a_n1992_n1088# 0.141267f
C225 source.n30 a_n1992_n1088# 0.307899f
C226 source.t13 a_n1992_n1088# 0.025381f
C227 source.t7 a_n1992_n1088# 0.025381f
C228 source.n31 a_n1992_n1088# 0.082314f
C229 source.n32 a_n1992_n1088# 0.300753f
C230 source.t38 a_n1992_n1088# 0.025381f
C231 source.t4 a_n1992_n1088# 0.025381f
C232 source.n33 a_n1992_n1088# 0.082314f
C233 source.n34 a_n1992_n1088# 0.300753f
C234 source.t1 a_n1992_n1088# 0.025381f
C235 source.t9 a_n1992_n1088# 0.025381f
C236 source.n35 a_n1992_n1088# 0.082314f
C237 source.n36 a_n1992_n1088# 0.300753f
C238 source.t11 a_n1992_n1088# 0.025381f
C239 source.t5 a_n1992_n1088# 0.025381f
C240 source.n37 a_n1992_n1088# 0.082314f
C241 source.n38 a_n1992_n1088# 0.300753f
C242 source.t2 a_n1992_n1088# 0.141267f
C243 source.n39 a_n1992_n1088# 0.485637f
C244 source.n40 a_n1992_n1088# 0.64867f
C245 plus.n0 a_n1992_n1088# 0.030894f
C246 plus.t12 a_n1992_n1088# 0.023809f
C247 plus.t3 a_n1992_n1088# 0.023809f
C248 plus.t6 a_n1992_n1088# 0.023809f
C249 plus.n1 a_n1992_n1088# 0.026118f
C250 plus.n2 a_n1992_n1088# 0.030894f
C251 plus.t18 a_n1992_n1088# 0.023809f
C252 plus.t7 a_n1992_n1088# 0.023809f
C253 plus.n3 a_n1992_n1088# 0.026118f
C254 plus.n4 a_n1992_n1088# 0.030894f
C255 plus.t0 a_n1992_n1088# 0.023809f
C256 plus.t8 a_n1992_n1088# 0.023809f
C257 plus.t1 a_n1992_n1088# 0.023809f
C258 plus.n5 a_n1992_n1088# 0.026118f
C259 plus.t4 a_n1992_n1088# 0.029218f
C260 plus.n6 a_n1992_n1088# 0.034624f
C261 plus.n7 a_n1992_n1088# 0.070693f
C262 plus.n8 a_n1992_n1088# 0.011772f
C263 plus.n9 a_n1992_n1088# 0.026118f
C264 plus.n10 a_n1992_n1088# 0.011772f
C265 plus.n11 a_n1992_n1088# 0.026118f
C266 plus.n12 a_n1992_n1088# 0.011772f
C267 plus.n13 a_n1992_n1088# 0.030894f
C268 plus.n14 a_n1992_n1088# 0.030894f
C269 plus.n15 a_n1992_n1088# 0.01101f
C270 plus.n16 a_n1992_n1088# 0.01101f
C271 plus.n17 a_n1992_n1088# 0.026118f
C272 plus.n18 a_n1992_n1088# 0.011772f
C273 plus.n19 a_n1992_n1088# 0.030894f
C274 plus.n20 a_n1992_n1088# 0.030894f
C275 plus.n21 a_n1992_n1088# 0.011772f
C276 plus.n22 a_n1992_n1088# 0.026118f
C277 plus.n23 a_n1992_n1088# 0.011772f
C278 plus.n24 a_n1992_n1088# 0.026118f
C279 plus.t2 a_n1992_n1088# 0.029218f
C280 plus.n25 a_n1992_n1088# 0.034577f
C281 plus.n26 a_n1992_n1088# 0.211556f
C282 plus.n27 a_n1992_n1088# 0.030894f
C283 plus.t17 a_n1992_n1088# 0.029218f
C284 plus.t19 a_n1992_n1088# 0.023809f
C285 plus.t15 a_n1992_n1088# 0.023809f
C286 plus.t11 a_n1992_n1088# 0.023809f
C287 plus.n28 a_n1992_n1088# 0.026118f
C288 plus.n29 a_n1992_n1088# 0.030894f
C289 plus.t14 a_n1992_n1088# 0.023809f
C290 plus.t9 a_n1992_n1088# 0.023809f
C291 plus.n30 a_n1992_n1088# 0.026118f
C292 plus.n31 a_n1992_n1088# 0.030894f
C293 plus.t16 a_n1992_n1088# 0.023809f
C294 plus.t13 a_n1992_n1088# 0.023809f
C295 plus.t5 a_n1992_n1088# 0.023809f
C296 plus.n32 a_n1992_n1088# 0.026118f
C297 plus.t10 a_n1992_n1088# 0.029218f
C298 plus.n33 a_n1992_n1088# 0.034624f
C299 plus.n34 a_n1992_n1088# 0.070693f
C300 plus.n35 a_n1992_n1088# 0.011772f
C301 plus.n36 a_n1992_n1088# 0.026118f
C302 plus.n37 a_n1992_n1088# 0.011772f
C303 plus.n38 a_n1992_n1088# 0.026118f
C304 plus.n39 a_n1992_n1088# 0.011772f
C305 plus.n40 a_n1992_n1088# 0.030894f
C306 plus.n41 a_n1992_n1088# 0.030894f
C307 plus.n42 a_n1992_n1088# 0.01101f
C308 plus.n43 a_n1992_n1088# 0.01101f
C309 plus.n44 a_n1992_n1088# 0.026118f
C310 plus.n45 a_n1992_n1088# 0.011772f
C311 plus.n46 a_n1992_n1088# 0.030894f
C312 plus.n47 a_n1992_n1088# 0.030894f
C313 plus.n48 a_n1992_n1088# 0.011772f
C314 plus.n49 a_n1992_n1088# 0.026118f
C315 plus.n50 a_n1992_n1088# 0.011772f
C316 plus.n51 a_n1992_n1088# 0.026118f
C317 plus.n52 a_n1992_n1088# 0.034577f
C318 plus.n53 a_n1992_n1088# 0.704592f
.ends

