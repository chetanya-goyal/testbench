* NGSPICE file created from diffpair590.ext - technology: sky130A

.subckt diffpair590 minus drain_right drain_left source plus
X0 a_n968_n4892# a_n968_n4892# a_n968_n4892# a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X1 drain_right minus source a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.3
X2 a_n968_n4892# a_n968_n4892# a_n968_n4892# a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X3 a_n968_n4892# a_n968_n4892# a_n968_n4892# a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X4 drain_left plus source a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.3
X5 drain_right minus source a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.3
X6 drain_left plus source a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.3
X7 a_n968_n4892# a_n968_n4892# a_n968_n4892# a_n968_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
.ends

