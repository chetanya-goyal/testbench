* NGSPICE file created from diffpair302.ext - technology: sky130A

.subckt diffpair302 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t6 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X1 source.t3 minus.t0 drain_right.t5 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X2 drain_left.t4 plus.t1 source.t10 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X3 a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X4 a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X5 drain_left.t3 plus.t2 source.t7 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X6 drain_left.t2 plus.t3 source.t9 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X7 drain_right.t4 minus.t1 source.t2 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X8 a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X9 drain_right.t3 minus.t2 source.t1 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X10 source.t8 plus.t4 drain_left.t1 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X11 drain_right.t2 minus.t3 source.t0 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X12 source.t11 plus.t5 drain_left.t0 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 drain_right.t1 minus.t4 source.t5 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X14 source.t4 minus.t5 drain_right.t0 a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# a_n1540_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
R0 plus.n1 plus.t1 284.284
R1 plus.n7 plus.t3 284.284
R2 plus.n4 plus.t0 262.69
R3 plus.n2 plus.t5 262.69
R4 plus.n10 plus.t2 262.69
R5 plus.n8 plus.t4 262.69
R6 plus.n3 plus.n0 161.3
R7 plus.n5 plus.n4 161.3
R8 plus.n9 plus.n6 161.3
R9 plus.n11 plus.n10 161.3
R10 plus.n1 plus.n0 44.8545
R11 plus.n7 plus.n6 44.8545
R12 plus plus.n11 26.6903
R13 plus.n4 plus.n3 26.2914
R14 plus.n10 plus.n9 26.2914
R15 plus.n3 plus.n2 21.9096
R16 plus.n9 plus.n8 21.9096
R17 plus.n2 plus.n1 20.3348
R18 plus.n8 plus.n7 20.3348
R19 plus plus.n5 9.99861
R20 plus.n5 plus.n0 0.189894
R21 plus.n11 plus.n6 0.189894
R22 source.n130 source.n104 289.615
R23 source.n96 source.n70 289.615
R24 source.n26 source.n0 289.615
R25 source.n60 source.n34 289.615
R26 source.n115 source.n114 185
R27 source.n112 source.n111 185
R28 source.n121 source.n120 185
R29 source.n123 source.n122 185
R30 source.n108 source.n107 185
R31 source.n129 source.n128 185
R32 source.n131 source.n130 185
R33 source.n81 source.n80 185
R34 source.n78 source.n77 185
R35 source.n87 source.n86 185
R36 source.n89 source.n88 185
R37 source.n74 source.n73 185
R38 source.n95 source.n94 185
R39 source.n97 source.n96 185
R40 source.n27 source.n26 185
R41 source.n25 source.n24 185
R42 source.n4 source.n3 185
R43 source.n19 source.n18 185
R44 source.n17 source.n16 185
R45 source.n8 source.n7 185
R46 source.n11 source.n10 185
R47 source.n61 source.n60 185
R48 source.n59 source.n58 185
R49 source.n38 source.n37 185
R50 source.n53 source.n52 185
R51 source.n51 source.n50 185
R52 source.n42 source.n41 185
R53 source.n45 source.n44 185
R54 source.t1 source.n113 147.661
R55 source.t9 source.n79 147.661
R56 source.t6 source.n9 147.661
R57 source.t0 source.n43 147.661
R58 source.n114 source.n111 104.615
R59 source.n121 source.n111 104.615
R60 source.n122 source.n121 104.615
R61 source.n122 source.n107 104.615
R62 source.n129 source.n107 104.615
R63 source.n130 source.n129 104.615
R64 source.n80 source.n77 104.615
R65 source.n87 source.n77 104.615
R66 source.n88 source.n87 104.615
R67 source.n88 source.n73 104.615
R68 source.n95 source.n73 104.615
R69 source.n96 source.n95 104.615
R70 source.n26 source.n25 104.615
R71 source.n25 source.n3 104.615
R72 source.n18 source.n3 104.615
R73 source.n18 source.n17 104.615
R74 source.n17 source.n7 104.615
R75 source.n10 source.n7 104.615
R76 source.n60 source.n59 104.615
R77 source.n59 source.n37 104.615
R78 source.n52 source.n37 104.615
R79 source.n52 source.n51 104.615
R80 source.n51 source.n41 104.615
R81 source.n44 source.n41 104.615
R82 source.n114 source.t1 52.3082
R83 source.n80 source.t9 52.3082
R84 source.n10 source.t6 52.3082
R85 source.n44 source.t0 52.3082
R86 source.n33 source.n32 50.512
R87 source.n67 source.n66 50.512
R88 source.n103 source.n102 50.5119
R89 source.n69 source.n68 50.5119
R90 source.n135 source.n134 32.1853
R91 source.n101 source.n100 32.1853
R92 source.n31 source.n30 32.1853
R93 source.n65 source.n64 32.1853
R94 source.n69 source.n67 18.5181
R95 source.n115 source.n113 15.6674
R96 source.n81 source.n79 15.6674
R97 source.n11 source.n9 15.6674
R98 source.n45 source.n43 15.6674
R99 source.n116 source.n112 12.8005
R100 source.n82 source.n78 12.8005
R101 source.n12 source.n8 12.8005
R102 source.n46 source.n42 12.8005
R103 source.n120 source.n119 12.0247
R104 source.n86 source.n85 12.0247
R105 source.n16 source.n15 12.0247
R106 source.n50 source.n49 12.0247
R107 source.n136 source.n31 11.9233
R108 source.n123 source.n110 11.249
R109 source.n89 source.n76 11.249
R110 source.n19 source.n6 11.249
R111 source.n53 source.n40 11.249
R112 source.n124 source.n108 10.4732
R113 source.n90 source.n74 10.4732
R114 source.n20 source.n4 10.4732
R115 source.n54 source.n38 10.4732
R116 source.n128 source.n127 9.69747
R117 source.n94 source.n93 9.69747
R118 source.n24 source.n23 9.69747
R119 source.n58 source.n57 9.69747
R120 source.n134 source.n133 9.45567
R121 source.n100 source.n99 9.45567
R122 source.n30 source.n29 9.45567
R123 source.n64 source.n63 9.45567
R124 source.n133 source.n132 9.3005
R125 source.n106 source.n105 9.3005
R126 source.n127 source.n126 9.3005
R127 source.n125 source.n124 9.3005
R128 source.n110 source.n109 9.3005
R129 source.n119 source.n118 9.3005
R130 source.n117 source.n116 9.3005
R131 source.n99 source.n98 9.3005
R132 source.n72 source.n71 9.3005
R133 source.n93 source.n92 9.3005
R134 source.n91 source.n90 9.3005
R135 source.n76 source.n75 9.3005
R136 source.n85 source.n84 9.3005
R137 source.n83 source.n82 9.3005
R138 source.n29 source.n28 9.3005
R139 source.n2 source.n1 9.3005
R140 source.n23 source.n22 9.3005
R141 source.n21 source.n20 9.3005
R142 source.n6 source.n5 9.3005
R143 source.n15 source.n14 9.3005
R144 source.n13 source.n12 9.3005
R145 source.n63 source.n62 9.3005
R146 source.n36 source.n35 9.3005
R147 source.n57 source.n56 9.3005
R148 source.n55 source.n54 9.3005
R149 source.n40 source.n39 9.3005
R150 source.n49 source.n48 9.3005
R151 source.n47 source.n46 9.3005
R152 source.n131 source.n106 8.92171
R153 source.n97 source.n72 8.92171
R154 source.n27 source.n2 8.92171
R155 source.n61 source.n36 8.92171
R156 source.n132 source.n104 8.14595
R157 source.n98 source.n70 8.14595
R158 source.n28 source.n0 8.14595
R159 source.n62 source.n34 8.14595
R160 source.n134 source.n104 5.81868
R161 source.n100 source.n70 5.81868
R162 source.n30 source.n0 5.81868
R163 source.n64 source.n34 5.81868
R164 source.n136 source.n135 5.7074
R165 source.n132 source.n131 5.04292
R166 source.n98 source.n97 5.04292
R167 source.n28 source.n27 5.04292
R168 source.n62 source.n61 5.04292
R169 source.n117 source.n113 4.38594
R170 source.n83 source.n79 4.38594
R171 source.n13 source.n9 4.38594
R172 source.n47 source.n43 4.38594
R173 source.n128 source.n106 4.26717
R174 source.n94 source.n72 4.26717
R175 source.n24 source.n2 4.26717
R176 source.n58 source.n36 4.26717
R177 source.n127 source.n108 3.49141
R178 source.n93 source.n74 3.49141
R179 source.n23 source.n4 3.49141
R180 source.n57 source.n38 3.49141
R181 source.n102 source.t5 3.3005
R182 source.n102 source.t4 3.3005
R183 source.n68 source.t7 3.3005
R184 source.n68 source.t8 3.3005
R185 source.n32 source.t10 3.3005
R186 source.n32 source.t11 3.3005
R187 source.n66 source.t2 3.3005
R188 source.n66 source.t3 3.3005
R189 source.n124 source.n123 2.71565
R190 source.n90 source.n89 2.71565
R191 source.n20 source.n19 2.71565
R192 source.n54 source.n53 2.71565
R193 source.n120 source.n110 1.93989
R194 source.n86 source.n76 1.93989
R195 source.n16 source.n6 1.93989
R196 source.n50 source.n40 1.93989
R197 source.n119 source.n112 1.16414
R198 source.n85 source.n78 1.16414
R199 source.n15 source.n8 1.16414
R200 source.n49 source.n42 1.16414
R201 source.n65 source.n33 0.914293
R202 source.n103 source.n101 0.914293
R203 source.n67 source.n65 0.888431
R204 source.n33 source.n31 0.888431
R205 source.n101 source.n69 0.888431
R206 source.n135 source.n103 0.888431
R207 source.n116 source.n115 0.388379
R208 source.n82 source.n81 0.388379
R209 source.n12 source.n11 0.388379
R210 source.n46 source.n45 0.388379
R211 source source.n136 0.188
R212 source.n118 source.n117 0.155672
R213 source.n118 source.n109 0.155672
R214 source.n125 source.n109 0.155672
R215 source.n126 source.n125 0.155672
R216 source.n126 source.n105 0.155672
R217 source.n133 source.n105 0.155672
R218 source.n84 source.n83 0.155672
R219 source.n84 source.n75 0.155672
R220 source.n91 source.n75 0.155672
R221 source.n92 source.n91 0.155672
R222 source.n92 source.n71 0.155672
R223 source.n99 source.n71 0.155672
R224 source.n29 source.n1 0.155672
R225 source.n22 source.n1 0.155672
R226 source.n22 source.n21 0.155672
R227 source.n21 source.n5 0.155672
R228 source.n14 source.n5 0.155672
R229 source.n14 source.n13 0.155672
R230 source.n63 source.n35 0.155672
R231 source.n56 source.n35 0.155672
R232 source.n56 source.n55 0.155672
R233 source.n55 source.n39 0.155672
R234 source.n48 source.n39 0.155672
R235 source.n48 source.n47 0.155672
R236 drain_left.n26 drain_left.n0 289.615
R237 drain_left.n59 drain_left.n33 289.615
R238 drain_left.n11 drain_left.n10 185
R239 drain_left.n8 drain_left.n7 185
R240 drain_left.n17 drain_left.n16 185
R241 drain_left.n19 drain_left.n18 185
R242 drain_left.n4 drain_left.n3 185
R243 drain_left.n25 drain_left.n24 185
R244 drain_left.n27 drain_left.n26 185
R245 drain_left.n60 drain_left.n59 185
R246 drain_left.n58 drain_left.n57 185
R247 drain_left.n37 drain_left.n36 185
R248 drain_left.n52 drain_left.n51 185
R249 drain_left.n50 drain_left.n49 185
R250 drain_left.n41 drain_left.n40 185
R251 drain_left.n44 drain_left.n43 185
R252 drain_left.t3 drain_left.n9 147.661
R253 drain_left.t4 drain_left.n42 147.661
R254 drain_left.n10 drain_left.n7 104.615
R255 drain_left.n17 drain_left.n7 104.615
R256 drain_left.n18 drain_left.n17 104.615
R257 drain_left.n18 drain_left.n3 104.615
R258 drain_left.n25 drain_left.n3 104.615
R259 drain_left.n26 drain_left.n25 104.615
R260 drain_left.n59 drain_left.n58 104.615
R261 drain_left.n58 drain_left.n36 104.615
R262 drain_left.n51 drain_left.n36 104.615
R263 drain_left.n51 drain_left.n50 104.615
R264 drain_left.n50 drain_left.n40 104.615
R265 drain_left.n43 drain_left.n40 104.615
R266 drain_left.n32 drain_left.n31 67.3573
R267 drain_left.n65 drain_left.n64 67.1907
R268 drain_left.n10 drain_left.t3 52.3082
R269 drain_left.n43 drain_left.t4 52.3082
R270 drain_left.n65 drain_left.n63 49.7521
R271 drain_left.n32 drain_left.n30 49.4747
R272 drain_left drain_left.n32 25.2634
R273 drain_left.n11 drain_left.n9 15.6674
R274 drain_left.n44 drain_left.n42 15.6674
R275 drain_left.n12 drain_left.n8 12.8005
R276 drain_left.n45 drain_left.n41 12.8005
R277 drain_left.n16 drain_left.n15 12.0247
R278 drain_left.n49 drain_left.n48 12.0247
R279 drain_left.n19 drain_left.n6 11.249
R280 drain_left.n52 drain_left.n39 11.249
R281 drain_left.n20 drain_left.n4 10.4732
R282 drain_left.n53 drain_left.n37 10.4732
R283 drain_left.n24 drain_left.n23 9.69747
R284 drain_left.n57 drain_left.n56 9.69747
R285 drain_left.n30 drain_left.n29 9.45567
R286 drain_left.n63 drain_left.n62 9.45567
R287 drain_left.n29 drain_left.n28 9.3005
R288 drain_left.n2 drain_left.n1 9.3005
R289 drain_left.n23 drain_left.n22 9.3005
R290 drain_left.n21 drain_left.n20 9.3005
R291 drain_left.n6 drain_left.n5 9.3005
R292 drain_left.n15 drain_left.n14 9.3005
R293 drain_left.n13 drain_left.n12 9.3005
R294 drain_left.n62 drain_left.n61 9.3005
R295 drain_left.n35 drain_left.n34 9.3005
R296 drain_left.n56 drain_left.n55 9.3005
R297 drain_left.n54 drain_left.n53 9.3005
R298 drain_left.n39 drain_left.n38 9.3005
R299 drain_left.n48 drain_left.n47 9.3005
R300 drain_left.n46 drain_left.n45 9.3005
R301 drain_left.n27 drain_left.n2 8.92171
R302 drain_left.n60 drain_left.n35 8.92171
R303 drain_left.n28 drain_left.n0 8.14595
R304 drain_left.n61 drain_left.n33 8.14595
R305 drain_left drain_left.n65 6.54115
R306 drain_left.n30 drain_left.n0 5.81868
R307 drain_left.n63 drain_left.n33 5.81868
R308 drain_left.n28 drain_left.n27 5.04292
R309 drain_left.n61 drain_left.n60 5.04292
R310 drain_left.n13 drain_left.n9 4.38594
R311 drain_left.n46 drain_left.n42 4.38594
R312 drain_left.n24 drain_left.n2 4.26717
R313 drain_left.n57 drain_left.n35 4.26717
R314 drain_left.n23 drain_left.n4 3.49141
R315 drain_left.n56 drain_left.n37 3.49141
R316 drain_left.n31 drain_left.t1 3.3005
R317 drain_left.n31 drain_left.t2 3.3005
R318 drain_left.n64 drain_left.t0 3.3005
R319 drain_left.n64 drain_left.t5 3.3005
R320 drain_left.n20 drain_left.n19 2.71565
R321 drain_left.n53 drain_left.n52 2.71565
R322 drain_left.n16 drain_left.n6 1.93989
R323 drain_left.n49 drain_left.n39 1.93989
R324 drain_left.n15 drain_left.n8 1.16414
R325 drain_left.n48 drain_left.n41 1.16414
R326 drain_left.n12 drain_left.n11 0.388379
R327 drain_left.n45 drain_left.n44 0.388379
R328 drain_left.n14 drain_left.n13 0.155672
R329 drain_left.n14 drain_left.n5 0.155672
R330 drain_left.n21 drain_left.n5 0.155672
R331 drain_left.n22 drain_left.n21 0.155672
R332 drain_left.n22 drain_left.n1 0.155672
R333 drain_left.n29 drain_left.n1 0.155672
R334 drain_left.n62 drain_left.n34 0.155672
R335 drain_left.n55 drain_left.n34 0.155672
R336 drain_left.n55 drain_left.n54 0.155672
R337 drain_left.n54 drain_left.n38 0.155672
R338 drain_left.n47 drain_left.n38 0.155672
R339 drain_left.n47 drain_left.n46 0.155672
R340 minus.n1 minus.t3 284.284
R341 minus.n7 minus.t4 284.284
R342 minus.n2 minus.t0 262.69
R343 minus.n4 minus.t1 262.69
R344 minus.n8 minus.t5 262.69
R345 minus.n10 minus.t2 262.69
R346 minus.n5 minus.n4 161.3
R347 minus.n3 minus.n0 161.3
R348 minus.n11 minus.n10 161.3
R349 minus.n9 minus.n6 161.3
R350 minus.n1 minus.n0 44.8545
R351 minus.n7 minus.n6 44.8545
R352 minus.n12 minus.n5 30.5365
R353 minus.n4 minus.n3 26.2914
R354 minus.n10 minus.n9 26.2914
R355 minus.n3 minus.n2 21.9096
R356 minus.n9 minus.n8 21.9096
R357 minus.n2 minus.n1 20.3348
R358 minus.n8 minus.n7 20.3348
R359 minus.n12 minus.n11 6.62739
R360 minus.n5 minus.n0 0.189894
R361 minus.n11 minus.n6 0.189894
R362 minus minus.n12 0.188
R363 drain_right.n26 drain_right.n0 289.615
R364 drain_right.n60 drain_right.n34 289.615
R365 drain_right.n11 drain_right.n10 185
R366 drain_right.n8 drain_right.n7 185
R367 drain_right.n17 drain_right.n16 185
R368 drain_right.n19 drain_right.n18 185
R369 drain_right.n4 drain_right.n3 185
R370 drain_right.n25 drain_right.n24 185
R371 drain_right.n27 drain_right.n26 185
R372 drain_right.n61 drain_right.n60 185
R373 drain_right.n59 drain_right.n58 185
R374 drain_right.n38 drain_right.n37 185
R375 drain_right.n53 drain_right.n52 185
R376 drain_right.n51 drain_right.n50 185
R377 drain_right.n42 drain_right.n41 185
R378 drain_right.n45 drain_right.n44 185
R379 drain_right.t1 drain_right.n9 147.661
R380 drain_right.t4 drain_right.n43 147.661
R381 drain_right.n10 drain_right.n7 104.615
R382 drain_right.n17 drain_right.n7 104.615
R383 drain_right.n18 drain_right.n17 104.615
R384 drain_right.n18 drain_right.n3 104.615
R385 drain_right.n25 drain_right.n3 104.615
R386 drain_right.n26 drain_right.n25 104.615
R387 drain_right.n60 drain_right.n59 104.615
R388 drain_right.n59 drain_right.n37 104.615
R389 drain_right.n52 drain_right.n37 104.615
R390 drain_right.n52 drain_right.n51 104.615
R391 drain_right.n51 drain_right.n41 104.615
R392 drain_right.n44 drain_right.n41 104.615
R393 drain_right.n65 drain_right.n33 68.0786
R394 drain_right.n32 drain_right.n31 67.3573
R395 drain_right.n10 drain_right.t1 52.3082
R396 drain_right.n44 drain_right.t4 52.3082
R397 drain_right.n32 drain_right.n30 49.4747
R398 drain_right.n65 drain_right.n64 48.8641
R399 drain_right drain_right.n32 24.7102
R400 drain_right.n11 drain_right.n9 15.6674
R401 drain_right.n45 drain_right.n43 15.6674
R402 drain_right.n12 drain_right.n8 12.8005
R403 drain_right.n46 drain_right.n42 12.8005
R404 drain_right.n16 drain_right.n15 12.0247
R405 drain_right.n50 drain_right.n49 12.0247
R406 drain_right.n19 drain_right.n6 11.249
R407 drain_right.n53 drain_right.n40 11.249
R408 drain_right.n20 drain_right.n4 10.4732
R409 drain_right.n54 drain_right.n38 10.4732
R410 drain_right.n24 drain_right.n23 9.69747
R411 drain_right.n58 drain_right.n57 9.69747
R412 drain_right.n30 drain_right.n29 9.45567
R413 drain_right.n64 drain_right.n63 9.45567
R414 drain_right.n29 drain_right.n28 9.3005
R415 drain_right.n2 drain_right.n1 9.3005
R416 drain_right.n23 drain_right.n22 9.3005
R417 drain_right.n21 drain_right.n20 9.3005
R418 drain_right.n6 drain_right.n5 9.3005
R419 drain_right.n15 drain_right.n14 9.3005
R420 drain_right.n13 drain_right.n12 9.3005
R421 drain_right.n63 drain_right.n62 9.3005
R422 drain_right.n36 drain_right.n35 9.3005
R423 drain_right.n57 drain_right.n56 9.3005
R424 drain_right.n55 drain_right.n54 9.3005
R425 drain_right.n40 drain_right.n39 9.3005
R426 drain_right.n49 drain_right.n48 9.3005
R427 drain_right.n47 drain_right.n46 9.3005
R428 drain_right.n27 drain_right.n2 8.92171
R429 drain_right.n61 drain_right.n36 8.92171
R430 drain_right.n28 drain_right.n0 8.14595
R431 drain_right.n62 drain_right.n34 8.14595
R432 drain_right drain_right.n65 6.09718
R433 drain_right.n30 drain_right.n0 5.81868
R434 drain_right.n64 drain_right.n34 5.81868
R435 drain_right.n28 drain_right.n27 5.04292
R436 drain_right.n62 drain_right.n61 5.04292
R437 drain_right.n13 drain_right.n9 4.38594
R438 drain_right.n47 drain_right.n43 4.38594
R439 drain_right.n24 drain_right.n2 4.26717
R440 drain_right.n58 drain_right.n36 4.26717
R441 drain_right.n23 drain_right.n4 3.49141
R442 drain_right.n57 drain_right.n38 3.49141
R443 drain_right.n31 drain_right.t0 3.3005
R444 drain_right.n31 drain_right.t3 3.3005
R445 drain_right.n33 drain_right.t5 3.3005
R446 drain_right.n33 drain_right.t2 3.3005
R447 drain_right.n20 drain_right.n19 2.71565
R448 drain_right.n54 drain_right.n53 2.71565
R449 drain_right.n16 drain_right.n6 1.93989
R450 drain_right.n50 drain_right.n40 1.93989
R451 drain_right.n15 drain_right.n8 1.16414
R452 drain_right.n49 drain_right.n42 1.16414
R453 drain_right.n12 drain_right.n11 0.388379
R454 drain_right.n46 drain_right.n45 0.388379
R455 drain_right.n14 drain_right.n13 0.155672
R456 drain_right.n14 drain_right.n5 0.155672
R457 drain_right.n21 drain_right.n5 0.155672
R458 drain_right.n22 drain_right.n21 0.155672
R459 drain_right.n22 drain_right.n1 0.155672
R460 drain_right.n29 drain_right.n1 0.155672
R461 drain_right.n63 drain_right.n35 0.155672
R462 drain_right.n56 drain_right.n35 0.155672
R463 drain_right.n56 drain_right.n55 0.155672
R464 drain_right.n55 drain_right.n39 0.155672
R465 drain_right.n48 drain_right.n39 0.155672
R466 drain_right.n48 drain_right.n47 0.155672
C0 plus minus 3.95061f
C1 source drain_right 6.00219f
C2 source drain_left 6.0054f
C3 drain_left drain_right 0.706716f
C4 source plus 2.34789f
C5 plus drain_right 0.302454f
C6 plus drain_left 2.49746f
C7 source minus 2.33363f
C8 minus drain_right 2.35126f
C9 minus drain_left 0.171172f
C10 drain_right a_n1540_n2088# 4.65749f
C11 drain_left a_n1540_n2088# 4.89355f
C12 source a_n1540_n2088# 4.049316f
C13 minus a_n1540_n2088# 5.415394f
C14 plus a_n1540_n2088# 6.80693f
C15 drain_right.n0 a_n1540_n2088# 0.032782f
C16 drain_right.n1 a_n1540_n2088# 0.023323f
C17 drain_right.n2 a_n1540_n2088# 0.012533f
C18 drain_right.n3 a_n1540_n2088# 0.029622f
C19 drain_right.n4 a_n1540_n2088# 0.01327f
C20 drain_right.n5 a_n1540_n2088# 0.023323f
C21 drain_right.n6 a_n1540_n2088# 0.012533f
C22 drain_right.n7 a_n1540_n2088# 0.029622f
C23 drain_right.n8 a_n1540_n2088# 0.01327f
C24 drain_right.n9 a_n1540_n2088# 0.099804f
C25 drain_right.t1 a_n1540_n2088# 0.048281f
C26 drain_right.n10 a_n1540_n2088# 0.022217f
C27 drain_right.n11 a_n1540_n2088# 0.017498f
C28 drain_right.n12 a_n1540_n2088# 0.012533f
C29 drain_right.n13 a_n1540_n2088# 0.554938f
C30 drain_right.n14 a_n1540_n2088# 0.023323f
C31 drain_right.n15 a_n1540_n2088# 0.012533f
C32 drain_right.n16 a_n1540_n2088# 0.01327f
C33 drain_right.n17 a_n1540_n2088# 0.029622f
C34 drain_right.n18 a_n1540_n2088# 0.029622f
C35 drain_right.n19 a_n1540_n2088# 0.01327f
C36 drain_right.n20 a_n1540_n2088# 0.012533f
C37 drain_right.n21 a_n1540_n2088# 0.023323f
C38 drain_right.n22 a_n1540_n2088# 0.023323f
C39 drain_right.n23 a_n1540_n2088# 0.012533f
C40 drain_right.n24 a_n1540_n2088# 0.01327f
C41 drain_right.n25 a_n1540_n2088# 0.029622f
C42 drain_right.n26 a_n1540_n2088# 0.064127f
C43 drain_right.n27 a_n1540_n2088# 0.01327f
C44 drain_right.n28 a_n1540_n2088# 0.012533f
C45 drain_right.n29 a_n1540_n2088# 0.053909f
C46 drain_right.n30 a_n1540_n2088# 0.053117f
C47 drain_right.t0 a_n1540_n2088# 0.110581f
C48 drain_right.t3 a_n1540_n2088# 0.110581f
C49 drain_right.n31 a_n1540_n2088# 0.922943f
C50 drain_right.n32 a_n1540_n2088# 1.10942f
C51 drain_right.t5 a_n1540_n2088# 0.110581f
C52 drain_right.t2 a_n1540_n2088# 0.110581f
C53 drain_right.n33 a_n1540_n2088# 0.926579f
C54 drain_right.n34 a_n1540_n2088# 0.032782f
C55 drain_right.n35 a_n1540_n2088# 0.023323f
C56 drain_right.n36 a_n1540_n2088# 0.012533f
C57 drain_right.n37 a_n1540_n2088# 0.029622f
C58 drain_right.n38 a_n1540_n2088# 0.01327f
C59 drain_right.n39 a_n1540_n2088# 0.023323f
C60 drain_right.n40 a_n1540_n2088# 0.012533f
C61 drain_right.n41 a_n1540_n2088# 0.029622f
C62 drain_right.n42 a_n1540_n2088# 0.01327f
C63 drain_right.n43 a_n1540_n2088# 0.099804f
C64 drain_right.t4 a_n1540_n2088# 0.048281f
C65 drain_right.n44 a_n1540_n2088# 0.022217f
C66 drain_right.n45 a_n1540_n2088# 0.017498f
C67 drain_right.n46 a_n1540_n2088# 0.012533f
C68 drain_right.n47 a_n1540_n2088# 0.554938f
C69 drain_right.n48 a_n1540_n2088# 0.023323f
C70 drain_right.n49 a_n1540_n2088# 0.012533f
C71 drain_right.n50 a_n1540_n2088# 0.01327f
C72 drain_right.n51 a_n1540_n2088# 0.029622f
C73 drain_right.n52 a_n1540_n2088# 0.029622f
C74 drain_right.n53 a_n1540_n2088# 0.01327f
C75 drain_right.n54 a_n1540_n2088# 0.012533f
C76 drain_right.n55 a_n1540_n2088# 0.023323f
C77 drain_right.n56 a_n1540_n2088# 0.023323f
C78 drain_right.n57 a_n1540_n2088# 0.012533f
C79 drain_right.n58 a_n1540_n2088# 0.01327f
C80 drain_right.n59 a_n1540_n2088# 0.029622f
C81 drain_right.n60 a_n1540_n2088# 0.064127f
C82 drain_right.n61 a_n1540_n2088# 0.01327f
C83 drain_right.n62 a_n1540_n2088# 0.012533f
C84 drain_right.n63 a_n1540_n2088# 0.053909f
C85 drain_right.n64 a_n1540_n2088# 0.051985f
C86 drain_right.n65 a_n1540_n2088# 0.653798f
C87 minus.n0 a_n1540_n2088# 0.196542f
C88 minus.t3 a_n1540_n2088# 0.598597f
C89 minus.n1 a_n1540_n2088# 0.251334f
C90 minus.t0 a_n1540_n2088# 0.578321f
C91 minus.n2 a_n1540_n2088# 0.271079f
C92 minus.n3 a_n1540_n2088# 0.010772f
C93 minus.t1 a_n1540_n2088# 0.578321f
C94 minus.n4 a_n1540_n2088# 0.263724f
C95 minus.n5 a_n1540_n2088# 1.27826f
C96 minus.n6 a_n1540_n2088# 0.196542f
C97 minus.t4 a_n1540_n2088# 0.598597f
C98 minus.n7 a_n1540_n2088# 0.251334f
C99 minus.t5 a_n1540_n2088# 0.578321f
C100 minus.n8 a_n1540_n2088# 0.271079f
C101 minus.n9 a_n1540_n2088# 0.010772f
C102 minus.t2 a_n1540_n2088# 0.578321f
C103 minus.n10 a_n1540_n2088# 0.263724f
C104 minus.n11 a_n1540_n2088# 0.324524f
C105 minus.n12 a_n1540_n2088# 1.56866f
C106 drain_left.n0 a_n1540_n2088# 0.032816f
C107 drain_left.n1 a_n1540_n2088# 0.023347f
C108 drain_left.n2 a_n1540_n2088# 0.012545f
C109 drain_left.n3 a_n1540_n2088# 0.029653f
C110 drain_left.n4 a_n1540_n2088# 0.013283f
C111 drain_left.n5 a_n1540_n2088# 0.023347f
C112 drain_left.n6 a_n1540_n2088# 0.012545f
C113 drain_left.n7 a_n1540_n2088# 0.029653f
C114 drain_left.n8 a_n1540_n2088# 0.013283f
C115 drain_left.n9 a_n1540_n2088# 0.099907f
C116 drain_left.t3 a_n1540_n2088# 0.04833f
C117 drain_left.n10 a_n1540_n2088# 0.02224f
C118 drain_left.n11 a_n1540_n2088# 0.017516f
C119 drain_left.n12 a_n1540_n2088# 0.012545f
C120 drain_left.n13 a_n1540_n2088# 0.55551f
C121 drain_left.n14 a_n1540_n2088# 0.023347f
C122 drain_left.n15 a_n1540_n2088# 0.012545f
C123 drain_left.n16 a_n1540_n2088# 0.013283f
C124 drain_left.n17 a_n1540_n2088# 0.029653f
C125 drain_left.n18 a_n1540_n2088# 0.029653f
C126 drain_left.n19 a_n1540_n2088# 0.013283f
C127 drain_left.n20 a_n1540_n2088# 0.012545f
C128 drain_left.n21 a_n1540_n2088# 0.023347f
C129 drain_left.n22 a_n1540_n2088# 0.023347f
C130 drain_left.n23 a_n1540_n2088# 0.012545f
C131 drain_left.n24 a_n1540_n2088# 0.013283f
C132 drain_left.n25 a_n1540_n2088# 0.029653f
C133 drain_left.n26 a_n1540_n2088# 0.064193f
C134 drain_left.n27 a_n1540_n2088# 0.013283f
C135 drain_left.n28 a_n1540_n2088# 0.012545f
C136 drain_left.n29 a_n1540_n2088# 0.053965f
C137 drain_left.n30 a_n1540_n2088# 0.053172f
C138 drain_left.t1 a_n1540_n2088# 0.110695f
C139 drain_left.t2 a_n1540_n2088# 0.110695f
C140 drain_left.n31 a_n1540_n2088# 0.923896f
C141 drain_left.n32 a_n1540_n2088# 1.15822f
C142 drain_left.n33 a_n1540_n2088# 0.032816f
C143 drain_left.n34 a_n1540_n2088# 0.023347f
C144 drain_left.n35 a_n1540_n2088# 0.012545f
C145 drain_left.n36 a_n1540_n2088# 0.029653f
C146 drain_left.n37 a_n1540_n2088# 0.013283f
C147 drain_left.n38 a_n1540_n2088# 0.023347f
C148 drain_left.n39 a_n1540_n2088# 0.012545f
C149 drain_left.n40 a_n1540_n2088# 0.029653f
C150 drain_left.n41 a_n1540_n2088# 0.013283f
C151 drain_left.n42 a_n1540_n2088# 0.099907f
C152 drain_left.t4 a_n1540_n2088# 0.04833f
C153 drain_left.n43 a_n1540_n2088# 0.02224f
C154 drain_left.n44 a_n1540_n2088# 0.017516f
C155 drain_left.n45 a_n1540_n2088# 0.012545f
C156 drain_left.n46 a_n1540_n2088# 0.55551f
C157 drain_left.n47 a_n1540_n2088# 0.023347f
C158 drain_left.n48 a_n1540_n2088# 0.012545f
C159 drain_left.n49 a_n1540_n2088# 0.013283f
C160 drain_left.n50 a_n1540_n2088# 0.029653f
C161 drain_left.n51 a_n1540_n2088# 0.029653f
C162 drain_left.n52 a_n1540_n2088# 0.013283f
C163 drain_left.n53 a_n1540_n2088# 0.012545f
C164 drain_left.n54 a_n1540_n2088# 0.023347f
C165 drain_left.n55 a_n1540_n2088# 0.023347f
C166 drain_left.n56 a_n1540_n2088# 0.012545f
C167 drain_left.n57 a_n1540_n2088# 0.013283f
C168 drain_left.n58 a_n1540_n2088# 0.029653f
C169 drain_left.n59 a_n1540_n2088# 0.064193f
C170 drain_left.n60 a_n1540_n2088# 0.013283f
C171 drain_left.n61 a_n1540_n2088# 0.012545f
C172 drain_left.n62 a_n1540_n2088# 0.053965f
C173 drain_left.n63 a_n1540_n2088# 0.054034f
C174 drain_left.t0 a_n1540_n2088# 0.110695f
C175 drain_left.t5 a_n1540_n2088# 0.110695f
C176 drain_left.n64 a_n1540_n2088# 0.923199f
C177 drain_left.n65 a_n1540_n2088# 0.639345f
C178 source.n0 a_n1540_n2088# 0.036161f
C179 source.n1 a_n1540_n2088# 0.025726f
C180 source.n2 a_n1540_n2088# 0.013824f
C181 source.n3 a_n1540_n2088# 0.032675f
C182 source.n4 a_n1540_n2088# 0.014637f
C183 source.n5 a_n1540_n2088# 0.025726f
C184 source.n6 a_n1540_n2088# 0.013824f
C185 source.n7 a_n1540_n2088# 0.032675f
C186 source.n8 a_n1540_n2088# 0.014637f
C187 source.n9 a_n1540_n2088# 0.110091f
C188 source.t6 a_n1540_n2088# 0.053257f
C189 source.n10 a_n1540_n2088# 0.024507f
C190 source.n11 a_n1540_n2088# 0.019301f
C191 source.n12 a_n1540_n2088# 0.013824f
C192 source.n13 a_n1540_n2088# 0.612133f
C193 source.n14 a_n1540_n2088# 0.025726f
C194 source.n15 a_n1540_n2088# 0.013824f
C195 source.n16 a_n1540_n2088# 0.014637f
C196 source.n17 a_n1540_n2088# 0.032675f
C197 source.n18 a_n1540_n2088# 0.032675f
C198 source.n19 a_n1540_n2088# 0.014637f
C199 source.n20 a_n1540_n2088# 0.013824f
C200 source.n21 a_n1540_n2088# 0.025726f
C201 source.n22 a_n1540_n2088# 0.025726f
C202 source.n23 a_n1540_n2088# 0.013824f
C203 source.n24 a_n1540_n2088# 0.014637f
C204 source.n25 a_n1540_n2088# 0.032675f
C205 source.n26 a_n1540_n2088# 0.070737f
C206 source.n27 a_n1540_n2088# 0.014637f
C207 source.n28 a_n1540_n2088# 0.013824f
C208 source.n29 a_n1540_n2088# 0.059465f
C209 source.n30 a_n1540_n2088# 0.03958f
C210 source.n31 a_n1540_n2088# 0.672064f
C211 source.t10 a_n1540_n2088# 0.121978f
C212 source.t11 a_n1540_n2088# 0.121978f
C213 source.n32 a_n1540_n2088# 0.949977f
C214 source.n33 a_n1540_n2088# 0.390515f
C215 source.n34 a_n1540_n2088# 0.036161f
C216 source.n35 a_n1540_n2088# 0.025726f
C217 source.n36 a_n1540_n2088# 0.013824f
C218 source.n37 a_n1540_n2088# 0.032675f
C219 source.n38 a_n1540_n2088# 0.014637f
C220 source.n39 a_n1540_n2088# 0.025726f
C221 source.n40 a_n1540_n2088# 0.013824f
C222 source.n41 a_n1540_n2088# 0.032675f
C223 source.n42 a_n1540_n2088# 0.014637f
C224 source.n43 a_n1540_n2088# 0.110091f
C225 source.t0 a_n1540_n2088# 0.053257f
C226 source.n44 a_n1540_n2088# 0.024507f
C227 source.n45 a_n1540_n2088# 0.019301f
C228 source.n46 a_n1540_n2088# 0.013824f
C229 source.n47 a_n1540_n2088# 0.612133f
C230 source.n48 a_n1540_n2088# 0.025726f
C231 source.n49 a_n1540_n2088# 0.013824f
C232 source.n50 a_n1540_n2088# 0.014637f
C233 source.n51 a_n1540_n2088# 0.032675f
C234 source.n52 a_n1540_n2088# 0.032675f
C235 source.n53 a_n1540_n2088# 0.014637f
C236 source.n54 a_n1540_n2088# 0.013824f
C237 source.n55 a_n1540_n2088# 0.025726f
C238 source.n56 a_n1540_n2088# 0.025726f
C239 source.n57 a_n1540_n2088# 0.013824f
C240 source.n58 a_n1540_n2088# 0.014637f
C241 source.n59 a_n1540_n2088# 0.032675f
C242 source.n60 a_n1540_n2088# 0.070737f
C243 source.n61 a_n1540_n2088# 0.014637f
C244 source.n62 a_n1540_n2088# 0.013824f
C245 source.n63 a_n1540_n2088# 0.059465f
C246 source.n64 a_n1540_n2088# 0.03958f
C247 source.n65 a_n1540_n2088# 0.171328f
C248 source.t2 a_n1540_n2088# 0.121978f
C249 source.t3 a_n1540_n2088# 0.121978f
C250 source.n66 a_n1540_n2088# 0.949977f
C251 source.n67 a_n1540_n2088# 1.30431f
C252 source.t7 a_n1540_n2088# 0.121978f
C253 source.t8 a_n1540_n2088# 0.121978f
C254 source.n68 a_n1540_n2088# 0.949971f
C255 source.n69 a_n1540_n2088# 1.30431f
C256 source.n70 a_n1540_n2088# 0.036161f
C257 source.n71 a_n1540_n2088# 0.025726f
C258 source.n72 a_n1540_n2088# 0.013824f
C259 source.n73 a_n1540_n2088# 0.032675f
C260 source.n74 a_n1540_n2088# 0.014637f
C261 source.n75 a_n1540_n2088# 0.025726f
C262 source.n76 a_n1540_n2088# 0.013824f
C263 source.n77 a_n1540_n2088# 0.032675f
C264 source.n78 a_n1540_n2088# 0.014637f
C265 source.n79 a_n1540_n2088# 0.110091f
C266 source.t9 a_n1540_n2088# 0.053257f
C267 source.n80 a_n1540_n2088# 0.024507f
C268 source.n81 a_n1540_n2088# 0.019301f
C269 source.n82 a_n1540_n2088# 0.013824f
C270 source.n83 a_n1540_n2088# 0.612133f
C271 source.n84 a_n1540_n2088# 0.025726f
C272 source.n85 a_n1540_n2088# 0.013824f
C273 source.n86 a_n1540_n2088# 0.014637f
C274 source.n87 a_n1540_n2088# 0.032675f
C275 source.n88 a_n1540_n2088# 0.032675f
C276 source.n89 a_n1540_n2088# 0.014637f
C277 source.n90 a_n1540_n2088# 0.013824f
C278 source.n91 a_n1540_n2088# 0.025726f
C279 source.n92 a_n1540_n2088# 0.025726f
C280 source.n93 a_n1540_n2088# 0.013824f
C281 source.n94 a_n1540_n2088# 0.014637f
C282 source.n95 a_n1540_n2088# 0.032675f
C283 source.n96 a_n1540_n2088# 0.070737f
C284 source.n97 a_n1540_n2088# 0.014637f
C285 source.n98 a_n1540_n2088# 0.013824f
C286 source.n99 a_n1540_n2088# 0.059465f
C287 source.n100 a_n1540_n2088# 0.03958f
C288 source.n101 a_n1540_n2088# 0.171328f
C289 source.t5 a_n1540_n2088# 0.121978f
C290 source.t4 a_n1540_n2088# 0.121978f
C291 source.n102 a_n1540_n2088# 0.949971f
C292 source.n103 a_n1540_n2088# 0.390522f
C293 source.n104 a_n1540_n2088# 0.036161f
C294 source.n105 a_n1540_n2088# 0.025726f
C295 source.n106 a_n1540_n2088# 0.013824f
C296 source.n107 a_n1540_n2088# 0.032675f
C297 source.n108 a_n1540_n2088# 0.014637f
C298 source.n109 a_n1540_n2088# 0.025726f
C299 source.n110 a_n1540_n2088# 0.013824f
C300 source.n111 a_n1540_n2088# 0.032675f
C301 source.n112 a_n1540_n2088# 0.014637f
C302 source.n113 a_n1540_n2088# 0.110091f
C303 source.t1 a_n1540_n2088# 0.053257f
C304 source.n114 a_n1540_n2088# 0.024507f
C305 source.n115 a_n1540_n2088# 0.019301f
C306 source.n116 a_n1540_n2088# 0.013824f
C307 source.n117 a_n1540_n2088# 0.612133f
C308 source.n118 a_n1540_n2088# 0.025726f
C309 source.n119 a_n1540_n2088# 0.013824f
C310 source.n120 a_n1540_n2088# 0.014637f
C311 source.n121 a_n1540_n2088# 0.032675f
C312 source.n122 a_n1540_n2088# 0.032675f
C313 source.n123 a_n1540_n2088# 0.014637f
C314 source.n124 a_n1540_n2088# 0.013824f
C315 source.n125 a_n1540_n2088# 0.025726f
C316 source.n126 a_n1540_n2088# 0.025726f
C317 source.n127 a_n1540_n2088# 0.013824f
C318 source.n128 a_n1540_n2088# 0.014637f
C319 source.n129 a_n1540_n2088# 0.032675f
C320 source.n130 a_n1540_n2088# 0.070737f
C321 source.n131 a_n1540_n2088# 0.014637f
C322 source.n132 a_n1540_n2088# 0.013824f
C323 source.n133 a_n1540_n2088# 0.059465f
C324 source.n134 a_n1540_n2088# 0.03958f
C325 source.n135 a_n1540_n2088# 0.302339f
C326 source.n136 a_n1540_n2088# 1.06692f
C327 plus.n0 a_n1540_n2088# 0.20102f
C328 plus.t0 a_n1540_n2088# 0.591496f
C329 plus.t5 a_n1540_n2088# 0.591496f
C330 plus.t1 a_n1540_n2088# 0.612233f
C331 plus.n1 a_n1540_n2088# 0.25706f
C332 plus.n2 a_n1540_n2088# 0.277254f
C333 plus.n3 a_n1540_n2088# 0.011018f
C334 plus.n4 a_n1540_n2088# 0.269732f
C335 plus.n5 a_n1540_n2088# 0.431187f
C336 plus.n6 a_n1540_n2088# 0.20102f
C337 plus.t2 a_n1540_n2088# 0.591496f
C338 plus.t3 a_n1540_n2088# 0.612233f
C339 plus.n7 a_n1540_n2088# 0.25706f
C340 plus.t4 a_n1540_n2088# 0.591496f
C341 plus.n8 a_n1540_n2088# 0.277254f
C342 plus.n9 a_n1540_n2088# 0.011018f
C343 plus.n10 a_n1540_n2088# 0.269732f
C344 plus.n11 a_n1540_n2088# 1.18274f
.ends

