* NGSPICE file created from diffpair33.ext - technology: sky130A

.subckt diffpair33 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t12 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 drain_right.t7 minus.t0 source.t2 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X2 source.t5 minus.t1 drain_right.t6 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 source.t11 plus.t1 drain_left.t6 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 source.t10 plus.t2 drain_left.t5 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X5 drain_right.t5 minus.t2 source.t7 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X6 a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X7 drain_left.t4 plus.t3 source.t9 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X8 drain_left.t3 plus.t4 source.t13 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X9 source.t6 minus.t3 drain_right.t4 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X10 drain_right.t3 minus.t4 source.t1 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X11 source.t3 minus.t5 drain_right.t2 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X12 source.t14 plus.t5 drain_left.t2 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X13 source.t8 plus.t6 drain_left.t1 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X15 drain_right.t1 minus.t6 source.t4 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X16 a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X17 source.t0 minus.t7 drain_right.t0 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X18 a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X19 drain_left.t0 plus.t7 source.t15 a_n1346_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
R0 plus.n2 plus.t2 213.25
R1 plus.n7 plus.t7 213.25
R2 plus.n11 plus.t4 213.25
R3 plus.n16 plus.t5 213.25
R4 plus.n1 plus.t3 184.768
R5 plus.n6 plus.t6 184.768
R6 plus.n10 plus.t1 184.768
R7 plus.n15 plus.t0 184.768
R8 plus.n3 plus.n2 161.489
R9 plus.n12 plus.n11 161.489
R10 plus.n4 plus.n3 161.3
R11 plus.n5 plus.n0 161.3
R12 plus.n8 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n14 plus.n9 161.3
R15 plus.n17 plus.n16 161.3
R16 plus.n5 plus.n4 73.0308
R17 plus.n14 plus.n13 73.0308
R18 plus.n2 plus.n1 63.5369
R19 plus.n7 plus.n6 63.5369
R20 plus.n16 plus.n15 63.5369
R21 plus.n11 plus.n10 63.5369
R22 plus plus.n17 23.8967
R23 plus.n4 plus.n1 9.49444
R24 plus.n6 plus.n5 9.49444
R25 plus.n15 plus.n14 9.49444
R26 plus.n13 plus.n10 9.49444
R27 plus plus.n8 7.93989
R28 plus.n3 plus.n0 0.189894
R29 plus.n8 plus.n0 0.189894
R30 plus.n17 plus.n9 0.189894
R31 plus.n12 plus.n9 0.189894
R32 source.n0 source.t15 243.255
R33 source.n3 source.t10 243.255
R34 source.n4 source.t1 243.255
R35 source.n7 source.t6 243.255
R36 source.n15 source.t4 243.254
R37 source.n12 source.t3 243.254
R38 source.n11 source.t13 243.254
R39 source.n8 source.t14 243.254
R40 source.n2 source.n1 223.454
R41 source.n6 source.n5 223.454
R42 source.n14 source.n13 223.453
R43 source.n10 source.n9 223.453
R44 source.n13 source.t7 19.8005
R45 source.n13 source.t5 19.8005
R46 source.n9 source.t12 19.8005
R47 source.n9 source.t11 19.8005
R48 source.n1 source.t9 19.8005
R49 source.n1 source.t8 19.8005
R50 source.n5 source.t2 19.8005
R51 source.n5 source.t0 19.8005
R52 source.n8 source.n7 13.4975
R53 source.n16 source.n0 7.96301
R54 source.n16 source.n15 5.53498
R55 source.n7 source.n6 0.543603
R56 source.n6 source.n4 0.543603
R57 source.n3 source.n2 0.543603
R58 source.n2 source.n0 0.543603
R59 source.n10 source.n8 0.543603
R60 source.n11 source.n10 0.543603
R61 source.n14 source.n12 0.543603
R62 source.n15 source.n14 0.543603
R63 source.n4 source.n3 0.470328
R64 source.n12 source.n11 0.470328
R65 source source.n16 0.188
R66 drain_left.n5 drain_left.n3 240.675
R67 drain_left.n2 drain_left.n1 240.349
R68 drain_left.n2 drain_left.n0 240.349
R69 drain_left.n5 drain_left.n4 240.132
R70 drain_left drain_left.n2 20.9346
R71 drain_left.n1 drain_left.t6 19.8005
R72 drain_left.n1 drain_left.t3 19.8005
R73 drain_left.n0 drain_left.t2 19.8005
R74 drain_left.n0 drain_left.t7 19.8005
R75 drain_left.n4 drain_left.t1 19.8005
R76 drain_left.n4 drain_left.t0 19.8005
R77 drain_left.n3 drain_left.t5 19.8005
R78 drain_left.n3 drain_left.t4 19.8005
R79 drain_left drain_left.n5 6.19632
R80 minus.n7 minus.t3 213.25
R81 minus.n2 minus.t4 213.25
R82 minus.n16 minus.t6 213.25
R83 minus.n11 minus.t5 213.25
R84 minus.n6 minus.t0 184.768
R85 minus.n1 minus.t7 184.768
R86 minus.n15 minus.t1 184.768
R87 minus.n10 minus.t2 184.768
R88 minus.n3 minus.n2 161.489
R89 minus.n12 minus.n11 161.489
R90 minus.n8 minus.n7 161.3
R91 minus.n5 minus.n0 161.3
R92 minus.n4 minus.n3 161.3
R93 minus.n17 minus.n16 161.3
R94 minus.n14 minus.n9 161.3
R95 minus.n13 minus.n12 161.3
R96 minus.n5 minus.n4 73.0308
R97 minus.n14 minus.n13 73.0308
R98 minus.n7 minus.n6 63.5369
R99 minus.n2 minus.n1 63.5369
R100 minus.n11 minus.n10 63.5369
R101 minus.n16 minus.n15 63.5369
R102 minus.n18 minus.n8 25.849
R103 minus.n6 minus.n5 9.49444
R104 minus.n4 minus.n1 9.49444
R105 minus.n13 minus.n10 9.49444
R106 minus.n15 minus.n14 9.49444
R107 minus.n18 minus.n17 6.46262
R108 minus.n8 minus.n0 0.189894
R109 minus.n3 minus.n0 0.189894
R110 minus.n12 minus.n9 0.189894
R111 minus.n17 minus.n9 0.189894
R112 minus minus.n18 0.188
R113 drain_right.n5 drain_right.n3 240.675
R114 drain_right.n2 drain_right.n1 240.349
R115 drain_right.n2 drain_right.n0 240.349
R116 drain_right.n5 drain_right.n4 240.132
R117 drain_right drain_right.n2 20.3814
R118 drain_right.n1 drain_right.t6 19.8005
R119 drain_right.n1 drain_right.t1 19.8005
R120 drain_right.n0 drain_right.t2 19.8005
R121 drain_right.n0 drain_right.t5 19.8005
R122 drain_right.n3 drain_right.t0 19.8005
R123 drain_right.n3 drain_right.t3 19.8005
R124 drain_right.n4 drain_right.t4 19.8005
R125 drain_right.n4 drain_right.t7 19.8005
R126 drain_right drain_right.n5 6.19632
C0 plus drain_right 0.288823f
C1 drain_right source 3.04867f
C2 drain_right drain_left 0.630134f
C3 plus minus 2.80431f
C4 source minus 0.762735f
C5 drain_left minus 0.177709f
C6 drain_right minus 0.60616f
C7 plus source 0.776599f
C8 plus drain_left 0.733309f
C9 drain_left source 3.04949f
C10 drain_right a_n1346_n1088# 2.836174f
C11 drain_left a_n1346_n1088# 2.99356f
C12 source a_n1346_n1088# 2.284312f
C13 minus a_n1346_n1088# 4.29638f
C14 plus a_n1346_n1088# 5.00257f
C15 drain_right.t2 a_n1346_n1088# 0.017973f
C16 drain_right.t5 a_n1346_n1088# 0.017973f
C17 drain_right.n0 a_n1346_n1088# 0.070041f
C18 drain_right.t6 a_n1346_n1088# 0.017973f
C19 drain_right.t1 a_n1346_n1088# 0.017973f
C20 drain_right.n1 a_n1346_n1088# 0.070041f
C21 drain_right.n2 a_n1346_n1088# 0.910282f
C22 drain_right.t0 a_n1346_n1088# 0.017973f
C23 drain_right.t3 a_n1346_n1088# 0.017973f
C24 drain_right.n3 a_n1346_n1088# 0.070396f
C25 drain_right.t4 a_n1346_n1088# 0.017973f
C26 drain_right.t7 a_n1346_n1088# 0.017973f
C27 drain_right.n4 a_n1346_n1088# 0.069837f
C28 drain_right.n5 a_n1346_n1088# 0.675217f
C29 minus.n0 a_n1346_n1088# 0.03682f
C30 minus.t3 a_n1346_n1088# 0.038723f
C31 minus.t0 a_n1346_n1088# 0.034052f
C32 minus.t7 a_n1346_n1088# 0.034052f
C33 minus.n1 a_n1346_n1088# 0.035084f
C34 minus.t4 a_n1346_n1088# 0.038723f
C35 minus.n2 a_n1346_n1088# 0.045513f
C36 minus.n3 a_n1346_n1088# 0.077905f
C37 minus.n4 a_n1346_n1088# 0.01369f
C38 minus.n5 a_n1346_n1088# 0.01369f
C39 minus.n6 a_n1346_n1088# 0.035084f
C40 minus.n7 a_n1346_n1088# 0.045465f
C41 minus.n8 a_n1346_n1088# 0.73366f
C42 minus.n9 a_n1346_n1088# 0.03682f
C43 minus.t1 a_n1346_n1088# 0.034052f
C44 minus.t2 a_n1346_n1088# 0.034052f
C45 minus.n10 a_n1346_n1088# 0.035084f
C46 minus.t5 a_n1346_n1088# 0.038723f
C47 minus.n11 a_n1346_n1088# 0.045513f
C48 minus.n12 a_n1346_n1088# 0.077905f
C49 minus.n13 a_n1346_n1088# 0.01369f
C50 minus.n14 a_n1346_n1088# 0.01369f
C51 minus.n15 a_n1346_n1088# 0.035084f
C52 minus.t6 a_n1346_n1088# 0.038723f
C53 minus.n16 a_n1346_n1088# 0.045465f
C54 minus.n17 a_n1346_n1088# 0.237473f
C55 minus.n18 a_n1346_n1088# 0.907086f
C56 drain_left.t2 a_n1346_n1088# 0.017455f
C57 drain_left.t7 a_n1346_n1088# 0.017455f
C58 drain_left.n0 a_n1346_n1088# 0.068023f
C59 drain_left.t6 a_n1346_n1088# 0.017455f
C60 drain_left.t3 a_n1346_n1088# 0.017455f
C61 drain_left.n1 a_n1346_n1088# 0.068023f
C62 drain_left.n2 a_n1346_n1088# 0.926896f
C63 drain_left.t5 a_n1346_n1088# 0.017455f
C64 drain_left.t4 a_n1346_n1088# 0.017455f
C65 drain_left.n3 a_n1346_n1088# 0.068369f
C66 drain_left.t1 a_n1346_n1088# 0.017455f
C67 drain_left.t0 a_n1346_n1088# 0.017455f
C68 drain_left.n4 a_n1346_n1088# 0.067826f
C69 drain_left.n5 a_n1346_n1088# 0.655769f
C70 source.t15 a_n1346_n1088# 0.110318f
C71 source.n0 a_n1346_n1088# 0.473687f
C72 source.t9 a_n1346_n1088# 0.019821f
C73 source.t8 a_n1346_n1088# 0.019821f
C74 source.n1 a_n1346_n1088# 0.064281f
C75 source.n2 a_n1346_n1088# 0.241831f
C76 source.t10 a_n1346_n1088# 0.110318f
C77 source.n3 a_n1346_n1088# 0.243928f
C78 source.t1 a_n1346_n1088# 0.110318f
C79 source.n4 a_n1346_n1088# 0.243928f
C80 source.t2 a_n1346_n1088# 0.019821f
C81 source.t0 a_n1346_n1088# 0.019821f
C82 source.n5 a_n1346_n1088# 0.064281f
C83 source.n6 a_n1346_n1088# 0.241831f
C84 source.t6 a_n1346_n1088# 0.110318f
C85 source.n7 a_n1346_n1088# 0.674668f
C86 source.t14 a_n1346_n1088# 0.110318f
C87 source.n8 a_n1346_n1088# 0.674669f
C88 source.t12 a_n1346_n1088# 0.019821f
C89 source.t11 a_n1346_n1088# 0.019821f
C90 source.n9 a_n1346_n1088# 0.064281f
C91 source.n10 a_n1346_n1088# 0.241831f
C92 source.t13 a_n1346_n1088# 0.110318f
C93 source.n11 a_n1346_n1088# 0.243928f
C94 source.t3 a_n1346_n1088# 0.110318f
C95 source.n12 a_n1346_n1088# 0.243928f
C96 source.t7 a_n1346_n1088# 0.019821f
C97 source.t5 a_n1346_n1088# 0.019821f
C98 source.n13 a_n1346_n1088# 0.064281f
C99 source.n14 a_n1346_n1088# 0.241831f
C100 source.t4 a_n1346_n1088# 0.110318f
C101 source.n15 a_n1346_n1088# 0.385515f
C102 source.n16 a_n1346_n1088# 0.507975f
C103 plus.n0 a_n1346_n1088# 0.037826f
C104 plus.t6 a_n1346_n1088# 0.034982f
C105 plus.t3 a_n1346_n1088# 0.034982f
C106 plus.n1 a_n1346_n1088# 0.036042f
C107 plus.t2 a_n1346_n1088# 0.03978f
C108 plus.n2 a_n1346_n1088# 0.046757f
C109 plus.n3 a_n1346_n1088# 0.080034f
C110 plus.n4 a_n1346_n1088# 0.014064f
C111 plus.n5 a_n1346_n1088# 0.014064f
C112 plus.n6 a_n1346_n1088# 0.036042f
C113 plus.t7 a_n1346_n1088# 0.03978f
C114 plus.n7 a_n1346_n1088# 0.046707f
C115 plus.n8 a_n1346_n1088# 0.25582f
C116 plus.n9 a_n1346_n1088# 0.037826f
C117 plus.t5 a_n1346_n1088# 0.03978f
C118 plus.t0 a_n1346_n1088# 0.034982f
C119 plus.t1 a_n1346_n1088# 0.034982f
C120 plus.n10 a_n1346_n1088# 0.036042f
C121 plus.t4 a_n1346_n1088# 0.03978f
C122 plus.n11 a_n1346_n1088# 0.046757f
C123 plus.n12 a_n1346_n1088# 0.080034f
C124 plus.n13 a_n1346_n1088# 0.014064f
C125 plus.n14 a_n1346_n1088# 0.014064f
C126 plus.n15 a_n1346_n1088# 0.036042f
C127 plus.n16 a_n1346_n1088# 0.046707f
C128 plus.n17 a_n1346_n1088# 0.736306f
.ends

