* NGSPICE file created from diffpair652.ext - technology: sky130A

.subckt diffpair652 minus drain_right drain_left source plus
X0 a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.2
X1 source plus drain_left a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X2 drain_right minus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X3 source plus drain_left a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X4 drain_right minus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X5 drain_right minus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X6 source minus drain_right a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X7 a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X8 source minus drain_right a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.2
X9 drain_left plus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
X10 a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X11 drain_right minus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X12 a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.2
X13 drain_left plus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X14 drain_left plus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.2
X15 drain_left plus source a_n1140_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.2
.ends

