* NGSPICE file created from diffpair476.ext - technology: sky130A

.subckt diffpair476 minus drain_right drain_left source plus
X0 a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X1 a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X2 source.t26 minus.t0 drain_right.t8 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X3 a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X4 source.t25 minus.t1 drain_right.t9 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X5 a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X6 source.t0 plus.t0 drain_left.t13 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X7 source.t7 plus.t1 drain_left.t12 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X8 source.t24 minus.t2 drain_right.t0 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X9 drain_left.t11 plus.t2 source.t5 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X10 drain_right.t6 minus.t3 source.t23 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X11 source.t22 minus.t4 drain_right.t7 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X12 drain_right.t3 minus.t5 source.t21 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X13 drain_right.t2 minus.t6 source.t20 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X14 source.t19 minus.t7 drain_right.t1 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X15 drain_left.t10 plus.t3 source.t12 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X16 source.t18 minus.t8 drain_right.t10 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X17 drain_left.t9 plus.t4 source.t4 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X18 drain_right.t5 minus.t9 source.t17 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X19 drain_right.t4 minus.t10 source.t16 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X20 drain_left.t8 plus.t5 source.t8 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X21 drain_right.t13 minus.t11 source.t15 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X22 source.t11 plus.t6 drain_left.t7 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X23 source.t10 plus.t7 drain_left.t6 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X24 drain_left.t5 plus.t8 source.t3 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X25 drain_left.t4 plus.t9 source.t6 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X26 drain_left.t3 plus.t10 source.t27 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X27 source.t2 plus.t11 drain_left.t2 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X28 drain_right.t12 minus.t12 source.t14 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X29 drain_left.t1 plus.t12 source.t9 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X30 drain_right.t11 minus.t13 source.t13 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X31 source.t1 plus.t13 drain_left.t0 a_n2524_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
R0 minus.n5 minus.t6 434.45
R1 minus.n23 minus.t13 434.45
R2 minus.n4 minus.t4 410.604
R3 minus.n8 minus.t3 410.604
R4 minus.n9 minus.t8 410.604
R5 minus.n10 minus.t9 410.604
R6 minus.n14 minus.t7 410.604
R7 minus.n16 minus.t5 410.604
R8 minus.n22 minus.t2 410.604
R9 minus.n26 minus.t11 410.604
R10 minus.n27 minus.t1 410.604
R11 minus.n28 minus.t12 410.604
R12 minus.n32 minus.t0 410.604
R13 minus.n34 minus.t10 410.604
R14 minus.n17 minus.n16 161.3
R15 minus.n15 minus.n0 161.3
R16 minus.n14 minus.n13 161.3
R17 minus.n12 minus.n1 161.3
R18 minus.n6 minus.n3 161.3
R19 minus.n35 minus.n34 161.3
R20 minus.n33 minus.n18 161.3
R21 minus.n32 minus.n31 161.3
R22 minus.n30 minus.n19 161.3
R23 minus.n24 minus.n21 161.3
R24 minus.n11 minus.n10 80.6037
R25 minus.n9 minus.n2 80.6037
R26 minus.n8 minus.n7 80.6037
R27 minus.n29 minus.n28 80.6037
R28 minus.n27 minus.n20 80.6037
R29 minus.n26 minus.n25 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n6 minus.n5 44.9119
R35 minus.n24 minus.n23 44.9119
R36 minus.n36 minus.n17 38.9077
R37 minus.n16 minus.n15 35.055
R38 minus.n34 minus.n33 35.055
R39 minus.n8 minus.n3 32.1338
R40 minus.n10 minus.n1 32.1338
R41 minus.n26 minus.n21 32.1338
R42 minus.n28 minus.n19 32.1338
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n4 minus.n3 16.0672
R46 minus.n14 minus.n1 16.0672
R47 minus.n22 minus.n21 16.0672
R48 minus.n32 minus.n19 16.0672
R49 minus.n15 minus.n14 13.146
R50 minus.n33 minus.n32 13.146
R51 minus.n36 minus.n35 6.72588
R52 minus.n11 minus.n2 0.380177
R53 minus.n7 minus.n2 0.380177
R54 minus.n25 minus.n20 0.380177
R55 minus.n29 minus.n20 0.380177
R56 minus.n12 minus.n11 0.285035
R57 minus.n7 minus.n6 0.285035
R58 minus.n25 minus.n24 0.285035
R59 minus.n30 minus.n29 0.285035
R60 minus.n17 minus.n0 0.189894
R61 minus.n13 minus.n0 0.189894
R62 minus.n13 minus.n12 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 drain_right.n60 drain_right.n0 289.615
R68 drain_right.n136 drain_right.n76 289.615
R69 drain_right.n20 drain_right.n19 185
R70 drain_right.n25 drain_right.n24 185
R71 drain_right.n27 drain_right.n26 185
R72 drain_right.n16 drain_right.n15 185
R73 drain_right.n33 drain_right.n32 185
R74 drain_right.n35 drain_right.n34 185
R75 drain_right.n12 drain_right.n11 185
R76 drain_right.n42 drain_right.n41 185
R77 drain_right.n43 drain_right.n10 185
R78 drain_right.n45 drain_right.n44 185
R79 drain_right.n8 drain_right.n7 185
R80 drain_right.n51 drain_right.n50 185
R81 drain_right.n53 drain_right.n52 185
R82 drain_right.n4 drain_right.n3 185
R83 drain_right.n59 drain_right.n58 185
R84 drain_right.n61 drain_right.n60 185
R85 drain_right.n137 drain_right.n136 185
R86 drain_right.n135 drain_right.n134 185
R87 drain_right.n80 drain_right.n79 185
R88 drain_right.n129 drain_right.n128 185
R89 drain_right.n127 drain_right.n126 185
R90 drain_right.n84 drain_right.n83 185
R91 drain_right.n121 drain_right.n120 185
R92 drain_right.n119 drain_right.n86 185
R93 drain_right.n118 drain_right.n117 185
R94 drain_right.n89 drain_right.n87 185
R95 drain_right.n112 drain_right.n111 185
R96 drain_right.n110 drain_right.n109 185
R97 drain_right.n93 drain_right.n92 185
R98 drain_right.n104 drain_right.n103 185
R99 drain_right.n102 drain_right.n101 185
R100 drain_right.n97 drain_right.n96 185
R101 drain_right.n21 drain_right.t11 149.524
R102 drain_right.n98 drain_right.t3 149.524
R103 drain_right.n25 drain_right.n19 104.615
R104 drain_right.n26 drain_right.n25 104.615
R105 drain_right.n26 drain_right.n15 104.615
R106 drain_right.n33 drain_right.n15 104.615
R107 drain_right.n34 drain_right.n33 104.615
R108 drain_right.n34 drain_right.n11 104.615
R109 drain_right.n42 drain_right.n11 104.615
R110 drain_right.n43 drain_right.n42 104.615
R111 drain_right.n44 drain_right.n43 104.615
R112 drain_right.n44 drain_right.n7 104.615
R113 drain_right.n51 drain_right.n7 104.615
R114 drain_right.n52 drain_right.n51 104.615
R115 drain_right.n52 drain_right.n3 104.615
R116 drain_right.n59 drain_right.n3 104.615
R117 drain_right.n60 drain_right.n59 104.615
R118 drain_right.n136 drain_right.n135 104.615
R119 drain_right.n135 drain_right.n79 104.615
R120 drain_right.n128 drain_right.n79 104.615
R121 drain_right.n128 drain_right.n127 104.615
R122 drain_right.n127 drain_right.n83 104.615
R123 drain_right.n120 drain_right.n83 104.615
R124 drain_right.n120 drain_right.n119 104.615
R125 drain_right.n119 drain_right.n118 104.615
R126 drain_right.n118 drain_right.n87 104.615
R127 drain_right.n111 drain_right.n87 104.615
R128 drain_right.n111 drain_right.n110 104.615
R129 drain_right.n110 drain_right.n92 104.615
R130 drain_right.n103 drain_right.n92 104.615
R131 drain_right.n103 drain_right.n102 104.615
R132 drain_right.n102 drain_right.n96 104.615
R133 drain_right.n69 drain_right.n67 60.5266
R134 drain_right.n73 drain_right.n71 60.5266
R135 drain_right.n73 drain_right.n72 59.5527
R136 drain_right.n75 drain_right.n74 59.5527
R137 drain_right.n69 drain_right.n68 59.5525
R138 drain_right.n66 drain_right.n65 59.5525
R139 drain_right.t11 drain_right.n19 52.3082
R140 drain_right.t3 drain_right.n96 52.3082
R141 drain_right.n66 drain_right.n64 47.511
R142 drain_right.n141 drain_right.n140 46.5369
R143 drain_right drain_right.n70 32.4151
R144 drain_right.n45 drain_right.n10 13.1884
R145 drain_right.n121 drain_right.n86 13.1884
R146 drain_right.n41 drain_right.n40 12.8005
R147 drain_right.n46 drain_right.n8 12.8005
R148 drain_right.n122 drain_right.n84 12.8005
R149 drain_right.n117 drain_right.n88 12.8005
R150 drain_right.n39 drain_right.n12 12.0247
R151 drain_right.n50 drain_right.n49 12.0247
R152 drain_right.n126 drain_right.n125 12.0247
R153 drain_right.n116 drain_right.n89 12.0247
R154 drain_right.n36 drain_right.n35 11.249
R155 drain_right.n53 drain_right.n6 11.249
R156 drain_right.n129 drain_right.n82 11.249
R157 drain_right.n113 drain_right.n112 11.249
R158 drain_right.n32 drain_right.n14 10.4732
R159 drain_right.n54 drain_right.n4 10.4732
R160 drain_right.n130 drain_right.n80 10.4732
R161 drain_right.n109 drain_right.n91 10.4732
R162 drain_right.n21 drain_right.n20 10.2747
R163 drain_right.n98 drain_right.n97 10.2747
R164 drain_right.n31 drain_right.n16 9.69747
R165 drain_right.n58 drain_right.n57 9.69747
R166 drain_right.n134 drain_right.n133 9.69747
R167 drain_right.n108 drain_right.n93 9.69747
R168 drain_right.n64 drain_right.n63 9.45567
R169 drain_right.n140 drain_right.n139 9.45567
R170 drain_right.n63 drain_right.n62 9.3005
R171 drain_right.n2 drain_right.n1 9.3005
R172 drain_right.n57 drain_right.n56 9.3005
R173 drain_right.n55 drain_right.n54 9.3005
R174 drain_right.n6 drain_right.n5 9.3005
R175 drain_right.n49 drain_right.n48 9.3005
R176 drain_right.n47 drain_right.n46 9.3005
R177 drain_right.n23 drain_right.n22 9.3005
R178 drain_right.n18 drain_right.n17 9.3005
R179 drain_right.n29 drain_right.n28 9.3005
R180 drain_right.n31 drain_right.n30 9.3005
R181 drain_right.n14 drain_right.n13 9.3005
R182 drain_right.n37 drain_right.n36 9.3005
R183 drain_right.n39 drain_right.n38 9.3005
R184 drain_right.n40 drain_right.n9 9.3005
R185 drain_right.n100 drain_right.n99 9.3005
R186 drain_right.n95 drain_right.n94 9.3005
R187 drain_right.n106 drain_right.n105 9.3005
R188 drain_right.n108 drain_right.n107 9.3005
R189 drain_right.n91 drain_right.n90 9.3005
R190 drain_right.n114 drain_right.n113 9.3005
R191 drain_right.n116 drain_right.n115 9.3005
R192 drain_right.n88 drain_right.n85 9.3005
R193 drain_right.n139 drain_right.n138 9.3005
R194 drain_right.n78 drain_right.n77 9.3005
R195 drain_right.n133 drain_right.n132 9.3005
R196 drain_right.n131 drain_right.n130 9.3005
R197 drain_right.n82 drain_right.n81 9.3005
R198 drain_right.n125 drain_right.n124 9.3005
R199 drain_right.n123 drain_right.n122 9.3005
R200 drain_right.n28 drain_right.n27 8.92171
R201 drain_right.n61 drain_right.n2 8.92171
R202 drain_right.n137 drain_right.n78 8.92171
R203 drain_right.n105 drain_right.n104 8.92171
R204 drain_right.n24 drain_right.n18 8.14595
R205 drain_right.n62 drain_right.n0 8.14595
R206 drain_right.n138 drain_right.n76 8.14595
R207 drain_right.n101 drain_right.n95 8.14595
R208 drain_right.n23 drain_right.n20 7.3702
R209 drain_right.n100 drain_right.n97 7.3702
R210 drain_right drain_right.n141 6.14028
R211 drain_right.n24 drain_right.n23 5.81868
R212 drain_right.n64 drain_right.n0 5.81868
R213 drain_right.n140 drain_right.n76 5.81868
R214 drain_right.n101 drain_right.n100 5.81868
R215 drain_right.n27 drain_right.n18 5.04292
R216 drain_right.n62 drain_right.n61 5.04292
R217 drain_right.n138 drain_right.n137 5.04292
R218 drain_right.n104 drain_right.n95 5.04292
R219 drain_right.n28 drain_right.n16 4.26717
R220 drain_right.n58 drain_right.n2 4.26717
R221 drain_right.n134 drain_right.n78 4.26717
R222 drain_right.n105 drain_right.n93 4.26717
R223 drain_right.n32 drain_right.n31 3.49141
R224 drain_right.n57 drain_right.n4 3.49141
R225 drain_right.n133 drain_right.n80 3.49141
R226 drain_right.n109 drain_right.n108 3.49141
R227 drain_right.n22 drain_right.n21 2.84303
R228 drain_right.n99 drain_right.n98 2.84303
R229 drain_right.n35 drain_right.n14 2.71565
R230 drain_right.n54 drain_right.n53 2.71565
R231 drain_right.n130 drain_right.n129 2.71565
R232 drain_right.n112 drain_right.n91 2.71565
R233 drain_right.n36 drain_right.n12 1.93989
R234 drain_right.n50 drain_right.n6 1.93989
R235 drain_right.n126 drain_right.n82 1.93989
R236 drain_right.n113 drain_right.n89 1.93989
R237 drain_right.n67 drain_right.t8 1.6505
R238 drain_right.n67 drain_right.t4 1.6505
R239 drain_right.n68 drain_right.t9 1.6505
R240 drain_right.n68 drain_right.t12 1.6505
R241 drain_right.n65 drain_right.t0 1.6505
R242 drain_right.n65 drain_right.t13 1.6505
R243 drain_right.n71 drain_right.t7 1.6505
R244 drain_right.n71 drain_right.t2 1.6505
R245 drain_right.n72 drain_right.t10 1.6505
R246 drain_right.n72 drain_right.t6 1.6505
R247 drain_right.n74 drain_right.t1 1.6505
R248 drain_right.n74 drain_right.t5 1.6505
R249 drain_right.n41 drain_right.n39 1.16414
R250 drain_right.n49 drain_right.n8 1.16414
R251 drain_right.n125 drain_right.n84 1.16414
R252 drain_right.n117 drain_right.n116 1.16414
R253 drain_right.n141 drain_right.n75 0.974638
R254 drain_right.n75 drain_right.n73 0.974638
R255 drain_right.n70 drain_right.n66 0.675757
R256 drain_right.n40 drain_right.n10 0.388379
R257 drain_right.n46 drain_right.n45 0.388379
R258 drain_right.n122 drain_right.n121 0.388379
R259 drain_right.n88 drain_right.n86 0.388379
R260 drain_right.n70 drain_right.n69 0.188688
R261 drain_right.n22 drain_right.n17 0.155672
R262 drain_right.n29 drain_right.n17 0.155672
R263 drain_right.n30 drain_right.n29 0.155672
R264 drain_right.n30 drain_right.n13 0.155672
R265 drain_right.n37 drain_right.n13 0.155672
R266 drain_right.n38 drain_right.n37 0.155672
R267 drain_right.n38 drain_right.n9 0.155672
R268 drain_right.n47 drain_right.n9 0.155672
R269 drain_right.n48 drain_right.n47 0.155672
R270 drain_right.n48 drain_right.n5 0.155672
R271 drain_right.n55 drain_right.n5 0.155672
R272 drain_right.n56 drain_right.n55 0.155672
R273 drain_right.n56 drain_right.n1 0.155672
R274 drain_right.n63 drain_right.n1 0.155672
R275 drain_right.n139 drain_right.n77 0.155672
R276 drain_right.n132 drain_right.n77 0.155672
R277 drain_right.n132 drain_right.n131 0.155672
R278 drain_right.n131 drain_right.n81 0.155672
R279 drain_right.n124 drain_right.n81 0.155672
R280 drain_right.n124 drain_right.n123 0.155672
R281 drain_right.n123 drain_right.n85 0.155672
R282 drain_right.n115 drain_right.n85 0.155672
R283 drain_right.n115 drain_right.n114 0.155672
R284 drain_right.n114 drain_right.n90 0.155672
R285 drain_right.n107 drain_right.n90 0.155672
R286 drain_right.n107 drain_right.n106 0.155672
R287 drain_right.n106 drain_right.n94 0.155672
R288 drain_right.n99 drain_right.n94 0.155672
R289 source.n282 source.n222 289.615
R290 source.n210 source.n150 289.615
R291 source.n60 source.n0 289.615
R292 source.n132 source.n72 289.615
R293 source.n242 source.n241 185
R294 source.n247 source.n246 185
R295 source.n249 source.n248 185
R296 source.n238 source.n237 185
R297 source.n255 source.n254 185
R298 source.n257 source.n256 185
R299 source.n234 source.n233 185
R300 source.n264 source.n263 185
R301 source.n265 source.n232 185
R302 source.n267 source.n266 185
R303 source.n230 source.n229 185
R304 source.n273 source.n272 185
R305 source.n275 source.n274 185
R306 source.n226 source.n225 185
R307 source.n281 source.n280 185
R308 source.n283 source.n282 185
R309 source.n170 source.n169 185
R310 source.n175 source.n174 185
R311 source.n177 source.n176 185
R312 source.n166 source.n165 185
R313 source.n183 source.n182 185
R314 source.n185 source.n184 185
R315 source.n162 source.n161 185
R316 source.n192 source.n191 185
R317 source.n193 source.n160 185
R318 source.n195 source.n194 185
R319 source.n158 source.n157 185
R320 source.n201 source.n200 185
R321 source.n203 source.n202 185
R322 source.n154 source.n153 185
R323 source.n209 source.n208 185
R324 source.n211 source.n210 185
R325 source.n61 source.n60 185
R326 source.n59 source.n58 185
R327 source.n4 source.n3 185
R328 source.n53 source.n52 185
R329 source.n51 source.n50 185
R330 source.n8 source.n7 185
R331 source.n45 source.n44 185
R332 source.n43 source.n10 185
R333 source.n42 source.n41 185
R334 source.n13 source.n11 185
R335 source.n36 source.n35 185
R336 source.n34 source.n33 185
R337 source.n17 source.n16 185
R338 source.n28 source.n27 185
R339 source.n26 source.n25 185
R340 source.n21 source.n20 185
R341 source.n133 source.n132 185
R342 source.n131 source.n130 185
R343 source.n76 source.n75 185
R344 source.n125 source.n124 185
R345 source.n123 source.n122 185
R346 source.n80 source.n79 185
R347 source.n117 source.n116 185
R348 source.n115 source.n82 185
R349 source.n114 source.n113 185
R350 source.n85 source.n83 185
R351 source.n108 source.n107 185
R352 source.n106 source.n105 185
R353 source.n89 source.n88 185
R354 source.n100 source.n99 185
R355 source.n98 source.n97 185
R356 source.n93 source.n92 185
R357 source.n243 source.t16 149.524
R358 source.n171 source.t6 149.524
R359 source.n22 source.t8 149.524
R360 source.n94 source.t20 149.524
R361 source.n247 source.n241 104.615
R362 source.n248 source.n247 104.615
R363 source.n248 source.n237 104.615
R364 source.n255 source.n237 104.615
R365 source.n256 source.n255 104.615
R366 source.n256 source.n233 104.615
R367 source.n264 source.n233 104.615
R368 source.n265 source.n264 104.615
R369 source.n266 source.n265 104.615
R370 source.n266 source.n229 104.615
R371 source.n273 source.n229 104.615
R372 source.n274 source.n273 104.615
R373 source.n274 source.n225 104.615
R374 source.n281 source.n225 104.615
R375 source.n282 source.n281 104.615
R376 source.n175 source.n169 104.615
R377 source.n176 source.n175 104.615
R378 source.n176 source.n165 104.615
R379 source.n183 source.n165 104.615
R380 source.n184 source.n183 104.615
R381 source.n184 source.n161 104.615
R382 source.n192 source.n161 104.615
R383 source.n193 source.n192 104.615
R384 source.n194 source.n193 104.615
R385 source.n194 source.n157 104.615
R386 source.n201 source.n157 104.615
R387 source.n202 source.n201 104.615
R388 source.n202 source.n153 104.615
R389 source.n209 source.n153 104.615
R390 source.n210 source.n209 104.615
R391 source.n60 source.n59 104.615
R392 source.n59 source.n3 104.615
R393 source.n52 source.n3 104.615
R394 source.n52 source.n51 104.615
R395 source.n51 source.n7 104.615
R396 source.n44 source.n7 104.615
R397 source.n44 source.n43 104.615
R398 source.n43 source.n42 104.615
R399 source.n42 source.n11 104.615
R400 source.n35 source.n11 104.615
R401 source.n35 source.n34 104.615
R402 source.n34 source.n16 104.615
R403 source.n27 source.n16 104.615
R404 source.n27 source.n26 104.615
R405 source.n26 source.n20 104.615
R406 source.n132 source.n131 104.615
R407 source.n131 source.n75 104.615
R408 source.n124 source.n75 104.615
R409 source.n124 source.n123 104.615
R410 source.n123 source.n79 104.615
R411 source.n116 source.n79 104.615
R412 source.n116 source.n115 104.615
R413 source.n115 source.n114 104.615
R414 source.n114 source.n83 104.615
R415 source.n107 source.n83 104.615
R416 source.n107 source.n106 104.615
R417 source.n106 source.n88 104.615
R418 source.n99 source.n88 104.615
R419 source.n99 source.n98 104.615
R420 source.n98 source.n92 104.615
R421 source.t16 source.n241 52.3082
R422 source.t6 source.n169 52.3082
R423 source.t8 source.n20 52.3082
R424 source.t20 source.n92 52.3082
R425 source.n67 source.n66 42.8739
R426 source.n69 source.n68 42.8739
R427 source.n71 source.n70 42.8739
R428 source.n139 source.n138 42.8739
R429 source.n141 source.n140 42.8739
R430 source.n143 source.n142 42.8739
R431 source.n221 source.n220 42.8737
R432 source.n219 source.n218 42.8737
R433 source.n217 source.n216 42.8737
R434 source.n149 source.n148 42.8737
R435 source.n147 source.n146 42.8737
R436 source.n145 source.n144 42.8737
R437 source.n287 source.n286 29.8581
R438 source.n215 source.n214 29.8581
R439 source.n65 source.n64 29.8581
R440 source.n137 source.n136 29.8581
R441 source.n145 source.n143 23.236
R442 source.n288 source.n65 16.5119
R443 source.n267 source.n232 13.1884
R444 source.n195 source.n160 13.1884
R445 source.n45 source.n10 13.1884
R446 source.n117 source.n82 13.1884
R447 source.n263 source.n262 12.8005
R448 source.n268 source.n230 12.8005
R449 source.n191 source.n190 12.8005
R450 source.n196 source.n158 12.8005
R451 source.n46 source.n8 12.8005
R452 source.n41 source.n12 12.8005
R453 source.n118 source.n80 12.8005
R454 source.n113 source.n84 12.8005
R455 source.n261 source.n234 12.0247
R456 source.n272 source.n271 12.0247
R457 source.n189 source.n162 12.0247
R458 source.n200 source.n199 12.0247
R459 source.n50 source.n49 12.0247
R460 source.n40 source.n13 12.0247
R461 source.n122 source.n121 12.0247
R462 source.n112 source.n85 12.0247
R463 source.n258 source.n257 11.249
R464 source.n275 source.n228 11.249
R465 source.n186 source.n185 11.249
R466 source.n203 source.n156 11.249
R467 source.n53 source.n6 11.249
R468 source.n37 source.n36 11.249
R469 source.n125 source.n78 11.249
R470 source.n109 source.n108 11.249
R471 source.n254 source.n236 10.4732
R472 source.n276 source.n226 10.4732
R473 source.n182 source.n164 10.4732
R474 source.n204 source.n154 10.4732
R475 source.n54 source.n4 10.4732
R476 source.n33 source.n15 10.4732
R477 source.n126 source.n76 10.4732
R478 source.n105 source.n87 10.4732
R479 source.n243 source.n242 10.2747
R480 source.n171 source.n170 10.2747
R481 source.n22 source.n21 10.2747
R482 source.n94 source.n93 10.2747
R483 source.n253 source.n238 9.69747
R484 source.n280 source.n279 9.69747
R485 source.n181 source.n166 9.69747
R486 source.n208 source.n207 9.69747
R487 source.n58 source.n57 9.69747
R488 source.n32 source.n17 9.69747
R489 source.n130 source.n129 9.69747
R490 source.n104 source.n89 9.69747
R491 source.n286 source.n285 9.45567
R492 source.n214 source.n213 9.45567
R493 source.n64 source.n63 9.45567
R494 source.n136 source.n135 9.45567
R495 source.n285 source.n284 9.3005
R496 source.n224 source.n223 9.3005
R497 source.n279 source.n278 9.3005
R498 source.n277 source.n276 9.3005
R499 source.n228 source.n227 9.3005
R500 source.n271 source.n270 9.3005
R501 source.n269 source.n268 9.3005
R502 source.n245 source.n244 9.3005
R503 source.n240 source.n239 9.3005
R504 source.n251 source.n250 9.3005
R505 source.n253 source.n252 9.3005
R506 source.n236 source.n235 9.3005
R507 source.n259 source.n258 9.3005
R508 source.n261 source.n260 9.3005
R509 source.n262 source.n231 9.3005
R510 source.n213 source.n212 9.3005
R511 source.n152 source.n151 9.3005
R512 source.n207 source.n206 9.3005
R513 source.n205 source.n204 9.3005
R514 source.n156 source.n155 9.3005
R515 source.n199 source.n198 9.3005
R516 source.n197 source.n196 9.3005
R517 source.n173 source.n172 9.3005
R518 source.n168 source.n167 9.3005
R519 source.n179 source.n178 9.3005
R520 source.n181 source.n180 9.3005
R521 source.n164 source.n163 9.3005
R522 source.n187 source.n186 9.3005
R523 source.n189 source.n188 9.3005
R524 source.n190 source.n159 9.3005
R525 source.n24 source.n23 9.3005
R526 source.n19 source.n18 9.3005
R527 source.n30 source.n29 9.3005
R528 source.n32 source.n31 9.3005
R529 source.n15 source.n14 9.3005
R530 source.n38 source.n37 9.3005
R531 source.n40 source.n39 9.3005
R532 source.n12 source.n9 9.3005
R533 source.n63 source.n62 9.3005
R534 source.n2 source.n1 9.3005
R535 source.n57 source.n56 9.3005
R536 source.n55 source.n54 9.3005
R537 source.n6 source.n5 9.3005
R538 source.n49 source.n48 9.3005
R539 source.n47 source.n46 9.3005
R540 source.n96 source.n95 9.3005
R541 source.n91 source.n90 9.3005
R542 source.n102 source.n101 9.3005
R543 source.n104 source.n103 9.3005
R544 source.n87 source.n86 9.3005
R545 source.n110 source.n109 9.3005
R546 source.n112 source.n111 9.3005
R547 source.n84 source.n81 9.3005
R548 source.n135 source.n134 9.3005
R549 source.n74 source.n73 9.3005
R550 source.n129 source.n128 9.3005
R551 source.n127 source.n126 9.3005
R552 source.n78 source.n77 9.3005
R553 source.n121 source.n120 9.3005
R554 source.n119 source.n118 9.3005
R555 source.n250 source.n249 8.92171
R556 source.n283 source.n224 8.92171
R557 source.n178 source.n177 8.92171
R558 source.n211 source.n152 8.92171
R559 source.n61 source.n2 8.92171
R560 source.n29 source.n28 8.92171
R561 source.n133 source.n74 8.92171
R562 source.n101 source.n100 8.92171
R563 source.n246 source.n240 8.14595
R564 source.n284 source.n222 8.14595
R565 source.n174 source.n168 8.14595
R566 source.n212 source.n150 8.14595
R567 source.n62 source.n0 8.14595
R568 source.n25 source.n19 8.14595
R569 source.n134 source.n72 8.14595
R570 source.n97 source.n91 8.14595
R571 source.n245 source.n242 7.3702
R572 source.n173 source.n170 7.3702
R573 source.n24 source.n21 7.3702
R574 source.n96 source.n93 7.3702
R575 source.n246 source.n245 5.81868
R576 source.n286 source.n222 5.81868
R577 source.n174 source.n173 5.81868
R578 source.n214 source.n150 5.81868
R579 source.n64 source.n0 5.81868
R580 source.n25 source.n24 5.81868
R581 source.n136 source.n72 5.81868
R582 source.n97 source.n96 5.81868
R583 source.n288 source.n287 5.7505
R584 source.n249 source.n240 5.04292
R585 source.n284 source.n283 5.04292
R586 source.n177 source.n168 5.04292
R587 source.n212 source.n211 5.04292
R588 source.n62 source.n61 5.04292
R589 source.n28 source.n19 5.04292
R590 source.n134 source.n133 5.04292
R591 source.n100 source.n91 5.04292
R592 source.n250 source.n238 4.26717
R593 source.n280 source.n224 4.26717
R594 source.n178 source.n166 4.26717
R595 source.n208 source.n152 4.26717
R596 source.n58 source.n2 4.26717
R597 source.n29 source.n17 4.26717
R598 source.n130 source.n74 4.26717
R599 source.n101 source.n89 4.26717
R600 source.n254 source.n253 3.49141
R601 source.n279 source.n226 3.49141
R602 source.n182 source.n181 3.49141
R603 source.n207 source.n154 3.49141
R604 source.n57 source.n4 3.49141
R605 source.n33 source.n32 3.49141
R606 source.n129 source.n76 3.49141
R607 source.n105 source.n104 3.49141
R608 source.n244 source.n243 2.84303
R609 source.n172 source.n171 2.84303
R610 source.n23 source.n22 2.84303
R611 source.n95 source.n94 2.84303
R612 source.n257 source.n236 2.71565
R613 source.n276 source.n275 2.71565
R614 source.n185 source.n164 2.71565
R615 source.n204 source.n203 2.71565
R616 source.n54 source.n53 2.71565
R617 source.n36 source.n15 2.71565
R618 source.n126 source.n125 2.71565
R619 source.n108 source.n87 2.71565
R620 source.n258 source.n234 1.93989
R621 source.n272 source.n228 1.93989
R622 source.n186 source.n162 1.93989
R623 source.n200 source.n156 1.93989
R624 source.n50 source.n6 1.93989
R625 source.n37 source.n13 1.93989
R626 source.n122 source.n78 1.93989
R627 source.n109 source.n85 1.93989
R628 source.n220 source.t14 1.6505
R629 source.n220 source.t26 1.6505
R630 source.n218 source.t15 1.6505
R631 source.n218 source.t25 1.6505
R632 source.n216 source.t13 1.6505
R633 source.n216 source.t24 1.6505
R634 source.n148 source.t4 1.6505
R635 source.n148 source.t7 1.6505
R636 source.n146 source.t12 1.6505
R637 source.n146 source.t0 1.6505
R638 source.n144 source.t5 1.6505
R639 source.n144 source.t1 1.6505
R640 source.n66 source.t27 1.6505
R641 source.n66 source.t11 1.6505
R642 source.n68 source.t3 1.6505
R643 source.n68 source.t10 1.6505
R644 source.n70 source.t9 1.6505
R645 source.n70 source.t2 1.6505
R646 source.n138 source.t23 1.6505
R647 source.n138 source.t22 1.6505
R648 source.n140 source.t17 1.6505
R649 source.n140 source.t18 1.6505
R650 source.n142 source.t21 1.6505
R651 source.n142 source.t19 1.6505
R652 source.n263 source.n261 1.16414
R653 source.n271 source.n230 1.16414
R654 source.n191 source.n189 1.16414
R655 source.n199 source.n158 1.16414
R656 source.n49 source.n8 1.16414
R657 source.n41 source.n40 1.16414
R658 source.n121 source.n80 1.16414
R659 source.n113 source.n112 1.16414
R660 source.n143 source.n141 0.974638
R661 source.n141 source.n139 0.974638
R662 source.n139 source.n137 0.974638
R663 source.n71 source.n69 0.974638
R664 source.n69 source.n67 0.974638
R665 source.n67 source.n65 0.974638
R666 source.n147 source.n145 0.974638
R667 source.n149 source.n147 0.974638
R668 source.n215 source.n149 0.974638
R669 source.n219 source.n217 0.974638
R670 source.n221 source.n219 0.974638
R671 source.n287 source.n221 0.974638
R672 source.n137 source.n71 0.957397
R673 source.n217 source.n215 0.957397
R674 source.n262 source.n232 0.388379
R675 source.n268 source.n267 0.388379
R676 source.n190 source.n160 0.388379
R677 source.n196 source.n195 0.388379
R678 source.n46 source.n45 0.388379
R679 source.n12 source.n10 0.388379
R680 source.n118 source.n117 0.388379
R681 source.n84 source.n82 0.388379
R682 source source.n288 0.188
R683 source.n244 source.n239 0.155672
R684 source.n251 source.n239 0.155672
R685 source.n252 source.n251 0.155672
R686 source.n252 source.n235 0.155672
R687 source.n259 source.n235 0.155672
R688 source.n260 source.n259 0.155672
R689 source.n260 source.n231 0.155672
R690 source.n269 source.n231 0.155672
R691 source.n270 source.n269 0.155672
R692 source.n270 source.n227 0.155672
R693 source.n277 source.n227 0.155672
R694 source.n278 source.n277 0.155672
R695 source.n278 source.n223 0.155672
R696 source.n285 source.n223 0.155672
R697 source.n172 source.n167 0.155672
R698 source.n179 source.n167 0.155672
R699 source.n180 source.n179 0.155672
R700 source.n180 source.n163 0.155672
R701 source.n187 source.n163 0.155672
R702 source.n188 source.n187 0.155672
R703 source.n188 source.n159 0.155672
R704 source.n197 source.n159 0.155672
R705 source.n198 source.n197 0.155672
R706 source.n198 source.n155 0.155672
R707 source.n205 source.n155 0.155672
R708 source.n206 source.n205 0.155672
R709 source.n206 source.n151 0.155672
R710 source.n213 source.n151 0.155672
R711 source.n63 source.n1 0.155672
R712 source.n56 source.n1 0.155672
R713 source.n56 source.n55 0.155672
R714 source.n55 source.n5 0.155672
R715 source.n48 source.n5 0.155672
R716 source.n48 source.n47 0.155672
R717 source.n47 source.n9 0.155672
R718 source.n39 source.n9 0.155672
R719 source.n39 source.n38 0.155672
R720 source.n38 source.n14 0.155672
R721 source.n31 source.n14 0.155672
R722 source.n31 source.n30 0.155672
R723 source.n30 source.n18 0.155672
R724 source.n23 source.n18 0.155672
R725 source.n135 source.n73 0.155672
R726 source.n128 source.n73 0.155672
R727 source.n128 source.n127 0.155672
R728 source.n127 source.n77 0.155672
R729 source.n120 source.n77 0.155672
R730 source.n120 source.n119 0.155672
R731 source.n119 source.n81 0.155672
R732 source.n111 source.n81 0.155672
R733 source.n111 source.n110 0.155672
R734 source.n110 source.n86 0.155672
R735 source.n103 source.n86 0.155672
R736 source.n103 source.n102 0.155672
R737 source.n102 source.n90 0.155672
R738 source.n95 source.n90 0.155672
R739 plus.n5 plus.t12 434.45
R740 plus.n23 plus.t9 434.45
R741 plus.n16 plus.t5 410.604
R742 plus.n14 plus.t6 410.604
R743 plus.n2 plus.t10 410.604
R744 plus.n9 plus.t7 410.604
R745 plus.n8 plus.t8 410.604
R746 plus.n4 plus.t11 410.604
R747 plus.n34 plus.t2 410.604
R748 plus.n32 plus.t13 410.604
R749 plus.n20 plus.t3 410.604
R750 plus.n27 plus.t0 410.604
R751 plus.n26 plus.t4 410.604
R752 plus.n22 plus.t1 410.604
R753 plus.n7 plus.n6 161.3
R754 plus.n13 plus.n12 161.3
R755 plus.n14 plus.n1 161.3
R756 plus.n15 plus.n0 161.3
R757 plus.n17 plus.n16 161.3
R758 plus.n25 plus.n24 161.3
R759 plus.n31 plus.n30 161.3
R760 plus.n32 plus.n19 161.3
R761 plus.n33 plus.n18 161.3
R762 plus.n35 plus.n34 161.3
R763 plus.n8 plus.n3 80.6037
R764 plus.n10 plus.n9 80.6037
R765 plus.n11 plus.n2 80.6037
R766 plus.n26 plus.n21 80.6037
R767 plus.n28 plus.n27 80.6037
R768 plus.n29 plus.n20 80.6037
R769 plus.n9 plus.n2 48.2005
R770 plus.n9 plus.n8 48.2005
R771 plus.n27 plus.n20 48.2005
R772 plus.n27 plus.n26 48.2005
R773 plus.n24 plus.n23 44.9119
R774 plus.n6 plus.n5 44.9119
R775 plus.n16 plus.n15 35.055
R776 plus.n34 plus.n33 35.055
R777 plus plus.n35 32.7888
R778 plus.n13 plus.n2 32.1338
R779 plus.n8 plus.n7 32.1338
R780 plus.n31 plus.n20 32.1338
R781 plus.n26 plus.n25 32.1338
R782 plus.n23 plus.n22 17.739
R783 plus.n5 plus.n4 17.739
R784 plus.n14 plus.n13 16.0672
R785 plus.n7 plus.n4 16.0672
R786 plus.n32 plus.n31 16.0672
R787 plus.n25 plus.n22 16.0672
R788 plus.n15 plus.n14 13.146
R789 plus.n33 plus.n32 13.146
R790 plus plus.n17 12.3698
R791 plus.n10 plus.n3 0.380177
R792 plus.n11 plus.n10 0.380177
R793 plus.n29 plus.n28 0.380177
R794 plus.n28 plus.n21 0.380177
R795 plus.n6 plus.n3 0.285035
R796 plus.n12 plus.n11 0.285035
R797 plus.n30 plus.n29 0.285035
R798 plus.n24 plus.n21 0.285035
R799 plus.n12 plus.n1 0.189894
R800 plus.n1 plus.n0 0.189894
R801 plus.n17 plus.n0 0.189894
R802 plus.n35 plus.n18 0.189894
R803 plus.n19 plus.n18 0.189894
R804 plus.n30 plus.n19 0.189894
R805 drain_left.n60 drain_left.n0 289.615
R806 drain_left.n131 drain_left.n71 289.615
R807 drain_left.n20 drain_left.n19 185
R808 drain_left.n25 drain_left.n24 185
R809 drain_left.n27 drain_left.n26 185
R810 drain_left.n16 drain_left.n15 185
R811 drain_left.n33 drain_left.n32 185
R812 drain_left.n35 drain_left.n34 185
R813 drain_left.n12 drain_left.n11 185
R814 drain_left.n42 drain_left.n41 185
R815 drain_left.n43 drain_left.n10 185
R816 drain_left.n45 drain_left.n44 185
R817 drain_left.n8 drain_left.n7 185
R818 drain_left.n51 drain_left.n50 185
R819 drain_left.n53 drain_left.n52 185
R820 drain_left.n4 drain_left.n3 185
R821 drain_left.n59 drain_left.n58 185
R822 drain_left.n61 drain_left.n60 185
R823 drain_left.n132 drain_left.n131 185
R824 drain_left.n130 drain_left.n129 185
R825 drain_left.n75 drain_left.n74 185
R826 drain_left.n124 drain_left.n123 185
R827 drain_left.n122 drain_left.n121 185
R828 drain_left.n79 drain_left.n78 185
R829 drain_left.n116 drain_left.n115 185
R830 drain_left.n114 drain_left.n81 185
R831 drain_left.n113 drain_left.n112 185
R832 drain_left.n84 drain_left.n82 185
R833 drain_left.n107 drain_left.n106 185
R834 drain_left.n105 drain_left.n104 185
R835 drain_left.n88 drain_left.n87 185
R836 drain_left.n99 drain_left.n98 185
R837 drain_left.n97 drain_left.n96 185
R838 drain_left.n92 drain_left.n91 185
R839 drain_left.n21 drain_left.t11 149.524
R840 drain_left.n93 drain_left.t1 149.524
R841 drain_left.n25 drain_left.n19 104.615
R842 drain_left.n26 drain_left.n25 104.615
R843 drain_left.n26 drain_left.n15 104.615
R844 drain_left.n33 drain_left.n15 104.615
R845 drain_left.n34 drain_left.n33 104.615
R846 drain_left.n34 drain_left.n11 104.615
R847 drain_left.n42 drain_left.n11 104.615
R848 drain_left.n43 drain_left.n42 104.615
R849 drain_left.n44 drain_left.n43 104.615
R850 drain_left.n44 drain_left.n7 104.615
R851 drain_left.n51 drain_left.n7 104.615
R852 drain_left.n52 drain_left.n51 104.615
R853 drain_left.n52 drain_left.n3 104.615
R854 drain_left.n59 drain_left.n3 104.615
R855 drain_left.n60 drain_left.n59 104.615
R856 drain_left.n131 drain_left.n130 104.615
R857 drain_left.n130 drain_left.n74 104.615
R858 drain_left.n123 drain_left.n74 104.615
R859 drain_left.n123 drain_left.n122 104.615
R860 drain_left.n122 drain_left.n78 104.615
R861 drain_left.n115 drain_left.n78 104.615
R862 drain_left.n115 drain_left.n114 104.615
R863 drain_left.n114 drain_left.n113 104.615
R864 drain_left.n113 drain_left.n82 104.615
R865 drain_left.n106 drain_left.n82 104.615
R866 drain_left.n106 drain_left.n105 104.615
R867 drain_left.n105 drain_left.n87 104.615
R868 drain_left.n98 drain_left.n87 104.615
R869 drain_left.n98 drain_left.n97 104.615
R870 drain_left.n97 drain_left.n91 104.615
R871 drain_left.n69 drain_left.n67 60.5266
R872 drain_left.n139 drain_left.n138 59.5527
R873 drain_left.n137 drain_left.n136 59.5527
R874 drain_left.n69 drain_left.n68 59.5525
R875 drain_left.n66 drain_left.n65 59.5525
R876 drain_left.n141 drain_left.n140 59.5525
R877 drain_left.t11 drain_left.n19 52.3082
R878 drain_left.t1 drain_left.n91 52.3082
R879 drain_left.n66 drain_left.n64 47.511
R880 drain_left.n137 drain_left.n135 47.511
R881 drain_left drain_left.n70 32.9684
R882 drain_left.n45 drain_left.n10 13.1884
R883 drain_left.n116 drain_left.n81 13.1884
R884 drain_left.n41 drain_left.n40 12.8005
R885 drain_left.n46 drain_left.n8 12.8005
R886 drain_left.n117 drain_left.n79 12.8005
R887 drain_left.n112 drain_left.n83 12.8005
R888 drain_left.n39 drain_left.n12 12.0247
R889 drain_left.n50 drain_left.n49 12.0247
R890 drain_left.n121 drain_left.n120 12.0247
R891 drain_left.n111 drain_left.n84 12.0247
R892 drain_left.n36 drain_left.n35 11.249
R893 drain_left.n53 drain_left.n6 11.249
R894 drain_left.n124 drain_left.n77 11.249
R895 drain_left.n108 drain_left.n107 11.249
R896 drain_left.n32 drain_left.n14 10.4732
R897 drain_left.n54 drain_left.n4 10.4732
R898 drain_left.n125 drain_left.n75 10.4732
R899 drain_left.n104 drain_left.n86 10.4732
R900 drain_left.n21 drain_left.n20 10.2747
R901 drain_left.n93 drain_left.n92 10.2747
R902 drain_left.n31 drain_left.n16 9.69747
R903 drain_left.n58 drain_left.n57 9.69747
R904 drain_left.n129 drain_left.n128 9.69747
R905 drain_left.n103 drain_left.n88 9.69747
R906 drain_left.n64 drain_left.n63 9.45567
R907 drain_left.n135 drain_left.n134 9.45567
R908 drain_left.n63 drain_left.n62 9.3005
R909 drain_left.n2 drain_left.n1 9.3005
R910 drain_left.n57 drain_left.n56 9.3005
R911 drain_left.n55 drain_left.n54 9.3005
R912 drain_left.n6 drain_left.n5 9.3005
R913 drain_left.n49 drain_left.n48 9.3005
R914 drain_left.n47 drain_left.n46 9.3005
R915 drain_left.n23 drain_left.n22 9.3005
R916 drain_left.n18 drain_left.n17 9.3005
R917 drain_left.n29 drain_left.n28 9.3005
R918 drain_left.n31 drain_left.n30 9.3005
R919 drain_left.n14 drain_left.n13 9.3005
R920 drain_left.n37 drain_left.n36 9.3005
R921 drain_left.n39 drain_left.n38 9.3005
R922 drain_left.n40 drain_left.n9 9.3005
R923 drain_left.n95 drain_left.n94 9.3005
R924 drain_left.n90 drain_left.n89 9.3005
R925 drain_left.n101 drain_left.n100 9.3005
R926 drain_left.n103 drain_left.n102 9.3005
R927 drain_left.n86 drain_left.n85 9.3005
R928 drain_left.n109 drain_left.n108 9.3005
R929 drain_left.n111 drain_left.n110 9.3005
R930 drain_left.n83 drain_left.n80 9.3005
R931 drain_left.n134 drain_left.n133 9.3005
R932 drain_left.n73 drain_left.n72 9.3005
R933 drain_left.n128 drain_left.n127 9.3005
R934 drain_left.n126 drain_left.n125 9.3005
R935 drain_left.n77 drain_left.n76 9.3005
R936 drain_left.n120 drain_left.n119 9.3005
R937 drain_left.n118 drain_left.n117 9.3005
R938 drain_left.n28 drain_left.n27 8.92171
R939 drain_left.n61 drain_left.n2 8.92171
R940 drain_left.n132 drain_left.n73 8.92171
R941 drain_left.n100 drain_left.n99 8.92171
R942 drain_left.n24 drain_left.n18 8.14595
R943 drain_left.n62 drain_left.n0 8.14595
R944 drain_left.n133 drain_left.n71 8.14595
R945 drain_left.n96 drain_left.n90 8.14595
R946 drain_left.n23 drain_left.n20 7.3702
R947 drain_left.n95 drain_left.n92 7.3702
R948 drain_left drain_left.n141 6.62735
R949 drain_left.n24 drain_left.n23 5.81868
R950 drain_left.n64 drain_left.n0 5.81868
R951 drain_left.n135 drain_left.n71 5.81868
R952 drain_left.n96 drain_left.n95 5.81868
R953 drain_left.n27 drain_left.n18 5.04292
R954 drain_left.n62 drain_left.n61 5.04292
R955 drain_left.n133 drain_left.n132 5.04292
R956 drain_left.n99 drain_left.n90 5.04292
R957 drain_left.n28 drain_left.n16 4.26717
R958 drain_left.n58 drain_left.n2 4.26717
R959 drain_left.n129 drain_left.n73 4.26717
R960 drain_left.n100 drain_left.n88 4.26717
R961 drain_left.n32 drain_left.n31 3.49141
R962 drain_left.n57 drain_left.n4 3.49141
R963 drain_left.n128 drain_left.n75 3.49141
R964 drain_left.n104 drain_left.n103 3.49141
R965 drain_left.n22 drain_left.n21 2.84303
R966 drain_left.n94 drain_left.n93 2.84303
R967 drain_left.n35 drain_left.n14 2.71565
R968 drain_left.n54 drain_left.n53 2.71565
R969 drain_left.n125 drain_left.n124 2.71565
R970 drain_left.n107 drain_left.n86 2.71565
R971 drain_left.n36 drain_left.n12 1.93989
R972 drain_left.n50 drain_left.n6 1.93989
R973 drain_left.n121 drain_left.n77 1.93989
R974 drain_left.n108 drain_left.n84 1.93989
R975 drain_left.n67 drain_left.t12 1.6505
R976 drain_left.n67 drain_left.t4 1.6505
R977 drain_left.n68 drain_left.t13 1.6505
R978 drain_left.n68 drain_left.t9 1.6505
R979 drain_left.n65 drain_left.t0 1.6505
R980 drain_left.n65 drain_left.t10 1.6505
R981 drain_left.n140 drain_left.t7 1.6505
R982 drain_left.n140 drain_left.t8 1.6505
R983 drain_left.n138 drain_left.t6 1.6505
R984 drain_left.n138 drain_left.t3 1.6505
R985 drain_left.n136 drain_left.t2 1.6505
R986 drain_left.n136 drain_left.t5 1.6505
R987 drain_left.n41 drain_left.n39 1.16414
R988 drain_left.n49 drain_left.n8 1.16414
R989 drain_left.n120 drain_left.n79 1.16414
R990 drain_left.n112 drain_left.n111 1.16414
R991 drain_left.n139 drain_left.n137 0.974638
R992 drain_left.n141 drain_left.n139 0.974638
R993 drain_left.n70 drain_left.n66 0.675757
R994 drain_left.n40 drain_left.n10 0.388379
R995 drain_left.n46 drain_left.n45 0.388379
R996 drain_left.n117 drain_left.n116 0.388379
R997 drain_left.n83 drain_left.n81 0.388379
R998 drain_left.n70 drain_left.n69 0.188688
R999 drain_left.n22 drain_left.n17 0.155672
R1000 drain_left.n29 drain_left.n17 0.155672
R1001 drain_left.n30 drain_left.n29 0.155672
R1002 drain_left.n30 drain_left.n13 0.155672
R1003 drain_left.n37 drain_left.n13 0.155672
R1004 drain_left.n38 drain_left.n37 0.155672
R1005 drain_left.n38 drain_left.n9 0.155672
R1006 drain_left.n47 drain_left.n9 0.155672
R1007 drain_left.n48 drain_left.n47 0.155672
R1008 drain_left.n48 drain_left.n5 0.155672
R1009 drain_left.n55 drain_left.n5 0.155672
R1010 drain_left.n56 drain_left.n55 0.155672
R1011 drain_left.n56 drain_left.n1 0.155672
R1012 drain_left.n63 drain_left.n1 0.155672
R1013 drain_left.n134 drain_left.n72 0.155672
R1014 drain_left.n127 drain_left.n72 0.155672
R1015 drain_left.n127 drain_left.n126 0.155672
R1016 drain_left.n126 drain_left.n76 0.155672
R1017 drain_left.n119 drain_left.n76 0.155672
R1018 drain_left.n119 drain_left.n118 0.155672
R1019 drain_left.n118 drain_left.n80 0.155672
R1020 drain_left.n110 drain_left.n80 0.155672
R1021 drain_left.n110 drain_left.n109 0.155672
R1022 drain_left.n109 drain_left.n85 0.155672
R1023 drain_left.n102 drain_left.n85 0.155672
R1024 drain_left.n102 drain_left.n101 0.155672
R1025 drain_left.n101 drain_left.n89 0.155672
R1026 drain_left.n94 drain_left.n89 0.155672
C0 plus source 9.76661f
C1 plus drain_right 0.408304f
C2 drain_left minus 0.173289f
C3 minus source 9.75211f
C4 minus drain_right 9.72201f
C5 drain_left source 17.5454f
C6 drain_left drain_right 1.31703f
C7 drain_right source 17.540098f
C8 plus minus 6.28665f
C9 drain_left plus 9.96961f
C10 drain_right a_n2524_n3288# 7.688139f
C11 drain_left a_n2524_n3288# 8.066219f
C12 source a_n2524_n3288# 6.807372f
C13 minus a_n2524_n3288# 10.034369f
C14 plus a_n2524_n3288# 11.719131f
C15 drain_left.n0 a_n2524_n3288# 0.032476f
C16 drain_left.n1 a_n2524_n3288# 0.024517f
C17 drain_left.n2 a_n2524_n3288# 0.013174f
C18 drain_left.n3 a_n2524_n3288# 0.031139f
C19 drain_left.n4 a_n2524_n3288# 0.013949f
C20 drain_left.n5 a_n2524_n3288# 0.024517f
C21 drain_left.n6 a_n2524_n3288# 0.013174f
C22 drain_left.n7 a_n2524_n3288# 0.031139f
C23 drain_left.n8 a_n2524_n3288# 0.013949f
C24 drain_left.n9 a_n2524_n3288# 0.024517f
C25 drain_left.n10 a_n2524_n3288# 0.013562f
C26 drain_left.n11 a_n2524_n3288# 0.031139f
C27 drain_left.n12 a_n2524_n3288# 0.013949f
C28 drain_left.n13 a_n2524_n3288# 0.024517f
C29 drain_left.n14 a_n2524_n3288# 0.013174f
C30 drain_left.n15 a_n2524_n3288# 0.031139f
C31 drain_left.n16 a_n2524_n3288# 0.013949f
C32 drain_left.n17 a_n2524_n3288# 0.024517f
C33 drain_left.n18 a_n2524_n3288# 0.013174f
C34 drain_left.n19 a_n2524_n3288# 0.023355f
C35 drain_left.n20 a_n2524_n3288# 0.022013f
C36 drain_left.t11 a_n2524_n3288# 0.052592f
C37 drain_left.n21 a_n2524_n3288# 0.176764f
C38 drain_left.n22 a_n2524_n3288# 1.23684f
C39 drain_left.n23 a_n2524_n3288# 0.013174f
C40 drain_left.n24 a_n2524_n3288# 0.013949f
C41 drain_left.n25 a_n2524_n3288# 0.031139f
C42 drain_left.n26 a_n2524_n3288# 0.031139f
C43 drain_left.n27 a_n2524_n3288# 0.013949f
C44 drain_left.n28 a_n2524_n3288# 0.013174f
C45 drain_left.n29 a_n2524_n3288# 0.024517f
C46 drain_left.n30 a_n2524_n3288# 0.024517f
C47 drain_left.n31 a_n2524_n3288# 0.013174f
C48 drain_left.n32 a_n2524_n3288# 0.013949f
C49 drain_left.n33 a_n2524_n3288# 0.031139f
C50 drain_left.n34 a_n2524_n3288# 0.031139f
C51 drain_left.n35 a_n2524_n3288# 0.013949f
C52 drain_left.n36 a_n2524_n3288# 0.013174f
C53 drain_left.n37 a_n2524_n3288# 0.024517f
C54 drain_left.n38 a_n2524_n3288# 0.024517f
C55 drain_left.n39 a_n2524_n3288# 0.013174f
C56 drain_left.n40 a_n2524_n3288# 0.013174f
C57 drain_left.n41 a_n2524_n3288# 0.013949f
C58 drain_left.n42 a_n2524_n3288# 0.031139f
C59 drain_left.n43 a_n2524_n3288# 0.031139f
C60 drain_left.n44 a_n2524_n3288# 0.031139f
C61 drain_left.n45 a_n2524_n3288# 0.013562f
C62 drain_left.n46 a_n2524_n3288# 0.013174f
C63 drain_left.n47 a_n2524_n3288# 0.024517f
C64 drain_left.n48 a_n2524_n3288# 0.024517f
C65 drain_left.n49 a_n2524_n3288# 0.013174f
C66 drain_left.n50 a_n2524_n3288# 0.013949f
C67 drain_left.n51 a_n2524_n3288# 0.031139f
C68 drain_left.n52 a_n2524_n3288# 0.031139f
C69 drain_left.n53 a_n2524_n3288# 0.013949f
C70 drain_left.n54 a_n2524_n3288# 0.013174f
C71 drain_left.n55 a_n2524_n3288# 0.024517f
C72 drain_left.n56 a_n2524_n3288# 0.024517f
C73 drain_left.n57 a_n2524_n3288# 0.013174f
C74 drain_left.n58 a_n2524_n3288# 0.013949f
C75 drain_left.n59 a_n2524_n3288# 0.031139f
C76 drain_left.n60 a_n2524_n3288# 0.063901f
C77 drain_left.n61 a_n2524_n3288# 0.013949f
C78 drain_left.n62 a_n2524_n3288# 0.013174f
C79 drain_left.n63 a_n2524_n3288# 0.052651f
C80 drain_left.n64 a_n2524_n3288# 0.054729f
C81 drain_left.t0 a_n2524_n3288# 0.232488f
C82 drain_left.t10 a_n2524_n3288# 0.232488f
C83 drain_left.n65 a_n2524_n3288# 2.06879f
C84 drain_left.n66 a_n2524_n3288# 0.45627f
C85 drain_left.t12 a_n2524_n3288# 0.232488f
C86 drain_left.t4 a_n2524_n3288# 0.232488f
C87 drain_left.n67 a_n2524_n3288# 2.07473f
C88 drain_left.t13 a_n2524_n3288# 0.232488f
C89 drain_left.t9 a_n2524_n3288# 0.232488f
C90 drain_left.n68 a_n2524_n3288# 2.06879f
C91 drain_left.n69 a_n2524_n3288# 0.664202f
C92 drain_left.n70 a_n2524_n3288# 1.40038f
C93 drain_left.n71 a_n2524_n3288# 0.032476f
C94 drain_left.n72 a_n2524_n3288# 0.024517f
C95 drain_left.n73 a_n2524_n3288# 0.013174f
C96 drain_left.n74 a_n2524_n3288# 0.031139f
C97 drain_left.n75 a_n2524_n3288# 0.013949f
C98 drain_left.n76 a_n2524_n3288# 0.024517f
C99 drain_left.n77 a_n2524_n3288# 0.013174f
C100 drain_left.n78 a_n2524_n3288# 0.031139f
C101 drain_left.n79 a_n2524_n3288# 0.013949f
C102 drain_left.n80 a_n2524_n3288# 0.024517f
C103 drain_left.n81 a_n2524_n3288# 0.013562f
C104 drain_left.n82 a_n2524_n3288# 0.031139f
C105 drain_left.n83 a_n2524_n3288# 0.013174f
C106 drain_left.n84 a_n2524_n3288# 0.013949f
C107 drain_left.n85 a_n2524_n3288# 0.024517f
C108 drain_left.n86 a_n2524_n3288# 0.013174f
C109 drain_left.n87 a_n2524_n3288# 0.031139f
C110 drain_left.n88 a_n2524_n3288# 0.013949f
C111 drain_left.n89 a_n2524_n3288# 0.024517f
C112 drain_left.n90 a_n2524_n3288# 0.013174f
C113 drain_left.n91 a_n2524_n3288# 0.023355f
C114 drain_left.n92 a_n2524_n3288# 0.022013f
C115 drain_left.t1 a_n2524_n3288# 0.052592f
C116 drain_left.n93 a_n2524_n3288# 0.176764f
C117 drain_left.n94 a_n2524_n3288# 1.23684f
C118 drain_left.n95 a_n2524_n3288# 0.013174f
C119 drain_left.n96 a_n2524_n3288# 0.013949f
C120 drain_left.n97 a_n2524_n3288# 0.031139f
C121 drain_left.n98 a_n2524_n3288# 0.031139f
C122 drain_left.n99 a_n2524_n3288# 0.013949f
C123 drain_left.n100 a_n2524_n3288# 0.013174f
C124 drain_left.n101 a_n2524_n3288# 0.024517f
C125 drain_left.n102 a_n2524_n3288# 0.024517f
C126 drain_left.n103 a_n2524_n3288# 0.013174f
C127 drain_left.n104 a_n2524_n3288# 0.013949f
C128 drain_left.n105 a_n2524_n3288# 0.031139f
C129 drain_left.n106 a_n2524_n3288# 0.031139f
C130 drain_left.n107 a_n2524_n3288# 0.013949f
C131 drain_left.n108 a_n2524_n3288# 0.013174f
C132 drain_left.n109 a_n2524_n3288# 0.024517f
C133 drain_left.n110 a_n2524_n3288# 0.024517f
C134 drain_left.n111 a_n2524_n3288# 0.013174f
C135 drain_left.n112 a_n2524_n3288# 0.013949f
C136 drain_left.n113 a_n2524_n3288# 0.031139f
C137 drain_left.n114 a_n2524_n3288# 0.031139f
C138 drain_left.n115 a_n2524_n3288# 0.031139f
C139 drain_left.n116 a_n2524_n3288# 0.013562f
C140 drain_left.n117 a_n2524_n3288# 0.013174f
C141 drain_left.n118 a_n2524_n3288# 0.024517f
C142 drain_left.n119 a_n2524_n3288# 0.024517f
C143 drain_left.n120 a_n2524_n3288# 0.013174f
C144 drain_left.n121 a_n2524_n3288# 0.013949f
C145 drain_left.n122 a_n2524_n3288# 0.031139f
C146 drain_left.n123 a_n2524_n3288# 0.031139f
C147 drain_left.n124 a_n2524_n3288# 0.013949f
C148 drain_left.n125 a_n2524_n3288# 0.013174f
C149 drain_left.n126 a_n2524_n3288# 0.024517f
C150 drain_left.n127 a_n2524_n3288# 0.024517f
C151 drain_left.n128 a_n2524_n3288# 0.013174f
C152 drain_left.n129 a_n2524_n3288# 0.013949f
C153 drain_left.n130 a_n2524_n3288# 0.031139f
C154 drain_left.n131 a_n2524_n3288# 0.063901f
C155 drain_left.n132 a_n2524_n3288# 0.013949f
C156 drain_left.n133 a_n2524_n3288# 0.013174f
C157 drain_left.n134 a_n2524_n3288# 0.052651f
C158 drain_left.n135 a_n2524_n3288# 0.054729f
C159 drain_left.t2 a_n2524_n3288# 0.232488f
C160 drain_left.t5 a_n2524_n3288# 0.232488f
C161 drain_left.n136 a_n2524_n3288# 2.0688f
C162 drain_left.n137 a_n2524_n3288# 0.479031f
C163 drain_left.t6 a_n2524_n3288# 0.232488f
C164 drain_left.t3 a_n2524_n3288# 0.232488f
C165 drain_left.n138 a_n2524_n3288# 2.0688f
C166 drain_left.n139 a_n2524_n3288# 0.359663f
C167 drain_left.t7 a_n2524_n3288# 0.232488f
C168 drain_left.t8 a_n2524_n3288# 0.232488f
C169 drain_left.n140 a_n2524_n3288# 2.06879f
C170 drain_left.n141 a_n2524_n3288# 0.579514f
C171 plus.n0 a_n2524_n3288# 0.039664f
C172 plus.t5 a_n2524_n3288# 1.08579f
C173 plus.t6 a_n2524_n3288# 1.08579f
C174 plus.n1 a_n2524_n3288# 0.039664f
C175 plus.t10 a_n2524_n3288# 1.08579f
C176 plus.n2 a_n2524_n3288# 0.438898f
C177 plus.n3 a_n2524_n3288# 0.066066f
C178 plus.t7 a_n2524_n3288# 1.08579f
C179 plus.t8 a_n2524_n3288# 1.08579f
C180 plus.t11 a_n2524_n3288# 1.08579f
C181 plus.n4 a_n2524_n3288# 0.434322f
C182 plus.t12 a_n2524_n3288# 1.1095f
C183 plus.n5 a_n2524_n3288# 0.411633f
C184 plus.n6 a_n2524_n3288# 0.185238f
C185 plus.n7 a_n2524_n3288# 0.009001f
C186 plus.n8 a_n2524_n3288# 0.438898f
C187 plus.n9 a_n2524_n3288# 0.441588f
C188 plus.n10 a_n2524_n3288# 0.079329f
C189 plus.n11 a_n2524_n3288# 0.066066f
C190 plus.n12 a_n2524_n3288# 0.052927f
C191 plus.n13 a_n2524_n3288# 0.009001f
C192 plus.n14 a_n2524_n3288# 0.429409f
C193 plus.n15 a_n2524_n3288# 0.009001f
C194 plus.n16 a_n2524_n3288# 0.430387f
C195 plus.n17 a_n2524_n3288# 0.465081f
C196 plus.n18 a_n2524_n3288# 0.039664f
C197 plus.t2 a_n2524_n3288# 1.08579f
C198 plus.n19 a_n2524_n3288# 0.039664f
C199 plus.t13 a_n2524_n3288# 1.08579f
C200 plus.t3 a_n2524_n3288# 1.08579f
C201 plus.n20 a_n2524_n3288# 0.438898f
C202 plus.n21 a_n2524_n3288# 0.066066f
C203 plus.t0 a_n2524_n3288# 1.08579f
C204 plus.t4 a_n2524_n3288# 1.08579f
C205 plus.t1 a_n2524_n3288# 1.08579f
C206 plus.n22 a_n2524_n3288# 0.434322f
C207 plus.t9 a_n2524_n3288# 1.1095f
C208 plus.n23 a_n2524_n3288# 0.411633f
C209 plus.n24 a_n2524_n3288# 0.185238f
C210 plus.n25 a_n2524_n3288# 0.009001f
C211 plus.n26 a_n2524_n3288# 0.438898f
C212 plus.n27 a_n2524_n3288# 0.441588f
C213 plus.n28 a_n2524_n3288# 0.079329f
C214 plus.n29 a_n2524_n3288# 0.066066f
C215 plus.n30 a_n2524_n3288# 0.052927f
C216 plus.n31 a_n2524_n3288# 0.009001f
C217 plus.n32 a_n2524_n3288# 0.429409f
C218 plus.n33 a_n2524_n3288# 0.009001f
C219 plus.n34 a_n2524_n3288# 0.430387f
C220 plus.n35 a_n2524_n3288# 1.34156f
C221 source.n0 a_n2524_n3288# 0.034287f
C222 source.n1 a_n2524_n3288# 0.025884f
C223 source.n2 a_n2524_n3288# 0.013909f
C224 source.n3 a_n2524_n3288# 0.032876f
C225 source.n4 a_n2524_n3288# 0.014727f
C226 source.n5 a_n2524_n3288# 0.025884f
C227 source.n6 a_n2524_n3288# 0.013909f
C228 source.n7 a_n2524_n3288# 0.032876f
C229 source.n8 a_n2524_n3288# 0.014727f
C230 source.n9 a_n2524_n3288# 0.025884f
C231 source.n10 a_n2524_n3288# 0.014318f
C232 source.n11 a_n2524_n3288# 0.032876f
C233 source.n12 a_n2524_n3288# 0.013909f
C234 source.n13 a_n2524_n3288# 0.014727f
C235 source.n14 a_n2524_n3288# 0.025884f
C236 source.n15 a_n2524_n3288# 0.013909f
C237 source.n16 a_n2524_n3288# 0.032876f
C238 source.n17 a_n2524_n3288# 0.014727f
C239 source.n18 a_n2524_n3288# 0.025884f
C240 source.n19 a_n2524_n3288# 0.013909f
C241 source.n20 a_n2524_n3288# 0.024657f
C242 source.n21 a_n2524_n3288# 0.023241f
C243 source.t8 a_n2524_n3288# 0.055525f
C244 source.n22 a_n2524_n3288# 0.186621f
C245 source.n23 a_n2524_n3288# 1.30581f
C246 source.n24 a_n2524_n3288# 0.013909f
C247 source.n25 a_n2524_n3288# 0.014727f
C248 source.n26 a_n2524_n3288# 0.032876f
C249 source.n27 a_n2524_n3288# 0.032876f
C250 source.n28 a_n2524_n3288# 0.014727f
C251 source.n29 a_n2524_n3288# 0.013909f
C252 source.n30 a_n2524_n3288# 0.025884f
C253 source.n31 a_n2524_n3288# 0.025884f
C254 source.n32 a_n2524_n3288# 0.013909f
C255 source.n33 a_n2524_n3288# 0.014727f
C256 source.n34 a_n2524_n3288# 0.032876f
C257 source.n35 a_n2524_n3288# 0.032876f
C258 source.n36 a_n2524_n3288# 0.014727f
C259 source.n37 a_n2524_n3288# 0.013909f
C260 source.n38 a_n2524_n3288# 0.025884f
C261 source.n39 a_n2524_n3288# 0.025884f
C262 source.n40 a_n2524_n3288# 0.013909f
C263 source.n41 a_n2524_n3288# 0.014727f
C264 source.n42 a_n2524_n3288# 0.032876f
C265 source.n43 a_n2524_n3288# 0.032876f
C266 source.n44 a_n2524_n3288# 0.032876f
C267 source.n45 a_n2524_n3288# 0.014318f
C268 source.n46 a_n2524_n3288# 0.013909f
C269 source.n47 a_n2524_n3288# 0.025884f
C270 source.n48 a_n2524_n3288# 0.025884f
C271 source.n49 a_n2524_n3288# 0.013909f
C272 source.n50 a_n2524_n3288# 0.014727f
C273 source.n51 a_n2524_n3288# 0.032876f
C274 source.n52 a_n2524_n3288# 0.032876f
C275 source.n53 a_n2524_n3288# 0.014727f
C276 source.n54 a_n2524_n3288# 0.013909f
C277 source.n55 a_n2524_n3288# 0.025884f
C278 source.n56 a_n2524_n3288# 0.025884f
C279 source.n57 a_n2524_n3288# 0.013909f
C280 source.n58 a_n2524_n3288# 0.014727f
C281 source.n59 a_n2524_n3288# 0.032876f
C282 source.n60 a_n2524_n3288# 0.067465f
C283 source.n61 a_n2524_n3288# 0.014727f
C284 source.n62 a_n2524_n3288# 0.013909f
C285 source.n63 a_n2524_n3288# 0.055587f
C286 source.n64 a_n2524_n3288# 0.037233f
C287 source.n65 a_n2524_n3288# 1.10062f
C288 source.t27 a_n2524_n3288# 0.245453f
C289 source.t11 a_n2524_n3288# 0.245453f
C290 source.n66 a_n2524_n3288# 2.10157f
C291 source.n67 a_n2524_n3288# 0.427126f
C292 source.t3 a_n2524_n3288# 0.245453f
C293 source.t10 a_n2524_n3288# 0.245453f
C294 source.n68 a_n2524_n3288# 2.10157f
C295 source.n69 a_n2524_n3288# 0.427126f
C296 source.t9 a_n2524_n3288# 0.245453f
C297 source.t2 a_n2524_n3288# 0.245453f
C298 source.n70 a_n2524_n3288# 2.10157f
C299 source.n71 a_n2524_n3288# 0.425688f
C300 source.n72 a_n2524_n3288# 0.034287f
C301 source.n73 a_n2524_n3288# 0.025884f
C302 source.n74 a_n2524_n3288# 0.013909f
C303 source.n75 a_n2524_n3288# 0.032876f
C304 source.n76 a_n2524_n3288# 0.014727f
C305 source.n77 a_n2524_n3288# 0.025884f
C306 source.n78 a_n2524_n3288# 0.013909f
C307 source.n79 a_n2524_n3288# 0.032876f
C308 source.n80 a_n2524_n3288# 0.014727f
C309 source.n81 a_n2524_n3288# 0.025884f
C310 source.n82 a_n2524_n3288# 0.014318f
C311 source.n83 a_n2524_n3288# 0.032876f
C312 source.n84 a_n2524_n3288# 0.013909f
C313 source.n85 a_n2524_n3288# 0.014727f
C314 source.n86 a_n2524_n3288# 0.025884f
C315 source.n87 a_n2524_n3288# 0.013909f
C316 source.n88 a_n2524_n3288# 0.032876f
C317 source.n89 a_n2524_n3288# 0.014727f
C318 source.n90 a_n2524_n3288# 0.025884f
C319 source.n91 a_n2524_n3288# 0.013909f
C320 source.n92 a_n2524_n3288# 0.024657f
C321 source.n93 a_n2524_n3288# 0.023241f
C322 source.t20 a_n2524_n3288# 0.055525f
C323 source.n94 a_n2524_n3288# 0.186621f
C324 source.n95 a_n2524_n3288# 1.30581f
C325 source.n96 a_n2524_n3288# 0.013909f
C326 source.n97 a_n2524_n3288# 0.014727f
C327 source.n98 a_n2524_n3288# 0.032876f
C328 source.n99 a_n2524_n3288# 0.032876f
C329 source.n100 a_n2524_n3288# 0.014727f
C330 source.n101 a_n2524_n3288# 0.013909f
C331 source.n102 a_n2524_n3288# 0.025884f
C332 source.n103 a_n2524_n3288# 0.025884f
C333 source.n104 a_n2524_n3288# 0.013909f
C334 source.n105 a_n2524_n3288# 0.014727f
C335 source.n106 a_n2524_n3288# 0.032876f
C336 source.n107 a_n2524_n3288# 0.032876f
C337 source.n108 a_n2524_n3288# 0.014727f
C338 source.n109 a_n2524_n3288# 0.013909f
C339 source.n110 a_n2524_n3288# 0.025884f
C340 source.n111 a_n2524_n3288# 0.025884f
C341 source.n112 a_n2524_n3288# 0.013909f
C342 source.n113 a_n2524_n3288# 0.014727f
C343 source.n114 a_n2524_n3288# 0.032876f
C344 source.n115 a_n2524_n3288# 0.032876f
C345 source.n116 a_n2524_n3288# 0.032876f
C346 source.n117 a_n2524_n3288# 0.014318f
C347 source.n118 a_n2524_n3288# 0.013909f
C348 source.n119 a_n2524_n3288# 0.025884f
C349 source.n120 a_n2524_n3288# 0.025884f
C350 source.n121 a_n2524_n3288# 0.013909f
C351 source.n122 a_n2524_n3288# 0.014727f
C352 source.n123 a_n2524_n3288# 0.032876f
C353 source.n124 a_n2524_n3288# 0.032876f
C354 source.n125 a_n2524_n3288# 0.014727f
C355 source.n126 a_n2524_n3288# 0.013909f
C356 source.n127 a_n2524_n3288# 0.025884f
C357 source.n128 a_n2524_n3288# 0.025884f
C358 source.n129 a_n2524_n3288# 0.013909f
C359 source.n130 a_n2524_n3288# 0.014727f
C360 source.n131 a_n2524_n3288# 0.032876f
C361 source.n132 a_n2524_n3288# 0.067465f
C362 source.n133 a_n2524_n3288# 0.014727f
C363 source.n134 a_n2524_n3288# 0.013909f
C364 source.n135 a_n2524_n3288# 0.055587f
C365 source.n136 a_n2524_n3288# 0.037233f
C366 source.n137 a_n2524_n3288# 0.180773f
C367 source.t23 a_n2524_n3288# 0.245453f
C368 source.t22 a_n2524_n3288# 0.245453f
C369 source.n138 a_n2524_n3288# 2.10157f
C370 source.n139 a_n2524_n3288# 0.427126f
C371 source.t17 a_n2524_n3288# 0.245453f
C372 source.t18 a_n2524_n3288# 0.245453f
C373 source.n140 a_n2524_n3288# 2.10157f
C374 source.n141 a_n2524_n3288# 0.427126f
C375 source.t21 a_n2524_n3288# 0.245453f
C376 source.t19 a_n2524_n3288# 0.245453f
C377 source.n142 a_n2524_n3288# 2.10157f
C378 source.n143 a_n2524_n3288# 1.84677f
C379 source.t5 a_n2524_n3288# 0.245453f
C380 source.t1 a_n2524_n3288# 0.245453f
C381 source.n144 a_n2524_n3288# 2.10156f
C382 source.n145 a_n2524_n3288# 1.84679f
C383 source.t12 a_n2524_n3288# 0.245453f
C384 source.t0 a_n2524_n3288# 0.245453f
C385 source.n146 a_n2524_n3288# 2.10156f
C386 source.n147 a_n2524_n3288# 0.427139f
C387 source.t4 a_n2524_n3288# 0.245453f
C388 source.t7 a_n2524_n3288# 0.245453f
C389 source.n148 a_n2524_n3288# 2.10156f
C390 source.n149 a_n2524_n3288# 0.427139f
C391 source.n150 a_n2524_n3288# 0.034287f
C392 source.n151 a_n2524_n3288# 0.025884f
C393 source.n152 a_n2524_n3288# 0.013909f
C394 source.n153 a_n2524_n3288# 0.032876f
C395 source.n154 a_n2524_n3288# 0.014727f
C396 source.n155 a_n2524_n3288# 0.025884f
C397 source.n156 a_n2524_n3288# 0.013909f
C398 source.n157 a_n2524_n3288# 0.032876f
C399 source.n158 a_n2524_n3288# 0.014727f
C400 source.n159 a_n2524_n3288# 0.025884f
C401 source.n160 a_n2524_n3288# 0.014318f
C402 source.n161 a_n2524_n3288# 0.032876f
C403 source.n162 a_n2524_n3288# 0.014727f
C404 source.n163 a_n2524_n3288# 0.025884f
C405 source.n164 a_n2524_n3288# 0.013909f
C406 source.n165 a_n2524_n3288# 0.032876f
C407 source.n166 a_n2524_n3288# 0.014727f
C408 source.n167 a_n2524_n3288# 0.025884f
C409 source.n168 a_n2524_n3288# 0.013909f
C410 source.n169 a_n2524_n3288# 0.024657f
C411 source.n170 a_n2524_n3288# 0.023241f
C412 source.t6 a_n2524_n3288# 0.055525f
C413 source.n171 a_n2524_n3288# 0.186621f
C414 source.n172 a_n2524_n3288# 1.30581f
C415 source.n173 a_n2524_n3288# 0.013909f
C416 source.n174 a_n2524_n3288# 0.014727f
C417 source.n175 a_n2524_n3288# 0.032876f
C418 source.n176 a_n2524_n3288# 0.032876f
C419 source.n177 a_n2524_n3288# 0.014727f
C420 source.n178 a_n2524_n3288# 0.013909f
C421 source.n179 a_n2524_n3288# 0.025884f
C422 source.n180 a_n2524_n3288# 0.025884f
C423 source.n181 a_n2524_n3288# 0.013909f
C424 source.n182 a_n2524_n3288# 0.014727f
C425 source.n183 a_n2524_n3288# 0.032876f
C426 source.n184 a_n2524_n3288# 0.032876f
C427 source.n185 a_n2524_n3288# 0.014727f
C428 source.n186 a_n2524_n3288# 0.013909f
C429 source.n187 a_n2524_n3288# 0.025884f
C430 source.n188 a_n2524_n3288# 0.025884f
C431 source.n189 a_n2524_n3288# 0.013909f
C432 source.n190 a_n2524_n3288# 0.013909f
C433 source.n191 a_n2524_n3288# 0.014727f
C434 source.n192 a_n2524_n3288# 0.032876f
C435 source.n193 a_n2524_n3288# 0.032876f
C436 source.n194 a_n2524_n3288# 0.032876f
C437 source.n195 a_n2524_n3288# 0.014318f
C438 source.n196 a_n2524_n3288# 0.013909f
C439 source.n197 a_n2524_n3288# 0.025884f
C440 source.n198 a_n2524_n3288# 0.025884f
C441 source.n199 a_n2524_n3288# 0.013909f
C442 source.n200 a_n2524_n3288# 0.014727f
C443 source.n201 a_n2524_n3288# 0.032876f
C444 source.n202 a_n2524_n3288# 0.032876f
C445 source.n203 a_n2524_n3288# 0.014727f
C446 source.n204 a_n2524_n3288# 0.013909f
C447 source.n205 a_n2524_n3288# 0.025884f
C448 source.n206 a_n2524_n3288# 0.025884f
C449 source.n207 a_n2524_n3288# 0.013909f
C450 source.n208 a_n2524_n3288# 0.014727f
C451 source.n209 a_n2524_n3288# 0.032876f
C452 source.n210 a_n2524_n3288# 0.067465f
C453 source.n211 a_n2524_n3288# 0.014727f
C454 source.n212 a_n2524_n3288# 0.013909f
C455 source.n213 a_n2524_n3288# 0.055587f
C456 source.n214 a_n2524_n3288# 0.037233f
C457 source.n215 a_n2524_n3288# 0.180773f
C458 source.t13 a_n2524_n3288# 0.245453f
C459 source.t24 a_n2524_n3288# 0.245453f
C460 source.n216 a_n2524_n3288# 2.10156f
C461 source.n217 a_n2524_n3288# 0.425701f
C462 source.t15 a_n2524_n3288# 0.245453f
C463 source.t25 a_n2524_n3288# 0.245453f
C464 source.n218 a_n2524_n3288# 2.10156f
C465 source.n219 a_n2524_n3288# 0.427139f
C466 source.t14 a_n2524_n3288# 0.245453f
C467 source.t26 a_n2524_n3288# 0.245453f
C468 source.n220 a_n2524_n3288# 2.10156f
C469 source.n221 a_n2524_n3288# 0.427139f
C470 source.n222 a_n2524_n3288# 0.034287f
C471 source.n223 a_n2524_n3288# 0.025884f
C472 source.n224 a_n2524_n3288# 0.013909f
C473 source.n225 a_n2524_n3288# 0.032876f
C474 source.n226 a_n2524_n3288# 0.014727f
C475 source.n227 a_n2524_n3288# 0.025884f
C476 source.n228 a_n2524_n3288# 0.013909f
C477 source.n229 a_n2524_n3288# 0.032876f
C478 source.n230 a_n2524_n3288# 0.014727f
C479 source.n231 a_n2524_n3288# 0.025884f
C480 source.n232 a_n2524_n3288# 0.014318f
C481 source.n233 a_n2524_n3288# 0.032876f
C482 source.n234 a_n2524_n3288# 0.014727f
C483 source.n235 a_n2524_n3288# 0.025884f
C484 source.n236 a_n2524_n3288# 0.013909f
C485 source.n237 a_n2524_n3288# 0.032876f
C486 source.n238 a_n2524_n3288# 0.014727f
C487 source.n239 a_n2524_n3288# 0.025884f
C488 source.n240 a_n2524_n3288# 0.013909f
C489 source.n241 a_n2524_n3288# 0.024657f
C490 source.n242 a_n2524_n3288# 0.023241f
C491 source.t16 a_n2524_n3288# 0.055525f
C492 source.n243 a_n2524_n3288# 0.186621f
C493 source.n244 a_n2524_n3288# 1.30581f
C494 source.n245 a_n2524_n3288# 0.013909f
C495 source.n246 a_n2524_n3288# 0.014727f
C496 source.n247 a_n2524_n3288# 0.032876f
C497 source.n248 a_n2524_n3288# 0.032876f
C498 source.n249 a_n2524_n3288# 0.014727f
C499 source.n250 a_n2524_n3288# 0.013909f
C500 source.n251 a_n2524_n3288# 0.025884f
C501 source.n252 a_n2524_n3288# 0.025884f
C502 source.n253 a_n2524_n3288# 0.013909f
C503 source.n254 a_n2524_n3288# 0.014727f
C504 source.n255 a_n2524_n3288# 0.032876f
C505 source.n256 a_n2524_n3288# 0.032876f
C506 source.n257 a_n2524_n3288# 0.014727f
C507 source.n258 a_n2524_n3288# 0.013909f
C508 source.n259 a_n2524_n3288# 0.025884f
C509 source.n260 a_n2524_n3288# 0.025884f
C510 source.n261 a_n2524_n3288# 0.013909f
C511 source.n262 a_n2524_n3288# 0.013909f
C512 source.n263 a_n2524_n3288# 0.014727f
C513 source.n264 a_n2524_n3288# 0.032876f
C514 source.n265 a_n2524_n3288# 0.032876f
C515 source.n266 a_n2524_n3288# 0.032876f
C516 source.n267 a_n2524_n3288# 0.014318f
C517 source.n268 a_n2524_n3288# 0.013909f
C518 source.n269 a_n2524_n3288# 0.025884f
C519 source.n270 a_n2524_n3288# 0.025884f
C520 source.n271 a_n2524_n3288# 0.013909f
C521 source.n272 a_n2524_n3288# 0.014727f
C522 source.n273 a_n2524_n3288# 0.032876f
C523 source.n274 a_n2524_n3288# 0.032876f
C524 source.n275 a_n2524_n3288# 0.014727f
C525 source.n276 a_n2524_n3288# 0.013909f
C526 source.n277 a_n2524_n3288# 0.025884f
C527 source.n278 a_n2524_n3288# 0.025884f
C528 source.n279 a_n2524_n3288# 0.013909f
C529 source.n280 a_n2524_n3288# 0.014727f
C530 source.n281 a_n2524_n3288# 0.032876f
C531 source.n282 a_n2524_n3288# 0.067465f
C532 source.n283 a_n2524_n3288# 0.014727f
C533 source.n284 a_n2524_n3288# 0.013909f
C534 source.n285 a_n2524_n3288# 0.055587f
C535 source.n286 a_n2524_n3288# 0.037233f
C536 source.n287 a_n2524_n3288# 0.314596f
C537 source.n288 a_n2524_n3288# 1.64441f
C538 drain_right.n0 a_n2524_n3288# 0.032234f
C539 drain_right.n1 a_n2524_n3288# 0.024334f
C540 drain_right.n2 a_n2524_n3288# 0.013076f
C541 drain_right.n3 a_n2524_n3288# 0.030907f
C542 drain_right.n4 a_n2524_n3288# 0.013845f
C543 drain_right.n5 a_n2524_n3288# 0.024334f
C544 drain_right.n6 a_n2524_n3288# 0.013076f
C545 drain_right.n7 a_n2524_n3288# 0.030907f
C546 drain_right.n8 a_n2524_n3288# 0.013845f
C547 drain_right.n9 a_n2524_n3288# 0.024334f
C548 drain_right.n10 a_n2524_n3288# 0.013461f
C549 drain_right.n11 a_n2524_n3288# 0.030907f
C550 drain_right.n12 a_n2524_n3288# 0.013845f
C551 drain_right.n13 a_n2524_n3288# 0.024334f
C552 drain_right.n14 a_n2524_n3288# 0.013076f
C553 drain_right.n15 a_n2524_n3288# 0.030907f
C554 drain_right.n16 a_n2524_n3288# 0.013845f
C555 drain_right.n17 a_n2524_n3288# 0.024334f
C556 drain_right.n18 a_n2524_n3288# 0.013076f
C557 drain_right.n19 a_n2524_n3288# 0.023181f
C558 drain_right.n20 a_n2524_n3288# 0.021849f
C559 drain_right.t11 a_n2524_n3288# 0.052201f
C560 drain_right.n21 a_n2524_n3288# 0.175448f
C561 drain_right.n22 a_n2524_n3288# 1.22763f
C562 drain_right.n23 a_n2524_n3288# 0.013076f
C563 drain_right.n24 a_n2524_n3288# 0.013845f
C564 drain_right.n25 a_n2524_n3288# 0.030907f
C565 drain_right.n26 a_n2524_n3288# 0.030907f
C566 drain_right.n27 a_n2524_n3288# 0.013845f
C567 drain_right.n28 a_n2524_n3288# 0.013076f
C568 drain_right.n29 a_n2524_n3288# 0.024334f
C569 drain_right.n30 a_n2524_n3288# 0.024334f
C570 drain_right.n31 a_n2524_n3288# 0.013076f
C571 drain_right.n32 a_n2524_n3288# 0.013845f
C572 drain_right.n33 a_n2524_n3288# 0.030907f
C573 drain_right.n34 a_n2524_n3288# 0.030907f
C574 drain_right.n35 a_n2524_n3288# 0.013845f
C575 drain_right.n36 a_n2524_n3288# 0.013076f
C576 drain_right.n37 a_n2524_n3288# 0.024334f
C577 drain_right.n38 a_n2524_n3288# 0.024334f
C578 drain_right.n39 a_n2524_n3288# 0.013076f
C579 drain_right.n40 a_n2524_n3288# 0.013076f
C580 drain_right.n41 a_n2524_n3288# 0.013845f
C581 drain_right.n42 a_n2524_n3288# 0.030907f
C582 drain_right.n43 a_n2524_n3288# 0.030907f
C583 drain_right.n44 a_n2524_n3288# 0.030907f
C584 drain_right.n45 a_n2524_n3288# 0.013461f
C585 drain_right.n46 a_n2524_n3288# 0.013076f
C586 drain_right.n47 a_n2524_n3288# 0.024334f
C587 drain_right.n48 a_n2524_n3288# 0.024334f
C588 drain_right.n49 a_n2524_n3288# 0.013076f
C589 drain_right.n50 a_n2524_n3288# 0.013845f
C590 drain_right.n51 a_n2524_n3288# 0.030907f
C591 drain_right.n52 a_n2524_n3288# 0.030907f
C592 drain_right.n53 a_n2524_n3288# 0.013845f
C593 drain_right.n54 a_n2524_n3288# 0.013076f
C594 drain_right.n55 a_n2524_n3288# 0.024334f
C595 drain_right.n56 a_n2524_n3288# 0.024334f
C596 drain_right.n57 a_n2524_n3288# 0.013076f
C597 drain_right.n58 a_n2524_n3288# 0.013845f
C598 drain_right.n59 a_n2524_n3288# 0.030907f
C599 drain_right.n60 a_n2524_n3288# 0.063425f
C600 drain_right.n61 a_n2524_n3288# 0.013845f
C601 drain_right.n62 a_n2524_n3288# 0.013076f
C602 drain_right.n63 a_n2524_n3288# 0.052258f
C603 drain_right.n64 a_n2524_n3288# 0.054321f
C604 drain_right.t0 a_n2524_n3288# 0.230757f
C605 drain_right.t13 a_n2524_n3288# 0.230757f
C606 drain_right.n65 a_n2524_n3288# 2.05338f
C607 drain_right.n66 a_n2524_n3288# 0.452871f
C608 drain_right.t8 a_n2524_n3288# 0.230757f
C609 drain_right.t4 a_n2524_n3288# 0.230757f
C610 drain_right.n67 a_n2524_n3288# 2.05928f
C611 drain_right.t9 a_n2524_n3288# 0.230757f
C612 drain_right.t12 a_n2524_n3288# 0.230757f
C613 drain_right.n68 a_n2524_n3288# 2.05338f
C614 drain_right.n69 a_n2524_n3288# 0.659255f
C615 drain_right.n70 a_n2524_n3288# 1.34003f
C616 drain_right.t7 a_n2524_n3288# 0.230757f
C617 drain_right.t2 a_n2524_n3288# 0.230757f
C618 drain_right.n71 a_n2524_n3288# 2.05928f
C619 drain_right.t10 a_n2524_n3288# 0.230757f
C620 drain_right.t6 a_n2524_n3288# 0.230757f
C621 drain_right.n72 a_n2524_n3288# 2.05339f
C622 drain_right.n73 a_n2524_n3288# 0.717876f
C623 drain_right.t1 a_n2524_n3288# 0.230757f
C624 drain_right.t5 a_n2524_n3288# 0.230757f
C625 drain_right.n74 a_n2524_n3288# 2.05339f
C626 drain_right.n75 a_n2524_n3288# 0.356985f
C627 drain_right.n76 a_n2524_n3288# 0.032234f
C628 drain_right.n77 a_n2524_n3288# 0.024334f
C629 drain_right.n78 a_n2524_n3288# 0.013076f
C630 drain_right.n79 a_n2524_n3288# 0.030907f
C631 drain_right.n80 a_n2524_n3288# 0.013845f
C632 drain_right.n81 a_n2524_n3288# 0.024334f
C633 drain_right.n82 a_n2524_n3288# 0.013076f
C634 drain_right.n83 a_n2524_n3288# 0.030907f
C635 drain_right.n84 a_n2524_n3288# 0.013845f
C636 drain_right.n85 a_n2524_n3288# 0.024334f
C637 drain_right.n86 a_n2524_n3288# 0.013461f
C638 drain_right.n87 a_n2524_n3288# 0.030907f
C639 drain_right.n88 a_n2524_n3288# 0.013076f
C640 drain_right.n89 a_n2524_n3288# 0.013845f
C641 drain_right.n90 a_n2524_n3288# 0.024334f
C642 drain_right.n91 a_n2524_n3288# 0.013076f
C643 drain_right.n92 a_n2524_n3288# 0.030907f
C644 drain_right.n93 a_n2524_n3288# 0.013845f
C645 drain_right.n94 a_n2524_n3288# 0.024334f
C646 drain_right.n95 a_n2524_n3288# 0.013076f
C647 drain_right.n96 a_n2524_n3288# 0.023181f
C648 drain_right.n97 a_n2524_n3288# 0.021849f
C649 drain_right.t3 a_n2524_n3288# 0.052201f
C650 drain_right.n98 a_n2524_n3288# 0.175448f
C651 drain_right.n99 a_n2524_n3288# 1.22763f
C652 drain_right.n100 a_n2524_n3288# 0.013076f
C653 drain_right.n101 a_n2524_n3288# 0.013845f
C654 drain_right.n102 a_n2524_n3288# 0.030907f
C655 drain_right.n103 a_n2524_n3288# 0.030907f
C656 drain_right.n104 a_n2524_n3288# 0.013845f
C657 drain_right.n105 a_n2524_n3288# 0.013076f
C658 drain_right.n106 a_n2524_n3288# 0.024334f
C659 drain_right.n107 a_n2524_n3288# 0.024334f
C660 drain_right.n108 a_n2524_n3288# 0.013076f
C661 drain_right.n109 a_n2524_n3288# 0.013845f
C662 drain_right.n110 a_n2524_n3288# 0.030907f
C663 drain_right.n111 a_n2524_n3288# 0.030907f
C664 drain_right.n112 a_n2524_n3288# 0.013845f
C665 drain_right.n113 a_n2524_n3288# 0.013076f
C666 drain_right.n114 a_n2524_n3288# 0.024334f
C667 drain_right.n115 a_n2524_n3288# 0.024334f
C668 drain_right.n116 a_n2524_n3288# 0.013076f
C669 drain_right.n117 a_n2524_n3288# 0.013845f
C670 drain_right.n118 a_n2524_n3288# 0.030907f
C671 drain_right.n119 a_n2524_n3288# 0.030907f
C672 drain_right.n120 a_n2524_n3288# 0.030907f
C673 drain_right.n121 a_n2524_n3288# 0.013461f
C674 drain_right.n122 a_n2524_n3288# 0.013076f
C675 drain_right.n123 a_n2524_n3288# 0.024334f
C676 drain_right.n124 a_n2524_n3288# 0.024334f
C677 drain_right.n125 a_n2524_n3288# 0.013076f
C678 drain_right.n126 a_n2524_n3288# 0.013845f
C679 drain_right.n127 a_n2524_n3288# 0.030907f
C680 drain_right.n128 a_n2524_n3288# 0.030907f
C681 drain_right.n129 a_n2524_n3288# 0.013845f
C682 drain_right.n130 a_n2524_n3288# 0.013076f
C683 drain_right.n131 a_n2524_n3288# 0.024334f
C684 drain_right.n132 a_n2524_n3288# 0.024334f
C685 drain_right.n133 a_n2524_n3288# 0.013076f
C686 drain_right.n134 a_n2524_n3288# 0.013845f
C687 drain_right.n135 a_n2524_n3288# 0.030907f
C688 drain_right.n136 a_n2524_n3288# 0.063425f
C689 drain_right.n137 a_n2524_n3288# 0.013845f
C690 drain_right.n138 a_n2524_n3288# 0.013076f
C691 drain_right.n139 a_n2524_n3288# 0.052258f
C692 drain_right.n140 a_n2524_n3288# 0.051841f
C693 drain_right.n141 a_n2524_n3288# 0.349702f
C694 minus.n0 a_n2524_n3288# 0.039088f
C695 minus.n1 a_n2524_n3288# 0.00887f
C696 minus.t7 a_n2524_n3288# 1.07002f
C697 minus.n2 a_n2524_n3288# 0.078177f
C698 minus.n3 a_n2524_n3288# 0.00887f
C699 minus.t3 a_n2524_n3288# 1.07002f
C700 minus.t6 a_n2524_n3288# 1.09339f
C701 minus.t4 a_n2524_n3288# 1.07002f
C702 minus.n4 a_n2524_n3288# 0.428014f
C703 minus.n5 a_n2524_n3288# 0.405655f
C704 minus.n6 a_n2524_n3288# 0.182548f
C705 minus.n7 a_n2524_n3288# 0.065107f
C706 minus.n8 a_n2524_n3288# 0.432524f
C707 minus.t8 a_n2524_n3288# 1.07002f
C708 minus.n9 a_n2524_n3288# 0.435175f
C709 minus.t9 a_n2524_n3288# 1.07002f
C710 minus.n10 a_n2524_n3288# 0.432524f
C711 minus.n11 a_n2524_n3288# 0.065107f
C712 minus.n12 a_n2524_n3288# 0.052159f
C713 minus.n13 a_n2524_n3288# 0.039088f
C714 minus.n14 a_n2524_n3288# 0.423172f
C715 minus.n15 a_n2524_n3288# 0.00887f
C716 minus.t5 a_n2524_n3288# 1.07002f
C717 minus.n16 a_n2524_n3288# 0.424136f
C718 minus.n17 a_n2524_n3288# 1.55046f
C719 minus.n18 a_n2524_n3288# 0.039088f
C720 minus.n19 a_n2524_n3288# 0.00887f
C721 minus.n20 a_n2524_n3288# 0.078177f
C722 minus.n21 a_n2524_n3288# 0.00887f
C723 minus.t13 a_n2524_n3288# 1.09339f
C724 minus.t2 a_n2524_n3288# 1.07002f
C725 minus.n22 a_n2524_n3288# 0.428014f
C726 minus.n23 a_n2524_n3288# 0.405655f
C727 minus.n24 a_n2524_n3288# 0.182548f
C728 minus.n25 a_n2524_n3288# 0.065107f
C729 minus.t11 a_n2524_n3288# 1.07002f
C730 minus.n26 a_n2524_n3288# 0.432524f
C731 minus.t1 a_n2524_n3288# 1.07002f
C732 minus.n27 a_n2524_n3288# 0.435175f
C733 minus.t12 a_n2524_n3288# 1.07002f
C734 minus.n28 a_n2524_n3288# 0.432524f
C735 minus.n29 a_n2524_n3288# 0.065107f
C736 minus.n30 a_n2524_n3288# 0.052159f
C737 minus.n31 a_n2524_n3288# 0.039088f
C738 minus.t0 a_n2524_n3288# 1.07002f
C739 minus.n32 a_n2524_n3288# 0.423172f
C740 minus.n33 a_n2524_n3288# 0.00887f
C741 minus.t10 a_n2524_n3288# 1.07002f
C742 minus.n34 a_n2524_n3288# 0.424136f
C743 minus.n35 a_n2524_n3288# 0.276134f
C744 minus.n36 a_n2524_n3288# 1.86249f
.ends

