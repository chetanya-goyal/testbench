* NGSPICE file created from diffpair445.ext - technology: sky130A

.subckt diffpair445 minus drain_right drain_left source plus
X0 a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.5
X1 source.t19 plus.t0 drain_left.t7 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X2 drain_left.t6 plus.t1 source.t18 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X3 drain_right.t11 minus.t0 source.t7 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X4 source.t1 minus.t1 drain_right.t10 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X5 source.t4 minus.t2 drain_right.t9 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X6 a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X7 source.t17 plus.t2 drain_left.t4 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X8 source.t6 minus.t3 drain_right.t8 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X9 drain_right.t7 minus.t4 source.t5 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X10 drain_left.t1 plus.t3 source.t16 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X11 drain_right.t6 minus.t5 source.t22 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X12 drain_left.t0 plus.t4 source.t15 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X13 source.t14 plus.t5 drain_left.t2 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X14 drain_right.t5 minus.t6 source.t0 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X15 source.t23 minus.t7 drain_right.t4 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X16 source.t3 minus.t8 drain_right.t3 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X17 a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X18 a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X19 drain_right.t2 minus.t9 source.t2 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X20 drain_right.t1 minus.t10 source.t20 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X21 drain_left.t3 plus.t6 source.t13 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X22 source.t21 minus.t11 drain_right.t0 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X23 source.t12 plus.t7 drain_left.t8 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X24 drain_left.t5 plus.t8 source.t11 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X25 source.t10 plus.t9 drain_left.t11 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X26 source.t9 plus.t10 drain_left.t10 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X27 drain_left.t9 plus.t11 source.t8 a_n1878_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
R0 plus.n5 plus.t2 683.635
R1 plus.n19 plus.t8 683.635
R2 plus.n12 plus.t11 656.966
R3 plus.n10 plus.t7 656.966
R4 plus.n9 plus.t4 656.966
R5 plus.n3 plus.t10 656.966
R6 plus.n4 plus.t6 656.966
R7 plus.n26 plus.t5 656.966
R8 plus.n24 plus.t1 656.966
R9 plus.n23 plus.t0 656.966
R10 plus.n17 plus.t3 656.966
R11 plus.n18 plus.t9 656.966
R12 plus.n6 plus.n3 161.3
R13 plus.n8 plus.n7 161.3
R14 plus.n9 plus.n2 161.3
R15 plus.n10 plus.n1 161.3
R16 plus.n11 plus.n0 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n20 plus.n17 161.3
R19 plus.n22 plus.n21 161.3
R20 plus.n23 plus.n16 161.3
R21 plus.n24 plus.n15 161.3
R22 plus.n25 plus.n14 161.3
R23 plus.n27 plus.n26 161.3
R24 plus.n10 plus.n9 48.2005
R25 plus.n4 plus.n3 48.2005
R26 plus.n24 plus.n23 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n12 plus.n11 47.4702
R29 plus.n26 plus.n25 47.4702
R30 plus.n6 plus.n5 45.1192
R31 plus.n20 plus.n19 45.1192
R32 plus plus.n27 30.1467
R33 plus.n8 plus.n3 24.1005
R34 plus.n9 plus.n8 24.1005
R35 plus.n23 plus.n22 24.1005
R36 plus.n22 plus.n17 24.1005
R37 plus.n5 plus.n4 13.6377
R38 plus.n19 plus.n18 13.6377
R39 plus plus.n13 12.1747
R40 plus.n11 plus.n10 0.730803
R41 plus.n25 plus.n24 0.730803
R42 plus.n7 plus.n6 0.189894
R43 plus.n7 plus.n2 0.189894
R44 plus.n2 plus.n1 0.189894
R45 plus.n1 plus.n0 0.189894
R46 plus.n13 plus.n0 0.189894
R47 plus.n27 plus.n14 0.189894
R48 plus.n15 plus.n14 0.189894
R49 plus.n16 plus.n15 0.189894
R50 plus.n21 plus.n16 0.189894
R51 plus.n21 plus.n20 0.189894
R52 drain_left.n6 drain_left.n4 60.2682
R53 drain_left.n3 drain_left.n2 60.2127
R54 drain_left.n3 drain_left.n0 60.2127
R55 drain_left.n6 drain_left.n5 59.5527
R56 drain_left.n3 drain_left.n1 59.5525
R57 drain_left.n8 drain_left.n7 59.5525
R58 drain_left drain_left.n3 30.9447
R59 drain_left drain_left.n8 6.36873
R60 drain_left.n1 drain_left.t7 1.6505
R61 drain_left.n1 drain_left.t1 1.6505
R62 drain_left.n2 drain_left.t11 1.6505
R63 drain_left.n2 drain_left.t5 1.6505
R64 drain_left.n0 drain_left.t2 1.6505
R65 drain_left.n0 drain_left.t6 1.6505
R66 drain_left.n7 drain_left.t8 1.6505
R67 drain_left.n7 drain_left.t9 1.6505
R68 drain_left.n5 drain_left.t10 1.6505
R69 drain_left.n5 drain_left.t0 1.6505
R70 drain_left.n4 drain_left.t4 1.6505
R71 drain_left.n4 drain_left.t3 1.6505
R72 drain_left.n8 drain_left.n6 0.716017
R73 source.n538 source.n478 289.615
R74 source.n468 source.n408 289.615
R75 source.n402 source.n342 289.615
R76 source.n332 source.n272 289.615
R77 source.n60 source.n0 289.615
R78 source.n130 source.n70 289.615
R79 source.n196 source.n136 289.615
R80 source.n266 source.n206 289.615
R81 source.n498 source.n497 185
R82 source.n503 source.n502 185
R83 source.n505 source.n504 185
R84 source.n494 source.n493 185
R85 source.n511 source.n510 185
R86 source.n513 source.n512 185
R87 source.n490 source.n489 185
R88 source.n520 source.n519 185
R89 source.n521 source.n488 185
R90 source.n523 source.n522 185
R91 source.n486 source.n485 185
R92 source.n529 source.n528 185
R93 source.n531 source.n530 185
R94 source.n482 source.n481 185
R95 source.n537 source.n536 185
R96 source.n539 source.n538 185
R97 source.n428 source.n427 185
R98 source.n433 source.n432 185
R99 source.n435 source.n434 185
R100 source.n424 source.n423 185
R101 source.n441 source.n440 185
R102 source.n443 source.n442 185
R103 source.n420 source.n419 185
R104 source.n450 source.n449 185
R105 source.n451 source.n418 185
R106 source.n453 source.n452 185
R107 source.n416 source.n415 185
R108 source.n459 source.n458 185
R109 source.n461 source.n460 185
R110 source.n412 source.n411 185
R111 source.n467 source.n466 185
R112 source.n469 source.n468 185
R113 source.n362 source.n361 185
R114 source.n367 source.n366 185
R115 source.n369 source.n368 185
R116 source.n358 source.n357 185
R117 source.n375 source.n374 185
R118 source.n377 source.n376 185
R119 source.n354 source.n353 185
R120 source.n384 source.n383 185
R121 source.n385 source.n352 185
R122 source.n387 source.n386 185
R123 source.n350 source.n349 185
R124 source.n393 source.n392 185
R125 source.n395 source.n394 185
R126 source.n346 source.n345 185
R127 source.n401 source.n400 185
R128 source.n403 source.n402 185
R129 source.n292 source.n291 185
R130 source.n297 source.n296 185
R131 source.n299 source.n298 185
R132 source.n288 source.n287 185
R133 source.n305 source.n304 185
R134 source.n307 source.n306 185
R135 source.n284 source.n283 185
R136 source.n314 source.n313 185
R137 source.n315 source.n282 185
R138 source.n317 source.n316 185
R139 source.n280 source.n279 185
R140 source.n323 source.n322 185
R141 source.n325 source.n324 185
R142 source.n276 source.n275 185
R143 source.n331 source.n330 185
R144 source.n333 source.n332 185
R145 source.n61 source.n60 185
R146 source.n59 source.n58 185
R147 source.n4 source.n3 185
R148 source.n53 source.n52 185
R149 source.n51 source.n50 185
R150 source.n8 source.n7 185
R151 source.n45 source.n44 185
R152 source.n43 source.n10 185
R153 source.n42 source.n41 185
R154 source.n13 source.n11 185
R155 source.n36 source.n35 185
R156 source.n34 source.n33 185
R157 source.n17 source.n16 185
R158 source.n28 source.n27 185
R159 source.n26 source.n25 185
R160 source.n21 source.n20 185
R161 source.n131 source.n130 185
R162 source.n129 source.n128 185
R163 source.n74 source.n73 185
R164 source.n123 source.n122 185
R165 source.n121 source.n120 185
R166 source.n78 source.n77 185
R167 source.n115 source.n114 185
R168 source.n113 source.n80 185
R169 source.n112 source.n111 185
R170 source.n83 source.n81 185
R171 source.n106 source.n105 185
R172 source.n104 source.n103 185
R173 source.n87 source.n86 185
R174 source.n98 source.n97 185
R175 source.n96 source.n95 185
R176 source.n91 source.n90 185
R177 source.n197 source.n196 185
R178 source.n195 source.n194 185
R179 source.n140 source.n139 185
R180 source.n189 source.n188 185
R181 source.n187 source.n186 185
R182 source.n144 source.n143 185
R183 source.n181 source.n180 185
R184 source.n179 source.n146 185
R185 source.n178 source.n177 185
R186 source.n149 source.n147 185
R187 source.n172 source.n171 185
R188 source.n170 source.n169 185
R189 source.n153 source.n152 185
R190 source.n164 source.n163 185
R191 source.n162 source.n161 185
R192 source.n157 source.n156 185
R193 source.n267 source.n266 185
R194 source.n265 source.n264 185
R195 source.n210 source.n209 185
R196 source.n259 source.n258 185
R197 source.n257 source.n256 185
R198 source.n214 source.n213 185
R199 source.n251 source.n250 185
R200 source.n249 source.n216 185
R201 source.n248 source.n247 185
R202 source.n219 source.n217 185
R203 source.n242 source.n241 185
R204 source.n240 source.n239 185
R205 source.n223 source.n222 185
R206 source.n234 source.n233 185
R207 source.n232 source.n231 185
R208 source.n227 source.n226 185
R209 source.n499 source.t2 149.524
R210 source.n429 source.t1 149.524
R211 source.n363 source.t11 149.524
R212 source.n293 source.t14 149.524
R213 source.n22 source.t8 149.524
R214 source.n92 source.t17 149.524
R215 source.n158 source.t20 149.524
R216 source.n228 source.t3 149.524
R217 source.n503 source.n497 104.615
R218 source.n504 source.n503 104.615
R219 source.n504 source.n493 104.615
R220 source.n511 source.n493 104.615
R221 source.n512 source.n511 104.615
R222 source.n512 source.n489 104.615
R223 source.n520 source.n489 104.615
R224 source.n521 source.n520 104.615
R225 source.n522 source.n521 104.615
R226 source.n522 source.n485 104.615
R227 source.n529 source.n485 104.615
R228 source.n530 source.n529 104.615
R229 source.n530 source.n481 104.615
R230 source.n537 source.n481 104.615
R231 source.n538 source.n537 104.615
R232 source.n433 source.n427 104.615
R233 source.n434 source.n433 104.615
R234 source.n434 source.n423 104.615
R235 source.n441 source.n423 104.615
R236 source.n442 source.n441 104.615
R237 source.n442 source.n419 104.615
R238 source.n450 source.n419 104.615
R239 source.n451 source.n450 104.615
R240 source.n452 source.n451 104.615
R241 source.n452 source.n415 104.615
R242 source.n459 source.n415 104.615
R243 source.n460 source.n459 104.615
R244 source.n460 source.n411 104.615
R245 source.n467 source.n411 104.615
R246 source.n468 source.n467 104.615
R247 source.n367 source.n361 104.615
R248 source.n368 source.n367 104.615
R249 source.n368 source.n357 104.615
R250 source.n375 source.n357 104.615
R251 source.n376 source.n375 104.615
R252 source.n376 source.n353 104.615
R253 source.n384 source.n353 104.615
R254 source.n385 source.n384 104.615
R255 source.n386 source.n385 104.615
R256 source.n386 source.n349 104.615
R257 source.n393 source.n349 104.615
R258 source.n394 source.n393 104.615
R259 source.n394 source.n345 104.615
R260 source.n401 source.n345 104.615
R261 source.n402 source.n401 104.615
R262 source.n297 source.n291 104.615
R263 source.n298 source.n297 104.615
R264 source.n298 source.n287 104.615
R265 source.n305 source.n287 104.615
R266 source.n306 source.n305 104.615
R267 source.n306 source.n283 104.615
R268 source.n314 source.n283 104.615
R269 source.n315 source.n314 104.615
R270 source.n316 source.n315 104.615
R271 source.n316 source.n279 104.615
R272 source.n323 source.n279 104.615
R273 source.n324 source.n323 104.615
R274 source.n324 source.n275 104.615
R275 source.n331 source.n275 104.615
R276 source.n332 source.n331 104.615
R277 source.n60 source.n59 104.615
R278 source.n59 source.n3 104.615
R279 source.n52 source.n3 104.615
R280 source.n52 source.n51 104.615
R281 source.n51 source.n7 104.615
R282 source.n44 source.n7 104.615
R283 source.n44 source.n43 104.615
R284 source.n43 source.n42 104.615
R285 source.n42 source.n11 104.615
R286 source.n35 source.n11 104.615
R287 source.n35 source.n34 104.615
R288 source.n34 source.n16 104.615
R289 source.n27 source.n16 104.615
R290 source.n27 source.n26 104.615
R291 source.n26 source.n20 104.615
R292 source.n130 source.n129 104.615
R293 source.n129 source.n73 104.615
R294 source.n122 source.n73 104.615
R295 source.n122 source.n121 104.615
R296 source.n121 source.n77 104.615
R297 source.n114 source.n77 104.615
R298 source.n114 source.n113 104.615
R299 source.n113 source.n112 104.615
R300 source.n112 source.n81 104.615
R301 source.n105 source.n81 104.615
R302 source.n105 source.n104 104.615
R303 source.n104 source.n86 104.615
R304 source.n97 source.n86 104.615
R305 source.n97 source.n96 104.615
R306 source.n96 source.n90 104.615
R307 source.n196 source.n195 104.615
R308 source.n195 source.n139 104.615
R309 source.n188 source.n139 104.615
R310 source.n188 source.n187 104.615
R311 source.n187 source.n143 104.615
R312 source.n180 source.n143 104.615
R313 source.n180 source.n179 104.615
R314 source.n179 source.n178 104.615
R315 source.n178 source.n147 104.615
R316 source.n171 source.n147 104.615
R317 source.n171 source.n170 104.615
R318 source.n170 source.n152 104.615
R319 source.n163 source.n152 104.615
R320 source.n163 source.n162 104.615
R321 source.n162 source.n156 104.615
R322 source.n266 source.n265 104.615
R323 source.n265 source.n209 104.615
R324 source.n258 source.n209 104.615
R325 source.n258 source.n257 104.615
R326 source.n257 source.n213 104.615
R327 source.n250 source.n213 104.615
R328 source.n250 source.n249 104.615
R329 source.n249 source.n248 104.615
R330 source.n248 source.n217 104.615
R331 source.n241 source.n217 104.615
R332 source.n241 source.n240 104.615
R333 source.n240 source.n222 104.615
R334 source.n233 source.n222 104.615
R335 source.n233 source.n232 104.615
R336 source.n232 source.n226 104.615
R337 source.t2 source.n497 52.3082
R338 source.t1 source.n427 52.3082
R339 source.t11 source.n361 52.3082
R340 source.t14 source.n291 52.3082
R341 source.t8 source.n20 52.3082
R342 source.t17 source.n90 52.3082
R343 source.t20 source.n156 52.3082
R344 source.t3 source.n226 52.3082
R345 source.n67 source.n66 42.8739
R346 source.n69 source.n68 42.8739
R347 source.n203 source.n202 42.8739
R348 source.n205 source.n204 42.8739
R349 source.n477 source.n476 42.8737
R350 source.n475 source.n474 42.8737
R351 source.n341 source.n340 42.8737
R352 source.n339 source.n338 42.8737
R353 source.n543 source.n542 29.8581
R354 source.n473 source.n472 29.8581
R355 source.n407 source.n406 29.8581
R356 source.n337 source.n336 29.8581
R357 source.n65 source.n64 29.8581
R358 source.n135 source.n134 29.8581
R359 source.n201 source.n200 29.8581
R360 source.n271 source.n270 29.8581
R361 source.n337 source.n271 22.0032
R362 source.n544 source.n65 16.3826
R363 source.n523 source.n488 13.1884
R364 source.n453 source.n418 13.1884
R365 source.n387 source.n352 13.1884
R366 source.n317 source.n282 13.1884
R367 source.n45 source.n10 13.1884
R368 source.n115 source.n80 13.1884
R369 source.n181 source.n146 13.1884
R370 source.n251 source.n216 13.1884
R371 source.n519 source.n518 12.8005
R372 source.n524 source.n486 12.8005
R373 source.n449 source.n448 12.8005
R374 source.n454 source.n416 12.8005
R375 source.n383 source.n382 12.8005
R376 source.n388 source.n350 12.8005
R377 source.n313 source.n312 12.8005
R378 source.n318 source.n280 12.8005
R379 source.n46 source.n8 12.8005
R380 source.n41 source.n12 12.8005
R381 source.n116 source.n78 12.8005
R382 source.n111 source.n82 12.8005
R383 source.n182 source.n144 12.8005
R384 source.n177 source.n148 12.8005
R385 source.n252 source.n214 12.8005
R386 source.n247 source.n218 12.8005
R387 source.n517 source.n490 12.0247
R388 source.n528 source.n527 12.0247
R389 source.n447 source.n420 12.0247
R390 source.n458 source.n457 12.0247
R391 source.n381 source.n354 12.0247
R392 source.n392 source.n391 12.0247
R393 source.n311 source.n284 12.0247
R394 source.n322 source.n321 12.0247
R395 source.n50 source.n49 12.0247
R396 source.n40 source.n13 12.0247
R397 source.n120 source.n119 12.0247
R398 source.n110 source.n83 12.0247
R399 source.n186 source.n185 12.0247
R400 source.n176 source.n149 12.0247
R401 source.n256 source.n255 12.0247
R402 source.n246 source.n219 12.0247
R403 source.n514 source.n513 11.249
R404 source.n531 source.n484 11.249
R405 source.n444 source.n443 11.249
R406 source.n461 source.n414 11.249
R407 source.n378 source.n377 11.249
R408 source.n395 source.n348 11.249
R409 source.n308 source.n307 11.249
R410 source.n325 source.n278 11.249
R411 source.n53 source.n6 11.249
R412 source.n37 source.n36 11.249
R413 source.n123 source.n76 11.249
R414 source.n107 source.n106 11.249
R415 source.n189 source.n142 11.249
R416 source.n173 source.n172 11.249
R417 source.n259 source.n212 11.249
R418 source.n243 source.n242 11.249
R419 source.n510 source.n492 10.4732
R420 source.n532 source.n482 10.4732
R421 source.n440 source.n422 10.4732
R422 source.n462 source.n412 10.4732
R423 source.n374 source.n356 10.4732
R424 source.n396 source.n346 10.4732
R425 source.n304 source.n286 10.4732
R426 source.n326 source.n276 10.4732
R427 source.n54 source.n4 10.4732
R428 source.n33 source.n15 10.4732
R429 source.n124 source.n74 10.4732
R430 source.n103 source.n85 10.4732
R431 source.n190 source.n140 10.4732
R432 source.n169 source.n151 10.4732
R433 source.n260 source.n210 10.4732
R434 source.n239 source.n221 10.4732
R435 source.n499 source.n498 10.2747
R436 source.n429 source.n428 10.2747
R437 source.n363 source.n362 10.2747
R438 source.n293 source.n292 10.2747
R439 source.n22 source.n21 10.2747
R440 source.n92 source.n91 10.2747
R441 source.n158 source.n157 10.2747
R442 source.n228 source.n227 10.2747
R443 source.n509 source.n494 9.69747
R444 source.n536 source.n535 9.69747
R445 source.n439 source.n424 9.69747
R446 source.n466 source.n465 9.69747
R447 source.n373 source.n358 9.69747
R448 source.n400 source.n399 9.69747
R449 source.n303 source.n288 9.69747
R450 source.n330 source.n329 9.69747
R451 source.n58 source.n57 9.69747
R452 source.n32 source.n17 9.69747
R453 source.n128 source.n127 9.69747
R454 source.n102 source.n87 9.69747
R455 source.n194 source.n193 9.69747
R456 source.n168 source.n153 9.69747
R457 source.n264 source.n263 9.69747
R458 source.n238 source.n223 9.69747
R459 source.n542 source.n541 9.45567
R460 source.n472 source.n471 9.45567
R461 source.n406 source.n405 9.45567
R462 source.n336 source.n335 9.45567
R463 source.n64 source.n63 9.45567
R464 source.n134 source.n133 9.45567
R465 source.n200 source.n199 9.45567
R466 source.n270 source.n269 9.45567
R467 source.n541 source.n540 9.3005
R468 source.n480 source.n479 9.3005
R469 source.n535 source.n534 9.3005
R470 source.n533 source.n532 9.3005
R471 source.n484 source.n483 9.3005
R472 source.n527 source.n526 9.3005
R473 source.n525 source.n524 9.3005
R474 source.n501 source.n500 9.3005
R475 source.n496 source.n495 9.3005
R476 source.n507 source.n506 9.3005
R477 source.n509 source.n508 9.3005
R478 source.n492 source.n491 9.3005
R479 source.n515 source.n514 9.3005
R480 source.n517 source.n516 9.3005
R481 source.n518 source.n487 9.3005
R482 source.n471 source.n470 9.3005
R483 source.n410 source.n409 9.3005
R484 source.n465 source.n464 9.3005
R485 source.n463 source.n462 9.3005
R486 source.n414 source.n413 9.3005
R487 source.n457 source.n456 9.3005
R488 source.n455 source.n454 9.3005
R489 source.n431 source.n430 9.3005
R490 source.n426 source.n425 9.3005
R491 source.n437 source.n436 9.3005
R492 source.n439 source.n438 9.3005
R493 source.n422 source.n421 9.3005
R494 source.n445 source.n444 9.3005
R495 source.n447 source.n446 9.3005
R496 source.n448 source.n417 9.3005
R497 source.n405 source.n404 9.3005
R498 source.n344 source.n343 9.3005
R499 source.n399 source.n398 9.3005
R500 source.n397 source.n396 9.3005
R501 source.n348 source.n347 9.3005
R502 source.n391 source.n390 9.3005
R503 source.n389 source.n388 9.3005
R504 source.n365 source.n364 9.3005
R505 source.n360 source.n359 9.3005
R506 source.n371 source.n370 9.3005
R507 source.n373 source.n372 9.3005
R508 source.n356 source.n355 9.3005
R509 source.n379 source.n378 9.3005
R510 source.n381 source.n380 9.3005
R511 source.n382 source.n351 9.3005
R512 source.n335 source.n334 9.3005
R513 source.n274 source.n273 9.3005
R514 source.n329 source.n328 9.3005
R515 source.n327 source.n326 9.3005
R516 source.n278 source.n277 9.3005
R517 source.n321 source.n320 9.3005
R518 source.n319 source.n318 9.3005
R519 source.n295 source.n294 9.3005
R520 source.n290 source.n289 9.3005
R521 source.n301 source.n300 9.3005
R522 source.n303 source.n302 9.3005
R523 source.n286 source.n285 9.3005
R524 source.n309 source.n308 9.3005
R525 source.n311 source.n310 9.3005
R526 source.n312 source.n281 9.3005
R527 source.n24 source.n23 9.3005
R528 source.n19 source.n18 9.3005
R529 source.n30 source.n29 9.3005
R530 source.n32 source.n31 9.3005
R531 source.n15 source.n14 9.3005
R532 source.n38 source.n37 9.3005
R533 source.n40 source.n39 9.3005
R534 source.n12 source.n9 9.3005
R535 source.n63 source.n62 9.3005
R536 source.n2 source.n1 9.3005
R537 source.n57 source.n56 9.3005
R538 source.n55 source.n54 9.3005
R539 source.n6 source.n5 9.3005
R540 source.n49 source.n48 9.3005
R541 source.n47 source.n46 9.3005
R542 source.n94 source.n93 9.3005
R543 source.n89 source.n88 9.3005
R544 source.n100 source.n99 9.3005
R545 source.n102 source.n101 9.3005
R546 source.n85 source.n84 9.3005
R547 source.n108 source.n107 9.3005
R548 source.n110 source.n109 9.3005
R549 source.n82 source.n79 9.3005
R550 source.n133 source.n132 9.3005
R551 source.n72 source.n71 9.3005
R552 source.n127 source.n126 9.3005
R553 source.n125 source.n124 9.3005
R554 source.n76 source.n75 9.3005
R555 source.n119 source.n118 9.3005
R556 source.n117 source.n116 9.3005
R557 source.n160 source.n159 9.3005
R558 source.n155 source.n154 9.3005
R559 source.n166 source.n165 9.3005
R560 source.n168 source.n167 9.3005
R561 source.n151 source.n150 9.3005
R562 source.n174 source.n173 9.3005
R563 source.n176 source.n175 9.3005
R564 source.n148 source.n145 9.3005
R565 source.n199 source.n198 9.3005
R566 source.n138 source.n137 9.3005
R567 source.n193 source.n192 9.3005
R568 source.n191 source.n190 9.3005
R569 source.n142 source.n141 9.3005
R570 source.n185 source.n184 9.3005
R571 source.n183 source.n182 9.3005
R572 source.n230 source.n229 9.3005
R573 source.n225 source.n224 9.3005
R574 source.n236 source.n235 9.3005
R575 source.n238 source.n237 9.3005
R576 source.n221 source.n220 9.3005
R577 source.n244 source.n243 9.3005
R578 source.n246 source.n245 9.3005
R579 source.n218 source.n215 9.3005
R580 source.n269 source.n268 9.3005
R581 source.n208 source.n207 9.3005
R582 source.n263 source.n262 9.3005
R583 source.n261 source.n260 9.3005
R584 source.n212 source.n211 9.3005
R585 source.n255 source.n254 9.3005
R586 source.n253 source.n252 9.3005
R587 source.n506 source.n505 8.92171
R588 source.n539 source.n480 8.92171
R589 source.n436 source.n435 8.92171
R590 source.n469 source.n410 8.92171
R591 source.n370 source.n369 8.92171
R592 source.n403 source.n344 8.92171
R593 source.n300 source.n299 8.92171
R594 source.n333 source.n274 8.92171
R595 source.n61 source.n2 8.92171
R596 source.n29 source.n28 8.92171
R597 source.n131 source.n72 8.92171
R598 source.n99 source.n98 8.92171
R599 source.n197 source.n138 8.92171
R600 source.n165 source.n164 8.92171
R601 source.n267 source.n208 8.92171
R602 source.n235 source.n234 8.92171
R603 source.n502 source.n496 8.14595
R604 source.n540 source.n478 8.14595
R605 source.n432 source.n426 8.14595
R606 source.n470 source.n408 8.14595
R607 source.n366 source.n360 8.14595
R608 source.n404 source.n342 8.14595
R609 source.n296 source.n290 8.14595
R610 source.n334 source.n272 8.14595
R611 source.n62 source.n0 8.14595
R612 source.n25 source.n19 8.14595
R613 source.n132 source.n70 8.14595
R614 source.n95 source.n89 8.14595
R615 source.n198 source.n136 8.14595
R616 source.n161 source.n155 8.14595
R617 source.n268 source.n206 8.14595
R618 source.n231 source.n225 8.14595
R619 source.n501 source.n498 7.3702
R620 source.n431 source.n428 7.3702
R621 source.n365 source.n362 7.3702
R622 source.n295 source.n292 7.3702
R623 source.n24 source.n21 7.3702
R624 source.n94 source.n91 7.3702
R625 source.n160 source.n157 7.3702
R626 source.n230 source.n227 7.3702
R627 source.n502 source.n501 5.81868
R628 source.n542 source.n478 5.81868
R629 source.n432 source.n431 5.81868
R630 source.n472 source.n408 5.81868
R631 source.n366 source.n365 5.81868
R632 source.n406 source.n342 5.81868
R633 source.n296 source.n295 5.81868
R634 source.n336 source.n272 5.81868
R635 source.n64 source.n0 5.81868
R636 source.n25 source.n24 5.81868
R637 source.n134 source.n70 5.81868
R638 source.n95 source.n94 5.81868
R639 source.n200 source.n136 5.81868
R640 source.n161 source.n160 5.81868
R641 source.n270 source.n206 5.81868
R642 source.n231 source.n230 5.81868
R643 source.n544 source.n543 5.62119
R644 source.n505 source.n496 5.04292
R645 source.n540 source.n539 5.04292
R646 source.n435 source.n426 5.04292
R647 source.n470 source.n469 5.04292
R648 source.n369 source.n360 5.04292
R649 source.n404 source.n403 5.04292
R650 source.n299 source.n290 5.04292
R651 source.n334 source.n333 5.04292
R652 source.n62 source.n61 5.04292
R653 source.n28 source.n19 5.04292
R654 source.n132 source.n131 5.04292
R655 source.n98 source.n89 5.04292
R656 source.n198 source.n197 5.04292
R657 source.n164 source.n155 5.04292
R658 source.n268 source.n267 5.04292
R659 source.n234 source.n225 5.04292
R660 source.n506 source.n494 4.26717
R661 source.n536 source.n480 4.26717
R662 source.n436 source.n424 4.26717
R663 source.n466 source.n410 4.26717
R664 source.n370 source.n358 4.26717
R665 source.n400 source.n344 4.26717
R666 source.n300 source.n288 4.26717
R667 source.n330 source.n274 4.26717
R668 source.n58 source.n2 4.26717
R669 source.n29 source.n17 4.26717
R670 source.n128 source.n72 4.26717
R671 source.n99 source.n87 4.26717
R672 source.n194 source.n138 4.26717
R673 source.n165 source.n153 4.26717
R674 source.n264 source.n208 4.26717
R675 source.n235 source.n223 4.26717
R676 source.n510 source.n509 3.49141
R677 source.n535 source.n482 3.49141
R678 source.n440 source.n439 3.49141
R679 source.n465 source.n412 3.49141
R680 source.n374 source.n373 3.49141
R681 source.n399 source.n346 3.49141
R682 source.n304 source.n303 3.49141
R683 source.n329 source.n276 3.49141
R684 source.n57 source.n4 3.49141
R685 source.n33 source.n32 3.49141
R686 source.n127 source.n74 3.49141
R687 source.n103 source.n102 3.49141
R688 source.n193 source.n140 3.49141
R689 source.n169 source.n168 3.49141
R690 source.n263 source.n210 3.49141
R691 source.n239 source.n238 3.49141
R692 source.n500 source.n499 2.84303
R693 source.n430 source.n429 2.84303
R694 source.n364 source.n363 2.84303
R695 source.n294 source.n293 2.84303
R696 source.n23 source.n22 2.84303
R697 source.n93 source.n92 2.84303
R698 source.n159 source.n158 2.84303
R699 source.n229 source.n228 2.84303
R700 source.n513 source.n492 2.71565
R701 source.n532 source.n531 2.71565
R702 source.n443 source.n422 2.71565
R703 source.n462 source.n461 2.71565
R704 source.n377 source.n356 2.71565
R705 source.n396 source.n395 2.71565
R706 source.n307 source.n286 2.71565
R707 source.n326 source.n325 2.71565
R708 source.n54 source.n53 2.71565
R709 source.n36 source.n15 2.71565
R710 source.n124 source.n123 2.71565
R711 source.n106 source.n85 2.71565
R712 source.n190 source.n189 2.71565
R713 source.n172 source.n151 2.71565
R714 source.n260 source.n259 2.71565
R715 source.n242 source.n221 2.71565
R716 source.n514 source.n490 1.93989
R717 source.n528 source.n484 1.93989
R718 source.n444 source.n420 1.93989
R719 source.n458 source.n414 1.93989
R720 source.n378 source.n354 1.93989
R721 source.n392 source.n348 1.93989
R722 source.n308 source.n284 1.93989
R723 source.n322 source.n278 1.93989
R724 source.n50 source.n6 1.93989
R725 source.n37 source.n13 1.93989
R726 source.n120 source.n76 1.93989
R727 source.n107 source.n83 1.93989
R728 source.n186 source.n142 1.93989
R729 source.n173 source.n149 1.93989
R730 source.n256 source.n212 1.93989
R731 source.n243 source.n219 1.93989
R732 source.n476 source.t0 1.6505
R733 source.n476 source.t6 1.6505
R734 source.n474 source.t7 1.6505
R735 source.n474 source.t23 1.6505
R736 source.n340 source.t16 1.6505
R737 source.n340 source.t10 1.6505
R738 source.n338 source.t18 1.6505
R739 source.n338 source.t19 1.6505
R740 source.n66 source.t15 1.6505
R741 source.n66 source.t12 1.6505
R742 source.n68 source.t13 1.6505
R743 source.n68 source.t9 1.6505
R744 source.n202 source.t22 1.6505
R745 source.n202 source.t4 1.6505
R746 source.n204 source.t5 1.6505
R747 source.n204 source.t21 1.6505
R748 source.n519 source.n517 1.16414
R749 source.n527 source.n486 1.16414
R750 source.n449 source.n447 1.16414
R751 source.n457 source.n416 1.16414
R752 source.n383 source.n381 1.16414
R753 source.n391 source.n350 1.16414
R754 source.n313 source.n311 1.16414
R755 source.n321 source.n280 1.16414
R756 source.n49 source.n8 1.16414
R757 source.n41 source.n40 1.16414
R758 source.n119 source.n78 1.16414
R759 source.n111 source.n110 1.16414
R760 source.n185 source.n144 1.16414
R761 source.n177 source.n176 1.16414
R762 source.n255 source.n214 1.16414
R763 source.n247 source.n246 1.16414
R764 source.n271 source.n205 0.716017
R765 source.n205 source.n203 0.716017
R766 source.n203 source.n201 0.716017
R767 source.n135 source.n69 0.716017
R768 source.n69 source.n67 0.716017
R769 source.n67 source.n65 0.716017
R770 source.n339 source.n337 0.716017
R771 source.n341 source.n339 0.716017
R772 source.n407 source.n341 0.716017
R773 source.n475 source.n473 0.716017
R774 source.n477 source.n475 0.716017
R775 source.n543 source.n477 0.716017
R776 source.n201 source.n135 0.470328
R777 source.n473 source.n407 0.470328
R778 source.n518 source.n488 0.388379
R779 source.n524 source.n523 0.388379
R780 source.n448 source.n418 0.388379
R781 source.n454 source.n453 0.388379
R782 source.n382 source.n352 0.388379
R783 source.n388 source.n387 0.388379
R784 source.n312 source.n282 0.388379
R785 source.n318 source.n317 0.388379
R786 source.n46 source.n45 0.388379
R787 source.n12 source.n10 0.388379
R788 source.n116 source.n115 0.388379
R789 source.n82 source.n80 0.388379
R790 source.n182 source.n181 0.388379
R791 source.n148 source.n146 0.388379
R792 source.n252 source.n251 0.388379
R793 source.n218 source.n216 0.388379
R794 source source.n544 0.188
R795 source.n500 source.n495 0.155672
R796 source.n507 source.n495 0.155672
R797 source.n508 source.n507 0.155672
R798 source.n508 source.n491 0.155672
R799 source.n515 source.n491 0.155672
R800 source.n516 source.n515 0.155672
R801 source.n516 source.n487 0.155672
R802 source.n525 source.n487 0.155672
R803 source.n526 source.n525 0.155672
R804 source.n526 source.n483 0.155672
R805 source.n533 source.n483 0.155672
R806 source.n534 source.n533 0.155672
R807 source.n534 source.n479 0.155672
R808 source.n541 source.n479 0.155672
R809 source.n430 source.n425 0.155672
R810 source.n437 source.n425 0.155672
R811 source.n438 source.n437 0.155672
R812 source.n438 source.n421 0.155672
R813 source.n445 source.n421 0.155672
R814 source.n446 source.n445 0.155672
R815 source.n446 source.n417 0.155672
R816 source.n455 source.n417 0.155672
R817 source.n456 source.n455 0.155672
R818 source.n456 source.n413 0.155672
R819 source.n463 source.n413 0.155672
R820 source.n464 source.n463 0.155672
R821 source.n464 source.n409 0.155672
R822 source.n471 source.n409 0.155672
R823 source.n364 source.n359 0.155672
R824 source.n371 source.n359 0.155672
R825 source.n372 source.n371 0.155672
R826 source.n372 source.n355 0.155672
R827 source.n379 source.n355 0.155672
R828 source.n380 source.n379 0.155672
R829 source.n380 source.n351 0.155672
R830 source.n389 source.n351 0.155672
R831 source.n390 source.n389 0.155672
R832 source.n390 source.n347 0.155672
R833 source.n397 source.n347 0.155672
R834 source.n398 source.n397 0.155672
R835 source.n398 source.n343 0.155672
R836 source.n405 source.n343 0.155672
R837 source.n294 source.n289 0.155672
R838 source.n301 source.n289 0.155672
R839 source.n302 source.n301 0.155672
R840 source.n302 source.n285 0.155672
R841 source.n309 source.n285 0.155672
R842 source.n310 source.n309 0.155672
R843 source.n310 source.n281 0.155672
R844 source.n319 source.n281 0.155672
R845 source.n320 source.n319 0.155672
R846 source.n320 source.n277 0.155672
R847 source.n327 source.n277 0.155672
R848 source.n328 source.n327 0.155672
R849 source.n328 source.n273 0.155672
R850 source.n335 source.n273 0.155672
R851 source.n63 source.n1 0.155672
R852 source.n56 source.n1 0.155672
R853 source.n56 source.n55 0.155672
R854 source.n55 source.n5 0.155672
R855 source.n48 source.n5 0.155672
R856 source.n48 source.n47 0.155672
R857 source.n47 source.n9 0.155672
R858 source.n39 source.n9 0.155672
R859 source.n39 source.n38 0.155672
R860 source.n38 source.n14 0.155672
R861 source.n31 source.n14 0.155672
R862 source.n31 source.n30 0.155672
R863 source.n30 source.n18 0.155672
R864 source.n23 source.n18 0.155672
R865 source.n133 source.n71 0.155672
R866 source.n126 source.n71 0.155672
R867 source.n126 source.n125 0.155672
R868 source.n125 source.n75 0.155672
R869 source.n118 source.n75 0.155672
R870 source.n118 source.n117 0.155672
R871 source.n117 source.n79 0.155672
R872 source.n109 source.n79 0.155672
R873 source.n109 source.n108 0.155672
R874 source.n108 source.n84 0.155672
R875 source.n101 source.n84 0.155672
R876 source.n101 source.n100 0.155672
R877 source.n100 source.n88 0.155672
R878 source.n93 source.n88 0.155672
R879 source.n199 source.n137 0.155672
R880 source.n192 source.n137 0.155672
R881 source.n192 source.n191 0.155672
R882 source.n191 source.n141 0.155672
R883 source.n184 source.n141 0.155672
R884 source.n184 source.n183 0.155672
R885 source.n183 source.n145 0.155672
R886 source.n175 source.n145 0.155672
R887 source.n175 source.n174 0.155672
R888 source.n174 source.n150 0.155672
R889 source.n167 source.n150 0.155672
R890 source.n167 source.n166 0.155672
R891 source.n166 source.n154 0.155672
R892 source.n159 source.n154 0.155672
R893 source.n269 source.n207 0.155672
R894 source.n262 source.n207 0.155672
R895 source.n262 source.n261 0.155672
R896 source.n261 source.n211 0.155672
R897 source.n254 source.n211 0.155672
R898 source.n254 source.n253 0.155672
R899 source.n253 source.n215 0.155672
R900 source.n245 source.n215 0.155672
R901 source.n245 source.n244 0.155672
R902 source.n244 source.n220 0.155672
R903 source.n237 source.n220 0.155672
R904 source.n237 source.n236 0.155672
R905 source.n236 source.n224 0.155672
R906 source.n229 source.n224 0.155672
R907 minus.n3 minus.t10 683.635
R908 minus.n17 minus.t1 683.635
R909 minus.n4 minus.t2 656.966
R910 minus.n5 minus.t5 656.966
R911 minus.n1 minus.t11 656.966
R912 minus.n10 minus.t4 656.966
R913 minus.n12 minus.t8 656.966
R914 minus.n18 minus.t0 656.966
R915 minus.n19 minus.t7 656.966
R916 minus.n15 minus.t6 656.966
R917 minus.n24 minus.t3 656.966
R918 minus.n26 minus.t9 656.966
R919 minus.n13 minus.n12 161.3
R920 minus.n11 minus.n0 161.3
R921 minus.n10 minus.n9 161.3
R922 minus.n8 minus.n1 161.3
R923 minus.n7 minus.n6 161.3
R924 minus.n5 minus.n2 161.3
R925 minus.n27 minus.n26 161.3
R926 minus.n25 minus.n14 161.3
R927 minus.n24 minus.n23 161.3
R928 minus.n22 minus.n15 161.3
R929 minus.n21 minus.n20 161.3
R930 minus.n19 minus.n16 161.3
R931 minus.n5 minus.n4 48.2005
R932 minus.n10 minus.n1 48.2005
R933 minus.n19 minus.n18 48.2005
R934 minus.n24 minus.n15 48.2005
R935 minus.n12 minus.n11 47.4702
R936 minus.n26 minus.n25 47.4702
R937 minus.n3 minus.n2 45.1192
R938 minus.n17 minus.n16 45.1192
R939 minus.n28 minus.n13 36.2656
R940 minus.n6 minus.n1 24.1005
R941 minus.n6 minus.n5 24.1005
R942 minus.n20 minus.n19 24.1005
R943 minus.n20 minus.n15 24.1005
R944 minus.n4 minus.n3 13.6377
R945 minus.n18 minus.n17 13.6377
R946 minus.n28 minus.n27 6.5308
R947 minus.n11 minus.n10 0.730803
R948 minus.n25 minus.n24 0.730803
R949 minus.n13 minus.n0 0.189894
R950 minus.n9 minus.n0 0.189894
R951 minus.n9 minus.n8 0.189894
R952 minus.n8 minus.n7 0.189894
R953 minus.n7 minus.n2 0.189894
R954 minus.n21 minus.n16 0.189894
R955 minus.n22 minus.n21 0.189894
R956 minus.n23 minus.n22 0.189894
R957 minus.n23 minus.n14 0.189894
R958 minus.n27 minus.n14 0.189894
R959 minus minus.n28 0.188
R960 drain_right.n6 drain_right.n4 60.268
R961 drain_right.n3 drain_right.n2 60.2127
R962 drain_right.n3 drain_right.n0 60.2127
R963 drain_right.n6 drain_right.n5 59.5527
R964 drain_right.n8 drain_right.n7 59.5527
R965 drain_right.n3 drain_right.n1 59.5525
R966 drain_right drain_right.n3 30.3914
R967 drain_right drain_right.n8 6.36873
R968 drain_right.n1 drain_right.t4 1.6505
R969 drain_right.n1 drain_right.t5 1.6505
R970 drain_right.n2 drain_right.t8 1.6505
R971 drain_right.n2 drain_right.t2 1.6505
R972 drain_right.n0 drain_right.t10 1.6505
R973 drain_right.n0 drain_right.t11 1.6505
R974 drain_right.n4 drain_right.t9 1.6505
R975 drain_right.n4 drain_right.t1 1.6505
R976 drain_right.n5 drain_right.t0 1.6505
R977 drain_right.n5 drain_right.t6 1.6505
R978 drain_right.n7 drain_right.t3 1.6505
R979 drain_right.n7 drain_right.t7 1.6505
R980 drain_right.n8 drain_right.n6 0.716017
C0 drain_right minus 6.4779f
C1 source drain_left 18.3029f
C2 source minus 6.24641f
C3 drain_right source 18.303902f
C4 plus drain_left 6.66049f
C5 minus plus 5.49323f
C6 drain_right plus 0.337327f
C7 source plus 6.26044f
C8 minus drain_left 0.171641f
C9 drain_right drain_left 0.936346f
C10 drain_right a_n1878_n3288# 6.08602f
C11 drain_left a_n1878_n3288# 6.36857f
C12 source a_n1878_n3288# 8.881788f
C13 minus a_n1878_n3288# 7.361398f
C14 plus a_n1878_n3288# 9.19608f
C15 drain_right.t10 a_n1878_n3288# 0.276564f
C16 drain_right.t11 a_n1878_n3288# 0.276564f
C17 drain_right.n0 a_n1878_n3288# 2.46524f
C18 drain_right.t4 a_n1878_n3288# 0.276564f
C19 drain_right.t5 a_n1878_n3288# 0.276564f
C20 drain_right.n1 a_n1878_n3288# 2.46099f
C21 drain_right.t8 a_n1878_n3288# 0.276564f
C22 drain_right.t2 a_n1878_n3288# 0.276564f
C23 drain_right.n2 a_n1878_n3288# 2.46524f
C24 drain_right.n3 a_n1878_n3288# 2.4711f
C25 drain_right.t9 a_n1878_n3288# 0.276564f
C26 drain_right.t1 a_n1878_n3288# 0.276564f
C27 drain_right.n4 a_n1878_n3288# 2.46564f
C28 drain_right.t0 a_n1878_n3288# 0.276564f
C29 drain_right.t6 a_n1878_n3288# 0.276564f
C30 drain_right.n5 a_n1878_n3288# 2.461f
C31 drain_right.n6 a_n1878_n3288# 0.765597f
C32 drain_right.t3 a_n1878_n3288# 0.276564f
C33 drain_right.t7 a_n1878_n3288# 0.276564f
C34 drain_right.n7 a_n1878_n3288# 2.461f
C35 drain_right.n8 a_n1878_n3288# 0.629809f
C36 minus.n0 a_n1878_n3288# 0.046443f
C37 minus.t11 a_n1878_n3288# 0.794595f
C38 minus.n1 a_n1878_n3288# 0.325249f
C39 minus.t4 a_n1878_n3288# 0.794595f
C40 minus.n2 a_n1878_n3288# 0.189145f
C41 minus.t10 a_n1878_n3288# 0.807101f
C42 minus.n3 a_n1878_n3288# 0.309156f
C43 minus.t2 a_n1878_n3288# 0.794595f
C44 minus.n4 a_n1878_n3288# 0.330847f
C45 minus.t5 a_n1878_n3288# 0.794595f
C46 minus.n5 a_n1878_n3288# 0.325249f
C47 minus.n6 a_n1878_n3288# 0.010539f
C48 minus.n7 a_n1878_n3288# 0.046443f
C49 minus.n8 a_n1878_n3288# 0.046443f
C50 minus.n9 a_n1878_n3288# 0.046443f
C51 minus.n10 a_n1878_n3288# 0.320667f
C52 minus.n11 a_n1878_n3288# 0.010539f
C53 minus.t8 a_n1878_n3288# 0.794595f
C54 minus.n12 a_n1878_n3288# 0.320381f
C55 minus.n13 a_n1878_n3288# 1.64754f
C56 minus.n14 a_n1878_n3288# 0.046443f
C57 minus.t6 a_n1878_n3288# 0.794595f
C58 minus.n15 a_n1878_n3288# 0.325249f
C59 minus.n16 a_n1878_n3288# 0.189145f
C60 minus.t1 a_n1878_n3288# 0.807101f
C61 minus.n17 a_n1878_n3288# 0.309156f
C62 minus.t0 a_n1878_n3288# 0.794595f
C63 minus.n18 a_n1878_n3288# 0.330847f
C64 minus.t7 a_n1878_n3288# 0.794595f
C65 minus.n19 a_n1878_n3288# 0.325249f
C66 minus.n20 a_n1878_n3288# 0.010539f
C67 minus.n21 a_n1878_n3288# 0.046443f
C68 minus.n22 a_n1878_n3288# 0.046443f
C69 minus.n23 a_n1878_n3288# 0.046443f
C70 minus.t3 a_n1878_n3288# 0.794595f
C71 minus.n24 a_n1878_n3288# 0.320667f
C72 minus.n25 a_n1878_n3288# 0.010539f
C73 minus.t9 a_n1878_n3288# 0.794595f
C74 minus.n26 a_n1878_n3288# 0.320381f
C75 minus.n27 a_n1878_n3288# 0.306997f
C76 minus.n28 a_n1878_n3288# 1.99972f
C77 source.n0 a_n1878_n3288# 0.030955f
C78 source.n1 a_n1878_n3288# 0.023369f
C79 source.n2 a_n1878_n3288# 0.012557f
C80 source.n3 a_n1878_n3288# 0.029681f
C81 source.n4 a_n1878_n3288# 0.013296f
C82 source.n5 a_n1878_n3288# 0.023369f
C83 source.n6 a_n1878_n3288# 0.012557f
C84 source.n7 a_n1878_n3288# 0.029681f
C85 source.n8 a_n1878_n3288# 0.013296f
C86 source.n9 a_n1878_n3288# 0.023369f
C87 source.n10 a_n1878_n3288# 0.012927f
C88 source.n11 a_n1878_n3288# 0.029681f
C89 source.n12 a_n1878_n3288# 0.012557f
C90 source.n13 a_n1878_n3288# 0.013296f
C91 source.n14 a_n1878_n3288# 0.023369f
C92 source.n15 a_n1878_n3288# 0.012557f
C93 source.n16 a_n1878_n3288# 0.029681f
C94 source.n17 a_n1878_n3288# 0.013296f
C95 source.n18 a_n1878_n3288# 0.023369f
C96 source.n19 a_n1878_n3288# 0.012557f
C97 source.n20 a_n1878_n3288# 0.022261f
C98 source.n21 a_n1878_n3288# 0.020982f
C99 source.t8 a_n1878_n3288# 0.050129f
C100 source.n22 a_n1878_n3288# 0.168486f
C101 source.n23 a_n1878_n3288# 1.17891f
C102 source.n24 a_n1878_n3288# 0.012557f
C103 source.n25 a_n1878_n3288# 0.013296f
C104 source.n26 a_n1878_n3288# 0.029681f
C105 source.n27 a_n1878_n3288# 0.029681f
C106 source.n28 a_n1878_n3288# 0.013296f
C107 source.n29 a_n1878_n3288# 0.012557f
C108 source.n30 a_n1878_n3288# 0.023369f
C109 source.n31 a_n1878_n3288# 0.023369f
C110 source.n32 a_n1878_n3288# 0.012557f
C111 source.n33 a_n1878_n3288# 0.013296f
C112 source.n34 a_n1878_n3288# 0.029681f
C113 source.n35 a_n1878_n3288# 0.029681f
C114 source.n36 a_n1878_n3288# 0.013296f
C115 source.n37 a_n1878_n3288# 0.012557f
C116 source.n38 a_n1878_n3288# 0.023369f
C117 source.n39 a_n1878_n3288# 0.023369f
C118 source.n40 a_n1878_n3288# 0.012557f
C119 source.n41 a_n1878_n3288# 0.013296f
C120 source.n42 a_n1878_n3288# 0.029681f
C121 source.n43 a_n1878_n3288# 0.029681f
C122 source.n44 a_n1878_n3288# 0.029681f
C123 source.n45 a_n1878_n3288# 0.012927f
C124 source.n46 a_n1878_n3288# 0.012557f
C125 source.n47 a_n1878_n3288# 0.023369f
C126 source.n48 a_n1878_n3288# 0.023369f
C127 source.n49 a_n1878_n3288# 0.012557f
C128 source.n50 a_n1878_n3288# 0.013296f
C129 source.n51 a_n1878_n3288# 0.029681f
C130 source.n52 a_n1878_n3288# 0.029681f
C131 source.n53 a_n1878_n3288# 0.013296f
C132 source.n54 a_n1878_n3288# 0.012557f
C133 source.n55 a_n1878_n3288# 0.023369f
C134 source.n56 a_n1878_n3288# 0.023369f
C135 source.n57 a_n1878_n3288# 0.012557f
C136 source.n58 a_n1878_n3288# 0.013296f
C137 source.n59 a_n1878_n3288# 0.029681f
C138 source.n60 a_n1878_n3288# 0.060908f
C139 source.n61 a_n1878_n3288# 0.013296f
C140 source.n62 a_n1878_n3288# 0.012557f
C141 source.n63 a_n1878_n3288# 0.050185f
C142 source.n64 a_n1878_n3288# 0.033615f
C143 source.n65 a_n1878_n3288# 0.961764f
C144 source.t15 a_n1878_n3288# 0.2216f
C145 source.t12 a_n1878_n3288# 0.2216f
C146 source.n66 a_n1878_n3288# 1.89734f
C147 source.n67 a_n1878_n3288# 0.346671f
C148 source.t13 a_n1878_n3288# 0.2216f
C149 source.t9 a_n1878_n3288# 0.2216f
C150 source.n68 a_n1878_n3288# 1.89734f
C151 source.n69 a_n1878_n3288# 0.346671f
C152 source.n70 a_n1878_n3288# 0.030955f
C153 source.n71 a_n1878_n3288# 0.023369f
C154 source.n72 a_n1878_n3288# 0.012557f
C155 source.n73 a_n1878_n3288# 0.029681f
C156 source.n74 a_n1878_n3288# 0.013296f
C157 source.n75 a_n1878_n3288# 0.023369f
C158 source.n76 a_n1878_n3288# 0.012557f
C159 source.n77 a_n1878_n3288# 0.029681f
C160 source.n78 a_n1878_n3288# 0.013296f
C161 source.n79 a_n1878_n3288# 0.023369f
C162 source.n80 a_n1878_n3288# 0.012927f
C163 source.n81 a_n1878_n3288# 0.029681f
C164 source.n82 a_n1878_n3288# 0.012557f
C165 source.n83 a_n1878_n3288# 0.013296f
C166 source.n84 a_n1878_n3288# 0.023369f
C167 source.n85 a_n1878_n3288# 0.012557f
C168 source.n86 a_n1878_n3288# 0.029681f
C169 source.n87 a_n1878_n3288# 0.013296f
C170 source.n88 a_n1878_n3288# 0.023369f
C171 source.n89 a_n1878_n3288# 0.012557f
C172 source.n90 a_n1878_n3288# 0.022261f
C173 source.n91 a_n1878_n3288# 0.020982f
C174 source.t17 a_n1878_n3288# 0.050129f
C175 source.n92 a_n1878_n3288# 0.168486f
C176 source.n93 a_n1878_n3288# 1.17891f
C177 source.n94 a_n1878_n3288# 0.012557f
C178 source.n95 a_n1878_n3288# 0.013296f
C179 source.n96 a_n1878_n3288# 0.029681f
C180 source.n97 a_n1878_n3288# 0.029681f
C181 source.n98 a_n1878_n3288# 0.013296f
C182 source.n99 a_n1878_n3288# 0.012557f
C183 source.n100 a_n1878_n3288# 0.023369f
C184 source.n101 a_n1878_n3288# 0.023369f
C185 source.n102 a_n1878_n3288# 0.012557f
C186 source.n103 a_n1878_n3288# 0.013296f
C187 source.n104 a_n1878_n3288# 0.029681f
C188 source.n105 a_n1878_n3288# 0.029681f
C189 source.n106 a_n1878_n3288# 0.013296f
C190 source.n107 a_n1878_n3288# 0.012557f
C191 source.n108 a_n1878_n3288# 0.023369f
C192 source.n109 a_n1878_n3288# 0.023369f
C193 source.n110 a_n1878_n3288# 0.012557f
C194 source.n111 a_n1878_n3288# 0.013296f
C195 source.n112 a_n1878_n3288# 0.029681f
C196 source.n113 a_n1878_n3288# 0.029681f
C197 source.n114 a_n1878_n3288# 0.029681f
C198 source.n115 a_n1878_n3288# 0.012927f
C199 source.n116 a_n1878_n3288# 0.012557f
C200 source.n117 a_n1878_n3288# 0.023369f
C201 source.n118 a_n1878_n3288# 0.023369f
C202 source.n119 a_n1878_n3288# 0.012557f
C203 source.n120 a_n1878_n3288# 0.013296f
C204 source.n121 a_n1878_n3288# 0.029681f
C205 source.n122 a_n1878_n3288# 0.029681f
C206 source.n123 a_n1878_n3288# 0.013296f
C207 source.n124 a_n1878_n3288# 0.012557f
C208 source.n125 a_n1878_n3288# 0.023369f
C209 source.n126 a_n1878_n3288# 0.023369f
C210 source.n127 a_n1878_n3288# 0.012557f
C211 source.n128 a_n1878_n3288# 0.013296f
C212 source.n129 a_n1878_n3288# 0.029681f
C213 source.n130 a_n1878_n3288# 0.060908f
C214 source.n131 a_n1878_n3288# 0.013296f
C215 source.n132 a_n1878_n3288# 0.012557f
C216 source.n133 a_n1878_n3288# 0.050185f
C217 source.n134 a_n1878_n3288# 0.033615f
C218 source.n135 a_n1878_n3288# 0.107056f
C219 source.n136 a_n1878_n3288# 0.030955f
C220 source.n137 a_n1878_n3288# 0.023369f
C221 source.n138 a_n1878_n3288# 0.012557f
C222 source.n139 a_n1878_n3288# 0.029681f
C223 source.n140 a_n1878_n3288# 0.013296f
C224 source.n141 a_n1878_n3288# 0.023369f
C225 source.n142 a_n1878_n3288# 0.012557f
C226 source.n143 a_n1878_n3288# 0.029681f
C227 source.n144 a_n1878_n3288# 0.013296f
C228 source.n145 a_n1878_n3288# 0.023369f
C229 source.n146 a_n1878_n3288# 0.012927f
C230 source.n147 a_n1878_n3288# 0.029681f
C231 source.n148 a_n1878_n3288# 0.012557f
C232 source.n149 a_n1878_n3288# 0.013296f
C233 source.n150 a_n1878_n3288# 0.023369f
C234 source.n151 a_n1878_n3288# 0.012557f
C235 source.n152 a_n1878_n3288# 0.029681f
C236 source.n153 a_n1878_n3288# 0.013296f
C237 source.n154 a_n1878_n3288# 0.023369f
C238 source.n155 a_n1878_n3288# 0.012557f
C239 source.n156 a_n1878_n3288# 0.022261f
C240 source.n157 a_n1878_n3288# 0.020982f
C241 source.t20 a_n1878_n3288# 0.050129f
C242 source.n158 a_n1878_n3288# 0.168486f
C243 source.n159 a_n1878_n3288# 1.17891f
C244 source.n160 a_n1878_n3288# 0.012557f
C245 source.n161 a_n1878_n3288# 0.013296f
C246 source.n162 a_n1878_n3288# 0.029681f
C247 source.n163 a_n1878_n3288# 0.029681f
C248 source.n164 a_n1878_n3288# 0.013296f
C249 source.n165 a_n1878_n3288# 0.012557f
C250 source.n166 a_n1878_n3288# 0.023369f
C251 source.n167 a_n1878_n3288# 0.023369f
C252 source.n168 a_n1878_n3288# 0.012557f
C253 source.n169 a_n1878_n3288# 0.013296f
C254 source.n170 a_n1878_n3288# 0.029681f
C255 source.n171 a_n1878_n3288# 0.029681f
C256 source.n172 a_n1878_n3288# 0.013296f
C257 source.n173 a_n1878_n3288# 0.012557f
C258 source.n174 a_n1878_n3288# 0.023369f
C259 source.n175 a_n1878_n3288# 0.023369f
C260 source.n176 a_n1878_n3288# 0.012557f
C261 source.n177 a_n1878_n3288# 0.013296f
C262 source.n178 a_n1878_n3288# 0.029681f
C263 source.n179 a_n1878_n3288# 0.029681f
C264 source.n180 a_n1878_n3288# 0.029681f
C265 source.n181 a_n1878_n3288# 0.012927f
C266 source.n182 a_n1878_n3288# 0.012557f
C267 source.n183 a_n1878_n3288# 0.023369f
C268 source.n184 a_n1878_n3288# 0.023369f
C269 source.n185 a_n1878_n3288# 0.012557f
C270 source.n186 a_n1878_n3288# 0.013296f
C271 source.n187 a_n1878_n3288# 0.029681f
C272 source.n188 a_n1878_n3288# 0.029681f
C273 source.n189 a_n1878_n3288# 0.013296f
C274 source.n190 a_n1878_n3288# 0.012557f
C275 source.n191 a_n1878_n3288# 0.023369f
C276 source.n192 a_n1878_n3288# 0.023369f
C277 source.n193 a_n1878_n3288# 0.012557f
C278 source.n194 a_n1878_n3288# 0.013296f
C279 source.n195 a_n1878_n3288# 0.029681f
C280 source.n196 a_n1878_n3288# 0.060908f
C281 source.n197 a_n1878_n3288# 0.013296f
C282 source.n198 a_n1878_n3288# 0.012557f
C283 source.n199 a_n1878_n3288# 0.050185f
C284 source.n200 a_n1878_n3288# 0.033615f
C285 source.n201 a_n1878_n3288# 0.107056f
C286 source.t22 a_n1878_n3288# 0.2216f
C287 source.t4 a_n1878_n3288# 0.2216f
C288 source.n202 a_n1878_n3288# 1.89734f
C289 source.n203 a_n1878_n3288# 0.346671f
C290 source.t5 a_n1878_n3288# 0.2216f
C291 source.t21 a_n1878_n3288# 0.2216f
C292 source.n204 a_n1878_n3288# 1.89734f
C293 source.n205 a_n1878_n3288# 0.346671f
C294 source.n206 a_n1878_n3288# 0.030955f
C295 source.n207 a_n1878_n3288# 0.023369f
C296 source.n208 a_n1878_n3288# 0.012557f
C297 source.n209 a_n1878_n3288# 0.029681f
C298 source.n210 a_n1878_n3288# 0.013296f
C299 source.n211 a_n1878_n3288# 0.023369f
C300 source.n212 a_n1878_n3288# 0.012557f
C301 source.n213 a_n1878_n3288# 0.029681f
C302 source.n214 a_n1878_n3288# 0.013296f
C303 source.n215 a_n1878_n3288# 0.023369f
C304 source.n216 a_n1878_n3288# 0.012927f
C305 source.n217 a_n1878_n3288# 0.029681f
C306 source.n218 a_n1878_n3288# 0.012557f
C307 source.n219 a_n1878_n3288# 0.013296f
C308 source.n220 a_n1878_n3288# 0.023369f
C309 source.n221 a_n1878_n3288# 0.012557f
C310 source.n222 a_n1878_n3288# 0.029681f
C311 source.n223 a_n1878_n3288# 0.013296f
C312 source.n224 a_n1878_n3288# 0.023369f
C313 source.n225 a_n1878_n3288# 0.012557f
C314 source.n226 a_n1878_n3288# 0.022261f
C315 source.n227 a_n1878_n3288# 0.020982f
C316 source.t3 a_n1878_n3288# 0.050129f
C317 source.n228 a_n1878_n3288# 0.168486f
C318 source.n229 a_n1878_n3288# 1.17891f
C319 source.n230 a_n1878_n3288# 0.012557f
C320 source.n231 a_n1878_n3288# 0.013296f
C321 source.n232 a_n1878_n3288# 0.029681f
C322 source.n233 a_n1878_n3288# 0.029681f
C323 source.n234 a_n1878_n3288# 0.013296f
C324 source.n235 a_n1878_n3288# 0.012557f
C325 source.n236 a_n1878_n3288# 0.023369f
C326 source.n237 a_n1878_n3288# 0.023369f
C327 source.n238 a_n1878_n3288# 0.012557f
C328 source.n239 a_n1878_n3288# 0.013296f
C329 source.n240 a_n1878_n3288# 0.029681f
C330 source.n241 a_n1878_n3288# 0.029681f
C331 source.n242 a_n1878_n3288# 0.013296f
C332 source.n243 a_n1878_n3288# 0.012557f
C333 source.n244 a_n1878_n3288# 0.023369f
C334 source.n245 a_n1878_n3288# 0.023369f
C335 source.n246 a_n1878_n3288# 0.012557f
C336 source.n247 a_n1878_n3288# 0.013296f
C337 source.n248 a_n1878_n3288# 0.029681f
C338 source.n249 a_n1878_n3288# 0.029681f
C339 source.n250 a_n1878_n3288# 0.029681f
C340 source.n251 a_n1878_n3288# 0.012927f
C341 source.n252 a_n1878_n3288# 0.012557f
C342 source.n253 a_n1878_n3288# 0.023369f
C343 source.n254 a_n1878_n3288# 0.023369f
C344 source.n255 a_n1878_n3288# 0.012557f
C345 source.n256 a_n1878_n3288# 0.013296f
C346 source.n257 a_n1878_n3288# 0.029681f
C347 source.n258 a_n1878_n3288# 0.029681f
C348 source.n259 a_n1878_n3288# 0.013296f
C349 source.n260 a_n1878_n3288# 0.012557f
C350 source.n261 a_n1878_n3288# 0.023369f
C351 source.n262 a_n1878_n3288# 0.023369f
C352 source.n263 a_n1878_n3288# 0.012557f
C353 source.n264 a_n1878_n3288# 0.013296f
C354 source.n265 a_n1878_n3288# 0.029681f
C355 source.n266 a_n1878_n3288# 0.060908f
C356 source.n267 a_n1878_n3288# 0.013296f
C357 source.n268 a_n1878_n3288# 0.012557f
C358 source.n269 a_n1878_n3288# 0.050185f
C359 source.n270 a_n1878_n3288# 0.033615f
C360 source.n271 a_n1878_n3288# 1.33389f
C361 source.n272 a_n1878_n3288# 0.030955f
C362 source.n273 a_n1878_n3288# 0.023369f
C363 source.n274 a_n1878_n3288# 0.012557f
C364 source.n275 a_n1878_n3288# 0.029681f
C365 source.n276 a_n1878_n3288# 0.013296f
C366 source.n277 a_n1878_n3288# 0.023369f
C367 source.n278 a_n1878_n3288# 0.012557f
C368 source.n279 a_n1878_n3288# 0.029681f
C369 source.n280 a_n1878_n3288# 0.013296f
C370 source.n281 a_n1878_n3288# 0.023369f
C371 source.n282 a_n1878_n3288# 0.012927f
C372 source.n283 a_n1878_n3288# 0.029681f
C373 source.n284 a_n1878_n3288# 0.013296f
C374 source.n285 a_n1878_n3288# 0.023369f
C375 source.n286 a_n1878_n3288# 0.012557f
C376 source.n287 a_n1878_n3288# 0.029681f
C377 source.n288 a_n1878_n3288# 0.013296f
C378 source.n289 a_n1878_n3288# 0.023369f
C379 source.n290 a_n1878_n3288# 0.012557f
C380 source.n291 a_n1878_n3288# 0.022261f
C381 source.n292 a_n1878_n3288# 0.020982f
C382 source.t14 a_n1878_n3288# 0.050129f
C383 source.n293 a_n1878_n3288# 0.168486f
C384 source.n294 a_n1878_n3288# 1.17891f
C385 source.n295 a_n1878_n3288# 0.012557f
C386 source.n296 a_n1878_n3288# 0.013296f
C387 source.n297 a_n1878_n3288# 0.029681f
C388 source.n298 a_n1878_n3288# 0.029681f
C389 source.n299 a_n1878_n3288# 0.013296f
C390 source.n300 a_n1878_n3288# 0.012557f
C391 source.n301 a_n1878_n3288# 0.023369f
C392 source.n302 a_n1878_n3288# 0.023369f
C393 source.n303 a_n1878_n3288# 0.012557f
C394 source.n304 a_n1878_n3288# 0.013296f
C395 source.n305 a_n1878_n3288# 0.029681f
C396 source.n306 a_n1878_n3288# 0.029681f
C397 source.n307 a_n1878_n3288# 0.013296f
C398 source.n308 a_n1878_n3288# 0.012557f
C399 source.n309 a_n1878_n3288# 0.023369f
C400 source.n310 a_n1878_n3288# 0.023369f
C401 source.n311 a_n1878_n3288# 0.012557f
C402 source.n312 a_n1878_n3288# 0.012557f
C403 source.n313 a_n1878_n3288# 0.013296f
C404 source.n314 a_n1878_n3288# 0.029681f
C405 source.n315 a_n1878_n3288# 0.029681f
C406 source.n316 a_n1878_n3288# 0.029681f
C407 source.n317 a_n1878_n3288# 0.012927f
C408 source.n318 a_n1878_n3288# 0.012557f
C409 source.n319 a_n1878_n3288# 0.023369f
C410 source.n320 a_n1878_n3288# 0.023369f
C411 source.n321 a_n1878_n3288# 0.012557f
C412 source.n322 a_n1878_n3288# 0.013296f
C413 source.n323 a_n1878_n3288# 0.029681f
C414 source.n324 a_n1878_n3288# 0.029681f
C415 source.n325 a_n1878_n3288# 0.013296f
C416 source.n326 a_n1878_n3288# 0.012557f
C417 source.n327 a_n1878_n3288# 0.023369f
C418 source.n328 a_n1878_n3288# 0.023369f
C419 source.n329 a_n1878_n3288# 0.012557f
C420 source.n330 a_n1878_n3288# 0.013296f
C421 source.n331 a_n1878_n3288# 0.029681f
C422 source.n332 a_n1878_n3288# 0.060908f
C423 source.n333 a_n1878_n3288# 0.013296f
C424 source.n334 a_n1878_n3288# 0.012557f
C425 source.n335 a_n1878_n3288# 0.050185f
C426 source.n336 a_n1878_n3288# 0.033615f
C427 source.n337 a_n1878_n3288# 1.33389f
C428 source.t18 a_n1878_n3288# 0.2216f
C429 source.t19 a_n1878_n3288# 0.2216f
C430 source.n338 a_n1878_n3288# 1.89733f
C431 source.n339 a_n1878_n3288# 0.346682f
C432 source.t16 a_n1878_n3288# 0.2216f
C433 source.t10 a_n1878_n3288# 0.2216f
C434 source.n340 a_n1878_n3288# 1.89733f
C435 source.n341 a_n1878_n3288# 0.346682f
C436 source.n342 a_n1878_n3288# 0.030955f
C437 source.n343 a_n1878_n3288# 0.023369f
C438 source.n344 a_n1878_n3288# 0.012557f
C439 source.n345 a_n1878_n3288# 0.029681f
C440 source.n346 a_n1878_n3288# 0.013296f
C441 source.n347 a_n1878_n3288# 0.023369f
C442 source.n348 a_n1878_n3288# 0.012557f
C443 source.n349 a_n1878_n3288# 0.029681f
C444 source.n350 a_n1878_n3288# 0.013296f
C445 source.n351 a_n1878_n3288# 0.023369f
C446 source.n352 a_n1878_n3288# 0.012927f
C447 source.n353 a_n1878_n3288# 0.029681f
C448 source.n354 a_n1878_n3288# 0.013296f
C449 source.n355 a_n1878_n3288# 0.023369f
C450 source.n356 a_n1878_n3288# 0.012557f
C451 source.n357 a_n1878_n3288# 0.029681f
C452 source.n358 a_n1878_n3288# 0.013296f
C453 source.n359 a_n1878_n3288# 0.023369f
C454 source.n360 a_n1878_n3288# 0.012557f
C455 source.n361 a_n1878_n3288# 0.022261f
C456 source.n362 a_n1878_n3288# 0.020982f
C457 source.t11 a_n1878_n3288# 0.050129f
C458 source.n363 a_n1878_n3288# 0.168486f
C459 source.n364 a_n1878_n3288# 1.17891f
C460 source.n365 a_n1878_n3288# 0.012557f
C461 source.n366 a_n1878_n3288# 0.013296f
C462 source.n367 a_n1878_n3288# 0.029681f
C463 source.n368 a_n1878_n3288# 0.029681f
C464 source.n369 a_n1878_n3288# 0.013296f
C465 source.n370 a_n1878_n3288# 0.012557f
C466 source.n371 a_n1878_n3288# 0.023369f
C467 source.n372 a_n1878_n3288# 0.023369f
C468 source.n373 a_n1878_n3288# 0.012557f
C469 source.n374 a_n1878_n3288# 0.013296f
C470 source.n375 a_n1878_n3288# 0.029681f
C471 source.n376 a_n1878_n3288# 0.029681f
C472 source.n377 a_n1878_n3288# 0.013296f
C473 source.n378 a_n1878_n3288# 0.012557f
C474 source.n379 a_n1878_n3288# 0.023369f
C475 source.n380 a_n1878_n3288# 0.023369f
C476 source.n381 a_n1878_n3288# 0.012557f
C477 source.n382 a_n1878_n3288# 0.012557f
C478 source.n383 a_n1878_n3288# 0.013296f
C479 source.n384 a_n1878_n3288# 0.029681f
C480 source.n385 a_n1878_n3288# 0.029681f
C481 source.n386 a_n1878_n3288# 0.029681f
C482 source.n387 a_n1878_n3288# 0.012927f
C483 source.n388 a_n1878_n3288# 0.012557f
C484 source.n389 a_n1878_n3288# 0.023369f
C485 source.n390 a_n1878_n3288# 0.023369f
C486 source.n391 a_n1878_n3288# 0.012557f
C487 source.n392 a_n1878_n3288# 0.013296f
C488 source.n393 a_n1878_n3288# 0.029681f
C489 source.n394 a_n1878_n3288# 0.029681f
C490 source.n395 a_n1878_n3288# 0.013296f
C491 source.n396 a_n1878_n3288# 0.012557f
C492 source.n397 a_n1878_n3288# 0.023369f
C493 source.n398 a_n1878_n3288# 0.023369f
C494 source.n399 a_n1878_n3288# 0.012557f
C495 source.n400 a_n1878_n3288# 0.013296f
C496 source.n401 a_n1878_n3288# 0.029681f
C497 source.n402 a_n1878_n3288# 0.060908f
C498 source.n403 a_n1878_n3288# 0.013296f
C499 source.n404 a_n1878_n3288# 0.012557f
C500 source.n405 a_n1878_n3288# 0.050185f
C501 source.n406 a_n1878_n3288# 0.033615f
C502 source.n407 a_n1878_n3288# 0.107056f
C503 source.n408 a_n1878_n3288# 0.030955f
C504 source.n409 a_n1878_n3288# 0.023369f
C505 source.n410 a_n1878_n3288# 0.012557f
C506 source.n411 a_n1878_n3288# 0.029681f
C507 source.n412 a_n1878_n3288# 0.013296f
C508 source.n413 a_n1878_n3288# 0.023369f
C509 source.n414 a_n1878_n3288# 0.012557f
C510 source.n415 a_n1878_n3288# 0.029681f
C511 source.n416 a_n1878_n3288# 0.013296f
C512 source.n417 a_n1878_n3288# 0.023369f
C513 source.n418 a_n1878_n3288# 0.012927f
C514 source.n419 a_n1878_n3288# 0.029681f
C515 source.n420 a_n1878_n3288# 0.013296f
C516 source.n421 a_n1878_n3288# 0.023369f
C517 source.n422 a_n1878_n3288# 0.012557f
C518 source.n423 a_n1878_n3288# 0.029681f
C519 source.n424 a_n1878_n3288# 0.013296f
C520 source.n425 a_n1878_n3288# 0.023369f
C521 source.n426 a_n1878_n3288# 0.012557f
C522 source.n427 a_n1878_n3288# 0.022261f
C523 source.n428 a_n1878_n3288# 0.020982f
C524 source.t1 a_n1878_n3288# 0.050129f
C525 source.n429 a_n1878_n3288# 0.168486f
C526 source.n430 a_n1878_n3288# 1.17891f
C527 source.n431 a_n1878_n3288# 0.012557f
C528 source.n432 a_n1878_n3288# 0.013296f
C529 source.n433 a_n1878_n3288# 0.029681f
C530 source.n434 a_n1878_n3288# 0.029681f
C531 source.n435 a_n1878_n3288# 0.013296f
C532 source.n436 a_n1878_n3288# 0.012557f
C533 source.n437 a_n1878_n3288# 0.023369f
C534 source.n438 a_n1878_n3288# 0.023369f
C535 source.n439 a_n1878_n3288# 0.012557f
C536 source.n440 a_n1878_n3288# 0.013296f
C537 source.n441 a_n1878_n3288# 0.029681f
C538 source.n442 a_n1878_n3288# 0.029681f
C539 source.n443 a_n1878_n3288# 0.013296f
C540 source.n444 a_n1878_n3288# 0.012557f
C541 source.n445 a_n1878_n3288# 0.023369f
C542 source.n446 a_n1878_n3288# 0.023369f
C543 source.n447 a_n1878_n3288# 0.012557f
C544 source.n448 a_n1878_n3288# 0.012557f
C545 source.n449 a_n1878_n3288# 0.013296f
C546 source.n450 a_n1878_n3288# 0.029681f
C547 source.n451 a_n1878_n3288# 0.029681f
C548 source.n452 a_n1878_n3288# 0.029681f
C549 source.n453 a_n1878_n3288# 0.012927f
C550 source.n454 a_n1878_n3288# 0.012557f
C551 source.n455 a_n1878_n3288# 0.023369f
C552 source.n456 a_n1878_n3288# 0.023369f
C553 source.n457 a_n1878_n3288# 0.012557f
C554 source.n458 a_n1878_n3288# 0.013296f
C555 source.n459 a_n1878_n3288# 0.029681f
C556 source.n460 a_n1878_n3288# 0.029681f
C557 source.n461 a_n1878_n3288# 0.013296f
C558 source.n462 a_n1878_n3288# 0.012557f
C559 source.n463 a_n1878_n3288# 0.023369f
C560 source.n464 a_n1878_n3288# 0.023369f
C561 source.n465 a_n1878_n3288# 0.012557f
C562 source.n466 a_n1878_n3288# 0.013296f
C563 source.n467 a_n1878_n3288# 0.029681f
C564 source.n468 a_n1878_n3288# 0.060908f
C565 source.n469 a_n1878_n3288# 0.013296f
C566 source.n470 a_n1878_n3288# 0.012557f
C567 source.n471 a_n1878_n3288# 0.050185f
C568 source.n472 a_n1878_n3288# 0.033615f
C569 source.n473 a_n1878_n3288# 0.107056f
C570 source.t7 a_n1878_n3288# 0.2216f
C571 source.t23 a_n1878_n3288# 0.2216f
C572 source.n474 a_n1878_n3288# 1.89733f
C573 source.n475 a_n1878_n3288# 0.346682f
C574 source.t0 a_n1878_n3288# 0.2216f
C575 source.t6 a_n1878_n3288# 0.2216f
C576 source.n476 a_n1878_n3288# 1.89733f
C577 source.n477 a_n1878_n3288# 0.346682f
C578 source.n478 a_n1878_n3288# 0.030955f
C579 source.n479 a_n1878_n3288# 0.023369f
C580 source.n480 a_n1878_n3288# 0.012557f
C581 source.n481 a_n1878_n3288# 0.029681f
C582 source.n482 a_n1878_n3288# 0.013296f
C583 source.n483 a_n1878_n3288# 0.023369f
C584 source.n484 a_n1878_n3288# 0.012557f
C585 source.n485 a_n1878_n3288# 0.029681f
C586 source.n486 a_n1878_n3288# 0.013296f
C587 source.n487 a_n1878_n3288# 0.023369f
C588 source.n488 a_n1878_n3288# 0.012927f
C589 source.n489 a_n1878_n3288# 0.029681f
C590 source.n490 a_n1878_n3288# 0.013296f
C591 source.n491 a_n1878_n3288# 0.023369f
C592 source.n492 a_n1878_n3288# 0.012557f
C593 source.n493 a_n1878_n3288# 0.029681f
C594 source.n494 a_n1878_n3288# 0.013296f
C595 source.n495 a_n1878_n3288# 0.023369f
C596 source.n496 a_n1878_n3288# 0.012557f
C597 source.n497 a_n1878_n3288# 0.022261f
C598 source.n498 a_n1878_n3288# 0.020982f
C599 source.t2 a_n1878_n3288# 0.050129f
C600 source.n499 a_n1878_n3288# 0.168486f
C601 source.n500 a_n1878_n3288# 1.17891f
C602 source.n501 a_n1878_n3288# 0.012557f
C603 source.n502 a_n1878_n3288# 0.013296f
C604 source.n503 a_n1878_n3288# 0.029681f
C605 source.n504 a_n1878_n3288# 0.029681f
C606 source.n505 a_n1878_n3288# 0.013296f
C607 source.n506 a_n1878_n3288# 0.012557f
C608 source.n507 a_n1878_n3288# 0.023369f
C609 source.n508 a_n1878_n3288# 0.023369f
C610 source.n509 a_n1878_n3288# 0.012557f
C611 source.n510 a_n1878_n3288# 0.013296f
C612 source.n511 a_n1878_n3288# 0.029681f
C613 source.n512 a_n1878_n3288# 0.029681f
C614 source.n513 a_n1878_n3288# 0.013296f
C615 source.n514 a_n1878_n3288# 0.012557f
C616 source.n515 a_n1878_n3288# 0.023369f
C617 source.n516 a_n1878_n3288# 0.023369f
C618 source.n517 a_n1878_n3288# 0.012557f
C619 source.n518 a_n1878_n3288# 0.012557f
C620 source.n519 a_n1878_n3288# 0.013296f
C621 source.n520 a_n1878_n3288# 0.029681f
C622 source.n521 a_n1878_n3288# 0.029681f
C623 source.n522 a_n1878_n3288# 0.029681f
C624 source.n523 a_n1878_n3288# 0.012927f
C625 source.n524 a_n1878_n3288# 0.012557f
C626 source.n525 a_n1878_n3288# 0.023369f
C627 source.n526 a_n1878_n3288# 0.023369f
C628 source.n527 a_n1878_n3288# 0.012557f
C629 source.n528 a_n1878_n3288# 0.013296f
C630 source.n529 a_n1878_n3288# 0.029681f
C631 source.n530 a_n1878_n3288# 0.029681f
C632 source.n531 a_n1878_n3288# 0.013296f
C633 source.n532 a_n1878_n3288# 0.012557f
C634 source.n533 a_n1878_n3288# 0.023369f
C635 source.n534 a_n1878_n3288# 0.023369f
C636 source.n535 a_n1878_n3288# 0.012557f
C637 source.n536 a_n1878_n3288# 0.013296f
C638 source.n537 a_n1878_n3288# 0.029681f
C639 source.n538 a_n1878_n3288# 0.060908f
C640 source.n539 a_n1878_n3288# 0.013296f
C641 source.n540 a_n1878_n3288# 0.012557f
C642 source.n541 a_n1878_n3288# 0.050185f
C643 source.n542 a_n1878_n3288# 0.033615f
C644 source.n543 a_n1878_n3288# 0.249289f
C645 source.n544 a_n1878_n3288# 1.47335f
C646 drain_left.t2 a_n1878_n3288# 0.277518f
C647 drain_left.t6 a_n1878_n3288# 0.277518f
C648 drain_left.n0 a_n1878_n3288# 2.47374f
C649 drain_left.t7 a_n1878_n3288# 0.277518f
C650 drain_left.t1 a_n1878_n3288# 0.277518f
C651 drain_left.n1 a_n1878_n3288# 2.46948f
C652 drain_left.t11 a_n1878_n3288# 0.277518f
C653 drain_left.t5 a_n1878_n3288# 0.277518f
C654 drain_left.n2 a_n1878_n3288# 2.47374f
C655 drain_left.n3 a_n1878_n3288# 2.5403f
C656 drain_left.t4 a_n1878_n3288# 0.277518f
C657 drain_left.t3 a_n1878_n3288# 0.277518f
C658 drain_left.n4 a_n1878_n3288# 2.47415f
C659 drain_left.t10 a_n1878_n3288# 0.277518f
C660 drain_left.t0 a_n1878_n3288# 0.277518f
C661 drain_left.n5 a_n1878_n3288# 2.46949f
C662 drain_left.n6 a_n1878_n3288# 0.768227f
C663 drain_left.t8 a_n1878_n3288# 0.277518f
C664 drain_left.t9 a_n1878_n3288# 0.277518f
C665 drain_left.n7 a_n1878_n3288# 2.46948f
C666 drain_left.n8 a_n1878_n3288# 0.631991f
C667 plus.n0 a_n1878_n3288# 0.047453f
C668 plus.t11 a_n1878_n3288# 0.811883f
C669 plus.t7 a_n1878_n3288# 0.811883f
C670 plus.n1 a_n1878_n3288# 0.047453f
C671 plus.t4 a_n1878_n3288# 0.811883f
C672 plus.n2 a_n1878_n3288# 0.047453f
C673 plus.t10 a_n1878_n3288# 0.811883f
C674 plus.n3 a_n1878_n3288# 0.332325f
C675 plus.t6 a_n1878_n3288# 0.811883f
C676 plus.n4 a_n1878_n3288# 0.338045f
C677 plus.t2 a_n1878_n3288# 0.824661f
C678 plus.n5 a_n1878_n3288# 0.315883f
C679 plus.n6 a_n1878_n3288# 0.19326f
C680 plus.n7 a_n1878_n3288# 0.047453f
C681 plus.n8 a_n1878_n3288# 0.010768f
C682 plus.n9 a_n1878_n3288# 0.332325f
C683 plus.n10 a_n1878_n3288# 0.327644f
C684 plus.n11 a_n1878_n3288# 0.010768f
C685 plus.n12 a_n1878_n3288# 0.327351f
C686 plus.n13 a_n1878_n3288# 0.534423f
C687 plus.n14 a_n1878_n3288# 0.047453f
C688 plus.t5 a_n1878_n3288# 0.811883f
C689 plus.n15 a_n1878_n3288# 0.047453f
C690 plus.t1 a_n1878_n3288# 0.811883f
C691 plus.n16 a_n1878_n3288# 0.047453f
C692 plus.t0 a_n1878_n3288# 0.811883f
C693 plus.t3 a_n1878_n3288# 0.811883f
C694 plus.n17 a_n1878_n3288# 0.332325f
C695 plus.t8 a_n1878_n3288# 0.824661f
C696 plus.t9 a_n1878_n3288# 0.811883f
C697 plus.n18 a_n1878_n3288# 0.338045f
C698 plus.n19 a_n1878_n3288# 0.315883f
C699 plus.n20 a_n1878_n3288# 0.19326f
C700 plus.n21 a_n1878_n3288# 0.047453f
C701 plus.n22 a_n1878_n3288# 0.010768f
C702 plus.n23 a_n1878_n3288# 0.332325f
C703 plus.n24 a_n1878_n3288# 0.327644f
C704 plus.n25 a_n1878_n3288# 0.010768f
C705 plus.n26 a_n1878_n3288# 0.327351f
C706 plus.n27 a_n1878_n3288# 1.4243f
.ends

