* NGSPICE file created from diffpair616.ext - technology: sky130A

.subckt diffpair616 minus drain_right drain_left source plus
X0 source.t24 minus.t0 drain_right.t8 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X1 drain_left.t13 plus.t0 source.t5 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X2 source.t1 plus.t1 drain_left.t12 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X3 drain_left.t11 plus.t2 source.t8 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X4 source.t10 plus.t3 drain_left.t10 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X5 source.t23 minus.t1 drain_right.t7 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X6 drain_right.t6 minus.t2 source.t22 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X7 drain_right.t3 minus.t3 source.t21 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X8 drain_left.t9 plus.t4 source.t9 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X9 source.t20 minus.t4 drain_right.t5 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X10 drain_right.t4 minus.t5 source.t19 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X11 source.t18 minus.t6 drain_right.t13 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X12 source.t2 plus.t5 drain_left.t8 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X13 drain_left.t7 plus.t6 source.t6 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X14 source.t17 minus.t7 drain_right.t2 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X15 drain_right.t1 minus.t8 source.t16 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X16 drain_right.t0 minus.t9 source.t15 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X17 source.t7 plus.t7 drain_left.t6 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X18 source.t0 plus.t8 drain_left.t5 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X19 source.t14 minus.t10 drain_right.t12 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X20 a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X21 drain_left.t4 plus.t9 source.t3 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X22 drain_right.t10 minus.t11 source.t13 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X23 drain_right.t9 minus.t12 source.t12 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X24 source.t25 plus.t10 drain_left.t3 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X25 drain_left.t2 plus.t11 source.t26 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X26 a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X27 drain_right.t11 minus.t13 source.t11 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X28 drain_left.t1 plus.t12 source.t27 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X29 drain_left.t0 plus.t13 source.t4 a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X30 a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X31 a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# a_n2204_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
R0 minus.n5 minus.t11 892.652
R1 minus.n23 minus.t13 892.652
R2 minus.n4 minus.t10 868.806
R3 minus.n8 minus.t9 868.806
R4 minus.n9 minus.t7 868.806
R5 minus.n10 minus.t2 868.806
R6 minus.n14 minus.t4 868.806
R7 minus.n16 minus.t3 868.806
R8 minus.n22 minus.t6 868.806
R9 minus.n26 minus.t8 868.806
R10 minus.n27 minus.t0 868.806
R11 minus.n28 minus.t5 868.806
R12 minus.n32 minus.t1 868.806
R13 minus.n34 minus.t12 868.806
R14 minus.n17 minus.n16 161.3
R15 minus.n15 minus.n0 161.3
R16 minus.n14 minus.n13 161.3
R17 minus.n12 minus.n1 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n6 minus.n3 161.3
R21 minus.n35 minus.n34 161.3
R22 minus.n33 minus.n18 161.3
R23 minus.n32 minus.n31 161.3
R24 minus.n30 minus.n19 161.3
R25 minus.n29 minus.n28 161.3
R26 minus.n26 minus.n25 161.3
R27 minus.n24 minus.n21 161.3
R28 minus.n9 minus.n2 80.6037
R29 minus.n27 minus.n20 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n4 minus.n3 45.2793
R35 minus.n14 minus.n1 45.2793
R36 minus.n22 minus.n21 45.2793
R37 minus.n32 minus.n19 45.2793
R38 minus.n6 minus.n5 44.9119
R39 minus.n24 minus.n23 44.9119
R40 minus.n36 minus.n17 43.6047
R41 minus.n16 minus.n15 35.055
R42 minus.n34 minus.n33 35.055
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n15 minus.n14 13.146
R46 minus.n33 minus.n32 13.146
R47 minus.n36 minus.n35 6.57436
R48 minus.n8 minus.n3 2.92171
R49 minus.n10 minus.n1 2.92171
R50 minus.n26 minus.n21 2.92171
R51 minus.n28 minus.n19 2.92171
R52 minus.n11 minus.n2 0.285035
R53 minus.n7 minus.n2 0.285035
R54 minus.n25 minus.n20 0.285035
R55 minus.n29 minus.n20 0.285035
R56 minus.n17 minus.n0 0.189894
R57 minus.n13 minus.n0 0.189894
R58 minus.n13 minus.n12 0.189894
R59 minus.n12 minus.n11 0.189894
R60 minus.n7 minus.n6 0.189894
R61 minus.n25 minus.n24 0.189894
R62 minus.n30 minus.n29 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 drain_right.n1 drain_right.t11 61.61
R68 drain_right.n11 drain_right.t3 60.8084
R69 drain_right.n8 drain_right.n6 60.6202
R70 drain_right.n4 drain_right.n2 60.6201
R71 drain_right.n8 drain_right.n7 59.8185
R72 drain_right.n10 drain_right.n9 59.8185
R73 drain_right.n4 drain_right.n3 59.8184
R74 drain_right.n1 drain_right.n0 59.8184
R75 drain_right drain_right.n5 37.4844
R76 drain_right drain_right.n11 6.05408
R77 drain_right.n2 drain_right.t7 0.9905
R78 drain_right.n2 drain_right.t9 0.9905
R79 drain_right.n3 drain_right.t8 0.9905
R80 drain_right.n3 drain_right.t4 0.9905
R81 drain_right.n0 drain_right.t13 0.9905
R82 drain_right.n0 drain_right.t1 0.9905
R83 drain_right.n6 drain_right.t12 0.9905
R84 drain_right.n6 drain_right.t10 0.9905
R85 drain_right.n7 drain_right.t2 0.9905
R86 drain_right.n7 drain_right.t0 0.9905
R87 drain_right.n9 drain_right.t5 0.9905
R88 drain_right.n9 drain_right.t6 0.9905
R89 drain_right.n11 drain_right.n10 0.802224
R90 drain_right.n10 drain_right.n8 0.802224
R91 drain_right.n5 drain_right.n1 0.546447
R92 drain_right.n5 drain_right.n4 0.145585
R93 source.n0 source.t8 44.1297
R94 source.n7 source.t13 44.1296
R95 source.n27 source.t12 44.1295
R96 source.n20 source.t5 44.1295
R97 source.n2 source.n1 43.1397
R98 source.n4 source.n3 43.1397
R99 source.n6 source.n5 43.1397
R100 source.n9 source.n8 43.1397
R101 source.n11 source.n10 43.1397
R102 source.n13 source.n12 43.1397
R103 source.n26 source.n25 43.1396
R104 source.n24 source.n23 43.1396
R105 source.n22 source.n21 43.1396
R106 source.n19 source.n18 43.1396
R107 source.n17 source.n16 43.1396
R108 source.n15 source.n14 43.1396
R109 source.n15 source.n13 28.9518
R110 source.n28 source.n0 22.4863
R111 source.n28 source.n27 5.66429
R112 source.n25 source.t19 0.9905
R113 source.n25 source.t23 0.9905
R114 source.n23 source.t16 0.9905
R115 source.n23 source.t24 0.9905
R116 source.n21 source.t11 0.9905
R117 source.n21 source.t18 0.9905
R118 source.n18 source.t27 0.9905
R119 source.n18 source.t7 0.9905
R120 source.n16 source.t9 0.9905
R121 source.n16 source.t1 0.9905
R122 source.n14 source.t4 0.9905
R123 source.n14 source.t2 0.9905
R124 source.n1 source.t6 0.9905
R125 source.n1 source.t10 0.9905
R126 source.n3 source.t3 0.9905
R127 source.n3 source.t0 0.9905
R128 source.n5 source.t26 0.9905
R129 source.n5 source.t25 0.9905
R130 source.n8 source.t15 0.9905
R131 source.n8 source.t14 0.9905
R132 source.n10 source.t22 0.9905
R133 source.n10 source.t17 0.9905
R134 source.n12 source.t21 0.9905
R135 source.n12 source.t20 0.9905
R136 source.n7 source.n6 0.87119
R137 source.n22 source.n20 0.87119
R138 source.n13 source.n11 0.802224
R139 source.n11 source.n9 0.802224
R140 source.n9 source.n7 0.802224
R141 source.n6 source.n4 0.802224
R142 source.n4 source.n2 0.802224
R143 source.n2 source.n0 0.802224
R144 source.n17 source.n15 0.802224
R145 source.n19 source.n17 0.802224
R146 source.n20 source.n19 0.802224
R147 source.n24 source.n22 0.802224
R148 source.n26 source.n24 0.802224
R149 source.n27 source.n26 0.802224
R150 source source.n28 0.188
R151 plus.n5 plus.t11 892.652
R152 plus.n23 plus.t0 892.652
R153 plus.n16 plus.t2 868.806
R154 plus.n14 plus.t3 868.806
R155 plus.n2 plus.t6 868.806
R156 plus.n9 plus.t8 868.806
R157 plus.n8 plus.t9 868.806
R158 plus.n4 plus.t10 868.806
R159 plus.n34 plus.t13 868.806
R160 plus.n32 plus.t5 868.806
R161 plus.n20 plus.t4 868.806
R162 plus.n27 plus.t1 868.806
R163 plus.n26 plus.t12 868.806
R164 plus.n22 plus.t7 868.806
R165 plus.n7 plus.n6 161.3
R166 plus.n8 plus.n3 161.3
R167 plus.n11 plus.n2 161.3
R168 plus.n13 plus.n12 161.3
R169 plus.n14 plus.n1 161.3
R170 plus.n15 plus.n0 161.3
R171 plus.n17 plus.n16 161.3
R172 plus.n25 plus.n24 161.3
R173 plus.n26 plus.n21 161.3
R174 plus.n29 plus.n20 161.3
R175 plus.n31 plus.n30 161.3
R176 plus.n32 plus.n19 161.3
R177 plus.n33 plus.n18 161.3
R178 plus.n35 plus.n34 161.3
R179 plus.n10 plus.n9 80.6037
R180 plus.n28 plus.n27 80.6037
R181 plus.n9 plus.n2 48.2005
R182 plus.n9 plus.n8 48.2005
R183 plus.n27 plus.n20 48.2005
R184 plus.n27 plus.n26 48.2005
R185 plus.n14 plus.n13 45.2793
R186 plus.n7 plus.n4 45.2793
R187 plus.n32 plus.n31 45.2793
R188 plus.n25 plus.n22 45.2793
R189 plus.n24 plus.n23 44.9119
R190 plus.n6 plus.n5 44.9119
R191 plus.n16 plus.n15 35.055
R192 plus.n34 plus.n33 35.055
R193 plus plus.n35 34.4555
R194 plus.n23 plus.n22 17.739
R195 plus.n5 plus.n4 17.739
R196 plus plus.n17 15.2486
R197 plus.n15 plus.n14 13.146
R198 plus.n33 plus.n32 13.146
R199 plus.n13 plus.n2 2.92171
R200 plus.n8 plus.n7 2.92171
R201 plus.n31 plus.n20 2.92171
R202 plus.n26 plus.n25 2.92171
R203 plus.n10 plus.n3 0.285035
R204 plus.n11 plus.n10 0.285035
R205 plus.n29 plus.n28 0.285035
R206 plus.n28 plus.n21 0.285035
R207 plus.n6 plus.n3 0.189894
R208 plus.n12 plus.n11 0.189894
R209 plus.n12 plus.n1 0.189894
R210 plus.n1 plus.n0 0.189894
R211 plus.n17 plus.n0 0.189894
R212 plus.n35 plus.n18 0.189894
R213 plus.n19 plus.n18 0.189894
R214 plus.n30 plus.n19 0.189894
R215 plus.n30 plus.n29 0.189894
R216 plus.n24 plus.n21 0.189894
R217 drain_left.n7 drain_left.t2 61.6101
R218 drain_left.n1 drain_left.t0 61.61
R219 drain_left.n4 drain_left.n2 60.6201
R220 drain_left.n11 drain_left.n10 59.8185
R221 drain_left.n9 drain_left.n8 59.8185
R222 drain_left.n7 drain_left.n6 59.8185
R223 drain_left.n4 drain_left.n3 59.8184
R224 drain_left.n1 drain_left.n0 59.8184
R225 drain_left drain_left.n5 38.0376
R226 drain_left drain_left.n11 6.45494
R227 drain_left.n2 drain_left.t6 0.9905
R228 drain_left.n2 drain_left.t13 0.9905
R229 drain_left.n3 drain_left.t12 0.9905
R230 drain_left.n3 drain_left.t1 0.9905
R231 drain_left.n0 drain_left.t8 0.9905
R232 drain_left.n0 drain_left.t9 0.9905
R233 drain_left.n10 drain_left.t10 0.9905
R234 drain_left.n10 drain_left.t11 0.9905
R235 drain_left.n8 drain_left.t5 0.9905
R236 drain_left.n8 drain_left.t7 0.9905
R237 drain_left.n6 drain_left.t3 0.9905
R238 drain_left.n6 drain_left.t4 0.9905
R239 drain_left.n9 drain_left.n7 0.802224
R240 drain_left.n11 drain_left.n9 0.802224
R241 drain_left.n5 drain_left.n1 0.546447
R242 drain_left.n5 drain_left.n4 0.145585
C0 plus minus 7.37972f
C1 source plus 13.083401f
C2 drain_left plus 13.6929f
C3 drain_right minus 13.480401f
C4 source drain_right 31.373999f
C5 drain_left drain_right 1.15099f
C6 source minus 13.068501f
C7 drain_left minus 0.172803f
C8 source drain_left 31.386702f
C9 drain_right plus 0.375748f
C10 drain_right a_n2204_n4888# 9.67959f
C11 drain_left a_n2204_n4888# 10.00932f
C12 source a_n2204_n4888# 9.449759f
C13 minus a_n2204_n4888# 9.258038f
C14 plus a_n2204_n4888# 11.46844f
C15 drain_left.t0 a_n2204_n4888# 4.76967f
C16 drain_left.t8 a_n2204_n4888# 0.407518f
C17 drain_left.t9 a_n2204_n4888# 0.407518f
C18 drain_left.n0 a_n2204_n4888# 3.72561f
C19 drain_left.n1 a_n2204_n4888# 0.692594f
C20 drain_left.t6 a_n2204_n4888# 0.407518f
C21 drain_left.t13 a_n2204_n4888# 0.407518f
C22 drain_left.n2 a_n2204_n4888# 3.73039f
C23 drain_left.t12 a_n2204_n4888# 0.407518f
C24 drain_left.t1 a_n2204_n4888# 0.407518f
C25 drain_left.n3 a_n2204_n4888# 3.72561f
C26 drain_left.n4 a_n2204_n4888# 0.656787f
C27 drain_left.n5 a_n2204_n4888# 1.88179f
C28 drain_left.t2 a_n2204_n4888# 4.76969f
C29 drain_left.t3 a_n2204_n4888# 0.407518f
C30 drain_left.t4 a_n2204_n4888# 0.407518f
C31 drain_left.n6 a_n2204_n4888# 3.72561f
C32 drain_left.n7 a_n2204_n4888# 0.712737f
C33 drain_left.t5 a_n2204_n4888# 0.407518f
C34 drain_left.t7 a_n2204_n4888# 0.407518f
C35 drain_left.n8 a_n2204_n4888# 3.72561f
C36 drain_left.n9 a_n2204_n4888# 0.350813f
C37 drain_left.t10 a_n2204_n4888# 0.407518f
C38 drain_left.t11 a_n2204_n4888# 0.407518f
C39 drain_left.n10 a_n2204_n4888# 3.72561f
C40 drain_left.n11 a_n2204_n4888# 0.575654f
C41 plus.n0 a_n2204_n4888# 0.043504f
C42 plus.t2 a_n2204_n4888# 1.47837f
C43 plus.t3 a_n2204_n4888# 1.47837f
C44 plus.n1 a_n2204_n4888# 0.043504f
C45 plus.t6 a_n2204_n4888# 1.47837f
C46 plus.n2 a_n2204_n4888# 0.553915f
C47 plus.n3 a_n2204_n4888# 0.05805f
C48 plus.t8 a_n2204_n4888# 1.47837f
C49 plus.t9 a_n2204_n4888# 1.47837f
C50 plus.t10 a_n2204_n4888# 1.47837f
C51 plus.n4 a_n2204_n4888# 0.560645f
C52 plus.t11 a_n2204_n4888# 1.49313f
C53 plus.n5 a_n2204_n4888# 0.54155f
C54 plus.n6 a_n2204_n4888# 0.177978f
C55 plus.n7 a_n2204_n4888# 0.009872f
C56 plus.n8 a_n2204_n4888# 0.553915f
C57 plus.n9 a_n2204_n4888# 0.563251f
C58 plus.n10 a_n2204_n4888# 0.057914f
C59 plus.n11 a_n2204_n4888# 0.05805f
C60 plus.n12 a_n2204_n4888# 0.043504f
C61 plus.n13 a_n2204_n4888# 0.009872f
C62 plus.n14 a_n2204_n4888# 0.555256f
C63 plus.n15 a_n2204_n4888# 0.009872f
C64 plus.n16 a_n2204_n4888# 0.550965f
C65 plus.n17 a_n2204_n4888# 0.668002f
C66 plus.n18 a_n2204_n4888# 0.043504f
C67 plus.t13 a_n2204_n4888# 1.47837f
C68 plus.n19 a_n2204_n4888# 0.043504f
C69 plus.t5 a_n2204_n4888# 1.47837f
C70 plus.t4 a_n2204_n4888# 1.47837f
C71 plus.n20 a_n2204_n4888# 0.553915f
C72 plus.n21 a_n2204_n4888# 0.05805f
C73 plus.t1 a_n2204_n4888# 1.47837f
C74 plus.t12 a_n2204_n4888# 1.47837f
C75 plus.t7 a_n2204_n4888# 1.47837f
C76 plus.n22 a_n2204_n4888# 0.560645f
C77 plus.t0 a_n2204_n4888# 1.49313f
C78 plus.n23 a_n2204_n4888# 0.54155f
C79 plus.n24 a_n2204_n4888# 0.177978f
C80 plus.n25 a_n2204_n4888# 0.009872f
C81 plus.n26 a_n2204_n4888# 0.553915f
C82 plus.n27 a_n2204_n4888# 0.563251f
C83 plus.n28 a_n2204_n4888# 0.057914f
C84 plus.n29 a_n2204_n4888# 0.05805f
C85 plus.n30 a_n2204_n4888# 0.043504f
C86 plus.n31 a_n2204_n4888# 0.009872f
C87 plus.n32 a_n2204_n4888# 0.555256f
C88 plus.n33 a_n2204_n4888# 0.009872f
C89 plus.n34 a_n2204_n4888# 0.550965f
C90 plus.n35 a_n2204_n4888# 1.62134f
C91 source.t8 a_n2204_n4888# 4.76175f
C92 source.n0 a_n2204_n4888# 2.05996f
C93 source.t6 a_n2204_n4888# 0.41666f
C94 source.t10 a_n2204_n4888# 0.41666f
C95 source.n1 a_n2204_n4888# 3.72512f
C96 source.n2 a_n2204_n4888# 0.406924f
C97 source.t3 a_n2204_n4888# 0.41666f
C98 source.t0 a_n2204_n4888# 0.41666f
C99 source.n3 a_n2204_n4888# 3.72512f
C100 source.n4 a_n2204_n4888# 0.406924f
C101 source.t26 a_n2204_n4888# 0.41666f
C102 source.t25 a_n2204_n4888# 0.41666f
C103 source.n5 a_n2204_n4888# 3.72512f
C104 source.n6 a_n2204_n4888# 0.412782f
C105 source.t13 a_n2204_n4888# 4.76176f
C106 source.n7 a_n2204_n4888# 0.512487f
C107 source.t15 a_n2204_n4888# 0.41666f
C108 source.t14 a_n2204_n4888# 0.41666f
C109 source.n8 a_n2204_n4888# 3.72512f
C110 source.n9 a_n2204_n4888# 0.406924f
C111 source.t22 a_n2204_n4888# 0.41666f
C112 source.t17 a_n2204_n4888# 0.41666f
C113 source.n10 a_n2204_n4888# 3.72512f
C114 source.n11 a_n2204_n4888# 0.406924f
C115 source.t21 a_n2204_n4888# 0.41666f
C116 source.t20 a_n2204_n4888# 0.41666f
C117 source.n12 a_n2204_n4888# 3.72512f
C118 source.n13 a_n2204_n4888# 2.50486f
C119 source.t4 a_n2204_n4888# 0.41666f
C120 source.t2 a_n2204_n4888# 0.41666f
C121 source.n14 a_n2204_n4888# 3.72513f
C122 source.n15 a_n2204_n4888# 2.50485f
C123 source.t9 a_n2204_n4888# 0.41666f
C124 source.t1 a_n2204_n4888# 0.41666f
C125 source.n16 a_n2204_n4888# 3.72513f
C126 source.n17 a_n2204_n4888# 0.406916f
C127 source.t27 a_n2204_n4888# 0.41666f
C128 source.t7 a_n2204_n4888# 0.41666f
C129 source.n18 a_n2204_n4888# 3.72513f
C130 source.n19 a_n2204_n4888# 0.406916f
C131 source.t5 a_n2204_n4888# 4.76173f
C132 source.n20 a_n2204_n4888# 0.512514f
C133 source.t11 a_n2204_n4888# 0.41666f
C134 source.t18 a_n2204_n4888# 0.41666f
C135 source.n21 a_n2204_n4888# 3.72513f
C136 source.n22 a_n2204_n4888# 0.412775f
C137 source.t16 a_n2204_n4888# 0.41666f
C138 source.t24 a_n2204_n4888# 0.41666f
C139 source.n23 a_n2204_n4888# 3.72513f
C140 source.n24 a_n2204_n4888# 0.406916f
C141 source.t19 a_n2204_n4888# 0.41666f
C142 source.t23 a_n2204_n4888# 0.41666f
C143 source.n25 a_n2204_n4888# 3.72513f
C144 source.n26 a_n2204_n4888# 0.406916f
C145 source.t12 a_n2204_n4888# 4.76173f
C146 source.n27 a_n2204_n4888# 0.644691f
C147 source.n28 a_n2204_n4888# 2.38706f
C148 drain_right.t11 a_n2204_n4888# 4.75916f
C149 drain_right.t13 a_n2204_n4888# 0.40662f
C150 drain_right.t1 a_n2204_n4888# 0.40662f
C151 drain_right.n0 a_n2204_n4888# 3.71741f
C152 drain_right.n1 a_n2204_n4888# 0.691068f
C153 drain_right.t7 a_n2204_n4888# 0.40662f
C154 drain_right.t9 a_n2204_n4888# 0.40662f
C155 drain_right.n2 a_n2204_n4888# 3.72217f
C156 drain_right.t8 a_n2204_n4888# 0.40662f
C157 drain_right.t4 a_n2204_n4888# 0.40662f
C158 drain_right.n3 a_n2204_n4888# 3.71741f
C159 drain_right.n4 a_n2204_n4888# 0.65534f
C160 drain_right.n5 a_n2204_n4888# 1.82437f
C161 drain_right.t12 a_n2204_n4888# 0.40662f
C162 drain_right.t10 a_n2204_n4888# 0.40662f
C163 drain_right.n6 a_n2204_n4888# 3.72217f
C164 drain_right.t2 a_n2204_n4888# 0.40662f
C165 drain_right.t0 a_n2204_n4888# 0.40662f
C166 drain_right.n7 a_n2204_n4888# 3.7174f
C167 drain_right.n8 a_n2204_n4888# 0.705676f
C168 drain_right.t5 a_n2204_n4888# 0.40662f
C169 drain_right.t6 a_n2204_n4888# 0.40662f
C170 drain_right.n9 a_n2204_n4888# 3.7174f
C171 drain_right.n10 a_n2204_n4888# 0.35004f
C172 drain_right.t3 a_n2204_n4888# 4.75442f
C173 drain_right.n11 a_n2204_n4888# 0.596927f
C174 minus.n0 a_n2204_n4888# 0.043138f
C175 minus.n1 a_n2204_n4888# 0.009789f
C176 minus.t4 a_n2204_n4888# 1.46595f
C177 minus.n2 a_n2204_n4888# 0.057428f
C178 minus.n3 a_n2204_n4888# 0.009789f
C179 minus.t9 a_n2204_n4888# 1.46595f
C180 minus.t11 a_n2204_n4888# 1.48059f
C181 minus.t10 a_n2204_n4888# 1.46595f
C182 minus.n4 a_n2204_n4888# 0.555936f
C183 minus.n5 a_n2204_n4888# 0.537001f
C184 minus.n6 a_n2204_n4888# 0.176483f
C185 minus.n7 a_n2204_n4888# 0.057562f
C186 minus.n8 a_n2204_n4888# 0.549263f
C187 minus.t7 a_n2204_n4888# 1.46595f
C188 minus.n9 a_n2204_n4888# 0.55852f
C189 minus.t2 a_n2204_n4888# 1.46595f
C190 minus.n10 a_n2204_n4888# 0.549263f
C191 minus.n11 a_n2204_n4888# 0.057562f
C192 minus.n12 a_n2204_n4888# 0.043138f
C193 minus.n13 a_n2204_n4888# 0.043138f
C194 minus.n14 a_n2204_n4888# 0.550593f
C195 minus.n15 a_n2204_n4888# 0.009789f
C196 minus.t3 a_n2204_n4888# 1.46595f
C197 minus.n16 a_n2204_n4888# 0.546337f
C198 minus.n17 a_n2204_n4888# 2.02016f
C199 minus.n18 a_n2204_n4888# 0.043138f
C200 minus.n19 a_n2204_n4888# 0.009789f
C201 minus.n20 a_n2204_n4888# 0.057428f
C202 minus.n21 a_n2204_n4888# 0.009789f
C203 minus.t13 a_n2204_n4888# 1.48059f
C204 minus.t6 a_n2204_n4888# 1.46595f
C205 minus.n22 a_n2204_n4888# 0.555936f
C206 minus.n23 a_n2204_n4888# 0.537001f
C207 minus.n24 a_n2204_n4888# 0.176483f
C208 minus.n25 a_n2204_n4888# 0.057562f
C209 minus.t8 a_n2204_n4888# 1.46595f
C210 minus.n26 a_n2204_n4888# 0.549263f
C211 minus.t0 a_n2204_n4888# 1.46595f
C212 minus.n27 a_n2204_n4888# 0.55852f
C213 minus.t5 a_n2204_n4888# 1.46595f
C214 minus.n28 a_n2204_n4888# 0.549263f
C215 minus.n29 a_n2204_n4888# 0.057562f
C216 minus.n30 a_n2204_n4888# 0.043138f
C217 minus.n31 a_n2204_n4888# 0.043138f
C218 minus.t1 a_n2204_n4888# 1.46595f
C219 minus.n32 a_n2204_n4888# 0.550593f
C220 minus.n33 a_n2204_n4888# 0.009789f
C221 minus.t12 a_n2204_n4888# 1.46595f
C222 minus.n34 a_n2204_n4888# 0.546337f
C223 minus.n35 a_n2204_n4888# 0.289557f
C224 minus.n36 a_n2204_n4888# 2.3999f
.ends

