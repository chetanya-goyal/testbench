* NGSPICE file created from diffpair518.ext - technology: sky130A

.subckt diffpair518 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t26 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X1 source.t15 minus.t0 drain_right.t19 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X2 drain_left.t18 plus.t1 source.t35 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X3 drain_left.t17 plus.t2 source.t24 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X4 drain_right.t18 minus.t1 source.t2 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X5 drain_right.t17 minus.t2 source.t8 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X6 source.t27 plus.t3 drain_left.t16 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X7 source.t1 minus.t3 drain_right.t16 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X8 source.t5 minus.t4 drain_right.t15 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X9 drain_right.t14 minus.t5 source.t3 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X10 drain_right.t13 minus.t6 source.t16 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X11 drain_left.t15 plus.t4 source.t22 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X12 source.t10 minus.t7 drain_right.t12 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X13 a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X14 drain_left.t14 plus.t5 source.t21 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X15 drain_left.t13 plus.t6 source.t29 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X16 source.t18 plus.t7 drain_left.t12 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 drain_left.t11 plus.t8 source.t37 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X18 source.t9 minus.t8 drain_right.t11 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X19 source.t38 minus.t9 drain_right.t10 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X20 source.t39 minus.t10 drain_right.t9 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X21 a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X22 source.t28 plus.t9 drain_left.t10 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X24 drain_right.t8 minus.t11 source.t4 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X25 drain_left.t9 plus.t10 source.t36 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X26 source.t34 plus.t11 drain_left.t8 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X27 source.t25 plus.t12 drain_left.t7 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X28 source.t23 plus.t13 drain_left.t6 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X29 source.t30 plus.t14 drain_left.t5 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X30 drain_left.t4 plus.t15 source.t19 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X31 drain_right.t7 minus.t12 source.t0 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X32 a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X33 drain_right.t6 minus.t13 source.t17 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X34 drain_right.t5 minus.t14 source.t12 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X35 source.t14 minus.t15 drain_right.t4 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X36 source.t7 minus.t16 drain_right.t3 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X37 source.t11 minus.t17 drain_right.t2 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X38 source.t20 plus.t16 drain_left.t3 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X39 drain_right.t1 minus.t18 source.t13 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X40 drain_right.t0 minus.t19 source.t6 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X41 source.t32 plus.t17 drain_left.t2 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X42 source.t31 plus.t18 drain_left.t1 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X43 drain_left.t0 plus.t19 source.t33 a_n2102_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 plus.n6 plus.t3 1358.36
R1 plus.n27 plus.t15 1358.36
R2 plus.n36 plus.t1 1358.36
R3 plus.n56 plus.t18 1358.36
R4 plus.n5 plus.t8 1309.43
R5 plus.n9 plus.t12 1309.43
R6 plus.n3 plus.t19 1309.43
R7 plus.n15 plus.t7 1309.43
R8 plus.n17 plus.t10 1309.43
R9 plus.n18 plus.t16 1309.43
R10 plus.n24 plus.t0 1309.43
R11 plus.n26 plus.t9 1309.43
R12 plus.n35 plus.t11 1309.43
R13 plus.n39 plus.t2 1309.43
R14 plus.n33 plus.t13 1309.43
R15 plus.n45 plus.t5 1309.43
R16 plus.n47 plus.t14 1309.43
R17 plus.n32 plus.t6 1309.43
R18 plus.n53 plus.t17 1309.43
R19 plus.n55 plus.t4 1309.43
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 64.9975
R47 plus.n19 plus.n18 64.9975
R48 plus.n48 plus.n32 64.9975
R49 plus.n44 plus.n33 64.9975
R50 plus.n9 plus.n8 62.0763
R51 plus.n25 plus.n24 62.0763
R52 plus.n54 plus.n53 62.0763
R53 plus.n39 plus.n38 62.0763
R54 plus.n16 plus.n15 46.0096
R55 plus.n17 plus.n16 46.0096
R56 plus.n47 plus.n46 46.0096
R57 plus.n46 plus.n45 46.0096
R58 plus.n6 plus.n5 43.0884
R59 plus.n27 plus.n26 43.0884
R60 plus.n56 plus.n55 43.0884
R61 plus.n36 plus.n35 43.0884
R62 plus plus.n57 32.1164
R63 plus.n8 plus.n5 29.9429
R64 plus.n26 plus.n25 29.9429
R65 plus.n55 plus.n54 29.9429
R66 plus.n38 plus.n35 29.9429
R67 plus.n15 plus.n14 27.0217
R68 plus.n19 plus.n17 27.0217
R69 plus.n48 plus.n47 27.0217
R70 plus.n45 plus.n44 27.0217
R71 plus plus.n28 13.296
R72 plus.n10 plus.n9 10.955
R73 plus.n24 plus.n23 10.955
R74 plus.n53 plus.n52 10.955
R75 plus.n40 plus.n39 10.955
R76 plus.n11 plus.n3 8.03383
R77 plus.n18 plus.n1 8.03383
R78 plus.n32 plus.n30 8.03383
R79 plus.n41 plus.n33 8.03383
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n9 source.t27 45.521
R99 source.n10 source.t4 45.521
R100 source.n19 source.t10 45.521
R101 source.n39 source.t3 45.5208
R102 source.n30 source.t5 45.5208
R103 source.n29 source.t35 45.5208
R104 source.n20 source.t31 45.5208
R105 source.n0 source.t19 45.5208
R106 source.n2 source.n1 44.201
R107 source.n4 source.n3 44.201
R108 source.n6 source.n5 44.201
R109 source.n8 source.n7 44.201
R110 source.n12 source.n11 44.201
R111 source.n14 source.n13 44.201
R112 source.n16 source.n15 44.201
R113 source.n18 source.n17 44.201
R114 source.n38 source.n37 44.2008
R115 source.n36 source.n35 44.2008
R116 source.n34 source.n33 44.2008
R117 source.n32 source.n31 44.2008
R118 source.n28 source.n27 44.2008
R119 source.n26 source.n25 44.2008
R120 source.n24 source.n23 44.2008
R121 source.n22 source.n21 44.2008
R122 source.n20 source.n19 24.1036
R123 source.n40 source.n0 18.5691
R124 source.n40 source.n39 5.53498
R125 source.n37 source.t13 1.3205
R126 source.n37 source.t11 1.3205
R127 source.n35 source.t6 1.3205
R128 source.n35 source.t38 1.3205
R129 source.n33 source.t17 1.3205
R130 source.n33 source.t39 1.3205
R131 source.n31 source.t12 1.3205
R132 source.n31 source.t1 1.3205
R133 source.n27 source.t24 1.3205
R134 source.n27 source.t34 1.3205
R135 source.n25 source.t21 1.3205
R136 source.n25 source.t23 1.3205
R137 source.n23 source.t29 1.3205
R138 source.n23 source.t30 1.3205
R139 source.n21 source.t22 1.3205
R140 source.n21 source.t32 1.3205
R141 source.n1 source.t26 1.3205
R142 source.n1 source.t28 1.3205
R143 source.n3 source.t36 1.3205
R144 source.n3 source.t20 1.3205
R145 source.n5 source.t33 1.3205
R146 source.n5 source.t18 1.3205
R147 source.n7 source.t37 1.3205
R148 source.n7 source.t25 1.3205
R149 source.n11 source.t2 1.3205
R150 source.n11 source.t14 1.3205
R151 source.n13 source.t0 1.3205
R152 source.n13 source.t9 1.3205
R153 source.n15 source.t16 1.3205
R154 source.n15 source.t15 1.3205
R155 source.n17 source.t8 1.3205
R156 source.n17 source.t7 1.3205
R157 source.n19 source.n18 0.543603
R158 source.n18 source.n16 0.543603
R159 source.n16 source.n14 0.543603
R160 source.n14 source.n12 0.543603
R161 source.n12 source.n10 0.543603
R162 source.n9 source.n8 0.543603
R163 source.n8 source.n6 0.543603
R164 source.n6 source.n4 0.543603
R165 source.n4 source.n2 0.543603
R166 source.n2 source.n0 0.543603
R167 source.n22 source.n20 0.543603
R168 source.n24 source.n22 0.543603
R169 source.n26 source.n24 0.543603
R170 source.n28 source.n26 0.543603
R171 source.n29 source.n28 0.543603
R172 source.n32 source.n30 0.543603
R173 source.n34 source.n32 0.543603
R174 source.n36 source.n34 0.543603
R175 source.n38 source.n36 0.543603
R176 source.n39 source.n38 0.543603
R177 source.n10 source.n9 0.470328
R178 source.n30 source.n29 0.470328
R179 source source.n40 0.188
R180 drain_left.n10 drain_left.n8 61.4229
R181 drain_left.n6 drain_left.n4 61.4227
R182 drain_left.n2 drain_left.n0 61.4227
R183 drain_left.n14 drain_left.n13 60.8798
R184 drain_left.n12 drain_left.n11 60.8798
R185 drain_left.n10 drain_left.n9 60.8798
R186 drain_left.n16 drain_left.n15 60.8796
R187 drain_left.n7 drain_left.n3 60.8796
R188 drain_left.n6 drain_left.n5 60.8796
R189 drain_left.n2 drain_left.n1 60.8796
R190 drain_left drain_left.n7 33.9846
R191 drain_left drain_left.n16 6.19632
R192 drain_left.n3 drain_left.t5 1.3205
R193 drain_left.n3 drain_left.t14 1.3205
R194 drain_left.n4 drain_left.t8 1.3205
R195 drain_left.n4 drain_left.t18 1.3205
R196 drain_left.n5 drain_left.t6 1.3205
R197 drain_left.n5 drain_left.t17 1.3205
R198 drain_left.n1 drain_left.t2 1.3205
R199 drain_left.n1 drain_left.t13 1.3205
R200 drain_left.n0 drain_left.t1 1.3205
R201 drain_left.n0 drain_left.t15 1.3205
R202 drain_left.n15 drain_left.t10 1.3205
R203 drain_left.n15 drain_left.t4 1.3205
R204 drain_left.n13 drain_left.t3 1.3205
R205 drain_left.n13 drain_left.t19 1.3205
R206 drain_left.n11 drain_left.t12 1.3205
R207 drain_left.n11 drain_left.t9 1.3205
R208 drain_left.n9 drain_left.t7 1.3205
R209 drain_left.n9 drain_left.t0 1.3205
R210 drain_left.n8 drain_left.t16 1.3205
R211 drain_left.n8 drain_left.t11 1.3205
R212 drain_left.n12 drain_left.n10 0.543603
R213 drain_left.n14 drain_left.n12 0.543603
R214 drain_left.n16 drain_left.n14 0.543603
R215 drain_left.n7 drain_left.n6 0.488257
R216 drain_left.n7 drain_left.n2 0.488257
R217 minus.n27 minus.t7 1358.36
R218 minus.n7 minus.t11 1358.36
R219 minus.n56 minus.t5 1358.36
R220 minus.n35 minus.t4 1358.36
R221 minus.n26 minus.t2 1309.43
R222 minus.n24 minus.t16 1309.43
R223 minus.n3 minus.t6 1309.43
R224 minus.n18 minus.t0 1309.43
R225 minus.n16 minus.t12 1309.43
R226 minus.n4 minus.t8 1309.43
R227 minus.n10 minus.t1 1309.43
R228 minus.n6 minus.t15 1309.43
R229 minus.n55 minus.t17 1309.43
R230 minus.n53 minus.t18 1309.43
R231 minus.n47 minus.t9 1309.43
R232 minus.n46 minus.t19 1309.43
R233 minus.n44 minus.t10 1309.43
R234 minus.n32 minus.t13 1309.43
R235 minus.n38 minus.t3 1309.43
R236 minus.n34 minus.t14 1309.43
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 64.9975
R264 minus.n15 minus.n4 64.9975
R265 minus.n43 minus.n32 64.9975
R266 minus.n48 minus.n47 64.9975
R267 minus.n25 minus.n24 62.0763
R268 minus.n10 minus.n9 62.0763
R269 minus.n38 minus.n37 62.0763
R270 minus.n54 minus.n53 62.0763
R271 minus.n18 minus.n17 46.0096
R272 minus.n17 minus.n16 46.0096
R273 minus.n45 minus.n44 46.0096
R274 minus.n46 minus.n45 46.0096
R275 minus.n27 minus.n26 43.0884
R276 minus.n7 minus.n6 43.0884
R277 minus.n35 minus.n34 43.0884
R278 minus.n56 minus.n55 43.0884
R279 minus.n58 minus.n28 39.3717
R280 minus.n26 minus.n25 29.9429
R281 minus.n9 minus.n6 29.9429
R282 minus.n37 minus.n34 29.9429
R283 minus.n55 minus.n54 29.9429
R284 minus.n19 minus.n18 27.0217
R285 minus.n16 minus.n15 27.0217
R286 minus.n44 minus.n43 27.0217
R287 minus.n48 minus.n46 27.0217
R288 minus.n24 minus.n23 10.955
R289 minus.n11 minus.n10 10.955
R290 minus.n39 minus.n38 10.955
R291 minus.n53 minus.n52 10.955
R292 minus.n3 minus.n1 8.03383
R293 minus.n12 minus.n4 8.03383
R294 minus.n40 minus.n32 8.03383
R295 minus.n47 minus.n30 8.03383
R296 minus.n58 minus.n57 6.51565
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 61.4227
R317 drain_right.n6 drain_right.n4 61.4227
R318 drain_right.n2 drain_right.n0 61.4227
R319 drain_right.n10 drain_right.n9 60.8798
R320 drain_right.n12 drain_right.n11 60.8798
R321 drain_right.n14 drain_right.n13 60.8798
R322 drain_right.n16 drain_right.n15 60.8798
R323 drain_right.n7 drain_right.n3 60.8796
R324 drain_right.n6 drain_right.n5 60.8796
R325 drain_right.n2 drain_right.n1 60.8796
R326 drain_right drain_right.n7 33.4314
R327 drain_right drain_right.n16 6.19632
R328 drain_right.n3 drain_right.t9 1.3205
R329 drain_right.n3 drain_right.t0 1.3205
R330 drain_right.n4 drain_right.t2 1.3205
R331 drain_right.n4 drain_right.t14 1.3205
R332 drain_right.n5 drain_right.t10 1.3205
R333 drain_right.n5 drain_right.t1 1.3205
R334 drain_right.n1 drain_right.t16 1.3205
R335 drain_right.n1 drain_right.t6 1.3205
R336 drain_right.n0 drain_right.t15 1.3205
R337 drain_right.n0 drain_right.t5 1.3205
R338 drain_right.n8 drain_right.t4 1.3205
R339 drain_right.n8 drain_right.t8 1.3205
R340 drain_right.n9 drain_right.t11 1.3205
R341 drain_right.n9 drain_right.t18 1.3205
R342 drain_right.n11 drain_right.t19 1.3205
R343 drain_right.n11 drain_right.t7 1.3205
R344 drain_right.n13 drain_right.t3 1.3205
R345 drain_right.n13 drain_right.t13 1.3205
R346 drain_right.n15 drain_right.t12 1.3205
R347 drain_right.n15 drain_right.t17 1.3205
R348 drain_right.n16 drain_right.n14 0.543603
R349 drain_right.n14 drain_right.n12 0.543603
R350 drain_right.n12 drain_right.n10 0.543603
R351 drain_right.n7 drain_right.n6 0.488257
R352 drain_right.n7 drain_right.n2 0.488257
C0 drain_left minus 0.171748f
C1 drain_right minus 8.82157f
C2 minus plus 6.33f
C3 drain_left drain_right 1.10832f
C4 drain_left plus 9.027519f
C5 drain_right plus 0.36079f
C6 minus source 8.447309f
C7 drain_left source 45.994102f
C8 drain_right source 45.9945f
C9 source plus 8.461349f
C10 drain_right a_n2102_n3888# 7.58873f
C11 drain_left a_n2102_n3888# 7.907589f
C12 source a_n2102_n3888# 10.417899f
C13 minus a_n2102_n3888# 8.447617f
C14 plus a_n2102_n3888# 10.66012f
C15 drain_right.t15 a_n2102_n3888# 0.405734f
C16 drain_right.t5 a_n2102_n3888# 0.405734f
C17 drain_right.n0 a_n2102_n3888# 3.67102f
C18 drain_right.t16 a_n2102_n3888# 0.405734f
C19 drain_right.t6 a_n2102_n3888# 0.405734f
C20 drain_right.n1 a_n2102_n3888# 3.66736f
C21 drain_right.n2 a_n2102_n3888# 0.805969f
C22 drain_right.t9 a_n2102_n3888# 0.405734f
C23 drain_right.t0 a_n2102_n3888# 0.405734f
C24 drain_right.n3 a_n2102_n3888# 3.66736f
C25 drain_right.t2 a_n2102_n3888# 0.405734f
C26 drain_right.t14 a_n2102_n3888# 0.405734f
C27 drain_right.n4 a_n2102_n3888# 3.67102f
C28 drain_right.t10 a_n2102_n3888# 0.405734f
C29 drain_right.t1 a_n2102_n3888# 0.405734f
C30 drain_right.n5 a_n2102_n3888# 3.66736f
C31 drain_right.n6 a_n2102_n3888# 0.805969f
C32 drain_right.n7 a_n2102_n3888# 2.28497f
C33 drain_right.t4 a_n2102_n3888# 0.405734f
C34 drain_right.t8 a_n2102_n3888# 0.405734f
C35 drain_right.n8 a_n2102_n3888# 3.67101f
C36 drain_right.t11 a_n2102_n3888# 0.405734f
C37 drain_right.t18 a_n2102_n3888# 0.405734f
C38 drain_right.n9 a_n2102_n3888# 3.66737f
C39 drain_right.n10 a_n2102_n3888# 0.810454f
C40 drain_right.t19 a_n2102_n3888# 0.405734f
C41 drain_right.t7 a_n2102_n3888# 0.405734f
C42 drain_right.n11 a_n2102_n3888# 3.66737f
C43 drain_right.n12 a_n2102_n3888# 0.400157f
C44 drain_right.t3 a_n2102_n3888# 0.405734f
C45 drain_right.t13 a_n2102_n3888# 0.405734f
C46 drain_right.n13 a_n2102_n3888# 3.66737f
C47 drain_right.n14 a_n2102_n3888# 0.400157f
C48 drain_right.t12 a_n2102_n3888# 0.405734f
C49 drain_right.t17 a_n2102_n3888# 0.405734f
C50 drain_right.n15 a_n2102_n3888# 3.66737f
C51 drain_right.n16 a_n2102_n3888# 0.685068f
C52 minus.n0 a_n2102_n3888# 0.049272f
C53 minus.t7 a_n2102_n3888# 0.63432f
C54 minus.t2 a_n2102_n3888# 0.625518f
C55 minus.t16 a_n2102_n3888# 0.625518f
C56 minus.n1 a_n2102_n3888# 0.018016f
C57 minus.n2 a_n2102_n3888# 0.049272f
C58 minus.t6 a_n2102_n3888# 0.625518f
C59 minus.n3 a_n2102_n3888# 0.240265f
C60 minus.t0 a_n2102_n3888# 0.625518f
C61 minus.t12 a_n2102_n3888# 0.625518f
C62 minus.t8 a_n2102_n3888# 0.625518f
C63 minus.n4 a_n2102_n3888# 0.240265f
C64 minus.n5 a_n2102_n3888# 0.049272f
C65 minus.t1 a_n2102_n3888# 0.625518f
C66 minus.t15 a_n2102_n3888# 0.625518f
C67 minus.n6 a_n2102_n3888# 0.240265f
C68 minus.t11 a_n2102_n3888# 0.63432f
C69 minus.n7 a_n2102_n3888# 0.255933f
C70 minus.n8 a_n2102_n3888# 0.112747f
C71 minus.n9 a_n2102_n3888# 0.020294f
C72 minus.n10 a_n2102_n3888# 0.240265f
C73 minus.n11 a_n2102_n3888# 0.018623f
C74 minus.n12 a_n2102_n3888# 0.018016f
C75 minus.n13 a_n2102_n3888# 0.049272f
C76 minus.n14 a_n2102_n3888# 0.049272f
C77 minus.n15 a_n2102_n3888# 0.020294f
C78 minus.n16 a_n2102_n3888# 0.240265f
C79 minus.n17 a_n2102_n3888# 0.020294f
C80 minus.n18 a_n2102_n3888# 0.240265f
C81 minus.n19 a_n2102_n3888# 0.020294f
C82 minus.n20 a_n2102_n3888# 0.049272f
C83 minus.n21 a_n2102_n3888# 0.049272f
C84 minus.n22 a_n2102_n3888# 0.049272f
C85 minus.n23 a_n2102_n3888# 0.018623f
C86 minus.n24 a_n2102_n3888# 0.240265f
C87 minus.n25 a_n2102_n3888# 0.020294f
C88 minus.n26 a_n2102_n3888# 0.240265f
C89 minus.n27 a_n2102_n3888# 0.255858f
C90 minus.n28 a_n2102_n3888# 1.9822f
C91 minus.n29 a_n2102_n3888# 0.049272f
C92 minus.t17 a_n2102_n3888# 0.625518f
C93 minus.t18 a_n2102_n3888# 0.625518f
C94 minus.n30 a_n2102_n3888# 0.018016f
C95 minus.n31 a_n2102_n3888# 0.049272f
C96 minus.t19 a_n2102_n3888# 0.625518f
C97 minus.t10 a_n2102_n3888# 0.625518f
C98 minus.t13 a_n2102_n3888# 0.625518f
C99 minus.n32 a_n2102_n3888# 0.240265f
C100 minus.n33 a_n2102_n3888# 0.049272f
C101 minus.t3 a_n2102_n3888# 0.625518f
C102 minus.t14 a_n2102_n3888# 0.625518f
C103 minus.n34 a_n2102_n3888# 0.240265f
C104 minus.t4 a_n2102_n3888# 0.63432f
C105 minus.n35 a_n2102_n3888# 0.255933f
C106 minus.n36 a_n2102_n3888# 0.112747f
C107 minus.n37 a_n2102_n3888# 0.020294f
C108 minus.n38 a_n2102_n3888# 0.240265f
C109 minus.n39 a_n2102_n3888# 0.018623f
C110 minus.n40 a_n2102_n3888# 0.018016f
C111 minus.n41 a_n2102_n3888# 0.049272f
C112 minus.n42 a_n2102_n3888# 0.049272f
C113 minus.n43 a_n2102_n3888# 0.020294f
C114 minus.n44 a_n2102_n3888# 0.240265f
C115 minus.n45 a_n2102_n3888# 0.020294f
C116 minus.n46 a_n2102_n3888# 0.240265f
C117 minus.t9 a_n2102_n3888# 0.625518f
C118 minus.n47 a_n2102_n3888# 0.240265f
C119 minus.n48 a_n2102_n3888# 0.020294f
C120 minus.n49 a_n2102_n3888# 0.049272f
C121 minus.n50 a_n2102_n3888# 0.049272f
C122 minus.n51 a_n2102_n3888# 0.049272f
C123 minus.n52 a_n2102_n3888# 0.018623f
C124 minus.n53 a_n2102_n3888# 0.240265f
C125 minus.n54 a_n2102_n3888# 0.020294f
C126 minus.n55 a_n2102_n3888# 0.240265f
C127 minus.t5 a_n2102_n3888# 0.63432f
C128 minus.n56 a_n2102_n3888# 0.255858f
C129 minus.n57 a_n2102_n3888# 0.323943f
C130 minus.n58 a_n2102_n3888# 2.38476f
C131 drain_left.t1 a_n2102_n3888# 0.406223f
C132 drain_left.t15 a_n2102_n3888# 0.406223f
C133 drain_left.n0 a_n2102_n3888# 3.67544f
C134 drain_left.t2 a_n2102_n3888# 0.406223f
C135 drain_left.t13 a_n2102_n3888# 0.406223f
C136 drain_left.n1 a_n2102_n3888# 3.67178f
C137 drain_left.n2 a_n2102_n3888# 0.806939f
C138 drain_left.t5 a_n2102_n3888# 0.406223f
C139 drain_left.t14 a_n2102_n3888# 0.406223f
C140 drain_left.n3 a_n2102_n3888# 3.67178f
C141 drain_left.t8 a_n2102_n3888# 0.406223f
C142 drain_left.t18 a_n2102_n3888# 0.406223f
C143 drain_left.n4 a_n2102_n3888# 3.67544f
C144 drain_left.t6 a_n2102_n3888# 0.406223f
C145 drain_left.t17 a_n2102_n3888# 0.406223f
C146 drain_left.n5 a_n2102_n3888# 3.67178f
C147 drain_left.n6 a_n2102_n3888# 0.806939f
C148 drain_left.n7 a_n2102_n3888# 2.35873f
C149 drain_left.t16 a_n2102_n3888# 0.406223f
C150 drain_left.t11 a_n2102_n3888# 0.406223f
C151 drain_left.n8 a_n2102_n3888# 3.67544f
C152 drain_left.t7 a_n2102_n3888# 0.406223f
C153 drain_left.t0 a_n2102_n3888# 0.406223f
C154 drain_left.n9 a_n2102_n3888# 3.67178f
C155 drain_left.n10 a_n2102_n3888# 0.811416f
C156 drain_left.t12 a_n2102_n3888# 0.406223f
C157 drain_left.t9 a_n2102_n3888# 0.406223f
C158 drain_left.n11 a_n2102_n3888# 3.67178f
C159 drain_left.n12 a_n2102_n3888# 0.400639f
C160 drain_left.t3 a_n2102_n3888# 0.406223f
C161 drain_left.t19 a_n2102_n3888# 0.406223f
C162 drain_left.n13 a_n2102_n3888# 3.67178f
C163 drain_left.n14 a_n2102_n3888# 0.400639f
C164 drain_left.t10 a_n2102_n3888# 0.406223f
C165 drain_left.t4 a_n2102_n3888# 0.406223f
C166 drain_left.n15 a_n2102_n3888# 3.67177f
C167 drain_left.n16 a_n2102_n3888# 0.685905f
C168 source.t19 a_n2102_n3888# 3.90603f
C169 source.n0 a_n2102_n3888# 1.8092f
C170 source.t26 a_n2102_n3888# 0.348547f
C171 source.t28 a_n2102_n3888# 0.348547f
C172 source.n1 a_n2102_n3888# 3.0617f
C173 source.n2 a_n2102_n3888# 0.392556f
C174 source.t36 a_n2102_n3888# 0.348547f
C175 source.t20 a_n2102_n3888# 0.348547f
C176 source.n3 a_n2102_n3888# 3.0617f
C177 source.n4 a_n2102_n3888# 0.392556f
C178 source.t33 a_n2102_n3888# 0.348547f
C179 source.t18 a_n2102_n3888# 0.348547f
C180 source.n5 a_n2102_n3888# 3.0617f
C181 source.n6 a_n2102_n3888# 0.392556f
C182 source.t37 a_n2102_n3888# 0.348547f
C183 source.t25 a_n2102_n3888# 0.348547f
C184 source.n7 a_n2102_n3888# 3.0617f
C185 source.n8 a_n2102_n3888# 0.392556f
C186 source.t27 a_n2102_n3888# 3.90604f
C187 source.n9 a_n2102_n3888# 0.491854f
C188 source.t4 a_n2102_n3888# 3.90604f
C189 source.n10 a_n2102_n3888# 0.491854f
C190 source.t2 a_n2102_n3888# 0.348547f
C191 source.t14 a_n2102_n3888# 0.348547f
C192 source.n11 a_n2102_n3888# 3.0617f
C193 source.n12 a_n2102_n3888# 0.392556f
C194 source.t0 a_n2102_n3888# 0.348547f
C195 source.t9 a_n2102_n3888# 0.348547f
C196 source.n13 a_n2102_n3888# 3.0617f
C197 source.n14 a_n2102_n3888# 0.392556f
C198 source.t16 a_n2102_n3888# 0.348547f
C199 source.t15 a_n2102_n3888# 0.348547f
C200 source.n15 a_n2102_n3888# 3.0617f
C201 source.n16 a_n2102_n3888# 0.392556f
C202 source.t8 a_n2102_n3888# 0.348547f
C203 source.t7 a_n2102_n3888# 0.348547f
C204 source.n17 a_n2102_n3888# 3.0617f
C205 source.n18 a_n2102_n3888# 0.392556f
C206 source.t10 a_n2102_n3888# 3.90604f
C207 source.n19 a_n2102_n3888# 2.29808f
C208 source.t31 a_n2102_n3888# 3.90603f
C209 source.n20 a_n2102_n3888# 2.29808f
C210 source.t22 a_n2102_n3888# 0.348547f
C211 source.t32 a_n2102_n3888# 0.348547f
C212 source.n21 a_n2102_n3888# 3.06169f
C213 source.n22 a_n2102_n3888# 0.39256f
C214 source.t29 a_n2102_n3888# 0.348547f
C215 source.t30 a_n2102_n3888# 0.348547f
C216 source.n23 a_n2102_n3888# 3.06169f
C217 source.n24 a_n2102_n3888# 0.39256f
C218 source.t21 a_n2102_n3888# 0.348547f
C219 source.t23 a_n2102_n3888# 0.348547f
C220 source.n25 a_n2102_n3888# 3.06169f
C221 source.n26 a_n2102_n3888# 0.39256f
C222 source.t24 a_n2102_n3888# 0.348547f
C223 source.t34 a_n2102_n3888# 0.348547f
C224 source.n27 a_n2102_n3888# 3.06169f
C225 source.n28 a_n2102_n3888# 0.39256f
C226 source.t35 a_n2102_n3888# 3.90603f
C227 source.n29 a_n2102_n3888# 0.491859f
C228 source.t5 a_n2102_n3888# 3.90603f
C229 source.n30 a_n2102_n3888# 0.491859f
C230 source.t12 a_n2102_n3888# 0.348547f
C231 source.t1 a_n2102_n3888# 0.348547f
C232 source.n31 a_n2102_n3888# 3.06169f
C233 source.n32 a_n2102_n3888# 0.39256f
C234 source.t17 a_n2102_n3888# 0.348547f
C235 source.t39 a_n2102_n3888# 0.348547f
C236 source.n33 a_n2102_n3888# 3.06169f
C237 source.n34 a_n2102_n3888# 0.39256f
C238 source.t6 a_n2102_n3888# 0.348547f
C239 source.t38 a_n2102_n3888# 0.348547f
C240 source.n35 a_n2102_n3888# 3.06169f
C241 source.n36 a_n2102_n3888# 0.39256f
C242 source.t13 a_n2102_n3888# 0.348547f
C243 source.t11 a_n2102_n3888# 0.348547f
C244 source.n37 a_n2102_n3888# 3.06169f
C245 source.n38 a_n2102_n3888# 0.39256f
C246 source.t3 a_n2102_n3888# 3.90603f
C247 source.n39 a_n2102_n3888# 0.657848f
C248 source.n40 a_n2102_n3888# 2.15003f
C249 plus.n0 a_n2102_n3888# 0.050113f
C250 plus.t9 a_n2102_n3888# 0.6362f
C251 plus.t0 a_n2102_n3888# 0.6362f
C252 plus.n1 a_n2102_n3888# 0.018324f
C253 plus.n2 a_n2102_n3888# 0.050113f
C254 plus.t10 a_n2102_n3888# 0.6362f
C255 plus.t7 a_n2102_n3888# 0.6362f
C256 plus.t19 a_n2102_n3888# 0.6362f
C257 plus.n3 a_n2102_n3888# 0.244368f
C258 plus.n4 a_n2102_n3888# 0.050113f
C259 plus.t12 a_n2102_n3888# 0.6362f
C260 plus.t8 a_n2102_n3888# 0.6362f
C261 plus.n5 a_n2102_n3888# 0.244368f
C262 plus.t3 a_n2102_n3888# 0.645153f
C263 plus.n6 a_n2102_n3888# 0.260303f
C264 plus.n7 a_n2102_n3888# 0.114673f
C265 plus.n8 a_n2102_n3888# 0.020641f
C266 plus.n9 a_n2102_n3888# 0.244368f
C267 plus.n10 a_n2102_n3888# 0.018942f
C268 plus.n11 a_n2102_n3888# 0.018324f
C269 plus.n12 a_n2102_n3888# 0.050113f
C270 plus.n13 a_n2102_n3888# 0.050113f
C271 plus.n14 a_n2102_n3888# 0.020641f
C272 plus.n15 a_n2102_n3888# 0.244368f
C273 plus.n16 a_n2102_n3888# 0.020641f
C274 plus.n17 a_n2102_n3888# 0.244368f
C275 plus.t16 a_n2102_n3888# 0.6362f
C276 plus.n18 a_n2102_n3888# 0.244368f
C277 plus.n19 a_n2102_n3888# 0.020641f
C278 plus.n20 a_n2102_n3888# 0.050113f
C279 plus.n21 a_n2102_n3888# 0.050113f
C280 plus.n22 a_n2102_n3888# 0.050113f
C281 plus.n23 a_n2102_n3888# 0.018942f
C282 plus.n24 a_n2102_n3888# 0.244368f
C283 plus.n25 a_n2102_n3888# 0.020641f
C284 plus.n26 a_n2102_n3888# 0.244368f
C285 plus.t15 a_n2102_n3888# 0.645153f
C286 plus.n27 a_n2102_n3888# 0.260228f
C287 plus.n28 a_n2102_n3888# 0.635124f
C288 plus.n29 a_n2102_n3888# 0.050113f
C289 plus.t18 a_n2102_n3888# 0.645153f
C290 plus.t4 a_n2102_n3888# 0.6362f
C291 plus.t17 a_n2102_n3888# 0.6362f
C292 plus.n30 a_n2102_n3888# 0.018324f
C293 plus.n31 a_n2102_n3888# 0.050113f
C294 plus.t6 a_n2102_n3888# 0.6362f
C295 plus.n32 a_n2102_n3888# 0.244368f
C296 plus.t14 a_n2102_n3888# 0.6362f
C297 plus.t5 a_n2102_n3888# 0.6362f
C298 plus.t13 a_n2102_n3888# 0.6362f
C299 plus.n33 a_n2102_n3888# 0.244368f
C300 plus.n34 a_n2102_n3888# 0.050113f
C301 plus.t2 a_n2102_n3888# 0.6362f
C302 plus.t11 a_n2102_n3888# 0.6362f
C303 plus.n35 a_n2102_n3888# 0.244368f
C304 plus.t1 a_n2102_n3888# 0.645153f
C305 plus.n36 a_n2102_n3888# 0.260303f
C306 plus.n37 a_n2102_n3888# 0.114673f
C307 plus.n38 a_n2102_n3888# 0.020641f
C308 plus.n39 a_n2102_n3888# 0.244368f
C309 plus.n40 a_n2102_n3888# 0.018942f
C310 plus.n41 a_n2102_n3888# 0.018324f
C311 plus.n42 a_n2102_n3888# 0.050113f
C312 plus.n43 a_n2102_n3888# 0.050113f
C313 plus.n44 a_n2102_n3888# 0.020641f
C314 plus.n45 a_n2102_n3888# 0.244368f
C315 plus.n46 a_n2102_n3888# 0.020641f
C316 plus.n47 a_n2102_n3888# 0.244368f
C317 plus.n48 a_n2102_n3888# 0.020641f
C318 plus.n49 a_n2102_n3888# 0.050113f
C319 plus.n50 a_n2102_n3888# 0.050113f
C320 plus.n51 a_n2102_n3888# 0.050113f
C321 plus.n52 a_n2102_n3888# 0.018942f
C322 plus.n53 a_n2102_n3888# 0.244368f
C323 plus.n54 a_n2102_n3888# 0.020641f
C324 plus.n55 a_n2102_n3888# 0.244368f
C325 plus.n56 a_n2102_n3888# 0.260228f
C326 plus.n57 a_n2102_n3888# 1.66379f
.ends

