* NGSPICE file created from diffpair409.ext - technology: sky130A

.subckt diffpair409 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t35 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X1 source.t34 minus.t1 drain_right.t22 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X2 source.t12 plus.t0 drain_left.t23 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X3 drain_left.t22 plus.t1 source.t5 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X4 drain_left.t21 plus.t2 source.t14 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X5 source.t6 plus.t3 drain_left.t20 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X6 drain_left.t19 plus.t4 source.t19 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X7 source.t23 plus.t5 drain_left.t18 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X8 drain_right.t21 minus.t2 source.t33 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X9 source.t13 plus.t6 drain_left.t17 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X10 a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X11 drain_left.t16 plus.t7 source.t0 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X12 a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X13 source.t45 minus.t3 drain_right.t20 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X14 a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X15 source.t26 minus.t4 drain_right.t19 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X16 drain_left.t15 plus.t8 source.t4 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X17 source.t29 minus.t5 drain_right.t18 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X18 drain_left.t14 plus.t9 source.t9 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 drain_right.t17 minus.t6 source.t36 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X20 drain_right.t16 minus.t7 source.t41 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X21 drain_right.t15 minus.t8 source.t30 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X22 source.t38 minus.t9 drain_right.t14 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X23 drain_right.t13 minus.t10 source.t24 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X24 drain_right.t12 minus.t11 source.t47 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X25 drain_right.t11 minus.t12 source.t37 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X26 source.t16 plus.t10 drain_left.t13 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X27 drain_left.t12 plus.t11 source.t21 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X28 source.t1 plus.t12 drain_left.t11 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X29 drain_right.t10 minus.t13 source.t46 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X30 drain_right.t9 minus.t14 source.t44 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X31 source.t8 plus.t13 drain_left.t10 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X32 source.t32 minus.t15 drain_right.t8 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X33 source.t31 minus.t16 drain_right.t7 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X34 drain_left.t9 plus.t14 source.t10 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X35 source.t39 minus.t17 drain_right.t6 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X36 source.t27 minus.t18 drain_right.t5 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X37 a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X38 drain_right.t4 minus.t19 source.t28 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X39 drain_left.t8 plus.t15 source.t15 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X40 source.t20 plus.t16 drain_left.t7 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X41 source.t11 plus.t17 drain_left.t6 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X42 source.t42 minus.t20 drain_right.t3 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X43 source.t40 minus.t21 drain_right.t2 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X44 source.t43 minus.t22 drain_right.t1 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X45 source.t18 plus.t18 drain_left.t5 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X46 drain_left.t4 plus.t19 source.t17 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X47 drain_left.t3 plus.t20 source.t22 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X48 drain_left.t2 plus.t21 source.t3 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X49 source.t7 plus.t22 drain_left.t1 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X50 drain_right.t0 minus.t23 source.t25 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X51 source.t2 plus.t23 drain_left.t0 a_n2406_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
R0 minus.n35 minus.t16 2184.34
R1 minus.n8 minus.t6 2184.34
R2 minus.n72 minus.t2 2184.34
R3 minus.n43 minus.t1 2184.34
R4 minus.n34 minus.t19 2136.87
R5 minus.n32 minus.t21 2136.87
R6 minus.n3 minus.t11 2136.87
R7 minus.n26 minus.t15 2136.87
R8 minus.n24 minus.t14 2136.87
R9 minus.n6 minus.t17 2136.87
R10 minus.n18 minus.t7 2136.87
R11 minus.n16 minus.t9 2136.87
R12 minus.n9 minus.t13 2136.87
R13 minus.n10 minus.t5 2136.87
R14 minus.n71 minus.t22 2136.87
R15 minus.n69 minus.t12 2136.87
R16 minus.n63 minus.t4 2136.87
R17 minus.n62 minus.t0 2136.87
R18 minus.n60 minus.t20 2136.87
R19 minus.n54 minus.t10 2136.87
R20 minus.n53 minus.t3 2136.87
R21 minus.n51 minus.t23 2136.87
R22 minus.n45 minus.t18 2136.87
R23 minus.n44 minus.t8 2136.87
R24 minus.n12 minus.n8 161.489
R25 minus.n47 minus.n43 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n31 minus.n30 161.3
R29 minus.n29 minus.n1 161.3
R30 minus.n28 minus.n27 161.3
R31 minus.n25 minus.n2 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n20 minus.n19 161.3
R35 minus.n17 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n7 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n68 minus.n67 161.3
R42 minus.n66 minus.n38 161.3
R43 minus.n65 minus.n64 161.3
R44 minus.n61 minus.n39 161.3
R45 minus.n59 minus.n58 161.3
R46 minus.n57 minus.n40 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n52 minus.n41 161.3
R49 minus.n50 minus.n49 161.3
R50 minus.n48 minus.n42 161.3
R51 minus.n47 minus.n46 161.3
R52 minus.n31 minus.n1 73.0308
R53 minus.n23 minus.n4 73.0308
R54 minus.n15 minus.n7 73.0308
R55 minus.n50 minus.n42 73.0308
R56 minus.n59 minus.n40 73.0308
R57 minus.n68 minus.n38 73.0308
R58 minus.n33 minus.n32 69.3793
R59 minus.n11 minus.n9 69.3793
R60 minus.n46 minus.n45 69.3793
R61 minus.n70 minus.n69 69.3793
R62 minus.n25 minus.n24 62.0763
R63 minus.n19 minus.n6 62.0763
R64 minus.n55 minus.n54 62.0763
R65 minus.n61 minus.n60 62.0763
R66 minus.n27 minus.n3 54.7732
R67 minus.n17 minus.n16 54.7732
R68 minus.n52 minus.n51 54.7732
R69 minus.n64 minus.n63 54.7732
R70 minus.n35 minus.n34 47.4702
R71 minus.n10 minus.n8 47.4702
R72 minus.n44 minus.n43 47.4702
R73 minus.n72 minus.n71 47.4702
R74 minus.n27 minus.n26 40.1672
R75 minus.n18 minus.n17 40.1672
R76 minus.n53 minus.n52 40.1672
R77 minus.n64 minus.n62 40.1672
R78 minus.n74 minus.n36 38.2581
R79 minus.n26 minus.n25 32.8641
R80 minus.n19 minus.n18 32.8641
R81 minus.n55 minus.n53 32.8641
R82 minus.n62 minus.n61 32.8641
R83 minus.n34 minus.n33 25.5611
R84 minus.n11 minus.n10 25.5611
R85 minus.n46 minus.n44 25.5611
R86 minus.n71 minus.n70 25.5611
R87 minus.n3 minus.n1 18.2581
R88 minus.n16 minus.n15 18.2581
R89 minus.n51 minus.n50 18.2581
R90 minus.n63 minus.n38 18.2581
R91 minus.n24 minus.n23 10.955
R92 minus.n6 minus.n4 10.955
R93 minus.n54 minus.n40 10.955
R94 minus.n60 minus.n59 10.955
R95 minus.n74 minus.n73 6.52323
R96 minus.n32 minus.n31 3.65202
R97 minus.n9 minus.n7 3.65202
R98 minus.n45 minus.n42 3.65202
R99 minus.n69 minus.n68 3.65202
R100 minus.n36 minus.n0 0.189894
R101 minus.n30 minus.n0 0.189894
R102 minus.n30 minus.n29 0.189894
R103 minus.n29 minus.n28 0.189894
R104 minus.n28 minus.n2 0.189894
R105 minus.n22 minus.n2 0.189894
R106 minus.n22 minus.n21 0.189894
R107 minus.n21 minus.n20 0.189894
R108 minus.n20 minus.n5 0.189894
R109 minus.n14 minus.n5 0.189894
R110 minus.n14 minus.n13 0.189894
R111 minus.n13 minus.n12 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n49 minus.n48 0.189894
R114 minus.n49 minus.n41 0.189894
R115 minus.n56 minus.n41 0.189894
R116 minus.n57 minus.n56 0.189894
R117 minus.n58 minus.n57 0.189894
R118 minus.n58 minus.n39 0.189894
R119 minus.n65 minus.n39 0.189894
R120 minus.n66 minus.n65 0.189894
R121 minus.n67 minus.n66 0.189894
R122 minus.n67 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 source.n11 source.t1 45.3739
R126 source.n12 source.t36 45.3739
R127 source.n23 source.t31 45.3739
R128 source.n47 source.t33 45.3737
R129 source.n36 source.t34 45.3737
R130 source.n35 source.t4 45.3737
R131 source.n24 source.t23 45.3737
R132 source.n0 source.t3 45.3737
R133 source.n2 source.n1 42.8739
R134 source.n4 source.n3 42.8739
R135 source.n6 source.n5 42.8739
R136 source.n8 source.n7 42.8739
R137 source.n10 source.n9 42.8739
R138 source.n14 source.n13 42.8739
R139 source.n16 source.n15 42.8739
R140 source.n18 source.n17 42.8739
R141 source.n20 source.n19 42.8739
R142 source.n22 source.n21 42.8739
R143 source.n46 source.n45 42.8737
R144 source.n44 source.n43 42.8737
R145 source.n42 source.n41 42.8737
R146 source.n40 source.n39 42.8737
R147 source.n38 source.n37 42.8737
R148 source.n34 source.n33 42.8737
R149 source.n32 source.n31 42.8737
R150 source.n30 source.n29 42.8737
R151 source.n28 source.n27 42.8737
R152 source.n26 source.n25 42.8737
R153 source.n24 source.n23 21.8481
R154 source.n48 source.n0 16.305
R155 source.n48 source.n47 5.5436
R156 source.n45 source.t37 2.5005
R157 source.n45 source.t43 2.5005
R158 source.n43 source.t35 2.5005
R159 source.n43 source.t26 2.5005
R160 source.n41 source.t24 2.5005
R161 source.n41 source.t42 2.5005
R162 source.n39 source.t25 2.5005
R163 source.n39 source.t45 2.5005
R164 source.n37 source.t30 2.5005
R165 source.n37 source.t27 2.5005
R166 source.n33 source.t14 2.5005
R167 source.n33 source.t16 2.5005
R168 source.n31 source.t9 2.5005
R169 source.n31 source.t13 2.5005
R170 source.n29 source.t19 2.5005
R171 source.n29 source.t12 2.5005
R172 source.n27 source.t0 2.5005
R173 source.n27 source.t6 2.5005
R174 source.n25 source.t5 2.5005
R175 source.n25 source.t2 2.5005
R176 source.n1 source.t15 2.5005
R177 source.n1 source.t8 2.5005
R178 source.n3 source.t21 2.5005
R179 source.n3 source.t18 2.5005
R180 source.n5 source.t17 2.5005
R181 source.n5 source.t20 2.5005
R182 source.n7 source.t10 2.5005
R183 source.n7 source.t7 2.5005
R184 source.n9 source.t22 2.5005
R185 source.n9 source.t11 2.5005
R186 source.n13 source.t46 2.5005
R187 source.n13 source.t29 2.5005
R188 source.n15 source.t41 2.5005
R189 source.n15 source.t38 2.5005
R190 source.n17 source.t44 2.5005
R191 source.n17 source.t39 2.5005
R192 source.n19 source.t47 2.5005
R193 source.n19 source.t32 2.5005
R194 source.n21 source.t28 2.5005
R195 source.n21 source.t40 2.5005
R196 source.n23 source.n22 0.560845
R197 source.n22 source.n20 0.560845
R198 source.n20 source.n18 0.560845
R199 source.n18 source.n16 0.560845
R200 source.n16 source.n14 0.560845
R201 source.n14 source.n12 0.560845
R202 source.n11 source.n10 0.560845
R203 source.n10 source.n8 0.560845
R204 source.n8 source.n6 0.560845
R205 source.n6 source.n4 0.560845
R206 source.n4 source.n2 0.560845
R207 source.n2 source.n0 0.560845
R208 source.n26 source.n24 0.560845
R209 source.n28 source.n26 0.560845
R210 source.n30 source.n28 0.560845
R211 source.n32 source.n30 0.560845
R212 source.n34 source.n32 0.560845
R213 source.n35 source.n34 0.560845
R214 source.n38 source.n36 0.560845
R215 source.n40 source.n38 0.560845
R216 source.n42 source.n40 0.560845
R217 source.n44 source.n42 0.560845
R218 source.n46 source.n44 0.560845
R219 source.n47 source.n46 0.560845
R220 source.n12 source.n11 0.470328
R221 source.n36 source.n35 0.470328
R222 source source.n48 0.188
R223 drain_right.n7 drain_right.n5 60.1128
R224 drain_right.n2 drain_right.n0 60.1128
R225 drain_right.n13 drain_right.n11 60.1128
R226 drain_right.n13 drain_right.n12 59.5527
R227 drain_right.n15 drain_right.n14 59.5527
R228 drain_right.n17 drain_right.n16 59.5527
R229 drain_right.n19 drain_right.n18 59.5527
R230 drain_right.n21 drain_right.n20 59.5527
R231 drain_right.n7 drain_right.n6 59.5525
R232 drain_right.n9 drain_right.n8 59.5525
R233 drain_right.n4 drain_right.n3 59.5525
R234 drain_right.n2 drain_right.n1 59.5525
R235 drain_right drain_right.n10 32.1371
R236 drain_right drain_right.n21 6.21356
R237 drain_right.n5 drain_right.t1 2.5005
R238 drain_right.n5 drain_right.t21 2.5005
R239 drain_right.n6 drain_right.t19 2.5005
R240 drain_right.n6 drain_right.t11 2.5005
R241 drain_right.n8 drain_right.t3 2.5005
R242 drain_right.n8 drain_right.t23 2.5005
R243 drain_right.n3 drain_right.t20 2.5005
R244 drain_right.n3 drain_right.t13 2.5005
R245 drain_right.n1 drain_right.t5 2.5005
R246 drain_right.n1 drain_right.t0 2.5005
R247 drain_right.n0 drain_right.t22 2.5005
R248 drain_right.n0 drain_right.t15 2.5005
R249 drain_right.n11 drain_right.t18 2.5005
R250 drain_right.n11 drain_right.t17 2.5005
R251 drain_right.n12 drain_right.t14 2.5005
R252 drain_right.n12 drain_right.t10 2.5005
R253 drain_right.n14 drain_right.t6 2.5005
R254 drain_right.n14 drain_right.t16 2.5005
R255 drain_right.n16 drain_right.t8 2.5005
R256 drain_right.n16 drain_right.t9 2.5005
R257 drain_right.n18 drain_right.t2 2.5005
R258 drain_right.n18 drain_right.t12 2.5005
R259 drain_right.n20 drain_right.t7 2.5005
R260 drain_right.n20 drain_right.t4 2.5005
R261 drain_right.n9 drain_right.n7 0.560845
R262 drain_right.n4 drain_right.n2 0.560845
R263 drain_right.n21 drain_right.n19 0.560845
R264 drain_right.n19 drain_right.n17 0.560845
R265 drain_right.n17 drain_right.n15 0.560845
R266 drain_right.n15 drain_right.n13 0.560845
R267 drain_right.n10 drain_right.n9 0.225326
R268 drain_right.n10 drain_right.n4 0.225326
R269 plus.n6 plus.t12 2184.34
R270 plus.n35 plus.t21 2184.34
R271 plus.n45 plus.t8 2184.34
R272 plus.n72 plus.t5 2184.34
R273 plus.n7 plus.t20 2136.87
R274 plus.n8 plus.t17 2136.87
R275 plus.n14 plus.t14 2136.87
R276 plus.n16 plus.t22 2136.87
R277 plus.n17 plus.t19 2136.87
R278 plus.n23 plus.t16 2136.87
R279 plus.n25 plus.t11 2136.87
R280 plus.n26 plus.t18 2136.87
R281 plus.n32 plus.t15 2136.87
R282 plus.n34 plus.t13 2136.87
R283 plus.n47 plus.t10 2136.87
R284 plus.n46 plus.t2 2136.87
R285 plus.n53 plus.t6 2136.87
R286 plus.n55 plus.t9 2136.87
R287 plus.n43 plus.t0 2136.87
R288 plus.n61 plus.t4 2136.87
R289 plus.n63 plus.t3 2136.87
R290 plus.n40 plus.t7 2136.87
R291 plus.n69 plus.t23 2136.87
R292 plus.n71 plus.t1 2136.87
R293 plus.n10 plus.n6 161.489
R294 plus.n49 plus.n45 161.489
R295 plus.n10 plus.n9 161.3
R296 plus.n11 plus.n5 161.3
R297 plus.n13 plus.n12 161.3
R298 plus.n15 plus.n4 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n3 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n24 plus.n2 161.3
R303 plus.n28 plus.n27 161.3
R304 plus.n29 plus.n1 161.3
R305 plus.n31 plus.n30 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n49 plus.n48 161.3
R309 plus.n50 plus.n44 161.3
R310 plus.n52 plus.n51 161.3
R311 plus.n54 plus.n42 161.3
R312 plus.n57 plus.n56 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n39 161.3
R316 plus.n65 plus.n64 161.3
R317 plus.n66 plus.n38 161.3
R318 plus.n68 plus.n67 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n13 plus.n5 73.0308
R322 plus.n22 plus.n3 73.0308
R323 plus.n31 plus.n1 73.0308
R324 plus.n68 plus.n38 73.0308
R325 plus.n60 plus.n41 73.0308
R326 plus.n52 plus.n44 73.0308
R327 plus.n9 plus.n8 69.3793
R328 plus.n33 plus.n32 69.3793
R329 plus.n70 plus.n69 69.3793
R330 plus.n48 plus.n46 69.3793
R331 plus.n18 plus.n17 62.0763
R332 plus.n24 plus.n23 62.0763
R333 plus.n62 plus.n61 62.0763
R334 plus.n56 plus.n43 62.0763
R335 plus.n15 plus.n14 54.7732
R336 plus.n27 plus.n26 54.7732
R337 plus.n64 plus.n40 54.7732
R338 plus.n54 plus.n53 54.7732
R339 plus.n7 plus.n6 47.4702
R340 plus.n35 plus.n34 47.4702
R341 plus.n72 plus.n71 47.4702
R342 plus.n47 plus.n45 47.4702
R343 plus.n16 plus.n15 40.1672
R344 plus.n27 plus.n25 40.1672
R345 plus.n64 plus.n63 40.1672
R346 plus.n55 plus.n54 40.1672
R347 plus.n18 plus.n16 32.8641
R348 plus.n25 plus.n24 32.8641
R349 plus.n63 plus.n62 32.8641
R350 plus.n56 plus.n55 32.8641
R351 plus plus.n73 32.1392
R352 plus.n9 plus.n7 25.5611
R353 plus.n34 plus.n33 25.5611
R354 plus.n71 plus.n70 25.5611
R355 plus.n48 plus.n47 25.5611
R356 plus.n14 plus.n13 18.2581
R357 plus.n26 plus.n1 18.2581
R358 plus.n40 plus.n38 18.2581
R359 plus.n53 plus.n52 18.2581
R360 plus plus.n36 12.1672
R361 plus.n17 plus.n3 10.955
R362 plus.n23 plus.n22 10.955
R363 plus.n61 plus.n60 10.955
R364 plus.n43 plus.n41 10.955
R365 plus.n8 plus.n5 3.65202
R366 plus.n32 plus.n31 3.65202
R367 plus.n69 plus.n68 3.65202
R368 plus.n46 plus.n44 3.65202
R369 plus.n11 plus.n10 0.189894
R370 plus.n12 plus.n11 0.189894
R371 plus.n12 plus.n4 0.189894
R372 plus.n19 plus.n4 0.189894
R373 plus.n20 plus.n19 0.189894
R374 plus.n21 plus.n20 0.189894
R375 plus.n21 plus.n2 0.189894
R376 plus.n28 plus.n2 0.189894
R377 plus.n29 plus.n28 0.189894
R378 plus.n30 plus.n29 0.189894
R379 plus.n30 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n67 plus.n37 0.189894
R383 plus.n67 plus.n66 0.189894
R384 plus.n66 plus.n65 0.189894
R385 plus.n65 plus.n39 0.189894
R386 plus.n59 plus.n39 0.189894
R387 plus.n59 plus.n58 0.189894
R388 plus.n58 plus.n57 0.189894
R389 plus.n57 plus.n42 0.189894
R390 plus.n51 plus.n42 0.189894
R391 plus.n51 plus.n50 0.189894
R392 plus.n50 plus.n49 0.189894
R393 drain_left.n13 drain_left.n11 60.113
R394 drain_left.n7 drain_left.n5 60.1128
R395 drain_left.n2 drain_left.n0 60.1128
R396 drain_left.n19 drain_left.n18 59.5527
R397 drain_left.n17 drain_left.n16 59.5527
R398 drain_left.n15 drain_left.n14 59.5527
R399 drain_left.n13 drain_left.n12 59.5527
R400 drain_left.n7 drain_left.n6 59.5525
R401 drain_left.n9 drain_left.n8 59.5525
R402 drain_left.n4 drain_left.n3 59.5525
R403 drain_left.n2 drain_left.n1 59.5525
R404 drain_left.n21 drain_left.n20 59.5525
R405 drain_left drain_left.n10 32.6903
R406 drain_left drain_left.n21 6.21356
R407 drain_left.n5 drain_left.t13 2.5005
R408 drain_left.n5 drain_left.t15 2.5005
R409 drain_left.n6 drain_left.t17 2.5005
R410 drain_left.n6 drain_left.t21 2.5005
R411 drain_left.n8 drain_left.t23 2.5005
R412 drain_left.n8 drain_left.t14 2.5005
R413 drain_left.n3 drain_left.t20 2.5005
R414 drain_left.n3 drain_left.t19 2.5005
R415 drain_left.n1 drain_left.t0 2.5005
R416 drain_left.n1 drain_left.t16 2.5005
R417 drain_left.n0 drain_left.t18 2.5005
R418 drain_left.n0 drain_left.t22 2.5005
R419 drain_left.n20 drain_left.t10 2.5005
R420 drain_left.n20 drain_left.t2 2.5005
R421 drain_left.n18 drain_left.t5 2.5005
R422 drain_left.n18 drain_left.t8 2.5005
R423 drain_left.n16 drain_left.t7 2.5005
R424 drain_left.n16 drain_left.t12 2.5005
R425 drain_left.n14 drain_left.t1 2.5005
R426 drain_left.n14 drain_left.t4 2.5005
R427 drain_left.n12 drain_left.t6 2.5005
R428 drain_left.n12 drain_left.t9 2.5005
R429 drain_left.n11 drain_left.t11 2.5005
R430 drain_left.n11 drain_left.t3 2.5005
R431 drain_left.n9 drain_left.n7 0.560845
R432 drain_left.n4 drain_left.n2 0.560845
R433 drain_left.n15 drain_left.n13 0.560845
R434 drain_left.n17 drain_left.n15 0.560845
R435 drain_left.n19 drain_left.n17 0.560845
R436 drain_left.n21 drain_left.n19 0.560845
R437 drain_left.n10 drain_left.n9 0.225326
R438 drain_left.n10 drain_left.n4 0.225326
C0 drain_left drain_right 1.29455f
C1 minus drain_left 0.171476f
C2 source drain_left 45.3833f
C3 minus drain_right 4.90476f
C4 source drain_right 45.384003f
C5 minus source 4.47084f
C6 plus drain_left 5.14254f
C7 plus drain_right 0.392113f
C8 minus plus 6.14151f
C9 source plus 4.48488f
C10 drain_right a_n2406_n3288# 6.8422f
C11 drain_left a_n2406_n3288# 7.1885f
C12 source a_n2406_n3288# 9.040753f
C13 minus a_n2406_n3288# 8.913962f
C14 plus a_n2406_n3288# 11.115701f
C15 drain_left.t18 a_n2406_n3288# 0.406351f
C16 drain_left.t22 a_n2406_n3288# 0.406351f
C17 drain_left.n0 a_n2406_n3288# 2.66608f
C18 drain_left.t0 a_n2406_n3288# 0.406351f
C19 drain_left.t16 a_n2406_n3288# 0.406351f
C20 drain_left.n1 a_n2406_n3288# 2.66281f
C21 drain_left.n2 a_n2406_n3288# 0.687096f
C22 drain_left.t20 a_n2406_n3288# 0.406351f
C23 drain_left.t19 a_n2406_n3288# 0.406351f
C24 drain_left.n3 a_n2406_n3288# 2.66281f
C25 drain_left.n4 a_n2406_n3288# 0.311828f
C26 drain_left.t13 a_n2406_n3288# 0.406351f
C27 drain_left.t15 a_n2406_n3288# 0.406351f
C28 drain_left.n5 a_n2406_n3288# 2.66608f
C29 drain_left.t17 a_n2406_n3288# 0.406351f
C30 drain_left.t21 a_n2406_n3288# 0.406351f
C31 drain_left.n6 a_n2406_n3288# 2.66281f
C32 drain_left.n7 a_n2406_n3288# 0.687096f
C33 drain_left.t23 a_n2406_n3288# 0.406351f
C34 drain_left.t14 a_n2406_n3288# 0.406351f
C35 drain_left.n8 a_n2406_n3288# 2.66281f
C36 drain_left.n9 a_n2406_n3288# 0.311828f
C37 drain_left.n10 a_n2406_n3288# 1.55107f
C38 drain_left.t11 a_n2406_n3288# 0.406351f
C39 drain_left.t3 a_n2406_n3288# 0.406351f
C40 drain_left.n11 a_n2406_n3288# 2.66609f
C41 drain_left.t6 a_n2406_n3288# 0.406351f
C42 drain_left.t9 a_n2406_n3288# 0.406351f
C43 drain_left.n12 a_n2406_n3288# 2.66282f
C44 drain_left.n13 a_n2406_n3288# 0.687077f
C45 drain_left.t1 a_n2406_n3288# 0.406351f
C46 drain_left.t4 a_n2406_n3288# 0.406351f
C47 drain_left.n14 a_n2406_n3288# 2.66282f
C48 drain_left.n15 a_n2406_n3288# 0.339478f
C49 drain_left.t7 a_n2406_n3288# 0.406351f
C50 drain_left.t12 a_n2406_n3288# 0.406351f
C51 drain_left.n16 a_n2406_n3288# 2.66282f
C52 drain_left.n17 a_n2406_n3288# 0.339478f
C53 drain_left.t5 a_n2406_n3288# 0.406351f
C54 drain_left.t8 a_n2406_n3288# 0.406351f
C55 drain_left.n18 a_n2406_n3288# 2.66282f
C56 drain_left.n19 a_n2406_n3288# 0.339478f
C57 drain_left.t10 a_n2406_n3288# 0.406351f
C58 drain_left.t2 a_n2406_n3288# 0.406351f
C59 drain_left.n20 a_n2406_n3288# 2.66281f
C60 drain_left.n21 a_n2406_n3288# 0.575673f
C61 plus.n0 a_n2406_n3288# 0.051974f
C62 plus.t13 a_n2406_n3288# 0.264367f
C63 plus.t15 a_n2406_n3288# 0.264367f
C64 plus.n1 a_n2406_n3288# 0.021247f
C65 plus.n2 a_n2406_n3288# 0.051974f
C66 plus.t11 a_n2406_n3288# 0.264367f
C67 plus.t16 a_n2406_n3288# 0.264367f
C68 plus.n3 a_n2406_n3288# 0.019645f
C69 plus.n4 a_n2406_n3288# 0.051974f
C70 plus.t22 a_n2406_n3288# 0.264367f
C71 plus.t14 a_n2406_n3288# 0.264367f
C72 plus.n5 a_n2406_n3288# 0.018043f
C73 plus.t12 a_n2406_n3288# 0.266803f
C74 plus.n6 a_n2406_n3288# 0.131768f
C75 plus.t20 a_n2406_n3288# 0.264367f
C76 plus.n7 a_n2406_n3288# 0.112884f
C77 plus.t17 a_n2406_n3288# 0.264367f
C78 plus.n8 a_n2406_n3288# 0.112884f
C79 plus.n9 a_n2406_n3288# 0.022048f
C80 plus.n10 a_n2406_n3288# 0.11349f
C81 plus.n11 a_n2406_n3288# 0.051974f
C82 plus.n12 a_n2406_n3288# 0.051974f
C83 plus.n13 a_n2406_n3288# 0.021247f
C84 plus.n14 a_n2406_n3288# 0.112884f
C85 plus.n15 a_n2406_n3288# 0.022048f
C86 plus.n16 a_n2406_n3288# 0.112884f
C87 plus.t19 a_n2406_n3288# 0.264367f
C88 plus.n17 a_n2406_n3288# 0.112884f
C89 plus.n18 a_n2406_n3288# 0.022048f
C90 plus.n19 a_n2406_n3288# 0.051974f
C91 plus.n20 a_n2406_n3288# 0.051974f
C92 plus.n21 a_n2406_n3288# 0.051974f
C93 plus.n22 a_n2406_n3288# 0.019645f
C94 plus.n23 a_n2406_n3288# 0.112884f
C95 plus.n24 a_n2406_n3288# 0.022048f
C96 plus.n25 a_n2406_n3288# 0.112884f
C97 plus.t18 a_n2406_n3288# 0.264367f
C98 plus.n26 a_n2406_n3288# 0.112884f
C99 plus.n27 a_n2406_n3288# 0.022048f
C100 plus.n28 a_n2406_n3288# 0.051974f
C101 plus.n29 a_n2406_n3288# 0.051974f
C102 plus.n30 a_n2406_n3288# 0.051974f
C103 plus.n31 a_n2406_n3288# 0.018043f
C104 plus.n32 a_n2406_n3288# 0.112884f
C105 plus.n33 a_n2406_n3288# 0.022048f
C106 plus.n34 a_n2406_n3288# 0.112884f
C107 plus.t21 a_n2406_n3288# 0.266803f
C108 plus.n35 a_n2406_n3288# 0.131696f
C109 plus.n36 a_n2406_n3288# 0.584401f
C110 plus.n37 a_n2406_n3288# 0.051974f
C111 plus.t5 a_n2406_n3288# 0.266803f
C112 plus.t1 a_n2406_n3288# 0.264367f
C113 plus.t23 a_n2406_n3288# 0.264367f
C114 plus.n38 a_n2406_n3288# 0.021247f
C115 plus.n39 a_n2406_n3288# 0.051974f
C116 plus.t7 a_n2406_n3288# 0.264367f
C117 plus.n40 a_n2406_n3288# 0.112884f
C118 plus.t3 a_n2406_n3288# 0.264367f
C119 plus.t4 a_n2406_n3288# 0.264367f
C120 plus.n41 a_n2406_n3288# 0.019645f
C121 plus.n42 a_n2406_n3288# 0.051974f
C122 plus.t0 a_n2406_n3288# 0.264367f
C123 plus.n43 a_n2406_n3288# 0.112884f
C124 plus.t9 a_n2406_n3288# 0.264367f
C125 plus.t6 a_n2406_n3288# 0.264367f
C126 plus.n44 a_n2406_n3288# 0.018043f
C127 plus.t8 a_n2406_n3288# 0.266803f
C128 plus.n45 a_n2406_n3288# 0.131768f
C129 plus.t2 a_n2406_n3288# 0.264367f
C130 plus.n46 a_n2406_n3288# 0.112884f
C131 plus.t10 a_n2406_n3288# 0.264367f
C132 plus.n47 a_n2406_n3288# 0.112884f
C133 plus.n48 a_n2406_n3288# 0.022048f
C134 plus.n49 a_n2406_n3288# 0.11349f
C135 plus.n50 a_n2406_n3288# 0.051974f
C136 plus.n51 a_n2406_n3288# 0.051974f
C137 plus.n52 a_n2406_n3288# 0.021247f
C138 plus.n53 a_n2406_n3288# 0.112884f
C139 plus.n54 a_n2406_n3288# 0.022048f
C140 plus.n55 a_n2406_n3288# 0.112884f
C141 plus.n56 a_n2406_n3288# 0.022048f
C142 plus.n57 a_n2406_n3288# 0.051974f
C143 plus.n58 a_n2406_n3288# 0.051974f
C144 plus.n59 a_n2406_n3288# 0.051974f
C145 plus.n60 a_n2406_n3288# 0.019645f
C146 plus.n61 a_n2406_n3288# 0.112884f
C147 plus.n62 a_n2406_n3288# 0.022048f
C148 plus.n63 a_n2406_n3288# 0.112884f
C149 plus.n64 a_n2406_n3288# 0.022048f
C150 plus.n65 a_n2406_n3288# 0.051974f
C151 plus.n66 a_n2406_n3288# 0.051974f
C152 plus.n67 a_n2406_n3288# 0.051974f
C153 plus.n68 a_n2406_n3288# 0.018043f
C154 plus.n69 a_n2406_n3288# 0.112884f
C155 plus.n70 a_n2406_n3288# 0.022048f
C156 plus.n71 a_n2406_n3288# 0.112884f
C157 plus.n72 a_n2406_n3288# 0.131696f
C158 plus.n73 a_n2406_n3288# 1.70189f
C159 drain_right.t22 a_n2406_n3288# 0.40563f
C160 drain_right.t15 a_n2406_n3288# 0.40563f
C161 drain_right.n0 a_n2406_n3288# 2.66135f
C162 drain_right.t5 a_n2406_n3288# 0.40563f
C163 drain_right.t0 a_n2406_n3288# 0.40563f
C164 drain_right.n1 a_n2406_n3288# 2.65809f
C165 drain_right.n2 a_n2406_n3288# 0.685878f
C166 drain_right.t20 a_n2406_n3288# 0.40563f
C167 drain_right.t13 a_n2406_n3288# 0.40563f
C168 drain_right.n3 a_n2406_n3288# 2.65809f
C169 drain_right.n4 a_n2406_n3288# 0.311275f
C170 drain_right.t1 a_n2406_n3288# 0.40563f
C171 drain_right.t21 a_n2406_n3288# 0.40563f
C172 drain_right.n5 a_n2406_n3288# 2.66135f
C173 drain_right.t19 a_n2406_n3288# 0.40563f
C174 drain_right.t11 a_n2406_n3288# 0.40563f
C175 drain_right.n6 a_n2406_n3288# 2.65809f
C176 drain_right.n7 a_n2406_n3288# 0.685878f
C177 drain_right.t3 a_n2406_n3288# 0.40563f
C178 drain_right.t23 a_n2406_n3288# 0.40563f
C179 drain_right.n8 a_n2406_n3288# 2.65809f
C180 drain_right.n9 a_n2406_n3288# 0.311275f
C181 drain_right.n10 a_n2406_n3288# 1.49033f
C182 drain_right.t18 a_n2406_n3288# 0.40563f
C183 drain_right.t17 a_n2406_n3288# 0.40563f
C184 drain_right.n11 a_n2406_n3288# 2.66135f
C185 drain_right.t14 a_n2406_n3288# 0.40563f
C186 drain_right.t10 a_n2406_n3288# 0.40563f
C187 drain_right.n12 a_n2406_n3288# 2.6581f
C188 drain_right.n13 a_n2406_n3288# 0.685868f
C189 drain_right.t6 a_n2406_n3288# 0.40563f
C190 drain_right.t16 a_n2406_n3288# 0.40563f
C191 drain_right.n14 a_n2406_n3288# 2.6581f
C192 drain_right.n15 a_n2406_n3288# 0.338876f
C193 drain_right.t8 a_n2406_n3288# 0.40563f
C194 drain_right.t9 a_n2406_n3288# 0.40563f
C195 drain_right.n16 a_n2406_n3288# 2.6581f
C196 drain_right.n17 a_n2406_n3288# 0.338876f
C197 drain_right.t2 a_n2406_n3288# 0.40563f
C198 drain_right.t12 a_n2406_n3288# 0.40563f
C199 drain_right.n18 a_n2406_n3288# 2.6581f
C200 drain_right.n19 a_n2406_n3288# 0.338876f
C201 drain_right.t7 a_n2406_n3288# 0.40563f
C202 drain_right.t4 a_n2406_n3288# 0.40563f
C203 drain_right.n20 a_n2406_n3288# 2.6581f
C204 drain_right.n21 a_n2406_n3288# 0.574642f
C205 source.t3 a_n2406_n3288# 2.82764f
C206 source.n0 a_n2406_n3288# 1.41012f
C207 source.t15 a_n2406_n3288# 0.365423f
C208 source.t8 a_n2406_n3288# 0.365423f
C209 source.n1 a_n2406_n3288# 2.31347f
C210 source.n2 a_n2406_n3288# 0.351867f
C211 source.t21 a_n2406_n3288# 0.365423f
C212 source.t18 a_n2406_n3288# 0.365423f
C213 source.n3 a_n2406_n3288# 2.31347f
C214 source.n4 a_n2406_n3288# 0.351867f
C215 source.t17 a_n2406_n3288# 0.365423f
C216 source.t20 a_n2406_n3288# 0.365423f
C217 source.n5 a_n2406_n3288# 2.31347f
C218 source.n6 a_n2406_n3288# 0.351867f
C219 source.t10 a_n2406_n3288# 0.365423f
C220 source.t7 a_n2406_n3288# 0.365423f
C221 source.n7 a_n2406_n3288# 2.31347f
C222 source.n8 a_n2406_n3288# 0.351867f
C223 source.t22 a_n2406_n3288# 0.365423f
C224 source.t11 a_n2406_n3288# 0.365423f
C225 source.n9 a_n2406_n3288# 2.31347f
C226 source.n10 a_n2406_n3288# 0.351867f
C227 source.t1 a_n2406_n3288# 2.82765f
C228 source.n11 a_n2406_n3288# 0.488025f
C229 source.t36 a_n2406_n3288# 2.82765f
C230 source.n12 a_n2406_n3288# 0.488025f
C231 source.t46 a_n2406_n3288# 0.365423f
C232 source.t29 a_n2406_n3288# 0.365423f
C233 source.n13 a_n2406_n3288# 2.31347f
C234 source.n14 a_n2406_n3288# 0.351867f
C235 source.t41 a_n2406_n3288# 0.365423f
C236 source.t38 a_n2406_n3288# 0.365423f
C237 source.n15 a_n2406_n3288# 2.31347f
C238 source.n16 a_n2406_n3288# 0.351867f
C239 source.t44 a_n2406_n3288# 0.365423f
C240 source.t39 a_n2406_n3288# 0.365423f
C241 source.n17 a_n2406_n3288# 2.31347f
C242 source.n18 a_n2406_n3288# 0.351867f
C243 source.t47 a_n2406_n3288# 0.365423f
C244 source.t32 a_n2406_n3288# 0.365423f
C245 source.n19 a_n2406_n3288# 2.31347f
C246 source.n20 a_n2406_n3288# 0.351867f
C247 source.t28 a_n2406_n3288# 0.365423f
C248 source.t40 a_n2406_n3288# 0.365423f
C249 source.n21 a_n2406_n3288# 2.31347f
C250 source.n22 a_n2406_n3288# 0.351867f
C251 source.t31 a_n2406_n3288# 2.82765f
C252 source.n23 a_n2406_n3288# 1.81054f
C253 source.t23 a_n2406_n3288# 2.82764f
C254 source.n24 a_n2406_n3288# 1.81055f
C255 source.t5 a_n2406_n3288# 0.365423f
C256 source.t2 a_n2406_n3288# 0.365423f
C257 source.n25 a_n2406_n3288# 2.31345f
C258 source.n26 a_n2406_n3288# 0.35188f
C259 source.t0 a_n2406_n3288# 0.365423f
C260 source.t6 a_n2406_n3288# 0.365423f
C261 source.n27 a_n2406_n3288# 2.31345f
C262 source.n28 a_n2406_n3288# 0.35188f
C263 source.t19 a_n2406_n3288# 0.365423f
C264 source.t12 a_n2406_n3288# 0.365423f
C265 source.n29 a_n2406_n3288# 2.31345f
C266 source.n30 a_n2406_n3288# 0.35188f
C267 source.t9 a_n2406_n3288# 0.365423f
C268 source.t13 a_n2406_n3288# 0.365423f
C269 source.n31 a_n2406_n3288# 2.31345f
C270 source.n32 a_n2406_n3288# 0.35188f
C271 source.t14 a_n2406_n3288# 0.365423f
C272 source.t16 a_n2406_n3288# 0.365423f
C273 source.n33 a_n2406_n3288# 2.31345f
C274 source.n34 a_n2406_n3288# 0.35188f
C275 source.t4 a_n2406_n3288# 2.82764f
C276 source.n35 a_n2406_n3288# 0.488037f
C277 source.t34 a_n2406_n3288# 2.82764f
C278 source.n36 a_n2406_n3288# 0.488037f
C279 source.t30 a_n2406_n3288# 0.365423f
C280 source.t27 a_n2406_n3288# 0.365423f
C281 source.n37 a_n2406_n3288# 2.31345f
C282 source.n38 a_n2406_n3288# 0.35188f
C283 source.t25 a_n2406_n3288# 0.365423f
C284 source.t45 a_n2406_n3288# 0.365423f
C285 source.n39 a_n2406_n3288# 2.31345f
C286 source.n40 a_n2406_n3288# 0.35188f
C287 source.t24 a_n2406_n3288# 0.365423f
C288 source.t42 a_n2406_n3288# 0.365423f
C289 source.n41 a_n2406_n3288# 2.31345f
C290 source.n42 a_n2406_n3288# 0.35188f
C291 source.t35 a_n2406_n3288# 0.365423f
C292 source.t26 a_n2406_n3288# 0.365423f
C293 source.n43 a_n2406_n3288# 2.31345f
C294 source.n44 a_n2406_n3288# 0.35188f
C295 source.t37 a_n2406_n3288# 0.365423f
C296 source.t43 a_n2406_n3288# 0.365423f
C297 source.n45 a_n2406_n3288# 2.31345f
C298 source.n46 a_n2406_n3288# 0.35188f
C299 source.t33 a_n2406_n3288# 2.82764f
C300 source.n47 a_n2406_n3288# 0.632737f
C301 source.n48 a_n2406_n3288# 1.59633f
C302 minus.n0 a_n2406_n3288# 0.050971f
C303 minus.t16 a_n2406_n3288# 0.261653f
C304 minus.t19 a_n2406_n3288# 0.259264f
C305 minus.t21 a_n2406_n3288# 0.259264f
C306 minus.n1 a_n2406_n3288# 0.020837f
C307 minus.n2 a_n2406_n3288# 0.050971f
C308 minus.t11 a_n2406_n3288# 0.259264f
C309 minus.n3 a_n2406_n3288# 0.110705f
C310 minus.t15 a_n2406_n3288# 0.259264f
C311 minus.t14 a_n2406_n3288# 0.259264f
C312 minus.n4 a_n2406_n3288# 0.019266f
C313 minus.n5 a_n2406_n3288# 0.050971f
C314 minus.t17 a_n2406_n3288# 0.259264f
C315 minus.n6 a_n2406_n3288# 0.110705f
C316 minus.t7 a_n2406_n3288# 0.259264f
C317 minus.t9 a_n2406_n3288# 0.259264f
C318 minus.n7 a_n2406_n3288# 0.017694f
C319 minus.t6 a_n2406_n3288# 0.261653f
C320 minus.n8 a_n2406_n3288# 0.129224f
C321 minus.t13 a_n2406_n3288# 0.259264f
C322 minus.n9 a_n2406_n3288# 0.110705f
C323 minus.t5 a_n2406_n3288# 0.259264f
C324 minus.n10 a_n2406_n3288# 0.110705f
C325 minus.n11 a_n2406_n3288# 0.021623f
C326 minus.n12 a_n2406_n3288# 0.111299f
C327 minus.n13 a_n2406_n3288# 0.050971f
C328 minus.n14 a_n2406_n3288# 0.050971f
C329 minus.n15 a_n2406_n3288# 0.020837f
C330 minus.n16 a_n2406_n3288# 0.110705f
C331 minus.n17 a_n2406_n3288# 0.021623f
C332 minus.n18 a_n2406_n3288# 0.110705f
C333 minus.n19 a_n2406_n3288# 0.021623f
C334 minus.n20 a_n2406_n3288# 0.050971f
C335 minus.n21 a_n2406_n3288# 0.050971f
C336 minus.n22 a_n2406_n3288# 0.050971f
C337 minus.n23 a_n2406_n3288# 0.019266f
C338 minus.n24 a_n2406_n3288# 0.110705f
C339 minus.n25 a_n2406_n3288# 0.021623f
C340 minus.n26 a_n2406_n3288# 0.110705f
C341 minus.n27 a_n2406_n3288# 0.021623f
C342 minus.n28 a_n2406_n3288# 0.050971f
C343 minus.n29 a_n2406_n3288# 0.050971f
C344 minus.n30 a_n2406_n3288# 0.050971f
C345 minus.n31 a_n2406_n3288# 0.017694f
C346 minus.n32 a_n2406_n3288# 0.110705f
C347 minus.n33 a_n2406_n3288# 0.021623f
C348 minus.n34 a_n2406_n3288# 0.110705f
C349 minus.n35 a_n2406_n3288# 0.129153f
C350 minus.n36 a_n2406_n3288# 1.96345f
C351 minus.n37 a_n2406_n3288# 0.050971f
C352 minus.t22 a_n2406_n3288# 0.259264f
C353 minus.t12 a_n2406_n3288# 0.259264f
C354 minus.n38 a_n2406_n3288# 0.020837f
C355 minus.n39 a_n2406_n3288# 0.050971f
C356 minus.t0 a_n2406_n3288# 0.259264f
C357 minus.t20 a_n2406_n3288# 0.259264f
C358 minus.n40 a_n2406_n3288# 0.019266f
C359 minus.n41 a_n2406_n3288# 0.050971f
C360 minus.t3 a_n2406_n3288# 0.259264f
C361 minus.t23 a_n2406_n3288# 0.259264f
C362 minus.n42 a_n2406_n3288# 0.017694f
C363 minus.t1 a_n2406_n3288# 0.261653f
C364 minus.n43 a_n2406_n3288# 0.129224f
C365 minus.t8 a_n2406_n3288# 0.259264f
C366 minus.n44 a_n2406_n3288# 0.110705f
C367 minus.t18 a_n2406_n3288# 0.259264f
C368 minus.n45 a_n2406_n3288# 0.110705f
C369 minus.n46 a_n2406_n3288# 0.021623f
C370 minus.n47 a_n2406_n3288# 0.111299f
C371 minus.n48 a_n2406_n3288# 0.050971f
C372 minus.n49 a_n2406_n3288# 0.050971f
C373 minus.n50 a_n2406_n3288# 0.020837f
C374 minus.n51 a_n2406_n3288# 0.110705f
C375 minus.n52 a_n2406_n3288# 0.021623f
C376 minus.n53 a_n2406_n3288# 0.110705f
C377 minus.t10 a_n2406_n3288# 0.259264f
C378 minus.n54 a_n2406_n3288# 0.110705f
C379 minus.n55 a_n2406_n3288# 0.021623f
C380 minus.n56 a_n2406_n3288# 0.050971f
C381 minus.n57 a_n2406_n3288# 0.050971f
C382 minus.n58 a_n2406_n3288# 0.050971f
C383 minus.n59 a_n2406_n3288# 0.019266f
C384 minus.n60 a_n2406_n3288# 0.110705f
C385 minus.n61 a_n2406_n3288# 0.021623f
C386 minus.n62 a_n2406_n3288# 0.110705f
C387 minus.t4 a_n2406_n3288# 0.259264f
C388 minus.n63 a_n2406_n3288# 0.110705f
C389 minus.n64 a_n2406_n3288# 0.021623f
C390 minus.n65 a_n2406_n3288# 0.050971f
C391 minus.n66 a_n2406_n3288# 0.050971f
C392 minus.n67 a_n2406_n3288# 0.050971f
C393 minus.n68 a_n2406_n3288# 0.017694f
C394 minus.n69 a_n2406_n3288# 0.110705f
C395 minus.n70 a_n2406_n3288# 0.021623f
C396 minus.n71 a_n2406_n3288# 0.110705f
C397 minus.t2 a_n2406_n3288# 0.261653f
C398 minus.n72 a_n2406_n3288# 0.129153f
C399 minus.n73 a_n2406_n3288# 0.336023f
C400 minus.n74 a_n2406_n3288# 2.36968f
.ends

