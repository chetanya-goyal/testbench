* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 drain_right.t13 minus.t0 source.t19 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X3 drain_right.t12 minus.t1 source.t15 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X4 drain_left.t13 plus.t0 source.t6 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X5 a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X6 drain_left.t12 plus.t1 source.t1 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X7 a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X8 drain_right.t11 minus.t2 source.t12 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X9 drain_right.t10 minus.t3 source.t22 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X10 drain_right.t9 minus.t4 source.t16 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X11 drain_left.t11 plus.t2 source.t2 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X12 drain_left.t10 plus.t3 source.t3 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X13 source.t13 minus.t5 drain_right.t8 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X14 drain_right.t7 minus.t6 source.t11 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X15 drain_right.t6 minus.t7 source.t17 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X16 source.t24 minus.t8 drain_right.t5 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X17 source.t23 minus.t9 drain_right.t4 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_right.t3 minus.t10 source.t14 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X19 drain_left.t9 plus.t4 source.t4 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X20 source.t5 plus.t5 drain_left.t8 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 source.t10 plus.t6 drain_left.t7 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 source.t20 minus.t11 drain_right.t2 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X23 source.t18 minus.t12 drain_right.t1 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X24 drain_left.t6 plus.t7 source.t0 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X25 drain_left.t5 plus.t8 source.t7 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X26 source.t27 plus.t9 drain_left.t4 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X27 source.t21 minus.t13 drain_right.t0 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X28 source.t26 plus.t10 drain_left.t3 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X29 drain_left.t2 plus.t11 source.t9 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X30 source.t8 plus.t12 drain_left.t1 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X31 source.t25 plus.t13 drain_left.t0 a_n2524_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n17 minus.n16 161.3
R1 minus.n15 minus.n0 161.3
R2 minus.n14 minus.n13 161.3
R3 minus.n12 minus.n1 161.3
R4 minus.n6 minus.n3 161.3
R5 minus.n35 minus.n34 161.3
R6 minus.n33 minus.n18 161.3
R7 minus.n32 minus.n31 161.3
R8 minus.n30 minus.n19 161.3
R9 minus.n24 minus.n21 161.3
R10 minus.n5 minus.t7 103.076
R11 minus.n23 minus.t3 103.076
R12 minus.n11 minus.n10 80.6037
R13 minus.n9 minus.n2 80.6037
R14 minus.n8 minus.n7 80.6037
R15 minus.n29 minus.n28 80.6037
R16 minus.n27 minus.n20 80.6037
R17 minus.n26 minus.n25 80.6037
R18 minus.n4 minus.t5 79.2293
R19 minus.n8 minus.t4 79.2293
R20 minus.n9 minus.t9 79.2293
R21 minus.n10 minus.t10 79.2293
R22 minus.n14 minus.t8 79.2293
R23 minus.n16 minus.t6 79.2293
R24 minus.n22 minus.t12 79.2293
R25 minus.n26 minus.t2 79.2293
R26 minus.n27 minus.t11 79.2293
R27 minus.n28 minus.t1 79.2293
R28 minus.n32 minus.t13 79.2293
R29 minus.n34 minus.t0 79.2293
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n6 minus.n5 44.9119
R35 minus.n24 minus.n23 44.9119
R36 minus.n16 minus.n15 35.055
R37 minus.n34 minus.n33 35.055
R38 minus.n8 minus.n3 32.1338
R39 minus.n10 minus.n1 32.1338
R40 minus.n26 minus.n21 32.1338
R41 minus.n28 minus.n19 32.1338
R42 minus.n36 minus.n17 30.5744
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n4 minus.n3 16.0672
R46 minus.n14 minus.n1 16.0672
R47 minus.n22 minus.n21 16.0672
R48 minus.n32 minus.n19 16.0672
R49 minus.n15 minus.n14 13.146
R50 minus.n33 minus.n32 13.146
R51 minus.n36 minus.n35 6.72588
R52 minus.n11 minus.n2 0.380177
R53 minus.n7 minus.n2 0.380177
R54 minus.n25 minus.n20 0.380177
R55 minus.n29 minus.n20 0.380177
R56 minus.n12 minus.n11 0.285035
R57 minus.n7 minus.n6 0.285035
R58 minus.n25 minus.n24 0.285035
R59 minus.n30 minus.n29 0.285035
R60 minus.n17 minus.n0 0.189894
R61 minus.n13 minus.n0 0.189894
R62 minus.n13 minus.n12 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 source.n0 source.t4 243.255
R68 source.n7 source.t17 243.255
R69 source.n27 source.t19 243.254
R70 source.n20 source.t2 243.254
R71 source.n2 source.n1 223.454
R72 source.n4 source.n3 223.454
R73 source.n6 source.n5 223.454
R74 source.n9 source.n8 223.454
R75 source.n11 source.n10 223.454
R76 source.n13 source.n12 223.454
R77 source.n26 source.n25 223.453
R78 source.n24 source.n23 223.453
R79 source.n22 source.n21 223.453
R80 source.n19 source.n18 223.453
R81 source.n17 source.n16 223.453
R82 source.n15 source.n14 223.453
R83 source.n25 source.t15 19.8005
R84 source.n25 source.t21 19.8005
R85 source.n23 source.t12 19.8005
R86 source.n23 source.t20 19.8005
R87 source.n21 source.t22 19.8005
R88 source.n21 source.t18 19.8005
R89 source.n18 source.t3 19.8005
R90 source.n18 source.t26 19.8005
R91 source.n16 source.t6 19.8005
R92 source.n16 source.t8 19.8005
R93 source.n14 source.t1 19.8005
R94 source.n14 source.t25 19.8005
R95 source.n1 source.t7 19.8005
R96 source.n1 source.t5 19.8005
R97 source.n3 source.t0 19.8005
R98 source.n3 source.t10 19.8005
R99 source.n5 source.t9 19.8005
R100 source.n5 source.t27 19.8005
R101 source.n8 source.t16 19.8005
R102 source.n8 source.t13 19.8005
R103 source.n10 source.t14 19.8005
R104 source.n10 source.t23 19.8005
R105 source.n12 source.t11 19.8005
R106 source.n12 source.t24 19.8005
R107 source.n15 source.n13 14.9027
R108 source.n28 source.n0 8.17853
R109 source.n28 source.n27 5.7505
R110 source.n13 source.n11 0.974638
R111 source.n11 source.n9 0.974638
R112 source.n9 source.n7 0.974638
R113 source.n6 source.n4 0.974638
R114 source.n4 source.n2 0.974638
R115 source.n2 source.n0 0.974638
R116 source.n17 source.n15 0.974638
R117 source.n19 source.n17 0.974638
R118 source.n20 source.n19 0.974638
R119 source.n24 source.n22 0.974638
R120 source.n26 source.n24 0.974638
R121 source.n27 source.n26 0.974638
R122 source.n7 source.n6 0.957397
R123 source.n22 source.n20 0.957397
R124 source source.n28 0.188
R125 drain_right.n1 drain_right.t10 260.906
R126 drain_right.n11 drain_right.t7 259.933
R127 drain_right.n8 drain_right.n6 241.107
R128 drain_right.n4 drain_right.n2 241.106
R129 drain_right.n8 drain_right.n7 240.132
R130 drain_right.n10 drain_right.n9 240.132
R131 drain_right.n4 drain_right.n3 240.131
R132 drain_right.n1 drain_right.n0 240.131
R133 drain_right drain_right.n5 24.0818
R134 drain_right.n2 drain_right.t0 19.8005
R135 drain_right.n2 drain_right.t13 19.8005
R136 drain_right.n3 drain_right.t2 19.8005
R137 drain_right.n3 drain_right.t12 19.8005
R138 drain_right.n0 drain_right.t1 19.8005
R139 drain_right.n0 drain_right.t11 19.8005
R140 drain_right.n6 drain_right.t8 19.8005
R141 drain_right.n6 drain_right.t6 19.8005
R142 drain_right.n7 drain_right.t4 19.8005
R143 drain_right.n7 drain_right.t9 19.8005
R144 drain_right.n9 drain_right.t5 19.8005
R145 drain_right.n9 drain_right.t3 19.8005
R146 drain_right drain_right.n11 6.14028
R147 drain_right.n11 drain_right.n10 0.974638
R148 drain_right.n10 drain_right.n8 0.974638
R149 drain_right.n5 drain_right.n1 0.675757
R150 drain_right.n5 drain_right.n4 0.188688
R151 plus.n7 plus.n6 161.3
R152 plus.n13 plus.n12 161.3
R153 plus.n14 plus.n1 161.3
R154 plus.n15 plus.n0 161.3
R155 plus.n17 plus.n16 161.3
R156 plus.n25 plus.n24 161.3
R157 plus.n31 plus.n30 161.3
R158 plus.n32 plus.n19 161.3
R159 plus.n33 plus.n18 161.3
R160 plus.n35 plus.n34 161.3
R161 plus.n5 plus.t11 103.076
R162 plus.n23 plus.t2 103.076
R163 plus.n8 plus.n3 80.6037
R164 plus.n10 plus.n9 80.6037
R165 plus.n11 plus.n2 80.6037
R166 plus.n26 plus.n21 80.6037
R167 plus.n28 plus.n27 80.6037
R168 plus.n29 plus.n20 80.6037
R169 plus.n16 plus.t4 79.2293
R170 plus.n14 plus.t5 79.2293
R171 plus.n2 plus.t8 79.2293
R172 plus.n9 plus.t6 79.2293
R173 plus.n8 plus.t7 79.2293
R174 plus.n4 plus.t9 79.2293
R175 plus.n34 plus.t1 79.2293
R176 plus.n32 plus.t13 79.2293
R177 plus.n20 plus.t0 79.2293
R178 plus.n27 plus.t12 79.2293
R179 plus.n26 plus.t3 79.2293
R180 plus.n22 plus.t10 79.2293
R181 plus.n9 plus.n2 48.2005
R182 plus.n9 plus.n8 48.2005
R183 plus.n27 plus.n20 48.2005
R184 plus.n27 plus.n26 48.2005
R185 plus.n24 plus.n23 44.9119
R186 plus.n6 plus.n5 44.9119
R187 plus.n16 plus.n15 35.055
R188 plus.n34 plus.n33 35.055
R189 plus.n13 plus.n2 32.1338
R190 plus.n8 plus.n7 32.1338
R191 plus.n31 plus.n20 32.1338
R192 plus.n26 plus.n25 32.1338
R193 plus plus.n35 28.6221
R194 plus.n23 plus.n22 17.739
R195 plus.n5 plus.n4 17.739
R196 plus.n14 plus.n13 16.0672
R197 plus.n7 plus.n4 16.0672
R198 plus.n32 plus.n31 16.0672
R199 plus.n25 plus.n22 16.0672
R200 plus.n15 plus.n14 13.146
R201 plus.n33 plus.n32 13.146
R202 plus plus.n17 8.20315
R203 plus.n10 plus.n3 0.380177
R204 plus.n11 plus.n10 0.380177
R205 plus.n29 plus.n28 0.380177
R206 plus.n28 plus.n21 0.380177
R207 plus.n6 plus.n3 0.285035
R208 plus.n12 plus.n11 0.285035
R209 plus.n30 plus.n29 0.285035
R210 plus.n24 plus.n21 0.285035
R211 plus.n12 plus.n1 0.189894
R212 plus.n1 plus.n0 0.189894
R213 plus.n17 plus.n0 0.189894
R214 plus.n35 plus.n18 0.189894
R215 plus.n19 plus.n18 0.189894
R216 plus.n30 plus.n19 0.189894
R217 drain_left.n7 drain_left.t2 260.906
R218 drain_left.n1 drain_left.t12 260.906
R219 drain_left.n4 drain_left.n2 241.106
R220 drain_left.n11 drain_left.n10 240.132
R221 drain_left.n9 drain_left.n8 240.132
R222 drain_left.n7 drain_left.n6 240.132
R223 drain_left.n4 drain_left.n3 240.131
R224 drain_left.n1 drain_left.n0 240.131
R225 drain_left drain_left.n5 24.635
R226 drain_left.n2 drain_left.t3 19.8005
R227 drain_left.n2 drain_left.t11 19.8005
R228 drain_left.n3 drain_left.t1 19.8005
R229 drain_left.n3 drain_left.t10 19.8005
R230 drain_left.n0 drain_left.t0 19.8005
R231 drain_left.n0 drain_left.t13 19.8005
R232 drain_left.n10 drain_left.t8 19.8005
R233 drain_left.n10 drain_left.t9 19.8005
R234 drain_left.n8 drain_left.t7 19.8005
R235 drain_left.n8 drain_left.t5 19.8005
R236 drain_left.n6 drain_left.t4 19.8005
R237 drain_left.n6 drain_left.t6 19.8005
R238 drain_left drain_left.n11 6.62735
R239 drain_left.n9 drain_left.n7 0.974638
R240 drain_left.n11 drain_left.n9 0.974638
R241 drain_left.n5 drain_left.n1 0.675757
R242 drain_left.n5 drain_left.n4 0.188688
C0 drain_right minus 1.31395f
C1 source drain_right 4.55394f
C2 drain_left drain_right 1.31379f
C3 source minus 2.00712f
C4 drain_left minus 0.181258f
C5 source drain_left 4.552721f
C6 drain_right plus 0.416062f
C7 plus minus 4.25911f
C8 source plus 2.02102f
C9 drain_left plus 1.56334f
C10 drain_right a_n2524_n1088# 4.28808f
C11 drain_left a_n2524_n1088# 4.61829f
C12 source a_n2524_n1088# 2.421517f
C13 minus a_n2524_n1088# 9.110234f
C14 plus a_n2524_n1088# 10.08821f
C15 drain_left.t12 a_n2524_n1088# 0.094968f
C16 drain_left.t0 a_n2524_n1088# 0.015227f
C17 drain_left.t13 a_n2524_n1088# 0.015227f
C18 drain_left.n0 a_n2524_n1088# 0.059168f
C19 drain_left.n1 a_n2524_n1088# 0.446549f
C20 drain_left.t3 a_n2524_n1088# 0.015227f
C21 drain_left.t11 a_n2524_n1088# 0.015227f
C22 drain_left.n2 a_n2524_n1088# 0.060233f
C23 drain_left.t1 a_n2524_n1088# 0.015227f
C24 drain_left.t10 a_n2524_n1088# 0.015227f
C25 drain_left.n3 a_n2524_n1088# 0.059168f
C26 drain_left.n4 a_n2524_n1088# 0.47171f
C27 drain_left.n5 a_n2524_n1088# 0.667385f
C28 drain_left.t2 a_n2524_n1088# 0.094968f
C29 drain_left.t4 a_n2524_n1088# 0.015227f
C30 drain_left.t6 a_n2524_n1088# 0.015227f
C31 drain_left.n6 a_n2524_n1088# 0.059168f
C32 drain_left.n7 a_n2524_n1088# 0.464444f
C33 drain_left.t7 a_n2524_n1088# 0.015227f
C34 drain_left.t5 a_n2524_n1088# 0.015227f
C35 drain_left.n8 a_n2524_n1088# 0.059168f
C36 drain_left.n9 a_n2524_n1088# 0.255719f
C37 drain_left.t8 a_n2524_n1088# 0.015227f
C38 drain_left.t9 a_n2524_n1088# 0.015227f
C39 drain_left.n10 a_n2524_n1088# 0.059168f
C40 drain_left.n11 a_n2524_n1088# 0.428505f
C41 plus.n0 a_n2524_n1088# 0.036941f
C42 plus.t4 a_n2524_n1088# 0.100214f
C43 plus.t5 a_n2524_n1088# 0.100214f
C44 plus.n1 a_n2524_n1088# 0.036941f
C45 plus.t8 a_n2524_n1088# 0.100214f
C46 plus.n2 a_n2524_n1088# 0.105088f
C47 plus.n3 a_n2524_n1088# 0.06153f
C48 plus.t6 a_n2524_n1088# 0.100214f
C49 plus.t7 a_n2524_n1088# 0.100214f
C50 plus.t9 a_n2524_n1088# 0.100214f
C51 plus.n4 a_n2524_n1088# 0.100825f
C52 plus.t11 a_n2524_n1088# 0.12302f
C53 plus.n5 a_n2524_n1088# 0.078968f
C54 plus.n6 a_n2524_n1088# 0.172521f
C55 plus.n7 a_n2524_n1088# 0.008383f
C56 plus.n8 a_n2524_n1088# 0.105088f
C57 plus.n9 a_n2524_n1088# 0.107593f
C58 plus.n10 a_n2524_n1088# 0.073883f
C59 plus.n11 a_n2524_n1088# 0.06153f
C60 plus.n12 a_n2524_n1088# 0.049294f
C61 plus.n13 a_n2524_n1088# 0.008383f
C62 plus.n14 a_n2524_n1088# 0.096249f
C63 plus.n15 a_n2524_n1088# 0.008383f
C64 plus.n16 a_n2524_n1088# 0.097161f
C65 plus.n17 a_n2524_n1088# 0.273788f
C66 plus.n18 a_n2524_n1088# 0.036941f
C67 plus.t1 a_n2524_n1088# 0.100214f
C68 plus.n19 a_n2524_n1088# 0.036941f
C69 plus.t13 a_n2524_n1088# 0.100214f
C70 plus.t0 a_n2524_n1088# 0.100214f
C71 plus.n20 a_n2524_n1088# 0.105088f
C72 plus.n21 a_n2524_n1088# 0.06153f
C73 plus.t12 a_n2524_n1088# 0.100214f
C74 plus.t3 a_n2524_n1088# 0.100214f
C75 plus.t10 a_n2524_n1088# 0.100214f
C76 plus.n22 a_n2524_n1088# 0.100825f
C77 plus.t2 a_n2524_n1088# 0.12302f
C78 plus.n23 a_n2524_n1088# 0.078968f
C79 plus.n24 a_n2524_n1088# 0.172521f
C80 plus.n25 a_n2524_n1088# 0.008383f
C81 plus.n26 a_n2524_n1088# 0.105088f
C82 plus.n27 a_n2524_n1088# 0.107593f
C83 plus.n28 a_n2524_n1088# 0.073883f
C84 plus.n29 a_n2524_n1088# 0.06153f
C85 plus.n30 a_n2524_n1088# 0.049294f
C86 plus.n31 a_n2524_n1088# 0.008383f
C87 plus.n32 a_n2524_n1088# 0.096249f
C88 plus.n33 a_n2524_n1088# 0.008383f
C89 plus.n34 a_n2524_n1088# 0.097161f
C90 plus.n35 a_n2524_n1088# 0.965158f
C91 drain_right.t10 a_n2524_n1088# 0.09655f
C92 drain_right.t1 a_n2524_n1088# 0.015481f
C93 drain_right.t11 a_n2524_n1088# 0.015481f
C94 drain_right.n0 a_n2524_n1088# 0.060154f
C95 drain_right.n1 a_n2524_n1088# 0.453988f
C96 drain_right.t0 a_n2524_n1088# 0.015481f
C97 drain_right.t13 a_n2524_n1088# 0.015481f
C98 drain_right.n2 a_n2524_n1088# 0.061236f
C99 drain_right.t2 a_n2524_n1088# 0.015481f
C100 drain_right.t12 a_n2524_n1088# 0.015481f
C101 drain_right.n3 a_n2524_n1088# 0.060154f
C102 drain_right.n4 a_n2524_n1088# 0.479569f
C103 drain_right.n5 a_n2524_n1088# 0.640811f
C104 drain_right.t8 a_n2524_n1088# 0.015481f
C105 drain_right.t6 a_n2524_n1088# 0.015481f
C106 drain_right.n6 a_n2524_n1088# 0.061236f
C107 drain_right.t4 a_n2524_n1088# 0.015481f
C108 drain_right.t9 a_n2524_n1088# 0.015481f
C109 drain_right.n7 a_n2524_n1088# 0.060154f
C110 drain_right.n8 a_n2524_n1088# 0.526767f
C111 drain_right.t5 a_n2524_n1088# 0.015481f
C112 drain_right.t3 a_n2524_n1088# 0.015481f
C113 drain_right.n9 a_n2524_n1088# 0.060154f
C114 drain_right.n10 a_n2524_n1088# 0.25998f
C115 drain_right.t7 a_n2524_n1088# 0.095755f
C116 drain_right.n11 a_n2524_n1088# 0.397146f
C117 source.t4 a_n2524_n1088# 0.169017f
C118 source.n0 a_n2524_n1088# 0.820963f
C119 source.t7 a_n2524_n1088# 0.030367f
C120 source.t5 a_n2524_n1088# 0.030367f
C121 source.n1 a_n2524_n1088# 0.098484f
C122 source.n2 a_n2524_n1088# 0.477251f
C123 source.t0 a_n2524_n1088# 0.030367f
C124 source.t10 a_n2524_n1088# 0.030367f
C125 source.n3 a_n2524_n1088# 0.098484f
C126 source.n4 a_n2524_n1088# 0.477251f
C127 source.t9 a_n2524_n1088# 0.030367f
C128 source.t27 a_n2524_n1088# 0.030367f
C129 source.n5 a_n2524_n1088# 0.098484f
C130 source.n6 a_n2524_n1088# 0.475116f
C131 source.t17 a_n2524_n1088# 0.169017f
C132 source.n7 a_n2524_n1088# 0.487402f
C133 source.t16 a_n2524_n1088# 0.030367f
C134 source.t13 a_n2524_n1088# 0.030367f
C135 source.n8 a_n2524_n1088# 0.098484f
C136 source.n9 a_n2524_n1088# 0.477251f
C137 source.t14 a_n2524_n1088# 0.030367f
C138 source.t23 a_n2524_n1088# 0.030367f
C139 source.n10 a_n2524_n1088# 0.098484f
C140 source.n11 a_n2524_n1088# 0.477251f
C141 source.t11 a_n2524_n1088# 0.030367f
C142 source.t24 a_n2524_n1088# 0.030367f
C143 source.n12 a_n2524_n1088# 0.098484f
C144 source.n13 a_n2524_n1088# 1.24873f
C145 source.t1 a_n2524_n1088# 0.030367f
C146 source.t25 a_n2524_n1088# 0.030367f
C147 source.n14 a_n2524_n1088# 0.098484f
C148 source.n15 a_n2524_n1088# 1.24873f
C149 source.t6 a_n2524_n1088# 0.030367f
C150 source.t8 a_n2524_n1088# 0.030367f
C151 source.n16 a_n2524_n1088# 0.098484f
C152 source.n17 a_n2524_n1088# 0.477251f
C153 source.t3 a_n2524_n1088# 0.030367f
C154 source.t26 a_n2524_n1088# 0.030367f
C155 source.n18 a_n2524_n1088# 0.098484f
C156 source.n19 a_n2524_n1088# 0.477251f
C157 source.t2 a_n2524_n1088# 0.169017f
C158 source.n20 a_n2524_n1088# 0.487402f
C159 source.t22 a_n2524_n1088# 0.030367f
C160 source.t18 a_n2524_n1088# 0.030367f
C161 source.n21 a_n2524_n1088# 0.098484f
C162 source.n22 a_n2524_n1088# 0.475116f
C163 source.t12 a_n2524_n1088# 0.030367f
C164 source.t20 a_n2524_n1088# 0.030367f
C165 source.n23 a_n2524_n1088# 0.098484f
C166 source.n24 a_n2524_n1088# 0.477251f
C167 source.t15 a_n2524_n1088# 0.030367f
C168 source.t21 a_n2524_n1088# 0.030367f
C169 source.n25 a_n2524_n1088# 0.098484f
C170 source.n26 a_n2524_n1088# 0.477251f
C171 source.t19 a_n2524_n1088# 0.169017f
C172 source.n27 a_n2524_n1088# 0.686076f
C173 source.n28 a_n2524_n1088# 0.801089f
C174 minus.n0 a_n2524_n1088# 0.036508f
C175 minus.n1 a_n2524_n1088# 0.008285f
C176 minus.t8 a_n2524_n1088# 0.09904f
C177 minus.n2 a_n2524_n1088# 0.073017f
C178 minus.n3 a_n2524_n1088# 0.008285f
C179 minus.t4 a_n2524_n1088# 0.09904f
C180 minus.t7 a_n2524_n1088# 0.121578f
C181 minus.t5 a_n2524_n1088# 0.09904f
C182 minus.n4 a_n2524_n1088# 0.099644f
C183 minus.n5 a_n2524_n1088# 0.078043f
C184 minus.n6 a_n2524_n1088# 0.170499f
C185 minus.n7 a_n2524_n1088# 0.060809f
C186 minus.n8 a_n2524_n1088# 0.103856f
C187 minus.t9 a_n2524_n1088# 0.09904f
C188 minus.n9 a_n2524_n1088# 0.106332f
C189 minus.t10 a_n2524_n1088# 0.09904f
C190 minus.n10 a_n2524_n1088# 0.103856f
C191 minus.n11 a_n2524_n1088# 0.060809f
C192 minus.n12 a_n2524_n1088# 0.048716f
C193 minus.n13 a_n2524_n1088# 0.036508f
C194 minus.n14 a_n2524_n1088# 0.095122f
C195 minus.n15 a_n2524_n1088# 0.008285f
C196 minus.t6 a_n2524_n1088# 0.09904f
C197 minus.n16 a_n2524_n1088# 0.096022f
C198 minus.n17 a_n2524_n1088# 0.988375f
C199 minus.n18 a_n2524_n1088# 0.036508f
C200 minus.n19 a_n2524_n1088# 0.008285f
C201 minus.n20 a_n2524_n1088# 0.073017f
C202 minus.n21 a_n2524_n1088# 0.008285f
C203 minus.t3 a_n2524_n1088# 0.121578f
C204 minus.t12 a_n2524_n1088# 0.09904f
C205 minus.n22 a_n2524_n1088# 0.099644f
C206 minus.n23 a_n2524_n1088# 0.078043f
C207 minus.n24 a_n2524_n1088# 0.170499f
C208 minus.n25 a_n2524_n1088# 0.060809f
C209 minus.t2 a_n2524_n1088# 0.09904f
C210 minus.n26 a_n2524_n1088# 0.103856f
C211 minus.t11 a_n2524_n1088# 0.09904f
C212 minus.n27 a_n2524_n1088# 0.106332f
C213 minus.t1 a_n2524_n1088# 0.09904f
C214 minus.n28 a_n2524_n1088# 0.103856f
C215 minus.n29 a_n2524_n1088# 0.060809f
C216 minus.n30 a_n2524_n1088# 0.048716f
C217 minus.n31 a_n2524_n1088# 0.036508f
C218 minus.t13 a_n2524_n1088# 0.09904f
C219 minus.n32 a_n2524_n1088# 0.095122f
C220 minus.n33 a_n2524_n1088# 0.008285f
C221 minus.t0 a_n2524_n1088# 0.09904f
C222 minus.n34 a_n2524_n1088# 0.096022f
C223 minus.n35 a_n2524_n1088# 0.257909f
C224 minus.n36 a_n2524_n1088# 1.20892f
.ends

