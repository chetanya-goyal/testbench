* NGSPICE file created from diffpair440.ext - technology: sky130A

.subckt diffpair440 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X1 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.5
X2 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X3 drain_left.t1 plus.t0 source.t1 a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X4 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X5 drain_right.t0 minus.t1 source.t3 a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X6 drain_left.t0 plus.t1 source.t0 a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X7 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
R0 minus.n0 minus.t0 851.375
R1 minus.n0 minus.t1 824.769
R2 minus minus.n0 0.188
R3 source.n258 source.n198 289.615
R4 source.n192 source.n132 289.615
R5 source.n60 source.n0 289.615
R6 source.n126 source.n66 289.615
R7 source.n218 source.n217 185
R8 source.n223 source.n222 185
R9 source.n225 source.n224 185
R10 source.n214 source.n213 185
R11 source.n231 source.n230 185
R12 source.n233 source.n232 185
R13 source.n210 source.n209 185
R14 source.n240 source.n239 185
R15 source.n241 source.n208 185
R16 source.n243 source.n242 185
R17 source.n206 source.n205 185
R18 source.n249 source.n248 185
R19 source.n251 source.n250 185
R20 source.n202 source.n201 185
R21 source.n257 source.n256 185
R22 source.n259 source.n258 185
R23 source.n152 source.n151 185
R24 source.n157 source.n156 185
R25 source.n159 source.n158 185
R26 source.n148 source.n147 185
R27 source.n165 source.n164 185
R28 source.n167 source.n166 185
R29 source.n144 source.n143 185
R30 source.n174 source.n173 185
R31 source.n175 source.n142 185
R32 source.n177 source.n176 185
R33 source.n140 source.n139 185
R34 source.n183 source.n182 185
R35 source.n185 source.n184 185
R36 source.n136 source.n135 185
R37 source.n191 source.n190 185
R38 source.n193 source.n192 185
R39 source.n61 source.n60 185
R40 source.n59 source.n58 185
R41 source.n4 source.n3 185
R42 source.n53 source.n52 185
R43 source.n51 source.n50 185
R44 source.n8 source.n7 185
R45 source.n45 source.n44 185
R46 source.n43 source.n10 185
R47 source.n42 source.n41 185
R48 source.n13 source.n11 185
R49 source.n36 source.n35 185
R50 source.n34 source.n33 185
R51 source.n17 source.n16 185
R52 source.n28 source.n27 185
R53 source.n26 source.n25 185
R54 source.n21 source.n20 185
R55 source.n127 source.n126 185
R56 source.n125 source.n124 185
R57 source.n70 source.n69 185
R58 source.n119 source.n118 185
R59 source.n117 source.n116 185
R60 source.n74 source.n73 185
R61 source.n111 source.n110 185
R62 source.n109 source.n76 185
R63 source.n108 source.n107 185
R64 source.n79 source.n77 185
R65 source.n102 source.n101 185
R66 source.n100 source.n99 185
R67 source.n83 source.n82 185
R68 source.n94 source.n93 185
R69 source.n92 source.n91 185
R70 source.n87 source.n86 185
R71 source.n219 source.t3 149.524
R72 source.n153 source.t1 149.524
R73 source.n22 source.t0 149.524
R74 source.n88 source.t2 149.524
R75 source.n223 source.n217 104.615
R76 source.n224 source.n223 104.615
R77 source.n224 source.n213 104.615
R78 source.n231 source.n213 104.615
R79 source.n232 source.n231 104.615
R80 source.n232 source.n209 104.615
R81 source.n240 source.n209 104.615
R82 source.n241 source.n240 104.615
R83 source.n242 source.n241 104.615
R84 source.n242 source.n205 104.615
R85 source.n249 source.n205 104.615
R86 source.n250 source.n249 104.615
R87 source.n250 source.n201 104.615
R88 source.n257 source.n201 104.615
R89 source.n258 source.n257 104.615
R90 source.n157 source.n151 104.615
R91 source.n158 source.n157 104.615
R92 source.n158 source.n147 104.615
R93 source.n165 source.n147 104.615
R94 source.n166 source.n165 104.615
R95 source.n166 source.n143 104.615
R96 source.n174 source.n143 104.615
R97 source.n175 source.n174 104.615
R98 source.n176 source.n175 104.615
R99 source.n176 source.n139 104.615
R100 source.n183 source.n139 104.615
R101 source.n184 source.n183 104.615
R102 source.n184 source.n135 104.615
R103 source.n191 source.n135 104.615
R104 source.n192 source.n191 104.615
R105 source.n60 source.n59 104.615
R106 source.n59 source.n3 104.615
R107 source.n52 source.n3 104.615
R108 source.n52 source.n51 104.615
R109 source.n51 source.n7 104.615
R110 source.n44 source.n7 104.615
R111 source.n44 source.n43 104.615
R112 source.n43 source.n42 104.615
R113 source.n42 source.n11 104.615
R114 source.n35 source.n11 104.615
R115 source.n35 source.n34 104.615
R116 source.n34 source.n16 104.615
R117 source.n27 source.n16 104.615
R118 source.n27 source.n26 104.615
R119 source.n26 source.n20 104.615
R120 source.n126 source.n125 104.615
R121 source.n125 source.n69 104.615
R122 source.n118 source.n69 104.615
R123 source.n118 source.n117 104.615
R124 source.n117 source.n73 104.615
R125 source.n110 source.n73 104.615
R126 source.n110 source.n109 104.615
R127 source.n109 source.n108 104.615
R128 source.n108 source.n77 104.615
R129 source.n101 source.n77 104.615
R130 source.n101 source.n100 104.615
R131 source.n100 source.n82 104.615
R132 source.n93 source.n82 104.615
R133 source.n93 source.n92 104.615
R134 source.n92 source.n86 104.615
R135 source.t3 source.n217 52.3082
R136 source.t1 source.n151 52.3082
R137 source.t0 source.n20 52.3082
R138 source.t2 source.n86 52.3082
R139 source.n263 source.n262 29.8581
R140 source.n197 source.n196 29.8581
R141 source.n65 source.n64 29.8581
R142 source.n131 source.n130 29.8581
R143 source.n197 source.n131 22.7339
R144 source.n264 source.n65 16.3977
R145 source.n243 source.n208 13.1884
R146 source.n177 source.n142 13.1884
R147 source.n45 source.n10 13.1884
R148 source.n111 source.n76 13.1884
R149 source.n239 source.n238 12.8005
R150 source.n244 source.n206 12.8005
R151 source.n173 source.n172 12.8005
R152 source.n178 source.n140 12.8005
R153 source.n46 source.n8 12.8005
R154 source.n41 source.n12 12.8005
R155 source.n112 source.n74 12.8005
R156 source.n107 source.n78 12.8005
R157 source.n237 source.n210 12.0247
R158 source.n248 source.n247 12.0247
R159 source.n171 source.n144 12.0247
R160 source.n182 source.n181 12.0247
R161 source.n50 source.n49 12.0247
R162 source.n40 source.n13 12.0247
R163 source.n116 source.n115 12.0247
R164 source.n106 source.n79 12.0247
R165 source.n234 source.n233 11.249
R166 source.n251 source.n204 11.249
R167 source.n168 source.n167 11.249
R168 source.n185 source.n138 11.249
R169 source.n53 source.n6 11.249
R170 source.n37 source.n36 11.249
R171 source.n119 source.n72 11.249
R172 source.n103 source.n102 11.249
R173 source.n230 source.n212 10.4732
R174 source.n252 source.n202 10.4732
R175 source.n164 source.n146 10.4732
R176 source.n186 source.n136 10.4732
R177 source.n54 source.n4 10.4732
R178 source.n33 source.n15 10.4732
R179 source.n120 source.n70 10.4732
R180 source.n99 source.n81 10.4732
R181 source.n219 source.n218 10.2747
R182 source.n153 source.n152 10.2747
R183 source.n22 source.n21 10.2747
R184 source.n88 source.n87 10.2747
R185 source.n229 source.n214 9.69747
R186 source.n256 source.n255 9.69747
R187 source.n163 source.n148 9.69747
R188 source.n190 source.n189 9.69747
R189 source.n58 source.n57 9.69747
R190 source.n32 source.n17 9.69747
R191 source.n124 source.n123 9.69747
R192 source.n98 source.n83 9.69747
R193 source.n262 source.n261 9.45567
R194 source.n196 source.n195 9.45567
R195 source.n64 source.n63 9.45567
R196 source.n130 source.n129 9.45567
R197 source.n261 source.n260 9.3005
R198 source.n200 source.n199 9.3005
R199 source.n255 source.n254 9.3005
R200 source.n253 source.n252 9.3005
R201 source.n204 source.n203 9.3005
R202 source.n247 source.n246 9.3005
R203 source.n245 source.n244 9.3005
R204 source.n221 source.n220 9.3005
R205 source.n216 source.n215 9.3005
R206 source.n227 source.n226 9.3005
R207 source.n229 source.n228 9.3005
R208 source.n212 source.n211 9.3005
R209 source.n235 source.n234 9.3005
R210 source.n237 source.n236 9.3005
R211 source.n238 source.n207 9.3005
R212 source.n195 source.n194 9.3005
R213 source.n134 source.n133 9.3005
R214 source.n189 source.n188 9.3005
R215 source.n187 source.n186 9.3005
R216 source.n138 source.n137 9.3005
R217 source.n181 source.n180 9.3005
R218 source.n179 source.n178 9.3005
R219 source.n155 source.n154 9.3005
R220 source.n150 source.n149 9.3005
R221 source.n161 source.n160 9.3005
R222 source.n163 source.n162 9.3005
R223 source.n146 source.n145 9.3005
R224 source.n169 source.n168 9.3005
R225 source.n171 source.n170 9.3005
R226 source.n172 source.n141 9.3005
R227 source.n24 source.n23 9.3005
R228 source.n19 source.n18 9.3005
R229 source.n30 source.n29 9.3005
R230 source.n32 source.n31 9.3005
R231 source.n15 source.n14 9.3005
R232 source.n38 source.n37 9.3005
R233 source.n40 source.n39 9.3005
R234 source.n12 source.n9 9.3005
R235 source.n63 source.n62 9.3005
R236 source.n2 source.n1 9.3005
R237 source.n57 source.n56 9.3005
R238 source.n55 source.n54 9.3005
R239 source.n6 source.n5 9.3005
R240 source.n49 source.n48 9.3005
R241 source.n47 source.n46 9.3005
R242 source.n90 source.n89 9.3005
R243 source.n85 source.n84 9.3005
R244 source.n96 source.n95 9.3005
R245 source.n98 source.n97 9.3005
R246 source.n81 source.n80 9.3005
R247 source.n104 source.n103 9.3005
R248 source.n106 source.n105 9.3005
R249 source.n78 source.n75 9.3005
R250 source.n129 source.n128 9.3005
R251 source.n68 source.n67 9.3005
R252 source.n123 source.n122 9.3005
R253 source.n121 source.n120 9.3005
R254 source.n72 source.n71 9.3005
R255 source.n115 source.n114 9.3005
R256 source.n113 source.n112 9.3005
R257 source.n226 source.n225 8.92171
R258 source.n259 source.n200 8.92171
R259 source.n160 source.n159 8.92171
R260 source.n193 source.n134 8.92171
R261 source.n61 source.n2 8.92171
R262 source.n29 source.n28 8.92171
R263 source.n127 source.n68 8.92171
R264 source.n95 source.n94 8.92171
R265 source.n222 source.n216 8.14595
R266 source.n260 source.n198 8.14595
R267 source.n156 source.n150 8.14595
R268 source.n194 source.n132 8.14595
R269 source.n62 source.n0 8.14595
R270 source.n25 source.n19 8.14595
R271 source.n128 source.n66 8.14595
R272 source.n91 source.n85 8.14595
R273 source.n221 source.n218 7.3702
R274 source.n155 source.n152 7.3702
R275 source.n24 source.n21 7.3702
R276 source.n90 source.n87 7.3702
R277 source.n222 source.n221 5.81868
R278 source.n262 source.n198 5.81868
R279 source.n156 source.n155 5.81868
R280 source.n196 source.n132 5.81868
R281 source.n64 source.n0 5.81868
R282 source.n25 source.n24 5.81868
R283 source.n130 source.n66 5.81868
R284 source.n91 source.n90 5.81868
R285 source.n264 source.n263 5.62119
R286 source.n225 source.n216 5.04292
R287 source.n260 source.n259 5.04292
R288 source.n159 source.n150 5.04292
R289 source.n194 source.n193 5.04292
R290 source.n62 source.n61 5.04292
R291 source.n28 source.n19 5.04292
R292 source.n128 source.n127 5.04292
R293 source.n94 source.n85 5.04292
R294 source.n226 source.n214 4.26717
R295 source.n256 source.n200 4.26717
R296 source.n160 source.n148 4.26717
R297 source.n190 source.n134 4.26717
R298 source.n58 source.n2 4.26717
R299 source.n29 source.n17 4.26717
R300 source.n124 source.n68 4.26717
R301 source.n95 source.n83 4.26717
R302 source.n230 source.n229 3.49141
R303 source.n255 source.n202 3.49141
R304 source.n164 source.n163 3.49141
R305 source.n189 source.n136 3.49141
R306 source.n57 source.n4 3.49141
R307 source.n33 source.n32 3.49141
R308 source.n123 source.n70 3.49141
R309 source.n99 source.n98 3.49141
R310 source.n220 source.n219 2.84303
R311 source.n154 source.n153 2.84303
R312 source.n23 source.n22 2.84303
R313 source.n89 source.n88 2.84303
R314 source.n233 source.n212 2.71565
R315 source.n252 source.n251 2.71565
R316 source.n167 source.n146 2.71565
R317 source.n186 source.n185 2.71565
R318 source.n54 source.n53 2.71565
R319 source.n36 source.n15 2.71565
R320 source.n120 source.n119 2.71565
R321 source.n102 source.n81 2.71565
R322 source.n234 source.n210 1.93989
R323 source.n248 source.n204 1.93989
R324 source.n168 source.n144 1.93989
R325 source.n182 source.n138 1.93989
R326 source.n50 source.n6 1.93989
R327 source.n37 source.n13 1.93989
R328 source.n116 source.n72 1.93989
R329 source.n103 source.n79 1.93989
R330 source.n239 source.n237 1.16414
R331 source.n247 source.n206 1.16414
R332 source.n173 source.n171 1.16414
R333 source.n181 source.n140 1.16414
R334 source.n49 source.n8 1.16414
R335 source.n41 source.n40 1.16414
R336 source.n115 source.n74 1.16414
R337 source.n107 source.n106 1.16414
R338 source.n131 source.n65 0.828086
R339 source.n263 source.n197 0.828086
R340 source.n238 source.n208 0.388379
R341 source.n244 source.n243 0.388379
R342 source.n172 source.n142 0.388379
R343 source.n178 source.n177 0.388379
R344 source.n46 source.n45 0.388379
R345 source.n12 source.n10 0.388379
R346 source.n112 source.n111 0.388379
R347 source.n78 source.n76 0.388379
R348 source source.n264 0.188
R349 source.n220 source.n215 0.155672
R350 source.n227 source.n215 0.155672
R351 source.n228 source.n227 0.155672
R352 source.n228 source.n211 0.155672
R353 source.n235 source.n211 0.155672
R354 source.n236 source.n235 0.155672
R355 source.n236 source.n207 0.155672
R356 source.n245 source.n207 0.155672
R357 source.n246 source.n245 0.155672
R358 source.n246 source.n203 0.155672
R359 source.n253 source.n203 0.155672
R360 source.n254 source.n253 0.155672
R361 source.n254 source.n199 0.155672
R362 source.n261 source.n199 0.155672
R363 source.n154 source.n149 0.155672
R364 source.n161 source.n149 0.155672
R365 source.n162 source.n161 0.155672
R366 source.n162 source.n145 0.155672
R367 source.n169 source.n145 0.155672
R368 source.n170 source.n169 0.155672
R369 source.n170 source.n141 0.155672
R370 source.n179 source.n141 0.155672
R371 source.n180 source.n179 0.155672
R372 source.n180 source.n137 0.155672
R373 source.n187 source.n137 0.155672
R374 source.n188 source.n187 0.155672
R375 source.n188 source.n133 0.155672
R376 source.n195 source.n133 0.155672
R377 source.n63 source.n1 0.155672
R378 source.n56 source.n1 0.155672
R379 source.n56 source.n55 0.155672
R380 source.n55 source.n5 0.155672
R381 source.n48 source.n5 0.155672
R382 source.n48 source.n47 0.155672
R383 source.n47 source.n9 0.155672
R384 source.n39 source.n9 0.155672
R385 source.n39 source.n38 0.155672
R386 source.n38 source.n14 0.155672
R387 source.n31 source.n14 0.155672
R388 source.n31 source.n30 0.155672
R389 source.n30 source.n18 0.155672
R390 source.n23 source.n18 0.155672
R391 source.n129 source.n67 0.155672
R392 source.n122 source.n67 0.155672
R393 source.n122 source.n121 0.155672
R394 source.n121 source.n71 0.155672
R395 source.n114 source.n71 0.155672
R396 source.n114 source.n113 0.155672
R397 source.n113 source.n75 0.155672
R398 source.n105 source.n75 0.155672
R399 source.n105 source.n104 0.155672
R400 source.n104 source.n80 0.155672
R401 source.n97 source.n80 0.155672
R402 source.n97 source.n96 0.155672
R403 source.n96 source.n84 0.155672
R404 source.n89 source.n84 0.155672
R405 drain_right.n60 drain_right.n0 289.615
R406 drain_right.n125 drain_right.n65 289.615
R407 drain_right.n20 drain_right.n19 185
R408 drain_right.n25 drain_right.n24 185
R409 drain_right.n27 drain_right.n26 185
R410 drain_right.n16 drain_right.n15 185
R411 drain_right.n33 drain_right.n32 185
R412 drain_right.n35 drain_right.n34 185
R413 drain_right.n12 drain_right.n11 185
R414 drain_right.n42 drain_right.n41 185
R415 drain_right.n43 drain_right.n10 185
R416 drain_right.n45 drain_right.n44 185
R417 drain_right.n8 drain_right.n7 185
R418 drain_right.n51 drain_right.n50 185
R419 drain_right.n53 drain_right.n52 185
R420 drain_right.n4 drain_right.n3 185
R421 drain_right.n59 drain_right.n58 185
R422 drain_right.n61 drain_right.n60 185
R423 drain_right.n126 drain_right.n125 185
R424 drain_right.n124 drain_right.n123 185
R425 drain_right.n69 drain_right.n68 185
R426 drain_right.n118 drain_right.n117 185
R427 drain_right.n116 drain_right.n115 185
R428 drain_right.n73 drain_right.n72 185
R429 drain_right.n110 drain_right.n109 185
R430 drain_right.n108 drain_right.n75 185
R431 drain_right.n107 drain_right.n106 185
R432 drain_right.n78 drain_right.n76 185
R433 drain_right.n101 drain_right.n100 185
R434 drain_right.n99 drain_right.n98 185
R435 drain_right.n82 drain_right.n81 185
R436 drain_right.n93 drain_right.n92 185
R437 drain_right.n91 drain_right.n90 185
R438 drain_right.n86 drain_right.n85 185
R439 drain_right.n21 drain_right.t0 149.524
R440 drain_right.n87 drain_right.t1 149.524
R441 drain_right.n25 drain_right.n19 104.615
R442 drain_right.n26 drain_right.n25 104.615
R443 drain_right.n26 drain_right.n15 104.615
R444 drain_right.n33 drain_right.n15 104.615
R445 drain_right.n34 drain_right.n33 104.615
R446 drain_right.n34 drain_right.n11 104.615
R447 drain_right.n42 drain_right.n11 104.615
R448 drain_right.n43 drain_right.n42 104.615
R449 drain_right.n44 drain_right.n43 104.615
R450 drain_right.n44 drain_right.n7 104.615
R451 drain_right.n51 drain_right.n7 104.615
R452 drain_right.n52 drain_right.n51 104.615
R453 drain_right.n52 drain_right.n3 104.615
R454 drain_right.n59 drain_right.n3 104.615
R455 drain_right.n60 drain_right.n59 104.615
R456 drain_right.n125 drain_right.n124 104.615
R457 drain_right.n124 drain_right.n68 104.615
R458 drain_right.n117 drain_right.n68 104.615
R459 drain_right.n117 drain_right.n116 104.615
R460 drain_right.n116 drain_right.n72 104.615
R461 drain_right.n109 drain_right.n72 104.615
R462 drain_right.n109 drain_right.n108 104.615
R463 drain_right.n108 drain_right.n107 104.615
R464 drain_right.n107 drain_right.n76 104.615
R465 drain_right.n100 drain_right.n76 104.615
R466 drain_right.n100 drain_right.n99 104.615
R467 drain_right.n99 drain_right.n81 104.615
R468 drain_right.n92 drain_right.n81 104.615
R469 drain_right.n92 drain_right.n91 104.615
R470 drain_right.n91 drain_right.n85 104.615
R471 drain_right drain_right.n64 74.3833
R472 drain_right drain_right.n129 52.5473
R473 drain_right.t0 drain_right.n19 52.3082
R474 drain_right.t1 drain_right.n85 52.3082
R475 drain_right.n45 drain_right.n10 13.1884
R476 drain_right.n110 drain_right.n75 13.1884
R477 drain_right.n41 drain_right.n40 12.8005
R478 drain_right.n46 drain_right.n8 12.8005
R479 drain_right.n111 drain_right.n73 12.8005
R480 drain_right.n106 drain_right.n77 12.8005
R481 drain_right.n39 drain_right.n12 12.0247
R482 drain_right.n50 drain_right.n49 12.0247
R483 drain_right.n115 drain_right.n114 12.0247
R484 drain_right.n105 drain_right.n78 12.0247
R485 drain_right.n36 drain_right.n35 11.249
R486 drain_right.n53 drain_right.n6 11.249
R487 drain_right.n118 drain_right.n71 11.249
R488 drain_right.n102 drain_right.n101 11.249
R489 drain_right.n32 drain_right.n14 10.4732
R490 drain_right.n54 drain_right.n4 10.4732
R491 drain_right.n119 drain_right.n69 10.4732
R492 drain_right.n98 drain_right.n80 10.4732
R493 drain_right.n21 drain_right.n20 10.2747
R494 drain_right.n87 drain_right.n86 10.2747
R495 drain_right.n31 drain_right.n16 9.69747
R496 drain_right.n58 drain_right.n57 9.69747
R497 drain_right.n123 drain_right.n122 9.69747
R498 drain_right.n97 drain_right.n82 9.69747
R499 drain_right.n64 drain_right.n63 9.45567
R500 drain_right.n129 drain_right.n128 9.45567
R501 drain_right.n63 drain_right.n62 9.3005
R502 drain_right.n2 drain_right.n1 9.3005
R503 drain_right.n57 drain_right.n56 9.3005
R504 drain_right.n55 drain_right.n54 9.3005
R505 drain_right.n6 drain_right.n5 9.3005
R506 drain_right.n49 drain_right.n48 9.3005
R507 drain_right.n47 drain_right.n46 9.3005
R508 drain_right.n23 drain_right.n22 9.3005
R509 drain_right.n18 drain_right.n17 9.3005
R510 drain_right.n29 drain_right.n28 9.3005
R511 drain_right.n31 drain_right.n30 9.3005
R512 drain_right.n14 drain_right.n13 9.3005
R513 drain_right.n37 drain_right.n36 9.3005
R514 drain_right.n39 drain_right.n38 9.3005
R515 drain_right.n40 drain_right.n9 9.3005
R516 drain_right.n89 drain_right.n88 9.3005
R517 drain_right.n84 drain_right.n83 9.3005
R518 drain_right.n95 drain_right.n94 9.3005
R519 drain_right.n97 drain_right.n96 9.3005
R520 drain_right.n80 drain_right.n79 9.3005
R521 drain_right.n103 drain_right.n102 9.3005
R522 drain_right.n105 drain_right.n104 9.3005
R523 drain_right.n77 drain_right.n74 9.3005
R524 drain_right.n128 drain_right.n127 9.3005
R525 drain_right.n67 drain_right.n66 9.3005
R526 drain_right.n122 drain_right.n121 9.3005
R527 drain_right.n120 drain_right.n119 9.3005
R528 drain_right.n71 drain_right.n70 9.3005
R529 drain_right.n114 drain_right.n113 9.3005
R530 drain_right.n112 drain_right.n111 9.3005
R531 drain_right.n28 drain_right.n27 8.92171
R532 drain_right.n61 drain_right.n2 8.92171
R533 drain_right.n126 drain_right.n67 8.92171
R534 drain_right.n94 drain_right.n93 8.92171
R535 drain_right.n24 drain_right.n18 8.14595
R536 drain_right.n62 drain_right.n0 8.14595
R537 drain_right.n127 drain_right.n65 8.14595
R538 drain_right.n90 drain_right.n84 8.14595
R539 drain_right.n23 drain_right.n20 7.3702
R540 drain_right.n89 drain_right.n86 7.3702
R541 drain_right.n24 drain_right.n23 5.81868
R542 drain_right.n64 drain_right.n0 5.81868
R543 drain_right.n129 drain_right.n65 5.81868
R544 drain_right.n90 drain_right.n89 5.81868
R545 drain_right.n27 drain_right.n18 5.04292
R546 drain_right.n62 drain_right.n61 5.04292
R547 drain_right.n127 drain_right.n126 5.04292
R548 drain_right.n93 drain_right.n84 5.04292
R549 drain_right.n28 drain_right.n16 4.26717
R550 drain_right.n58 drain_right.n2 4.26717
R551 drain_right.n123 drain_right.n67 4.26717
R552 drain_right.n94 drain_right.n82 4.26717
R553 drain_right.n32 drain_right.n31 3.49141
R554 drain_right.n57 drain_right.n4 3.49141
R555 drain_right.n122 drain_right.n69 3.49141
R556 drain_right.n98 drain_right.n97 3.49141
R557 drain_right.n22 drain_right.n21 2.84303
R558 drain_right.n88 drain_right.n87 2.84303
R559 drain_right.n35 drain_right.n14 2.71565
R560 drain_right.n54 drain_right.n53 2.71565
R561 drain_right.n119 drain_right.n118 2.71565
R562 drain_right.n101 drain_right.n80 2.71565
R563 drain_right.n36 drain_right.n12 1.93989
R564 drain_right.n50 drain_right.n6 1.93989
R565 drain_right.n115 drain_right.n71 1.93989
R566 drain_right.n102 drain_right.n78 1.93989
R567 drain_right.n41 drain_right.n39 1.16414
R568 drain_right.n49 drain_right.n8 1.16414
R569 drain_right.n114 drain_right.n73 1.16414
R570 drain_right.n106 drain_right.n105 1.16414
R571 drain_right.n40 drain_right.n10 0.388379
R572 drain_right.n46 drain_right.n45 0.388379
R573 drain_right.n111 drain_right.n110 0.388379
R574 drain_right.n77 drain_right.n75 0.388379
R575 drain_right.n22 drain_right.n17 0.155672
R576 drain_right.n29 drain_right.n17 0.155672
R577 drain_right.n30 drain_right.n29 0.155672
R578 drain_right.n30 drain_right.n13 0.155672
R579 drain_right.n37 drain_right.n13 0.155672
R580 drain_right.n38 drain_right.n37 0.155672
R581 drain_right.n38 drain_right.n9 0.155672
R582 drain_right.n47 drain_right.n9 0.155672
R583 drain_right.n48 drain_right.n47 0.155672
R584 drain_right.n48 drain_right.n5 0.155672
R585 drain_right.n55 drain_right.n5 0.155672
R586 drain_right.n56 drain_right.n55 0.155672
R587 drain_right.n56 drain_right.n1 0.155672
R588 drain_right.n63 drain_right.n1 0.155672
R589 drain_right.n128 drain_right.n66 0.155672
R590 drain_right.n121 drain_right.n66 0.155672
R591 drain_right.n121 drain_right.n120 0.155672
R592 drain_right.n120 drain_right.n70 0.155672
R593 drain_right.n113 drain_right.n70 0.155672
R594 drain_right.n113 drain_right.n112 0.155672
R595 drain_right.n112 drain_right.n74 0.155672
R596 drain_right.n104 drain_right.n74 0.155672
R597 drain_right.n104 drain_right.n103 0.155672
R598 drain_right.n103 drain_right.n79 0.155672
R599 drain_right.n96 drain_right.n79 0.155672
R600 drain_right.n96 drain_right.n95 0.155672
R601 drain_right.n95 drain_right.n83 0.155672
R602 drain_right.n88 drain_right.n83 0.155672
R603 plus plus.t0 845.255
R604 plus plus.t1 830.413
R605 drain_left.n60 drain_left.n0 289.615
R606 drain_left.n125 drain_left.n65 289.615
R607 drain_left.n20 drain_left.n19 185
R608 drain_left.n25 drain_left.n24 185
R609 drain_left.n27 drain_left.n26 185
R610 drain_left.n16 drain_left.n15 185
R611 drain_left.n33 drain_left.n32 185
R612 drain_left.n35 drain_left.n34 185
R613 drain_left.n12 drain_left.n11 185
R614 drain_left.n42 drain_left.n41 185
R615 drain_left.n43 drain_left.n10 185
R616 drain_left.n45 drain_left.n44 185
R617 drain_left.n8 drain_left.n7 185
R618 drain_left.n51 drain_left.n50 185
R619 drain_left.n53 drain_left.n52 185
R620 drain_left.n4 drain_left.n3 185
R621 drain_left.n59 drain_left.n58 185
R622 drain_left.n61 drain_left.n60 185
R623 drain_left.n126 drain_left.n125 185
R624 drain_left.n124 drain_left.n123 185
R625 drain_left.n69 drain_left.n68 185
R626 drain_left.n118 drain_left.n117 185
R627 drain_left.n116 drain_left.n115 185
R628 drain_left.n73 drain_left.n72 185
R629 drain_left.n110 drain_left.n109 185
R630 drain_left.n108 drain_left.n75 185
R631 drain_left.n107 drain_left.n106 185
R632 drain_left.n78 drain_left.n76 185
R633 drain_left.n101 drain_left.n100 185
R634 drain_left.n99 drain_left.n98 185
R635 drain_left.n82 drain_left.n81 185
R636 drain_left.n93 drain_left.n92 185
R637 drain_left.n91 drain_left.n90 185
R638 drain_left.n86 drain_left.n85 185
R639 drain_left.n21 drain_left.t1 149.524
R640 drain_left.n87 drain_left.t0 149.524
R641 drain_left.n25 drain_left.n19 104.615
R642 drain_left.n26 drain_left.n25 104.615
R643 drain_left.n26 drain_left.n15 104.615
R644 drain_left.n33 drain_left.n15 104.615
R645 drain_left.n34 drain_left.n33 104.615
R646 drain_left.n34 drain_left.n11 104.615
R647 drain_left.n42 drain_left.n11 104.615
R648 drain_left.n43 drain_left.n42 104.615
R649 drain_left.n44 drain_left.n43 104.615
R650 drain_left.n44 drain_left.n7 104.615
R651 drain_left.n51 drain_left.n7 104.615
R652 drain_left.n52 drain_left.n51 104.615
R653 drain_left.n52 drain_left.n3 104.615
R654 drain_left.n59 drain_left.n3 104.615
R655 drain_left.n60 drain_left.n59 104.615
R656 drain_left.n125 drain_left.n124 104.615
R657 drain_left.n124 drain_left.n68 104.615
R658 drain_left.n117 drain_left.n68 104.615
R659 drain_left.n117 drain_left.n116 104.615
R660 drain_left.n116 drain_left.n72 104.615
R661 drain_left.n109 drain_left.n72 104.615
R662 drain_left.n109 drain_left.n108 104.615
R663 drain_left.n108 drain_left.n107 104.615
R664 drain_left.n107 drain_left.n76 104.615
R665 drain_left.n100 drain_left.n76 104.615
R666 drain_left.n100 drain_left.n99 104.615
R667 drain_left.n99 drain_left.n81 104.615
R668 drain_left.n92 drain_left.n81 104.615
R669 drain_left.n92 drain_left.n91 104.615
R670 drain_left.n91 drain_left.n85 104.615
R671 drain_left drain_left.n64 74.9365
R672 drain_left drain_left.n129 52.9051
R673 drain_left.t1 drain_left.n19 52.3082
R674 drain_left.t0 drain_left.n85 52.3082
R675 drain_left.n45 drain_left.n10 13.1884
R676 drain_left.n110 drain_left.n75 13.1884
R677 drain_left.n41 drain_left.n40 12.8005
R678 drain_left.n46 drain_left.n8 12.8005
R679 drain_left.n111 drain_left.n73 12.8005
R680 drain_left.n106 drain_left.n77 12.8005
R681 drain_left.n39 drain_left.n12 12.0247
R682 drain_left.n50 drain_left.n49 12.0247
R683 drain_left.n115 drain_left.n114 12.0247
R684 drain_left.n105 drain_left.n78 12.0247
R685 drain_left.n36 drain_left.n35 11.249
R686 drain_left.n53 drain_left.n6 11.249
R687 drain_left.n118 drain_left.n71 11.249
R688 drain_left.n102 drain_left.n101 11.249
R689 drain_left.n32 drain_left.n14 10.4732
R690 drain_left.n54 drain_left.n4 10.4732
R691 drain_left.n119 drain_left.n69 10.4732
R692 drain_left.n98 drain_left.n80 10.4732
R693 drain_left.n21 drain_left.n20 10.2747
R694 drain_left.n87 drain_left.n86 10.2747
R695 drain_left.n31 drain_left.n16 9.69747
R696 drain_left.n58 drain_left.n57 9.69747
R697 drain_left.n123 drain_left.n122 9.69747
R698 drain_left.n97 drain_left.n82 9.69747
R699 drain_left.n64 drain_left.n63 9.45567
R700 drain_left.n129 drain_left.n128 9.45567
R701 drain_left.n63 drain_left.n62 9.3005
R702 drain_left.n2 drain_left.n1 9.3005
R703 drain_left.n57 drain_left.n56 9.3005
R704 drain_left.n55 drain_left.n54 9.3005
R705 drain_left.n6 drain_left.n5 9.3005
R706 drain_left.n49 drain_left.n48 9.3005
R707 drain_left.n47 drain_left.n46 9.3005
R708 drain_left.n23 drain_left.n22 9.3005
R709 drain_left.n18 drain_left.n17 9.3005
R710 drain_left.n29 drain_left.n28 9.3005
R711 drain_left.n31 drain_left.n30 9.3005
R712 drain_left.n14 drain_left.n13 9.3005
R713 drain_left.n37 drain_left.n36 9.3005
R714 drain_left.n39 drain_left.n38 9.3005
R715 drain_left.n40 drain_left.n9 9.3005
R716 drain_left.n89 drain_left.n88 9.3005
R717 drain_left.n84 drain_left.n83 9.3005
R718 drain_left.n95 drain_left.n94 9.3005
R719 drain_left.n97 drain_left.n96 9.3005
R720 drain_left.n80 drain_left.n79 9.3005
R721 drain_left.n103 drain_left.n102 9.3005
R722 drain_left.n105 drain_left.n104 9.3005
R723 drain_left.n77 drain_left.n74 9.3005
R724 drain_left.n128 drain_left.n127 9.3005
R725 drain_left.n67 drain_left.n66 9.3005
R726 drain_left.n122 drain_left.n121 9.3005
R727 drain_left.n120 drain_left.n119 9.3005
R728 drain_left.n71 drain_left.n70 9.3005
R729 drain_left.n114 drain_left.n113 9.3005
R730 drain_left.n112 drain_left.n111 9.3005
R731 drain_left.n28 drain_left.n27 8.92171
R732 drain_left.n61 drain_left.n2 8.92171
R733 drain_left.n126 drain_left.n67 8.92171
R734 drain_left.n94 drain_left.n93 8.92171
R735 drain_left.n24 drain_left.n18 8.14595
R736 drain_left.n62 drain_left.n0 8.14595
R737 drain_left.n127 drain_left.n65 8.14595
R738 drain_left.n90 drain_left.n84 8.14595
R739 drain_left.n23 drain_left.n20 7.3702
R740 drain_left.n89 drain_left.n86 7.3702
R741 drain_left.n24 drain_left.n23 5.81868
R742 drain_left.n64 drain_left.n0 5.81868
R743 drain_left.n129 drain_left.n65 5.81868
R744 drain_left.n90 drain_left.n89 5.81868
R745 drain_left.n27 drain_left.n18 5.04292
R746 drain_left.n62 drain_left.n61 5.04292
R747 drain_left.n127 drain_left.n126 5.04292
R748 drain_left.n93 drain_left.n84 5.04292
R749 drain_left.n28 drain_left.n16 4.26717
R750 drain_left.n58 drain_left.n2 4.26717
R751 drain_left.n123 drain_left.n67 4.26717
R752 drain_left.n94 drain_left.n82 4.26717
R753 drain_left.n32 drain_left.n31 3.49141
R754 drain_left.n57 drain_left.n4 3.49141
R755 drain_left.n122 drain_left.n69 3.49141
R756 drain_left.n98 drain_left.n97 3.49141
R757 drain_left.n22 drain_left.n21 2.84303
R758 drain_left.n88 drain_left.n87 2.84303
R759 drain_left.n35 drain_left.n14 2.71565
R760 drain_left.n54 drain_left.n53 2.71565
R761 drain_left.n119 drain_left.n118 2.71565
R762 drain_left.n101 drain_left.n80 2.71565
R763 drain_left.n36 drain_left.n12 1.93989
R764 drain_left.n50 drain_left.n6 1.93989
R765 drain_left.n115 drain_left.n71 1.93989
R766 drain_left.n102 drain_left.n78 1.93989
R767 drain_left.n41 drain_left.n39 1.16414
R768 drain_left.n49 drain_left.n8 1.16414
R769 drain_left.n114 drain_left.n73 1.16414
R770 drain_left.n106 drain_left.n105 1.16414
R771 drain_left.n40 drain_left.n10 0.388379
R772 drain_left.n46 drain_left.n45 0.388379
R773 drain_left.n111 drain_left.n110 0.388379
R774 drain_left.n77 drain_left.n75 0.388379
R775 drain_left.n22 drain_left.n17 0.155672
R776 drain_left.n29 drain_left.n17 0.155672
R777 drain_left.n30 drain_left.n29 0.155672
R778 drain_left.n30 drain_left.n13 0.155672
R779 drain_left.n37 drain_left.n13 0.155672
R780 drain_left.n38 drain_left.n37 0.155672
R781 drain_left.n38 drain_left.n9 0.155672
R782 drain_left.n47 drain_left.n9 0.155672
R783 drain_left.n48 drain_left.n47 0.155672
R784 drain_left.n48 drain_left.n5 0.155672
R785 drain_left.n55 drain_left.n5 0.155672
R786 drain_left.n56 drain_left.n55 0.155672
R787 drain_left.n56 drain_left.n1 0.155672
R788 drain_left.n63 drain_left.n1 0.155672
R789 drain_left.n128 drain_left.n66 0.155672
R790 drain_left.n121 drain_left.n66 0.155672
R791 drain_left.n121 drain_left.n120 0.155672
R792 drain_left.n120 drain_left.n70 0.155672
R793 drain_left.n113 drain_left.n70 0.155672
R794 drain_left.n113 drain_left.n112 0.155672
R795 drain_left.n112 drain_left.n74 0.155672
R796 drain_left.n104 drain_left.n74 0.155672
R797 drain_left.n104 drain_left.n103 0.155672
R798 drain_left.n103 drain_left.n79 0.155672
R799 drain_left.n96 drain_left.n79 0.155672
R800 drain_left.n96 drain_left.n95 0.155672
R801 drain_left.n95 drain_left.n83 0.155672
R802 drain_left.n88 drain_left.n83 0.155672
C0 plus source 1.23411f
C1 plus minus 4.45179f
C2 drain_right source 6.2474f
C3 drain_right minus 1.76769f
C4 drain_left source 6.257451f
C5 drain_left minus 0.171767f
C6 plus drain_right 0.252683f
C7 plus drain_left 1.86128f
C8 drain_left drain_right 0.443275f
C9 minus source 1.2195f
C10 drain_right a_n1048_n3292# 5.71202f
C11 drain_left a_n1048_n3292# 5.87008f
C12 source a_n1048_n3292# 5.846318f
C13 minus a_n1048_n3292# 3.898337f
C14 plus a_n1048_n3292# 6.83266f
C15 drain_left.n0 a_n1048_n3292# 0.022022f
C16 drain_left.n1 a_n1048_n3292# 0.016625f
C17 drain_left.n2 a_n1048_n3292# 0.008934f
C18 drain_left.n3 a_n1048_n3292# 0.021116f
C19 drain_left.n4 a_n1048_n3292# 0.009459f
C20 drain_left.n5 a_n1048_n3292# 0.016625f
C21 drain_left.n6 a_n1048_n3292# 0.008934f
C22 drain_left.n7 a_n1048_n3292# 0.021116f
C23 drain_left.n8 a_n1048_n3292# 0.009459f
C24 drain_left.n9 a_n1048_n3292# 0.016625f
C25 drain_left.n10 a_n1048_n3292# 0.009196f
C26 drain_left.n11 a_n1048_n3292# 0.021116f
C27 drain_left.n12 a_n1048_n3292# 0.009459f
C28 drain_left.n13 a_n1048_n3292# 0.016625f
C29 drain_left.n14 a_n1048_n3292# 0.008934f
C30 drain_left.n15 a_n1048_n3292# 0.021116f
C31 drain_left.n16 a_n1048_n3292# 0.009459f
C32 drain_left.n17 a_n1048_n3292# 0.016625f
C33 drain_left.n18 a_n1048_n3292# 0.008934f
C34 drain_left.n19 a_n1048_n3292# 0.015837f
C35 drain_left.n20 a_n1048_n3292# 0.014927f
C36 drain_left.t1 a_n1048_n3292# 0.035663f
C37 drain_left.n21 a_n1048_n3292# 0.119866f
C38 drain_left.n22 a_n1048_n3292# 0.838712f
C39 drain_left.n23 a_n1048_n3292# 0.008934f
C40 drain_left.n24 a_n1048_n3292# 0.009459f
C41 drain_left.n25 a_n1048_n3292# 0.021116f
C42 drain_left.n26 a_n1048_n3292# 0.021116f
C43 drain_left.n27 a_n1048_n3292# 0.009459f
C44 drain_left.n28 a_n1048_n3292# 0.008934f
C45 drain_left.n29 a_n1048_n3292# 0.016625f
C46 drain_left.n30 a_n1048_n3292# 0.016625f
C47 drain_left.n31 a_n1048_n3292# 0.008934f
C48 drain_left.n32 a_n1048_n3292# 0.009459f
C49 drain_left.n33 a_n1048_n3292# 0.021116f
C50 drain_left.n34 a_n1048_n3292# 0.021116f
C51 drain_left.n35 a_n1048_n3292# 0.009459f
C52 drain_left.n36 a_n1048_n3292# 0.008934f
C53 drain_left.n37 a_n1048_n3292# 0.016625f
C54 drain_left.n38 a_n1048_n3292# 0.016625f
C55 drain_left.n39 a_n1048_n3292# 0.008934f
C56 drain_left.n40 a_n1048_n3292# 0.008934f
C57 drain_left.n41 a_n1048_n3292# 0.009459f
C58 drain_left.n42 a_n1048_n3292# 0.021116f
C59 drain_left.n43 a_n1048_n3292# 0.021116f
C60 drain_left.n44 a_n1048_n3292# 0.021116f
C61 drain_left.n45 a_n1048_n3292# 0.009196f
C62 drain_left.n46 a_n1048_n3292# 0.008934f
C63 drain_left.n47 a_n1048_n3292# 0.016625f
C64 drain_left.n48 a_n1048_n3292# 0.016625f
C65 drain_left.n49 a_n1048_n3292# 0.008934f
C66 drain_left.n50 a_n1048_n3292# 0.009459f
C67 drain_left.n51 a_n1048_n3292# 0.021116f
C68 drain_left.n52 a_n1048_n3292# 0.021116f
C69 drain_left.n53 a_n1048_n3292# 0.009459f
C70 drain_left.n54 a_n1048_n3292# 0.008934f
C71 drain_left.n55 a_n1048_n3292# 0.016625f
C72 drain_left.n56 a_n1048_n3292# 0.016625f
C73 drain_left.n57 a_n1048_n3292# 0.008934f
C74 drain_left.n58 a_n1048_n3292# 0.009459f
C75 drain_left.n59 a_n1048_n3292# 0.021116f
C76 drain_left.n60 a_n1048_n3292# 0.043332f
C77 drain_left.n61 a_n1048_n3292# 0.009459f
C78 drain_left.n62 a_n1048_n3292# 0.008934f
C79 drain_left.n63 a_n1048_n3292# 0.035703f
C80 drain_left.n64 a_n1048_n3292# 0.294725f
C81 drain_left.n65 a_n1048_n3292# 0.022022f
C82 drain_left.n66 a_n1048_n3292# 0.016625f
C83 drain_left.n67 a_n1048_n3292# 0.008934f
C84 drain_left.n68 a_n1048_n3292# 0.021116f
C85 drain_left.n69 a_n1048_n3292# 0.009459f
C86 drain_left.n70 a_n1048_n3292# 0.016625f
C87 drain_left.n71 a_n1048_n3292# 0.008934f
C88 drain_left.n72 a_n1048_n3292# 0.021116f
C89 drain_left.n73 a_n1048_n3292# 0.009459f
C90 drain_left.n74 a_n1048_n3292# 0.016625f
C91 drain_left.n75 a_n1048_n3292# 0.009196f
C92 drain_left.n76 a_n1048_n3292# 0.021116f
C93 drain_left.n77 a_n1048_n3292# 0.008934f
C94 drain_left.n78 a_n1048_n3292# 0.009459f
C95 drain_left.n79 a_n1048_n3292# 0.016625f
C96 drain_left.n80 a_n1048_n3292# 0.008934f
C97 drain_left.n81 a_n1048_n3292# 0.021116f
C98 drain_left.n82 a_n1048_n3292# 0.009459f
C99 drain_left.n83 a_n1048_n3292# 0.016625f
C100 drain_left.n84 a_n1048_n3292# 0.008934f
C101 drain_left.n85 a_n1048_n3292# 0.015837f
C102 drain_left.n86 a_n1048_n3292# 0.014927f
C103 drain_left.t0 a_n1048_n3292# 0.035663f
C104 drain_left.n87 a_n1048_n3292# 0.119866f
C105 drain_left.n88 a_n1048_n3292# 0.838712f
C106 drain_left.n89 a_n1048_n3292# 0.008934f
C107 drain_left.n90 a_n1048_n3292# 0.009459f
C108 drain_left.n91 a_n1048_n3292# 0.021116f
C109 drain_left.n92 a_n1048_n3292# 0.021116f
C110 drain_left.n93 a_n1048_n3292# 0.009459f
C111 drain_left.n94 a_n1048_n3292# 0.008934f
C112 drain_left.n95 a_n1048_n3292# 0.016625f
C113 drain_left.n96 a_n1048_n3292# 0.016625f
C114 drain_left.n97 a_n1048_n3292# 0.008934f
C115 drain_left.n98 a_n1048_n3292# 0.009459f
C116 drain_left.n99 a_n1048_n3292# 0.021116f
C117 drain_left.n100 a_n1048_n3292# 0.021116f
C118 drain_left.n101 a_n1048_n3292# 0.009459f
C119 drain_left.n102 a_n1048_n3292# 0.008934f
C120 drain_left.n103 a_n1048_n3292# 0.016625f
C121 drain_left.n104 a_n1048_n3292# 0.016625f
C122 drain_left.n105 a_n1048_n3292# 0.008934f
C123 drain_left.n106 a_n1048_n3292# 0.009459f
C124 drain_left.n107 a_n1048_n3292# 0.021116f
C125 drain_left.n108 a_n1048_n3292# 0.021116f
C126 drain_left.n109 a_n1048_n3292# 0.021116f
C127 drain_left.n110 a_n1048_n3292# 0.009196f
C128 drain_left.n111 a_n1048_n3292# 0.008934f
C129 drain_left.n112 a_n1048_n3292# 0.016625f
C130 drain_left.n113 a_n1048_n3292# 0.016625f
C131 drain_left.n114 a_n1048_n3292# 0.008934f
C132 drain_left.n115 a_n1048_n3292# 0.009459f
C133 drain_left.n116 a_n1048_n3292# 0.021116f
C134 drain_left.n117 a_n1048_n3292# 0.021116f
C135 drain_left.n118 a_n1048_n3292# 0.009459f
C136 drain_left.n119 a_n1048_n3292# 0.008934f
C137 drain_left.n120 a_n1048_n3292# 0.016625f
C138 drain_left.n121 a_n1048_n3292# 0.016625f
C139 drain_left.n122 a_n1048_n3292# 0.008934f
C140 drain_left.n123 a_n1048_n3292# 0.009459f
C141 drain_left.n124 a_n1048_n3292# 0.021116f
C142 drain_left.n125 a_n1048_n3292# 0.043332f
C143 drain_left.n126 a_n1048_n3292# 0.009459f
C144 drain_left.n127 a_n1048_n3292# 0.008934f
C145 drain_left.n128 a_n1048_n3292# 0.035703f
C146 drain_left.n129 a_n1048_n3292# 0.06089f
C147 plus.t1 a_n1048_n3292# 0.694287f
C148 plus.t0 a_n1048_n3292# 0.722303f
C149 drain_right.n0 a_n1048_n3292# 0.021899f
C150 drain_right.n1 a_n1048_n3292# 0.016532f
C151 drain_right.n2 a_n1048_n3292# 0.008884f
C152 drain_right.n3 a_n1048_n3292# 0.020998f
C153 drain_right.n4 a_n1048_n3292# 0.009406f
C154 drain_right.n5 a_n1048_n3292# 0.016532f
C155 drain_right.n6 a_n1048_n3292# 0.008884f
C156 drain_right.n7 a_n1048_n3292# 0.020998f
C157 drain_right.n8 a_n1048_n3292# 0.009406f
C158 drain_right.n9 a_n1048_n3292# 0.016532f
C159 drain_right.n10 a_n1048_n3292# 0.009145f
C160 drain_right.n11 a_n1048_n3292# 0.020998f
C161 drain_right.n12 a_n1048_n3292# 0.009406f
C162 drain_right.n13 a_n1048_n3292# 0.016532f
C163 drain_right.n14 a_n1048_n3292# 0.008884f
C164 drain_right.n15 a_n1048_n3292# 0.020998f
C165 drain_right.n16 a_n1048_n3292# 0.009406f
C166 drain_right.n17 a_n1048_n3292# 0.016532f
C167 drain_right.n18 a_n1048_n3292# 0.008884f
C168 drain_right.n19 a_n1048_n3292# 0.015748f
C169 drain_right.n20 a_n1048_n3292# 0.014844f
C170 drain_right.t0 a_n1048_n3292# 0.035463f
C171 drain_right.n21 a_n1048_n3292# 0.119193f
C172 drain_right.n22 a_n1048_n3292# 0.834009f
C173 drain_right.n23 a_n1048_n3292# 0.008884f
C174 drain_right.n24 a_n1048_n3292# 0.009406f
C175 drain_right.n25 a_n1048_n3292# 0.020998f
C176 drain_right.n26 a_n1048_n3292# 0.020998f
C177 drain_right.n27 a_n1048_n3292# 0.009406f
C178 drain_right.n28 a_n1048_n3292# 0.008884f
C179 drain_right.n29 a_n1048_n3292# 0.016532f
C180 drain_right.n30 a_n1048_n3292# 0.016532f
C181 drain_right.n31 a_n1048_n3292# 0.008884f
C182 drain_right.n32 a_n1048_n3292# 0.009406f
C183 drain_right.n33 a_n1048_n3292# 0.020998f
C184 drain_right.n34 a_n1048_n3292# 0.020998f
C185 drain_right.n35 a_n1048_n3292# 0.009406f
C186 drain_right.n36 a_n1048_n3292# 0.008884f
C187 drain_right.n37 a_n1048_n3292# 0.016532f
C188 drain_right.n38 a_n1048_n3292# 0.016532f
C189 drain_right.n39 a_n1048_n3292# 0.008884f
C190 drain_right.n40 a_n1048_n3292# 0.008884f
C191 drain_right.n41 a_n1048_n3292# 0.009406f
C192 drain_right.n42 a_n1048_n3292# 0.020998f
C193 drain_right.n43 a_n1048_n3292# 0.020998f
C194 drain_right.n44 a_n1048_n3292# 0.020998f
C195 drain_right.n45 a_n1048_n3292# 0.009145f
C196 drain_right.n46 a_n1048_n3292# 0.008884f
C197 drain_right.n47 a_n1048_n3292# 0.016532f
C198 drain_right.n48 a_n1048_n3292# 0.016532f
C199 drain_right.n49 a_n1048_n3292# 0.008884f
C200 drain_right.n50 a_n1048_n3292# 0.009406f
C201 drain_right.n51 a_n1048_n3292# 0.020998f
C202 drain_right.n52 a_n1048_n3292# 0.020998f
C203 drain_right.n53 a_n1048_n3292# 0.009406f
C204 drain_right.n54 a_n1048_n3292# 0.008884f
C205 drain_right.n55 a_n1048_n3292# 0.016532f
C206 drain_right.n56 a_n1048_n3292# 0.016532f
C207 drain_right.n57 a_n1048_n3292# 0.008884f
C208 drain_right.n58 a_n1048_n3292# 0.009406f
C209 drain_right.n59 a_n1048_n3292# 0.020998f
C210 drain_right.n60 a_n1048_n3292# 0.043089f
C211 drain_right.n61 a_n1048_n3292# 0.009406f
C212 drain_right.n62 a_n1048_n3292# 0.008884f
C213 drain_right.n63 a_n1048_n3292# 0.035503f
C214 drain_right.n64 a_n1048_n3292# 0.276926f
C215 drain_right.n65 a_n1048_n3292# 0.021899f
C216 drain_right.n66 a_n1048_n3292# 0.016532f
C217 drain_right.n67 a_n1048_n3292# 0.008884f
C218 drain_right.n68 a_n1048_n3292# 0.020998f
C219 drain_right.n69 a_n1048_n3292# 0.009406f
C220 drain_right.n70 a_n1048_n3292# 0.016532f
C221 drain_right.n71 a_n1048_n3292# 0.008884f
C222 drain_right.n72 a_n1048_n3292# 0.020998f
C223 drain_right.n73 a_n1048_n3292# 0.009406f
C224 drain_right.n74 a_n1048_n3292# 0.016532f
C225 drain_right.n75 a_n1048_n3292# 0.009145f
C226 drain_right.n76 a_n1048_n3292# 0.020998f
C227 drain_right.n77 a_n1048_n3292# 0.008884f
C228 drain_right.n78 a_n1048_n3292# 0.009406f
C229 drain_right.n79 a_n1048_n3292# 0.016532f
C230 drain_right.n80 a_n1048_n3292# 0.008884f
C231 drain_right.n81 a_n1048_n3292# 0.020998f
C232 drain_right.n82 a_n1048_n3292# 0.009406f
C233 drain_right.n83 a_n1048_n3292# 0.016532f
C234 drain_right.n84 a_n1048_n3292# 0.008884f
C235 drain_right.n85 a_n1048_n3292# 0.015748f
C236 drain_right.n86 a_n1048_n3292# 0.014844f
C237 drain_right.t1 a_n1048_n3292# 0.035463f
C238 drain_right.n87 a_n1048_n3292# 0.119193f
C239 drain_right.n88 a_n1048_n3292# 0.834009f
C240 drain_right.n89 a_n1048_n3292# 0.008884f
C241 drain_right.n90 a_n1048_n3292# 0.009406f
C242 drain_right.n91 a_n1048_n3292# 0.020998f
C243 drain_right.n92 a_n1048_n3292# 0.020998f
C244 drain_right.n93 a_n1048_n3292# 0.009406f
C245 drain_right.n94 a_n1048_n3292# 0.008884f
C246 drain_right.n95 a_n1048_n3292# 0.016532f
C247 drain_right.n96 a_n1048_n3292# 0.016532f
C248 drain_right.n97 a_n1048_n3292# 0.008884f
C249 drain_right.n98 a_n1048_n3292# 0.009406f
C250 drain_right.n99 a_n1048_n3292# 0.020998f
C251 drain_right.n100 a_n1048_n3292# 0.020998f
C252 drain_right.n101 a_n1048_n3292# 0.009406f
C253 drain_right.n102 a_n1048_n3292# 0.008884f
C254 drain_right.n103 a_n1048_n3292# 0.016532f
C255 drain_right.n104 a_n1048_n3292# 0.016532f
C256 drain_right.n105 a_n1048_n3292# 0.008884f
C257 drain_right.n106 a_n1048_n3292# 0.009406f
C258 drain_right.n107 a_n1048_n3292# 0.020998f
C259 drain_right.n108 a_n1048_n3292# 0.020998f
C260 drain_right.n109 a_n1048_n3292# 0.020998f
C261 drain_right.n110 a_n1048_n3292# 0.009145f
C262 drain_right.n111 a_n1048_n3292# 0.008884f
C263 drain_right.n112 a_n1048_n3292# 0.016532f
C264 drain_right.n113 a_n1048_n3292# 0.016532f
C265 drain_right.n114 a_n1048_n3292# 0.008884f
C266 drain_right.n115 a_n1048_n3292# 0.009406f
C267 drain_right.n116 a_n1048_n3292# 0.020998f
C268 drain_right.n117 a_n1048_n3292# 0.020998f
C269 drain_right.n118 a_n1048_n3292# 0.009406f
C270 drain_right.n119 a_n1048_n3292# 0.008884f
C271 drain_right.n120 a_n1048_n3292# 0.016532f
C272 drain_right.n121 a_n1048_n3292# 0.016532f
C273 drain_right.n122 a_n1048_n3292# 0.008884f
C274 drain_right.n123 a_n1048_n3292# 0.009406f
C275 drain_right.n124 a_n1048_n3292# 0.020998f
C276 drain_right.n125 a_n1048_n3292# 0.043089f
C277 drain_right.n126 a_n1048_n3292# 0.009406f
C278 drain_right.n127 a_n1048_n3292# 0.008884f
C279 drain_right.n128 a_n1048_n3292# 0.035503f
C280 drain_right.n129 a_n1048_n3292# 0.060386f
C281 source.n0 a_n1048_n3292# 0.02355f
C282 source.n1 a_n1048_n3292# 0.017779f
C283 source.n2 a_n1048_n3292# 0.009554f
C284 source.n3 a_n1048_n3292# 0.022581f
C285 source.n4 a_n1048_n3292# 0.010116f
C286 source.n5 a_n1048_n3292# 0.017779f
C287 source.n6 a_n1048_n3292# 0.009554f
C288 source.n7 a_n1048_n3292# 0.022581f
C289 source.n8 a_n1048_n3292# 0.010116f
C290 source.n9 a_n1048_n3292# 0.017779f
C291 source.n10 a_n1048_n3292# 0.009835f
C292 source.n11 a_n1048_n3292# 0.022581f
C293 source.n12 a_n1048_n3292# 0.009554f
C294 source.n13 a_n1048_n3292# 0.010116f
C295 source.n14 a_n1048_n3292# 0.017779f
C296 source.n15 a_n1048_n3292# 0.009554f
C297 source.n16 a_n1048_n3292# 0.022581f
C298 source.n17 a_n1048_n3292# 0.010116f
C299 source.n18 a_n1048_n3292# 0.017779f
C300 source.n19 a_n1048_n3292# 0.009554f
C301 source.n20 a_n1048_n3292# 0.016936f
C302 source.n21 a_n1048_n3292# 0.015963f
C303 source.t0 a_n1048_n3292# 0.038138f
C304 source.n22 a_n1048_n3292# 0.128183f
C305 source.n23 a_n1048_n3292# 0.896907f
C306 source.n24 a_n1048_n3292# 0.009554f
C307 source.n25 a_n1048_n3292# 0.010116f
C308 source.n26 a_n1048_n3292# 0.022581f
C309 source.n27 a_n1048_n3292# 0.022581f
C310 source.n28 a_n1048_n3292# 0.010116f
C311 source.n29 a_n1048_n3292# 0.009554f
C312 source.n30 a_n1048_n3292# 0.017779f
C313 source.n31 a_n1048_n3292# 0.017779f
C314 source.n32 a_n1048_n3292# 0.009554f
C315 source.n33 a_n1048_n3292# 0.010116f
C316 source.n34 a_n1048_n3292# 0.022581f
C317 source.n35 a_n1048_n3292# 0.022581f
C318 source.n36 a_n1048_n3292# 0.010116f
C319 source.n37 a_n1048_n3292# 0.009554f
C320 source.n38 a_n1048_n3292# 0.017779f
C321 source.n39 a_n1048_n3292# 0.017779f
C322 source.n40 a_n1048_n3292# 0.009554f
C323 source.n41 a_n1048_n3292# 0.010116f
C324 source.n42 a_n1048_n3292# 0.022581f
C325 source.n43 a_n1048_n3292# 0.022581f
C326 source.n44 a_n1048_n3292# 0.022581f
C327 source.n45 a_n1048_n3292# 0.009835f
C328 source.n46 a_n1048_n3292# 0.009554f
C329 source.n47 a_n1048_n3292# 0.017779f
C330 source.n48 a_n1048_n3292# 0.017779f
C331 source.n49 a_n1048_n3292# 0.009554f
C332 source.n50 a_n1048_n3292# 0.010116f
C333 source.n51 a_n1048_n3292# 0.022581f
C334 source.n52 a_n1048_n3292# 0.022581f
C335 source.n53 a_n1048_n3292# 0.010116f
C336 source.n54 a_n1048_n3292# 0.009554f
C337 source.n55 a_n1048_n3292# 0.017779f
C338 source.n56 a_n1048_n3292# 0.017779f
C339 source.n57 a_n1048_n3292# 0.009554f
C340 source.n58 a_n1048_n3292# 0.010116f
C341 source.n59 a_n1048_n3292# 0.022581f
C342 source.n60 a_n1048_n3292# 0.046339f
C343 source.n61 a_n1048_n3292# 0.010116f
C344 source.n62 a_n1048_n3292# 0.009554f
C345 source.n63 a_n1048_n3292# 0.03818f
C346 source.n64 a_n1048_n3292# 0.025574f
C347 source.n65 a_n1048_n3292# 0.739124f
C348 source.n66 a_n1048_n3292# 0.02355f
C349 source.n67 a_n1048_n3292# 0.017779f
C350 source.n68 a_n1048_n3292# 0.009554f
C351 source.n69 a_n1048_n3292# 0.022581f
C352 source.n70 a_n1048_n3292# 0.010116f
C353 source.n71 a_n1048_n3292# 0.017779f
C354 source.n72 a_n1048_n3292# 0.009554f
C355 source.n73 a_n1048_n3292# 0.022581f
C356 source.n74 a_n1048_n3292# 0.010116f
C357 source.n75 a_n1048_n3292# 0.017779f
C358 source.n76 a_n1048_n3292# 0.009835f
C359 source.n77 a_n1048_n3292# 0.022581f
C360 source.n78 a_n1048_n3292# 0.009554f
C361 source.n79 a_n1048_n3292# 0.010116f
C362 source.n80 a_n1048_n3292# 0.017779f
C363 source.n81 a_n1048_n3292# 0.009554f
C364 source.n82 a_n1048_n3292# 0.022581f
C365 source.n83 a_n1048_n3292# 0.010116f
C366 source.n84 a_n1048_n3292# 0.017779f
C367 source.n85 a_n1048_n3292# 0.009554f
C368 source.n86 a_n1048_n3292# 0.016936f
C369 source.n87 a_n1048_n3292# 0.015963f
C370 source.t2 a_n1048_n3292# 0.038138f
C371 source.n88 a_n1048_n3292# 0.128183f
C372 source.n89 a_n1048_n3292# 0.896907f
C373 source.n90 a_n1048_n3292# 0.009554f
C374 source.n91 a_n1048_n3292# 0.010116f
C375 source.n92 a_n1048_n3292# 0.022581f
C376 source.n93 a_n1048_n3292# 0.022581f
C377 source.n94 a_n1048_n3292# 0.010116f
C378 source.n95 a_n1048_n3292# 0.009554f
C379 source.n96 a_n1048_n3292# 0.017779f
C380 source.n97 a_n1048_n3292# 0.017779f
C381 source.n98 a_n1048_n3292# 0.009554f
C382 source.n99 a_n1048_n3292# 0.010116f
C383 source.n100 a_n1048_n3292# 0.022581f
C384 source.n101 a_n1048_n3292# 0.022581f
C385 source.n102 a_n1048_n3292# 0.010116f
C386 source.n103 a_n1048_n3292# 0.009554f
C387 source.n104 a_n1048_n3292# 0.017779f
C388 source.n105 a_n1048_n3292# 0.017779f
C389 source.n106 a_n1048_n3292# 0.009554f
C390 source.n107 a_n1048_n3292# 0.010116f
C391 source.n108 a_n1048_n3292# 0.022581f
C392 source.n109 a_n1048_n3292# 0.022581f
C393 source.n110 a_n1048_n3292# 0.022581f
C394 source.n111 a_n1048_n3292# 0.009835f
C395 source.n112 a_n1048_n3292# 0.009554f
C396 source.n113 a_n1048_n3292# 0.017779f
C397 source.n114 a_n1048_n3292# 0.017779f
C398 source.n115 a_n1048_n3292# 0.009554f
C399 source.n116 a_n1048_n3292# 0.010116f
C400 source.n117 a_n1048_n3292# 0.022581f
C401 source.n118 a_n1048_n3292# 0.022581f
C402 source.n119 a_n1048_n3292# 0.010116f
C403 source.n120 a_n1048_n3292# 0.009554f
C404 source.n121 a_n1048_n3292# 0.017779f
C405 source.n122 a_n1048_n3292# 0.017779f
C406 source.n123 a_n1048_n3292# 0.009554f
C407 source.n124 a_n1048_n3292# 0.010116f
C408 source.n125 a_n1048_n3292# 0.022581f
C409 source.n126 a_n1048_n3292# 0.046339f
C410 source.n127 a_n1048_n3292# 0.010116f
C411 source.n128 a_n1048_n3292# 0.009554f
C412 source.n129 a_n1048_n3292# 0.03818f
C413 source.n130 a_n1048_n3292# 0.025574f
C414 source.n131 a_n1048_n3292# 1.06335f
C415 source.n132 a_n1048_n3292# 0.02355f
C416 source.n133 a_n1048_n3292# 0.017779f
C417 source.n134 a_n1048_n3292# 0.009554f
C418 source.n135 a_n1048_n3292# 0.022581f
C419 source.n136 a_n1048_n3292# 0.010116f
C420 source.n137 a_n1048_n3292# 0.017779f
C421 source.n138 a_n1048_n3292# 0.009554f
C422 source.n139 a_n1048_n3292# 0.022581f
C423 source.n140 a_n1048_n3292# 0.010116f
C424 source.n141 a_n1048_n3292# 0.017779f
C425 source.n142 a_n1048_n3292# 0.009835f
C426 source.n143 a_n1048_n3292# 0.022581f
C427 source.n144 a_n1048_n3292# 0.010116f
C428 source.n145 a_n1048_n3292# 0.017779f
C429 source.n146 a_n1048_n3292# 0.009554f
C430 source.n147 a_n1048_n3292# 0.022581f
C431 source.n148 a_n1048_n3292# 0.010116f
C432 source.n149 a_n1048_n3292# 0.017779f
C433 source.n150 a_n1048_n3292# 0.009554f
C434 source.n151 a_n1048_n3292# 0.016936f
C435 source.n152 a_n1048_n3292# 0.015963f
C436 source.t1 a_n1048_n3292# 0.038138f
C437 source.n153 a_n1048_n3292# 0.128183f
C438 source.n154 a_n1048_n3292# 0.896907f
C439 source.n155 a_n1048_n3292# 0.009554f
C440 source.n156 a_n1048_n3292# 0.010116f
C441 source.n157 a_n1048_n3292# 0.022581f
C442 source.n158 a_n1048_n3292# 0.022581f
C443 source.n159 a_n1048_n3292# 0.010116f
C444 source.n160 a_n1048_n3292# 0.009554f
C445 source.n161 a_n1048_n3292# 0.017779f
C446 source.n162 a_n1048_n3292# 0.017779f
C447 source.n163 a_n1048_n3292# 0.009554f
C448 source.n164 a_n1048_n3292# 0.010116f
C449 source.n165 a_n1048_n3292# 0.022581f
C450 source.n166 a_n1048_n3292# 0.022581f
C451 source.n167 a_n1048_n3292# 0.010116f
C452 source.n168 a_n1048_n3292# 0.009554f
C453 source.n169 a_n1048_n3292# 0.017779f
C454 source.n170 a_n1048_n3292# 0.017779f
C455 source.n171 a_n1048_n3292# 0.009554f
C456 source.n172 a_n1048_n3292# 0.009554f
C457 source.n173 a_n1048_n3292# 0.010116f
C458 source.n174 a_n1048_n3292# 0.022581f
C459 source.n175 a_n1048_n3292# 0.022581f
C460 source.n176 a_n1048_n3292# 0.022581f
C461 source.n177 a_n1048_n3292# 0.009835f
C462 source.n178 a_n1048_n3292# 0.009554f
C463 source.n179 a_n1048_n3292# 0.017779f
C464 source.n180 a_n1048_n3292# 0.017779f
C465 source.n181 a_n1048_n3292# 0.009554f
C466 source.n182 a_n1048_n3292# 0.010116f
C467 source.n183 a_n1048_n3292# 0.022581f
C468 source.n184 a_n1048_n3292# 0.022581f
C469 source.n185 a_n1048_n3292# 0.010116f
C470 source.n186 a_n1048_n3292# 0.009554f
C471 source.n187 a_n1048_n3292# 0.017779f
C472 source.n188 a_n1048_n3292# 0.017779f
C473 source.n189 a_n1048_n3292# 0.009554f
C474 source.n190 a_n1048_n3292# 0.010116f
C475 source.n191 a_n1048_n3292# 0.022581f
C476 source.n192 a_n1048_n3292# 0.046339f
C477 source.n193 a_n1048_n3292# 0.010116f
C478 source.n194 a_n1048_n3292# 0.009554f
C479 source.n195 a_n1048_n3292# 0.03818f
C480 source.n196 a_n1048_n3292# 0.025574f
C481 source.n197 a_n1048_n3292# 1.06335f
C482 source.n198 a_n1048_n3292# 0.02355f
C483 source.n199 a_n1048_n3292# 0.017779f
C484 source.n200 a_n1048_n3292# 0.009554f
C485 source.n201 a_n1048_n3292# 0.022581f
C486 source.n202 a_n1048_n3292# 0.010116f
C487 source.n203 a_n1048_n3292# 0.017779f
C488 source.n204 a_n1048_n3292# 0.009554f
C489 source.n205 a_n1048_n3292# 0.022581f
C490 source.n206 a_n1048_n3292# 0.010116f
C491 source.n207 a_n1048_n3292# 0.017779f
C492 source.n208 a_n1048_n3292# 0.009835f
C493 source.n209 a_n1048_n3292# 0.022581f
C494 source.n210 a_n1048_n3292# 0.010116f
C495 source.n211 a_n1048_n3292# 0.017779f
C496 source.n212 a_n1048_n3292# 0.009554f
C497 source.n213 a_n1048_n3292# 0.022581f
C498 source.n214 a_n1048_n3292# 0.010116f
C499 source.n215 a_n1048_n3292# 0.017779f
C500 source.n216 a_n1048_n3292# 0.009554f
C501 source.n217 a_n1048_n3292# 0.016936f
C502 source.n218 a_n1048_n3292# 0.015963f
C503 source.t3 a_n1048_n3292# 0.038138f
C504 source.n219 a_n1048_n3292# 0.128183f
C505 source.n220 a_n1048_n3292# 0.896907f
C506 source.n221 a_n1048_n3292# 0.009554f
C507 source.n222 a_n1048_n3292# 0.010116f
C508 source.n223 a_n1048_n3292# 0.022581f
C509 source.n224 a_n1048_n3292# 0.022581f
C510 source.n225 a_n1048_n3292# 0.010116f
C511 source.n226 a_n1048_n3292# 0.009554f
C512 source.n227 a_n1048_n3292# 0.017779f
C513 source.n228 a_n1048_n3292# 0.017779f
C514 source.n229 a_n1048_n3292# 0.009554f
C515 source.n230 a_n1048_n3292# 0.010116f
C516 source.n231 a_n1048_n3292# 0.022581f
C517 source.n232 a_n1048_n3292# 0.022581f
C518 source.n233 a_n1048_n3292# 0.010116f
C519 source.n234 a_n1048_n3292# 0.009554f
C520 source.n235 a_n1048_n3292# 0.017779f
C521 source.n236 a_n1048_n3292# 0.017779f
C522 source.n237 a_n1048_n3292# 0.009554f
C523 source.n238 a_n1048_n3292# 0.009554f
C524 source.n239 a_n1048_n3292# 0.010116f
C525 source.n240 a_n1048_n3292# 0.022581f
C526 source.n241 a_n1048_n3292# 0.022581f
C527 source.n242 a_n1048_n3292# 0.022581f
C528 source.n243 a_n1048_n3292# 0.009835f
C529 source.n244 a_n1048_n3292# 0.009554f
C530 source.n245 a_n1048_n3292# 0.017779f
C531 source.n246 a_n1048_n3292# 0.017779f
C532 source.n247 a_n1048_n3292# 0.009554f
C533 source.n248 a_n1048_n3292# 0.010116f
C534 source.n249 a_n1048_n3292# 0.022581f
C535 source.n250 a_n1048_n3292# 0.022581f
C536 source.n251 a_n1048_n3292# 0.010116f
C537 source.n252 a_n1048_n3292# 0.009554f
C538 source.n253 a_n1048_n3292# 0.017779f
C539 source.n254 a_n1048_n3292# 0.017779f
C540 source.n255 a_n1048_n3292# 0.009554f
C541 source.n256 a_n1048_n3292# 0.010116f
C542 source.n257 a_n1048_n3292# 0.022581f
C543 source.n258 a_n1048_n3292# 0.046339f
C544 source.n259 a_n1048_n3292# 0.010116f
C545 source.n260 a_n1048_n3292# 0.009554f
C546 source.n261 a_n1048_n3292# 0.03818f
C547 source.n262 a_n1048_n3292# 0.025574f
C548 source.n263 a_n1048_n3292# 0.196078f
C549 source.n264 a_n1048_n3292# 1.12216f
C550 minus.t0 a_n1048_n3292# 0.725258f
C551 minus.t1 a_n1048_n3292# 0.677448f
C552 minus.n0 a_n1048_n3292# 3.07328f
.ends

