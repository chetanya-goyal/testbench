* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t19 plus.t0 drain_left.t7 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 source.t18 plus.t1 drain_left.t9 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 source.t1 minus.t0 drain_right.t9 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X3 source.t0 minus.t1 drain_right.t8 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X4 drain_left.t3 plus.t2 source.t17 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X5 source.t16 plus.t3 drain_left.t4 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X6 a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X7 drain_left.t5 plus.t4 source.t15 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X8 drain_left.t0 plus.t5 source.t14 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X9 drain_left.t8 plus.t6 source.t13 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X10 drain_left.t1 plus.t7 source.t12 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X11 drain_left.t6 plus.t8 source.t11 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X12 a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X13 source.t10 plus.t9 drain_left.t2 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X14 drain_right.t7 minus.t2 source.t3 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X15 drain_right.t6 minus.t3 source.t6 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X16 source.t8 minus.t4 drain_right.t5 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X17 source.t7 minus.t5 drain_right.t4 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 drain_right.t3 minus.t6 source.t2 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X19 drain_right.t2 minus.t7 source.t4 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X20 a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X21 a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X22 drain_right.t1 minus.t8 source.t5 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X23 drain_right.t0 minus.t9 source.t9 a_n1412_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n2 plus.t2 474.406
R1 plus.n8 plus.t7 474.406
R2 plus.n12 plus.t5 474.406
R3 plus.n18 plus.t4 474.406
R4 plus.n1 plus.t1 414.521
R5 plus.n5 plus.t8 414.521
R6 plus.n7 plus.t0 414.521
R7 plus.n11 plus.t3 414.521
R8 plus.n15 plus.t6 414.521
R9 plus.n17 plus.t9 414.521
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 24.9574
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 8.7505
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n5 drain_left.t3 86.8731
R37 drain_left.n1 drain_left.t5 86.873
R38 drain_left.n3 drain_left.n2 80.0927
R39 drain_left.n7 drain_left.n6 79.7731
R40 drain_left.n5 drain_left.n4 79.7731
R41 drain_left.n1 drain_left.n0 79.773
R42 drain_left drain_left.n3 22.6739
R43 drain_left.n2 drain_left.t4 6.6005
R44 drain_left.n2 drain_left.t0 6.6005
R45 drain_left.n0 drain_left.t2 6.6005
R46 drain_left.n0 drain_left.t8 6.6005
R47 drain_left.n6 drain_left.t7 6.6005
R48 drain_left.n6 drain_left.t1 6.6005
R49 drain_left.n4 drain_left.t9 6.6005
R50 drain_left.n4 drain_left.t6 6.6005
R51 drain_left drain_left.n7 6.15322
R52 drain_left.n7 drain_left.n5 0.5005
R53 drain_left.n3 drain_left.n1 0.070154
R54 source.n0 source.t12 69.6943
R55 source.n5 source.t6 69.6943
R56 source.n19 source.t5 69.6942
R57 source.n14 source.t14 69.6942
R58 source.n2 source.n1 63.0943
R59 source.n4 source.n3 63.0943
R60 source.n7 source.n6 63.0943
R61 source.n9 source.n8 63.0943
R62 source.n18 source.n17 63.0942
R63 source.n16 source.n15 63.0942
R64 source.n13 source.n12 63.0942
R65 source.n11 source.n10 63.0942
R66 source.n11 source.n9 15.4695
R67 source.n20 source.n0 9.45661
R68 source.n17 source.t2 6.6005
R69 source.n17 source.t7 6.6005
R70 source.n15 source.t9 6.6005
R71 source.n15 source.t8 6.6005
R72 source.n12 source.t13 6.6005
R73 source.n12 source.t16 6.6005
R74 source.n10 source.t15 6.6005
R75 source.n10 source.t10 6.6005
R76 source.n1 source.t11 6.6005
R77 source.n1 source.t19 6.6005
R78 source.n3 source.t17 6.6005
R79 source.n3 source.t18 6.6005
R80 source.n6 source.t3 6.6005
R81 source.n6 source.t0 6.6005
R82 source.n8 source.t4 6.6005
R83 source.n8 source.t1 6.6005
R84 source.n20 source.n19 5.51343
R85 source.n5 source.n4 0.720328
R86 source.n16 source.n14 0.720328
R87 source.n9 source.n7 0.5005
R88 source.n7 source.n5 0.5005
R89 source.n4 source.n2 0.5005
R90 source.n2 source.n0 0.5005
R91 source.n13 source.n11 0.5005
R92 source.n14 source.n13 0.5005
R93 source.n18 source.n16 0.5005
R94 source.n19 source.n18 0.5005
R95 source source.n20 0.188
R96 minus.n8 minus.t7 474.406
R97 minus.n2 minus.t3 474.406
R98 minus.n18 minus.t8 474.406
R99 minus.n12 minus.t9 474.406
R100 minus.n7 minus.t0 414.521
R101 minus.n5 minus.t2 414.521
R102 minus.n1 minus.t1 414.521
R103 minus.n17 minus.t5 414.521
R104 minus.n15 minus.t6 414.521
R105 minus.n11 minus.t4 414.521
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 48.2005
R115 minus.n4 minus.n1 48.2005
R116 minus.n14 minus.n11 48.2005
R117 minus.n17 minus.n16 48.2005
R118 minus.n6 minus.n5 36.5157
R119 minus.n5 minus.n4 36.5157
R120 minus.n15 minus.n14 36.5157
R121 minus.n16 minus.n15 36.5157
R122 minus.n20 minus.n9 27.6672
R123 minus.n8 minus.n7 24.8308
R124 minus.n2 minus.n1 24.8308
R125 minus.n12 minus.n11 24.8308
R126 minus.n18 minus.n17 24.8308
R127 minus.n20 minus.n19 6.51565
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t0 86.873
R134 drain_right.n7 drain_right.t2 86.3731
R135 drain_right.n6 drain_right.n4 80.2731
R136 drain_right.n3 drain_right.n2 80.0927
R137 drain_right.n6 drain_right.n5 79.7731
R138 drain_right.n1 drain_right.n0 79.773
R139 drain_right drain_right.n3 22.1207
R140 drain_right.n2 drain_right.t4 6.6005
R141 drain_right.n2 drain_right.t1 6.6005
R142 drain_right.n0 drain_right.t5 6.6005
R143 drain_right.n0 drain_right.t3 6.6005
R144 drain_right.n4 drain_right.t8 6.6005
R145 drain_right.n4 drain_right.t6 6.6005
R146 drain_right.n5 drain_right.t9 6.6005
R147 drain_right.n5 drain_right.t7 6.6005
R148 drain_right drain_right.n7 5.90322
R149 drain_right.n7 drain_right.n6 0.5005
R150 drain_right.n3 drain_right.n1 0.070154
C0 plus source 1.22077f
C1 drain_left minus 0.176151f
C2 drain_right minus 1.17714f
C3 drain_left source 7.27319f
C4 drain_right source 7.26904f
C5 drain_left plus 1.31057f
C6 drain_right plus 0.294086f
C7 drain_left drain_right 0.690178f
C8 minus source 1.20661f
C9 plus minus 3.24993f
C10 drain_right a_n1412_n1488# 3.84388f
C11 drain_left a_n1412_n1488# 4.05153f
C12 source a_n1412_n1488# 2.775574f
C13 minus a_n1412_n1488# 4.726942f
C14 plus a_n1412_n1488# 5.409138f
C15 drain_right.t0 a_n1412_n1488# 0.565964f
C16 drain_right.t5 a_n1412_n1488# 0.060959f
C17 drain_right.t3 a_n1412_n1488# 0.060959f
C18 drain_right.n0 a_n1412_n1488# 0.43963f
C19 drain_right.n1 a_n1412_n1488# 0.559125f
C20 drain_right.t4 a_n1412_n1488# 0.060959f
C21 drain_right.t1 a_n1412_n1488# 0.060959f
C22 drain_right.n2 a_n1412_n1488# 0.440771f
C23 drain_right.n3 a_n1412_n1488# 0.893396f
C24 drain_right.t8 a_n1412_n1488# 0.060959f
C25 drain_right.t6 a_n1412_n1488# 0.060959f
C26 drain_right.n4 a_n1412_n1488# 0.441494f
C27 drain_right.t9 a_n1412_n1488# 0.060959f
C28 drain_right.t7 a_n1412_n1488# 0.060959f
C29 drain_right.n5 a_n1412_n1488# 0.439632f
C30 drain_right.n6 a_n1412_n1488# 0.585866f
C31 drain_right.t2 a_n1412_n1488# 0.564244f
C32 drain_right.n7 a_n1412_n1488# 0.511013f
C33 minus.n0 a_n1412_n1488# 0.031144f
C34 minus.t7 a_n1412_n1488# 0.07319f
C35 minus.t0 a_n1412_n1488# 0.067642f
C36 minus.t2 a_n1412_n1488# 0.067642f
C37 minus.t1 a_n1412_n1488# 0.067642f
C38 minus.n1 a_n1412_n1488# 0.040876f
C39 minus.t3 a_n1412_n1488# 0.07319f
C40 minus.n2 a_n1412_n1488# 0.050318f
C41 minus.n3 a_n1412_n1488# 0.073183f
C42 minus.n4 a_n1412_n1488# 0.011868f
C43 minus.n5 a_n1412_n1488# 0.040876f
C44 minus.n6 a_n1412_n1488# 0.011868f
C45 minus.n7 a_n1412_n1488# 0.040876f
C46 minus.n8 a_n1412_n1488# 0.050268f
C47 minus.n9 a_n1412_n1488# 0.704001f
C48 minus.n10 a_n1412_n1488# 0.031144f
C49 minus.t5 a_n1412_n1488# 0.067642f
C50 minus.t6 a_n1412_n1488# 0.067642f
C51 minus.t4 a_n1412_n1488# 0.067642f
C52 minus.n11 a_n1412_n1488# 0.040876f
C53 minus.t9 a_n1412_n1488# 0.07319f
C54 minus.n12 a_n1412_n1488# 0.050318f
C55 minus.n13 a_n1412_n1488# 0.073183f
C56 minus.n14 a_n1412_n1488# 0.011868f
C57 minus.n15 a_n1412_n1488# 0.040876f
C58 minus.n16 a_n1412_n1488# 0.011868f
C59 minus.n17 a_n1412_n1488# 0.040876f
C60 minus.t8 a_n1412_n1488# 0.07319f
C61 minus.n18 a_n1412_n1488# 0.050268f
C62 minus.n19 a_n1412_n1488# 0.204759f
C63 minus.n20 a_n1412_n1488# 0.869623f
C64 source.t12 a_n1412_n1488# 0.587924f
C65 source.n0 a_n1412_n1488# 0.794817f
C66 source.t11 a_n1412_n1488# 0.070802f
C67 source.t19 a_n1412_n1488# 0.070802f
C68 source.n1 a_n1412_n1488# 0.448923f
C69 source.n2 a_n1412_n1488# 0.356399f
C70 source.t17 a_n1412_n1488# 0.070802f
C71 source.t18 a_n1412_n1488# 0.070802f
C72 source.n3 a_n1412_n1488# 0.448923f
C73 source.n4 a_n1412_n1488# 0.377553f
C74 source.t6 a_n1412_n1488# 0.587924f
C75 source.n5 a_n1412_n1488# 0.431648f
C76 source.t3 a_n1412_n1488# 0.070802f
C77 source.t0 a_n1412_n1488# 0.070802f
C78 source.n6 a_n1412_n1488# 0.448923f
C79 source.n7 a_n1412_n1488# 0.356399f
C80 source.t4 a_n1412_n1488# 0.070802f
C81 source.t1 a_n1412_n1488# 0.070802f
C82 source.n8 a_n1412_n1488# 0.448923f
C83 source.n9 a_n1412_n1488# 1.09916f
C84 source.t15 a_n1412_n1488# 0.070802f
C85 source.t10 a_n1412_n1488# 0.070802f
C86 source.n10 a_n1412_n1488# 0.448919f
C87 source.n11 a_n1412_n1488# 1.09916f
C88 source.t13 a_n1412_n1488# 0.070802f
C89 source.t16 a_n1412_n1488# 0.070802f
C90 source.n12 a_n1412_n1488# 0.448919f
C91 source.n13 a_n1412_n1488# 0.356402f
C92 source.t14 a_n1412_n1488# 0.587921f
C93 source.n14 a_n1412_n1488# 0.431651f
C94 source.t9 a_n1412_n1488# 0.070802f
C95 source.t8 a_n1412_n1488# 0.070802f
C96 source.n15 a_n1412_n1488# 0.448919f
C97 source.n16 a_n1412_n1488# 0.377557f
C98 source.t2 a_n1412_n1488# 0.070802f
C99 source.t7 a_n1412_n1488# 0.070802f
C100 source.n17 a_n1412_n1488# 0.448919f
C101 source.n18 a_n1412_n1488# 0.356402f
C102 source.t5 a_n1412_n1488# 0.587921f
C103 source.n19 a_n1412_n1488# 0.572862f
C104 source.n20 a_n1412_n1488# 0.863837f
C105 drain_left.t5 a_n1412_n1488# 0.558272f
C106 drain_left.t2 a_n1412_n1488# 0.06013f
C107 drain_left.t8 a_n1412_n1488# 0.06013f
C108 drain_left.n0 a_n1412_n1488# 0.433654f
C109 drain_left.n1 a_n1412_n1488# 0.551525f
C110 drain_left.t4 a_n1412_n1488# 0.06013f
C111 drain_left.t0 a_n1412_n1488# 0.06013f
C112 drain_left.n2 a_n1412_n1488# 0.43478f
C113 drain_left.n3 a_n1412_n1488# 0.931787f
C114 drain_left.t3 a_n1412_n1488# 0.558274f
C115 drain_left.t9 a_n1412_n1488# 0.06013f
C116 drain_left.t6 a_n1412_n1488# 0.06013f
C117 drain_left.n4 a_n1412_n1488# 0.433656f
C118 drain_left.n5 a_n1412_n1488# 0.578251f
C119 drain_left.t7 a_n1412_n1488# 0.06013f
C120 drain_left.t1 a_n1412_n1488# 0.06013f
C121 drain_left.n6 a_n1412_n1488# 0.433656f
C122 drain_left.n7 a_n1412_n1488# 0.494126f
C123 plus.n0 a_n1412_n1488# 0.031769f
C124 plus.t0 a_n1412_n1488# 0.069f
C125 plus.t8 a_n1412_n1488# 0.069f
C126 plus.t1 a_n1412_n1488# 0.069f
C127 plus.n1 a_n1412_n1488# 0.041697f
C128 plus.t2 a_n1412_n1488# 0.074659f
C129 plus.n2 a_n1412_n1488# 0.051328f
C130 plus.n3 a_n1412_n1488# 0.074653f
C131 plus.n4 a_n1412_n1488# 0.012106f
C132 plus.n5 a_n1412_n1488# 0.041697f
C133 plus.n6 a_n1412_n1488# 0.012106f
C134 plus.n7 a_n1412_n1488# 0.041697f
C135 plus.t7 a_n1412_n1488# 0.074659f
C136 plus.n8 a_n1412_n1488# 0.051278f
C137 plus.n9 a_n1412_n1488# 0.238545f
C138 plus.n10 a_n1412_n1488# 0.031769f
C139 plus.t4 a_n1412_n1488# 0.074659f
C140 plus.t9 a_n1412_n1488# 0.069f
C141 plus.t6 a_n1412_n1488# 0.069f
C142 plus.t3 a_n1412_n1488# 0.069f
C143 plus.n11 a_n1412_n1488# 0.041697f
C144 plus.t5 a_n1412_n1488# 0.074659f
C145 plus.n12 a_n1412_n1488# 0.051328f
C146 plus.n13 a_n1412_n1488# 0.074653f
C147 plus.n14 a_n1412_n1488# 0.012106f
C148 plus.n15 a_n1412_n1488# 0.041697f
C149 plus.n16 a_n1412_n1488# 0.012106f
C150 plus.n17 a_n1412_n1488# 0.041697f
C151 plus.n18 a_n1412_n1488# 0.051278f
C152 plus.n19 a_n1412_n1488# 0.678071f
.ends

