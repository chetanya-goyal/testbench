* NGSPICE file created from diffpair278.ext - technology: sky130A

.subckt diffpair278 minus drain_right drain_left source plus
X0 source.t39 minus.t0 drain_right.t9 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t38 minus.t1 drain_right.t2 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X3 drain_left.t19 plus.t0 source.t15 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X4 source.t37 minus.t2 drain_right.t1 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X5 drain_right.t0 minus.t3 source.t36 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X6 drain_right.t12 minus.t4 source.t35 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 source.t2 plus.t1 drain_left.t18 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X8 source.t8 plus.t2 drain_left.t17 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X9 source.t1 plus.t3 drain_left.t16 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 source.t5 plus.t4 drain_left.t15 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X11 a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X12 drain_right.t14 minus.t5 source.t34 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X13 drain_right.t7 minus.t6 source.t33 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 drain_right.t6 minus.t7 source.t32 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X15 source.t31 minus.t8 drain_right.t18 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X16 source.t30 minus.t9 drain_right.t17 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X17 a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X18 drain_right.t16 minus.t10 source.t29 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X19 source.t3 plus.t5 drain_left.t14 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X20 source.t16 plus.t6 drain_left.t13 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X21 drain_right.t8 minus.t11 source.t28 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X22 source.t10 plus.t7 drain_left.t12 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X23 drain_left.t11 plus.t8 source.t9 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X24 drain_left.t10 plus.t9 source.t18 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X25 drain_left.t9 plus.t10 source.t19 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X26 source.t27 minus.t12 drain_right.t19 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X27 a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X28 source.t4 plus.t11 drain_left.t8 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X29 drain_right.t10 minus.t13 source.t26 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X30 drain_left.t7 plus.t12 source.t0 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X31 source.t25 minus.t14 drain_right.t11 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X32 source.t24 minus.t15 drain_right.t4 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X33 source.t17 plus.t13 drain_left.t6 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X34 drain_right.t5 minus.t16 source.t23 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X35 drain_left.t5 plus.t14 source.t12 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X36 drain_left.t4 plus.t15 source.t14 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X37 drain_right.t3 minus.t17 source.t22 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X38 drain_left.t3 plus.t16 source.t7 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X39 drain_left.t2 plus.t17 source.t11 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X40 source.t21 minus.t18 drain_right.t13 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X41 source.t20 minus.t19 drain_right.t15 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X42 source.t13 plus.t18 drain_left.t1 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X43 drain_left.t0 plus.t19 source.t6 a_n2102_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n27 minus.t8 635.365
R1 minus.n7 minus.t13 635.365
R2 minus.n56 minus.t16 635.365
R3 minus.n35 minus.t15 635.365
R4 minus.n26 minus.t4 586.433
R5 minus.n24 minus.t19 586.433
R6 minus.n3 minus.t5 586.433
R7 minus.n18 minus.t2 586.433
R8 minus.n16 minus.t17 586.433
R9 minus.n4 minus.t12 586.433
R10 minus.n10 minus.t3 586.433
R11 minus.n6 minus.t18 586.433
R12 minus.n55 minus.t9 586.433
R13 minus.n53 minus.t10 586.433
R14 minus.n47 minus.t0 586.433
R15 minus.n46 minus.t11 586.433
R16 minus.n44 minus.t1 586.433
R17 minus.n32 minus.t6 586.433
R18 minus.n38 minus.t14 586.433
R19 minus.n34 minus.t7 586.433
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 64.9975
R47 minus.n15 minus.n4 64.9975
R48 minus.n43 minus.n32 64.9975
R49 minus.n48 minus.n47 64.9975
R50 minus.n25 minus.n24 62.0763
R51 minus.n10 minus.n9 62.0763
R52 minus.n38 minus.n37 62.0763
R53 minus.n54 minus.n53 62.0763
R54 minus.n18 minus.n17 46.0096
R55 minus.n17 minus.n16 46.0096
R56 minus.n45 minus.n44 46.0096
R57 minus.n46 minus.n45 46.0096
R58 minus.n27 minus.n26 43.0884
R59 minus.n7 minus.n6 43.0884
R60 minus.n35 minus.n34 43.0884
R61 minus.n56 minus.n55 43.0884
R62 minus.n58 minus.n28 32.5535
R63 minus.n26 minus.n25 29.9429
R64 minus.n9 minus.n6 29.9429
R65 minus.n37 minus.n34 29.9429
R66 minus.n55 minus.n54 29.9429
R67 minus.n19 minus.n18 27.0217
R68 minus.n16 minus.n15 27.0217
R69 minus.n44 minus.n43 27.0217
R70 minus.n48 minus.n46 27.0217
R71 minus.n24 minus.n23 10.955
R72 minus.n11 minus.n10 10.955
R73 minus.n39 minus.n38 10.955
R74 minus.n53 minus.n52 10.955
R75 minus.n3 minus.n1 8.03383
R76 minus.n12 minus.n4 8.03383
R77 minus.n40 minus.n32 8.03383
R78 minus.n47 minus.n30 8.03383
R79 minus.n58 minus.n57 6.51565
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 drain_right.n6 drain_right.n4 67.7338
R100 drain_right.n2 drain_right.n0 67.7338
R101 drain_right.n10 drain_right.n8 67.7338
R102 drain_right.n10 drain_right.n9 67.1908
R103 drain_right.n12 drain_right.n11 67.1908
R104 drain_right.n14 drain_right.n13 67.1908
R105 drain_right.n16 drain_right.n15 67.1908
R106 drain_right.n7 drain_right.n3 67.1907
R107 drain_right.n6 drain_right.n5 67.1907
R108 drain_right.n2 drain_right.n1 67.1907
R109 drain_right drain_right.n7 26.6132
R110 drain_right drain_right.n16 6.19632
R111 drain_right.n3 drain_right.t2 3.3005
R112 drain_right.n3 drain_right.t8 3.3005
R113 drain_right.n4 drain_right.t17 3.3005
R114 drain_right.n4 drain_right.t5 3.3005
R115 drain_right.n5 drain_right.t9 3.3005
R116 drain_right.n5 drain_right.t16 3.3005
R117 drain_right.n1 drain_right.t11 3.3005
R118 drain_right.n1 drain_right.t7 3.3005
R119 drain_right.n0 drain_right.t4 3.3005
R120 drain_right.n0 drain_right.t6 3.3005
R121 drain_right.n8 drain_right.t13 3.3005
R122 drain_right.n8 drain_right.t10 3.3005
R123 drain_right.n9 drain_right.t19 3.3005
R124 drain_right.n9 drain_right.t0 3.3005
R125 drain_right.n11 drain_right.t1 3.3005
R126 drain_right.n11 drain_right.t3 3.3005
R127 drain_right.n13 drain_right.t15 3.3005
R128 drain_right.n13 drain_right.t14 3.3005
R129 drain_right.n15 drain_right.t18 3.3005
R130 drain_right.n15 drain_right.t12 3.3005
R131 drain_right.n16 drain_right.n14 0.543603
R132 drain_right.n14 drain_right.n12 0.543603
R133 drain_right.n12 drain_right.n10 0.543603
R134 drain_right.n7 drain_right.n6 0.488257
R135 drain_right.n7 drain_right.n2 0.488257
R136 source.n282 source.n256 289.615
R137 source.n242 source.n216 289.615
R138 source.n210 source.n184 289.615
R139 source.n170 source.n144 289.615
R140 source.n26 source.n0 289.615
R141 source.n66 source.n40 289.615
R142 source.n98 source.n72 289.615
R143 source.n138 source.n112 289.615
R144 source.n267 source.n266 185
R145 source.n264 source.n263 185
R146 source.n273 source.n272 185
R147 source.n275 source.n274 185
R148 source.n260 source.n259 185
R149 source.n281 source.n280 185
R150 source.n283 source.n282 185
R151 source.n227 source.n226 185
R152 source.n224 source.n223 185
R153 source.n233 source.n232 185
R154 source.n235 source.n234 185
R155 source.n220 source.n219 185
R156 source.n241 source.n240 185
R157 source.n243 source.n242 185
R158 source.n195 source.n194 185
R159 source.n192 source.n191 185
R160 source.n201 source.n200 185
R161 source.n203 source.n202 185
R162 source.n188 source.n187 185
R163 source.n209 source.n208 185
R164 source.n211 source.n210 185
R165 source.n155 source.n154 185
R166 source.n152 source.n151 185
R167 source.n161 source.n160 185
R168 source.n163 source.n162 185
R169 source.n148 source.n147 185
R170 source.n169 source.n168 185
R171 source.n171 source.n170 185
R172 source.n27 source.n26 185
R173 source.n25 source.n24 185
R174 source.n4 source.n3 185
R175 source.n19 source.n18 185
R176 source.n17 source.n16 185
R177 source.n8 source.n7 185
R178 source.n11 source.n10 185
R179 source.n67 source.n66 185
R180 source.n65 source.n64 185
R181 source.n44 source.n43 185
R182 source.n59 source.n58 185
R183 source.n57 source.n56 185
R184 source.n48 source.n47 185
R185 source.n51 source.n50 185
R186 source.n99 source.n98 185
R187 source.n97 source.n96 185
R188 source.n76 source.n75 185
R189 source.n91 source.n90 185
R190 source.n89 source.n88 185
R191 source.n80 source.n79 185
R192 source.n83 source.n82 185
R193 source.n139 source.n138 185
R194 source.n137 source.n136 185
R195 source.n116 source.n115 185
R196 source.n131 source.n130 185
R197 source.n129 source.n128 185
R198 source.n120 source.n119 185
R199 source.n123 source.n122 185
R200 source.t23 source.n265 147.661
R201 source.t24 source.n225 147.661
R202 source.t18 source.n193 147.661
R203 source.t16 source.n153 147.661
R204 source.t14 source.n9 147.661
R205 source.t8 source.n49 147.661
R206 source.t26 source.n81 147.661
R207 source.t31 source.n121 147.661
R208 source.n266 source.n263 104.615
R209 source.n273 source.n263 104.615
R210 source.n274 source.n273 104.615
R211 source.n274 source.n259 104.615
R212 source.n281 source.n259 104.615
R213 source.n282 source.n281 104.615
R214 source.n226 source.n223 104.615
R215 source.n233 source.n223 104.615
R216 source.n234 source.n233 104.615
R217 source.n234 source.n219 104.615
R218 source.n241 source.n219 104.615
R219 source.n242 source.n241 104.615
R220 source.n194 source.n191 104.615
R221 source.n201 source.n191 104.615
R222 source.n202 source.n201 104.615
R223 source.n202 source.n187 104.615
R224 source.n209 source.n187 104.615
R225 source.n210 source.n209 104.615
R226 source.n154 source.n151 104.615
R227 source.n161 source.n151 104.615
R228 source.n162 source.n161 104.615
R229 source.n162 source.n147 104.615
R230 source.n169 source.n147 104.615
R231 source.n170 source.n169 104.615
R232 source.n26 source.n25 104.615
R233 source.n25 source.n3 104.615
R234 source.n18 source.n3 104.615
R235 source.n18 source.n17 104.615
R236 source.n17 source.n7 104.615
R237 source.n10 source.n7 104.615
R238 source.n66 source.n65 104.615
R239 source.n65 source.n43 104.615
R240 source.n58 source.n43 104.615
R241 source.n58 source.n57 104.615
R242 source.n57 source.n47 104.615
R243 source.n50 source.n47 104.615
R244 source.n98 source.n97 104.615
R245 source.n97 source.n75 104.615
R246 source.n90 source.n75 104.615
R247 source.n90 source.n89 104.615
R248 source.n89 source.n79 104.615
R249 source.n82 source.n79 104.615
R250 source.n138 source.n137 104.615
R251 source.n137 source.n115 104.615
R252 source.n130 source.n115 104.615
R253 source.n130 source.n129 104.615
R254 source.n129 source.n119 104.615
R255 source.n122 source.n119 104.615
R256 source.n266 source.t23 52.3082
R257 source.n226 source.t24 52.3082
R258 source.n194 source.t18 52.3082
R259 source.n154 source.t16 52.3082
R260 source.n10 source.t14 52.3082
R261 source.n50 source.t8 52.3082
R262 source.n82 source.t26 52.3082
R263 source.n122 source.t31 52.3082
R264 source.n33 source.n32 50.512
R265 source.n35 source.n34 50.512
R266 source.n37 source.n36 50.512
R267 source.n39 source.n38 50.512
R268 source.n105 source.n104 50.512
R269 source.n107 source.n106 50.512
R270 source.n109 source.n108 50.512
R271 source.n111 source.n110 50.512
R272 source.n255 source.n254 50.5119
R273 source.n253 source.n252 50.5119
R274 source.n251 source.n250 50.5119
R275 source.n249 source.n248 50.5119
R276 source.n183 source.n182 50.5119
R277 source.n181 source.n180 50.5119
R278 source.n179 source.n178 50.5119
R279 source.n177 source.n176 50.5119
R280 source.n287 source.n286 32.1853
R281 source.n247 source.n246 32.1853
R282 source.n215 source.n214 32.1853
R283 source.n175 source.n174 32.1853
R284 source.n31 source.n30 32.1853
R285 source.n71 source.n70 32.1853
R286 source.n103 source.n102 32.1853
R287 source.n143 source.n142 32.1853
R288 source.n175 source.n143 17.2854
R289 source.n267 source.n265 15.6674
R290 source.n227 source.n225 15.6674
R291 source.n195 source.n193 15.6674
R292 source.n155 source.n153 15.6674
R293 source.n11 source.n9 15.6674
R294 source.n51 source.n49 15.6674
R295 source.n83 source.n81 15.6674
R296 source.n123 source.n121 15.6674
R297 source.n268 source.n264 12.8005
R298 source.n228 source.n224 12.8005
R299 source.n196 source.n192 12.8005
R300 source.n156 source.n152 12.8005
R301 source.n12 source.n8 12.8005
R302 source.n52 source.n48 12.8005
R303 source.n84 source.n80 12.8005
R304 source.n124 source.n120 12.8005
R305 source.n272 source.n271 12.0247
R306 source.n232 source.n231 12.0247
R307 source.n200 source.n199 12.0247
R308 source.n160 source.n159 12.0247
R309 source.n16 source.n15 12.0247
R310 source.n56 source.n55 12.0247
R311 source.n88 source.n87 12.0247
R312 source.n128 source.n127 12.0247
R313 source.n288 source.n31 11.7509
R314 source.n275 source.n262 11.249
R315 source.n235 source.n222 11.249
R316 source.n203 source.n190 11.249
R317 source.n163 source.n150 11.249
R318 source.n19 source.n6 11.249
R319 source.n59 source.n46 11.249
R320 source.n91 source.n78 11.249
R321 source.n131 source.n118 11.249
R322 source.n276 source.n260 10.4732
R323 source.n236 source.n220 10.4732
R324 source.n204 source.n188 10.4732
R325 source.n164 source.n148 10.4732
R326 source.n20 source.n4 10.4732
R327 source.n60 source.n44 10.4732
R328 source.n92 source.n76 10.4732
R329 source.n132 source.n116 10.4732
R330 source.n280 source.n279 9.69747
R331 source.n240 source.n239 9.69747
R332 source.n208 source.n207 9.69747
R333 source.n168 source.n167 9.69747
R334 source.n24 source.n23 9.69747
R335 source.n64 source.n63 9.69747
R336 source.n96 source.n95 9.69747
R337 source.n136 source.n135 9.69747
R338 source.n286 source.n285 9.45567
R339 source.n246 source.n245 9.45567
R340 source.n214 source.n213 9.45567
R341 source.n174 source.n173 9.45567
R342 source.n30 source.n29 9.45567
R343 source.n70 source.n69 9.45567
R344 source.n102 source.n101 9.45567
R345 source.n142 source.n141 9.45567
R346 source.n285 source.n284 9.3005
R347 source.n258 source.n257 9.3005
R348 source.n279 source.n278 9.3005
R349 source.n277 source.n276 9.3005
R350 source.n262 source.n261 9.3005
R351 source.n271 source.n270 9.3005
R352 source.n269 source.n268 9.3005
R353 source.n245 source.n244 9.3005
R354 source.n218 source.n217 9.3005
R355 source.n239 source.n238 9.3005
R356 source.n237 source.n236 9.3005
R357 source.n222 source.n221 9.3005
R358 source.n231 source.n230 9.3005
R359 source.n229 source.n228 9.3005
R360 source.n213 source.n212 9.3005
R361 source.n186 source.n185 9.3005
R362 source.n207 source.n206 9.3005
R363 source.n205 source.n204 9.3005
R364 source.n190 source.n189 9.3005
R365 source.n199 source.n198 9.3005
R366 source.n197 source.n196 9.3005
R367 source.n173 source.n172 9.3005
R368 source.n146 source.n145 9.3005
R369 source.n167 source.n166 9.3005
R370 source.n165 source.n164 9.3005
R371 source.n150 source.n149 9.3005
R372 source.n159 source.n158 9.3005
R373 source.n157 source.n156 9.3005
R374 source.n29 source.n28 9.3005
R375 source.n2 source.n1 9.3005
R376 source.n23 source.n22 9.3005
R377 source.n21 source.n20 9.3005
R378 source.n6 source.n5 9.3005
R379 source.n15 source.n14 9.3005
R380 source.n13 source.n12 9.3005
R381 source.n69 source.n68 9.3005
R382 source.n42 source.n41 9.3005
R383 source.n63 source.n62 9.3005
R384 source.n61 source.n60 9.3005
R385 source.n46 source.n45 9.3005
R386 source.n55 source.n54 9.3005
R387 source.n53 source.n52 9.3005
R388 source.n101 source.n100 9.3005
R389 source.n74 source.n73 9.3005
R390 source.n95 source.n94 9.3005
R391 source.n93 source.n92 9.3005
R392 source.n78 source.n77 9.3005
R393 source.n87 source.n86 9.3005
R394 source.n85 source.n84 9.3005
R395 source.n141 source.n140 9.3005
R396 source.n114 source.n113 9.3005
R397 source.n135 source.n134 9.3005
R398 source.n133 source.n132 9.3005
R399 source.n118 source.n117 9.3005
R400 source.n127 source.n126 9.3005
R401 source.n125 source.n124 9.3005
R402 source.n283 source.n258 8.92171
R403 source.n243 source.n218 8.92171
R404 source.n211 source.n186 8.92171
R405 source.n171 source.n146 8.92171
R406 source.n27 source.n2 8.92171
R407 source.n67 source.n42 8.92171
R408 source.n99 source.n74 8.92171
R409 source.n139 source.n114 8.92171
R410 source.n284 source.n256 8.14595
R411 source.n244 source.n216 8.14595
R412 source.n212 source.n184 8.14595
R413 source.n172 source.n144 8.14595
R414 source.n28 source.n0 8.14595
R415 source.n68 source.n40 8.14595
R416 source.n100 source.n72 8.14595
R417 source.n140 source.n112 8.14595
R418 source.n286 source.n256 5.81868
R419 source.n246 source.n216 5.81868
R420 source.n214 source.n184 5.81868
R421 source.n174 source.n144 5.81868
R422 source.n30 source.n0 5.81868
R423 source.n70 source.n40 5.81868
R424 source.n102 source.n72 5.81868
R425 source.n142 source.n112 5.81868
R426 source.n288 source.n287 5.53498
R427 source.n284 source.n283 5.04292
R428 source.n244 source.n243 5.04292
R429 source.n212 source.n211 5.04292
R430 source.n172 source.n171 5.04292
R431 source.n28 source.n27 5.04292
R432 source.n68 source.n67 5.04292
R433 source.n100 source.n99 5.04292
R434 source.n140 source.n139 5.04292
R435 source.n269 source.n265 4.38594
R436 source.n229 source.n225 4.38594
R437 source.n197 source.n193 4.38594
R438 source.n157 source.n153 4.38594
R439 source.n13 source.n9 4.38594
R440 source.n53 source.n49 4.38594
R441 source.n85 source.n81 4.38594
R442 source.n125 source.n121 4.38594
R443 source.n280 source.n258 4.26717
R444 source.n240 source.n218 4.26717
R445 source.n208 source.n186 4.26717
R446 source.n168 source.n146 4.26717
R447 source.n24 source.n2 4.26717
R448 source.n64 source.n42 4.26717
R449 source.n96 source.n74 4.26717
R450 source.n136 source.n114 4.26717
R451 source.n279 source.n260 3.49141
R452 source.n239 source.n220 3.49141
R453 source.n207 source.n188 3.49141
R454 source.n167 source.n148 3.49141
R455 source.n23 source.n4 3.49141
R456 source.n63 source.n44 3.49141
R457 source.n95 source.n76 3.49141
R458 source.n135 source.n116 3.49141
R459 source.n254 source.t29 3.3005
R460 source.n254 source.t30 3.3005
R461 source.n252 source.t28 3.3005
R462 source.n252 source.t39 3.3005
R463 source.n250 source.t33 3.3005
R464 source.n250 source.t38 3.3005
R465 source.n248 source.t32 3.3005
R466 source.n248 source.t25 3.3005
R467 source.n182 source.t19 3.3005
R468 source.n182 source.t2 3.3005
R469 source.n180 source.t7 3.3005
R470 source.n180 source.t1 3.3005
R471 source.n178 source.t11 3.3005
R472 source.n178 source.t5 3.3005
R473 source.n176 source.t12 3.3005
R474 source.n176 source.t3 3.3005
R475 source.n32 source.t15 3.3005
R476 source.n32 source.t4 3.3005
R477 source.n34 source.t0 3.3005
R478 source.n34 source.t13 3.3005
R479 source.n36 source.t6 3.3005
R480 source.n36 source.t10 3.3005
R481 source.n38 source.t9 3.3005
R482 source.n38 source.t17 3.3005
R483 source.n104 source.t36 3.3005
R484 source.n104 source.t21 3.3005
R485 source.n106 source.t22 3.3005
R486 source.n106 source.t27 3.3005
R487 source.n108 source.t34 3.3005
R488 source.n108 source.t37 3.3005
R489 source.n110 source.t35 3.3005
R490 source.n110 source.t20 3.3005
R491 source.n276 source.n275 2.71565
R492 source.n236 source.n235 2.71565
R493 source.n204 source.n203 2.71565
R494 source.n164 source.n163 2.71565
R495 source.n20 source.n19 2.71565
R496 source.n60 source.n59 2.71565
R497 source.n92 source.n91 2.71565
R498 source.n132 source.n131 2.71565
R499 source.n272 source.n262 1.93989
R500 source.n232 source.n222 1.93989
R501 source.n200 source.n190 1.93989
R502 source.n160 source.n150 1.93989
R503 source.n16 source.n6 1.93989
R504 source.n56 source.n46 1.93989
R505 source.n88 source.n78 1.93989
R506 source.n128 source.n118 1.93989
R507 source.n271 source.n264 1.16414
R508 source.n231 source.n224 1.16414
R509 source.n199 source.n192 1.16414
R510 source.n159 source.n152 1.16414
R511 source.n15 source.n8 1.16414
R512 source.n55 source.n48 1.16414
R513 source.n87 source.n80 1.16414
R514 source.n127 source.n120 1.16414
R515 source.n143 source.n111 0.543603
R516 source.n111 source.n109 0.543603
R517 source.n109 source.n107 0.543603
R518 source.n107 source.n105 0.543603
R519 source.n105 source.n103 0.543603
R520 source.n71 source.n39 0.543603
R521 source.n39 source.n37 0.543603
R522 source.n37 source.n35 0.543603
R523 source.n35 source.n33 0.543603
R524 source.n33 source.n31 0.543603
R525 source.n177 source.n175 0.543603
R526 source.n179 source.n177 0.543603
R527 source.n181 source.n179 0.543603
R528 source.n183 source.n181 0.543603
R529 source.n215 source.n183 0.543603
R530 source.n249 source.n247 0.543603
R531 source.n251 source.n249 0.543603
R532 source.n253 source.n251 0.543603
R533 source.n255 source.n253 0.543603
R534 source.n287 source.n255 0.543603
R535 source.n103 source.n71 0.470328
R536 source.n247 source.n215 0.470328
R537 source.n268 source.n267 0.388379
R538 source.n228 source.n227 0.388379
R539 source.n196 source.n195 0.388379
R540 source.n156 source.n155 0.388379
R541 source.n12 source.n11 0.388379
R542 source.n52 source.n51 0.388379
R543 source.n84 source.n83 0.388379
R544 source.n124 source.n123 0.388379
R545 source source.n288 0.188
R546 source.n270 source.n269 0.155672
R547 source.n270 source.n261 0.155672
R548 source.n277 source.n261 0.155672
R549 source.n278 source.n277 0.155672
R550 source.n278 source.n257 0.155672
R551 source.n285 source.n257 0.155672
R552 source.n230 source.n229 0.155672
R553 source.n230 source.n221 0.155672
R554 source.n237 source.n221 0.155672
R555 source.n238 source.n237 0.155672
R556 source.n238 source.n217 0.155672
R557 source.n245 source.n217 0.155672
R558 source.n198 source.n197 0.155672
R559 source.n198 source.n189 0.155672
R560 source.n205 source.n189 0.155672
R561 source.n206 source.n205 0.155672
R562 source.n206 source.n185 0.155672
R563 source.n213 source.n185 0.155672
R564 source.n158 source.n157 0.155672
R565 source.n158 source.n149 0.155672
R566 source.n165 source.n149 0.155672
R567 source.n166 source.n165 0.155672
R568 source.n166 source.n145 0.155672
R569 source.n173 source.n145 0.155672
R570 source.n29 source.n1 0.155672
R571 source.n22 source.n1 0.155672
R572 source.n22 source.n21 0.155672
R573 source.n21 source.n5 0.155672
R574 source.n14 source.n5 0.155672
R575 source.n14 source.n13 0.155672
R576 source.n69 source.n41 0.155672
R577 source.n62 source.n41 0.155672
R578 source.n62 source.n61 0.155672
R579 source.n61 source.n45 0.155672
R580 source.n54 source.n45 0.155672
R581 source.n54 source.n53 0.155672
R582 source.n101 source.n73 0.155672
R583 source.n94 source.n73 0.155672
R584 source.n94 source.n93 0.155672
R585 source.n93 source.n77 0.155672
R586 source.n86 source.n77 0.155672
R587 source.n86 source.n85 0.155672
R588 source.n141 source.n113 0.155672
R589 source.n134 source.n113 0.155672
R590 source.n134 source.n133 0.155672
R591 source.n133 source.n117 0.155672
R592 source.n126 source.n117 0.155672
R593 source.n126 source.n125 0.155672
R594 plus.n6 plus.t2 635.365
R595 plus.n27 plus.t15 635.365
R596 plus.n36 plus.t9 635.365
R597 plus.n56 plus.t6 635.365
R598 plus.n5 plus.t8 586.433
R599 plus.n9 plus.t13 586.433
R600 plus.n3 plus.t19 586.433
R601 plus.n15 plus.t7 586.433
R602 plus.n17 plus.t12 586.433
R603 plus.n18 plus.t18 586.433
R604 plus.n24 plus.t0 586.433
R605 plus.n26 plus.t11 586.433
R606 plus.n35 plus.t1 586.433
R607 plus.n39 plus.t10 586.433
R608 plus.n33 plus.t3 586.433
R609 plus.n45 plus.t16 586.433
R610 plus.n47 plus.t4 586.433
R611 plus.n32 plus.t17 586.433
R612 plus.n53 plus.t5 586.433
R613 plus.n55 plus.t14 586.433
R614 plus.n7 plus.n6 161.489
R615 plus.n37 plus.n36 161.489
R616 plus.n8 plus.n7 161.3
R617 plus.n10 plus.n4 161.3
R618 plus.n12 plus.n11 161.3
R619 plus.n14 plus.n13 161.3
R620 plus.n16 plus.n2 161.3
R621 plus.n20 plus.n19 161.3
R622 plus.n21 plus.n1 161.3
R623 plus.n23 plus.n22 161.3
R624 plus.n25 plus.n0 161.3
R625 plus.n28 plus.n27 161.3
R626 plus.n38 plus.n37 161.3
R627 plus.n40 plus.n34 161.3
R628 plus.n42 plus.n41 161.3
R629 plus.n44 plus.n43 161.3
R630 plus.n46 plus.n31 161.3
R631 plus.n49 plus.n48 161.3
R632 plus.n50 plus.n30 161.3
R633 plus.n52 plus.n51 161.3
R634 plus.n54 plus.n29 161.3
R635 plus.n57 plus.n56 161.3
R636 plus.n11 plus.n10 73.0308
R637 plus.n23 plus.n1 73.0308
R638 plus.n52 plus.n30 73.0308
R639 plus.n41 plus.n40 73.0308
R640 plus.n14 plus.n3 64.9975
R641 plus.n19 plus.n18 64.9975
R642 plus.n48 plus.n32 64.9975
R643 plus.n44 plus.n33 64.9975
R644 plus.n9 plus.n8 62.0763
R645 plus.n25 plus.n24 62.0763
R646 plus.n54 plus.n53 62.0763
R647 plus.n39 plus.n38 62.0763
R648 plus.n16 plus.n15 46.0096
R649 plus.n17 plus.n16 46.0096
R650 plus.n47 plus.n46 46.0096
R651 plus.n46 plus.n45 46.0096
R652 plus.n6 plus.n5 43.0884
R653 plus.n27 plus.n26 43.0884
R654 plus.n56 plus.n55 43.0884
R655 plus.n36 plus.n35 43.0884
R656 plus.n8 plus.n5 29.9429
R657 plus.n26 plus.n25 29.9429
R658 plus.n55 plus.n54 29.9429
R659 plus.n38 plus.n35 29.9429
R660 plus plus.n57 28.7074
R661 plus.n15 plus.n14 27.0217
R662 plus.n19 plus.n17 27.0217
R663 plus.n48 plus.n47 27.0217
R664 plus.n45 plus.n44 27.0217
R665 plus.n10 plus.n9 10.955
R666 plus.n24 plus.n23 10.955
R667 plus.n53 plus.n52 10.955
R668 plus.n40 plus.n39 10.955
R669 plus plus.n28 9.88686
R670 plus.n11 plus.n3 8.03383
R671 plus.n18 plus.n1 8.03383
R672 plus.n32 plus.n30 8.03383
R673 plus.n41 plus.n33 8.03383
R674 plus.n7 plus.n4 0.189894
R675 plus.n12 plus.n4 0.189894
R676 plus.n13 plus.n12 0.189894
R677 plus.n13 plus.n2 0.189894
R678 plus.n20 plus.n2 0.189894
R679 plus.n21 plus.n20 0.189894
R680 plus.n22 plus.n21 0.189894
R681 plus.n22 plus.n0 0.189894
R682 plus.n28 plus.n0 0.189894
R683 plus.n57 plus.n29 0.189894
R684 plus.n51 plus.n29 0.189894
R685 plus.n51 plus.n50 0.189894
R686 plus.n50 plus.n49 0.189894
R687 plus.n49 plus.n31 0.189894
R688 plus.n43 plus.n31 0.189894
R689 plus.n43 plus.n42 0.189894
R690 plus.n42 plus.n34 0.189894
R691 plus.n37 plus.n34 0.189894
R692 drain_left.n10 drain_left.n8 67.7339
R693 drain_left.n6 drain_left.n4 67.7338
R694 drain_left.n2 drain_left.n0 67.7338
R695 drain_left.n14 drain_left.n13 67.1908
R696 drain_left.n12 drain_left.n11 67.1908
R697 drain_left.n10 drain_left.n9 67.1908
R698 drain_left.n16 drain_left.n15 67.1907
R699 drain_left.n7 drain_left.n3 67.1907
R700 drain_left.n6 drain_left.n5 67.1907
R701 drain_left.n2 drain_left.n1 67.1907
R702 drain_left drain_left.n7 27.1664
R703 drain_left drain_left.n16 6.19632
R704 drain_left.n3 drain_left.t15 3.3005
R705 drain_left.n3 drain_left.t3 3.3005
R706 drain_left.n4 drain_left.t18 3.3005
R707 drain_left.n4 drain_left.t10 3.3005
R708 drain_left.n5 drain_left.t16 3.3005
R709 drain_left.n5 drain_left.t9 3.3005
R710 drain_left.n1 drain_left.t14 3.3005
R711 drain_left.n1 drain_left.t2 3.3005
R712 drain_left.n0 drain_left.t13 3.3005
R713 drain_left.n0 drain_left.t5 3.3005
R714 drain_left.n15 drain_left.t8 3.3005
R715 drain_left.n15 drain_left.t4 3.3005
R716 drain_left.n13 drain_left.t1 3.3005
R717 drain_left.n13 drain_left.t19 3.3005
R718 drain_left.n11 drain_left.t12 3.3005
R719 drain_left.n11 drain_left.t7 3.3005
R720 drain_left.n9 drain_left.t6 3.3005
R721 drain_left.n9 drain_left.t0 3.3005
R722 drain_left.n8 drain_left.t17 3.3005
R723 drain_left.n8 drain_left.t11 3.3005
R724 drain_left.n12 drain_left.n10 0.543603
R725 drain_left.n14 drain_left.n12 0.543603
R726 drain_left.n16 drain_left.n14 0.543603
R727 drain_left.n7 drain_left.n6 0.488257
R728 drain_left.n7 drain_left.n2 0.488257
C0 drain_left minus 0.171748f
C1 plus drain_right 0.36079f
C2 plus source 3.96573f
C3 drain_right source 20.3851f
C4 drain_left plus 4.09834f
C5 drain_left drain_right 1.10832f
C6 minus plus 4.66333f
C7 drain_left source 20.3846f
C8 minus drain_right 3.89238f
C9 minus source 3.95171f
C10 drain_right a_n2102_n2088# 5.59581f
C11 drain_left a_n2102_n2088# 5.91761f
C12 source a_n2102_n2088# 5.43897f
C13 minus a_n2102_n2088# 7.761909f
C14 plus a_n2102_n2088# 9.4104f
C15 drain_left.t13 a_n2102_n2088# 0.159342f
C16 drain_left.t5 a_n2102_n2088# 0.159342f
C17 drain_left.n0 a_n2102_n2088# 1.33215f
C18 drain_left.t14 a_n2102_n2088# 0.159342f
C19 drain_left.t2 a_n2102_n2088# 0.159342f
C20 drain_left.n1 a_n2102_n2088# 1.32891f
C21 drain_left.n2 a_n2102_n2088# 0.786676f
C22 drain_left.t15 a_n2102_n2088# 0.159342f
C23 drain_left.t3 a_n2102_n2088# 0.159342f
C24 drain_left.n3 a_n2102_n2088# 1.32891f
C25 drain_left.t18 a_n2102_n2088# 0.159342f
C26 drain_left.t10 a_n2102_n2088# 0.159342f
C27 drain_left.n4 a_n2102_n2088# 1.33215f
C28 drain_left.t16 a_n2102_n2088# 0.159342f
C29 drain_left.t9 a_n2102_n2088# 0.159342f
C30 drain_left.n5 a_n2102_n2088# 1.32891f
C31 drain_left.n6 a_n2102_n2088# 0.786676f
C32 drain_left.n7 a_n2102_n2088# 1.63104f
C33 drain_left.t17 a_n2102_n2088# 0.159342f
C34 drain_left.t11 a_n2102_n2088# 0.159342f
C35 drain_left.n8 a_n2102_n2088# 1.33216f
C36 drain_left.t6 a_n2102_n2088# 0.159342f
C37 drain_left.t0 a_n2102_n2088# 0.159342f
C38 drain_left.n9 a_n2102_n2088# 1.32892f
C39 drain_left.n10 a_n2102_n2088# 0.791059f
C40 drain_left.t12 a_n2102_n2088# 0.159342f
C41 drain_left.t7 a_n2102_n2088# 0.159342f
C42 drain_left.n11 a_n2102_n2088# 1.32892f
C43 drain_left.n12 a_n2102_n2088# 0.390381f
C44 drain_left.t1 a_n2102_n2088# 0.159342f
C45 drain_left.t19 a_n2102_n2088# 0.159342f
C46 drain_left.n13 a_n2102_n2088# 1.32892f
C47 drain_left.n14 a_n2102_n2088# 0.390381f
C48 drain_left.t8 a_n2102_n2088# 0.159342f
C49 drain_left.t4 a_n2102_n2088# 0.159342f
C50 drain_left.n15 a_n2102_n2088# 1.32891f
C51 drain_left.n16 a_n2102_n2088# 0.670116f
C52 plus.n0 a_n2102_n2088# 0.051006f
C53 plus.t11 a_n2102_n2088# 0.261588f
C54 plus.t0 a_n2102_n2088# 0.261588f
C55 plus.n1 a_n2102_n2088# 0.01865f
C56 plus.n2 a_n2102_n2088# 0.051006f
C57 plus.t12 a_n2102_n2088# 0.261588f
C58 plus.t7 a_n2102_n2088# 0.261588f
C59 plus.t19 a_n2102_n2088# 0.261588f
C60 plus.n3 a_n2102_n2088# 0.120073f
C61 plus.n4 a_n2102_n2088# 0.051006f
C62 plus.t13 a_n2102_n2088# 0.261588f
C63 plus.t8 a_n2102_n2088# 0.261588f
C64 plus.n5 a_n2102_n2088# 0.120073f
C65 plus.t2 a_n2102_n2088# 0.271162f
C66 plus.n6 a_n2102_n2088# 0.13583f
C67 plus.n7 a_n2102_n2088# 0.116716f
C68 plus.n8 a_n2102_n2088# 0.021009f
C69 plus.n9 a_n2102_n2088# 0.120073f
C70 plus.n10 a_n2102_n2088# 0.019279f
C71 plus.n11 a_n2102_n2088# 0.01865f
C72 plus.n12 a_n2102_n2088# 0.051006f
C73 plus.n13 a_n2102_n2088# 0.051006f
C74 plus.n14 a_n2102_n2088# 0.021009f
C75 plus.n15 a_n2102_n2088# 0.120073f
C76 plus.n16 a_n2102_n2088# 0.021009f
C77 plus.n17 a_n2102_n2088# 0.120073f
C78 plus.t18 a_n2102_n2088# 0.261588f
C79 plus.n18 a_n2102_n2088# 0.120073f
C80 plus.n19 a_n2102_n2088# 0.021009f
C81 plus.n20 a_n2102_n2088# 0.051006f
C82 plus.n21 a_n2102_n2088# 0.051006f
C83 plus.n22 a_n2102_n2088# 0.051006f
C84 plus.n23 a_n2102_n2088# 0.019279f
C85 plus.n24 a_n2102_n2088# 0.120073f
C86 plus.n25 a_n2102_n2088# 0.021009f
C87 plus.n26 a_n2102_n2088# 0.120073f
C88 plus.t15 a_n2102_n2088# 0.271162f
C89 plus.n27 a_n2102_n2088# 0.135753f
C90 plus.n28 a_n2102_n2088# 0.439033f
C91 plus.n29 a_n2102_n2088# 0.051006f
C92 plus.t6 a_n2102_n2088# 0.271162f
C93 plus.t14 a_n2102_n2088# 0.261588f
C94 plus.t5 a_n2102_n2088# 0.261588f
C95 plus.n30 a_n2102_n2088# 0.01865f
C96 plus.n31 a_n2102_n2088# 0.051006f
C97 plus.t17 a_n2102_n2088# 0.261588f
C98 plus.n32 a_n2102_n2088# 0.120073f
C99 plus.t4 a_n2102_n2088# 0.261588f
C100 plus.t16 a_n2102_n2088# 0.261588f
C101 plus.t3 a_n2102_n2088# 0.261588f
C102 plus.n33 a_n2102_n2088# 0.120073f
C103 plus.n34 a_n2102_n2088# 0.051006f
C104 plus.t10 a_n2102_n2088# 0.261588f
C105 plus.t1 a_n2102_n2088# 0.261588f
C106 plus.n35 a_n2102_n2088# 0.120073f
C107 plus.t9 a_n2102_n2088# 0.271162f
C108 plus.n36 a_n2102_n2088# 0.13583f
C109 plus.n37 a_n2102_n2088# 0.116716f
C110 plus.n38 a_n2102_n2088# 0.021009f
C111 plus.n39 a_n2102_n2088# 0.120073f
C112 plus.n40 a_n2102_n2088# 0.019279f
C113 plus.n41 a_n2102_n2088# 0.01865f
C114 plus.n42 a_n2102_n2088# 0.051006f
C115 plus.n43 a_n2102_n2088# 0.051006f
C116 plus.n44 a_n2102_n2088# 0.021009f
C117 plus.n45 a_n2102_n2088# 0.120073f
C118 plus.n46 a_n2102_n2088# 0.021009f
C119 plus.n47 a_n2102_n2088# 0.120073f
C120 plus.n48 a_n2102_n2088# 0.021009f
C121 plus.n49 a_n2102_n2088# 0.051006f
C122 plus.n50 a_n2102_n2088# 0.051006f
C123 plus.n51 a_n2102_n2088# 0.051006f
C124 plus.n52 a_n2102_n2088# 0.019279f
C125 plus.n53 a_n2102_n2088# 0.120073f
C126 plus.n54 a_n2102_n2088# 0.021009f
C127 plus.n55 a_n2102_n2088# 0.120073f
C128 plus.n56 a_n2102_n2088# 0.135753f
C129 plus.n57 a_n2102_n2088# 1.37523f
C130 source.n0 a_n2102_n2088# 0.043336f
C131 source.n1 a_n2102_n2088# 0.030831f
C132 source.n2 a_n2102_n2088# 0.016568f
C133 source.n3 a_n2102_n2088# 0.03916f
C134 source.n4 a_n2102_n2088# 0.017542f
C135 source.n5 a_n2102_n2088# 0.030831f
C136 source.n6 a_n2102_n2088# 0.016568f
C137 source.n7 a_n2102_n2088# 0.03916f
C138 source.n8 a_n2102_n2088# 0.017542f
C139 source.n9 a_n2102_n2088# 0.131937f
C140 source.t14 a_n2102_n2088# 0.063825f
C141 source.n10 a_n2102_n2088# 0.02937f
C142 source.n11 a_n2102_n2088# 0.023131f
C143 source.n12 a_n2102_n2088# 0.016568f
C144 source.n13 a_n2102_n2088# 0.733605f
C145 source.n14 a_n2102_n2088# 0.030831f
C146 source.n15 a_n2102_n2088# 0.016568f
C147 source.n16 a_n2102_n2088# 0.017542f
C148 source.n17 a_n2102_n2088# 0.03916f
C149 source.n18 a_n2102_n2088# 0.03916f
C150 source.n19 a_n2102_n2088# 0.017542f
C151 source.n20 a_n2102_n2088# 0.016568f
C152 source.n21 a_n2102_n2088# 0.030831f
C153 source.n22 a_n2102_n2088# 0.030831f
C154 source.n23 a_n2102_n2088# 0.016568f
C155 source.n24 a_n2102_n2088# 0.017542f
C156 source.n25 a_n2102_n2088# 0.03916f
C157 source.n26 a_n2102_n2088# 0.084774f
C158 source.n27 a_n2102_n2088# 0.017542f
C159 source.n28 a_n2102_n2088# 0.016568f
C160 source.n29 a_n2102_n2088# 0.071266f
C161 source.n30 a_n2102_n2088# 0.047434f
C162 source.n31 a_n2102_n2088# 0.7468f
C163 source.t15 a_n2102_n2088# 0.146184f
C164 source.t4 a_n2102_n2088# 0.146184f
C165 source.n32 a_n2102_n2088# 1.13849f
C166 source.n33 a_n2102_n2088# 0.396926f
C167 source.t0 a_n2102_n2088# 0.146184f
C168 source.t13 a_n2102_n2088# 0.146184f
C169 source.n34 a_n2102_n2088# 1.13849f
C170 source.n35 a_n2102_n2088# 0.396926f
C171 source.t6 a_n2102_n2088# 0.146184f
C172 source.t10 a_n2102_n2088# 0.146184f
C173 source.n36 a_n2102_n2088# 1.13849f
C174 source.n37 a_n2102_n2088# 0.396926f
C175 source.t9 a_n2102_n2088# 0.146184f
C176 source.t17 a_n2102_n2088# 0.146184f
C177 source.n38 a_n2102_n2088# 1.13849f
C178 source.n39 a_n2102_n2088# 0.396926f
C179 source.n40 a_n2102_n2088# 0.043336f
C180 source.n41 a_n2102_n2088# 0.030831f
C181 source.n42 a_n2102_n2088# 0.016568f
C182 source.n43 a_n2102_n2088# 0.03916f
C183 source.n44 a_n2102_n2088# 0.017542f
C184 source.n45 a_n2102_n2088# 0.030831f
C185 source.n46 a_n2102_n2088# 0.016568f
C186 source.n47 a_n2102_n2088# 0.03916f
C187 source.n48 a_n2102_n2088# 0.017542f
C188 source.n49 a_n2102_n2088# 0.131937f
C189 source.t8 a_n2102_n2088# 0.063825f
C190 source.n50 a_n2102_n2088# 0.02937f
C191 source.n51 a_n2102_n2088# 0.023131f
C192 source.n52 a_n2102_n2088# 0.016568f
C193 source.n53 a_n2102_n2088# 0.733605f
C194 source.n54 a_n2102_n2088# 0.030831f
C195 source.n55 a_n2102_n2088# 0.016568f
C196 source.n56 a_n2102_n2088# 0.017542f
C197 source.n57 a_n2102_n2088# 0.03916f
C198 source.n58 a_n2102_n2088# 0.03916f
C199 source.n59 a_n2102_n2088# 0.017542f
C200 source.n60 a_n2102_n2088# 0.016568f
C201 source.n61 a_n2102_n2088# 0.030831f
C202 source.n62 a_n2102_n2088# 0.030831f
C203 source.n63 a_n2102_n2088# 0.016568f
C204 source.n64 a_n2102_n2088# 0.017542f
C205 source.n65 a_n2102_n2088# 0.03916f
C206 source.n66 a_n2102_n2088# 0.084774f
C207 source.n67 a_n2102_n2088# 0.017542f
C208 source.n68 a_n2102_n2088# 0.016568f
C209 source.n69 a_n2102_n2088# 0.071266f
C210 source.n70 a_n2102_n2088# 0.047434f
C211 source.n71 a_n2102_n2088# 0.126963f
C212 source.n72 a_n2102_n2088# 0.043336f
C213 source.n73 a_n2102_n2088# 0.030831f
C214 source.n74 a_n2102_n2088# 0.016568f
C215 source.n75 a_n2102_n2088# 0.03916f
C216 source.n76 a_n2102_n2088# 0.017542f
C217 source.n77 a_n2102_n2088# 0.030831f
C218 source.n78 a_n2102_n2088# 0.016568f
C219 source.n79 a_n2102_n2088# 0.03916f
C220 source.n80 a_n2102_n2088# 0.017542f
C221 source.n81 a_n2102_n2088# 0.131937f
C222 source.t26 a_n2102_n2088# 0.063825f
C223 source.n82 a_n2102_n2088# 0.02937f
C224 source.n83 a_n2102_n2088# 0.023131f
C225 source.n84 a_n2102_n2088# 0.016568f
C226 source.n85 a_n2102_n2088# 0.733605f
C227 source.n86 a_n2102_n2088# 0.030831f
C228 source.n87 a_n2102_n2088# 0.016568f
C229 source.n88 a_n2102_n2088# 0.017542f
C230 source.n89 a_n2102_n2088# 0.03916f
C231 source.n90 a_n2102_n2088# 0.03916f
C232 source.n91 a_n2102_n2088# 0.017542f
C233 source.n92 a_n2102_n2088# 0.016568f
C234 source.n93 a_n2102_n2088# 0.030831f
C235 source.n94 a_n2102_n2088# 0.030831f
C236 source.n95 a_n2102_n2088# 0.016568f
C237 source.n96 a_n2102_n2088# 0.017542f
C238 source.n97 a_n2102_n2088# 0.03916f
C239 source.n98 a_n2102_n2088# 0.084774f
C240 source.n99 a_n2102_n2088# 0.017542f
C241 source.n100 a_n2102_n2088# 0.016568f
C242 source.n101 a_n2102_n2088# 0.071266f
C243 source.n102 a_n2102_n2088# 0.047434f
C244 source.n103 a_n2102_n2088# 0.126963f
C245 source.t36 a_n2102_n2088# 0.146184f
C246 source.t21 a_n2102_n2088# 0.146184f
C247 source.n104 a_n2102_n2088# 1.13849f
C248 source.n105 a_n2102_n2088# 0.396926f
C249 source.t22 a_n2102_n2088# 0.146184f
C250 source.t27 a_n2102_n2088# 0.146184f
C251 source.n106 a_n2102_n2088# 1.13849f
C252 source.n107 a_n2102_n2088# 0.396926f
C253 source.t34 a_n2102_n2088# 0.146184f
C254 source.t37 a_n2102_n2088# 0.146184f
C255 source.n108 a_n2102_n2088# 1.13849f
C256 source.n109 a_n2102_n2088# 0.396926f
C257 source.t35 a_n2102_n2088# 0.146184f
C258 source.t20 a_n2102_n2088# 0.146184f
C259 source.n110 a_n2102_n2088# 1.13849f
C260 source.n111 a_n2102_n2088# 0.396926f
C261 source.n112 a_n2102_n2088# 0.043336f
C262 source.n113 a_n2102_n2088# 0.030831f
C263 source.n114 a_n2102_n2088# 0.016568f
C264 source.n115 a_n2102_n2088# 0.03916f
C265 source.n116 a_n2102_n2088# 0.017542f
C266 source.n117 a_n2102_n2088# 0.030831f
C267 source.n118 a_n2102_n2088# 0.016568f
C268 source.n119 a_n2102_n2088# 0.03916f
C269 source.n120 a_n2102_n2088# 0.017542f
C270 source.n121 a_n2102_n2088# 0.131937f
C271 source.t31 a_n2102_n2088# 0.063825f
C272 source.n122 a_n2102_n2088# 0.02937f
C273 source.n123 a_n2102_n2088# 0.023131f
C274 source.n124 a_n2102_n2088# 0.016568f
C275 source.n125 a_n2102_n2088# 0.733605f
C276 source.n126 a_n2102_n2088# 0.030831f
C277 source.n127 a_n2102_n2088# 0.016568f
C278 source.n128 a_n2102_n2088# 0.017542f
C279 source.n129 a_n2102_n2088# 0.03916f
C280 source.n130 a_n2102_n2088# 0.03916f
C281 source.n131 a_n2102_n2088# 0.017542f
C282 source.n132 a_n2102_n2088# 0.016568f
C283 source.n133 a_n2102_n2088# 0.030831f
C284 source.n134 a_n2102_n2088# 0.030831f
C285 source.n135 a_n2102_n2088# 0.016568f
C286 source.n136 a_n2102_n2088# 0.017542f
C287 source.n137 a_n2102_n2088# 0.03916f
C288 source.n138 a_n2102_n2088# 0.084774f
C289 source.n139 a_n2102_n2088# 0.017542f
C290 source.n140 a_n2102_n2088# 0.016568f
C291 source.n141 a_n2102_n2088# 0.071266f
C292 source.n142 a_n2102_n2088# 0.047434f
C293 source.n143 a_n2102_n2088# 1.14372f
C294 source.n144 a_n2102_n2088# 0.043336f
C295 source.n145 a_n2102_n2088# 0.030831f
C296 source.n146 a_n2102_n2088# 0.016568f
C297 source.n147 a_n2102_n2088# 0.03916f
C298 source.n148 a_n2102_n2088# 0.017542f
C299 source.n149 a_n2102_n2088# 0.030831f
C300 source.n150 a_n2102_n2088# 0.016568f
C301 source.n151 a_n2102_n2088# 0.03916f
C302 source.n152 a_n2102_n2088# 0.017542f
C303 source.n153 a_n2102_n2088# 0.131937f
C304 source.t16 a_n2102_n2088# 0.063825f
C305 source.n154 a_n2102_n2088# 0.02937f
C306 source.n155 a_n2102_n2088# 0.023131f
C307 source.n156 a_n2102_n2088# 0.016568f
C308 source.n157 a_n2102_n2088# 0.733605f
C309 source.n158 a_n2102_n2088# 0.030831f
C310 source.n159 a_n2102_n2088# 0.016568f
C311 source.n160 a_n2102_n2088# 0.017542f
C312 source.n161 a_n2102_n2088# 0.03916f
C313 source.n162 a_n2102_n2088# 0.03916f
C314 source.n163 a_n2102_n2088# 0.017542f
C315 source.n164 a_n2102_n2088# 0.016568f
C316 source.n165 a_n2102_n2088# 0.030831f
C317 source.n166 a_n2102_n2088# 0.030831f
C318 source.n167 a_n2102_n2088# 0.016568f
C319 source.n168 a_n2102_n2088# 0.017542f
C320 source.n169 a_n2102_n2088# 0.03916f
C321 source.n170 a_n2102_n2088# 0.084774f
C322 source.n171 a_n2102_n2088# 0.017542f
C323 source.n172 a_n2102_n2088# 0.016568f
C324 source.n173 a_n2102_n2088# 0.071266f
C325 source.n174 a_n2102_n2088# 0.047434f
C326 source.n175 a_n2102_n2088# 1.14372f
C327 source.t12 a_n2102_n2088# 0.146184f
C328 source.t3 a_n2102_n2088# 0.146184f
C329 source.n176 a_n2102_n2088# 1.13848f
C330 source.n177 a_n2102_n2088# 0.396934f
C331 source.t11 a_n2102_n2088# 0.146184f
C332 source.t5 a_n2102_n2088# 0.146184f
C333 source.n178 a_n2102_n2088# 1.13848f
C334 source.n179 a_n2102_n2088# 0.396934f
C335 source.t7 a_n2102_n2088# 0.146184f
C336 source.t1 a_n2102_n2088# 0.146184f
C337 source.n180 a_n2102_n2088# 1.13848f
C338 source.n181 a_n2102_n2088# 0.396934f
C339 source.t19 a_n2102_n2088# 0.146184f
C340 source.t2 a_n2102_n2088# 0.146184f
C341 source.n182 a_n2102_n2088# 1.13848f
C342 source.n183 a_n2102_n2088# 0.396934f
C343 source.n184 a_n2102_n2088# 0.043336f
C344 source.n185 a_n2102_n2088# 0.030831f
C345 source.n186 a_n2102_n2088# 0.016568f
C346 source.n187 a_n2102_n2088# 0.03916f
C347 source.n188 a_n2102_n2088# 0.017542f
C348 source.n189 a_n2102_n2088# 0.030831f
C349 source.n190 a_n2102_n2088# 0.016568f
C350 source.n191 a_n2102_n2088# 0.03916f
C351 source.n192 a_n2102_n2088# 0.017542f
C352 source.n193 a_n2102_n2088# 0.131937f
C353 source.t18 a_n2102_n2088# 0.063825f
C354 source.n194 a_n2102_n2088# 0.02937f
C355 source.n195 a_n2102_n2088# 0.023131f
C356 source.n196 a_n2102_n2088# 0.016568f
C357 source.n197 a_n2102_n2088# 0.733605f
C358 source.n198 a_n2102_n2088# 0.030831f
C359 source.n199 a_n2102_n2088# 0.016568f
C360 source.n200 a_n2102_n2088# 0.017542f
C361 source.n201 a_n2102_n2088# 0.03916f
C362 source.n202 a_n2102_n2088# 0.03916f
C363 source.n203 a_n2102_n2088# 0.017542f
C364 source.n204 a_n2102_n2088# 0.016568f
C365 source.n205 a_n2102_n2088# 0.030831f
C366 source.n206 a_n2102_n2088# 0.030831f
C367 source.n207 a_n2102_n2088# 0.016568f
C368 source.n208 a_n2102_n2088# 0.017542f
C369 source.n209 a_n2102_n2088# 0.03916f
C370 source.n210 a_n2102_n2088# 0.084774f
C371 source.n211 a_n2102_n2088# 0.017542f
C372 source.n212 a_n2102_n2088# 0.016568f
C373 source.n213 a_n2102_n2088# 0.071266f
C374 source.n214 a_n2102_n2088# 0.047434f
C375 source.n215 a_n2102_n2088# 0.126963f
C376 source.n216 a_n2102_n2088# 0.043336f
C377 source.n217 a_n2102_n2088# 0.030831f
C378 source.n218 a_n2102_n2088# 0.016568f
C379 source.n219 a_n2102_n2088# 0.03916f
C380 source.n220 a_n2102_n2088# 0.017542f
C381 source.n221 a_n2102_n2088# 0.030831f
C382 source.n222 a_n2102_n2088# 0.016568f
C383 source.n223 a_n2102_n2088# 0.03916f
C384 source.n224 a_n2102_n2088# 0.017542f
C385 source.n225 a_n2102_n2088# 0.131937f
C386 source.t24 a_n2102_n2088# 0.063825f
C387 source.n226 a_n2102_n2088# 0.02937f
C388 source.n227 a_n2102_n2088# 0.023131f
C389 source.n228 a_n2102_n2088# 0.016568f
C390 source.n229 a_n2102_n2088# 0.733605f
C391 source.n230 a_n2102_n2088# 0.030831f
C392 source.n231 a_n2102_n2088# 0.016568f
C393 source.n232 a_n2102_n2088# 0.017542f
C394 source.n233 a_n2102_n2088# 0.03916f
C395 source.n234 a_n2102_n2088# 0.03916f
C396 source.n235 a_n2102_n2088# 0.017542f
C397 source.n236 a_n2102_n2088# 0.016568f
C398 source.n237 a_n2102_n2088# 0.030831f
C399 source.n238 a_n2102_n2088# 0.030831f
C400 source.n239 a_n2102_n2088# 0.016568f
C401 source.n240 a_n2102_n2088# 0.017542f
C402 source.n241 a_n2102_n2088# 0.03916f
C403 source.n242 a_n2102_n2088# 0.084774f
C404 source.n243 a_n2102_n2088# 0.017542f
C405 source.n244 a_n2102_n2088# 0.016568f
C406 source.n245 a_n2102_n2088# 0.071266f
C407 source.n246 a_n2102_n2088# 0.047434f
C408 source.n247 a_n2102_n2088# 0.126963f
C409 source.t32 a_n2102_n2088# 0.146184f
C410 source.t25 a_n2102_n2088# 0.146184f
C411 source.n248 a_n2102_n2088# 1.13848f
C412 source.n249 a_n2102_n2088# 0.396934f
C413 source.t33 a_n2102_n2088# 0.146184f
C414 source.t38 a_n2102_n2088# 0.146184f
C415 source.n250 a_n2102_n2088# 1.13848f
C416 source.n251 a_n2102_n2088# 0.396934f
C417 source.t28 a_n2102_n2088# 0.146184f
C418 source.t39 a_n2102_n2088# 0.146184f
C419 source.n252 a_n2102_n2088# 1.13848f
C420 source.n253 a_n2102_n2088# 0.396934f
C421 source.t29 a_n2102_n2088# 0.146184f
C422 source.t30 a_n2102_n2088# 0.146184f
C423 source.n254 a_n2102_n2088# 1.13848f
C424 source.n255 a_n2102_n2088# 0.396934f
C425 source.n256 a_n2102_n2088# 0.043336f
C426 source.n257 a_n2102_n2088# 0.030831f
C427 source.n258 a_n2102_n2088# 0.016568f
C428 source.n259 a_n2102_n2088# 0.03916f
C429 source.n260 a_n2102_n2088# 0.017542f
C430 source.n261 a_n2102_n2088# 0.030831f
C431 source.n262 a_n2102_n2088# 0.016568f
C432 source.n263 a_n2102_n2088# 0.03916f
C433 source.n264 a_n2102_n2088# 0.017542f
C434 source.n265 a_n2102_n2088# 0.131937f
C435 source.t23 a_n2102_n2088# 0.063825f
C436 source.n266 a_n2102_n2088# 0.02937f
C437 source.n267 a_n2102_n2088# 0.023131f
C438 source.n268 a_n2102_n2088# 0.016568f
C439 source.n269 a_n2102_n2088# 0.733605f
C440 source.n270 a_n2102_n2088# 0.030831f
C441 source.n271 a_n2102_n2088# 0.016568f
C442 source.n272 a_n2102_n2088# 0.017542f
C443 source.n273 a_n2102_n2088# 0.03916f
C444 source.n274 a_n2102_n2088# 0.03916f
C445 source.n275 a_n2102_n2088# 0.017542f
C446 source.n276 a_n2102_n2088# 0.016568f
C447 source.n277 a_n2102_n2088# 0.030831f
C448 source.n278 a_n2102_n2088# 0.030831f
C449 source.n279 a_n2102_n2088# 0.016568f
C450 source.n280 a_n2102_n2088# 0.017542f
C451 source.n281 a_n2102_n2088# 0.03916f
C452 source.n282 a_n2102_n2088# 0.084774f
C453 source.n283 a_n2102_n2088# 0.017542f
C454 source.n284 a_n2102_n2088# 0.016568f
C455 source.n285 a_n2102_n2088# 0.071266f
C456 source.n286 a_n2102_n2088# 0.047434f
C457 source.n287 a_n2102_n2088# 0.301006f
C458 source.n288 a_n2102_n2088# 1.26157f
C459 drain_right.t4 a_n2102_n2088# 0.158894f
C460 drain_right.t6 a_n2102_n2088# 0.158894f
C461 drain_right.n0 a_n2102_n2088# 1.32841f
C462 drain_right.t11 a_n2102_n2088# 0.158894f
C463 drain_right.t7 a_n2102_n2088# 0.158894f
C464 drain_right.n1 a_n2102_n2088# 1.32518f
C465 drain_right.n2 a_n2102_n2088# 0.784463f
C466 drain_right.t2 a_n2102_n2088# 0.158894f
C467 drain_right.t8 a_n2102_n2088# 0.158894f
C468 drain_right.n3 a_n2102_n2088# 1.32518f
C469 drain_right.t17 a_n2102_n2088# 0.158894f
C470 drain_right.t5 a_n2102_n2088# 0.158894f
C471 drain_right.n4 a_n2102_n2088# 1.32841f
C472 drain_right.t9 a_n2102_n2088# 0.158894f
C473 drain_right.t16 a_n2102_n2088# 0.158894f
C474 drain_right.n5 a_n2102_n2088# 1.32518f
C475 drain_right.n6 a_n2102_n2088# 0.784463f
C476 drain_right.n7 a_n2102_n2088# 1.55872f
C477 drain_right.t13 a_n2102_n2088# 0.158894f
C478 drain_right.t10 a_n2102_n2088# 0.158894f
C479 drain_right.n8 a_n2102_n2088# 1.32841f
C480 drain_right.t19 a_n2102_n2088# 0.158894f
C481 drain_right.t0 a_n2102_n2088# 0.158894f
C482 drain_right.n9 a_n2102_n2088# 1.32518f
C483 drain_right.n10 a_n2102_n2088# 0.788841f
C484 drain_right.t1 a_n2102_n2088# 0.158894f
C485 drain_right.t3 a_n2102_n2088# 0.158894f
C486 drain_right.n11 a_n2102_n2088# 1.32518f
C487 drain_right.n12 a_n2102_n2088# 0.389283f
C488 drain_right.t15 a_n2102_n2088# 0.158894f
C489 drain_right.t14 a_n2102_n2088# 0.158894f
C490 drain_right.n13 a_n2102_n2088# 1.32518f
C491 drain_right.n14 a_n2102_n2088# 0.389283f
C492 drain_right.t18 a_n2102_n2088# 0.158894f
C493 drain_right.t12 a_n2102_n2088# 0.158894f
C494 drain_right.n15 a_n2102_n2088# 1.32518f
C495 drain_right.n16 a_n2102_n2088# 0.668225f
C496 minus.n0 a_n2102_n2088# 0.049808f
C497 minus.t8 a_n2102_n2088# 0.264791f
C498 minus.t4 a_n2102_n2088# 0.255442f
C499 minus.t19 a_n2102_n2088# 0.255442f
C500 minus.n1 a_n2102_n2088# 0.018212f
C501 minus.n2 a_n2102_n2088# 0.049808f
C502 minus.t5 a_n2102_n2088# 0.255442f
C503 minus.n3 a_n2102_n2088# 0.117252f
C504 minus.t2 a_n2102_n2088# 0.255442f
C505 minus.t17 a_n2102_n2088# 0.255442f
C506 minus.t12 a_n2102_n2088# 0.255442f
C507 minus.n4 a_n2102_n2088# 0.117252f
C508 minus.n5 a_n2102_n2088# 0.049808f
C509 minus.t3 a_n2102_n2088# 0.255442f
C510 minus.t18 a_n2102_n2088# 0.255442f
C511 minus.n6 a_n2102_n2088# 0.117252f
C512 minus.t13 a_n2102_n2088# 0.264791f
C513 minus.n7 a_n2102_n2088# 0.132639f
C514 minus.n8 a_n2102_n2088# 0.113974f
C515 minus.n9 a_n2102_n2088# 0.020515f
C516 minus.n10 a_n2102_n2088# 0.117252f
C517 minus.n11 a_n2102_n2088# 0.018826f
C518 minus.n12 a_n2102_n2088# 0.018212f
C519 minus.n13 a_n2102_n2088# 0.049808f
C520 minus.n14 a_n2102_n2088# 0.049808f
C521 minus.n15 a_n2102_n2088# 0.020515f
C522 minus.n16 a_n2102_n2088# 0.117252f
C523 minus.n17 a_n2102_n2088# 0.020515f
C524 minus.n18 a_n2102_n2088# 0.117252f
C525 minus.n19 a_n2102_n2088# 0.020515f
C526 minus.n20 a_n2102_n2088# 0.049808f
C527 minus.n21 a_n2102_n2088# 0.049808f
C528 minus.n22 a_n2102_n2088# 0.049808f
C529 minus.n23 a_n2102_n2088# 0.018826f
C530 minus.n24 a_n2102_n2088# 0.117252f
C531 minus.n25 a_n2102_n2088# 0.020515f
C532 minus.n26 a_n2102_n2088# 0.117252f
C533 minus.n27 a_n2102_n2088# 0.132564f
C534 minus.n28 a_n2102_n2088# 1.48618f
C535 minus.n29 a_n2102_n2088# 0.049808f
C536 minus.t9 a_n2102_n2088# 0.255442f
C537 minus.t10 a_n2102_n2088# 0.255442f
C538 minus.n30 a_n2102_n2088# 0.018212f
C539 minus.n31 a_n2102_n2088# 0.049808f
C540 minus.t11 a_n2102_n2088# 0.255442f
C541 minus.t1 a_n2102_n2088# 0.255442f
C542 minus.t6 a_n2102_n2088# 0.255442f
C543 minus.n32 a_n2102_n2088# 0.117252f
C544 minus.n33 a_n2102_n2088# 0.049808f
C545 minus.t14 a_n2102_n2088# 0.255442f
C546 minus.t7 a_n2102_n2088# 0.255442f
C547 minus.n34 a_n2102_n2088# 0.117252f
C548 minus.t15 a_n2102_n2088# 0.264791f
C549 minus.n35 a_n2102_n2088# 0.132639f
C550 minus.n36 a_n2102_n2088# 0.113974f
C551 minus.n37 a_n2102_n2088# 0.020515f
C552 minus.n38 a_n2102_n2088# 0.117252f
C553 minus.n39 a_n2102_n2088# 0.018826f
C554 minus.n40 a_n2102_n2088# 0.018212f
C555 minus.n41 a_n2102_n2088# 0.049808f
C556 minus.n42 a_n2102_n2088# 0.049808f
C557 minus.n43 a_n2102_n2088# 0.020515f
C558 minus.n44 a_n2102_n2088# 0.117252f
C559 minus.n45 a_n2102_n2088# 0.020515f
C560 minus.n46 a_n2102_n2088# 0.117252f
C561 minus.t0 a_n2102_n2088# 0.255442f
C562 minus.n47 a_n2102_n2088# 0.117252f
C563 minus.n48 a_n2102_n2088# 0.020515f
C564 minus.n49 a_n2102_n2088# 0.049808f
C565 minus.n50 a_n2102_n2088# 0.049808f
C566 minus.n51 a_n2102_n2088# 0.049808f
C567 minus.n52 a_n2102_n2088# 0.018826f
C568 minus.n53 a_n2102_n2088# 0.117252f
C569 minus.n54 a_n2102_n2088# 0.020515f
C570 minus.n55 a_n2102_n2088# 0.117252f
C571 minus.t16 a_n2102_n2088# 0.264791f
C572 minus.n56 a_n2102_n2088# 0.132564f
C573 minus.n57 a_n2102_n2088# 0.327468f
C574 minus.n58 a_n2102_n2088# 1.82279f
.ends

