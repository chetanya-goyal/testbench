* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t25 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X1 drain_right.t13 minus.t0 source.t12 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 source.t1 minus.t1 drain_right.t12 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_left.t12 plus.t1 source.t19 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X5 drain_right.t11 minus.t2 source.t4 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X6 drain_right.t10 minus.t3 source.t6 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 drain_right.t9 minus.t4 source.t9 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 source.t26 plus.t2 drain_left.t11 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 drain_left.t10 plus.t3 source.t23 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X11 drain_right.t8 minus.t5 source.t11 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X12 drain_left.t9 plus.t4 source.t18 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X13 source.t5 minus.t6 drain_right.t7 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 source.t8 minus.t7 drain_right.t6 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X15 drain_left.t8 plus.t5 source.t24 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X16 drain_right.t5 minus.t8 source.t3 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X17 source.t10 minus.t9 drain_right.t4 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 source.t13 minus.t10 drain_right.t3 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 source.t14 plus.t6 drain_left.t7 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X20 a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X21 source.t22 plus.t7 drain_left.t6 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 source.t21 plus.t8 drain_left.t5 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X24 source.t7 minus.t11 drain_right.t2 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 source.t20 plus.t9 drain_left.t4 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 drain_left.t3 plus.t10 source.t17 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 drain_right.t1 minus.t12 source.t0 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X28 drain_left.t2 plus.t11 source.t15 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X29 drain_left.t1 plus.t12 source.t16 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 drain_right.t0 minus.t13 source.t2 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 source.t27 plus.t13 drain_left.t0 a_n2044_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
R0 plus.n6 plus.n5 161.3
R1 plus.n7 plus.n2 161.3
R2 plus.n10 plus.n1 161.3
R3 plus.n12 plus.n11 161.3
R4 plus.n13 plus.n0 161.3
R5 plus.n15 plus.n14 161.3
R6 plus.n22 plus.n21 161.3
R7 plus.n23 plus.n18 161.3
R8 plus.n26 plus.n17 161.3
R9 plus.n28 plus.n27 161.3
R10 plus.n29 plus.n16 161.3
R11 plus.n31 plus.n30 161.3
R12 plus.n4 plus.t1 147.749
R13 plus.n20 plus.t5 147.749
R14 plus.n14 plus.t4 126.766
R15 plus.n13 plus.t13 126.766
R16 plus.n1 plus.t10 126.766
R17 plus.n8 plus.t2 126.766
R18 plus.n7 plus.t12 126.766
R19 plus.n3 plus.t6 126.766
R20 plus.n30 plus.t11 126.766
R21 plus.n29 plus.t8 126.766
R22 plus.n17 plus.t0 126.766
R23 plus.n24 plus.t9 126.766
R24 plus.n23 plus.t3 126.766
R25 plus.n19 plus.t7 126.766
R26 plus.n9 plus.n8 80.6037
R27 plus.n25 plus.n24 80.6037
R28 plus.n5 plus.n4 70.4033
R29 plus.n21 plus.n20 70.4033
R30 plus.n14 plus.n13 48.2005
R31 plus.n8 plus.n1 48.2005
R32 plus.n8 plus.n7 48.2005
R33 plus.n30 plus.n29 48.2005
R34 plus.n24 plus.n17 48.2005
R35 plus.n24 plus.n23 48.2005
R36 plus plus.n31 26.6714
R37 plus.n12 plus.n1 24.8308
R38 plus.n7 plus.n6 24.8308
R39 plus.n28 plus.n17 24.8308
R40 plus.n23 plus.n22 24.8308
R41 plus.n13 plus.n12 23.3702
R42 plus.n6 plus.n3 23.3702
R43 plus.n29 plus.n28 23.3702
R44 plus.n22 plus.n19 23.3702
R45 plus.n4 plus.n3 20.9576
R46 plus.n20 plus.n19 20.9576
R47 plus plus.n15 8.07058
R48 plus.n9 plus.n2 0.285035
R49 plus.n10 plus.n9 0.285035
R50 plus.n26 plus.n25 0.285035
R51 plus.n25 plus.n18 0.285035
R52 plus.n5 plus.n2 0.189894
R53 plus.n11 plus.n10 0.189894
R54 plus.n11 plus.n0 0.189894
R55 plus.n15 plus.n0 0.189894
R56 plus.n31 plus.n16 0.189894
R57 plus.n27 plus.n16 0.189894
R58 plus.n27 plus.n26 0.189894
R59 plus.n21 plus.n18 0.189894
R60 source.n0 source.t18 243.255
R61 source.n7 source.t3 243.255
R62 source.n27 source.t0 243.254
R63 source.n20 source.t24 243.254
R64 source.n2 source.n1 223.454
R65 source.n4 source.n3 223.454
R66 source.n6 source.n5 223.454
R67 source.n9 source.n8 223.454
R68 source.n11 source.n10 223.454
R69 source.n13 source.n12 223.454
R70 source.n26 source.n25 223.453
R71 source.n24 source.n23 223.453
R72 source.n22 source.n21 223.453
R73 source.n19 source.n18 223.453
R74 source.n17 source.n16 223.453
R75 source.n15 source.n14 223.453
R76 source.n25 source.t2 19.8005
R77 source.n25 source.t13 19.8005
R78 source.n23 source.t9 19.8005
R79 source.n23 source.t8 19.8005
R80 source.n21 source.t11 19.8005
R81 source.n21 source.t10 19.8005
R82 source.n18 source.t23 19.8005
R83 source.n18 source.t22 19.8005
R84 source.n16 source.t25 19.8005
R85 source.n16 source.t20 19.8005
R86 source.n14 source.t15 19.8005
R87 source.n14 source.t21 19.8005
R88 source.n1 source.t17 19.8005
R89 source.n1 source.t27 19.8005
R90 source.n3 source.t16 19.8005
R91 source.n3 source.t26 19.8005
R92 source.n5 source.t19 19.8005
R93 source.n5 source.t14 19.8005
R94 source.n8 source.t6 19.8005
R95 source.n8 source.t1 19.8005
R96 source.n10 source.t4 19.8005
R97 source.n10 source.t7 19.8005
R98 source.n12 source.t12 19.8005
R99 source.n12 source.t5 19.8005
R100 source.n15 source.n13 14.3854
R101 source.n28 source.n0 8.04922
R102 source.n28 source.n27 5.62119
R103 source.n7 source.n6 0.828086
R104 source.n22 source.n20 0.828086
R105 source.n13 source.n11 0.716017
R106 source.n11 source.n9 0.716017
R107 source.n9 source.n7 0.716017
R108 source.n6 source.n4 0.716017
R109 source.n4 source.n2 0.716017
R110 source.n2 source.n0 0.716017
R111 source.n17 source.n15 0.716017
R112 source.n19 source.n17 0.716017
R113 source.n20 source.n19 0.716017
R114 source.n24 source.n22 0.716017
R115 source.n26 source.n24 0.716017
R116 source.n27 source.n26 0.716017
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t12 260.649
R119 drain_left.n1 drain_left.t2 260.647
R120 drain_left.n4 drain_left.n2 240.847
R121 drain_left.n11 drain_left.n10 240.132
R122 drain_left.n9 drain_left.n8 240.132
R123 drain_left.n7 drain_left.n6 240.132
R124 drain_left.n4 drain_left.n3 240.131
R125 drain_left.n1 drain_left.n0 240.131
R126 drain_left drain_left.n5 23.148
R127 drain_left.n2 drain_left.t6 19.8005
R128 drain_left.n2 drain_left.t8 19.8005
R129 drain_left.n3 drain_left.t4 19.8005
R130 drain_left.n3 drain_left.t10 19.8005
R131 drain_left.n0 drain_left.t5 19.8005
R132 drain_left.n0 drain_left.t13 19.8005
R133 drain_left.n10 drain_left.t0 19.8005
R134 drain_left.n10 drain_left.t9 19.8005
R135 drain_left.n8 drain_left.t11 19.8005
R136 drain_left.n8 drain_left.t3 19.8005
R137 drain_left.n6 drain_left.t7 19.8005
R138 drain_left.n6 drain_left.t1 19.8005
R139 drain_left drain_left.n11 6.36873
R140 drain_left.n9 drain_left.n7 0.716017
R141 drain_left.n11 drain_left.n9 0.716017
R142 drain_left.n5 drain_left.n1 0.481792
R143 drain_left.n5 drain_left.n4 0.124033
R144 minus.n15 minus.n14 161.3
R145 minus.n13 minus.n0 161.3
R146 minus.n12 minus.n11 161.3
R147 minus.n10 minus.n1 161.3
R148 minus.n7 minus.n2 161.3
R149 minus.n6 minus.n5 161.3
R150 minus.n31 minus.n30 161.3
R151 minus.n29 minus.n16 161.3
R152 minus.n28 minus.n27 161.3
R153 minus.n26 minus.n17 161.3
R154 minus.n23 minus.n18 161.3
R155 minus.n22 minus.n21 161.3
R156 minus.n4 minus.t8 147.749
R157 minus.n20 minus.t5 147.749
R158 minus.n3 minus.t1 126.766
R159 minus.n7 minus.t3 126.766
R160 minus.n8 minus.t11 126.766
R161 minus.n1 minus.t2 126.766
R162 minus.n13 minus.t6 126.766
R163 minus.n14 minus.t0 126.766
R164 minus.n19 minus.t9 126.766
R165 minus.n23 minus.t4 126.766
R166 minus.n24 minus.t7 126.766
R167 minus.n17 minus.t13 126.766
R168 minus.n29 minus.t10 126.766
R169 minus.n30 minus.t12 126.766
R170 minus.n9 minus.n8 80.6037
R171 minus.n25 minus.n24 80.6037
R172 minus.n5 minus.n4 70.4033
R173 minus.n21 minus.n20 70.4033
R174 minus.n8 minus.n7 48.2005
R175 minus.n8 minus.n1 48.2005
R176 minus.n14 minus.n13 48.2005
R177 minus.n24 minus.n23 48.2005
R178 minus.n24 minus.n17 48.2005
R179 minus.n30 minus.n29 48.2005
R180 minus.n32 minus.n15 28.6236
R181 minus.n7 minus.n6 24.8308
R182 minus.n12 minus.n1 24.8308
R183 minus.n23 minus.n22 24.8308
R184 minus.n28 minus.n17 24.8308
R185 minus.n6 minus.n3 23.3702
R186 minus.n13 minus.n12 23.3702
R187 minus.n22 minus.n19 23.3702
R188 minus.n29 minus.n28 23.3702
R189 minus.n4 minus.n3 20.9576
R190 minus.n20 minus.n19 20.9576
R191 minus.n32 minus.n31 6.5933
R192 minus.n10 minus.n9 0.285035
R193 minus.n9 minus.n2 0.285035
R194 minus.n25 minus.n18 0.285035
R195 minus.n26 minus.n25 0.285035
R196 minus.n15 minus.n0 0.189894
R197 minus.n11 minus.n0 0.189894
R198 minus.n11 minus.n10 0.189894
R199 minus.n5 minus.n2 0.189894
R200 minus.n21 minus.n18 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n16 0.189894
R203 minus.n31 minus.n16 0.189894
R204 minus minus.n32 0.188
R205 drain_right.n1 drain_right.t8 260.647
R206 drain_right.n11 drain_right.t13 259.933
R207 drain_right.n8 drain_right.n6 240.849
R208 drain_right.n4 drain_right.n2 240.847
R209 drain_right.n8 drain_right.n7 240.132
R210 drain_right.n10 drain_right.n9 240.132
R211 drain_right.n4 drain_right.n3 240.131
R212 drain_right.n1 drain_right.n0 240.131
R213 drain_right drain_right.n5 22.5947
R214 drain_right.n2 drain_right.t3 19.8005
R215 drain_right.n2 drain_right.t1 19.8005
R216 drain_right.n3 drain_right.t6 19.8005
R217 drain_right.n3 drain_right.t0 19.8005
R218 drain_right.n0 drain_right.t4 19.8005
R219 drain_right.n0 drain_right.t9 19.8005
R220 drain_right.n6 drain_right.t12 19.8005
R221 drain_right.n6 drain_right.t5 19.8005
R222 drain_right.n7 drain_right.t2 19.8005
R223 drain_right.n7 drain_right.t10 19.8005
R224 drain_right.n9 drain_right.t7 19.8005
R225 drain_right.n9 drain_right.t11 19.8005
R226 drain_right drain_right.n11 6.01097
R227 drain_right.n11 drain_right.n10 0.716017
R228 drain_right.n10 drain_right.n8 0.716017
R229 drain_right.n5 drain_right.n1 0.481792
R230 drain_right.n5 drain_right.n4 0.124033
C0 drain_right drain_left 1.05542f
C1 drain_right minus 1.08565f
C2 drain_left minus 0.180362f
C3 drain_right source 4.49135f
C4 drain_left source 4.49185f
C5 source minus 1.53109f
C6 drain_right plus 0.364786f
C7 drain_left plus 1.28514f
C8 plus minus 3.66829f
C9 plus source 1.54501f
C10 drain_right a_n2044_n1088# 3.82913f
C11 drain_left a_n2044_n1088# 4.10381f
C12 source a_n2044_n1088# 2.248037f
C13 minus a_n2044_n1088# 7.128135f
C14 plus a_n2044_n1088# 7.759729f
C15 drain_right.t8 a_n2044_n1088# 0.103981f
C16 drain_right.t4 a_n2044_n1088# 0.016716f
C17 drain_right.t9 a_n2044_n1088# 0.016716f
C18 drain_right.n0 a_n2044_n1088# 0.064955f
C19 drain_right.n1 a_n2044_n1088# 0.442314f
C20 drain_right.t3 a_n2044_n1088# 0.016716f
C21 drain_right.t1 a_n2044_n1088# 0.016716f
C22 drain_right.n2 a_n2044_n1088# 0.06571f
C23 drain_right.t6 a_n2044_n1088# 0.016716f
C24 drain_right.t0 a_n2044_n1088# 0.016716f
C25 drain_right.n3 a_n2044_n1088# 0.064955f
C26 drain_right.n4 a_n2044_n1088# 0.462332f
C27 drain_right.n5 a_n2044_n1088# 0.577448f
C28 drain_right.t12 a_n2044_n1088# 0.016716f
C29 drain_right.t5 a_n2044_n1088# 0.016716f
C30 drain_right.n6 a_n2044_n1088# 0.06571f
C31 drain_right.t2 a_n2044_n1088# 0.016716f
C32 drain_right.t10 a_n2044_n1088# 0.016716f
C33 drain_right.n7 a_n2044_n1088# 0.064955f
C34 drain_right.n8 a_n2044_n1088# 0.498712f
C35 drain_right.t7 a_n2044_n1088# 0.016716f
C36 drain_right.t11 a_n2044_n1088# 0.016716f
C37 drain_right.n9 a_n2044_n1088# 0.064955f
C38 drain_right.n10 a_n2044_n1088# 0.245473f
C39 drain_right.t13 a_n2044_n1088# 0.103398f
C40 drain_right.n11 a_n2044_n1088# 0.397859f
C41 minus.n0 a_n2044_n1088# 0.028392f
C42 minus.t2 a_n2044_n1088# 0.048138f
C43 minus.n1 a_n2044_n1088# 0.053048f
C44 minus.n2 a_n2044_n1088# 0.037885f
C45 minus.t1 a_n2044_n1088# 0.048138f
C46 minus.n3 a_n2044_n1088# 0.052873f
C47 minus.t8 a_n2044_n1088# 0.055255f
C48 minus.n4 a_n2044_n1088# 0.043173f
C49 minus.n5 a_n2044_n1088# 0.093359f
C50 minus.n6 a_n2044_n1088# 0.006443f
C51 minus.t3 a_n2044_n1088# 0.048138f
C52 minus.n7 a_n2044_n1088# 0.053048f
C53 minus.t11 a_n2044_n1088# 0.048138f
C54 minus.n8 a_n2044_n1088# 0.056515f
C55 minus.n9 a_n2044_n1088# 0.037797f
C56 minus.n10 a_n2044_n1088# 0.037885f
C57 minus.n11 a_n2044_n1088# 0.028392f
C58 minus.n12 a_n2044_n1088# 0.006443f
C59 minus.t6 a_n2044_n1088# 0.048138f
C60 minus.n13 a_n2044_n1088# 0.052873f
C61 minus.t0 a_n2044_n1088# 0.048138f
C62 minus.n14 a_n2044_n1088# 0.050072f
C63 minus.n15 a_n2044_n1088# 0.683586f
C64 minus.n16 a_n2044_n1088# 0.028392f
C65 minus.t13 a_n2044_n1088# 0.048138f
C66 minus.n17 a_n2044_n1088# 0.053048f
C67 minus.n18 a_n2044_n1088# 0.037885f
C68 minus.t9 a_n2044_n1088# 0.048138f
C69 minus.n19 a_n2044_n1088# 0.052873f
C70 minus.t5 a_n2044_n1088# 0.055255f
C71 minus.n20 a_n2044_n1088# 0.043173f
C72 minus.n21 a_n2044_n1088# 0.093359f
C73 minus.n22 a_n2044_n1088# 0.006443f
C74 minus.t4 a_n2044_n1088# 0.048138f
C75 minus.n23 a_n2044_n1088# 0.053048f
C76 minus.t7 a_n2044_n1088# 0.048138f
C77 minus.n24 a_n2044_n1088# 0.056515f
C78 minus.n25 a_n2044_n1088# 0.037797f
C79 minus.n26 a_n2044_n1088# 0.037885f
C80 minus.n27 a_n2044_n1088# 0.028392f
C81 minus.n28 a_n2044_n1088# 0.006443f
C82 minus.t10 a_n2044_n1088# 0.048138f
C83 minus.n29 a_n2044_n1088# 0.052873f
C84 minus.t12 a_n2044_n1088# 0.048138f
C85 minus.n30 a_n2044_n1088# 0.050072f
C86 minus.n31 a_n2044_n1088# 0.191831f
C87 minus.n32 a_n2044_n1088# 0.841383f
C88 drain_left.t2 a_n2044_n1088# 0.102103f
C89 drain_left.t5 a_n2044_n1088# 0.016414f
C90 drain_left.t13 a_n2044_n1088# 0.016414f
C91 drain_left.n0 a_n2044_n1088# 0.063782f
C92 drain_left.n1 a_n2044_n1088# 0.434327f
C93 drain_left.t6 a_n2044_n1088# 0.016414f
C94 drain_left.t8 a_n2044_n1088# 0.016414f
C95 drain_left.n2 a_n2044_n1088# 0.064523f
C96 drain_left.t4 a_n2044_n1088# 0.016414f
C97 drain_left.t10 a_n2044_n1088# 0.016414f
C98 drain_left.n3 a_n2044_n1088# 0.063782f
C99 drain_left.n4 a_n2044_n1088# 0.453983f
C100 drain_left.n5 a_n2044_n1088# 0.607116f
C101 drain_left.t12 a_n2044_n1088# 0.102103f
C102 drain_left.t7 a_n2044_n1088# 0.016414f
C103 drain_left.t1 a_n2044_n1088# 0.016414f
C104 drain_left.n6 a_n2044_n1088# 0.063782f
C105 drain_left.n7 a_n2044_n1088# 0.449003f
C106 drain_left.t11 a_n2044_n1088# 0.016414f
C107 drain_left.t3 a_n2044_n1088# 0.016414f
C108 drain_left.n8 a_n2044_n1088# 0.063782f
C109 drain_left.n9 a_n2044_n1088# 0.241041f
C110 drain_left.t0 a_n2044_n1088# 0.016414f
C111 drain_left.t9 a_n2044_n1088# 0.016414f
C112 drain_left.n10 a_n2044_n1088# 0.063782f
C113 drain_left.n11 a_n2044_n1088# 0.4195f
C114 source.t18 a_n2044_n1088# 0.124938f
C115 source.n0 a_n2044_n1088# 0.564694f
C116 source.t17 a_n2044_n1088# 0.022447f
C117 source.t27 a_n2044_n1088# 0.022447f
C118 source.n1 a_n2044_n1088# 0.0728f
C119 source.n2 a_n2044_n1088# 0.305442f
C120 source.t16 a_n2044_n1088# 0.022447f
C121 source.t26 a_n2044_n1088# 0.022447f
C122 source.n3 a_n2044_n1088# 0.0728f
C123 source.n4 a_n2044_n1088# 0.305442f
C124 source.t19 a_n2044_n1088# 0.022447f
C125 source.t14 a_n2044_n1088# 0.022447f
C126 source.n5 a_n2044_n1088# 0.0728f
C127 source.n6 a_n2044_n1088# 0.3157f
C128 source.t3 a_n2044_n1088# 0.124938f
C129 source.n7 a_n2044_n1088# 0.324782f
C130 source.t6 a_n2044_n1088# 0.022447f
C131 source.t1 a_n2044_n1088# 0.022447f
C132 source.n8 a_n2044_n1088# 0.0728f
C133 source.n9 a_n2044_n1088# 0.305442f
C134 source.t4 a_n2044_n1088# 0.022447f
C135 source.t7 a_n2044_n1088# 0.022447f
C136 source.n10 a_n2044_n1088# 0.0728f
C137 source.n11 a_n2044_n1088# 0.305442f
C138 source.t12 a_n2044_n1088# 0.022447f
C139 source.t5 a_n2044_n1088# 0.022447f
C140 source.n12 a_n2044_n1088# 0.0728f
C141 source.n13 a_n2044_n1088# 0.852053f
C142 source.t15 a_n2044_n1088# 0.022447f
C143 source.t21 a_n2044_n1088# 0.022447f
C144 source.n14 a_n2044_n1088# 0.0728f
C145 source.n15 a_n2044_n1088# 0.852053f
C146 source.t25 a_n2044_n1088# 0.022447f
C147 source.t20 a_n2044_n1088# 0.022447f
C148 source.n16 a_n2044_n1088# 0.0728f
C149 source.n17 a_n2044_n1088# 0.305443f
C150 source.t23 a_n2044_n1088# 0.022447f
C151 source.t22 a_n2044_n1088# 0.022447f
C152 source.n18 a_n2044_n1088# 0.0728f
C153 source.n19 a_n2044_n1088# 0.305443f
C154 source.t24 a_n2044_n1088# 0.124938f
C155 source.n20 a_n2044_n1088# 0.324782f
C156 source.t11 a_n2044_n1088# 0.022447f
C157 source.t10 a_n2044_n1088# 0.022447f
C158 source.n21 a_n2044_n1088# 0.0728f
C159 source.n22 a_n2044_n1088# 0.3157f
C160 source.t9 a_n2044_n1088# 0.022447f
C161 source.t8 a_n2044_n1088# 0.022447f
C162 source.n23 a_n2044_n1088# 0.0728f
C163 source.n24 a_n2044_n1088# 0.305443f
C164 source.t2 a_n2044_n1088# 0.022447f
C165 source.t13 a_n2044_n1088# 0.022447f
C166 source.n25 a_n2044_n1088# 0.0728f
C167 source.n26 a_n2044_n1088# 0.305443f
C168 source.t0 a_n2044_n1088# 0.124938f
C169 source.n27 a_n2044_n1088# 0.464928f
C170 source.n28 a_n2044_n1088# 0.581868f
C171 plus.n0 a_n2044_n1088# 0.028839f
C172 plus.t4 a_n2044_n1088# 0.048897f
C173 plus.t13 a_n2044_n1088# 0.048897f
C174 plus.t10 a_n2044_n1088# 0.048897f
C175 plus.n1 a_n2044_n1088# 0.053884f
C176 plus.n2 a_n2044_n1088# 0.038482f
C177 plus.t2 a_n2044_n1088# 0.048897f
C178 plus.t12 a_n2044_n1088# 0.048897f
C179 plus.t6 a_n2044_n1088# 0.048897f
C180 plus.n3 a_n2044_n1088# 0.053706f
C181 plus.t1 a_n2044_n1088# 0.056126f
C182 plus.n4 a_n2044_n1088# 0.043854f
C183 plus.n5 a_n2044_n1088# 0.094831f
C184 plus.n6 a_n2044_n1088# 0.006544f
C185 plus.n7 a_n2044_n1088# 0.053884f
C186 plus.n8 a_n2044_n1088# 0.057405f
C187 plus.n9 a_n2044_n1088# 0.038392f
C188 plus.n10 a_n2044_n1088# 0.038482f
C189 plus.n11 a_n2044_n1088# 0.028839f
C190 plus.n12 a_n2044_n1088# 0.006544f
C191 plus.n13 a_n2044_n1088# 0.053706f
C192 plus.n14 a_n2044_n1088# 0.050861f
C193 plus.n15 a_n2044_n1088# 0.204375f
C194 plus.n16 a_n2044_n1088# 0.028839f
C195 plus.t11 a_n2044_n1088# 0.048897f
C196 plus.t8 a_n2044_n1088# 0.048897f
C197 plus.t0 a_n2044_n1088# 0.048897f
C198 plus.n17 a_n2044_n1088# 0.053884f
C199 plus.n18 a_n2044_n1088# 0.038482f
C200 plus.t9 a_n2044_n1088# 0.048897f
C201 plus.t3 a_n2044_n1088# 0.048897f
C202 plus.t7 a_n2044_n1088# 0.048897f
C203 plus.n19 a_n2044_n1088# 0.053706f
C204 plus.t5 a_n2044_n1088# 0.056126f
C205 plus.n20 a_n2044_n1088# 0.043854f
C206 plus.n21 a_n2044_n1088# 0.094831f
C207 plus.n22 a_n2044_n1088# 0.006544f
C208 plus.n23 a_n2044_n1088# 0.053884f
C209 plus.n24 a_n2044_n1088# 0.057405f
C210 plus.n25 a_n2044_n1088# 0.038392f
C211 plus.n26 a_n2044_n1088# 0.038482f
C212 plus.n27 a_n2044_n1088# 0.028839f
C213 plus.n28 a_n2044_n1088# 0.006544f
C214 plus.n29 a_n2044_n1088# 0.053706f
C215 plus.n30 a_n2044_n1088# 0.050861f
C216 plus.n31 a_n2044_n1088# 0.672174f
.ends

