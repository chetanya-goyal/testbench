* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X3 a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X4 drain_right.t5 minus.t0 source.t6 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X5 drain_right.t4 minus.t1 source.t9 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X6 drain_right.t3 minus.t2 source.t10 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X7 drain_left.t5 plus.t0 source.t1 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X8 drain_left.t4 plus.t1 source.t5 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X9 source.t8 minus.t3 drain_right.t2 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X10 drain_right.t1 minus.t4 source.t11 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X11 source.t7 minus.t5 drain_right.t0 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X12 drain_left.t3 plus.t2 source.t0 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X13 source.t2 plus.t3 drain_left.t2 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X14 source.t4 plus.t4 drain_left.t1 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X15 drain_left.t0 plus.t5 source.t3 a_n1620_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n5 minus.n4 161.3
R1 minus.n3 minus.n0 161.3
R2 minus.n11 minus.n10 161.3
R3 minus.n9 minus.n6 161.3
R4 minus.n1 minus.t4 102.716
R5 minus.n7 minus.t1 102.716
R6 minus.n2 minus.t3 79.2293
R7 minus.n4 minus.t2 79.2293
R8 minus.n8 minus.t5 79.2293
R9 minus.n10 minus.t0 79.2293
R10 minus.n1 minus.n0 44.8973
R11 minus.n7 minus.n6 44.8973
R12 minus.n4 minus.n3 33.5944
R13 minus.n10 minus.n9 33.5944
R14 minus.n12 minus.n5 27.1463
R15 minus.n2 minus.n1 18.1882
R16 minus.n8 minus.n7 18.1882
R17 minus.n3 minus.n2 14.6066
R18 minus.n9 minus.n8 14.6066
R19 minus.n12 minus.n11 6.72209
R20 minus.n5 minus.n0 0.189894
R21 minus.n11 minus.n6 0.189894
R22 minus minus.n12 0.188
R23 source.n0 source.t0 243.255
R24 source.n3 source.t11 243.255
R25 source.n11 source.t6 243.254
R26 source.n8 source.t1 243.254
R27 source.n2 source.n1 223.454
R28 source.n5 source.n4 223.454
R29 source.n10 source.n9 223.453
R30 source.n7 source.n6 223.453
R31 source.n9 source.t9 19.8005
R32 source.n9 source.t7 19.8005
R33 source.n6 source.t5 19.8005
R34 source.n6 source.t4 19.8005
R35 source.n1 source.t3 19.8005
R36 source.n1 source.t2 19.8005
R37 source.n4 source.t10 19.8005
R38 source.n4 source.t8 19.8005
R39 source.n7 source.n5 14.9027
R40 source.n12 source.n0 8.17853
R41 source.n12 source.n11 5.7505
R42 source.n5 source.n3 0.974638
R43 source.n2 source.n0 0.974638
R44 source.n8 source.n7 0.974638
R45 source.n11 source.n10 0.974638
R46 source.n3 source.n2 0.957397
R47 source.n10 source.n8 0.957397
R48 source source.n12 0.188
R49 drain_right.n1 drain_right.t4 260.608
R50 drain_right.n3 drain_right.t3 259.933
R51 drain_right.n3 drain_right.n2 241.107
R52 drain_right.n1 drain_right.n0 240.321
R53 drain_right drain_right.n1 21.1594
R54 drain_right.n0 drain_right.t0 19.8005
R55 drain_right.n0 drain_right.t5 19.8005
R56 drain_right.n2 drain_right.t2 19.8005
R57 drain_right.n2 drain_right.t1 19.8005
R58 drain_right drain_right.n3 6.14028
R59 plus.n3 plus.n0 161.3
R60 plus.n5 plus.n4 161.3
R61 plus.n9 plus.n6 161.3
R62 plus.n11 plus.n10 161.3
R63 plus.n1 plus.t5 102.716
R64 plus.n7 plus.t0 102.716
R65 plus.n4 plus.t2 79.2293
R66 plus.n2 plus.t3 79.2293
R67 plus.n10 plus.t1 79.2293
R68 plus.n8 plus.t4 79.2293
R69 plus.n7 plus.n6 44.8973
R70 plus.n1 plus.n0 44.8973
R71 plus.n4 plus.n3 33.5944
R72 plus.n10 plus.n9 33.5944
R73 plus plus.n11 25.1941
R74 plus.n8 plus.n7 18.1882
R75 plus.n2 plus.n1 18.1882
R76 plus.n3 plus.n2 14.6066
R77 plus.n9 plus.n8 14.6066
R78 plus plus.n5 8.19936
R79 plus.n5 plus.n0 0.189894
R80 plus.n11 plus.n6 0.189894
R81 drain_left.n3 drain_left.t0 260.906
R82 drain_left.n1 drain_left.t4 260.608
R83 drain_left.n1 drain_left.n0 240.321
R84 drain_left.n3 drain_left.n2 240.132
R85 drain_left drain_left.n1 21.7126
R86 drain_left.n0 drain_left.t1 19.8005
R87 drain_left.n0 drain_left.t5 19.8005
R88 drain_left.n2 drain_left.t2 19.8005
R89 drain_left.n2 drain_left.t3 19.8005
R90 drain_left drain_left.n3 6.62735
C0 drain_left source 2.63229f
C1 drain_right source 2.63296f
C2 plus source 1.04551f
C3 drain_left minus 0.179156f
C4 drain_right minus 0.704773f
C5 plus minus 3.12593f
C6 source minus 1.03161f
C7 drain_right drain_left 0.742213f
C8 drain_left plus 0.860234f
C9 drain_right plus 0.31914f
C10 drain_right a_n1620_n1088# 3.050789f
C11 drain_left a_n1620_n1088# 3.259773f
C12 source a_n1620_n1088# 2.086656f
C13 minus a_n1620_n1088# 5.261596f
C14 plus a_n1620_n1088# 5.908962f
C15 drain_left.t4 a_n1620_n1088# 0.086204f
C16 drain_left.t1 a_n1620_n1088# 0.013864f
C17 drain_left.t5 a_n1620_n1088# 0.013864f
C18 drain_left.n0 a_n1620_n1088# 0.054024f
C19 drain_left.n1 a_n1620_n1088# 0.824775f
C20 drain_left.t0 a_n1620_n1088# 0.086464f
C21 drain_left.t2 a_n1620_n1088# 0.013864f
C22 drain_left.t3 a_n1620_n1088# 0.013864f
C23 drain_left.n2 a_n1620_n1088# 0.05387f
C24 drain_left.n3 a_n1620_n1088# 0.580166f
C25 plus.n0 a_n1620_n1088# 0.139187f
C26 plus.t2 a_n1620_n1088# 0.087332f
C27 plus.t3 a_n1620_n1088# 0.087332f
C28 plus.t5 a_n1620_n1088# 0.106963f
C29 plus.n1 a_n1620_n1088# 0.069121f
C30 plus.n2 a_n1620_n1088# 0.087604f
C31 plus.n3 a_n1620_n1088# 0.007305f
C32 plus.n4 a_n1620_n1088# 0.084473f
C33 plus.n5 a_n1620_n1088# 0.238298f
C34 plus.n6 a_n1620_n1088# 0.139187f
C35 plus.t1 a_n1620_n1088# 0.087332f
C36 plus.t0 a_n1620_n1088# 0.106963f
C37 plus.n7 a_n1620_n1088# 0.069121f
C38 plus.t4 a_n1620_n1088# 0.087332f
C39 plus.n8 a_n1620_n1088# 0.087604f
C40 plus.n9 a_n1620_n1088# 0.007305f
C41 plus.n10 a_n1620_n1088# 0.084473f
C42 plus.n11 a_n1620_n1088# 0.690966f
C43 drain_right.t4 a_n1620_n1088# 0.088541f
C44 drain_right.t0 a_n1620_n1088# 0.014239f
C45 drain_right.t5 a_n1620_n1088# 0.014239f
C46 drain_right.n0 a_n1620_n1088# 0.055489f
C47 drain_right.n1 a_n1620_n1088# 0.812249f
C48 drain_right.t2 a_n1620_n1088# 0.014239f
C49 drain_right.t1 a_n1620_n1088# 0.014239f
C50 drain_right.n2 a_n1620_n1088# 0.056326f
C51 drain_right.t3 a_n1620_n1088# 0.088077f
C52 drain_right.n3 a_n1620_n1088# 0.610693f
C53 source.t0 a_n1620_n1088# 0.108394f
C54 source.n0 a_n1620_n1088# 0.526501f
C55 source.t3 a_n1620_n1088# 0.019475f
C56 source.t2 a_n1620_n1088# 0.019475f
C57 source.n1 a_n1620_n1088# 0.06316f
C58 source.n2 a_n1620_n1088# 0.304702f
C59 source.t11 a_n1620_n1088# 0.108394f
C60 source.n3 a_n1620_n1088# 0.312581f
C61 source.t10 a_n1620_n1088# 0.019475f
C62 source.t8 a_n1620_n1088# 0.019475f
C63 source.n4 a_n1620_n1088# 0.06316f
C64 source.n5 a_n1620_n1088# 0.800839f
C65 source.t5 a_n1620_n1088# 0.019475f
C66 source.t4 a_n1620_n1088# 0.019475f
C67 source.n6 a_n1620_n1088# 0.06316f
C68 source.n7 a_n1620_n1088# 0.800839f
C69 source.t1 a_n1620_n1088# 0.108394f
C70 source.n8 a_n1620_n1088# 0.312581f
C71 source.t9 a_n1620_n1088# 0.019475f
C72 source.t7 a_n1620_n1088# 0.019475f
C73 source.n9 a_n1620_n1088# 0.06316f
C74 source.n10 a_n1620_n1088# 0.304702f
C75 source.t6 a_n1620_n1088# 0.108394f
C76 source.n11 a_n1620_n1088# 0.439996f
C77 source.n12 a_n1620_n1088# 0.513756f
C78 minus.n0 a_n1620_n1088# 0.136324f
C79 minus.t4 a_n1620_n1088# 0.104763f
C80 minus.n1 a_n1620_n1088# 0.067699f
C81 minus.t3 a_n1620_n1088# 0.085536f
C82 minus.n2 a_n1620_n1088# 0.085802f
C83 minus.n3 a_n1620_n1088# 0.007155f
C84 minus.t2 a_n1620_n1088# 0.085536f
C85 minus.n4 a_n1620_n1088# 0.082735f
C86 minus.n5 a_n1620_n1088# 0.695608f
C87 minus.n6 a_n1620_n1088# 0.136324f
C88 minus.t1 a_n1620_n1088# 0.104763f
C89 minus.n7 a_n1620_n1088# 0.067699f
C90 minus.t5 a_n1620_n1088# 0.085536f
C91 minus.n8 a_n1620_n1088# 0.085802f
C92 minus.n9 a_n1620_n1088# 0.007155f
C93 minus.t0 a_n1620_n1088# 0.085536f
C94 minus.n10 a_n1620_n1088# 0.082735f
C95 minus.n11 a_n1620_n1088# 0.222469f
C96 minus.n12 a_n1620_n1088# 0.850117f
.ends

