* NGSPICE file created from diffpair505.ext - technology: sky130A

.subckt diffpair505 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t23 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X1 drain_left.t10 plus.t1 source.t20 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X2 source.t16 plus.t2 drain_left.t9 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X3 drain_right.t11 minus.t0 source.t9 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X4 drain_left.t8 plus.t3 source.t21 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X5 source.t0 minus.t1 drain_right.t10 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X6 source.t8 minus.t2 drain_right.t9 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X7 source.t11 minus.t3 drain_right.t8 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 source.t13 plus.t4 drain_left.t7 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X9 a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X10 a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X11 source.t18 plus.t5 drain_left.t6 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X12 source.t1 minus.t4 drain_right.t7 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X13 drain_right.t6 minus.t5 source.t2 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X14 drain_left.t5 plus.t6 source.t22 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X15 source.t3 minus.t6 drain_right.t5 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X16 source.t19 plus.t7 drain_left.t4 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X17 source.t17 plus.t8 drain_left.t3 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X18 a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X19 drain_left.t2 plus.t9 source.t15 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X20 drain_right.t4 minus.t7 source.t7 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X21 a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X22 drain_right.t3 minus.t8 source.t10 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X23 drain_right.t2 minus.t9 source.t4 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X24 drain_right.t1 minus.t10 source.t6 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X25 source.t14 plus.t10 drain_left.t1 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X26 drain_left.t0 plus.t11 source.t12 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X27 source.t5 minus.t11 drain_right.t0 a_n1528_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
R0 plus.n2 plus.t5 1600.53
R1 plus.n13 plus.t11 1600.53
R2 plus.n17 plus.t3 1600.53
R3 plus.n28 plus.t2 1600.53
R4 plus.n3 plus.t1 1571.32
R5 plus.n4 plus.t8 1571.32
R6 plus.n10 plus.t0 1571.32
R7 plus.n12 plus.t7 1571.32
R8 plus.n19 plus.t10 1571.32
R9 plus.n18 plus.t9 1571.32
R10 plus.n25 plus.t4 1571.32
R11 plus.n27 plus.t6 1571.32
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 29.8627
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 13.2164
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n5 source.t18 45.521
R53 source.n6 source.t10 45.521
R54 source.n11 source.t1 45.521
R55 source.n23 source.t9 45.5208
R56 source.n18 source.t11 45.5208
R57 source.n17 source.t21 45.5208
R58 source.n12 source.t16 45.5208
R59 source.n0 source.t12 45.5208
R60 source.n2 source.n1 44.201
R61 source.n4 source.n3 44.201
R62 source.n8 source.n7 44.201
R63 source.n10 source.n9 44.201
R64 source.n22 source.n21 44.2008
R65 source.n20 source.n19 44.2008
R66 source.n16 source.n15 44.2008
R67 source.n14 source.n13 44.2008
R68 source.n12 source.n11 24.0605
R69 source.n24 source.n0 18.5475
R70 source.n24 source.n23 5.51343
R71 source.n21 source.t4 1.3205
R72 source.n21 source.t3 1.3205
R73 source.n19 source.t2 1.3205
R74 source.n19 source.t5 1.3205
R75 source.n15 source.t15 1.3205
R76 source.n15 source.t14 1.3205
R77 source.n13 source.t22 1.3205
R78 source.n13 source.t13 1.3205
R79 source.n1 source.t23 1.3205
R80 source.n1 source.t19 1.3205
R81 source.n3 source.t20 1.3205
R82 source.n3 source.t17 1.3205
R83 source.n7 source.t7 1.3205
R84 source.n7 source.t8 1.3205
R85 source.n9 source.t6 1.3205
R86 source.n9 source.t0 1.3205
R87 source.n11 source.n10 0.5005
R88 source.n10 source.n8 0.5005
R89 source.n8 source.n6 0.5005
R90 source.n5 source.n4 0.5005
R91 source.n4 source.n2 0.5005
R92 source.n2 source.n0 0.5005
R93 source.n14 source.n12 0.5005
R94 source.n16 source.n14 0.5005
R95 source.n17 source.n16 0.5005
R96 source.n20 source.n18 0.5005
R97 source.n22 source.n20 0.5005
R98 source.n23 source.n22 0.5005
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 61.3798
R103 drain_left.n3 drain_left.n2 61.3242
R104 drain_left.n3 drain_left.n0 61.3242
R105 drain_left.n6 drain_left.n5 60.8798
R106 drain_left.n8 drain_left.n7 60.8796
R107 drain_left.n3 drain_left.n1 60.8796
R108 drain_left drain_left.n3 32.1398
R109 drain_left drain_left.n8 6.15322
R110 drain_left.n1 drain_left.t7 1.3205
R111 drain_left.n1 drain_left.t2 1.3205
R112 drain_left.n2 drain_left.t1 1.3205
R113 drain_left.n2 drain_left.t8 1.3205
R114 drain_left.n0 drain_left.t9 1.3205
R115 drain_left.n0 drain_left.t5 1.3205
R116 drain_left.n7 drain_left.t4 1.3205
R117 drain_left.n7 drain_left.t0 1.3205
R118 drain_left.n5 drain_left.t3 1.3205
R119 drain_left.n5 drain_left.t11 1.3205
R120 drain_left.n4 drain_left.t6 1.3205
R121 drain_left.n4 drain_left.t10 1.3205
R122 drain_left.n8 drain_left.n6 0.5005
R123 minus.n13 minus.t4 1600.53
R124 minus.n2 minus.t8 1600.53
R125 minus.n28 minus.t0 1600.53
R126 minus.n17 minus.t3 1600.53
R127 minus.n12 minus.t10 1571.32
R128 minus.n10 minus.t1 1571.32
R129 minus.n3 minus.t7 1571.32
R130 minus.n4 minus.t2 1571.32
R131 minus.n27 minus.t6 1571.32
R132 minus.n25 minus.t9 1571.32
R133 minus.n19 minus.t11 1571.32
R134 minus.n18 minus.t5 1571.32
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 67.1884
R150 minus.n5 minus.n3 67.1884
R151 minus.n20 minus.n19 67.1884
R152 minus.n26 minus.n25 67.1884
R153 minus.n13 minus.n12 55.5035
R154 minus.n4 minus.n2 55.5035
R155 minus.n18 minus.n17 55.5035
R156 minus.n28 minus.n27 55.5035
R157 minus.n30 minus.n14 37.1179
R158 minus.n12 minus.n11 17.5278
R159 minus.n5 minus.n4 17.5278
R160 minus.n20 minus.n18 17.5278
R161 minus.n27 minus.n26 17.5278
R162 minus.n30 minus.n29 6.43611
R163 minus.n10 minus.n9 5.84292
R164 minus.n3 minus.n1 5.84292
R165 minus.n19 minus.n16 5.84292
R166 minus.n25 minus.n24 5.84292
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 61.3796
R177 drain_right.n3 drain_right.n2 61.3242
R178 drain_right.n3 drain_right.n0 61.3242
R179 drain_right.n6 drain_right.n5 60.8798
R180 drain_right.n8 drain_right.n7 60.8798
R181 drain_right.n3 drain_right.n1 60.8796
R182 drain_right drain_right.n3 31.5866
R183 drain_right drain_right.n8 6.15322
R184 drain_right.n1 drain_right.t0 1.3205
R185 drain_right.n1 drain_right.t2 1.3205
R186 drain_right.n2 drain_right.t5 1.3205
R187 drain_right.n2 drain_right.t11 1.3205
R188 drain_right.n0 drain_right.t8 1.3205
R189 drain_right.n0 drain_right.t6 1.3205
R190 drain_right.n4 drain_right.t9 1.3205
R191 drain_right.n4 drain_right.t3 1.3205
R192 drain_right.n5 drain_right.t10 1.3205
R193 drain_right.n5 drain_right.t4 1.3205
R194 drain_right.n7 drain_right.t7 1.3205
R195 drain_right.n7 drain_right.t1 1.3205
R196 drain_right.n8 drain_right.n6 0.5005
C0 drain_right drain_left 0.751086f
C1 minus drain_left 0.171004f
C2 plus drain_left 5.15185f
C3 minus drain_right 5.00568f
C4 plus drain_right 0.300071f
C5 source drain_left 31.4093f
C6 minus plus 5.61778f
C7 source drain_right 31.408699f
C8 source minus 4.46395f
C9 source plus 4.47799f
C10 drain_right a_n1528_n3888# 6.93378f
C11 drain_left a_n1528_n3888# 7.186201f
C12 source a_n1528_n3888# 10.173927f
C13 minus a_n1528_n3888# 6.124974f
C14 plus a_n1528_n3888# 8.360909f
C15 drain_right.t8 a_n1528_n3888# 0.424203f
C16 drain_right.t6 a_n1528_n3888# 0.424203f
C17 drain_right.n0 a_n1528_n3888# 3.83733f
C18 drain_right.t0 a_n1528_n3888# 0.424203f
C19 drain_right.t2 a_n1528_n3888# 0.424203f
C20 drain_right.n1 a_n1528_n3888# 3.83429f
C21 drain_right.t5 a_n1528_n3888# 0.424203f
C22 drain_right.t11 a_n1528_n3888# 0.424203f
C23 drain_right.n2 a_n1528_n3888# 3.83733f
C24 drain_right.n3 a_n1528_n3888# 2.99597f
C25 drain_right.t9 a_n1528_n3888# 0.424203f
C26 drain_right.t3 a_n1528_n3888# 0.424203f
C27 drain_right.n4 a_n1528_n3888# 3.83773f
C28 drain_right.t10 a_n1528_n3888# 0.424203f
C29 drain_right.t4 a_n1528_n3888# 0.424203f
C30 drain_right.n5 a_n1528_n3888# 3.8343f
C31 drain_right.n6 a_n1528_n3888# 0.827844f
C32 drain_right.t7 a_n1528_n3888# 0.424203f
C33 drain_right.t1 a_n1528_n3888# 0.424203f
C34 drain_right.n7 a_n1528_n3888# 3.8343f
C35 drain_right.n8 a_n1528_n3888# 0.70383f
C36 minus.n0 a_n1528_n3888# 0.054096f
C37 minus.t4 a_n1528_n3888# 0.576334f
C38 minus.t10 a_n1528_n3888# 0.572301f
C39 minus.t1 a_n1528_n3888# 0.572301f
C40 minus.n1 a_n1528_n3888# 0.01928f
C41 minus.t8 a_n1528_n3888# 0.576334f
C42 minus.n2 a_n1528_n3888# 0.237587f
C43 minus.t7 a_n1528_n3888# 0.572301f
C44 minus.n3 a_n1528_n3888# 0.222604f
C45 minus.t2 a_n1528_n3888# 0.572301f
C46 minus.n4 a_n1528_n3888# 0.222604f
C47 minus.n5 a_n1528_n3888# 0.020614f
C48 minus.n6 a_n1528_n3888# 0.113126f
C49 minus.n7 a_n1528_n3888# 0.054096f
C50 minus.n8 a_n1528_n3888# 0.054096f
C51 minus.n9 a_n1528_n3888# 0.01928f
C52 minus.n10 a_n1528_n3888# 0.222604f
C53 minus.n11 a_n1528_n3888# 0.020614f
C54 minus.n12 a_n1528_n3888# 0.222604f
C55 minus.n13 a_n1528_n3888# 0.237517f
C56 minus.n14 a_n1528_n3888# 1.98567f
C57 minus.n15 a_n1528_n3888# 0.054096f
C58 minus.t6 a_n1528_n3888# 0.572301f
C59 minus.t9 a_n1528_n3888# 0.572301f
C60 minus.n16 a_n1528_n3888# 0.01928f
C61 minus.t3 a_n1528_n3888# 0.576334f
C62 minus.n17 a_n1528_n3888# 0.237587f
C63 minus.t5 a_n1528_n3888# 0.572301f
C64 minus.n18 a_n1528_n3888# 0.222604f
C65 minus.t11 a_n1528_n3888# 0.572301f
C66 minus.n19 a_n1528_n3888# 0.222604f
C67 minus.n20 a_n1528_n3888# 0.020614f
C68 minus.n21 a_n1528_n3888# 0.113126f
C69 minus.n22 a_n1528_n3888# 0.054096f
C70 minus.n23 a_n1528_n3888# 0.054096f
C71 minus.n24 a_n1528_n3888# 0.01928f
C72 minus.n25 a_n1528_n3888# 0.222604f
C73 minus.n26 a_n1528_n3888# 0.020614f
C74 minus.n27 a_n1528_n3888# 0.222604f
C75 minus.t0 a_n1528_n3888# 0.576334f
C76 minus.n28 a_n1528_n3888# 0.237517f
C77 minus.n29 a_n1528_n3888# 0.345499f
C78 minus.n30 a_n1528_n3888# 2.40812f
C79 drain_left.t9 a_n1528_n3888# 0.424899f
C80 drain_left.t5 a_n1528_n3888# 0.424899f
C81 drain_left.n0 a_n1528_n3888# 3.84363f
C82 drain_left.t7 a_n1528_n3888# 0.424899f
C83 drain_left.t2 a_n1528_n3888# 0.424899f
C84 drain_left.n1 a_n1528_n3888# 3.84059f
C85 drain_left.t1 a_n1528_n3888# 0.424899f
C86 drain_left.t8 a_n1528_n3888# 0.424899f
C87 drain_left.n2 a_n1528_n3888# 3.84363f
C88 drain_left.n3 a_n1528_n3888# 3.0759f
C89 drain_left.t6 a_n1528_n3888# 0.424899f
C90 drain_left.t10 a_n1528_n3888# 0.424899f
C91 drain_left.n4 a_n1528_n3888# 3.84404f
C92 drain_left.t3 a_n1528_n3888# 0.424899f
C93 drain_left.t11 a_n1528_n3888# 0.424899f
C94 drain_left.n5 a_n1528_n3888# 3.84059f
C95 drain_left.n6 a_n1528_n3888# 0.82919f
C96 drain_left.t4 a_n1528_n3888# 0.424899f
C97 drain_left.t0 a_n1528_n3888# 0.424899f
C98 drain_left.n7 a_n1528_n3888# 3.84058f
C99 drain_left.n8 a_n1528_n3888# 0.704999f
C100 source.t12 a_n1528_n3888# 3.71093f
C101 source.n0 a_n1528_n3888# 1.71257f
C102 source.t23 a_n1528_n3888# 0.331138f
C103 source.t19 a_n1528_n3888# 0.331138f
C104 source.n1 a_n1528_n3888# 2.90877f
C105 source.n2 a_n1528_n3888# 0.365189f
C106 source.t20 a_n1528_n3888# 0.331138f
C107 source.t17 a_n1528_n3888# 0.331138f
C108 source.n3 a_n1528_n3888# 2.90877f
C109 source.n4 a_n1528_n3888# 0.365189f
C110 source.t18 a_n1528_n3888# 3.71094f
C111 source.n5 a_n1528_n3888# 0.463407f
C112 source.t10 a_n1528_n3888# 3.71094f
C113 source.n6 a_n1528_n3888# 0.463407f
C114 source.t7 a_n1528_n3888# 0.331138f
C115 source.t8 a_n1528_n3888# 0.331138f
C116 source.n7 a_n1528_n3888# 2.90877f
C117 source.n8 a_n1528_n3888# 0.365189f
C118 source.t6 a_n1528_n3888# 0.331138f
C119 source.t0 a_n1528_n3888# 0.331138f
C120 source.n9 a_n1528_n3888# 2.90877f
C121 source.n10 a_n1528_n3888# 0.365189f
C122 source.t1 a_n1528_n3888# 3.71094f
C123 source.n11 a_n1528_n3888# 2.17553f
C124 source.t16 a_n1528_n3888# 3.71093f
C125 source.n12 a_n1528_n3888# 2.17553f
C126 source.t22 a_n1528_n3888# 0.331138f
C127 source.t13 a_n1528_n3888# 0.331138f
C128 source.n13 a_n1528_n3888# 2.90876f
C129 source.n14 a_n1528_n3888# 0.365192f
C130 source.t15 a_n1528_n3888# 0.331138f
C131 source.t14 a_n1528_n3888# 0.331138f
C132 source.n15 a_n1528_n3888# 2.90876f
C133 source.n16 a_n1528_n3888# 0.365192f
C134 source.t21 a_n1528_n3888# 3.71093f
C135 source.n17 a_n1528_n3888# 0.463411f
C136 source.t11 a_n1528_n3888# 3.71093f
C137 source.n18 a_n1528_n3888# 0.463411f
C138 source.t2 a_n1528_n3888# 0.331138f
C139 source.t5 a_n1528_n3888# 0.331138f
C140 source.n19 a_n1528_n3888# 2.90876f
C141 source.n20 a_n1528_n3888# 0.365192f
C142 source.t4 a_n1528_n3888# 0.331138f
C143 source.t3 a_n1528_n3888# 0.331138f
C144 source.n21 a_n1528_n3888# 2.90876f
C145 source.n22 a_n1528_n3888# 0.365192f
C146 source.t9 a_n1528_n3888# 3.71093f
C147 source.n23 a_n1528_n3888# 0.618004f
C148 source.n24 a_n1528_n3888# 2.04036f
C149 plus.n0 a_n1528_n3888# 0.055213f
C150 plus.t7 a_n1528_n3888# 0.584113f
C151 plus.t0 a_n1528_n3888# 0.584113f
C152 plus.n1 a_n1528_n3888# 0.019677f
C153 plus.t5 a_n1528_n3888# 0.588229f
C154 plus.n2 a_n1528_n3888# 0.24249f
C155 plus.t1 a_n1528_n3888# 0.584113f
C156 plus.n3 a_n1528_n3888# 0.227198f
C157 plus.t8 a_n1528_n3888# 0.584113f
C158 plus.n4 a_n1528_n3888# 0.227198f
C159 plus.n5 a_n1528_n3888# 0.021039f
C160 plus.n6 a_n1528_n3888# 0.115461f
C161 plus.n7 a_n1528_n3888# 0.055213f
C162 plus.n8 a_n1528_n3888# 0.055213f
C163 plus.n9 a_n1528_n3888# 0.019677f
C164 plus.n10 a_n1528_n3888# 0.227198f
C165 plus.n11 a_n1528_n3888# 0.021039f
C166 plus.n12 a_n1528_n3888# 0.227198f
C167 plus.t11 a_n1528_n3888# 0.588229f
C168 plus.n13 a_n1528_n3888# 0.24242f
C169 plus.n14 a_n1528_n3888# 0.689391f
C170 plus.n15 a_n1528_n3888# 0.055213f
C171 plus.t2 a_n1528_n3888# 0.588229f
C172 plus.t6 a_n1528_n3888# 0.584113f
C173 plus.t4 a_n1528_n3888# 0.584113f
C174 plus.n16 a_n1528_n3888# 0.019677f
C175 plus.t3 a_n1528_n3888# 0.588229f
C176 plus.n17 a_n1528_n3888# 0.24249f
C177 plus.t9 a_n1528_n3888# 0.584113f
C178 plus.n18 a_n1528_n3888# 0.227198f
C179 plus.t10 a_n1528_n3888# 0.584113f
C180 plus.n19 a_n1528_n3888# 0.227198f
C181 plus.n20 a_n1528_n3888# 0.021039f
C182 plus.n21 a_n1528_n3888# 0.115461f
C183 plus.n22 a_n1528_n3888# 0.055213f
C184 plus.n23 a_n1528_n3888# 0.055213f
C185 plus.n24 a_n1528_n3888# 0.019677f
C186 plus.n25 a_n1528_n3888# 0.227198f
C187 plus.n26 a_n1528_n3888# 0.021039f
C188 plus.n27 a_n1528_n3888# 0.227198f
C189 plus.n28 a_n1528_n3888# 0.24242f
C190 plus.n29 a_n1528_n3888# 1.6604f
.ends

