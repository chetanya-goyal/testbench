* NGSPICE file created from diffpair193.ext - technology: sky130A

.subckt diffpair193 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t14 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 drain_right.t6 minus.t1 source.t13 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X2 source.t15 plus.t0 drain_left.t7 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X3 drain_left.t6 plus.t1 source.t0 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X4 a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X5 source.t12 minus.t2 drain_right.t5 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X6 source.t1 plus.t2 drain_left.t5 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X7 a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X8 drain_left.t4 plus.t3 source.t6 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X9 drain_right.t4 minus.t3 source.t11 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X10 source.t7 minus.t4 drain_right.t3 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X11 a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X12 drain_right.t2 minus.t5 source.t10 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X13 source.t5 plus.t4 drain_left.t3 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X14 drain_left.t2 plus.t5 source.t2 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X15 source.t8 minus.t6 drain_right.t1 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X16 source.t9 minus.t7 drain_right.t0 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X17 source.t4 plus.t6 drain_left.t1 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X18 a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X19 drain_left.t0 plus.t7 source.t3 a_n1346_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
R0 minus.n7 minus.t4 373.916
R1 minus.n2 minus.t5 373.916
R2 minus.n16 minus.t3 373.916
R3 minus.n11 minus.t2 373.916
R4 minus.n6 minus.t1 345.433
R5 minus.n1 minus.t6 345.433
R6 minus.n15 minus.t7 345.433
R7 minus.n10 minus.t0 345.433
R8 minus.n3 minus.n2 161.489
R9 minus.n12 minus.n11 161.489
R10 minus.n8 minus.n7 161.3
R11 minus.n5 minus.n0 161.3
R12 minus.n4 minus.n3 161.3
R13 minus.n17 minus.n16 161.3
R14 minus.n14 minus.n9 161.3
R15 minus.n13 minus.n12 161.3
R16 minus.n5 minus.n4 73.0308
R17 minus.n14 minus.n13 73.0308
R18 minus.n7 minus.n6 63.5369
R19 minus.n2 minus.n1 63.5369
R20 minus.n11 minus.n10 63.5369
R21 minus.n16 minus.n15 63.5369
R22 minus.n18 minus.n8 27.3641
R23 minus.n6 minus.n5 9.49444
R24 minus.n4 minus.n1 9.49444
R25 minus.n13 minus.n10 9.49444
R26 minus.n15 minus.n14 9.49444
R27 minus.n18 minus.n17 6.46262
R28 minus.n8 minus.n0 0.189894
R29 minus.n3 minus.n0 0.189894
R30 minus.n12 minus.n9 0.189894
R31 minus.n17 minus.n9 0.189894
R32 minus minus.n18 0.188
R33 source.n0 source.t3 69.6943
R34 source.n3 source.t15 69.6943
R35 source.n4 source.t10 69.6943
R36 source.n7 source.t7 69.6943
R37 source.n15 source.t11 69.6942
R38 source.n12 source.t12 69.6942
R39 source.n11 source.t0 69.6942
R40 source.n8 source.t1 69.6942
R41 source.n2 source.n1 63.0943
R42 source.n6 source.n5 63.0943
R43 source.n14 source.n13 63.0942
R44 source.n10 source.n9 63.0942
R45 source.n8 source.n7 15.0126
R46 source.n16 source.n0 9.47816
R47 source.n13 source.t14 6.6005
R48 source.n13 source.t9 6.6005
R49 source.n9 source.t2 6.6005
R50 source.n9 source.t4 6.6005
R51 source.n1 source.t6 6.6005
R52 source.n1 source.t5 6.6005
R53 source.n5 source.t13 6.6005
R54 source.n5 source.t8 6.6005
R55 source.n16 source.n15 5.53498
R56 source.n7 source.n6 0.543603
R57 source.n6 source.n4 0.543603
R58 source.n3 source.n2 0.543603
R59 source.n2 source.n0 0.543603
R60 source.n10 source.n8 0.543603
R61 source.n11 source.n10 0.543603
R62 source.n14 source.n12 0.543603
R63 source.n15 source.n14 0.543603
R64 source.n4 source.n3 0.470328
R65 source.n12 source.n11 0.470328
R66 source source.n16 0.188
R67 drain_right.n5 drain_right.n3 80.3162
R68 drain_right.n2 drain_right.n1 79.9892
R69 drain_right.n2 drain_right.n0 79.9892
R70 drain_right.n5 drain_right.n4 79.7731
R71 drain_right drain_right.n2 21.8965
R72 drain_right.n1 drain_right.t0 6.6005
R73 drain_right.n1 drain_right.t4 6.6005
R74 drain_right.n0 drain_right.t5 6.6005
R75 drain_right.n0 drain_right.t7 6.6005
R76 drain_right.n3 drain_right.t1 6.6005
R77 drain_right.n3 drain_right.t2 6.6005
R78 drain_right.n4 drain_right.t3 6.6005
R79 drain_right.n4 drain_right.t6 6.6005
R80 drain_right drain_right.n5 6.19632
R81 plus.n2 plus.t0 373.916
R82 plus.n7 plus.t7 373.916
R83 plus.n11 plus.t1 373.916
R84 plus.n16 plus.t2 373.916
R85 plus.n1 plus.t3 345.433
R86 plus.n6 plus.t4 345.433
R87 plus.n10 plus.t6 345.433
R88 plus.n15 plus.t5 345.433
R89 plus.n3 plus.n2 161.489
R90 plus.n12 plus.n11 161.489
R91 plus.n4 plus.n3 161.3
R92 plus.n5 plus.n0 161.3
R93 plus.n8 plus.n7 161.3
R94 plus.n13 plus.n12 161.3
R95 plus.n14 plus.n9 161.3
R96 plus.n17 plus.n16 161.3
R97 plus.n5 plus.n4 73.0308
R98 plus.n14 plus.n13 73.0308
R99 plus.n2 plus.n1 63.5369
R100 plus.n7 plus.n6 63.5369
R101 plus.n16 plus.n15 63.5369
R102 plus.n11 plus.n10 63.5369
R103 plus plus.n17 24.6543
R104 plus.n4 plus.n1 9.49444
R105 plus.n6 plus.n5 9.49444
R106 plus.n15 plus.n14 9.49444
R107 plus.n13 plus.n10 9.49444
R108 plus plus.n8 8.69747
R109 plus.n3 plus.n0 0.189894
R110 plus.n8 plus.n0 0.189894
R111 plus.n17 plus.n9 0.189894
R112 plus.n12 plus.n9 0.189894
R113 drain_left.n5 drain_left.n3 80.3162
R114 drain_left.n2 drain_left.n1 79.9892
R115 drain_left.n2 drain_left.n0 79.9892
R116 drain_left.n5 drain_left.n4 79.7731
R117 drain_left drain_left.n2 22.4498
R118 drain_left.n1 drain_left.t1 6.6005
R119 drain_left.n1 drain_left.t6 6.6005
R120 drain_left.n0 drain_left.t5 6.6005
R121 drain_left.n0 drain_left.t2 6.6005
R122 drain_left.n4 drain_left.t3 6.6005
R123 drain_left.n4 drain_left.t0 6.6005
R124 drain_left.n3 drain_left.t7 6.6005
R125 drain_left.n3 drain_left.t4 6.6005
R126 drain_left drain_left.n5 6.19632
C0 source minus 1.11997f
C1 drain_left minus 0.175592f
C2 drain_right minus 1.10491f
C3 plus source 1.13397f
C4 plus drain_left 1.2321f
C5 drain_left source 5.5088f
C6 plus drain_right 0.286118f
C7 drain_right source 5.50799f
C8 drain_right drain_left 0.630082f
C9 plus minus 3.17198f
C10 drain_right a_n1346_n1488# 3.35206f
C11 drain_left a_n1346_n1488# 3.51793f
C12 source a_n1346_n1488# 3.458569f
C13 minus a_n1346_n1488# 4.476064f
C14 plus a_n1346_n1488# 5.174556f
C15 drain_left.t5 a_n1346_n1488# 0.058931f
C16 drain_left.t2 a_n1346_n1488# 0.058931f
C17 drain_left.n0 a_n1346_n1488# 0.425738f
C18 drain_left.t1 a_n1346_n1488# 0.058931f
C19 drain_left.t6 a_n1346_n1488# 0.058931f
C20 drain_left.n1 a_n1346_n1488# 0.425738f
C21 drain_left.n2 a_n1346_n1488# 1.17251f
C22 drain_left.t7 a_n1346_n1488# 0.058931f
C23 drain_left.t4 a_n1346_n1488# 0.058931f
C24 drain_left.n3 a_n1346_n1488# 0.427005f
C25 drain_left.t3 a_n1346_n1488# 0.058931f
C26 drain_left.t0 a_n1346_n1488# 0.058931f
C27 drain_left.n4 a_n1346_n1488# 0.425004f
C28 drain_left.n5 a_n1346_n1488# 0.78689f
C29 plus.n0 a_n1346_n1488# 0.033027f
C30 plus.t4 a_n1346_n1488# 0.086078f
C31 plus.t3 a_n1346_n1488# 0.086078f
C32 plus.n1 a_n1346_n1488# 0.04998f
C33 plus.t0 a_n1346_n1488# 0.089877f
C34 plus.n2 a_n1346_n1488# 0.059726f
C35 plus.n3 a_n1346_n1488# 0.069879f
C36 plus.n4 a_n1346_n1488# 0.01228f
C37 plus.n5 a_n1346_n1488# 0.01228f
C38 plus.n6 a_n1346_n1488# 0.04998f
C39 plus.t7 a_n1346_n1488# 0.089877f
C40 plus.n7 a_n1346_n1488# 0.059682f
C41 plus.n8 a_n1346_n1488# 0.243641f
C42 plus.n9 a_n1346_n1488# 0.033027f
C43 plus.t2 a_n1346_n1488# 0.089877f
C44 plus.t5 a_n1346_n1488# 0.086078f
C45 plus.t6 a_n1346_n1488# 0.086078f
C46 plus.n10 a_n1346_n1488# 0.04998f
C47 plus.t1 a_n1346_n1488# 0.089877f
C48 plus.n11 a_n1346_n1488# 0.059726f
C49 plus.n12 a_n1346_n1488# 0.069879f
C50 plus.n13 a_n1346_n1488# 0.01228f
C51 plus.n14 a_n1346_n1488# 0.01228f
C52 plus.n15 a_n1346_n1488# 0.04998f
C53 plus.n16 a_n1346_n1488# 0.059682f
C54 plus.n17 a_n1346_n1488# 0.689864f
C55 drain_right.t5 a_n1346_n1488# 0.059991f
C56 drain_right.t7 a_n1346_n1488# 0.059991f
C57 drain_right.n0 a_n1346_n1488# 0.433401f
C58 drain_right.t0 a_n1346_n1488# 0.059991f
C59 drain_right.t4 a_n1346_n1488# 0.059991f
C60 drain_right.n1 a_n1346_n1488# 0.433401f
C61 drain_right.n2 a_n1346_n1488# 1.14315f
C62 drain_right.t1 a_n1346_n1488# 0.059991f
C63 drain_right.t2 a_n1346_n1488# 0.059991f
C64 drain_right.n3 a_n1346_n1488# 0.434691f
C65 drain_right.t3 a_n1346_n1488# 0.059991f
C66 drain_right.t6 a_n1346_n1488# 0.059991f
C67 drain_right.n4 a_n1346_n1488# 0.432653f
C68 drain_right.n5 a_n1346_n1488# 0.801052f
C69 source.t3 a_n1346_n1488# 0.440049f
C70 source.n0 a_n1346_n1488# 0.600374f
C71 source.t6 a_n1346_n1488# 0.052994f
C72 source.t5 a_n1346_n1488# 0.052994f
C73 source.n1 a_n1346_n1488# 0.336009f
C74 source.n2 a_n1346_n1488# 0.272966f
C75 source.t15 a_n1346_n1488# 0.440049f
C76 source.n3 a_n1346_n1488# 0.308177f
C77 source.t10 a_n1346_n1488# 0.440049f
C78 source.n4 a_n1346_n1488# 0.308177f
C79 source.t13 a_n1346_n1488# 0.052994f
C80 source.t8 a_n1346_n1488# 0.052994f
C81 source.n5 a_n1346_n1488# 0.336009f
C82 source.n6 a_n1346_n1488# 0.272966f
C83 source.t7 a_n1346_n1488# 0.440049f
C84 source.n7 a_n1346_n1488# 0.83338f
C85 source.t1 a_n1346_n1488# 0.440047f
C86 source.n8 a_n1346_n1488# 0.833383f
C87 source.t2 a_n1346_n1488# 0.052994f
C88 source.t4 a_n1346_n1488# 0.052994f
C89 source.n9 a_n1346_n1488# 0.336007f
C90 source.n10 a_n1346_n1488# 0.272969f
C91 source.t0 a_n1346_n1488# 0.440047f
C92 source.n11 a_n1346_n1488# 0.308179f
C93 source.t12 a_n1346_n1488# 0.440047f
C94 source.n12 a_n1346_n1488# 0.308179f
C95 source.t14 a_n1346_n1488# 0.052994f
C96 source.t9 a_n1346_n1488# 0.052994f
C97 source.n13 a_n1346_n1488# 0.336007f
C98 source.n14 a_n1346_n1488# 0.272969f
C99 source.t11 a_n1346_n1488# 0.440047f
C100 source.n15 a_n1346_n1488# 0.434365f
C101 source.n16 a_n1346_n1488# 0.647923f
C102 minus.n0 a_n1346_n1488# 0.032352f
C103 minus.t4 a_n1346_n1488# 0.088039f
C104 minus.t1 a_n1346_n1488# 0.084318f
C105 minus.t6 a_n1346_n1488# 0.084318f
C106 minus.n1 a_n1346_n1488# 0.048959f
C107 minus.t5 a_n1346_n1488# 0.088039f
C108 minus.n2 a_n1346_n1488# 0.058505f
C109 minus.n3 a_n1346_n1488# 0.06845f
C110 minus.n4 a_n1346_n1488# 0.012029f
C111 minus.n5 a_n1346_n1488# 0.012029f
C112 minus.n6 a_n1346_n1488# 0.048959f
C113 minus.n7 a_n1346_n1488# 0.058462f
C114 minus.n8 a_n1346_n1488# 0.715309f
C115 minus.n9 a_n1346_n1488# 0.032352f
C116 minus.t7 a_n1346_n1488# 0.084318f
C117 minus.t0 a_n1346_n1488# 0.084318f
C118 minus.n10 a_n1346_n1488# 0.048959f
C119 minus.t2 a_n1346_n1488# 0.088039f
C120 minus.n11 a_n1346_n1488# 0.058505f
C121 minus.n12 a_n1346_n1488# 0.06845f
C122 minus.n13 a_n1346_n1488# 0.012029f
C123 minus.n14 a_n1346_n1488# 0.012029f
C124 minus.n15 a_n1346_n1488# 0.048959f
C125 minus.t3 a_n1346_n1488# 0.088039f
C126 minus.n16 a_n1346_n1488# 0.058462f
C127 minus.n17 a_n1346_n1488# 0.208652f
C128 minus.n18 a_n1346_n1488# 0.885878f
.ends

