* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t11 minus.t0 drain_right.t0 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X1 a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X2 source.t0 plus.t0 drain_left.t5 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X4 a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X5 drain_right.t4 minus.t1 source.t10 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X6 source.t9 minus.t2 drain_right.t3 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X7 drain_right.t2 minus.t3 source.t8 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X8 a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X9 drain_right.t1 minus.t4 source.t7 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X10 drain_left.t4 plus.t1 source.t2 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X11 drain_right.t5 minus.t5 source.t6 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X12 source.t5 plus.t2 drain_left.t3 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X13 drain_left.t2 plus.t3 source.t3 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X14 drain_left.t1 plus.t4 source.t1 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X15 drain_left.t0 plus.t5 source.t4 a_n1620_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n5 minus.n4 161.3
R1 minus.n3 minus.n0 161.3
R2 minus.n11 minus.n10 161.3
R3 minus.n9 minus.n6 161.3
R4 minus.n1 minus.t3 132.84
R5 minus.n7 minus.t4 132.84
R6 minus.n2 minus.t2 109.355
R7 minus.n4 minus.t1 109.355
R8 minus.n8 minus.t0 109.355
R9 minus.n10 minus.t5 109.355
R10 minus.n1 minus.n0 44.8973
R11 minus.n7 minus.n6 44.8973
R12 minus.n4 minus.n3 33.5944
R13 minus.n10 minus.n9 33.5944
R14 minus.n12 minus.n5 27.9039
R15 minus.n2 minus.n1 18.1882
R16 minus.n8 minus.n7 18.1882
R17 minus.n3 minus.n2 14.6066
R18 minus.n9 minus.n8 14.6066
R19 minus.n12 minus.n11 6.72209
R20 minus.n5 minus.n0 0.189894
R21 minus.n11 minus.n6 0.189894
R22 minus minus.n12 0.188
R23 drain_right.n2 drain_right.n0 289.615
R24 drain_right.n12 drain_right.n10 289.615
R25 drain_right.n3 drain_right.n2 185
R26 drain_right.n13 drain_right.n12 185
R27 drain_right.t1 drain_right.n1 167.117
R28 drain_right.t4 drain_right.n11 167.117
R29 drain_right.n17 drain_right.n9 101.769
R30 drain_right.n8 drain_right.n7 100.984
R31 drain_right.n2 drain_right.t1 52.3082
R32 drain_right.n12 drain_right.t4 52.3082
R33 drain_right.n8 drain_right.n6 48.7636
R34 drain_right.n17 drain_right.n16 48.0884
R35 drain_right drain_right.n8 21.917
R36 drain_right.n7 drain_right.t0 9.9005
R37 drain_right.n7 drain_right.t5 9.9005
R38 drain_right.n9 drain_right.t3 9.9005
R39 drain_right.n9 drain_right.t2 9.9005
R40 drain_right.n3 drain_right.n1 9.71174
R41 drain_right.n13 drain_right.n11 9.71174
R42 drain_right.n6 drain_right.n5 9.45567
R43 drain_right.n16 drain_right.n15 9.45567
R44 drain_right.n5 drain_right.n4 9.3005
R45 drain_right.n15 drain_right.n14 9.3005
R46 drain_right.n6 drain_right.n0 8.14595
R47 drain_right.n16 drain_right.n10 8.14595
R48 drain_right.n4 drain_right.n3 7.3702
R49 drain_right.n14 drain_right.n13 7.3702
R50 drain_right drain_right.n17 6.14028
R51 drain_right.n4 drain_right.n0 5.81868
R52 drain_right.n14 drain_right.n10 5.81868
R53 drain_right.n5 drain_right.n1 3.44771
R54 drain_right.n15 drain_right.n11 3.44771
R55 source.n34 source.n32 289.615
R56 source.n24 source.n22 289.615
R57 source.n2 source.n0 289.615
R58 source.n12 source.n10 289.615
R59 source.n35 source.n34 185
R60 source.n25 source.n24 185
R61 source.n3 source.n2 185
R62 source.n13 source.n12 185
R63 source.t6 source.n33 167.117
R64 source.t3 source.n23 167.117
R65 source.t2 source.n1 167.117
R66 source.t8 source.n11 167.117
R67 source.n9 source.n8 84.1169
R68 source.n19 source.n18 84.1169
R69 source.n31 source.n30 84.1168
R70 source.n21 source.n20 84.1168
R71 source.n34 source.t6 52.3082
R72 source.n24 source.t3 52.3082
R73 source.n2 source.t2 52.3082
R74 source.n12 source.t8 52.3082
R75 source.n39 source.n38 31.4096
R76 source.n29 source.n28 31.4096
R77 source.n7 source.n6 31.4096
R78 source.n17 source.n16 31.4096
R79 source.n21 source.n19 15.6602
R80 source.n30 source.t7 9.9005
R81 source.n30 source.t11 9.9005
R82 source.n20 source.t4 9.9005
R83 source.n20 source.t0 9.9005
R84 source.n8 source.t1 9.9005
R85 source.n8 source.t5 9.9005
R86 source.n18 source.t10 9.9005
R87 source.n18 source.t9 9.9005
R88 source.n35 source.n33 9.71174
R89 source.n25 source.n23 9.71174
R90 source.n3 source.n1 9.71174
R91 source.n13 source.n11 9.71174
R92 source.n38 source.n37 9.45567
R93 source.n28 source.n27 9.45567
R94 source.n6 source.n5 9.45567
R95 source.n16 source.n15 9.45567
R96 source.n37 source.n36 9.3005
R97 source.n27 source.n26 9.3005
R98 source.n5 source.n4 9.3005
R99 source.n15 source.n14 9.3005
R100 source.n40 source.n7 8.93611
R101 source.n38 source.n32 8.14595
R102 source.n28 source.n22 8.14595
R103 source.n6 source.n0 8.14595
R104 source.n16 source.n10 8.14595
R105 source.n36 source.n35 7.3702
R106 source.n26 source.n25 7.3702
R107 source.n4 source.n3 7.3702
R108 source.n14 source.n13 7.3702
R109 source.n36 source.n32 5.81868
R110 source.n26 source.n22 5.81868
R111 source.n4 source.n0 5.81868
R112 source.n14 source.n10 5.81868
R113 source.n40 source.n39 5.7505
R114 source.n37 source.n33 3.44771
R115 source.n27 source.n23 3.44771
R116 source.n5 source.n1 3.44771
R117 source.n15 source.n11 3.44771
R118 source.n19 source.n17 0.974638
R119 source.n9 source.n7 0.974638
R120 source.n29 source.n21 0.974638
R121 source.n39 source.n31 0.974638
R122 source.n17 source.n9 0.957397
R123 source.n31 source.n29 0.957397
R124 source source.n40 0.188
R125 plus.n3 plus.n0 161.3
R126 plus.n5 plus.n4 161.3
R127 plus.n9 plus.n6 161.3
R128 plus.n11 plus.n10 161.3
R129 plus.n7 plus.t3 132.84
R130 plus.n1 plus.t4 132.84
R131 plus.n4 plus.t1 109.355
R132 plus.n2 plus.t2 109.355
R133 plus.n10 plus.t5 109.355
R134 plus.n8 plus.t0 109.355
R135 plus.n7 plus.n6 44.8973
R136 plus.n1 plus.n0 44.8973
R137 plus.n4 plus.n3 33.5944
R138 plus.n10 plus.n9 33.5944
R139 plus plus.n11 25.5729
R140 plus.n8 plus.n7 18.1882
R141 plus.n2 plus.n1 18.1882
R142 plus.n3 plus.n2 14.6066
R143 plus.n9 plus.n8 14.6066
R144 plus plus.n5 8.57815
R145 plus.n5 plus.n0 0.189894
R146 plus.n11 plus.n6 0.189894
R147 drain_left.n2 drain_left.n0 289.615
R148 drain_left.n11 drain_left.n9 289.615
R149 drain_left.n3 drain_left.n2 185
R150 drain_left.n12 drain_left.n11 185
R151 drain_left.t0 drain_left.n1 167.117
R152 drain_left.t1 drain_left.n10 167.117
R153 drain_left.n8 drain_left.n7 100.984
R154 drain_left.n17 drain_left.n16 100.796
R155 drain_left.n2 drain_left.t0 52.3082
R156 drain_left.n11 drain_left.t1 52.3082
R157 drain_left.n17 drain_left.n15 49.0625
R158 drain_left.n8 drain_left.n6 48.7636
R159 drain_left drain_left.n8 22.4702
R160 drain_left.n7 drain_left.t5 9.9005
R161 drain_left.n7 drain_left.t2 9.9005
R162 drain_left.n16 drain_left.t3 9.9005
R163 drain_left.n16 drain_left.t4 9.9005
R164 drain_left.n3 drain_left.n1 9.71174
R165 drain_left.n12 drain_left.n10 9.71174
R166 drain_left.n6 drain_left.n5 9.45567
R167 drain_left.n15 drain_left.n14 9.45567
R168 drain_left.n5 drain_left.n4 9.3005
R169 drain_left.n14 drain_left.n13 9.3005
R170 drain_left.n6 drain_left.n0 8.14595
R171 drain_left.n15 drain_left.n9 8.14595
R172 drain_left.n4 drain_left.n3 7.3702
R173 drain_left.n13 drain_left.n12 7.3702
R174 drain_left drain_left.n17 6.62735
R175 drain_left.n4 drain_left.n0 5.81868
R176 drain_left.n13 drain_left.n9 5.81868
R177 drain_left.n5 drain_left.n1 3.44771
R178 drain_left.n14 drain_left.n10 3.44771
C0 source drain_left 3.26904f
C1 plus minus 3.30956f
C2 source drain_right 3.26912f
C3 drain_left drain_right 0.74246f
C4 source plus 1.3115f
C5 drain_left plus 1.21679f
C6 source minus 1.29746f
C7 drain_left minus 0.177716f
C8 drain_right plus 0.317445f
C9 drain_right minus 1.06149f
C10 drain_right a_n1620_n1288# 3.297284f
C11 drain_left a_n1620_n1288# 3.508325f
C12 source a_n1620_n1288# 2.52452f
C13 minus a_n1620_n1288# 5.362693f
C14 plus a_n1620_n1288# 5.94926f
C15 drain_left.n0 a_n1620_n1288# 0.025077f
C16 drain_left.n1 a_n1620_n1288# 0.055486f
C17 drain_left.t0 a_n1620_n1288# 0.041639f
C18 drain_left.n2 a_n1620_n1288# 0.043425f
C19 drain_left.n3 a_n1620_n1288# 0.013999f
C20 drain_left.n4 a_n1620_n1288# 0.009232f
C21 drain_left.n5 a_n1620_n1288# 0.122304f
C22 drain_left.n6 a_n1620_n1288# 0.040338f
C23 drain_left.t5 a_n1620_n1288# 0.027154f
C24 drain_left.t2 a_n1620_n1288# 0.027154f
C25 drain_left.n7 a_n1620_n1288# 0.170972f
C26 drain_left.n8 a_n1620_n1288# 0.745393f
C27 drain_left.n9 a_n1620_n1288# 0.025077f
C28 drain_left.n10 a_n1620_n1288# 0.055486f
C29 drain_left.t1 a_n1620_n1288# 0.041639f
C30 drain_left.n11 a_n1620_n1288# 0.043425f
C31 drain_left.n12 a_n1620_n1288# 0.013999f
C32 drain_left.n13 a_n1620_n1288# 0.009232f
C33 drain_left.n14 a_n1620_n1288# 0.122304f
C34 drain_left.n15 a_n1620_n1288# 0.041078f
C35 drain_left.t3 a_n1620_n1288# 0.027154f
C36 drain_left.t4 a_n1620_n1288# 0.027154f
C37 drain_left.n16 a_n1620_n1288# 0.170591f
C38 drain_left.n17 a_n1620_n1288# 0.478182f
C39 plus.n0 a_n1620_n1288# 0.122263f
C40 plus.t1 a_n1620_n1288# 0.140113f
C41 plus.t2 a_n1620_n1288# 0.140113f
C42 plus.t4 a_n1620_n1288# 0.157182f
C43 plus.n1 a_n1620_n1288# 0.082024f
C44 plus.n2 a_n1620_n1288# 0.098085f
C45 plus.n3 a_n1620_n1288# 0.006417f
C46 plus.n4 a_n1620_n1288# 0.095335f
C47 plus.n5 a_n1620_n1288# 0.217612f
C48 plus.n6 a_n1620_n1288# 0.122263f
C49 plus.t5 a_n1620_n1288# 0.140113f
C50 plus.t3 a_n1620_n1288# 0.157182f
C51 plus.n7 a_n1620_n1288# 0.082024f
C52 plus.t0 a_n1620_n1288# 0.140113f
C53 plus.n8 a_n1620_n1288# 0.098085f
C54 plus.n9 a_n1620_n1288# 0.006417f
C55 plus.n10 a_n1620_n1288# 0.095335f
C56 plus.n11 a_n1620_n1288# 0.627014f
C57 source.n0 a_n1620_n1288# 0.032246f
C58 source.n1 a_n1620_n1288# 0.071348f
C59 source.t2 a_n1620_n1288# 0.053543f
C60 source.n2 a_n1620_n1288# 0.05584f
C61 source.n3 a_n1620_n1288# 0.018001f
C62 source.n4 a_n1620_n1288# 0.011872f
C63 source.n5 a_n1620_n1288# 0.157268f
C64 source.n6 a_n1620_n1288# 0.035349f
C65 source.n7 a_n1620_n1288# 0.387891f
C66 source.t1 a_n1620_n1288# 0.034917f
C67 source.t5 a_n1620_n1288# 0.034917f
C68 source.n8 a_n1620_n1288# 0.186665f
C69 source.n9 a_n1620_n1288# 0.309228f
C70 source.n10 a_n1620_n1288# 0.032246f
C71 source.n11 a_n1620_n1288# 0.071348f
C72 source.t8 a_n1620_n1288# 0.053543f
C73 source.n12 a_n1620_n1288# 0.05584f
C74 source.n13 a_n1620_n1288# 0.018001f
C75 source.n14 a_n1620_n1288# 0.011872f
C76 source.n15 a_n1620_n1288# 0.157268f
C77 source.n16 a_n1620_n1288# 0.035349f
C78 source.n17 a_n1620_n1288# 0.155654f
C79 source.t10 a_n1620_n1288# 0.034917f
C80 source.t9 a_n1620_n1288# 0.034917f
C81 source.n18 a_n1620_n1288# 0.186665f
C82 source.n19 a_n1620_n1288# 0.823828f
C83 source.t4 a_n1620_n1288# 0.034917f
C84 source.t0 a_n1620_n1288# 0.034917f
C85 source.n20 a_n1620_n1288# 0.186664f
C86 source.n21 a_n1620_n1288# 0.82383f
C87 source.n22 a_n1620_n1288# 0.032246f
C88 source.n23 a_n1620_n1288# 0.071348f
C89 source.t3 a_n1620_n1288# 0.053543f
C90 source.n24 a_n1620_n1288# 0.05584f
C91 source.n25 a_n1620_n1288# 0.018001f
C92 source.n26 a_n1620_n1288# 0.011872f
C93 source.n27 a_n1620_n1288# 0.157268f
C94 source.n28 a_n1620_n1288# 0.035349f
C95 source.n29 a_n1620_n1288# 0.155654f
C96 source.t7 a_n1620_n1288# 0.034917f
C97 source.t11 a_n1620_n1288# 0.034917f
C98 source.n30 a_n1620_n1288# 0.186664f
C99 source.n31 a_n1620_n1288# 0.30923f
C100 source.n32 a_n1620_n1288# 0.032246f
C101 source.n33 a_n1620_n1288# 0.071348f
C102 source.t6 a_n1620_n1288# 0.053543f
C103 source.n34 a_n1620_n1288# 0.05584f
C104 source.n35 a_n1620_n1288# 0.018001f
C105 source.n36 a_n1620_n1288# 0.011872f
C106 source.n37 a_n1620_n1288# 0.157268f
C107 source.n38 a_n1620_n1288# 0.035349f
C108 source.n39 a_n1620_n1288# 0.269876f
C109 source.n40 a_n1620_n1288# 0.559762f
C110 drain_right.n0 a_n1620_n1288# 0.025598f
C111 drain_right.n1 a_n1620_n1288# 0.056639f
C112 drain_right.t1 a_n1620_n1288# 0.042505f
C113 drain_right.n2 a_n1620_n1288# 0.044328f
C114 drain_right.n3 a_n1620_n1288# 0.01429f
C115 drain_right.n4 a_n1620_n1288# 0.009424f
C116 drain_right.n5 a_n1620_n1288# 0.124847f
C117 drain_right.n6 a_n1620_n1288# 0.041176f
C118 drain_right.t0 a_n1620_n1288# 0.027719f
C119 drain_right.t5 a_n1620_n1288# 0.027719f
C120 drain_right.n7 a_n1620_n1288# 0.174527f
C121 drain_right.n8 a_n1620_n1288# 0.726442f
C122 drain_right.t3 a_n1620_n1288# 0.027719f
C123 drain_right.t2 a_n1620_n1288# 0.027719f
C124 drain_right.n9 a_n1620_n1288# 0.176544f
C125 drain_right.n10 a_n1620_n1288# 0.025598f
C126 drain_right.n11 a_n1620_n1288# 0.056639f
C127 drain_right.t4 a_n1620_n1288# 0.042505f
C128 drain_right.n12 a_n1620_n1288# 0.044328f
C129 drain_right.n13 a_n1620_n1288# 0.01429f
C130 drain_right.n14 a_n1620_n1288# 0.009424f
C131 drain_right.n15 a_n1620_n1288# 0.124847f
C132 drain_right.n16 a_n1620_n1288# 0.040179f
C133 drain_right.n17 a_n1620_n1288# 0.502129f
C134 minus.n0 a_n1620_n1288# 0.120181f
C135 minus.t3 a_n1620_n1288# 0.154505f
C136 minus.n1 a_n1620_n1288# 0.080626f
C137 minus.t2 a_n1620_n1288# 0.137726f
C138 minus.n2 a_n1620_n1288# 0.096414f
C139 minus.n3 a_n1620_n1288# 0.006308f
C140 minus.t1 a_n1620_n1288# 0.137726f
C141 minus.n4 a_n1620_n1288# 0.093711f
C142 minus.n5 a_n1620_n1288# 0.643659f
C143 minus.n6 a_n1620_n1288# 0.120181f
C144 minus.t4 a_n1620_n1288# 0.154505f
C145 minus.n7 a_n1620_n1288# 0.080626f
C146 minus.t0 a_n1620_n1288# 0.137726f
C147 minus.n8 a_n1620_n1288# 0.096414f
C148 minus.n9 a_n1620_n1288# 0.006308f
C149 minus.t5 a_n1620_n1288# 0.137726f
C150 minus.n10 a_n1620_n1288# 0.093711f
C151 minus.n11 a_n1620_n1288# 0.196123f
C152 minus.n12 a_n1620_n1288# 0.78757f
.ends

