* NGSPICE file created from diffpair242.ext - technology: sky130A

.subckt diffpair242 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t10 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X1 a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X2 source.t4 minus.t0 drain_right.t5 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X3 a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X4 source.t6 plus.t1 drain_left.t4 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X5 drain_right.t4 minus.t1 source.t5 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X6 source.t0 minus.t2 drain_right.t3 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X8 drain_right.t2 minus.t3 source.t1 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X9 drain_left.t3 plus.t2 source.t11 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X10 drain_right.t1 minus.t4 source.t3 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X11 drain_right.t0 minus.t5 source.t2 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X12 drain_left.t2 plus.t3 source.t7 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X13 drain_left.t1 plus.t4 source.t9 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X14 source.t8 plus.t5 drain_left.t0 a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# a_n1236_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
R0 plus.n0 plus.t2 1231.29
R1 plus.n2 plus.t3 1231.29
R2 plus.n4 plus.t0 1231.29
R3 plus.n6 plus.t4 1231.29
R4 plus.n1 plus.t5 1172.87
R5 plus.n5 plus.t1 1172.87
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 25.463
R15 plus plus.n3 9.92285
R16 source.n3 source.t1 55.512
R17 source.n0 source.t7 55.5119
R18 source.n11 source.t5 55.5119
R19 source.n8 source.t10 55.5119
R20 source.n2 source.n1 50.512
R21 source.n5 source.n4 50.512
R22 source.n10 source.n9 50.5119
R23 source.n7 source.n6 50.5119
R24 source.n7 source.n5 17.863
R25 source.n12 source.n0 11.7595
R26 source.n12 source.n11 5.5436
R27 source.n9 source.t2 5.0005
R28 source.n9 source.t4 5.0005
R29 source.n6 source.t9 5.0005
R30 source.n6 source.t6 5.0005
R31 source.n1 source.t11 5.0005
R32 source.n1 source.t8 5.0005
R33 source.n4 source.t3 5.0005
R34 source.n4 source.t0 5.0005
R35 source.n3 source.n2 0.7505
R36 source.n10 source.n8 0.7505
R37 source.n5 source.n3 0.560845
R38 source.n2 source.n0 0.560845
R39 source.n8 source.n7 0.560845
R40 source.n11 source.n10 0.560845
R41 source source.n12 0.188
R42 drain_left.n3 drain_left.t3 72.7512
R43 drain_left.n1 drain_left.t1 72.5556
R44 drain_left.n1 drain_left.n0 67.2754
R45 drain_left.n3 drain_left.n2 67.1907
R46 drain_left drain_left.n1 24.3626
R47 drain_left drain_left.n3 6.21356
R48 drain_left.n0 drain_left.t4 5.0005
R49 drain_left.n0 drain_left.t5 5.0005
R50 drain_left.n2 drain_left.t0 5.0005
R51 drain_left.n2 drain_left.t2 5.0005
R52 minus.n2 minus.t4 1231.29
R53 minus.n0 minus.t3 1231.29
R54 minus.n6 minus.t1 1231.29
R55 minus.n4 minus.t5 1231.29
R56 minus.n1 minus.t2 1172.87
R57 minus.n5 minus.t0 1172.87
R58 minus.n3 minus.n0 161.489
R59 minus.n7 minus.n4 161.489
R60 minus.n3 minus.n2 161.3
R61 minus.n7 minus.n6 161.3
R62 minus.n2 minus.n1 36.5157
R63 minus.n1 minus.n0 36.5157
R64 minus.n5 minus.n4 36.5157
R65 minus.n6 minus.n5 36.5157
R66 minus.n8 minus.n3 29.3092
R67 minus.n8 minus.n7 6.55164
R68 minus minus.n8 0.188
R69 drain_right.n1 drain_right.t0 72.5556
R70 drain_right.n3 drain_right.t1 72.1908
R71 drain_right.n3 drain_right.n2 67.751
R72 drain_right.n1 drain_right.n0 67.2754
R73 drain_right drain_right.n1 23.8093
R74 drain_right drain_right.n3 5.93339
R75 drain_right.n0 drain_right.t5 5.0005
R76 drain_right.n0 drain_right.t4 5.0005
R77 drain_right.n2 drain_right.t3 5.0005
R78 drain_right.n2 drain_right.t2 5.0005
C0 minus plus 3.56375f
C1 source drain_right 8.00688f
C2 minus drain_right 1.07202f
C3 minus source 0.836291f
C4 drain_left plus 1.18648f
C5 drain_left drain_right 0.573457f
C6 drain_left source 8.01349f
C7 drain_right plus 0.27008f
C8 minus drain_left 0.170478f
C9 source plus 0.850631f
C10 drain_right a_n1236_n2088# 4.18814f
C11 drain_left a_n1236_n2088# 4.34982f
C12 source a_n1236_n2088# 3.851546f
C13 minus a_n1236_n2088# 4.044858f
C14 plus a_n1236_n2088# 5.09511f
C15 drain_right.t0 a_n1236_n2088# 1.14702f
C16 drain_right.t5 a_n1236_n2088# 0.152735f
C17 drain_right.t4 a_n1236_n2088# 0.152735f
C18 drain_right.n0 a_n1236_n2088# 0.944863f
C19 drain_right.n1 a_n1236_n2088# 1.09763f
C20 drain_right.t3 a_n1236_n2088# 0.152735f
C21 drain_right.t2 a_n1236_n2088# 0.152735f
C22 drain_right.n2 a_n1236_n2088# 0.946705f
C23 drain_right.t1 a_n1236_n2088# 1.14561f
C24 drain_right.n3 a_n1236_n2088# 0.727431f
C25 minus.t3 a_n1236_n2088# 0.104035f
C26 minus.n0 a_n1236_n2088# 0.068189f
C27 minus.t4 a_n1236_n2088# 0.104035f
C28 minus.t2 a_n1236_n2088# 0.101478f
C29 minus.n1 a_n1236_n2088# 0.05268f
C30 minus.n2 a_n1236_n2088# 0.06813f
C31 minus.n3 a_n1236_n2088# 1.04154f
C32 minus.t5 a_n1236_n2088# 0.104035f
C33 minus.n4 a_n1236_n2088# 0.068189f
C34 minus.t0 a_n1236_n2088# 0.101478f
C35 minus.n5 a_n1236_n2088# 0.05268f
C36 minus.t1 a_n1236_n2088# 0.104035f
C37 minus.n6 a_n1236_n2088# 0.06813f
C38 minus.n7 a_n1236_n2088# 0.314021f
C39 minus.n8 a_n1236_n2088# 1.22135f
C40 drain_left.t1 a_n1236_n2088# 1.13522f
C41 drain_left.t4 a_n1236_n2088# 0.151163f
C42 drain_left.t5 a_n1236_n2088# 0.151163f
C43 drain_left.n0 a_n1236_n2088# 0.935141f
C44 drain_left.n1 a_n1236_n2088# 1.12951f
C45 drain_left.t3 a_n1236_n2088# 1.13606f
C46 drain_left.t0 a_n1236_n2088# 0.151163f
C47 drain_left.t2 a_n1236_n2088# 0.151163f
C48 drain_left.n2 a_n1236_n2088# 0.934853f
C49 drain_left.n3 a_n1236_n2088# 0.710626f
C50 source.t7 a_n1236_n2088# 1.17519f
C51 source.n0 a_n1236_n2088# 0.864557f
C52 source.t11 a_n1236_n2088# 0.167315f
C53 source.t8 a_n1236_n2088# 0.167315f
C54 source.n1 a_n1236_n2088# 0.973793f
C55 source.n2 a_n1236_n2088# 0.316659f
C56 source.t1 a_n1236_n2088# 1.17519f
C57 source.n3 a_n1236_n2088# 0.416426f
C58 source.t3 a_n1236_n2088# 0.167315f
C59 source.t0 a_n1236_n2088# 0.167315f
C60 source.n4 a_n1236_n2088# 0.973793f
C61 source.n5 a_n1236_n2088# 1.10704f
C62 source.t9 a_n1236_n2088# 0.167315f
C63 source.t6 a_n1236_n2088# 0.167315f
C64 source.n6 a_n1236_n2088# 0.973787f
C65 source.n7 a_n1236_n2088# 1.10705f
C66 source.t10 a_n1236_n2088# 1.17519f
C67 source.n8 a_n1236_n2088# 0.416432f
C68 source.t2 a_n1236_n2088# 0.167315f
C69 source.t4 a_n1236_n2088# 0.167315f
C70 source.n9 a_n1236_n2088# 0.973787f
C71 source.n10 a_n1236_n2088# 0.316665f
C72 source.t5 a_n1236_n2088# 1.17519f
C73 source.n11 a_n1236_n2088# 0.527913f
C74 source.n12 a_n1236_n2088# 0.953623f
C75 plus.t2 a_n1236_n2088# 0.106401f
C76 plus.n0 a_n1236_n2088# 0.06974f
C77 plus.t5 a_n1236_n2088# 0.103785f
C78 plus.n1 a_n1236_n2088# 0.053877f
C79 plus.t3 a_n1236_n2088# 0.106401f
C80 plus.n2 a_n1236_n2088# 0.069679f
C81 plus.n3 a_n1236_n2088# 0.403586f
C82 plus.t0 a_n1236_n2088# 0.106401f
C83 plus.n4 a_n1236_n2088# 0.06974f
C84 plus.t4 a_n1236_n2088# 0.106401f
C85 plus.t1 a_n1236_n2088# 0.103785f
C86 plus.n5 a_n1236_n2088# 0.053877f
C87 plus.n6 a_n1236_n2088# 0.069679f
C88 plus.n7 a_n1236_n2088# 0.969234f
.ends

