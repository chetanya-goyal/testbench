* NGSPICE file created from diffpair239.ext - technology: sky130A

.subckt diffpair239 minus drain_right drain_left source plus
X0 source.t41 minus.t0 drain_right.t0 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X1 a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X2 source.t40 minus.t1 drain_right.t1 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X3 drain_left.t23 plus.t0 source.t3 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X4 drain_left.t22 plus.t1 source.t45 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X5 drain_left.t21 plus.t2 source.t47 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X6 source.t39 minus.t2 drain_right.t2 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X7 source.t38 minus.t3 drain_right.t3 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X8 source.t37 minus.t4 drain_right.t4 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X9 drain_left.t20 plus.t3 source.t6 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X10 drain_left.t19 plus.t4 source.t42 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X11 drain_left.t18 plus.t5 source.t0 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X12 source.t36 minus.t5 drain_right.t5 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X13 source.t35 minus.t6 drain_right.t6 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X14 drain_left.t17 plus.t6 source.t12 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X15 source.t1 plus.t7 drain_left.t16 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X16 source.t9 plus.t8 drain_left.t15 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X17 drain_right.t7 minus.t7 source.t34 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X18 drain_right.t8 minus.t8 source.t33 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 drain_left.t14 plus.t9 source.t4 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X20 source.t32 minus.t9 drain_right.t12 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X21 source.t31 minus.t10 drain_right.t13 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X22 drain_right.t9 minus.t11 source.t30 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X23 drain_right.t14 minus.t12 source.t29 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X24 drain_right.t10 minus.t13 source.t28 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X25 source.t14 plus.t10 drain_left.t13 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X26 drain_right.t11 minus.t14 source.t27 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X27 source.t10 plus.t11 drain_left.t12 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X28 source.t26 minus.t15 drain_right.t15 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X29 drain_right.t16 minus.t16 source.t25 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X30 drain_right.t17 minus.t17 source.t24 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X31 source.t8 plus.t12 drain_left.t11 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X32 drain_left.t10 plus.t13 source.t11 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X33 source.t23 minus.t18 drain_right.t18 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X34 drain_right.t19 minus.t19 source.t22 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X35 source.t7 plus.t14 drain_left.t9 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X36 source.t17 plus.t15 drain_left.t8 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X37 drain_right.t20 minus.t20 source.t21 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X38 source.t13 plus.t16 drain_left.t7 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X39 a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X40 drain_left.t6 plus.t17 source.t15 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X41 drain_left.t5 plus.t18 source.t44 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X42 source.t20 minus.t21 drain_right.t21 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X43 drain_right.t22 minus.t22 source.t19 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X44 source.t46 plus.t19 drain_left.t4 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X45 drain_right.t23 minus.t23 source.t18 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X46 source.t5 plus.t20 drain_left.t3 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X47 source.t2 plus.t21 drain_left.t2 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X48 drain_left.t1 plus.t22 source.t43 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X49 a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X50 source.t16 plus.t23 drain_left.t0 a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X51 a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# a_n3654_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
R0 minus.n35 minus.n34 161.3
R1 minus.n33 minus.n0 161.3
R2 minus.n29 minus.n28 161.3
R3 minus.n27 minus.n2 161.3
R4 minus.n26 minus.n25 161.3
R5 minus.n24 minus.n3 161.3
R6 minus.n23 minus.n22 161.3
R7 minus.n18 minus.n5 161.3
R8 minus.n17 minus.n16 161.3
R9 minus.n15 minus.n6 161.3
R10 minus.n14 minus.n13 161.3
R11 minus.n12 minus.n7 161.3
R12 minus.n71 minus.n70 161.3
R13 minus.n69 minus.n36 161.3
R14 minus.n65 minus.n64 161.3
R15 minus.n63 minus.n38 161.3
R16 minus.n62 minus.n61 161.3
R17 minus.n60 minus.n39 161.3
R18 minus.n59 minus.n58 161.3
R19 minus.n54 minus.n41 161.3
R20 minus.n53 minus.n52 161.3
R21 minus.n51 minus.n42 161.3
R22 minus.n50 minus.n49 161.3
R23 minus.n48 minus.n43 161.3
R24 minus.n8 minus.t14 160.916
R25 minus.n44 minus.t3 160.916
R26 minus.n9 minus.t9 139.48
R27 minus.n10 minus.t7 139.48
R28 minus.n14 minus.t18 139.48
R29 minus.n16 minus.t20 139.48
R30 minus.n20 minus.t15 139.48
R31 minus.n21 minus.t12 139.48
R32 minus.n3 minus.t21 139.48
R33 minus.n27 minus.t19 139.48
R34 minus.n1 minus.t5 139.48
R35 minus.n32 minus.t13 139.48
R36 minus.n34 minus.t10 139.48
R37 minus.n45 minus.t8 139.48
R38 minus.n46 minus.t4 139.48
R39 minus.n50 minus.t11 139.48
R40 minus.n52 minus.t0 139.48
R41 minus.n56 minus.t17 139.48
R42 minus.n57 minus.t1 139.48
R43 minus.n39 minus.t16 139.48
R44 minus.n63 minus.t2 139.48
R45 minus.n37 minus.t22 139.48
R46 minus.n68 minus.t6 139.48
R47 minus.n70 minus.t23 139.48
R48 minus.n32 minus.n31 80.6037
R49 minus.n30 minus.n1 80.6037
R50 minus.n21 minus.n4 80.6037
R51 minus.n20 minus.n19 80.6037
R52 minus.n11 minus.n10 80.6037
R53 minus.n68 minus.n67 80.6037
R54 minus.n66 minus.n37 80.6037
R55 minus.n57 minus.n40 80.6037
R56 minus.n56 minus.n55 80.6037
R57 minus.n47 minus.n46 80.6037
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n20 minus.n5 41.6278
R69 minus.n22 minus.n21 41.6278
R70 minus.n56 minus.n41 41.6278
R71 minus.n58 minus.n57 41.6278
R72 minus.n33 minus.n32 38.7066
R73 minus.n69 minus.n68 38.7066
R74 minus.n72 minus.n35 36.3035
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 drain_right.n13 drain_right.n11 80.7472
R132 drain_right.n7 drain_right.n5 80.7471
R133 drain_right.n2 drain_right.n0 80.7471
R134 drain_right.n13 drain_right.n12 79.7731
R135 drain_right.n15 drain_right.n14 79.7731
R136 drain_right.n17 drain_right.n16 79.7731
R137 drain_right.n19 drain_right.n18 79.7731
R138 drain_right.n21 drain_right.n20 79.7731
R139 drain_right.n7 drain_right.n6 79.773
R140 drain_right.n9 drain_right.n8 79.773
R141 drain_right.n4 drain_right.n3 79.773
R142 drain_right.n2 drain_right.n1 79.773
R143 drain_right drain_right.n10 29.25
R144 drain_right drain_right.n21 6.62735
R145 drain_right.n5 drain_right.t6 6.6005
R146 drain_right.n5 drain_right.t23 6.6005
R147 drain_right.n6 drain_right.t2 6.6005
R148 drain_right.n6 drain_right.t22 6.6005
R149 drain_right.n8 drain_right.t1 6.6005
R150 drain_right.n8 drain_right.t16 6.6005
R151 drain_right.n3 drain_right.t0 6.6005
R152 drain_right.n3 drain_right.t17 6.6005
R153 drain_right.n1 drain_right.t4 6.6005
R154 drain_right.n1 drain_right.t9 6.6005
R155 drain_right.n0 drain_right.t3 6.6005
R156 drain_right.n0 drain_right.t8 6.6005
R157 drain_right.n11 drain_right.t12 6.6005
R158 drain_right.n11 drain_right.t11 6.6005
R159 drain_right.n12 drain_right.t18 6.6005
R160 drain_right.n12 drain_right.t7 6.6005
R161 drain_right.n14 drain_right.t15 6.6005
R162 drain_right.n14 drain_right.t20 6.6005
R163 drain_right.n16 drain_right.t21 6.6005
R164 drain_right.n16 drain_right.t14 6.6005
R165 drain_right.n18 drain_right.t5 6.6005
R166 drain_right.n18 drain_right.t19 6.6005
R167 drain_right.n20 drain_right.t13 6.6005
R168 drain_right.n20 drain_right.t10 6.6005
R169 drain_right.n9 drain_right.n7 0.974638
R170 drain_right.n4 drain_right.n2 0.974638
R171 drain_right.n21 drain_right.n19 0.974638
R172 drain_right.n19 drain_right.n17 0.974638
R173 drain_right.n17 drain_right.n15 0.974638
R174 drain_right.n15 drain_right.n13 0.974638
R175 drain_right.n10 drain_right.n9 0.432223
R176 drain_right.n10 drain_right.n4 0.432223
R177 source.n0 source.t12 69.6943
R178 source.n11 source.t16 69.6943
R179 source.n12 source.t27 69.6943
R180 source.n23 source.t31 69.6943
R181 source.n47 source.t18 69.6942
R182 source.n36 source.t38 69.6942
R183 source.n35 source.t42 69.6942
R184 source.n24 source.t14 69.6942
R185 source.n2 source.n1 63.0943
R186 source.n4 source.n3 63.0943
R187 source.n6 source.n5 63.0943
R188 source.n8 source.n7 63.0943
R189 source.n10 source.n9 63.0943
R190 source.n14 source.n13 63.0943
R191 source.n16 source.n15 63.0943
R192 source.n18 source.n17 63.0943
R193 source.n20 source.n19 63.0943
R194 source.n22 source.n21 63.0943
R195 source.n46 source.n45 63.0942
R196 source.n44 source.n43 63.0942
R197 source.n42 source.n41 63.0942
R198 source.n40 source.n39 63.0942
R199 source.n38 source.n37 63.0942
R200 source.n34 source.n33 63.0942
R201 source.n32 source.n31 63.0942
R202 source.n30 source.n29 63.0942
R203 source.n28 source.n27 63.0942
R204 source.n26 source.n25 63.0942
R205 source.n24 source.n23 15.4437
R206 source.n48 source.n0 9.69368
R207 source.n45 source.t19 6.6005
R208 source.n45 source.t35 6.6005
R209 source.n43 source.t25 6.6005
R210 source.n43 source.t39 6.6005
R211 source.n41 source.t24 6.6005
R212 source.n41 source.t40 6.6005
R213 source.n39 source.t30 6.6005
R214 source.n39 source.t41 6.6005
R215 source.n37 source.t33 6.6005
R216 source.n37 source.t37 6.6005
R217 source.n33 source.t0 6.6005
R218 source.n33 source.t8 6.6005
R219 source.n31 source.t3 6.6005
R220 source.n31 source.t7 6.6005
R221 source.n29 source.t45 6.6005
R222 source.n29 source.t17 6.6005
R223 source.n27 source.t47 6.6005
R224 source.n27 source.t1 6.6005
R225 source.n25 source.t6 6.6005
R226 source.n25 source.t5 6.6005
R227 source.n1 source.t4 6.6005
R228 source.n1 source.t9 6.6005
R229 source.n3 source.t11 6.6005
R230 source.n3 source.t10 6.6005
R231 source.n5 source.t15 6.6005
R232 source.n5 source.t13 6.6005
R233 source.n7 source.t44 6.6005
R234 source.n7 source.t2 6.6005
R235 source.n9 source.t43 6.6005
R236 source.n9 source.t46 6.6005
R237 source.n13 source.t34 6.6005
R238 source.n13 source.t32 6.6005
R239 source.n15 source.t21 6.6005
R240 source.n15 source.t23 6.6005
R241 source.n17 source.t29 6.6005
R242 source.n17 source.t26 6.6005
R243 source.n19 source.t22 6.6005
R244 source.n19 source.t20 6.6005
R245 source.n21 source.t28 6.6005
R246 source.n21 source.t36 6.6005
R247 source.n48 source.n47 5.7505
R248 source.n23 source.n22 0.974638
R249 source.n22 source.n20 0.974638
R250 source.n20 source.n18 0.974638
R251 source.n18 source.n16 0.974638
R252 source.n16 source.n14 0.974638
R253 source.n14 source.n12 0.974638
R254 source.n11 source.n10 0.974638
R255 source.n10 source.n8 0.974638
R256 source.n8 source.n6 0.974638
R257 source.n6 source.n4 0.974638
R258 source.n4 source.n2 0.974638
R259 source.n2 source.n0 0.974638
R260 source.n26 source.n24 0.974638
R261 source.n28 source.n26 0.974638
R262 source.n30 source.n28 0.974638
R263 source.n32 source.n30 0.974638
R264 source.n34 source.n32 0.974638
R265 source.n35 source.n34 0.974638
R266 source.n38 source.n36 0.974638
R267 source.n40 source.n38 0.974638
R268 source.n42 source.n40 0.974638
R269 source.n44 source.n42 0.974638
R270 source.n46 source.n44 0.974638
R271 source.n47 source.n46 0.974638
R272 source.n12 source.n11 0.470328
R273 source.n36 source.n35 0.470328
R274 source source.n48 0.188
R275 plus.n14 plus.n13 161.3
R276 plus.n15 plus.n8 161.3
R277 plus.n17 plus.n16 161.3
R278 plus.n18 plus.n7 161.3
R279 plus.n19 plus.n6 161.3
R280 plus.n24 plus.n23 161.3
R281 plus.n25 plus.n4 161.3
R282 plus.n27 plus.n26 161.3
R283 plus.n28 plus.n3 161.3
R284 plus.n30 plus.n29 161.3
R285 plus.n33 plus.n0 161.3
R286 plus.n35 plus.n34 161.3
R287 plus.n50 plus.n49 161.3
R288 plus.n51 plus.n44 161.3
R289 plus.n53 plus.n52 161.3
R290 plus.n54 plus.n43 161.3
R291 plus.n55 plus.n42 161.3
R292 plus.n60 plus.n59 161.3
R293 plus.n61 plus.n40 161.3
R294 plus.n63 plus.n62 161.3
R295 plus.n64 plus.n39 161.3
R296 plus.n66 plus.n65 161.3
R297 plus.n69 plus.n36 161.3
R298 plus.n71 plus.n70 161.3
R299 plus.n10 plus.t23 160.916
R300 plus.n46 plus.t4 160.916
R301 plus.n34 plus.t6 139.48
R302 plus.n32 plus.t8 139.48
R303 plus.n31 plus.t9 139.48
R304 plus.n3 plus.t11 139.48
R305 plus.n25 plus.t13 139.48
R306 plus.n5 plus.t16 139.48
R307 plus.n20 plus.t17 139.48
R308 plus.n18 plus.t21 139.48
R309 plus.n8 plus.t18 139.48
R310 plus.n12 plus.t19 139.48
R311 plus.n11 plus.t22 139.48
R312 plus.n70 plus.t10 139.48
R313 plus.n68 plus.t3 139.48
R314 plus.n67 plus.t20 139.48
R315 plus.n39 plus.t2 139.48
R316 plus.n61 plus.t7 139.48
R317 plus.n41 plus.t1 139.48
R318 plus.n56 plus.t15 139.48
R319 plus.n54 plus.t0 139.48
R320 plus.n44 plus.t14 139.48
R321 plus.n48 plus.t5 139.48
R322 plus.n47 plus.t12 139.48
R323 plus.n12 plus.n9 80.6037
R324 plus.n21 plus.n20 80.6037
R325 plus.n22 plus.n5 80.6037
R326 plus.n31 plus.n2 80.6037
R327 plus.n32 plus.n1 80.6037
R328 plus.n48 plus.n45 80.6037
R329 plus.n57 plus.n56 80.6037
R330 plus.n58 plus.n41 80.6037
R331 plus.n67 plus.n38 80.6037
R332 plus.n68 plus.n37 80.6037
R333 plus.n32 plus.n31 48.2005
R334 plus.n20 plus.n5 48.2005
R335 plus.n12 plus.n11 48.2005
R336 plus.n68 plus.n67 48.2005
R337 plus.n56 plus.n41 48.2005
R338 plus.n48 plus.n47 48.2005
R339 plus.n31 plus.n30 44.549
R340 plus.n13 plus.n12 44.549
R341 plus.n67 plus.n66 44.549
R342 plus.n49 plus.n48 44.549
R343 plus.n24 plus.n5 41.6278
R344 plus.n20 plus.n19 41.6278
R345 plus.n60 plus.n41 41.6278
R346 plus.n56 plus.n55 41.6278
R347 plus.n33 plus.n32 38.7066
R348 plus.n69 plus.n68 38.7066
R349 plus plus.n71 33.5937
R350 plus.n10 plus.n9 31.6825
R351 plus.n46 plus.n45 31.6825
R352 plus.n26 plus.n3 25.5611
R353 plus.n17 plus.n8 25.5611
R354 plus.n62 plus.n39 25.5611
R355 plus.n53 plus.n44 25.5611
R356 plus.n26 plus.n25 22.6399
R357 plus.n18 plus.n17 22.6399
R358 plus.n62 plus.n61 22.6399
R359 plus.n54 plus.n53 22.6399
R360 plus.n11 plus.n10 17.2341
R361 plus.n47 plus.n46 17.2341
R362 plus.n34 plus.n33 9.49444
R363 plus.n70 plus.n69 9.49444
R364 plus plus.n35 8.89444
R365 plus.n25 plus.n24 6.57323
R366 plus.n19 plus.n18 6.57323
R367 plus.n61 plus.n60 6.57323
R368 plus.n55 plus.n54 6.57323
R369 plus.n30 plus.n3 3.65202
R370 plus.n13 plus.n8 3.65202
R371 plus.n66 plus.n39 3.65202
R372 plus.n49 plus.n44 3.65202
R373 plus.n22 plus.n21 0.380177
R374 plus.n2 plus.n1 0.380177
R375 plus.n38 plus.n37 0.380177
R376 plus.n58 plus.n57 0.380177
R377 plus.n14 plus.n9 0.285035
R378 plus.n21 plus.n6 0.285035
R379 plus.n23 plus.n22 0.285035
R380 plus.n29 plus.n2 0.285035
R381 plus.n1 plus.n0 0.285035
R382 plus.n37 plus.n36 0.285035
R383 plus.n65 plus.n38 0.285035
R384 plus.n59 plus.n58 0.285035
R385 plus.n57 plus.n42 0.285035
R386 plus.n50 plus.n45 0.285035
R387 plus.n15 plus.n14 0.189894
R388 plus.n16 plus.n15 0.189894
R389 plus.n16 plus.n7 0.189894
R390 plus.n7 plus.n6 0.189894
R391 plus.n23 plus.n4 0.189894
R392 plus.n27 plus.n4 0.189894
R393 plus.n28 plus.n27 0.189894
R394 plus.n29 plus.n28 0.189894
R395 plus.n35 plus.n0 0.189894
R396 plus.n71 plus.n36 0.189894
R397 plus.n65 plus.n64 0.189894
R398 plus.n64 plus.n63 0.189894
R399 plus.n63 plus.n40 0.189894
R400 plus.n59 plus.n40 0.189894
R401 plus.n43 plus.n42 0.189894
R402 plus.n52 plus.n43 0.189894
R403 plus.n52 plus.n51 0.189894
R404 plus.n51 plus.n50 0.189894
R405 drain_left.n13 drain_left.n11 80.7472
R406 drain_left.n7 drain_left.n5 80.7471
R407 drain_left.n2 drain_left.n0 80.7471
R408 drain_left.n21 drain_left.n20 79.7731
R409 drain_left.n19 drain_left.n18 79.7731
R410 drain_left.n17 drain_left.n16 79.7731
R411 drain_left.n15 drain_left.n14 79.7731
R412 drain_left.n13 drain_left.n12 79.7731
R413 drain_left.n7 drain_left.n6 79.773
R414 drain_left.n9 drain_left.n8 79.773
R415 drain_left.n4 drain_left.n3 79.773
R416 drain_left.n2 drain_left.n1 79.773
R417 drain_left drain_left.n10 29.8032
R418 drain_left drain_left.n21 6.62735
R419 drain_left.n5 drain_left.t11 6.6005
R420 drain_left.n5 drain_left.t19 6.6005
R421 drain_left.n6 drain_left.t9 6.6005
R422 drain_left.n6 drain_left.t18 6.6005
R423 drain_left.n8 drain_left.t8 6.6005
R424 drain_left.n8 drain_left.t23 6.6005
R425 drain_left.n3 drain_left.t16 6.6005
R426 drain_left.n3 drain_left.t22 6.6005
R427 drain_left.n1 drain_left.t3 6.6005
R428 drain_left.n1 drain_left.t21 6.6005
R429 drain_left.n0 drain_left.t13 6.6005
R430 drain_left.n0 drain_left.t20 6.6005
R431 drain_left.n20 drain_left.t15 6.6005
R432 drain_left.n20 drain_left.t17 6.6005
R433 drain_left.n18 drain_left.t12 6.6005
R434 drain_left.n18 drain_left.t14 6.6005
R435 drain_left.n16 drain_left.t7 6.6005
R436 drain_left.n16 drain_left.t10 6.6005
R437 drain_left.n14 drain_left.t2 6.6005
R438 drain_left.n14 drain_left.t6 6.6005
R439 drain_left.n12 drain_left.t4 6.6005
R440 drain_left.n12 drain_left.t5 6.6005
R441 drain_left.n11 drain_left.t0 6.6005
R442 drain_left.n11 drain_left.t1 6.6005
R443 drain_left.n9 drain_left.n7 0.974638
R444 drain_left.n4 drain_left.n2 0.974638
R445 drain_left.n15 drain_left.n13 0.974638
R446 drain_left.n17 drain_left.n15 0.974638
R447 drain_left.n19 drain_left.n17 0.974638
R448 drain_left.n21 drain_left.n19 0.974638
R449 drain_left.n10 drain_left.n9 0.432223
R450 drain_left.n10 drain_left.n4 0.432223
C0 source plus 5.57721f
C1 drain_left drain_right 2.02887f
C2 minus source 5.56321f
C3 drain_right plus 0.532688f
C4 drain_right minus 4.61784f
C5 drain_left plus 4.98517f
C6 drain_left minus 0.180512f
C7 drain_right source 10.383699f
C8 minus plus 6.04905f
C9 drain_left source 10.3806f
C10 drain_right a_n3654_n1488# 6.71806f
C11 drain_left a_n3654_n1488# 7.25026f
C12 source a_n3654_n1488# 4.334909f
C13 minus a_n3654_n1488# 14.078671f
C14 plus a_n3654_n1488# 15.56008f
C15 drain_left.t13 a_n3654_n1488# 0.072354f
C16 drain_left.t20 a_n3654_n1488# 0.072354f
C17 drain_left.n0 a_n3654_n1488# 0.527216f
C18 drain_left.t3 a_n3654_n1488# 0.072354f
C19 drain_left.t21 a_n3654_n1488# 0.072354f
C20 drain_left.n1 a_n3654_n1488# 0.521808f
C21 drain_left.n2 a_n3654_n1488# 0.878701f
C22 drain_left.t16 a_n3654_n1488# 0.072354f
C23 drain_left.t22 a_n3654_n1488# 0.072354f
C24 drain_left.n3 a_n3654_n1488# 0.521808f
C25 drain_left.n4 a_n3654_n1488# 0.384204f
C26 drain_left.t11 a_n3654_n1488# 0.072354f
C27 drain_left.t19 a_n3654_n1488# 0.072354f
C28 drain_left.n5 a_n3654_n1488# 0.527216f
C29 drain_left.t9 a_n3654_n1488# 0.072354f
C30 drain_left.t18 a_n3654_n1488# 0.072354f
C31 drain_left.n6 a_n3654_n1488# 0.521808f
C32 drain_left.n7 a_n3654_n1488# 0.878701f
C33 drain_left.t8 a_n3654_n1488# 0.072354f
C34 drain_left.t23 a_n3654_n1488# 0.072354f
C35 drain_left.n8 a_n3654_n1488# 0.521808f
C36 drain_left.n9 a_n3654_n1488# 0.384204f
C37 drain_left.n10 a_n3654_n1488# 1.51272f
C38 drain_left.t0 a_n3654_n1488# 0.072354f
C39 drain_left.t1 a_n3654_n1488# 0.072354f
C40 drain_left.n11 a_n3654_n1488# 0.527218f
C41 drain_left.t4 a_n3654_n1488# 0.072354f
C42 drain_left.t5 a_n3654_n1488# 0.072354f
C43 drain_left.n12 a_n3654_n1488# 0.521811f
C44 drain_left.n13 a_n3654_n1488# 0.878696f
C45 drain_left.t2 a_n3654_n1488# 0.072354f
C46 drain_left.t6 a_n3654_n1488# 0.072354f
C47 drain_left.n14 a_n3654_n1488# 0.521811f
C48 drain_left.n15 a_n3654_n1488# 0.435905f
C49 drain_left.t7 a_n3654_n1488# 0.072354f
C50 drain_left.t10 a_n3654_n1488# 0.072354f
C51 drain_left.n16 a_n3654_n1488# 0.521811f
C52 drain_left.n17 a_n3654_n1488# 0.435905f
C53 drain_left.t12 a_n3654_n1488# 0.072354f
C54 drain_left.t14 a_n3654_n1488# 0.072354f
C55 drain_left.n18 a_n3654_n1488# 0.521811f
C56 drain_left.n19 a_n3654_n1488# 0.435905f
C57 drain_left.t15 a_n3654_n1488# 0.072354f
C58 drain_left.t17 a_n3654_n1488# 0.072354f
C59 drain_left.n20 a_n3654_n1488# 0.521811f
C60 drain_left.n21 a_n3654_n1488# 0.709578f
C61 plus.n0 a_n3654_n1488# 0.053715f
C62 plus.t6 a_n3654_n1488# 0.2897f
C63 plus.t8 a_n3654_n1488# 0.2897f
C64 plus.n1 a_n3654_n1488# 0.067049f
C65 plus.t9 a_n3654_n1488# 0.2897f
C66 plus.n2 a_n3654_n1488# 0.067049f
C67 plus.t11 a_n3654_n1488# 0.2897f
C68 plus.n3 a_n3654_n1488# 0.165048f
C69 plus.n4 a_n3654_n1488# 0.040254f
C70 plus.t13 a_n3654_n1488# 0.2897f
C71 plus.t16 a_n3654_n1488# 0.2897f
C72 plus.n5 a_n3654_n1488# 0.176292f
C73 plus.n6 a_n3654_n1488# 0.053715f
C74 plus.t17 a_n3654_n1488# 0.2897f
C75 plus.t21 a_n3654_n1488# 0.2897f
C76 plus.n7 a_n3654_n1488# 0.040254f
C77 plus.t18 a_n3654_n1488# 0.2897f
C78 plus.n8 a_n3654_n1488# 0.165048f
C79 plus.n9 a_n3654_n1488# 0.231367f
C80 plus.t19 a_n3654_n1488# 0.2897f
C81 plus.t22 a_n3654_n1488# 0.2897f
C82 plus.t23 a_n3654_n1488# 0.312139f
C83 plus.n10 a_n3654_n1488# 0.149829f
C84 plus.n11 a_n3654_n1488# 0.176768f
C85 plus.n12 a_n3654_n1488# 0.176788f
C86 plus.n13 a_n3654_n1488# 0.009135f
C87 plus.n14 a_n3654_n1488# 0.053715f
C88 plus.n15 a_n3654_n1488# 0.040254f
C89 plus.n16 a_n3654_n1488# 0.040254f
C90 plus.n17 a_n3654_n1488# 0.009135f
C91 plus.n18 a_n3654_n1488# 0.165048f
C92 plus.n19 a_n3654_n1488# 0.009135f
C93 plus.n20 a_n3654_n1488# 0.176292f
C94 plus.n21 a_n3654_n1488# 0.067049f
C95 plus.n22 a_n3654_n1488# 0.067049f
C96 plus.n23 a_n3654_n1488# 0.053715f
C97 plus.n24 a_n3654_n1488# 0.009135f
C98 plus.n25 a_n3654_n1488# 0.165048f
C99 plus.n26 a_n3654_n1488# 0.009135f
C100 plus.n27 a_n3654_n1488# 0.040254f
C101 plus.n28 a_n3654_n1488# 0.040254f
C102 plus.n29 a_n3654_n1488# 0.053715f
C103 plus.n30 a_n3654_n1488# 0.009135f
C104 plus.n31 a_n3654_n1488# 0.176788f
C105 plus.n32 a_n3654_n1488# 0.175796f
C106 plus.n33 a_n3654_n1488# 0.009135f
C107 plus.n34 a_n3654_n1488# 0.161697f
C108 plus.n35 a_n3654_n1488# 0.316525f
C109 plus.n36 a_n3654_n1488# 0.053715f
C110 plus.t10 a_n3654_n1488# 0.2897f
C111 plus.n37 a_n3654_n1488# 0.067049f
C112 plus.t3 a_n3654_n1488# 0.2897f
C113 plus.n38 a_n3654_n1488# 0.067049f
C114 plus.t20 a_n3654_n1488# 0.2897f
C115 plus.t2 a_n3654_n1488# 0.2897f
C116 plus.n39 a_n3654_n1488# 0.165048f
C117 plus.n40 a_n3654_n1488# 0.040254f
C118 plus.t7 a_n3654_n1488# 0.2897f
C119 plus.t1 a_n3654_n1488# 0.2897f
C120 plus.n41 a_n3654_n1488# 0.176292f
C121 plus.n42 a_n3654_n1488# 0.053715f
C122 plus.t15 a_n3654_n1488# 0.2897f
C123 plus.n43 a_n3654_n1488# 0.040254f
C124 plus.t0 a_n3654_n1488# 0.2897f
C125 plus.t14 a_n3654_n1488# 0.2897f
C126 plus.n44 a_n3654_n1488# 0.165048f
C127 plus.n45 a_n3654_n1488# 0.231367f
C128 plus.t5 a_n3654_n1488# 0.2897f
C129 plus.t4 a_n3654_n1488# 0.312139f
C130 plus.n46 a_n3654_n1488# 0.149829f
C131 plus.t12 a_n3654_n1488# 0.2897f
C132 plus.n47 a_n3654_n1488# 0.176768f
C133 plus.n48 a_n3654_n1488# 0.176788f
C134 plus.n49 a_n3654_n1488# 0.009135f
C135 plus.n50 a_n3654_n1488# 0.053715f
C136 plus.n51 a_n3654_n1488# 0.040254f
C137 plus.n52 a_n3654_n1488# 0.040254f
C138 plus.n53 a_n3654_n1488# 0.009135f
C139 plus.n54 a_n3654_n1488# 0.165048f
C140 plus.n55 a_n3654_n1488# 0.009135f
C141 plus.n56 a_n3654_n1488# 0.176292f
C142 plus.n57 a_n3654_n1488# 0.067049f
C143 plus.n58 a_n3654_n1488# 0.067049f
C144 plus.n59 a_n3654_n1488# 0.053715f
C145 plus.n60 a_n3654_n1488# 0.009135f
C146 plus.n61 a_n3654_n1488# 0.165048f
C147 plus.n62 a_n3654_n1488# 0.009135f
C148 plus.n63 a_n3654_n1488# 0.040254f
C149 plus.n64 a_n3654_n1488# 0.040254f
C150 plus.n65 a_n3654_n1488# 0.053715f
C151 plus.n66 a_n3654_n1488# 0.009135f
C152 plus.n67 a_n3654_n1488# 0.176788f
C153 plus.n68 a_n3654_n1488# 0.175796f
C154 plus.n69 a_n3654_n1488# 0.009135f
C155 plus.n70 a_n3654_n1488# 0.161697f
C156 plus.n71 a_n3654_n1488# 1.34762f
C157 source.t12 a_n3654_n1488# 0.585419f
C158 source.n0 a_n3654_n1488# 0.87121f
C159 source.t4 a_n3654_n1488# 0.0705f
C160 source.t9 a_n3654_n1488# 0.0705f
C161 source.n1 a_n3654_n1488# 0.44701f
C162 source.n2 a_n3654_n1488# 0.445747f
C163 source.t11 a_n3654_n1488# 0.0705f
C164 source.t10 a_n3654_n1488# 0.0705f
C165 source.n3 a_n3654_n1488# 0.44701f
C166 source.n4 a_n3654_n1488# 0.445747f
C167 source.t15 a_n3654_n1488# 0.0705f
C168 source.t13 a_n3654_n1488# 0.0705f
C169 source.n5 a_n3654_n1488# 0.44701f
C170 source.n6 a_n3654_n1488# 0.445747f
C171 source.t44 a_n3654_n1488# 0.0705f
C172 source.t2 a_n3654_n1488# 0.0705f
C173 source.n7 a_n3654_n1488# 0.44701f
C174 source.n8 a_n3654_n1488# 0.445747f
C175 source.t43 a_n3654_n1488# 0.0705f
C176 source.t46 a_n3654_n1488# 0.0705f
C177 source.n9 a_n3654_n1488# 0.44701f
C178 source.n10 a_n3654_n1488# 0.445747f
C179 source.t16 a_n3654_n1488# 0.585419f
C180 source.n11 a_n3654_n1488# 0.451286f
C181 source.t27 a_n3654_n1488# 0.585419f
C182 source.n12 a_n3654_n1488# 0.451286f
C183 source.t34 a_n3654_n1488# 0.0705f
C184 source.t32 a_n3654_n1488# 0.0705f
C185 source.n13 a_n3654_n1488# 0.44701f
C186 source.n14 a_n3654_n1488# 0.445747f
C187 source.t21 a_n3654_n1488# 0.0705f
C188 source.t23 a_n3654_n1488# 0.0705f
C189 source.n15 a_n3654_n1488# 0.44701f
C190 source.n16 a_n3654_n1488# 0.445747f
C191 source.t29 a_n3654_n1488# 0.0705f
C192 source.t26 a_n3654_n1488# 0.0705f
C193 source.n17 a_n3654_n1488# 0.44701f
C194 source.n18 a_n3654_n1488# 0.445747f
C195 source.t22 a_n3654_n1488# 0.0705f
C196 source.t20 a_n3654_n1488# 0.0705f
C197 source.n19 a_n3654_n1488# 0.44701f
C198 source.n20 a_n3654_n1488# 0.445747f
C199 source.t28 a_n3654_n1488# 0.0705f
C200 source.t36 a_n3654_n1488# 0.0705f
C201 source.n21 a_n3654_n1488# 0.44701f
C202 source.n22 a_n3654_n1488# 0.445747f
C203 source.t31 a_n3654_n1488# 0.585419f
C204 source.n23 a_n3654_n1488# 1.19129f
C205 source.t14 a_n3654_n1488# 0.585416f
C206 source.n24 a_n3654_n1488# 1.1913f
C207 source.t6 a_n3654_n1488# 0.0705f
C208 source.t5 a_n3654_n1488# 0.0705f
C209 source.n25 a_n3654_n1488# 0.447007f
C210 source.n26 a_n3654_n1488# 0.44575f
C211 source.t47 a_n3654_n1488# 0.0705f
C212 source.t1 a_n3654_n1488# 0.0705f
C213 source.n27 a_n3654_n1488# 0.447007f
C214 source.n28 a_n3654_n1488# 0.44575f
C215 source.t45 a_n3654_n1488# 0.0705f
C216 source.t17 a_n3654_n1488# 0.0705f
C217 source.n29 a_n3654_n1488# 0.447007f
C218 source.n30 a_n3654_n1488# 0.44575f
C219 source.t3 a_n3654_n1488# 0.0705f
C220 source.t7 a_n3654_n1488# 0.0705f
C221 source.n31 a_n3654_n1488# 0.447007f
C222 source.n32 a_n3654_n1488# 0.44575f
C223 source.t0 a_n3654_n1488# 0.0705f
C224 source.t8 a_n3654_n1488# 0.0705f
C225 source.n33 a_n3654_n1488# 0.447007f
C226 source.n34 a_n3654_n1488# 0.44575f
C227 source.t42 a_n3654_n1488# 0.585416f
C228 source.n35 a_n3654_n1488# 0.451289f
C229 source.t38 a_n3654_n1488# 0.585416f
C230 source.n36 a_n3654_n1488# 0.451289f
C231 source.t33 a_n3654_n1488# 0.0705f
C232 source.t37 a_n3654_n1488# 0.0705f
C233 source.n37 a_n3654_n1488# 0.447007f
C234 source.n38 a_n3654_n1488# 0.44575f
C235 source.t30 a_n3654_n1488# 0.0705f
C236 source.t41 a_n3654_n1488# 0.0705f
C237 source.n39 a_n3654_n1488# 0.447007f
C238 source.n40 a_n3654_n1488# 0.44575f
C239 source.t24 a_n3654_n1488# 0.0705f
C240 source.t40 a_n3654_n1488# 0.0705f
C241 source.n41 a_n3654_n1488# 0.447007f
C242 source.n42 a_n3654_n1488# 0.44575f
C243 source.t25 a_n3654_n1488# 0.0705f
C244 source.t39 a_n3654_n1488# 0.0705f
C245 source.n43 a_n3654_n1488# 0.447007f
C246 source.n44 a_n3654_n1488# 0.44575f
C247 source.t19 a_n3654_n1488# 0.0705f
C248 source.t35 a_n3654_n1488# 0.0705f
C249 source.n45 a_n3654_n1488# 0.447007f
C250 source.n46 a_n3654_n1488# 0.44575f
C251 source.t18 a_n3654_n1488# 0.585416f
C252 source.n47 a_n3654_n1488# 0.65171f
C253 source.n48 a_n3654_n1488# 0.880821f
C254 drain_right.t3 a_n3654_n1488# 0.071179f
C255 drain_right.t8 a_n3654_n1488# 0.071179f
C256 drain_right.n0 a_n3654_n1488# 0.518654f
C257 drain_right.t4 a_n3654_n1488# 0.071179f
C258 drain_right.t9 a_n3654_n1488# 0.071179f
C259 drain_right.n1 a_n3654_n1488# 0.513335f
C260 drain_right.n2 a_n3654_n1488# 0.864433f
C261 drain_right.t0 a_n3654_n1488# 0.071179f
C262 drain_right.t17 a_n3654_n1488# 0.071179f
C263 drain_right.n3 a_n3654_n1488# 0.513335f
C264 drain_right.n4 a_n3654_n1488# 0.377965f
C265 drain_right.t6 a_n3654_n1488# 0.071179f
C266 drain_right.t23 a_n3654_n1488# 0.071179f
C267 drain_right.n5 a_n3654_n1488# 0.518654f
C268 drain_right.t2 a_n3654_n1488# 0.071179f
C269 drain_right.t22 a_n3654_n1488# 0.071179f
C270 drain_right.n6 a_n3654_n1488# 0.513335f
C271 drain_right.n7 a_n3654_n1488# 0.864433f
C272 drain_right.t1 a_n3654_n1488# 0.071179f
C273 drain_right.t16 a_n3654_n1488# 0.071179f
C274 drain_right.n8 a_n3654_n1488# 0.513335f
C275 drain_right.n9 a_n3654_n1488# 0.377965f
C276 drain_right.n10 a_n3654_n1488# 1.42983f
C277 drain_right.t12 a_n3654_n1488# 0.071179f
C278 drain_right.t11 a_n3654_n1488# 0.071179f
C279 drain_right.n11 a_n3654_n1488# 0.518657f
C280 drain_right.t18 a_n3654_n1488# 0.071179f
C281 drain_right.t7 a_n3654_n1488# 0.071179f
C282 drain_right.n12 a_n3654_n1488# 0.513338f
C283 drain_right.n13 a_n3654_n1488# 0.864428f
C284 drain_right.t15 a_n3654_n1488# 0.071179f
C285 drain_right.t20 a_n3654_n1488# 0.071179f
C286 drain_right.n14 a_n3654_n1488# 0.513338f
C287 drain_right.n15 a_n3654_n1488# 0.428827f
C288 drain_right.t21 a_n3654_n1488# 0.071179f
C289 drain_right.t14 a_n3654_n1488# 0.071179f
C290 drain_right.n16 a_n3654_n1488# 0.513338f
C291 drain_right.n17 a_n3654_n1488# 0.428827f
C292 drain_right.t5 a_n3654_n1488# 0.071179f
C293 drain_right.t19 a_n3654_n1488# 0.071179f
C294 drain_right.n18 a_n3654_n1488# 0.513338f
C295 drain_right.n19 a_n3654_n1488# 0.428827f
C296 drain_right.t13 a_n3654_n1488# 0.071179f
C297 drain_right.t10 a_n3654_n1488# 0.071179f
C298 drain_right.n20 a_n3654_n1488# 0.513338f
C299 drain_right.n21 a_n3654_n1488# 0.698055f
C300 minus.n0 a_n3654_n1488# 0.052164f
C301 minus.t5 a_n3654_n1488# 0.28134f
C302 minus.n1 a_n3654_n1488# 0.171686f
C303 minus.t13 a_n3654_n1488# 0.28134f
C304 minus.n2 a_n3654_n1488# 0.039093f
C305 minus.t21 a_n3654_n1488# 0.28134f
C306 minus.n3 a_n3654_n1488# 0.160285f
C307 minus.n4 a_n3654_n1488# 0.065114f
C308 minus.n5 a_n3654_n1488# 0.008871f
C309 minus.t15 a_n3654_n1488# 0.28134f
C310 minus.n6 a_n3654_n1488# 0.039093f
C311 minus.n7 a_n3654_n1488# 0.008871f
C312 minus.t18 a_n3654_n1488# 0.28134f
C313 minus.t14 a_n3654_n1488# 0.303131f
C314 minus.n8 a_n3654_n1488# 0.145505f
C315 minus.t9 a_n3654_n1488# 0.28134f
C316 minus.n9 a_n3654_n1488# 0.171666f
C317 minus.t7 a_n3654_n1488# 0.28134f
C318 minus.n10 a_n3654_n1488# 0.171686f
C319 minus.n11 a_n3654_n1488# 0.22469f
C320 minus.n12 a_n3654_n1488# 0.052164f
C321 minus.n13 a_n3654_n1488# 0.039093f
C322 minus.n14 a_n3654_n1488# 0.160285f
C323 minus.n15 a_n3654_n1488# 0.008871f
C324 minus.t20 a_n3654_n1488# 0.28134f
C325 minus.n16 a_n3654_n1488# 0.160285f
C326 minus.n17 a_n3654_n1488# 0.039093f
C327 minus.n18 a_n3654_n1488# 0.052164f
C328 minus.n19 a_n3654_n1488# 0.065114f
C329 minus.n20 a_n3654_n1488# 0.171204f
C330 minus.t12 a_n3654_n1488# 0.28134f
C331 minus.n21 a_n3654_n1488# 0.171204f
C332 minus.n22 a_n3654_n1488# 0.008871f
C333 minus.n23 a_n3654_n1488# 0.052164f
C334 minus.n24 a_n3654_n1488# 0.039093f
C335 minus.n25 a_n3654_n1488# 0.039093f
C336 minus.n26 a_n3654_n1488# 0.008871f
C337 minus.t19 a_n3654_n1488# 0.28134f
C338 minus.n27 a_n3654_n1488# 0.160285f
C339 minus.n28 a_n3654_n1488# 0.008871f
C340 minus.n29 a_n3654_n1488# 0.052164f
C341 minus.n30 a_n3654_n1488# 0.065114f
C342 minus.n31 a_n3654_n1488# 0.065114f
C343 minus.n32 a_n3654_n1488# 0.170722f
C344 minus.n33 a_n3654_n1488# 0.008871f
C345 minus.t10 a_n3654_n1488# 0.28134f
C346 minus.n34 a_n3654_n1488# 0.157031f
C347 minus.n35 a_n3654_n1488# 1.39293f
C348 minus.n36 a_n3654_n1488# 0.052164f
C349 minus.t22 a_n3654_n1488# 0.28134f
C350 minus.n37 a_n3654_n1488# 0.171686f
C351 minus.n38 a_n3654_n1488# 0.039093f
C352 minus.t16 a_n3654_n1488# 0.28134f
C353 minus.n39 a_n3654_n1488# 0.160285f
C354 minus.n40 a_n3654_n1488# 0.065114f
C355 minus.n41 a_n3654_n1488# 0.008871f
C356 minus.n42 a_n3654_n1488# 0.039093f
C357 minus.n43 a_n3654_n1488# 0.008871f
C358 minus.t3 a_n3654_n1488# 0.303131f
C359 minus.n44 a_n3654_n1488# 0.145505f
C360 minus.t8 a_n3654_n1488# 0.28134f
C361 minus.n45 a_n3654_n1488# 0.171666f
C362 minus.t4 a_n3654_n1488# 0.28134f
C363 minus.n46 a_n3654_n1488# 0.171686f
C364 minus.n47 a_n3654_n1488# 0.22469f
C365 minus.n48 a_n3654_n1488# 0.052164f
C366 minus.n49 a_n3654_n1488# 0.039093f
C367 minus.t11 a_n3654_n1488# 0.28134f
C368 minus.n50 a_n3654_n1488# 0.160285f
C369 minus.n51 a_n3654_n1488# 0.008871f
C370 minus.t0 a_n3654_n1488# 0.28134f
C371 minus.n52 a_n3654_n1488# 0.160285f
C372 minus.n53 a_n3654_n1488# 0.039093f
C373 minus.n54 a_n3654_n1488# 0.052164f
C374 minus.n55 a_n3654_n1488# 0.065114f
C375 minus.t17 a_n3654_n1488# 0.28134f
C376 minus.n56 a_n3654_n1488# 0.171204f
C377 minus.t1 a_n3654_n1488# 0.28134f
C378 minus.n57 a_n3654_n1488# 0.171204f
C379 minus.n58 a_n3654_n1488# 0.008871f
C380 minus.n59 a_n3654_n1488# 0.052164f
C381 minus.n60 a_n3654_n1488# 0.039093f
C382 minus.n61 a_n3654_n1488# 0.039093f
C383 minus.n62 a_n3654_n1488# 0.008871f
C384 minus.t2 a_n3654_n1488# 0.28134f
C385 minus.n63 a_n3654_n1488# 0.160285f
C386 minus.n64 a_n3654_n1488# 0.008871f
C387 minus.n65 a_n3654_n1488# 0.052164f
C388 minus.n66 a_n3654_n1488# 0.065114f
C389 minus.n67 a_n3654_n1488# 0.065114f
C390 minus.t6 a_n3654_n1488# 0.28134f
C391 minus.n68 a_n3654_n1488# 0.170722f
C392 minus.n69 a_n3654_n1488# 0.008871f
C393 minus.t23 a_n3654_n1488# 0.28134f
C394 minus.n70 a_n3654_n1488# 0.157031f
C395 minus.n71 a_n3654_n1488# 0.270167f
C396 minus.n72 a_n3654_n1488# 1.68656f
.ends

