* NGSPICE file created from diffpair185.ext - technology: sky130A

.subckt diffpair185 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t20 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 drain_left.t10 plus.t1 source.t16 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 source.t4 minus.t0 drain_right.t11 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X3 drain_right.t10 minus.t1 source.t5 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X4 source.t8 minus.t2 drain_right.t9 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X5 a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X6 source.t12 plus.t2 drain_left.t9 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X7 source.t14 plus.t3 drain_left.t8 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X8 a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X9 drain_left.t7 plus.t4 source.t21 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X10 drain_left.t6 plus.t5 source.t13 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X11 source.t3 minus.t3 drain_right.t8 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X12 drain_left.t5 plus.t6 source.t18 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X13 source.t15 plus.t7 drain_left.t4 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X14 source.t11 plus.t8 drain_left.t3 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X15 source.t17 plus.t9 drain_left.t2 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X16 a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X17 source.t19 plus.t10 drain_left.t1 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 drain_right.t7 minus.t4 source.t6 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X19 drain_right.t6 minus.t5 source.t7 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X20 drain_right.t5 minus.t6 source.t0 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X21 drain_right.t4 minus.t7 source.t1 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X22 a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X23 source.t2 minus.t8 drain_right.t3 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X24 drain_right.t2 minus.t9 source.t9 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X25 source.t22 minus.t10 drain_right.t1 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X26 drain_left.t0 plus.t11 source.t10 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X27 source.t23 minus.t11 drain_right.t0 a_n1528_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n2 plus.t2 443.733
R1 plus.n13 plus.t11 443.733
R2 plus.n17 plus.t5 443.733
R3 plus.n28 plus.t7 443.733
R4 plus.n3 plus.t1 414.521
R5 plus.n4 plus.t9 414.521
R6 plus.n10 plus.t0 414.521
R7 plus.n12 plus.t8 414.521
R8 plus.n19 plus.t3 414.521
R9 plus.n18 plus.t6 414.521
R10 plus.n25 plus.t10 414.521
R11 plus.n27 plus.t4 414.521
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 25.3172
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 8.67095
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n0 source.t10 69.6943
R53 source.n5 source.t12 69.6943
R54 source.n6 source.t7 69.6943
R55 source.n11 source.t3 69.6943
R56 source.n23 source.t5 69.6942
R57 source.n18 source.t23 69.6942
R58 source.n17 source.t13 69.6942
R59 source.n12 source.t15 69.6942
R60 source.n2 source.n1 63.0943
R61 source.n4 source.n3 63.0943
R62 source.n8 source.n7 63.0943
R63 source.n10 source.n9 63.0943
R64 source.n22 source.n21 63.0942
R65 source.n20 source.n19 63.0942
R66 source.n16 source.n15 63.0942
R67 source.n14 source.n13 63.0942
R68 source.n12 source.n11 14.9695
R69 source.n24 source.n0 9.45661
R70 source.n21 source.t1 6.6005
R71 source.n21 source.t22 6.6005
R72 source.n19 source.t0 6.6005
R73 source.n19 source.t2 6.6005
R74 source.n15 source.t18 6.6005
R75 source.n15 source.t14 6.6005
R76 source.n13 source.t21 6.6005
R77 source.n13 source.t19 6.6005
R78 source.n1 source.t20 6.6005
R79 source.n1 source.t11 6.6005
R80 source.n3 source.t16 6.6005
R81 source.n3 source.t17 6.6005
R82 source.n7 source.t6 6.6005
R83 source.n7 source.t8 6.6005
R84 source.n9 source.t9 6.6005
R85 source.n9 source.t4 6.6005
R86 source.n24 source.n23 5.51343
R87 source.n11 source.n10 0.5005
R88 source.n10 source.n8 0.5005
R89 source.n8 source.n6 0.5005
R90 source.n5 source.n4 0.5005
R91 source.n4 source.n2 0.5005
R92 source.n2 source.n0 0.5005
R93 source.n14 source.n12 0.5005
R94 source.n16 source.n14 0.5005
R95 source.n17 source.n16 0.5005
R96 source.n20 source.n18 0.5005
R97 source.n22 source.n20 0.5005
R98 source.n23 source.n22 0.5005
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 80.2731
R103 drain_left.n3 drain_left.n2 80.2177
R104 drain_left.n3 drain_left.n0 80.2177
R105 drain_left.n8 drain_left.n7 79.7731
R106 drain_left.n6 drain_left.n5 79.7731
R107 drain_left.n3 drain_left.n1 79.773
R108 drain_left drain_left.n3 23.0489
R109 drain_left.n1 drain_left.t1 6.6005
R110 drain_left.n1 drain_left.t5 6.6005
R111 drain_left.n2 drain_left.t8 6.6005
R112 drain_left.n2 drain_left.t6 6.6005
R113 drain_left.n0 drain_left.t4 6.6005
R114 drain_left.n0 drain_left.t7 6.6005
R115 drain_left.n7 drain_left.t3 6.6005
R116 drain_left.n7 drain_left.t0 6.6005
R117 drain_left.n5 drain_left.t2 6.6005
R118 drain_left.n5 drain_left.t11 6.6005
R119 drain_left.n4 drain_left.t9 6.6005
R120 drain_left.n4 drain_left.t10 6.6005
R121 drain_left drain_left.n8 6.15322
R122 drain_left.n8 drain_left.n6 0.5005
R123 minus.n13 minus.t3 443.733
R124 minus.n2 minus.t5 443.733
R125 minus.n28 minus.t1 443.733
R126 minus.n17 minus.t11 443.733
R127 minus.n12 minus.t9 414.521
R128 minus.n10 minus.t0 414.521
R129 minus.n3 minus.t4 414.521
R130 minus.n4 minus.t2 414.521
R131 minus.n27 minus.t10 414.521
R132 minus.n25 minus.t7 414.521
R133 minus.n19 minus.t8 414.521
R134 minus.n18 minus.t6 414.521
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 67.1884
R150 minus.n5 minus.n3 67.1884
R151 minus.n20 minus.n19 67.1884
R152 minus.n26 minus.n25 67.1884
R153 minus.n13 minus.n12 55.5035
R154 minus.n4 minus.n2 55.5035
R155 minus.n18 minus.n17 55.5035
R156 minus.n28 minus.n27 55.5035
R157 minus.n30 minus.n14 28.027
R158 minus.n12 minus.n11 17.5278
R159 minus.n5 minus.n4 17.5278
R160 minus.n20 minus.n18 17.5278
R161 minus.n27 minus.n26 17.5278
R162 minus.n30 minus.n29 6.43611
R163 minus.n10 minus.n9 5.84292
R164 minus.n3 minus.n1 5.84292
R165 minus.n19 minus.n16 5.84292
R166 minus.n25 minus.n24 5.84292
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 80.2731
R177 drain_right.n3 drain_right.n2 80.2177
R178 drain_right.n3 drain_right.n0 80.2177
R179 drain_right.n6 drain_right.n5 79.7731
R180 drain_right.n8 drain_right.n7 79.7731
R181 drain_right.n3 drain_right.n1 79.773
R182 drain_right drain_right.n3 22.4957
R183 drain_right.n1 drain_right.t3 6.6005
R184 drain_right.n1 drain_right.t4 6.6005
R185 drain_right.n2 drain_right.t1 6.6005
R186 drain_right.n2 drain_right.t10 6.6005
R187 drain_right.n0 drain_right.t0 6.6005
R188 drain_right.n0 drain_right.t5 6.6005
R189 drain_right.n4 drain_right.t9 6.6005
R190 drain_right.n4 drain_right.t6 6.6005
R191 drain_right.n5 drain_right.t11 6.6005
R192 drain_right.n5 drain_right.t7 6.6005
R193 drain_right.n7 drain_right.t8 6.6005
R194 drain_right.n7 drain_right.t2 6.6005
R195 drain_right drain_right.n8 6.15322
R196 drain_right.n8 drain_right.n6 0.5005
C0 minus plus 3.40215f
C1 source drain_right 8.09615f
C2 source minus 1.38541f
C3 source plus 1.39941f
C4 drain_right drain_left 0.751108f
C5 minus drain_left 0.175975f
C6 plus drain_left 1.48743f
C7 minus drain_right 1.34128f
C8 plus drain_right 0.305514f
C9 source drain_left 8.0967f
C10 drain_right a_n1528_n1488# 3.78461f
C11 drain_left a_n1528_n1488# 3.99875f
C12 source a_n1528_n1488# 3.5418f
C13 minus a_n1528_n1488# 5.208692f
C14 plus a_n1528_n1488# 5.864906f
C15 drain_right.t0 a_n1528_n1488# 0.067121f
C16 drain_right.t5 a_n1528_n1488# 0.067121f
C17 drain_right.n0 a_n1528_n1488# 0.485878f
C18 drain_right.t3 a_n1528_n1488# 0.067121f
C19 drain_right.t4 a_n1528_n1488# 0.067121f
C20 drain_right.n1 a_n1528_n1488# 0.484073f
C21 drain_right.t1 a_n1528_n1488# 0.067121f
C22 drain_right.t10 a_n1528_n1488# 0.067121f
C23 drain_right.n2 a_n1528_n1488# 0.485878f
C24 drain_right.n3 a_n1528_n1488# 1.63125f
C25 drain_right.t9 a_n1528_n1488# 0.067121f
C26 drain_right.t6 a_n1528_n1488# 0.067121f
C27 drain_right.n4 a_n1528_n1488# 0.486126f
C28 drain_right.t11 a_n1528_n1488# 0.067121f
C29 drain_right.t7 a_n1528_n1488# 0.067121f
C30 drain_right.n5 a_n1528_n1488# 0.484075f
C31 drain_right.n6 a_n1528_n1488# 0.645093f
C32 drain_right.t8 a_n1528_n1488# 0.067121f
C33 drain_right.t2 a_n1528_n1488# 0.067121f
C34 drain_right.n7 a_n1528_n1488# 0.484075f
C35 drain_right.n8 a_n1528_n1488# 0.551575f
C36 minus.n0 a_n1528_n1488# 0.02956f
C37 minus.t3 a_n1528_n1488# 0.066696f
C38 minus.t9 a_n1528_n1488# 0.064202f
C39 minus.t0 a_n1528_n1488# 0.064202f
C40 minus.n1 a_n1528_n1488# 0.010535f
C41 minus.t5 a_n1528_n1488# 0.066696f
C42 minus.n2 a_n1528_n1488# 0.046694f
C43 minus.t4 a_n1528_n1488# 0.064202f
C44 minus.n3 a_n1528_n1488# 0.038797f
C45 minus.t2 a_n1528_n1488# 0.064202f
C46 minus.n4 a_n1528_n1488# 0.038797f
C47 minus.n5 a_n1528_n1488# 0.011264f
C48 minus.n6 a_n1528_n1488# 0.061816f
C49 minus.n7 a_n1528_n1488# 0.02956f
C50 minus.n8 a_n1528_n1488# 0.02956f
C51 minus.n9 a_n1528_n1488# 0.010535f
C52 minus.n10 a_n1528_n1488# 0.038797f
C53 minus.n11 a_n1528_n1488# 0.011264f
C54 minus.n12 a_n1528_n1488# 0.038797f
C55 minus.n13 a_n1528_n1488# 0.046656f
C56 minus.n14 a_n1528_n1488# 0.68135f
C57 minus.n15 a_n1528_n1488# 0.02956f
C58 minus.t10 a_n1528_n1488# 0.064202f
C59 minus.t7 a_n1528_n1488# 0.064202f
C60 minus.n16 a_n1528_n1488# 0.010535f
C61 minus.t11 a_n1528_n1488# 0.066696f
C62 minus.n17 a_n1528_n1488# 0.046694f
C63 minus.t6 a_n1528_n1488# 0.064202f
C64 minus.n18 a_n1528_n1488# 0.038797f
C65 minus.t8 a_n1528_n1488# 0.064202f
C66 minus.n19 a_n1528_n1488# 0.038797f
C67 minus.n20 a_n1528_n1488# 0.011264f
C68 minus.n21 a_n1528_n1488# 0.061816f
C69 minus.n22 a_n1528_n1488# 0.02956f
C70 minus.n23 a_n1528_n1488# 0.02956f
C71 minus.n24 a_n1528_n1488# 0.010535f
C72 minus.n25 a_n1528_n1488# 0.038797f
C73 minus.n26 a_n1528_n1488# 0.011264f
C74 minus.n27 a_n1528_n1488# 0.038797f
C75 minus.t1 a_n1528_n1488# 0.066696f
C76 minus.n28 a_n1528_n1488# 0.046656f
C77 minus.n29 a_n1528_n1488# 0.188794f
C78 minus.n30 a_n1528_n1488# 0.844773f
C79 drain_left.t4 a_n1528_n1488# 0.066216f
C80 drain_left.t7 a_n1528_n1488# 0.066216f
C81 drain_left.n0 a_n1528_n1488# 0.479324f
C82 drain_left.t1 a_n1528_n1488# 0.066216f
C83 drain_left.t5 a_n1528_n1488# 0.066216f
C84 drain_left.n1 a_n1528_n1488# 0.477543f
C85 drain_left.t8 a_n1528_n1488# 0.066216f
C86 drain_left.t6 a_n1528_n1488# 0.066216f
C87 drain_left.n2 a_n1528_n1488# 0.479324f
C88 drain_left.n3 a_n1528_n1488# 1.66481f
C89 drain_left.t9 a_n1528_n1488# 0.066216f
C90 drain_left.t10 a_n1528_n1488# 0.066216f
C91 drain_left.n4 a_n1528_n1488# 0.479569f
C92 drain_left.t2 a_n1528_n1488# 0.066216f
C93 drain_left.t11 a_n1528_n1488# 0.066216f
C94 drain_left.n5 a_n1528_n1488# 0.477546f
C95 drain_left.n6 a_n1528_n1488# 0.636391f
C96 drain_left.t3 a_n1528_n1488# 0.066216f
C97 drain_left.t0 a_n1528_n1488# 0.066216f
C98 drain_left.n7 a_n1528_n1488# 0.477546f
C99 drain_left.n8 a_n1528_n1488# 0.544135f
C100 source.t10 a_n1528_n1488# 0.517595f
C101 source.n0 a_n1528_n1488# 0.699739f
C102 source.t20 a_n1528_n1488# 0.062332f
C103 source.t11 a_n1528_n1488# 0.062332f
C104 source.n1 a_n1528_n1488# 0.395221f
C105 source.n2 a_n1528_n1488# 0.313765f
C106 source.t16 a_n1528_n1488# 0.062332f
C107 source.t17 a_n1528_n1488# 0.062332f
C108 source.n3 a_n1528_n1488# 0.395221f
C109 source.n4 a_n1528_n1488# 0.313765f
C110 source.t12 a_n1528_n1488# 0.517595f
C111 source.n5 a_n1528_n1488# 0.358832f
C112 source.t7 a_n1528_n1488# 0.517595f
C113 source.n6 a_n1528_n1488# 0.358832f
C114 source.t6 a_n1528_n1488# 0.062332f
C115 source.t8 a_n1528_n1488# 0.062332f
C116 source.n7 a_n1528_n1488# 0.395221f
C117 source.n8 a_n1528_n1488# 0.313765f
C118 source.t9 a_n1528_n1488# 0.062332f
C119 source.t4 a_n1528_n1488# 0.062332f
C120 source.n9 a_n1528_n1488# 0.395221f
C121 source.n10 a_n1528_n1488# 0.313765f
C122 source.t3 a_n1528_n1488# 0.517595f
C123 source.n11 a_n1528_n1488# 0.972936f
C124 source.t15 a_n1528_n1488# 0.517592f
C125 source.n12 a_n1528_n1488# 0.972939f
C126 source.t21 a_n1528_n1488# 0.062332f
C127 source.t19 a_n1528_n1488# 0.062332f
C128 source.n13 a_n1528_n1488# 0.395218f
C129 source.n14 a_n1528_n1488# 0.313768f
C130 source.t18 a_n1528_n1488# 0.062332f
C131 source.t14 a_n1528_n1488# 0.062332f
C132 source.n15 a_n1528_n1488# 0.395218f
C133 source.n16 a_n1528_n1488# 0.313768f
C134 source.t13 a_n1528_n1488# 0.517592f
C135 source.n17 a_n1528_n1488# 0.358835f
C136 source.t23 a_n1528_n1488# 0.517592f
C137 source.n18 a_n1528_n1488# 0.358835f
C138 source.t0 a_n1528_n1488# 0.062332f
C139 source.t2 a_n1528_n1488# 0.062332f
C140 source.n19 a_n1528_n1488# 0.395218f
C141 source.n20 a_n1528_n1488# 0.313768f
C142 source.t1 a_n1528_n1488# 0.062332f
C143 source.t22 a_n1528_n1488# 0.062332f
C144 source.n21 a_n1528_n1488# 0.395218f
C145 source.n22 a_n1528_n1488# 0.313768f
C146 source.t5 a_n1528_n1488# 0.517592f
C147 source.n23 a_n1528_n1488# 0.504335f
C148 source.n24 a_n1528_n1488# 0.760503f
C149 plus.n0 a_n1528_n1488# 0.030089f
C150 plus.t8 a_n1528_n1488# 0.065351f
C151 plus.t0 a_n1528_n1488# 0.065351f
C152 plus.n1 a_n1528_n1488# 0.010724f
C153 plus.t2 a_n1528_n1488# 0.06789f
C154 plus.n2 a_n1528_n1488# 0.04753f
C155 plus.t1 a_n1528_n1488# 0.065351f
C156 plus.n3 a_n1528_n1488# 0.039492f
C157 plus.t9 a_n1528_n1488# 0.065351f
C158 plus.n4 a_n1528_n1488# 0.039492f
C159 plus.n5 a_n1528_n1488# 0.011466f
C160 plus.n6 a_n1528_n1488# 0.062923f
C161 plus.n7 a_n1528_n1488# 0.030089f
C162 plus.n8 a_n1528_n1488# 0.030089f
C163 plus.n9 a_n1528_n1488# 0.010724f
C164 plus.n10 a_n1528_n1488# 0.039492f
C165 plus.n11 a_n1528_n1488# 0.011466f
C166 plus.n12 a_n1528_n1488# 0.039492f
C167 plus.t11 a_n1528_n1488# 0.06789f
C168 plus.n13 a_n1528_n1488# 0.047491f
C169 plus.n14 a_n1528_n1488# 0.219984f
C170 plus.n15 a_n1528_n1488# 0.030089f
C171 plus.t7 a_n1528_n1488# 0.06789f
C172 plus.t4 a_n1528_n1488# 0.065351f
C173 plus.t10 a_n1528_n1488# 0.065351f
C174 plus.n16 a_n1528_n1488# 0.010724f
C175 plus.t5 a_n1528_n1488# 0.06789f
C176 plus.n17 a_n1528_n1488# 0.04753f
C177 plus.t6 a_n1528_n1488# 0.065351f
C178 plus.n18 a_n1528_n1488# 0.039492f
C179 plus.t3 a_n1528_n1488# 0.065351f
C180 plus.n19 a_n1528_n1488# 0.039492f
C181 plus.n20 a_n1528_n1488# 0.011466f
C182 plus.n21 a_n1528_n1488# 0.062923f
C183 plus.n22 a_n1528_n1488# 0.030089f
C184 plus.n23 a_n1528_n1488# 0.030089f
C185 plus.n24 a_n1528_n1488# 0.010724f
C186 plus.n25 a_n1528_n1488# 0.039492f
C187 plus.n26 a_n1528_n1488# 0.011466f
C188 plus.n27 a_n1528_n1488# 0.039492f
C189 plus.n28 a_n1528_n1488# 0.047491f
C190 plus.n29 a_n1528_n1488# 0.653798f
.ends

