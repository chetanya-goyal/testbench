* NGSPICE file created from diffpair227.ext - technology: sky130A

.subckt diffpair227 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t20 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 source.t23 minus.t1 drain_right.t14 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 source.t4 plus.t0 drain_left.t15 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X3 source.t7 plus.t1 drain_left.t14 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X4 source.t18 minus.t2 drain_right.t13 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 source.t0 plus.t2 drain_left.t13 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X6 source.t13 plus.t3 drain_left.t12 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X7 source.t2 plus.t4 drain_left.t11 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X8 drain_right.t12 minus.t3 source.t17 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X9 source.t16 minus.t4 drain_right.t11 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X10 a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X11 source.t30 minus.t5 drain_right.t10 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X12 drain_left.t10 plus.t5 source.t1 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X13 source.t9 plus.t6 drain_left.t9 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X14 drain_right.t9 minus.t6 source.t22 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X15 drain_right.t8 minus.t7 source.t26 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X17 source.t28 minus.t8 drain_right.t7 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X18 drain_left.t8 plus.t7 source.t14 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X19 drain_right.t6 minus.t9 source.t21 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X20 drain_left.t7 plus.t8 source.t3 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X21 drain_right.t5 minus.t10 source.t29 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X22 drain_left.t6 plus.t9 source.t5 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 drain_left.t5 plus.t10 source.t8 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X24 drain_right.t4 minus.t11 source.t24 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X25 drain_left.t4 plus.t11 source.t10 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X26 a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X27 drain_right.t3 minus.t12 source.t19 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X28 drain_left.t3 plus.t12 source.t11 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X29 source.t12 plus.t13 drain_left.t2 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X30 source.t27 minus.t13 drain_right.t2 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X31 a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X32 drain_left.t1 plus.t14 source.t6 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X33 source.t31 minus.t14 drain_right.t1 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X34 source.t25 minus.t15 drain_right.t0 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X35 source.t15 plus.t15 drain_left.t0 a_n2570_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n7 minus.t11 183.78
R1 minus.n33 minus.t1 183.78
R2 minus.n25 minus.n24 161.3
R3 minus.n23 minus.n0 161.3
R4 minus.n22 minus.n21 161.3
R5 minus.n20 minus.n1 161.3
R6 minus.n19 minus.n18 161.3
R7 minus.n17 minus.n2 161.3
R8 minus.n16 minus.n15 161.3
R9 minus.n14 minus.n3 161.3
R10 minus.n13 minus.n12 161.3
R11 minus.n11 minus.n4 161.3
R12 minus.n10 minus.n9 161.3
R13 minus.n8 minus.n5 161.3
R14 minus.n51 minus.n50 161.3
R15 minus.n49 minus.n26 161.3
R16 minus.n48 minus.n47 161.3
R17 minus.n46 minus.n27 161.3
R18 minus.n45 minus.n44 161.3
R19 minus.n43 minus.n28 161.3
R20 minus.n42 minus.n41 161.3
R21 minus.n40 minus.n29 161.3
R22 minus.n39 minus.n38 161.3
R23 minus.n37 minus.n30 161.3
R24 minus.n36 minus.n35 161.3
R25 minus.n34 minus.n31 161.3
R26 minus.n6 minus.t2 159.405
R27 minus.n10 minus.t10 159.405
R28 minus.n12 minus.t14 159.405
R29 minus.n16 minus.t7 159.405
R30 minus.n18 minus.t15 159.405
R31 minus.n22 minus.t6 159.405
R32 minus.n24 minus.t13 159.405
R33 minus.n32 minus.t0 159.405
R34 minus.n36 minus.t4 159.405
R35 minus.n38 minus.t3 159.405
R36 minus.n42 minus.t5 159.405
R37 minus.n44 minus.t9 159.405
R38 minus.n48 minus.t8 159.405
R39 minus.n50 minus.t12 159.405
R40 minus.n8 minus.n7 44.9377
R41 minus.n34 minus.n33 44.9377
R42 minus.n24 minus.n23 37.246
R43 minus.n50 minus.n49 37.246
R44 minus.n6 minus.n5 32.8641
R45 minus.n22 minus.n1 32.8641
R46 minus.n32 minus.n31 32.8641
R47 minus.n48 minus.n27 32.8641
R48 minus.n52 minus.n25 32.1937
R49 minus.n11 minus.n10 28.4823
R50 minus.n18 minus.n17 28.4823
R51 minus.n37 minus.n36 28.4823
R52 minus.n44 minus.n43 28.4823
R53 minus.n16 minus.n3 24.1005
R54 minus.n12 minus.n3 24.1005
R55 minus.n38 minus.n29 24.1005
R56 minus.n42 minus.n29 24.1005
R57 minus.n12 minus.n11 19.7187
R58 minus.n17 minus.n16 19.7187
R59 minus.n38 minus.n37 19.7187
R60 minus.n43 minus.n42 19.7187
R61 minus.n7 minus.n6 17.0522
R62 minus.n33 minus.n32 17.0522
R63 minus.n10 minus.n5 15.3369
R64 minus.n18 minus.n1 15.3369
R65 minus.n36 minus.n31 15.3369
R66 minus.n44 minus.n27 15.3369
R67 minus.n23 minus.n22 10.955
R68 minus.n49 minus.n48 10.955
R69 minus.n52 minus.n51 6.6558
R70 minus.n25 minus.n0 0.189894
R71 minus.n21 minus.n0 0.189894
R72 minus.n21 minus.n20 0.189894
R73 minus.n20 minus.n19 0.189894
R74 minus.n19 minus.n2 0.189894
R75 minus.n15 minus.n2 0.189894
R76 minus.n15 minus.n14 0.189894
R77 minus.n14 minus.n13 0.189894
R78 minus.n13 minus.n4 0.189894
R79 minus.n9 minus.n4 0.189894
R80 minus.n9 minus.n8 0.189894
R81 minus.n35 minus.n34 0.189894
R82 minus.n35 minus.n30 0.189894
R83 minus.n39 minus.n30 0.189894
R84 minus.n40 minus.n39 0.189894
R85 minus.n41 minus.n40 0.189894
R86 minus.n41 minus.n28 0.189894
R87 minus.n45 minus.n28 0.189894
R88 minus.n46 minus.n45 0.189894
R89 minus.n47 minus.n46 0.189894
R90 minus.n47 minus.n26 0.189894
R91 minus.n51 minus.n26 0.189894
R92 minus minus.n52 0.188
R93 source.n0 source.t14 69.6943
R94 source.n7 source.t2 69.6943
R95 source.n8 source.t24 69.6943
R96 source.n15 source.t27 69.6943
R97 source.n31 source.t19 69.6942
R98 source.n24 source.t23 69.6942
R99 source.n23 source.t1 69.6942
R100 source.n16 source.t0 69.6942
R101 source.n2 source.n1 63.0943
R102 source.n4 source.n3 63.0943
R103 source.n6 source.n5 63.0943
R104 source.n10 source.n9 63.0943
R105 source.n12 source.n11 63.0943
R106 source.n14 source.n13 63.0943
R107 source.n30 source.n29 63.0942
R108 source.n28 source.n27 63.0942
R109 source.n26 source.n25 63.0942
R110 source.n22 source.n21 63.0942
R111 source.n20 source.n19 63.0942
R112 source.n18 source.n17 63.0942
R113 source.n16 source.n15 15.3575
R114 source.n32 source.n0 9.65058
R115 source.n29 source.t21 6.6005
R116 source.n29 source.t28 6.6005
R117 source.n27 source.t17 6.6005
R118 source.n27 source.t30 6.6005
R119 source.n25 source.t20 6.6005
R120 source.n25 source.t16 6.6005
R121 source.n21 source.t3 6.6005
R122 source.n21 source.t9 6.6005
R123 source.n19 source.t11 6.6005
R124 source.n19 source.t12 6.6005
R125 source.n17 source.t6 6.6005
R126 source.n17 source.t15 6.6005
R127 source.n1 source.t8 6.6005
R128 source.n1 source.t4 6.6005
R129 source.n3 source.t5 6.6005
R130 source.n3 source.t13 6.6005
R131 source.n5 source.t10 6.6005
R132 source.n5 source.t7 6.6005
R133 source.n9 source.t29 6.6005
R134 source.n9 source.t18 6.6005
R135 source.n11 source.t26 6.6005
R136 source.n11 source.t31 6.6005
R137 source.n13 source.t22 6.6005
R138 source.n13 source.t25 6.6005
R139 source.n32 source.n31 5.7074
R140 source.n15 source.n14 0.888431
R141 source.n14 source.n12 0.888431
R142 source.n12 source.n10 0.888431
R143 source.n10 source.n8 0.888431
R144 source.n7 source.n6 0.888431
R145 source.n6 source.n4 0.888431
R146 source.n4 source.n2 0.888431
R147 source.n2 source.n0 0.888431
R148 source.n18 source.n16 0.888431
R149 source.n20 source.n18 0.888431
R150 source.n22 source.n20 0.888431
R151 source.n23 source.n22 0.888431
R152 source.n26 source.n24 0.888431
R153 source.n28 source.n26 0.888431
R154 source.n30 source.n28 0.888431
R155 source.n31 source.n30 0.888431
R156 source.n8 source.n7 0.470328
R157 source.n24 source.n23 0.470328
R158 source source.n32 0.188
R159 drain_right.n9 drain_right.n7 80.661
R160 drain_right.n5 drain_right.n3 80.6609
R161 drain_right.n2 drain_right.n0 80.6609
R162 drain_right.n9 drain_right.n8 79.7731
R163 drain_right.n11 drain_right.n10 79.7731
R164 drain_right.n13 drain_right.n12 79.7731
R165 drain_right.n5 drain_right.n4 79.773
R166 drain_right.n2 drain_right.n1 79.773
R167 drain_right drain_right.n6 25.7672
R168 drain_right.n3 drain_right.t7 6.6005
R169 drain_right.n3 drain_right.t3 6.6005
R170 drain_right.n4 drain_right.t10 6.6005
R171 drain_right.n4 drain_right.t6 6.6005
R172 drain_right.n1 drain_right.t11 6.6005
R173 drain_right.n1 drain_right.t12 6.6005
R174 drain_right.n0 drain_right.t14 6.6005
R175 drain_right.n0 drain_right.t15 6.6005
R176 drain_right.n7 drain_right.t13 6.6005
R177 drain_right.n7 drain_right.t4 6.6005
R178 drain_right.n8 drain_right.t1 6.6005
R179 drain_right.n8 drain_right.t5 6.6005
R180 drain_right.n10 drain_right.t0 6.6005
R181 drain_right.n10 drain_right.t8 6.6005
R182 drain_right.n12 drain_right.t2 6.6005
R183 drain_right.n12 drain_right.t9 6.6005
R184 drain_right drain_right.n13 6.54115
R185 drain_right.n13 drain_right.n11 0.888431
R186 drain_right.n11 drain_right.n9 0.888431
R187 drain_right.n6 drain_right.n5 0.389119
R188 drain_right.n6 drain_right.n2 0.389119
R189 plus.n7 plus.t4 183.78
R190 plus.n33 plus.t5 183.78
R191 plus.n9 plus.n8 161.3
R192 plus.n10 plus.n5 161.3
R193 plus.n12 plus.n11 161.3
R194 plus.n13 plus.n4 161.3
R195 plus.n15 plus.n14 161.3
R196 plus.n16 plus.n3 161.3
R197 plus.n18 plus.n17 161.3
R198 plus.n19 plus.n2 161.3
R199 plus.n21 plus.n20 161.3
R200 plus.n22 plus.n1 161.3
R201 plus.n23 plus.n0 161.3
R202 plus.n25 plus.n24 161.3
R203 plus.n35 plus.n34 161.3
R204 plus.n36 plus.n31 161.3
R205 plus.n38 plus.n37 161.3
R206 plus.n39 plus.n30 161.3
R207 plus.n41 plus.n40 161.3
R208 plus.n42 plus.n29 161.3
R209 plus.n44 plus.n43 161.3
R210 plus.n45 plus.n28 161.3
R211 plus.n47 plus.n46 161.3
R212 plus.n48 plus.n27 161.3
R213 plus.n49 plus.n26 161.3
R214 plus.n51 plus.n50 161.3
R215 plus.n24 plus.t7 159.405
R216 plus.n22 plus.t0 159.405
R217 plus.n2 plus.t10 159.405
R218 plus.n16 plus.t3 159.405
R219 plus.n4 plus.t9 159.405
R220 plus.n10 plus.t1 159.405
R221 plus.n6 plus.t11 159.405
R222 plus.n50 plus.t2 159.405
R223 plus.n48 plus.t14 159.405
R224 plus.n28 plus.t15 159.405
R225 plus.n42 plus.t12 159.405
R226 plus.n30 plus.t13 159.405
R227 plus.n36 plus.t8 159.405
R228 plus.n32 plus.t6 159.405
R229 plus.n8 plus.n7 44.9377
R230 plus.n34 plus.n33 44.9377
R231 plus.n24 plus.n23 37.246
R232 plus.n50 plus.n49 37.246
R233 plus.n22 plus.n21 32.8641
R234 plus.n9 plus.n6 32.8641
R235 plus.n48 plus.n47 32.8641
R236 plus.n35 plus.n32 32.8641
R237 plus plus.n51 29.4839
R238 plus.n17 plus.n2 28.4823
R239 plus.n11 plus.n10 28.4823
R240 plus.n43 plus.n28 28.4823
R241 plus.n37 plus.n36 28.4823
R242 plus.n15 plus.n4 24.1005
R243 plus.n16 plus.n15 24.1005
R244 plus.n42 plus.n41 24.1005
R245 plus.n41 plus.n30 24.1005
R246 plus.n17 plus.n16 19.7187
R247 plus.n11 plus.n4 19.7187
R248 plus.n43 plus.n42 19.7187
R249 plus.n37 plus.n30 19.7187
R250 plus.n7 plus.n6 17.0522
R251 plus.n33 plus.n32 17.0522
R252 plus.n21 plus.n2 15.3369
R253 plus.n10 plus.n9 15.3369
R254 plus.n47 plus.n28 15.3369
R255 plus.n36 plus.n35 15.3369
R256 plus.n23 plus.n22 10.955
R257 plus.n49 plus.n48 10.955
R258 plus plus.n25 8.89065
R259 plus.n8 plus.n5 0.189894
R260 plus.n12 plus.n5 0.189894
R261 plus.n13 plus.n12 0.189894
R262 plus.n14 plus.n13 0.189894
R263 plus.n14 plus.n3 0.189894
R264 plus.n18 plus.n3 0.189894
R265 plus.n19 plus.n18 0.189894
R266 plus.n20 plus.n19 0.189894
R267 plus.n20 plus.n1 0.189894
R268 plus.n1 plus.n0 0.189894
R269 plus.n25 plus.n0 0.189894
R270 plus.n51 plus.n26 0.189894
R271 plus.n27 plus.n26 0.189894
R272 plus.n46 plus.n27 0.189894
R273 plus.n46 plus.n45 0.189894
R274 plus.n45 plus.n44 0.189894
R275 plus.n44 plus.n29 0.189894
R276 plus.n40 plus.n29 0.189894
R277 plus.n40 plus.n39 0.189894
R278 plus.n39 plus.n38 0.189894
R279 plus.n38 plus.n31 0.189894
R280 plus.n34 plus.n31 0.189894
R281 drain_left.n9 drain_left.n7 80.661
R282 drain_left.n5 drain_left.n3 80.6609
R283 drain_left.n2 drain_left.n0 80.6609
R284 drain_left.n13 drain_left.n12 79.7731
R285 drain_left.n11 drain_left.n10 79.7731
R286 drain_left.n9 drain_left.n8 79.7731
R287 drain_left.n5 drain_left.n4 79.773
R288 drain_left.n2 drain_left.n1 79.773
R289 drain_left drain_left.n6 26.3204
R290 drain_left.n3 drain_left.t9 6.6005
R291 drain_left.n3 drain_left.t10 6.6005
R292 drain_left.n4 drain_left.t2 6.6005
R293 drain_left.n4 drain_left.t7 6.6005
R294 drain_left.n1 drain_left.t0 6.6005
R295 drain_left.n1 drain_left.t3 6.6005
R296 drain_left.n0 drain_left.t13 6.6005
R297 drain_left.n0 drain_left.t1 6.6005
R298 drain_left.n12 drain_left.t15 6.6005
R299 drain_left.n12 drain_left.t8 6.6005
R300 drain_left.n10 drain_left.t12 6.6005
R301 drain_left.n10 drain_left.t5 6.6005
R302 drain_left.n8 drain_left.t14 6.6005
R303 drain_left.n8 drain_left.t6 6.6005
R304 drain_left.n7 drain_left.t11 6.6005
R305 drain_left.n7 drain_left.t4 6.6005
R306 drain_left drain_left.n13 6.54115
R307 drain_left.n11 drain_left.n9 0.888431
R308 drain_left.n13 drain_left.n11 0.888431
R309 drain_left.n6 drain_left.n5 0.389119
R310 drain_left.n6 drain_left.n2 0.389119
C0 source drain_left 7.54678f
C1 source drain_right 7.549029f
C2 minus drain_left 0.17772f
C3 minus drain_right 3.00649f
C4 drain_left drain_right 1.34352f
C5 source plus 3.53182f
C6 minus plus 4.6902f
C7 minus source 3.51782f
C8 plus drain_left 3.26107f
C9 plus drain_right 0.416359f
C10 drain_right a_n2570_n1488# 5.01699f
C11 drain_left a_n2570_n1488# 5.40332f
C12 source a_n2570_n1488# 3.950219f
C13 minus a_n2570_n1488# 9.502752f
C14 plus a_n2570_n1488# 10.842971f
C15 drain_left.t13 a_n2570_n1488# 0.064255f
C16 drain_left.t1 a_n2570_n1488# 0.064255f
C17 drain_left.n0 a_n2570_n1488# 0.467619f
C18 drain_left.t0 a_n2570_n1488# 0.064255f
C19 drain_left.t3 a_n2570_n1488# 0.064255f
C20 drain_left.n1 a_n2570_n1488# 0.463404f
C21 drain_left.n2 a_n2570_n1488# 0.70883f
C22 drain_left.t9 a_n2570_n1488# 0.064255f
C23 drain_left.t10 a_n2570_n1488# 0.064255f
C24 drain_left.n3 a_n2570_n1488# 0.467619f
C25 drain_left.t2 a_n2570_n1488# 0.064255f
C26 drain_left.t7 a_n2570_n1488# 0.064255f
C27 drain_left.n4 a_n2570_n1488# 0.463404f
C28 drain_left.n5 a_n2570_n1488# 0.70883f
C29 drain_left.n6 a_n2570_n1488# 1.04157f
C30 drain_left.t11 a_n2570_n1488# 0.064255f
C31 drain_left.t4 a_n2570_n1488# 0.064255f
C32 drain_left.n7 a_n2570_n1488# 0.467622f
C33 drain_left.t14 a_n2570_n1488# 0.064255f
C34 drain_left.t6 a_n2570_n1488# 0.064255f
C35 drain_left.n8 a_n2570_n1488# 0.463406f
C36 drain_left.n9 a_n2570_n1488# 0.750816f
C37 drain_left.t12 a_n2570_n1488# 0.064255f
C38 drain_left.t5 a_n2570_n1488# 0.064255f
C39 drain_left.n10 a_n2570_n1488# 0.463406f
C40 drain_left.n11 a_n2570_n1488# 0.372058f
C41 drain_left.t15 a_n2570_n1488# 0.064255f
C42 drain_left.t8 a_n2570_n1488# 0.064255f
C43 drain_left.n12 a_n2570_n1488# 0.463406f
C44 drain_left.n13 a_n2570_n1488# 0.611795f
C45 plus.n0 a_n2570_n1488# 0.043904f
C46 plus.t7 a_n2570_n1488# 0.276469f
C47 plus.t0 a_n2570_n1488# 0.276469f
C48 plus.n1 a_n2570_n1488# 0.043904f
C49 plus.t10 a_n2570_n1488# 0.276469f
C50 plus.n2 a_n2570_n1488# 0.161022f
C51 plus.n3 a_n2570_n1488# 0.043904f
C52 plus.t3 a_n2570_n1488# 0.276469f
C53 plus.t9 a_n2570_n1488# 0.276469f
C54 plus.n4 a_n2570_n1488# 0.161022f
C55 plus.n5 a_n2570_n1488# 0.043904f
C56 plus.t1 a_n2570_n1488# 0.276469f
C57 plus.t11 a_n2570_n1488# 0.276469f
C58 plus.n6 a_n2570_n1488# 0.167037f
C59 plus.t4 a_n2570_n1488# 0.297849f
C60 plus.n7 a_n2570_n1488# 0.143296f
C61 plus.n8 a_n2570_n1488# 0.185791f
C62 plus.n9 a_n2570_n1488# 0.009963f
C63 plus.n10 a_n2570_n1488# 0.161022f
C64 plus.n11 a_n2570_n1488# 0.009963f
C65 plus.n12 a_n2570_n1488# 0.043904f
C66 plus.n13 a_n2570_n1488# 0.043904f
C67 plus.n14 a_n2570_n1488# 0.043904f
C68 plus.n15 a_n2570_n1488# 0.009963f
C69 plus.n16 a_n2570_n1488# 0.161022f
C70 plus.n17 a_n2570_n1488# 0.009963f
C71 plus.n18 a_n2570_n1488# 0.043904f
C72 plus.n19 a_n2570_n1488# 0.043904f
C73 plus.n20 a_n2570_n1488# 0.043904f
C74 plus.n21 a_n2570_n1488# 0.009963f
C75 plus.n22 a_n2570_n1488# 0.161022f
C76 plus.n23 a_n2570_n1488# 0.009963f
C77 plus.n24 a_n2570_n1488# 0.159804f
C78 plus.n25 a_n2570_n1488# 0.344815f
C79 plus.n26 a_n2570_n1488# 0.043904f
C80 plus.t2 a_n2570_n1488# 0.276469f
C81 plus.n27 a_n2570_n1488# 0.043904f
C82 plus.t14 a_n2570_n1488# 0.276469f
C83 plus.t15 a_n2570_n1488# 0.276469f
C84 plus.n28 a_n2570_n1488# 0.161022f
C85 plus.n29 a_n2570_n1488# 0.043904f
C86 plus.t12 a_n2570_n1488# 0.276469f
C87 plus.t13 a_n2570_n1488# 0.276469f
C88 plus.n30 a_n2570_n1488# 0.161022f
C89 plus.n31 a_n2570_n1488# 0.043904f
C90 plus.t8 a_n2570_n1488# 0.276469f
C91 plus.t6 a_n2570_n1488# 0.276469f
C92 plus.n32 a_n2570_n1488# 0.167037f
C93 plus.t5 a_n2570_n1488# 0.297849f
C94 plus.n33 a_n2570_n1488# 0.143296f
C95 plus.n34 a_n2570_n1488# 0.185791f
C96 plus.n35 a_n2570_n1488# 0.009963f
C97 plus.n36 a_n2570_n1488# 0.161022f
C98 plus.n37 a_n2570_n1488# 0.009963f
C99 plus.n38 a_n2570_n1488# 0.043904f
C100 plus.n39 a_n2570_n1488# 0.043904f
C101 plus.n40 a_n2570_n1488# 0.043904f
C102 plus.n41 a_n2570_n1488# 0.009963f
C103 plus.n42 a_n2570_n1488# 0.161022f
C104 plus.n43 a_n2570_n1488# 0.009963f
C105 plus.n44 a_n2570_n1488# 0.043904f
C106 plus.n45 a_n2570_n1488# 0.043904f
C107 plus.n46 a_n2570_n1488# 0.043904f
C108 plus.n47 a_n2570_n1488# 0.009963f
C109 plus.n48 a_n2570_n1488# 0.161022f
C110 plus.n49 a_n2570_n1488# 0.009963f
C111 plus.n50 a_n2570_n1488# 0.159804f
C112 plus.n51 a_n2570_n1488# 1.2128f
C113 drain_right.t14 a_n2570_n1488# 0.06309f
C114 drain_right.t15 a_n2570_n1488# 0.06309f
C115 drain_right.n0 a_n2570_n1488# 0.459137f
C116 drain_right.t11 a_n2570_n1488# 0.06309f
C117 drain_right.t12 a_n2570_n1488# 0.06309f
C118 drain_right.n1 a_n2570_n1488# 0.454998f
C119 drain_right.n2 a_n2570_n1488# 0.695973f
C120 drain_right.t7 a_n2570_n1488# 0.06309f
C121 drain_right.t3 a_n2570_n1488# 0.06309f
C122 drain_right.n3 a_n2570_n1488# 0.459137f
C123 drain_right.t10 a_n2570_n1488# 0.06309f
C124 drain_right.t6 a_n2570_n1488# 0.06309f
C125 drain_right.n4 a_n2570_n1488# 0.454998f
C126 drain_right.n5 a_n2570_n1488# 0.695973f
C127 drain_right.n6 a_n2570_n1488# 0.97039f
C128 drain_right.t13 a_n2570_n1488# 0.06309f
C129 drain_right.t4 a_n2570_n1488# 0.06309f
C130 drain_right.n7 a_n2570_n1488# 0.45914f
C131 drain_right.t1 a_n2570_n1488# 0.06309f
C132 drain_right.t5 a_n2570_n1488# 0.06309f
C133 drain_right.n8 a_n2570_n1488# 0.455f
C134 drain_right.n9 a_n2570_n1488# 0.737198f
C135 drain_right.t0 a_n2570_n1488# 0.06309f
C136 drain_right.t8 a_n2570_n1488# 0.06309f
C137 drain_right.n10 a_n2570_n1488# 0.455f
C138 drain_right.n11 a_n2570_n1488# 0.365309f
C139 drain_right.t2 a_n2570_n1488# 0.06309f
C140 drain_right.t9 a_n2570_n1488# 0.06309f
C141 drain_right.n12 a_n2570_n1488# 0.455f
C142 drain_right.n13 a_n2570_n1488# 0.600698f
C143 source.t14 a_n2570_n1488# 0.549629f
C144 source.n0 a_n2570_n1488# 0.804369f
C145 source.t8 a_n2570_n1488# 0.06619f
C146 source.t4 a_n2570_n1488# 0.06619f
C147 source.n1 a_n2570_n1488# 0.419682f
C148 source.n2 a_n2570_n1488# 0.402984f
C149 source.t5 a_n2570_n1488# 0.06619f
C150 source.t13 a_n2570_n1488# 0.06619f
C151 source.n3 a_n2570_n1488# 0.419682f
C152 source.n4 a_n2570_n1488# 0.402984f
C153 source.t10 a_n2570_n1488# 0.06619f
C154 source.t7 a_n2570_n1488# 0.06619f
C155 source.n5 a_n2570_n1488# 0.419682f
C156 source.n6 a_n2570_n1488# 0.402984f
C157 source.t2 a_n2570_n1488# 0.549629f
C158 source.n7 a_n2570_n1488# 0.415941f
C159 source.t24 a_n2570_n1488# 0.549629f
C160 source.n8 a_n2570_n1488# 0.415941f
C161 source.t29 a_n2570_n1488# 0.06619f
C162 source.t18 a_n2570_n1488# 0.06619f
C163 source.n9 a_n2570_n1488# 0.419682f
C164 source.n10 a_n2570_n1488# 0.402984f
C165 source.t26 a_n2570_n1488# 0.06619f
C166 source.t31 a_n2570_n1488# 0.06619f
C167 source.n11 a_n2570_n1488# 0.419682f
C168 source.n12 a_n2570_n1488# 0.402984f
C169 source.t22 a_n2570_n1488# 0.06619f
C170 source.t25 a_n2570_n1488# 0.06619f
C171 source.n13 a_n2570_n1488# 0.419682f
C172 source.n14 a_n2570_n1488# 0.402984f
C173 source.t27 a_n2570_n1488# 0.549629f
C174 source.n15 a_n2570_n1488# 1.10295f
C175 source.t0 a_n2570_n1488# 0.549626f
C176 source.n16 a_n2570_n1488# 1.10295f
C177 source.t6 a_n2570_n1488# 0.06619f
C178 source.t15 a_n2570_n1488# 0.06619f
C179 source.n17 a_n2570_n1488# 0.419678f
C180 source.n18 a_n2570_n1488# 0.402987f
C181 source.t11 a_n2570_n1488# 0.06619f
C182 source.t12 a_n2570_n1488# 0.06619f
C183 source.n19 a_n2570_n1488# 0.419678f
C184 source.n20 a_n2570_n1488# 0.402987f
C185 source.t3 a_n2570_n1488# 0.06619f
C186 source.t9 a_n2570_n1488# 0.06619f
C187 source.n21 a_n2570_n1488# 0.419678f
C188 source.n22 a_n2570_n1488# 0.402987f
C189 source.t1 a_n2570_n1488# 0.549626f
C190 source.n23 a_n2570_n1488# 0.415943f
C191 source.t23 a_n2570_n1488# 0.549626f
C192 source.n24 a_n2570_n1488# 0.415943f
C193 source.t20 a_n2570_n1488# 0.06619f
C194 source.t16 a_n2570_n1488# 0.06619f
C195 source.n25 a_n2570_n1488# 0.419678f
C196 source.n26 a_n2570_n1488# 0.402987f
C197 source.t17 a_n2570_n1488# 0.06619f
C198 source.t30 a_n2570_n1488# 0.06619f
C199 source.n27 a_n2570_n1488# 0.419678f
C200 source.n28 a_n2570_n1488# 0.402987f
C201 source.t21 a_n2570_n1488# 0.06619f
C202 source.t28 a_n2570_n1488# 0.06619f
C203 source.n29 a_n2570_n1488# 0.419678f
C204 source.n30 a_n2570_n1488# 0.402987f
C205 source.t19 a_n2570_n1488# 0.549626f
C206 source.n31 a_n2570_n1488# 0.598067f
C207 source.n32 a_n2570_n1488# 0.823327f
C208 minus.n0 a_n2570_n1488# 0.042431f
C209 minus.n1 a_n2570_n1488# 0.009628f
C210 minus.t6 a_n2570_n1488# 0.267194f
C211 minus.n2 a_n2570_n1488# 0.042431f
C212 minus.n3 a_n2570_n1488# 0.009628f
C213 minus.t7 a_n2570_n1488# 0.267194f
C214 minus.n4 a_n2570_n1488# 0.042431f
C215 minus.n5 a_n2570_n1488# 0.009628f
C216 minus.t10 a_n2570_n1488# 0.267194f
C217 minus.t11 a_n2570_n1488# 0.287857f
C218 minus.t2 a_n2570_n1488# 0.267194f
C219 minus.n6 a_n2570_n1488# 0.161433f
C220 minus.n7 a_n2570_n1488# 0.138489f
C221 minus.n8 a_n2570_n1488# 0.179558f
C222 minus.n9 a_n2570_n1488# 0.042431f
C223 minus.n10 a_n2570_n1488# 0.15562f
C224 minus.n11 a_n2570_n1488# 0.009628f
C225 minus.t14 a_n2570_n1488# 0.267194f
C226 minus.n12 a_n2570_n1488# 0.15562f
C227 minus.n13 a_n2570_n1488# 0.042431f
C228 minus.n14 a_n2570_n1488# 0.042431f
C229 minus.n15 a_n2570_n1488# 0.042431f
C230 minus.n16 a_n2570_n1488# 0.15562f
C231 minus.n17 a_n2570_n1488# 0.009628f
C232 minus.t15 a_n2570_n1488# 0.267194f
C233 minus.n18 a_n2570_n1488# 0.15562f
C234 minus.n19 a_n2570_n1488# 0.042431f
C235 minus.n20 a_n2570_n1488# 0.042431f
C236 minus.n21 a_n2570_n1488# 0.042431f
C237 minus.n22 a_n2570_n1488# 0.15562f
C238 minus.n23 a_n2570_n1488# 0.009628f
C239 minus.t13 a_n2570_n1488# 0.267194f
C240 minus.n24 a_n2570_n1488# 0.154443f
C241 minus.n25 a_n2570_n1488# 1.2483f
C242 minus.n26 a_n2570_n1488# 0.042431f
C243 minus.n27 a_n2570_n1488# 0.009628f
C244 minus.n28 a_n2570_n1488# 0.042431f
C245 minus.n29 a_n2570_n1488# 0.009628f
C246 minus.n30 a_n2570_n1488# 0.042431f
C247 minus.n31 a_n2570_n1488# 0.009628f
C248 minus.t1 a_n2570_n1488# 0.287857f
C249 minus.t0 a_n2570_n1488# 0.267194f
C250 minus.n32 a_n2570_n1488# 0.161433f
C251 minus.n33 a_n2570_n1488# 0.138489f
C252 minus.n34 a_n2570_n1488# 0.179558f
C253 minus.n35 a_n2570_n1488# 0.042431f
C254 minus.t4 a_n2570_n1488# 0.267194f
C255 minus.n36 a_n2570_n1488# 0.15562f
C256 minus.n37 a_n2570_n1488# 0.009628f
C257 minus.t3 a_n2570_n1488# 0.267194f
C258 minus.n38 a_n2570_n1488# 0.15562f
C259 minus.n39 a_n2570_n1488# 0.042431f
C260 minus.n40 a_n2570_n1488# 0.042431f
C261 minus.n41 a_n2570_n1488# 0.042431f
C262 minus.t5 a_n2570_n1488# 0.267194f
C263 minus.n42 a_n2570_n1488# 0.15562f
C264 minus.n43 a_n2570_n1488# 0.009628f
C265 minus.t9 a_n2570_n1488# 0.267194f
C266 minus.n44 a_n2570_n1488# 0.15562f
C267 minus.n45 a_n2570_n1488# 0.042431f
C268 minus.n46 a_n2570_n1488# 0.042431f
C269 minus.n47 a_n2570_n1488# 0.042431f
C270 minus.t8 a_n2570_n1488# 0.267194f
C271 minus.n48 a_n2570_n1488# 0.15562f
C272 minus.n49 a_n2570_n1488# 0.009628f
C273 minus.t12 a_n2570_n1488# 0.267194f
C274 minus.n50 a_n2570_n1488# 0.154443f
C275 minus.n51 a_n2570_n1488# 0.292865f
C276 minus.n52 a_n2570_n1488# 1.52633f
.ends

