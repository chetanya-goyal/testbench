* NGSPICE file created from diffpair401.ext - technology: sky130A

.subckt diffpair401 minus drain_right drain_left source plus
X0 drain_right minus source a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X1 drain_right minus source a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X2 source plus drain_left a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X3 a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X4 source plus drain_left a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X5 drain_left plus source a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X6 source minus drain_right a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X7 a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X8 a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X9 a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X10 drain_left plus source a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X11 source minus drain_right a_n1106_n3292# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
.ends

