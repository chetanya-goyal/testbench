* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t9 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X1 drain_right.t4 minus.t1 source.t8 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X2 drain_left.t5 plus.t0 source.t3 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X3 source.t2 plus.t1 drain_left.t4 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X4 source.t10 minus.t2 drain_right.t3 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X5 a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.2
X6 drain_left.t3 plus.t2 source.t0 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X7 drain_right.t2 minus.t3 source.t6 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X8 a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X9 drain_left.t2 plus.t3 source.t5 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X10 a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X11 drain_right.t1 minus.t4 source.t7 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X12 source.t11 minus.t5 drain_right.t0 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X13 source.t1 plus.t4 drain_left.t1 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X14 a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X15 drain_left.t0 plus.t5 source.t4 a_n1140_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
R0 minus.n2 minus.t0 318.048
R1 minus.n0 minus.t4 318.048
R2 minus.n6 minus.t1 318.048
R3 minus.n4 minus.t3 318.048
R4 minus.n1 minus.t2 277.151
R5 minus.n5 minus.t5 277.151
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 25.0441
R15 minus.n8 minus.n7 6.438
R16 minus minus.n8 0.188
R17 source.n0 source.t4 243.255
R18 source.n3 source.t7 243.255
R19 source.n11 source.t8 243.254
R20 source.n8 source.t5 243.254
R21 source.n2 source.n1 223.454
R22 source.n5 source.n4 223.454
R23 source.n10 source.n9 223.453
R24 source.n7 source.n6 223.453
R25 source.n9 source.t6 19.8005
R26 source.n9 source.t11 19.8005
R27 source.n6 source.t3 19.8005
R28 source.n6 source.t1 19.8005
R29 source.n1 source.t0 19.8005
R30 source.n1 source.t2 19.8005
R31 source.n4 source.t9 19.8005
R32 source.n4 source.t10 19.8005
R33 source.n7 source.n5 13.8682
R34 source.n12 source.n0 7.91991
R35 source.n12 source.n11 5.49188
R36 source.n3 source.n2 0.698776
R37 source.n10 source.n8 0.698776
R38 source.n5 source.n3 0.457397
R39 source.n2 source.n0 0.457397
R40 source.n8 source.n7 0.457397
R41 source.n11 source.n10 0.457397
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t2 260.219
R44 drain_right.n3 drain_right.t5 259.933
R45 drain_right.n3 drain_right.n2 240.589
R46 drain_right.n1 drain_right.n0 240.19
R47 drain_right.n0 drain_right.t0 19.8005
R48 drain_right.n0 drain_right.t4 19.8005
R49 drain_right.n2 drain_right.t3 19.8005
R50 drain_right.n2 drain_right.t1 19.8005
R51 drain_right drain_right.n1 19.737
R52 drain_right drain_right.n3 5.88166
R53 plus.n0 plus.t2 318.048
R54 plus.n2 plus.t5 318.048
R55 plus.n4 plus.t3 318.048
R56 plus.n6 plus.t0 318.048
R57 plus.n1 plus.t1 277.151
R58 plus.n5 plus.t4 277.151
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 23.0918
R68 plus plus.n3 7.91527
R69 drain_left.n3 drain_left.t3 260.389
R70 drain_left.n1 drain_left.t5 260.219
R71 drain_left.n1 drain_left.n0 240.19
R72 drain_left.n3 drain_left.n2 240.132
R73 drain_left drain_left.n1 20.2902
R74 drain_left.n0 drain_left.t1 19.8005
R75 drain_left.n0 drain_left.t2 19.8005
R76 drain_left.n2 drain_left.t4 19.8005
R77 drain_left.n2 drain_left.t0 19.8005
R78 drain_left drain_left.n3 6.11011
C0 drain_left source 2.83381f
C1 drain_right plus 0.267611f
C2 minus drain_left 0.177937f
C3 source plus 0.566968f
C4 minus plus 2.54817f
C5 source drain_right 2.83036f
C6 minus drain_right 0.461065f
C7 minus source 0.553046f
C8 drain_left plus 0.566637f
C9 drain_left drain_right 0.530412f
C10 drain_right a_n1140_n1088# 2.716167f
C11 drain_left a_n1140_n1088# 2.85691f
C12 source a_n1140_n1088# 1.88208f
C13 minus a_n1140_n1088# 3.483217f
C14 plus a_n1140_n1088# 4.237042f
C15 drain_left.t5 a_n1140_n1088# 0.107665f
C16 drain_left.t1 a_n1140_n1088# 0.017372f
C17 drain_left.t2 a_n1140_n1088# 0.017372f
C18 drain_left.n0 a_n1140_n1088# 0.067553f
C19 drain_left.n1 a_n1140_n1088# 0.831393f
C20 drain_left.t3 a_n1140_n1088# 0.107808f
C21 drain_left.t4 a_n1140_n1088# 0.017372f
C22 drain_left.t0 a_n1140_n1088# 0.017372f
C23 drain_left.n2 a_n1140_n1088# 0.067503f
C24 drain_left.n3 a_n1140_n1088# 0.6004f
C25 plus.t2 a_n1140_n1088# 0.03021f
C26 plus.n0 a_n1140_n1088# 0.041874f
C27 plus.t1 a_n1140_n1088# 0.026239f
C28 plus.n1 a_n1140_n1088# 0.031407f
C29 plus.t5 a_n1140_n1088# 0.03021f
C30 plus.n2 a_n1140_n1088# 0.041816f
C31 plus.n3 a_n1140_n1088# 0.334529f
C32 plus.t3 a_n1140_n1088# 0.03021f
C33 plus.n4 a_n1140_n1088# 0.041874f
C34 plus.t0 a_n1140_n1088# 0.03021f
C35 plus.t4 a_n1140_n1088# 0.026239f
C36 plus.n5 a_n1140_n1088# 0.031407f
C37 plus.n6 a_n1140_n1088# 0.041816f
C38 plus.n7 a_n1140_n1088# 0.83227f
C39 drain_right.t2 a_n1140_n1088# 0.111077f
C40 drain_right.t0 a_n1140_n1088# 0.017923f
C41 drain_right.t4 a_n1140_n1088# 0.017923f
C42 drain_right.n0 a_n1140_n1088# 0.069694f
C43 drain_right.n1 a_n1140_n1088# 0.813704f
C44 drain_right.t3 a_n1140_n1088# 0.017923f
C45 drain_right.t1 a_n1140_n1088# 0.017923f
C46 drain_right.n2 a_n1140_n1088# 0.070087f
C47 drain_right.t5 a_n1140_n1088# 0.110858f
C48 drain_right.n3 a_n1140_n1088# 0.627204f
C49 source.t4 a_n1140_n1088# 0.133619f
C50 source.n0 a_n1140_n1088# 0.558605f
C51 source.t0 a_n1140_n1088# 0.024007f
C52 source.t2 a_n1140_n1088# 0.024007f
C53 source.n1 a_n1140_n1088# 0.077859f
C54 source.n2 a_n1140_n1088# 0.299662f
C55 source.t7 a_n1140_n1088# 0.133619f
C56 source.n3 a_n1140_n1088# 0.309375f
C57 source.t9 a_n1140_n1088# 0.024007f
C58 source.t10 a_n1140_n1088# 0.024007f
C59 source.n4 a_n1140_n1088# 0.077859f
C60 source.n5 a_n1140_n1088# 0.835309f
C61 source.t3 a_n1140_n1088# 0.024007f
C62 source.t1 a_n1140_n1088# 0.024007f
C63 source.n6 a_n1140_n1088# 0.077858f
C64 source.n7 a_n1140_n1088# 0.835309f
C65 source.t5 a_n1140_n1088# 0.133619f
C66 source.n8 a_n1140_n1088# 0.309375f
C67 source.t6 a_n1140_n1088# 0.024007f
C68 source.t11 a_n1140_n1088# 0.024007f
C69 source.n9 a_n1140_n1088# 0.077858f
C70 source.n10 a_n1140_n1088# 0.299662f
C71 source.t8 a_n1140_n1088# 0.133619f
C72 source.n11 a_n1140_n1088# 0.451741f
C73 source.n12 a_n1140_n1088# 0.611855f
C74 minus.t4 a_n1140_n1088# 0.029204f
C75 minus.n0 a_n1140_n1088# 0.04048f
C76 minus.t0 a_n1140_n1088# 0.029204f
C77 minus.t2 a_n1140_n1088# 0.025365f
C78 minus.n1 a_n1140_n1088# 0.030362f
C79 minus.n2 a_n1140_n1088# 0.040424f
C80 minus.n3 a_n1140_n1088# 0.819124f
C81 minus.t3 a_n1140_n1088# 0.029204f
C82 minus.n4 a_n1140_n1088# 0.04048f
C83 minus.t5 a_n1140_n1088# 0.025365f
C84 minus.n5 a_n1140_n1088# 0.030362f
C85 minus.t1 a_n1140_n1088# 0.029204f
C86 minus.n6 a_n1140_n1088# 0.040424f
C87 minus.n7 a_n1140_n1088# 0.310625f
C88 minus.n8 a_n1140_n1088# 0.953154f
.ends

