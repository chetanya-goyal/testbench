* NGSPICE file created from diffpair358.ext - technology: sky130A

.subckt diffpair358 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t30 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X1 source.t5 minus.t0 drain_right.t19 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 drain_left.t18 plus.t1 source.t32 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X3 drain_left.t17 plus.t2 source.t21 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 drain_right.t18 minus.t1 source.t9 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X5 drain_right.t17 minus.t2 source.t10 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X6 source.t33 plus.t3 drain_left.t16 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X7 source.t14 minus.t3 drain_right.t16 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X8 source.t1 minus.t4 drain_right.t15 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X10 drain_right.t14 minus.t5 source.t2 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 source.t39 minus.t6 drain_right.t13 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X12 source.t26 plus.t4 drain_left.t15 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X13 a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X14 source.t36 plus.t5 drain_left.t14 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 source.t27 plus.t6 drain_left.t13 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X16 source.t24 plus.t7 drain_left.t12 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X17 a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X18 drain_left.t11 plus.t8 source.t20 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X19 drain_right.t12 minus.t7 source.t4 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X20 drain_right.t11 minus.t8 source.t0 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X21 source.t3 minus.t9 drain_right.t10 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X22 source.t13 minus.t10 drain_right.t9 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X23 a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X24 source.t28 plus.t9 drain_left.t10 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X25 drain_right.t8 minus.t11 source.t11 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X26 drain_right.t7 minus.t12 source.t15 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X27 source.t37 plus.t10 drain_left.t9 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X28 source.t35 plus.t11 drain_left.t8 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X29 drain_right.t6 minus.t13 source.t38 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X30 drain_left.t7 plus.t12 source.t31 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X31 drain_left.t6 plus.t13 source.t22 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X32 source.t29 plus.t14 drain_left.t5 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X33 drain_left.t4 plus.t15 source.t23 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X34 drain_left.t3 plus.t16 source.t19 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X35 drain_right.t5 minus.t14 source.t12 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X36 source.t6 minus.t15 drain_right.t4 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X37 source.t7 minus.t16 drain_right.t3 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X38 source.t17 minus.t17 drain_right.t2 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X39 source.t16 minus.t18 drain_right.t1 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X40 source.t18 plus.t17 drain_left.t2 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X41 drain_right.t0 minus.t19 source.t8 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X42 drain_left.t1 plus.t18 source.t34 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X43 drain_left.t0 plus.t19 source.t25 a_n2102_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 plus.n6 plus.t3 876.365
R1 plus.n27 plus.t16 876.365
R2 plus.n36 plus.t13 876.365
R3 plus.n56 plus.t11 876.365
R4 plus.n5 plus.t8 827.433
R5 plus.n9 plus.t14 827.433
R6 plus.n3 plus.t18 827.433
R7 plus.n15 plus.t5 827.433
R8 plus.n17 plus.t12 827.433
R9 plus.n18 plus.t17 827.433
R10 plus.n24 plus.t0 827.433
R11 plus.n26 plus.t9 827.433
R12 plus.n35 plus.t4 827.433
R13 plus.n39 plus.t15 827.433
R14 plus.n33 plus.t6 827.433
R15 plus.n45 plus.t1 827.433
R16 plus.n47 plus.t7 827.433
R17 plus.n32 plus.t2 827.433
R18 plus.n53 plus.t10 827.433
R19 plus.n55 plus.t19 827.433
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 64.9975
R47 plus.n19 plus.n18 64.9975
R48 plus.n48 plus.n32 64.9975
R49 plus.n44 plus.n33 64.9975
R50 plus.n9 plus.n8 62.0763
R51 plus.n25 plus.n24 62.0763
R52 plus.n54 plus.n53 62.0763
R53 plus.n39 plus.n38 62.0763
R54 plus.n16 plus.n15 46.0096
R55 plus.n17 plus.n16 46.0096
R56 plus.n47 plus.n46 46.0096
R57 plus.n46 plus.n45 46.0096
R58 plus.n6 plus.n5 43.0884
R59 plus.n27 plus.n26 43.0884
R60 plus.n56 plus.n55 43.0884
R61 plus.n36 plus.n35 43.0884
R62 plus.n8 plus.n5 29.9429
R63 plus.n26 plus.n25 29.9429
R64 plus.n55 plus.n54 29.9429
R65 plus.n38 plus.n35 29.9429
R66 plus plus.n57 29.8437
R67 plus.n15 plus.n14 27.0217
R68 plus.n19 plus.n17 27.0217
R69 plus.n48 plus.n47 27.0217
R70 plus.n45 plus.n44 27.0217
R71 plus plus.n28 11.0232
R72 plus.n10 plus.n9 10.955
R73 plus.n24 plus.n23 10.955
R74 plus.n53 plus.n52 10.955
R75 plus.n40 plus.n39 10.955
R76 plus.n11 plus.n3 8.03383
R77 plus.n18 plus.n1 8.03383
R78 plus.n32 plus.n30 8.03383
R79 plus.n41 plus.n33 8.03383
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n9 source.t33 51.0588
R99 source.n10 source.t38 51.0588
R100 source.n19 source.t39 51.0588
R101 source.n39 source.t8 51.0586
R102 source.n30 source.t16 51.0586
R103 source.n29 source.t22 51.0586
R104 source.n20 source.t35 51.0586
R105 source.n0 source.t19 51.0586
R106 source.n2 source.n1 48.8588
R107 source.n4 source.n3 48.8588
R108 source.n6 source.n5 48.8588
R109 source.n8 source.n7 48.8588
R110 source.n12 source.n11 48.8588
R111 source.n14 source.n13 48.8588
R112 source.n16 source.n15 48.8588
R113 source.n18 source.n17 48.8588
R114 source.n38 source.n37 48.8586
R115 source.n36 source.n35 48.8586
R116 source.n34 source.n33 48.8586
R117 source.n32 source.n31 48.8586
R118 source.n28 source.n27 48.8586
R119 source.n26 source.n25 48.8586
R120 source.n24 source.n23 48.8586
R121 source.n22 source.n21 48.8586
R122 source.n20 source.n19 19.5581
R123 source.n40 source.n0 14.0236
R124 source.n40 source.n39 5.53498
R125 source.n37 source.t11 2.2005
R126 source.n37 source.t13 2.2005
R127 source.n35 source.t15 2.2005
R128 source.n35 source.t14 2.2005
R129 source.n33 source.t4 2.2005
R130 source.n33 source.t1 2.2005
R131 source.n31 source.t0 2.2005
R132 source.n31 source.t17 2.2005
R133 source.n27 source.t23 2.2005
R134 source.n27 source.t26 2.2005
R135 source.n25 source.t32 2.2005
R136 source.n25 source.t27 2.2005
R137 source.n23 source.t21 2.2005
R138 source.n23 source.t24 2.2005
R139 source.n21 source.t25 2.2005
R140 source.n21 source.t37 2.2005
R141 source.n1 source.t30 2.2005
R142 source.n1 source.t28 2.2005
R143 source.n3 source.t31 2.2005
R144 source.n3 source.t18 2.2005
R145 source.n5 source.t34 2.2005
R146 source.n5 source.t36 2.2005
R147 source.n7 source.t20 2.2005
R148 source.n7 source.t29 2.2005
R149 source.n11 source.t9 2.2005
R150 source.n11 source.t6 2.2005
R151 source.n13 source.t12 2.2005
R152 source.n13 source.t3 2.2005
R153 source.n15 source.t2 2.2005
R154 source.n15 source.t5 2.2005
R155 source.n17 source.t10 2.2005
R156 source.n17 source.t7 2.2005
R157 source.n19 source.n18 0.543603
R158 source.n18 source.n16 0.543603
R159 source.n16 source.n14 0.543603
R160 source.n14 source.n12 0.543603
R161 source.n12 source.n10 0.543603
R162 source.n9 source.n8 0.543603
R163 source.n8 source.n6 0.543603
R164 source.n6 source.n4 0.543603
R165 source.n4 source.n2 0.543603
R166 source.n2 source.n0 0.543603
R167 source.n22 source.n20 0.543603
R168 source.n24 source.n22 0.543603
R169 source.n26 source.n24 0.543603
R170 source.n28 source.n26 0.543603
R171 source.n29 source.n28 0.543603
R172 source.n32 source.n30 0.543603
R173 source.n34 source.n32 0.543603
R174 source.n36 source.n34 0.543603
R175 source.n38 source.n36 0.543603
R176 source.n39 source.n38 0.543603
R177 source.n10 source.n9 0.470328
R178 source.n30 source.n29 0.470328
R179 source source.n40 0.188
R180 drain_left.n10 drain_left.n8 66.0807
R181 drain_left.n6 drain_left.n4 66.0804
R182 drain_left.n2 drain_left.n0 66.0804
R183 drain_left.n14 drain_left.n13 65.5376
R184 drain_left.n12 drain_left.n11 65.5376
R185 drain_left.n10 drain_left.n9 65.5376
R186 drain_left.n16 drain_left.n15 65.5374
R187 drain_left.n7 drain_left.n3 65.5373
R188 drain_left.n6 drain_left.n5 65.5373
R189 drain_left.n2 drain_left.n1 65.5373
R190 drain_left drain_left.n7 29.4392
R191 drain_left drain_left.n16 6.19632
R192 drain_left.n3 drain_left.t12 2.2005
R193 drain_left.n3 drain_left.t18 2.2005
R194 drain_left.n4 drain_left.t15 2.2005
R195 drain_left.n4 drain_left.t6 2.2005
R196 drain_left.n5 drain_left.t13 2.2005
R197 drain_left.n5 drain_left.t4 2.2005
R198 drain_left.n1 drain_left.t9 2.2005
R199 drain_left.n1 drain_left.t17 2.2005
R200 drain_left.n0 drain_left.t8 2.2005
R201 drain_left.n0 drain_left.t0 2.2005
R202 drain_left.n15 drain_left.t10 2.2005
R203 drain_left.n15 drain_left.t3 2.2005
R204 drain_left.n13 drain_left.t2 2.2005
R205 drain_left.n13 drain_left.t19 2.2005
R206 drain_left.n11 drain_left.t14 2.2005
R207 drain_left.n11 drain_left.t7 2.2005
R208 drain_left.n9 drain_left.t5 2.2005
R209 drain_left.n9 drain_left.t1 2.2005
R210 drain_left.n8 drain_left.t16 2.2005
R211 drain_left.n8 drain_left.t11 2.2005
R212 drain_left.n12 drain_left.n10 0.543603
R213 drain_left.n14 drain_left.n12 0.543603
R214 drain_left.n16 drain_left.n14 0.543603
R215 drain_left.n7 drain_left.n6 0.488257
R216 drain_left.n7 drain_left.n2 0.488257
R217 minus.n27 minus.t6 876.365
R218 minus.n7 minus.t13 876.365
R219 minus.n56 minus.t19 876.365
R220 minus.n35 minus.t18 876.365
R221 minus.n26 minus.t2 827.433
R222 minus.n24 minus.t16 827.433
R223 minus.n3 minus.t5 827.433
R224 minus.n18 minus.t0 827.433
R225 minus.n16 minus.t14 827.433
R226 minus.n4 minus.t9 827.433
R227 minus.n10 minus.t1 827.433
R228 minus.n6 minus.t15 827.433
R229 minus.n55 minus.t10 827.433
R230 minus.n53 minus.t11 827.433
R231 minus.n47 minus.t3 827.433
R232 minus.n46 minus.t12 827.433
R233 minus.n44 minus.t4 827.433
R234 minus.n32 minus.t7 827.433
R235 minus.n38 minus.t17 827.433
R236 minus.n34 minus.t8 827.433
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 64.9975
R264 minus.n15 minus.n4 64.9975
R265 minus.n43 minus.n32 64.9975
R266 minus.n48 minus.n47 64.9975
R267 minus.n25 minus.n24 62.0763
R268 minus.n10 minus.n9 62.0763
R269 minus.n38 minus.n37 62.0763
R270 minus.n54 minus.n53 62.0763
R271 minus.n18 minus.n17 46.0096
R272 minus.n17 minus.n16 46.0096
R273 minus.n45 minus.n44 46.0096
R274 minus.n46 minus.n45 46.0096
R275 minus.n27 minus.n26 43.0884
R276 minus.n7 minus.n6 43.0884
R277 minus.n35 minus.n34 43.0884
R278 minus.n56 minus.n55 43.0884
R279 minus.n58 minus.n28 34.8263
R280 minus.n26 minus.n25 29.9429
R281 minus.n9 minus.n6 29.9429
R282 minus.n37 minus.n34 29.9429
R283 minus.n55 minus.n54 29.9429
R284 minus.n19 minus.n18 27.0217
R285 minus.n16 minus.n15 27.0217
R286 minus.n44 minus.n43 27.0217
R287 minus.n48 minus.n46 27.0217
R288 minus.n24 minus.n23 10.955
R289 minus.n11 minus.n10 10.955
R290 minus.n39 minus.n38 10.955
R291 minus.n53 minus.n52 10.955
R292 minus.n3 minus.n1 8.03383
R293 minus.n12 minus.n4 8.03383
R294 minus.n40 minus.n32 8.03383
R295 minus.n47 minus.n30 8.03383
R296 minus.n58 minus.n57 6.51565
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 66.0805
R317 drain_right.n6 drain_right.n4 66.0804
R318 drain_right.n2 drain_right.n0 66.0804
R319 drain_right.n10 drain_right.n9 65.5376
R320 drain_right.n12 drain_right.n11 65.5376
R321 drain_right.n14 drain_right.n13 65.5376
R322 drain_right.n16 drain_right.n15 65.5376
R323 drain_right.n7 drain_right.n3 65.5373
R324 drain_right.n6 drain_right.n5 65.5373
R325 drain_right.n2 drain_right.n1 65.5373
R326 drain_right drain_right.n7 28.8859
R327 drain_right drain_right.n16 6.19632
R328 drain_right.n3 drain_right.t15 2.2005
R329 drain_right.n3 drain_right.t7 2.2005
R330 drain_right.n4 drain_right.t9 2.2005
R331 drain_right.n4 drain_right.t0 2.2005
R332 drain_right.n5 drain_right.t16 2.2005
R333 drain_right.n5 drain_right.t8 2.2005
R334 drain_right.n1 drain_right.t2 2.2005
R335 drain_right.n1 drain_right.t12 2.2005
R336 drain_right.n0 drain_right.t1 2.2005
R337 drain_right.n0 drain_right.t11 2.2005
R338 drain_right.n8 drain_right.t4 2.2005
R339 drain_right.n8 drain_right.t6 2.2005
R340 drain_right.n9 drain_right.t10 2.2005
R341 drain_right.n9 drain_right.t18 2.2005
R342 drain_right.n11 drain_right.t19 2.2005
R343 drain_right.n11 drain_right.t5 2.2005
R344 drain_right.n13 drain_right.t3 2.2005
R345 drain_right.n13 drain_right.t14 2.2005
R346 drain_right.n15 drain_right.t13 2.2005
R347 drain_right.n15 drain_right.t17 2.2005
R348 drain_right.n16 drain_right.n14 0.543603
R349 drain_right.n14 drain_right.n12 0.543603
R350 drain_right.n12 drain_right.n10 0.543603
R351 drain_right.n7 drain_right.n6 0.488257
R352 drain_right.n7 drain_right.n2 0.488257
C0 drain_right plus 0.36079f
C1 drain_right minus 5.53266f
C2 drain_right source 28.9217f
C3 drain_left plus 5.73862f
C4 drain_left minus 0.171748f
C5 plus minus 5.21889f
C6 drain_left source 28.921299f
C7 plus source 5.4182f
C8 minus source 5.40416f
C9 drain_left drain_right 1.10832f
C10 drain_right a_n2102_n2688# 6.27777f
C11 drain_left a_n2102_n2688# 6.59791f
C12 source a_n2102_n2688# 7.198724f
C13 minus a_n2102_n2688# 8.04309f
C14 plus a_n2102_n2688# 9.860529f
C15 drain_right.t1 a_n2102_n2688# 0.240551f
C16 drain_right.t11 a_n2102_n2688# 0.240551f
C17 drain_right.n0 a_n2102_n2688# 2.10733f
C18 drain_right.t2 a_n2102_n2688# 0.240551f
C19 drain_right.t12 a_n2102_n2688# 0.240551f
C20 drain_right.n1 a_n2102_n2688# 2.10401f
C21 drain_right.n2 a_n2102_n2688# 0.784497f
C22 drain_right.t15 a_n2102_n2688# 0.240551f
C23 drain_right.t7 a_n2102_n2688# 0.240551f
C24 drain_right.n3 a_n2102_n2688# 2.10401f
C25 drain_right.t9 a_n2102_n2688# 0.240551f
C26 drain_right.t0 a_n2102_n2688# 0.240551f
C27 drain_right.n4 a_n2102_n2688# 2.10733f
C28 drain_right.t16 a_n2102_n2688# 0.240551f
C29 drain_right.t8 a_n2102_n2688# 0.240551f
C30 drain_right.n5 a_n2102_n2688# 2.10401f
C31 drain_right.n6 a_n2102_n2688# 0.784497f
C32 drain_right.n7 a_n2102_n2688# 1.78228f
C33 drain_right.t4 a_n2102_n2688# 0.240551f
C34 drain_right.t6 a_n2102_n2688# 0.240551f
C35 drain_right.n8 a_n2102_n2688# 2.10732f
C36 drain_right.t10 a_n2102_n2688# 0.240551f
C37 drain_right.t18 a_n2102_n2688# 0.240551f
C38 drain_right.n9 a_n2102_n2688# 2.10402f
C39 drain_right.n10 a_n2102_n2688# 0.788922f
C40 drain_right.t19 a_n2102_n2688# 0.240551f
C41 drain_right.t5 a_n2102_n2688# 0.240551f
C42 drain_right.n11 a_n2102_n2688# 2.10402f
C43 drain_right.n12 a_n2102_n2688# 0.389301f
C44 drain_right.t3 a_n2102_n2688# 0.240551f
C45 drain_right.t14 a_n2102_n2688# 0.240551f
C46 drain_right.n13 a_n2102_n2688# 2.10402f
C47 drain_right.n14 a_n2102_n2688# 0.389301f
C48 drain_right.t13 a_n2102_n2688# 0.240551f
C49 drain_right.t17 a_n2102_n2688# 0.240551f
C50 drain_right.n15 a_n2102_n2688# 2.10402f
C51 drain_right.n16 a_n2102_n2688# 0.670829f
C52 minus.n0 a_n2102_n2688# 0.049141f
C53 minus.t6 a_n2102_n2688# 0.384959f
C54 minus.t2 a_n2102_n2688# 0.375965f
C55 minus.t16 a_n2102_n2688# 0.375965f
C56 minus.n1 a_n2102_n2688# 0.017968f
C57 minus.n2 a_n2102_n2688# 0.049141f
C58 minus.t5 a_n2102_n2688# 0.375965f
C59 minus.n3 a_n2102_n2688# 0.156996f
C60 minus.t0 a_n2102_n2688# 0.375965f
C61 minus.t14 a_n2102_n2688# 0.375965f
C62 minus.t9 a_n2102_n2688# 0.375965f
C63 minus.n4 a_n2102_n2688# 0.156996f
C64 minus.n5 a_n2102_n2688# 0.049141f
C65 minus.t1 a_n2102_n2688# 0.375965f
C66 minus.t15 a_n2102_n2688# 0.375965f
C67 minus.n6 a_n2102_n2688# 0.156996f
C68 minus.t13 a_n2102_n2688# 0.384959f
C69 minus.n7 a_n2102_n2688# 0.172407f
C70 minus.n8 a_n2102_n2688# 0.112448f
C71 minus.n9 a_n2102_n2688# 0.02024f
C72 minus.n10 a_n2102_n2688# 0.156996f
C73 minus.n11 a_n2102_n2688# 0.018574f
C74 minus.n12 a_n2102_n2688# 0.017968f
C75 minus.n13 a_n2102_n2688# 0.049141f
C76 minus.n14 a_n2102_n2688# 0.049141f
C77 minus.n15 a_n2102_n2688# 0.02024f
C78 minus.n16 a_n2102_n2688# 0.156996f
C79 minus.n17 a_n2102_n2688# 0.02024f
C80 minus.n18 a_n2102_n2688# 0.156996f
C81 minus.n19 a_n2102_n2688# 0.02024f
C82 minus.n20 a_n2102_n2688# 0.049141f
C83 minus.n21 a_n2102_n2688# 0.049141f
C84 minus.n22 a_n2102_n2688# 0.049141f
C85 minus.n23 a_n2102_n2688# 0.018574f
C86 minus.n24 a_n2102_n2688# 0.156996f
C87 minus.n25 a_n2102_n2688# 0.02024f
C88 minus.n26 a_n2102_n2688# 0.156996f
C89 minus.n27 a_n2102_n2688# 0.172333f
C90 minus.n28 a_n2102_n2688# 1.63498f
C91 minus.n29 a_n2102_n2688# 0.049141f
C92 minus.t10 a_n2102_n2688# 0.375965f
C93 minus.t11 a_n2102_n2688# 0.375965f
C94 minus.n30 a_n2102_n2688# 0.017968f
C95 minus.n31 a_n2102_n2688# 0.049141f
C96 minus.t12 a_n2102_n2688# 0.375965f
C97 minus.t4 a_n2102_n2688# 0.375965f
C98 minus.t7 a_n2102_n2688# 0.375965f
C99 minus.n32 a_n2102_n2688# 0.156996f
C100 minus.n33 a_n2102_n2688# 0.049141f
C101 minus.t17 a_n2102_n2688# 0.375965f
C102 minus.t8 a_n2102_n2688# 0.375965f
C103 minus.n34 a_n2102_n2688# 0.156996f
C104 minus.t18 a_n2102_n2688# 0.384959f
C105 minus.n35 a_n2102_n2688# 0.172407f
C106 minus.n36 a_n2102_n2688# 0.112448f
C107 minus.n37 a_n2102_n2688# 0.02024f
C108 minus.n38 a_n2102_n2688# 0.156996f
C109 minus.n39 a_n2102_n2688# 0.018574f
C110 minus.n40 a_n2102_n2688# 0.017968f
C111 minus.n41 a_n2102_n2688# 0.049141f
C112 minus.n42 a_n2102_n2688# 0.049141f
C113 minus.n43 a_n2102_n2688# 0.02024f
C114 minus.n44 a_n2102_n2688# 0.156996f
C115 minus.n45 a_n2102_n2688# 0.02024f
C116 minus.n46 a_n2102_n2688# 0.156996f
C117 minus.t3 a_n2102_n2688# 0.375965f
C118 minus.n47 a_n2102_n2688# 0.156996f
C119 minus.n48 a_n2102_n2688# 0.02024f
C120 minus.n49 a_n2102_n2688# 0.049141f
C121 minus.n50 a_n2102_n2688# 0.049141f
C122 minus.n51 a_n2102_n2688# 0.049141f
C123 minus.n52 a_n2102_n2688# 0.018574f
C124 minus.n53 a_n2102_n2688# 0.156996f
C125 minus.n54 a_n2102_n2688# 0.02024f
C126 minus.n55 a_n2102_n2688# 0.156996f
C127 minus.t19 a_n2102_n2688# 0.384959f
C128 minus.n56 a_n2102_n2688# 0.172333f
C129 minus.n57 a_n2102_n2688# 0.323082f
C130 minus.n58 a_n2102_n2688# 1.99323f
C131 drain_left.t8 a_n2102_n2688# 0.241022f
C132 drain_left.t0 a_n2102_n2688# 0.241022f
C133 drain_left.n0 a_n2102_n2688# 2.11146f
C134 drain_left.t9 a_n2102_n2688# 0.241022f
C135 drain_left.t17 a_n2102_n2688# 0.241022f
C136 drain_left.n1 a_n2102_n2688# 2.10814f
C137 drain_left.n2 a_n2102_n2688# 0.786035f
C138 drain_left.t12 a_n2102_n2688# 0.241022f
C139 drain_left.t18 a_n2102_n2688# 0.241022f
C140 drain_left.n3 a_n2102_n2688# 2.10814f
C141 drain_left.t15 a_n2102_n2688# 0.241022f
C142 drain_left.t6 a_n2102_n2688# 0.241022f
C143 drain_left.n4 a_n2102_n2688# 2.11146f
C144 drain_left.t13 a_n2102_n2688# 0.241022f
C145 drain_left.t4 a_n2102_n2688# 0.241022f
C146 drain_left.n5 a_n2102_n2688# 2.10814f
C147 drain_left.n6 a_n2102_n2688# 0.786035f
C148 drain_left.n7 a_n2102_n2688# 1.85521f
C149 drain_left.t16 a_n2102_n2688# 0.241022f
C150 drain_left.t11 a_n2102_n2688# 0.241022f
C151 drain_left.n8 a_n2102_n2688# 2.11146f
C152 drain_left.t5 a_n2102_n2688# 0.241022f
C153 drain_left.t1 a_n2102_n2688# 0.241022f
C154 drain_left.n9 a_n2102_n2688# 2.10814f
C155 drain_left.n10 a_n2102_n2688# 0.790459f
C156 drain_left.t14 a_n2102_n2688# 0.241022f
C157 drain_left.t7 a_n2102_n2688# 0.241022f
C158 drain_left.n11 a_n2102_n2688# 2.10814f
C159 drain_left.n12 a_n2102_n2688# 0.390064f
C160 drain_left.t2 a_n2102_n2688# 0.241022f
C161 drain_left.t19 a_n2102_n2688# 0.241022f
C162 drain_left.n13 a_n2102_n2688# 2.10814f
C163 drain_left.n14 a_n2102_n2688# 0.390064f
C164 drain_left.t10 a_n2102_n2688# 0.241022f
C165 drain_left.t3 a_n2102_n2688# 0.241022f
C166 drain_left.n15 a_n2102_n2688# 2.10813f
C167 drain_left.n16 a_n2102_n2688# 0.672153f
C168 source.t19 a_n2102_n2688# 2.27217f
C169 source.n0 a_n2102_n2688# 1.30656f
C170 source.t30 a_n2102_n2688# 0.21308f
C171 source.t28 a_n2102_n2688# 0.21308f
C172 source.n1 a_n2102_n2688# 1.78377f
C173 source.n2 a_n2102_n2688# 0.384097f
C174 source.t31 a_n2102_n2688# 0.21308f
C175 source.t18 a_n2102_n2688# 0.21308f
C176 source.n3 a_n2102_n2688# 1.78377f
C177 source.n4 a_n2102_n2688# 0.384097f
C178 source.t34 a_n2102_n2688# 0.21308f
C179 source.t36 a_n2102_n2688# 0.21308f
C180 source.n5 a_n2102_n2688# 1.78377f
C181 source.n6 a_n2102_n2688# 0.384097f
C182 source.t20 a_n2102_n2688# 0.21308f
C183 source.t29 a_n2102_n2688# 0.21308f
C184 source.n7 a_n2102_n2688# 1.78377f
C185 source.n8 a_n2102_n2688# 0.384097f
C186 source.t33 a_n2102_n2688# 2.27218f
C187 source.n9 a_n2102_n2688# 0.46974f
C188 source.t38 a_n2102_n2688# 2.27218f
C189 source.n10 a_n2102_n2688# 0.46974f
C190 source.t9 a_n2102_n2688# 0.21308f
C191 source.t6 a_n2102_n2688# 0.21308f
C192 source.n11 a_n2102_n2688# 1.78377f
C193 source.n12 a_n2102_n2688# 0.384097f
C194 source.t12 a_n2102_n2688# 0.21308f
C195 source.t3 a_n2102_n2688# 0.21308f
C196 source.n13 a_n2102_n2688# 1.78377f
C197 source.n14 a_n2102_n2688# 0.384097f
C198 source.t2 a_n2102_n2688# 0.21308f
C199 source.t5 a_n2102_n2688# 0.21308f
C200 source.n15 a_n2102_n2688# 1.78377f
C201 source.n16 a_n2102_n2688# 0.384097f
C202 source.t10 a_n2102_n2688# 0.21308f
C203 source.t7 a_n2102_n2688# 0.21308f
C204 source.n17 a_n2102_n2688# 1.78377f
C205 source.n18 a_n2102_n2688# 0.384097f
C206 source.t39 a_n2102_n2688# 2.27218f
C207 source.n19 a_n2102_n2688# 1.74188f
C208 source.t35 a_n2102_n2688# 2.27217f
C209 source.n20 a_n2102_n2688# 1.74188f
C210 source.t25 a_n2102_n2688# 0.21308f
C211 source.t37 a_n2102_n2688# 0.21308f
C212 source.n21 a_n2102_n2688# 1.78376f
C213 source.n22 a_n2102_n2688# 0.384102f
C214 source.t21 a_n2102_n2688# 0.21308f
C215 source.t24 a_n2102_n2688# 0.21308f
C216 source.n23 a_n2102_n2688# 1.78376f
C217 source.n24 a_n2102_n2688# 0.384102f
C218 source.t32 a_n2102_n2688# 0.21308f
C219 source.t27 a_n2102_n2688# 0.21308f
C220 source.n25 a_n2102_n2688# 1.78376f
C221 source.n26 a_n2102_n2688# 0.384102f
C222 source.t23 a_n2102_n2688# 0.21308f
C223 source.t26 a_n2102_n2688# 0.21308f
C224 source.n27 a_n2102_n2688# 1.78376f
C225 source.n28 a_n2102_n2688# 0.384102f
C226 source.t22 a_n2102_n2688# 2.27217f
C227 source.n29 a_n2102_n2688# 0.469745f
C228 source.t16 a_n2102_n2688# 2.27217f
C229 source.n30 a_n2102_n2688# 0.469745f
C230 source.t0 a_n2102_n2688# 0.21308f
C231 source.t17 a_n2102_n2688# 0.21308f
C232 source.n31 a_n2102_n2688# 1.78376f
C233 source.n32 a_n2102_n2688# 0.384102f
C234 source.t4 a_n2102_n2688# 0.21308f
C235 source.t1 a_n2102_n2688# 0.21308f
C236 source.n33 a_n2102_n2688# 1.78376f
C237 source.n34 a_n2102_n2688# 0.384102f
C238 source.t15 a_n2102_n2688# 0.21308f
C239 source.t14 a_n2102_n2688# 0.21308f
C240 source.n35 a_n2102_n2688# 1.78376f
C241 source.n36 a_n2102_n2688# 0.384102f
C242 source.t11 a_n2102_n2688# 0.21308f
C243 source.t13 a_n2102_n2688# 0.21308f
C244 source.n37 a_n2102_n2688# 1.78376f
C245 source.n38 a_n2102_n2688# 0.384102f
C246 source.t8 a_n2102_n2688# 2.27217f
C247 source.n39 a_n2102_n2688# 0.638871f
C248 source.n40 a_n2102_n2688# 1.55965f
C249 plus.n0 a_n2102_n2688# 0.05006f
C250 plus.t9 a_n2102_n2688# 0.383f
C251 plus.t0 a_n2102_n2688# 0.383f
C252 plus.n1 a_n2102_n2688# 0.018304f
C253 plus.n2 a_n2102_n2688# 0.05006f
C254 plus.t12 a_n2102_n2688# 0.383f
C255 plus.t5 a_n2102_n2688# 0.383f
C256 plus.t18 a_n2102_n2688# 0.383f
C257 plus.n3 a_n2102_n2688# 0.159934f
C258 plus.n4 a_n2102_n2688# 0.05006f
C259 plus.t14 a_n2102_n2688# 0.383f
C260 plus.t8 a_n2102_n2688# 0.383f
C261 plus.n5 a_n2102_n2688# 0.159934f
C262 plus.t3 a_n2102_n2688# 0.392162f
C263 plus.n6 a_n2102_n2688# 0.175633f
C264 plus.n7 a_n2102_n2688# 0.114552f
C265 plus.n8 a_n2102_n2688# 0.020619f
C266 plus.n9 a_n2102_n2688# 0.159934f
C267 plus.n10 a_n2102_n2688# 0.018921f
C268 plus.n11 a_n2102_n2688# 0.018304f
C269 plus.n12 a_n2102_n2688# 0.05006f
C270 plus.n13 a_n2102_n2688# 0.05006f
C271 plus.n14 a_n2102_n2688# 0.020619f
C272 plus.n15 a_n2102_n2688# 0.159934f
C273 plus.n16 a_n2102_n2688# 0.020619f
C274 plus.n17 a_n2102_n2688# 0.159934f
C275 plus.t17 a_n2102_n2688# 0.383f
C276 plus.n18 a_n2102_n2688# 0.159934f
C277 plus.n19 a_n2102_n2688# 0.020619f
C278 plus.n20 a_n2102_n2688# 0.05006f
C279 plus.n21 a_n2102_n2688# 0.05006f
C280 plus.n22 a_n2102_n2688# 0.05006f
C281 plus.n23 a_n2102_n2688# 0.018921f
C282 plus.n24 a_n2102_n2688# 0.159934f
C283 plus.n25 a_n2102_n2688# 0.020619f
C284 plus.n26 a_n2102_n2688# 0.159934f
C285 plus.t16 a_n2102_n2688# 0.392162f
C286 plus.n27 a_n2102_n2688# 0.175557f
C287 plus.n28 a_n2102_n2688# 0.493643f
C288 plus.n29 a_n2102_n2688# 0.05006f
C289 plus.t11 a_n2102_n2688# 0.392162f
C290 plus.t19 a_n2102_n2688# 0.383f
C291 plus.t10 a_n2102_n2688# 0.383f
C292 plus.n30 a_n2102_n2688# 0.018304f
C293 plus.n31 a_n2102_n2688# 0.05006f
C294 plus.t2 a_n2102_n2688# 0.383f
C295 plus.n32 a_n2102_n2688# 0.159934f
C296 plus.t7 a_n2102_n2688# 0.383f
C297 plus.t1 a_n2102_n2688# 0.383f
C298 plus.t6 a_n2102_n2688# 0.383f
C299 plus.n33 a_n2102_n2688# 0.159934f
C300 plus.n34 a_n2102_n2688# 0.05006f
C301 plus.t15 a_n2102_n2688# 0.383f
C302 plus.t4 a_n2102_n2688# 0.383f
C303 plus.n35 a_n2102_n2688# 0.159934f
C304 plus.t13 a_n2102_n2688# 0.392162f
C305 plus.n36 a_n2102_n2688# 0.175633f
C306 plus.n37 a_n2102_n2688# 0.114552f
C307 plus.n38 a_n2102_n2688# 0.020619f
C308 plus.n39 a_n2102_n2688# 0.159934f
C309 plus.n40 a_n2102_n2688# 0.018921f
C310 plus.n41 a_n2102_n2688# 0.018304f
C311 plus.n42 a_n2102_n2688# 0.05006f
C312 plus.n43 a_n2102_n2688# 0.05006f
C313 plus.n44 a_n2102_n2688# 0.020619f
C314 plus.n45 a_n2102_n2688# 0.159934f
C315 plus.n46 a_n2102_n2688# 0.020619f
C316 plus.n47 a_n2102_n2688# 0.159934f
C317 plus.n48 a_n2102_n2688# 0.020619f
C318 plus.n49 a_n2102_n2688# 0.05006f
C319 plus.n50 a_n2102_n2688# 0.05006f
C320 plus.n51 a_n2102_n2688# 0.05006f
C321 plus.n52 a_n2102_n2688# 0.018921f
C322 plus.n53 a_n2102_n2688# 0.159934f
C323 plus.n54 a_n2102_n2688# 0.020619f
C324 plus.n55 a_n2102_n2688# 0.159934f
C325 plus.n56 a_n2102_n2688# 0.175557f
C326 plus.n57 a_n2102_n2688# 1.4547f
.ends

