* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t11 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 source.t26 plus.t1 drain_left.t9 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 drain_right.t13 minus.t0 source.t6 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X3 source.t8 minus.t1 drain_right.t12 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X4 source.t2 minus.t2 drain_right.t11 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X5 source.t0 minus.t3 drain_right.t10 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X6 drain_left.t12 plus.t2 source.t25 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X7 source.t24 plus.t3 drain_left.t4 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X8 drain_left.t5 plus.t4 source.t23 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X9 drain_left.t6 plus.t5 source.t22 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X10 source.t1 minus.t4 drain_right.t9 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X11 drain_left.t0 plus.t6 source.t21 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X12 drain_left.t10 plus.t7 source.t20 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X13 a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X14 source.t19 plus.t8 drain_left.t1 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X15 drain_left.t8 plus.t9 source.t18 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X16 drain_left.t2 plus.t10 source.t17 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X17 drain_left.t3 plus.t11 source.t16 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 source.t15 plus.t12 drain_left.t7 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X19 drain_right.t8 minus.t5 source.t3 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X20 drain_right.t7 minus.t6 source.t10 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X21 source.t5 minus.t7 drain_right.t6 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X22 a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X23 source.t12 minus.t8 drain_right.t5 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X24 drain_right.t4 minus.t9 source.t13 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X25 drain_right.t3 minus.t10 source.t4 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X26 drain_right.t2 minus.t11 source.t9 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X27 drain_right.t1 minus.t12 source.t11 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X28 source.t14 plus.t13 drain_left.t13 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X29 a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X30 a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X31 drain_right.t0 minus.t13 source.t7 a_n1644_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n3 plus.t2 449.575
R1 plus.n15 plus.t9 449.575
R2 plus.n20 plus.t5 449.575
R3 plus.n32 plus.t6 449.575
R4 plus.n1 plus.t0 414.521
R5 plus.n4 plus.t1 414.521
R6 plus.n6 plus.t11 414.521
R7 plus.n12 plus.t10 414.521
R8 plus.n14 plus.t13 414.521
R9 plus.n18 plus.t12 414.521
R10 plus.n21 plus.t3 414.521
R11 plus.n23 plus.t7 414.521
R12 plus.n29 plus.t4 414.521
R13 plus.n31 plus.t8 414.521
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 25.7717
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus.n7 plus.n6 11.6853
R46 plus.n12 plus.n11 11.6853
R47 plus.n29 plus.n28 11.6853
R48 plus.n24 plus.n23 11.6853
R49 plus plus.n16 8.68611
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t12 86.8731
R61 drain_left.n1 drain_left.t0 86.873
R62 drain_left.n4 drain_left.n2 80.273
R63 drain_left.n11 drain_left.n10 79.7731
R64 drain_left.n9 drain_left.n8 79.7731
R65 drain_left.n7 drain_left.n6 79.7731
R66 drain_left.n4 drain_left.n3 79.773
R67 drain_left.n1 drain_left.n0 79.773
R68 drain_left drain_left.n5 23.4239
R69 drain_left.n2 drain_left.t4 6.6005
R70 drain_left.n2 drain_left.t6 6.6005
R71 drain_left.n3 drain_left.t7 6.6005
R72 drain_left.n3 drain_left.t10 6.6005
R73 drain_left.n0 drain_left.t1 6.6005
R74 drain_left.n0 drain_left.t5 6.6005
R75 drain_left.n10 drain_left.t13 6.6005
R76 drain_left.n10 drain_left.t8 6.6005
R77 drain_left.n8 drain_left.t11 6.6005
R78 drain_left.n8 drain_left.t2 6.6005
R79 drain_left.n6 drain_left.t9 6.6005
R80 drain_left.n6 drain_left.t3 6.6005
R81 drain_left drain_left.n11 6.15322
R82 drain_left.n9 drain_left.n7 0.5005
R83 drain_left.n11 drain_left.n9 0.5005
R84 drain_left.n5 drain_left.n1 0.320154
R85 drain_left.n5 drain_left.n4 0.070154
R86 source.n0 source.t18 69.6943
R87 source.n7 source.t10 69.6943
R88 source.n27 source.t6 69.6942
R89 source.n20 source.t22 69.6942
R90 source.n2 source.n1 63.0943
R91 source.n4 source.n3 63.0943
R92 source.n6 source.n5 63.0943
R93 source.n9 source.n8 63.0943
R94 source.n11 source.n10 63.0943
R95 source.n13 source.n12 63.0943
R96 source.n26 source.n25 63.0942
R97 source.n24 source.n23 63.0942
R98 source.n22 source.n21 63.0942
R99 source.n19 source.n18 63.0942
R100 source.n17 source.n16 63.0942
R101 source.n15 source.n14 63.0942
R102 source.n15 source.n13 15.4695
R103 source.n28 source.n0 9.45661
R104 source.n25 source.t11 6.6005
R105 source.n25 source.t2 6.6005
R106 source.n23 source.t13 6.6005
R107 source.n23 source.t12 6.6005
R108 source.n21 source.t7 6.6005
R109 source.n21 source.t5 6.6005
R110 source.n18 source.t20 6.6005
R111 source.n18 source.t24 6.6005
R112 source.n16 source.t23 6.6005
R113 source.n16 source.t15 6.6005
R114 source.n14 source.t21 6.6005
R115 source.n14 source.t19 6.6005
R116 source.n1 source.t17 6.6005
R117 source.n1 source.t14 6.6005
R118 source.n3 source.t16 6.6005
R119 source.n3 source.t27 6.6005
R120 source.n5 source.t25 6.6005
R121 source.n5 source.t26 6.6005
R122 source.n8 source.t3 6.6005
R123 source.n8 source.t0 6.6005
R124 source.n10 source.t4 6.6005
R125 source.n10 source.t8 6.6005
R126 source.n12 source.t9 6.6005
R127 source.n12 source.t1 6.6005
R128 source.n28 source.n27 5.51343
R129 source.n7 source.n6 0.720328
R130 source.n22 source.n20 0.720328
R131 source.n13 source.n11 0.5005
R132 source.n11 source.n9 0.5005
R133 source.n9 source.n7 0.5005
R134 source.n6 source.n4 0.5005
R135 source.n4 source.n2 0.5005
R136 source.n2 source.n0 0.5005
R137 source.n17 source.n15 0.5005
R138 source.n19 source.n17 0.5005
R139 source.n20 source.n19 0.5005
R140 source.n24 source.n22 0.5005
R141 source.n26 source.n24 0.5005
R142 source.n27 source.n26 0.5005
R143 source source.n28 0.188
R144 minus.n15 minus.t11 449.575
R145 minus.n3 minus.t6 449.575
R146 minus.n32 minus.t0 449.575
R147 minus.n20 minus.t13 449.575
R148 minus.n1 minus.t1 414.521
R149 minus.n14 minus.t4 414.521
R150 minus.n12 minus.t10 414.521
R151 minus.n6 minus.t5 414.521
R152 minus.n4 minus.t3 414.521
R153 minus.n18 minus.t8 414.521
R154 minus.n31 minus.t2 414.521
R155 minus.n29 minus.t12 414.521
R156 minus.n23 minus.t9 414.521
R157 minus.n21 minus.t7 414.521
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 61.346
R177 minus.n6 minus.n5 61.346
R178 minus.n23 minus.n22 61.346
R179 minus.n30 minus.n29 61.346
R180 minus.n15 minus.n14 49.6611
R181 minus.n4 minus.n3 49.6611
R182 minus.n21 minus.n20 49.6611
R183 minus.n32 minus.n31 49.6611
R184 minus.n34 minus.n16 28.4816
R185 minus.n14 minus.n13 23.3702
R186 minus.n5 minus.n4 23.3702
R187 minus.n22 minus.n21 23.3702
R188 minus.n31 minus.n30 23.3702
R189 minus.n12 minus.n11 11.6853
R190 minus.n7 minus.n6 11.6853
R191 minus.n24 minus.n23 11.6853
R192 minus.n29 minus.n28 11.6853
R193 minus.n34 minus.n33 6.45126
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t0 86.873
R206 drain_right.n11 drain_right.t2 86.3731
R207 drain_right.n8 drain_right.n6 80.2731
R208 drain_right.n4 drain_right.n2 80.273
R209 drain_right.n8 drain_right.n7 79.7731
R210 drain_right.n10 drain_right.n9 79.7731
R211 drain_right.n4 drain_right.n3 79.773
R212 drain_right.n1 drain_right.n0 79.773
R213 drain_right drain_right.n5 22.8707
R214 drain_right.n2 drain_right.t11 6.6005
R215 drain_right.n2 drain_right.t13 6.6005
R216 drain_right.n3 drain_right.t5 6.6005
R217 drain_right.n3 drain_right.t1 6.6005
R218 drain_right.n0 drain_right.t6 6.6005
R219 drain_right.n0 drain_right.t4 6.6005
R220 drain_right.n6 drain_right.t10 6.6005
R221 drain_right.n6 drain_right.t7 6.6005
R222 drain_right.n7 drain_right.t12 6.6005
R223 drain_right.n7 drain_right.t8 6.6005
R224 drain_right.n9 drain_right.t9 6.6005
R225 drain_right.n9 drain_right.t3 6.6005
R226 drain_right drain_right.n11 5.90322
R227 drain_right.n11 drain_right.n10 0.5005
R228 drain_right.n10 drain_right.n8 0.5005
R229 drain_right.n5 drain_right.n1 0.320154
R230 drain_right.n5 drain_right.n4 0.070154
C0 drain_right drain_left 0.83729f
C1 drain_right source 9.545889f
C2 minus drain_left 0.176767f
C3 plus drain_left 1.66235f
C4 minus source 1.59073f
C5 plus source 1.6049f
C6 source drain_left 9.54951f
C7 drain_right minus 1.50477f
C8 drain_right plus 0.318971f
C9 plus minus 3.54619f
C10 drain_right a_n1644_n1488# 4.24343f
C11 drain_left a_n1644_n1488# 4.48474f
C12 source a_n1644_n1488# 2.885928f
C13 minus a_n1644_n1488# 5.668163f
C14 plus a_n1644_n1488# 6.292076f
C15 drain_right.t0 a_n1644_n1488# 0.589239f
C16 drain_right.t6 a_n1644_n1488# 0.063466f
C17 drain_right.t4 a_n1644_n1488# 0.063466f
C18 drain_right.n0 a_n1644_n1488# 0.457709f
C19 drain_right.n1 a_n1644_n1488# 0.596715f
C20 drain_right.t11 a_n1644_n1488# 0.063466f
C21 drain_right.t13 a_n1644_n1488# 0.063466f
C22 drain_right.n2 a_n1644_n1488# 0.459648f
C23 drain_right.t5 a_n1644_n1488# 0.063466f
C24 drain_right.t1 a_n1644_n1488# 0.063466f
C25 drain_right.n3 a_n1644_n1488# 0.457709f
C26 drain_right.n4 a_n1644_n1488# 0.581752f
C27 drain_right.n5 a_n1644_n1488# 0.695257f
C28 drain_right.t10 a_n1644_n1488# 0.063466f
C29 drain_right.t7 a_n1644_n1488# 0.063466f
C30 drain_right.n6 a_n1644_n1488# 0.45965f
C31 drain_right.t12 a_n1644_n1488# 0.063466f
C32 drain_right.t8 a_n1644_n1488# 0.063466f
C33 drain_right.n7 a_n1644_n1488# 0.457711f
C34 drain_right.n8 a_n1644_n1488# 0.609959f
C35 drain_right.t9 a_n1644_n1488# 0.063466f
C36 drain_right.t3 a_n1644_n1488# 0.063466f
C37 drain_right.n9 a_n1644_n1488# 0.457711f
C38 drain_right.n10 a_n1644_n1488# 0.300558f
C39 drain_right.t2 a_n1644_n1488# 0.587448f
C40 drain_right.n11 a_n1644_n1488# 0.532028f
C41 minus.n0 a_n1644_n1488# 0.027673f
C42 minus.t11 a_n1644_n1488# 0.062922f
C43 minus.t4 a_n1644_n1488# 0.060103f
C44 minus.t10 a_n1644_n1488# 0.060103f
C45 minus.t1 a_n1644_n1488# 0.060103f
C46 minus.n1 a_n1644_n1488# 0.045501f
C47 minus.n2 a_n1644_n1488# 0.059233f
C48 minus.t5 a_n1644_n1488# 0.060103f
C49 minus.t3 a_n1644_n1488# 0.060103f
C50 minus.t6 a_n1644_n1488# 0.062922f
C51 minus.n3 a_n1644_n1488# 0.043913f
C52 minus.n4 a_n1644_n1488# 0.036321f
C53 minus.n5 a_n1644_n1488# 0.010545f
C54 minus.n6 a_n1644_n1488# 0.036321f
C55 minus.n7 a_n1644_n1488# 0.010545f
C56 minus.n8 a_n1644_n1488# 0.027673f
C57 minus.n9 a_n1644_n1488# 0.027673f
C58 minus.n10 a_n1644_n1488# 0.027673f
C59 minus.n11 a_n1644_n1488# 0.010545f
C60 minus.n12 a_n1644_n1488# 0.036321f
C61 minus.n13 a_n1644_n1488# 0.010545f
C62 minus.n14 a_n1644_n1488# 0.036321f
C63 minus.n15 a_n1644_n1488# 0.043876f
C64 minus.n16 a_n1644_n1488# 0.656681f
C65 minus.n17 a_n1644_n1488# 0.027673f
C66 minus.t2 a_n1644_n1488# 0.060103f
C67 minus.t12 a_n1644_n1488# 0.060103f
C68 minus.t8 a_n1644_n1488# 0.060103f
C69 minus.n18 a_n1644_n1488# 0.045501f
C70 minus.n19 a_n1644_n1488# 0.059233f
C71 minus.t9 a_n1644_n1488# 0.060103f
C72 minus.t7 a_n1644_n1488# 0.060103f
C73 minus.t13 a_n1644_n1488# 0.062922f
C74 minus.n20 a_n1644_n1488# 0.043913f
C75 minus.n21 a_n1644_n1488# 0.036321f
C76 minus.n22 a_n1644_n1488# 0.010545f
C77 minus.n23 a_n1644_n1488# 0.036321f
C78 minus.n24 a_n1644_n1488# 0.010545f
C79 minus.n25 a_n1644_n1488# 0.027673f
C80 minus.n26 a_n1644_n1488# 0.027673f
C81 minus.n27 a_n1644_n1488# 0.027673f
C82 minus.n28 a_n1644_n1488# 0.010545f
C83 minus.n29 a_n1644_n1488# 0.036321f
C84 minus.n30 a_n1644_n1488# 0.010545f
C85 minus.n31 a_n1644_n1488# 0.036321f
C86 minus.t0 a_n1644_n1488# 0.062922f
C87 minus.n32 a_n1644_n1488# 0.043876f
C88 minus.n33 a_n1644_n1488# 0.177734f
C89 minus.n34 a_n1644_n1488# 0.813334f
C90 source.t18 a_n1644_n1488# 0.607501f
C91 source.n0 a_n1644_n1488# 0.821284f
C92 source.t17 a_n1644_n1488# 0.073159f
C93 source.t14 a_n1644_n1488# 0.073159f
C94 source.n1 a_n1644_n1488# 0.463872f
C95 source.n2 a_n1644_n1488# 0.368267f
C96 source.t16 a_n1644_n1488# 0.073159f
C97 source.t27 a_n1644_n1488# 0.073159f
C98 source.n3 a_n1644_n1488# 0.463872f
C99 source.n4 a_n1644_n1488# 0.368267f
C100 source.t25 a_n1644_n1488# 0.073159f
C101 source.t26 a_n1644_n1488# 0.073159f
C102 source.n5 a_n1644_n1488# 0.463872f
C103 source.n6 a_n1644_n1488# 0.390126f
C104 source.t10 a_n1644_n1488# 0.607501f
C105 source.n7 a_n1644_n1488# 0.446021f
C106 source.t3 a_n1644_n1488# 0.073159f
C107 source.t0 a_n1644_n1488# 0.073159f
C108 source.n8 a_n1644_n1488# 0.463872f
C109 source.n9 a_n1644_n1488# 0.368267f
C110 source.t4 a_n1644_n1488# 0.073159f
C111 source.t8 a_n1644_n1488# 0.073159f
C112 source.n10 a_n1644_n1488# 0.463872f
C113 source.n11 a_n1644_n1488# 0.368267f
C114 source.t9 a_n1644_n1488# 0.073159f
C115 source.t1 a_n1644_n1488# 0.073159f
C116 source.n12 a_n1644_n1488# 0.463872f
C117 source.n13 a_n1644_n1488# 1.13576f
C118 source.t21 a_n1644_n1488# 0.073159f
C119 source.t19 a_n1644_n1488# 0.073159f
C120 source.n14 a_n1644_n1488# 0.463868f
C121 source.n15 a_n1644_n1488# 1.13576f
C122 source.t23 a_n1644_n1488# 0.073159f
C123 source.t15 a_n1644_n1488# 0.073159f
C124 source.n16 a_n1644_n1488# 0.463868f
C125 source.n17 a_n1644_n1488# 0.36827f
C126 source.t20 a_n1644_n1488# 0.073159f
C127 source.t24 a_n1644_n1488# 0.073159f
C128 source.n18 a_n1644_n1488# 0.463868f
C129 source.n19 a_n1644_n1488# 0.36827f
C130 source.t22 a_n1644_n1488# 0.607498f
C131 source.n20 a_n1644_n1488# 0.446024f
C132 source.t7 a_n1644_n1488# 0.073159f
C133 source.t5 a_n1644_n1488# 0.073159f
C134 source.n21 a_n1644_n1488# 0.463868f
C135 source.n22 a_n1644_n1488# 0.390129f
C136 source.t13 a_n1644_n1488# 0.073159f
C137 source.t12 a_n1644_n1488# 0.073159f
C138 source.n23 a_n1644_n1488# 0.463868f
C139 source.n24 a_n1644_n1488# 0.36827f
C140 source.t11 a_n1644_n1488# 0.073159f
C141 source.t2 a_n1644_n1488# 0.073159f
C142 source.n25 a_n1644_n1488# 0.463868f
C143 source.n26 a_n1644_n1488# 0.36827f
C144 source.t6 a_n1644_n1488# 0.607498f
C145 source.n27 a_n1644_n1488# 0.591938f
C146 source.n28 a_n1644_n1488# 0.892602f
C147 drain_left.t0 a_n1644_n1488# 0.582814f
C148 drain_left.t1 a_n1644_n1488# 0.062774f
C149 drain_left.t5 a_n1644_n1488# 0.062774f
C150 drain_left.n0 a_n1644_n1488# 0.452718f
C151 drain_left.n1 a_n1644_n1488# 0.590209f
C152 drain_left.t4 a_n1644_n1488# 0.062774f
C153 drain_left.t6 a_n1644_n1488# 0.062774f
C154 drain_left.n2 a_n1644_n1488# 0.454636f
C155 drain_left.t7 a_n1644_n1488# 0.062774f
C156 drain_left.t10 a_n1644_n1488# 0.062774f
C157 drain_left.n3 a_n1644_n1488# 0.452718f
C158 drain_left.n4 a_n1644_n1488# 0.575409f
C159 drain_left.n5 a_n1644_n1488# 0.74027f
C160 drain_left.t12 a_n1644_n1488# 0.582816f
C161 drain_left.t9 a_n1644_n1488# 0.062774f
C162 drain_left.t3 a_n1644_n1488# 0.062774f
C163 drain_left.n6 a_n1644_n1488# 0.452721f
C164 drain_left.n7 a_n1644_n1488# 0.603671f
C165 drain_left.t11 a_n1644_n1488# 0.062774f
C166 drain_left.t2 a_n1644_n1488# 0.062774f
C167 drain_left.n8 a_n1644_n1488# 0.452721f
C168 drain_left.n9 a_n1644_n1488# 0.297281f
C169 drain_left.t13 a_n1644_n1488# 0.062774f
C170 drain_left.t8 a_n1644_n1488# 0.062774f
C171 drain_left.n10 a_n1644_n1488# 0.452721f
C172 drain_left.n11 a_n1644_n1488# 0.515848f
C173 plus.n0 a_n1644_n1488# 0.028123f
C174 plus.t13 a_n1644_n1488# 0.06108f
C175 plus.t10 a_n1644_n1488# 0.06108f
C176 plus.t0 a_n1644_n1488# 0.06108f
C177 plus.n1 a_n1644_n1488# 0.04624f
C178 plus.n2 a_n1644_n1488# 0.060196f
C179 plus.t11 a_n1644_n1488# 0.06108f
C180 plus.t1 a_n1644_n1488# 0.06108f
C181 plus.t2 a_n1644_n1488# 0.063945f
C182 plus.n3 a_n1644_n1488# 0.044627f
C183 plus.n4 a_n1644_n1488# 0.036911f
C184 plus.n5 a_n1644_n1488# 0.010716f
C185 plus.n6 a_n1644_n1488# 0.036911f
C186 plus.n7 a_n1644_n1488# 0.010716f
C187 plus.n8 a_n1644_n1488# 0.028123f
C188 plus.n9 a_n1644_n1488# 0.028123f
C189 plus.n10 a_n1644_n1488# 0.028123f
C190 plus.n11 a_n1644_n1488# 0.010716f
C191 plus.n12 a_n1644_n1488# 0.036911f
C192 plus.n13 a_n1644_n1488# 0.010716f
C193 plus.n14 a_n1644_n1488# 0.036911f
C194 plus.t9 a_n1644_n1488# 0.063945f
C195 plus.n15 a_n1644_n1488# 0.044589f
C196 plus.n16 a_n1644_n1488# 0.206668f
C197 plus.n17 a_n1644_n1488# 0.028123f
C198 plus.t6 a_n1644_n1488# 0.063945f
C199 plus.t8 a_n1644_n1488# 0.06108f
C200 plus.t4 a_n1644_n1488# 0.06108f
C201 plus.t12 a_n1644_n1488# 0.06108f
C202 plus.n18 a_n1644_n1488# 0.04624f
C203 plus.n19 a_n1644_n1488# 0.060196f
C204 plus.t7 a_n1644_n1488# 0.06108f
C205 plus.t3 a_n1644_n1488# 0.06108f
C206 plus.t5 a_n1644_n1488# 0.063945f
C207 plus.n20 a_n1644_n1488# 0.044627f
C208 plus.n21 a_n1644_n1488# 0.036911f
C209 plus.n22 a_n1644_n1488# 0.010716f
C210 plus.n23 a_n1644_n1488# 0.036911f
C211 plus.n24 a_n1644_n1488# 0.010716f
C212 plus.n25 a_n1644_n1488# 0.028123f
C213 plus.n26 a_n1644_n1488# 0.028123f
C214 plus.n27 a_n1644_n1488# 0.028123f
C215 plus.n28 a_n1644_n1488# 0.010716f
C216 plus.n29 a_n1644_n1488# 0.036911f
C217 plus.n30 a_n1644_n1488# 0.010716f
C218 plus.n31 a_n1644_n1488# 0.036911f
C219 plus.n32 a_n1644_n1488# 0.044589f
C220 plus.n33 a_n1644_n1488# 0.628495f
.ends

