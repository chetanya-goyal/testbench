* NGSPICE file created from diffpair262.ext - technology: sky130A

.subckt diffpair262 minus drain_right drain_left source plus
X0 source.t11 plus.t0 drain_left.t3 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_left.t1 plus.t1 source.t10 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X2 source.t0 minus.t0 drain_right.t5 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X4 drain_left.t4 plus.t2 source.t9 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X5 a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X6 source.t8 plus.t3 drain_left.t5 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X7 drain_right.t4 minus.t1 source.t2 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X8 drain_left.t2 plus.t4 source.t7 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X9 drain_left.t0 plus.t5 source.t6 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X10 a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X11 drain_right.t3 minus.t2 source.t5 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X12 drain_right.t2 minus.t3 source.t1 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X13 drain_right.t1 minus.t4 source.t4 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X14 source.t3 minus.t5 drain_right.t0 a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# a_n1180_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
R0 plus.n0 plus.t2 751.92
R1 plus.n2 plus.t4 751.92
R2 plus.n4 plus.t5 751.92
R3 plus.n6 plus.t1 751.92
R4 plus.n1 plus.t0 703.721
R5 plus.n5 plus.t3 703.721
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 25.1846
R15 plus plus.n3 9.85656
R16 drain_left.n26 drain_left.n0 289.615
R17 drain_left.n59 drain_left.n33 289.615
R18 drain_left.n11 drain_left.n10 185
R19 drain_left.n8 drain_left.n7 185
R20 drain_left.n17 drain_left.n16 185
R21 drain_left.n19 drain_left.n18 185
R22 drain_left.n4 drain_left.n3 185
R23 drain_left.n25 drain_left.n24 185
R24 drain_left.n27 drain_left.n26 185
R25 drain_left.n60 drain_left.n59 185
R26 drain_left.n58 drain_left.n57 185
R27 drain_left.n37 drain_left.n36 185
R28 drain_left.n52 drain_left.n51 185
R29 drain_left.n50 drain_left.n49 185
R30 drain_left.n41 drain_left.n40 185
R31 drain_left.n44 drain_left.n43 185
R32 drain_left.t1 drain_left.n9 147.661
R33 drain_left.t4 drain_left.n42 147.661
R34 drain_left.n10 drain_left.n7 104.615
R35 drain_left.n17 drain_left.n7 104.615
R36 drain_left.n18 drain_left.n17 104.615
R37 drain_left.n18 drain_left.n3 104.615
R38 drain_left.n25 drain_left.n3 104.615
R39 drain_left.n26 drain_left.n25 104.615
R40 drain_left.n59 drain_left.n58 104.615
R41 drain_left.n58 drain_left.n36 104.615
R42 drain_left.n51 drain_left.n36 104.615
R43 drain_left.n51 drain_left.n50 104.615
R44 drain_left.n50 drain_left.n40 104.615
R45 drain_left.n43 drain_left.n40 104.615
R46 drain_left.n32 drain_left.n31 67.2603
R47 drain_left.n65 drain_left.n64 67.1907
R48 drain_left.n10 drain_left.t1 52.3082
R49 drain_left.n43 drain_left.t4 52.3082
R50 drain_left.n65 drain_left.n63 49.3641
R51 drain_left.n32 drain_left.n30 49.1838
R52 drain_left drain_left.n32 24.1966
R53 drain_left.n11 drain_left.n9 15.6674
R54 drain_left.n44 drain_left.n42 15.6674
R55 drain_left.n12 drain_left.n8 12.8005
R56 drain_left.n45 drain_left.n41 12.8005
R57 drain_left.n16 drain_left.n15 12.0247
R58 drain_left.n49 drain_left.n48 12.0247
R59 drain_left.n19 drain_left.n6 11.249
R60 drain_left.n52 drain_left.n39 11.249
R61 drain_left.n20 drain_left.n4 10.4732
R62 drain_left.n53 drain_left.n37 10.4732
R63 drain_left.n24 drain_left.n23 9.69747
R64 drain_left.n57 drain_left.n56 9.69747
R65 drain_left.n30 drain_left.n29 9.45567
R66 drain_left.n63 drain_left.n62 9.45567
R67 drain_left.n29 drain_left.n28 9.3005
R68 drain_left.n2 drain_left.n1 9.3005
R69 drain_left.n23 drain_left.n22 9.3005
R70 drain_left.n21 drain_left.n20 9.3005
R71 drain_left.n6 drain_left.n5 9.3005
R72 drain_left.n15 drain_left.n14 9.3005
R73 drain_left.n13 drain_left.n12 9.3005
R74 drain_left.n62 drain_left.n61 9.3005
R75 drain_left.n35 drain_left.n34 9.3005
R76 drain_left.n56 drain_left.n55 9.3005
R77 drain_left.n54 drain_left.n53 9.3005
R78 drain_left.n39 drain_left.n38 9.3005
R79 drain_left.n48 drain_left.n47 9.3005
R80 drain_left.n46 drain_left.n45 9.3005
R81 drain_left.n27 drain_left.n2 8.92171
R82 drain_left.n60 drain_left.n35 8.92171
R83 drain_left.n28 drain_left.n0 8.14595
R84 drain_left.n61 drain_left.n33 8.14595
R85 drain_left drain_left.n65 6.15322
R86 drain_left.n30 drain_left.n0 5.81868
R87 drain_left.n63 drain_left.n33 5.81868
R88 drain_left.n28 drain_left.n27 5.04292
R89 drain_left.n61 drain_left.n60 5.04292
R90 drain_left.n13 drain_left.n9 4.38594
R91 drain_left.n46 drain_left.n42 4.38594
R92 drain_left.n24 drain_left.n2 4.26717
R93 drain_left.n57 drain_left.n35 4.26717
R94 drain_left.n23 drain_left.n4 3.49141
R95 drain_left.n56 drain_left.n37 3.49141
R96 drain_left.n31 drain_left.t5 3.3005
R97 drain_left.n31 drain_left.t0 3.3005
R98 drain_left.n64 drain_left.t3 3.3005
R99 drain_left.n64 drain_left.t2 3.3005
R100 drain_left.n20 drain_left.n19 2.71565
R101 drain_left.n53 drain_left.n52 2.71565
R102 drain_left.n16 drain_left.n6 1.93989
R103 drain_left.n49 drain_left.n39 1.93989
R104 drain_left.n15 drain_left.n8 1.16414
R105 drain_left.n48 drain_left.n41 1.16414
R106 drain_left.n12 drain_left.n11 0.388379
R107 drain_left.n45 drain_left.n44 0.388379
R108 drain_left.n14 drain_left.n13 0.155672
R109 drain_left.n14 drain_left.n5 0.155672
R110 drain_left.n21 drain_left.n5 0.155672
R111 drain_left.n22 drain_left.n21 0.155672
R112 drain_left.n22 drain_left.n1 0.155672
R113 drain_left.n29 drain_left.n1 0.155672
R114 drain_left.n62 drain_left.n34 0.155672
R115 drain_left.n55 drain_left.n34 0.155672
R116 drain_left.n55 drain_left.n54 0.155672
R117 drain_left.n54 drain_left.n38 0.155672
R118 drain_left.n47 drain_left.n38 0.155672
R119 drain_left.n47 drain_left.n46 0.155672
R120 source.n130 source.n104 289.615
R121 source.n96 source.n70 289.615
R122 source.n26 source.n0 289.615
R123 source.n60 source.n34 289.615
R124 source.n115 source.n114 185
R125 source.n112 source.n111 185
R126 source.n121 source.n120 185
R127 source.n123 source.n122 185
R128 source.n108 source.n107 185
R129 source.n129 source.n128 185
R130 source.n131 source.n130 185
R131 source.n81 source.n80 185
R132 source.n78 source.n77 185
R133 source.n87 source.n86 185
R134 source.n89 source.n88 185
R135 source.n74 source.n73 185
R136 source.n95 source.n94 185
R137 source.n97 source.n96 185
R138 source.n27 source.n26 185
R139 source.n25 source.n24 185
R140 source.n4 source.n3 185
R141 source.n19 source.n18 185
R142 source.n17 source.n16 185
R143 source.n8 source.n7 185
R144 source.n11 source.n10 185
R145 source.n61 source.n60 185
R146 source.n59 source.n58 185
R147 source.n38 source.n37 185
R148 source.n53 source.n52 185
R149 source.n51 source.n50 185
R150 source.n42 source.n41 185
R151 source.n45 source.n44 185
R152 source.t2 source.n113 147.661
R153 source.t6 source.n79 147.661
R154 source.t7 source.n9 147.661
R155 source.t4 source.n43 147.661
R156 source.n114 source.n111 104.615
R157 source.n121 source.n111 104.615
R158 source.n122 source.n121 104.615
R159 source.n122 source.n107 104.615
R160 source.n129 source.n107 104.615
R161 source.n130 source.n129 104.615
R162 source.n80 source.n77 104.615
R163 source.n87 source.n77 104.615
R164 source.n88 source.n87 104.615
R165 source.n88 source.n73 104.615
R166 source.n95 source.n73 104.615
R167 source.n96 source.n95 104.615
R168 source.n26 source.n25 104.615
R169 source.n25 source.n3 104.615
R170 source.n18 source.n3 104.615
R171 source.n18 source.n17 104.615
R172 source.n17 source.n7 104.615
R173 source.n10 source.n7 104.615
R174 source.n60 source.n59 104.615
R175 source.n59 source.n37 104.615
R176 source.n52 source.n37 104.615
R177 source.n52 source.n51 104.615
R178 source.n51 source.n41 104.615
R179 source.n44 source.n41 104.615
R180 source.n114 source.t2 52.3082
R181 source.n80 source.t6 52.3082
R182 source.n10 source.t7 52.3082
R183 source.n44 source.t4 52.3082
R184 source.n33 source.n32 50.512
R185 source.n67 source.n66 50.512
R186 source.n103 source.n102 50.5119
R187 source.n69 source.n68 50.5119
R188 source.n135 source.n134 32.1853
R189 source.n101 source.n100 32.1853
R190 source.n31 source.n30 32.1853
R191 source.n65 source.n64 32.1853
R192 source.n69 source.n67 17.7423
R193 source.n115 source.n113 15.6674
R194 source.n81 source.n79 15.6674
R195 source.n11 source.n9 15.6674
R196 source.n45 source.n43 15.6674
R197 source.n116 source.n112 12.8005
R198 source.n82 source.n78 12.8005
R199 source.n12 source.n8 12.8005
R200 source.n46 source.n42 12.8005
R201 source.n120 source.n119 12.0247
R202 source.n86 source.n85 12.0247
R203 source.n16 source.n15 12.0247
R204 source.n50 source.n49 12.0247
R205 source.n136 source.n31 11.7293
R206 source.n123 source.n110 11.249
R207 source.n89 source.n76 11.249
R208 source.n19 source.n6 11.249
R209 source.n53 source.n40 11.249
R210 source.n124 source.n108 10.4732
R211 source.n90 source.n74 10.4732
R212 source.n20 source.n4 10.4732
R213 source.n54 source.n38 10.4732
R214 source.n128 source.n127 9.69747
R215 source.n94 source.n93 9.69747
R216 source.n24 source.n23 9.69747
R217 source.n58 source.n57 9.69747
R218 source.n134 source.n133 9.45567
R219 source.n100 source.n99 9.45567
R220 source.n30 source.n29 9.45567
R221 source.n64 source.n63 9.45567
R222 source.n133 source.n132 9.3005
R223 source.n106 source.n105 9.3005
R224 source.n127 source.n126 9.3005
R225 source.n125 source.n124 9.3005
R226 source.n110 source.n109 9.3005
R227 source.n119 source.n118 9.3005
R228 source.n117 source.n116 9.3005
R229 source.n99 source.n98 9.3005
R230 source.n72 source.n71 9.3005
R231 source.n93 source.n92 9.3005
R232 source.n91 source.n90 9.3005
R233 source.n76 source.n75 9.3005
R234 source.n85 source.n84 9.3005
R235 source.n83 source.n82 9.3005
R236 source.n29 source.n28 9.3005
R237 source.n2 source.n1 9.3005
R238 source.n23 source.n22 9.3005
R239 source.n21 source.n20 9.3005
R240 source.n6 source.n5 9.3005
R241 source.n15 source.n14 9.3005
R242 source.n13 source.n12 9.3005
R243 source.n63 source.n62 9.3005
R244 source.n36 source.n35 9.3005
R245 source.n57 source.n56 9.3005
R246 source.n55 source.n54 9.3005
R247 source.n40 source.n39 9.3005
R248 source.n49 source.n48 9.3005
R249 source.n47 source.n46 9.3005
R250 source.n131 source.n106 8.92171
R251 source.n97 source.n72 8.92171
R252 source.n27 source.n2 8.92171
R253 source.n61 source.n36 8.92171
R254 source.n132 source.n104 8.14595
R255 source.n98 source.n70 8.14595
R256 source.n28 source.n0 8.14595
R257 source.n62 source.n34 8.14595
R258 source.n134 source.n104 5.81868
R259 source.n100 source.n70 5.81868
R260 source.n30 source.n0 5.81868
R261 source.n64 source.n34 5.81868
R262 source.n136 source.n135 5.51343
R263 source.n132 source.n131 5.04292
R264 source.n98 source.n97 5.04292
R265 source.n28 source.n27 5.04292
R266 source.n62 source.n61 5.04292
R267 source.n117 source.n113 4.38594
R268 source.n83 source.n79 4.38594
R269 source.n13 source.n9 4.38594
R270 source.n47 source.n43 4.38594
R271 source.n128 source.n106 4.26717
R272 source.n94 source.n72 4.26717
R273 source.n24 source.n2 4.26717
R274 source.n58 source.n36 4.26717
R275 source.n127 source.n108 3.49141
R276 source.n93 source.n74 3.49141
R277 source.n23 source.n4 3.49141
R278 source.n57 source.n38 3.49141
R279 source.n102 source.t1 3.3005
R280 source.n102 source.t3 3.3005
R281 source.n68 source.t10 3.3005
R282 source.n68 source.t8 3.3005
R283 source.n32 source.t9 3.3005
R284 source.n32 source.t11 3.3005
R285 source.n66 source.t5 3.3005
R286 source.n66 source.t0 3.3005
R287 source.n124 source.n123 2.71565
R288 source.n90 source.n89 2.71565
R289 source.n20 source.n19 2.71565
R290 source.n54 source.n53 2.71565
R291 source.n120 source.n110 1.93989
R292 source.n86 source.n76 1.93989
R293 source.n16 source.n6 1.93989
R294 source.n50 source.n40 1.93989
R295 source.n119 source.n112 1.16414
R296 source.n85 source.n78 1.16414
R297 source.n15 source.n8 1.16414
R298 source.n49 source.n42 1.16414
R299 source.n65 source.n33 0.720328
R300 source.n103 source.n101 0.720328
R301 source.n67 source.n65 0.5005
R302 source.n33 source.n31 0.5005
R303 source.n101 source.n69 0.5005
R304 source.n135 source.n103 0.5005
R305 source.n116 source.n115 0.388379
R306 source.n82 source.n81 0.388379
R307 source.n12 source.n11 0.388379
R308 source.n46 source.n45 0.388379
R309 source source.n136 0.188
R310 source.n118 source.n117 0.155672
R311 source.n118 source.n109 0.155672
R312 source.n125 source.n109 0.155672
R313 source.n126 source.n125 0.155672
R314 source.n126 source.n105 0.155672
R315 source.n133 source.n105 0.155672
R316 source.n84 source.n83 0.155672
R317 source.n84 source.n75 0.155672
R318 source.n91 source.n75 0.155672
R319 source.n92 source.n91 0.155672
R320 source.n92 source.n71 0.155672
R321 source.n99 source.n71 0.155672
R322 source.n29 source.n1 0.155672
R323 source.n22 source.n1 0.155672
R324 source.n22 source.n21 0.155672
R325 source.n21 source.n5 0.155672
R326 source.n14 source.n5 0.155672
R327 source.n14 source.n13 0.155672
R328 source.n63 source.n35 0.155672
R329 source.n56 source.n35 0.155672
R330 source.n56 source.n55 0.155672
R331 source.n55 source.n39 0.155672
R332 source.n48 source.n39 0.155672
R333 source.n48 source.n47 0.155672
R334 minus.n2 minus.t2 751.92
R335 minus.n0 minus.t4 751.92
R336 minus.n6 minus.t1 751.92
R337 minus.n4 minus.t3 751.92
R338 minus.n1 minus.t0 703.721
R339 minus.n5 minus.t5 703.721
R340 minus.n3 minus.n0 161.489
R341 minus.n7 minus.n4 161.489
R342 minus.n3 minus.n2 161.3
R343 minus.n7 minus.n6 161.3
R344 minus.n2 minus.n1 36.5157
R345 minus.n1 minus.n0 36.5157
R346 minus.n5 minus.n4 36.5157
R347 minus.n6 minus.n5 36.5157
R348 minus.n8 minus.n3 29.0308
R349 minus.n8 minus.n7 6.48535
R350 minus minus.n8 0.188
R351 drain_right.n26 drain_right.n0 289.615
R352 drain_right.n60 drain_right.n34 289.615
R353 drain_right.n11 drain_right.n10 185
R354 drain_right.n8 drain_right.n7 185
R355 drain_right.n17 drain_right.n16 185
R356 drain_right.n19 drain_right.n18 185
R357 drain_right.n4 drain_right.n3 185
R358 drain_right.n25 drain_right.n24 185
R359 drain_right.n27 drain_right.n26 185
R360 drain_right.n61 drain_right.n60 185
R361 drain_right.n59 drain_right.n58 185
R362 drain_right.n38 drain_right.n37 185
R363 drain_right.n53 drain_right.n52 185
R364 drain_right.n51 drain_right.n50 185
R365 drain_right.n42 drain_right.n41 185
R366 drain_right.n45 drain_right.n44 185
R367 drain_right.t2 drain_right.n9 147.661
R368 drain_right.t3 drain_right.n43 147.661
R369 drain_right.n10 drain_right.n7 104.615
R370 drain_right.n17 drain_right.n7 104.615
R371 drain_right.n18 drain_right.n17 104.615
R372 drain_right.n18 drain_right.n3 104.615
R373 drain_right.n25 drain_right.n3 104.615
R374 drain_right.n26 drain_right.n25 104.615
R375 drain_right.n60 drain_right.n59 104.615
R376 drain_right.n59 drain_right.n37 104.615
R377 drain_right.n52 drain_right.n37 104.615
R378 drain_right.n52 drain_right.n51 104.615
R379 drain_right.n51 drain_right.n41 104.615
R380 drain_right.n44 drain_right.n41 104.615
R381 drain_right.n65 drain_right.n33 67.6907
R382 drain_right.n32 drain_right.n31 67.2603
R383 drain_right.n10 drain_right.t2 52.3082
R384 drain_right.n44 drain_right.t3 52.3082
R385 drain_right.n32 drain_right.n30 49.1838
R386 drain_right.n65 drain_right.n64 48.8641
R387 drain_right drain_right.n32 23.6434
R388 drain_right.n11 drain_right.n9 15.6674
R389 drain_right.n45 drain_right.n43 15.6674
R390 drain_right.n12 drain_right.n8 12.8005
R391 drain_right.n46 drain_right.n42 12.8005
R392 drain_right.n16 drain_right.n15 12.0247
R393 drain_right.n50 drain_right.n49 12.0247
R394 drain_right.n19 drain_right.n6 11.249
R395 drain_right.n53 drain_right.n40 11.249
R396 drain_right.n20 drain_right.n4 10.4732
R397 drain_right.n54 drain_right.n38 10.4732
R398 drain_right.n24 drain_right.n23 9.69747
R399 drain_right.n58 drain_right.n57 9.69747
R400 drain_right.n30 drain_right.n29 9.45567
R401 drain_right.n64 drain_right.n63 9.45567
R402 drain_right.n29 drain_right.n28 9.3005
R403 drain_right.n2 drain_right.n1 9.3005
R404 drain_right.n23 drain_right.n22 9.3005
R405 drain_right.n21 drain_right.n20 9.3005
R406 drain_right.n6 drain_right.n5 9.3005
R407 drain_right.n15 drain_right.n14 9.3005
R408 drain_right.n13 drain_right.n12 9.3005
R409 drain_right.n63 drain_right.n62 9.3005
R410 drain_right.n36 drain_right.n35 9.3005
R411 drain_right.n57 drain_right.n56 9.3005
R412 drain_right.n55 drain_right.n54 9.3005
R413 drain_right.n40 drain_right.n39 9.3005
R414 drain_right.n49 drain_right.n48 9.3005
R415 drain_right.n47 drain_right.n46 9.3005
R416 drain_right.n27 drain_right.n2 8.92171
R417 drain_right.n61 drain_right.n36 8.92171
R418 drain_right.n28 drain_right.n0 8.14595
R419 drain_right.n62 drain_right.n34 8.14595
R420 drain_right drain_right.n65 5.90322
R421 drain_right.n30 drain_right.n0 5.81868
R422 drain_right.n64 drain_right.n34 5.81868
R423 drain_right.n28 drain_right.n27 5.04292
R424 drain_right.n62 drain_right.n61 5.04292
R425 drain_right.n13 drain_right.n9 4.38594
R426 drain_right.n47 drain_right.n43 4.38594
R427 drain_right.n24 drain_right.n2 4.26717
R428 drain_right.n58 drain_right.n36 4.26717
R429 drain_right.n23 drain_right.n4 3.49141
R430 drain_right.n57 drain_right.n38 3.49141
R431 drain_right.n31 drain_right.t0 3.3005
R432 drain_right.n31 drain_right.t4 3.3005
R433 drain_right.n33 drain_right.t5 3.3005
R434 drain_right.n33 drain_right.t1 3.3005
R435 drain_right.n20 drain_right.n19 2.71565
R436 drain_right.n54 drain_right.n53 2.71565
R437 drain_right.n16 drain_right.n6 1.93989
R438 drain_right.n50 drain_right.n40 1.93989
R439 drain_right.n15 drain_right.n8 1.16414
R440 drain_right.n49 drain_right.n42 1.16414
R441 drain_right.n12 drain_right.n11 0.388379
R442 drain_right.n46 drain_right.n45 0.388379
R443 drain_right.n14 drain_right.n13 0.155672
R444 drain_right.n14 drain_right.n5 0.155672
R445 drain_right.n21 drain_right.n5 0.155672
R446 drain_right.n22 drain_right.n21 0.155672
R447 drain_right.n22 drain_right.n1 0.155672
R448 drain_right.n29 drain_right.n1 0.155672
R449 drain_right.n63 drain_right.n35 0.155672
R450 drain_right.n56 drain_right.n35 0.155672
R451 drain_right.n56 drain_right.n55 0.155672
R452 drain_right.n55 drain_right.n39 0.155672
R453 drain_right.n48 drain_right.n39 0.155672
R454 drain_right.n48 drain_right.n47 0.155672
C0 drain_right plus 0.264418f
C1 drain_left minus 0.170597f
C2 drain_left source 8.3689f
C3 drain_right minus 1.38515f
C4 source drain_right 8.361629f
C5 drain_left drain_right 0.549358f
C6 minus plus 3.51111f
C7 source plus 1.20902f
C8 drain_left plus 1.4937f
C9 source minus 1.19467f
C10 drain_right a_n1180_n2088# 4.31461f
C11 drain_left a_n1180_n2088# 4.47271f
C12 source a_n1180_n2088# 3.79786f
C13 minus a_n1180_n2088# 4.04558f
C14 plus a_n1180_n2088# 4.89948f
C15 drain_right.n0 a_n1180_n2088# 0.034269f
C16 drain_right.n1 a_n1180_n2088# 0.02438f
C17 drain_right.n2 a_n1180_n2088# 0.013101f
C18 drain_right.n3 a_n1180_n2088# 0.030966f
C19 drain_right.n4 a_n1180_n2088# 0.013872f
C20 drain_right.n5 a_n1180_n2088# 0.02438f
C21 drain_right.n6 a_n1180_n2088# 0.013101f
C22 drain_right.n7 a_n1180_n2088# 0.030966f
C23 drain_right.n8 a_n1180_n2088# 0.013872f
C24 drain_right.n9 a_n1180_n2088# 0.10433f
C25 drain_right.t2 a_n1180_n2088# 0.05047f
C26 drain_right.n10 a_n1180_n2088# 0.023224f
C27 drain_right.n11 a_n1180_n2088# 0.018291f
C28 drain_right.n12 a_n1180_n2088# 0.013101f
C29 drain_right.n13 a_n1180_n2088# 0.580104f
C30 drain_right.n14 a_n1180_n2088# 0.02438f
C31 drain_right.n15 a_n1180_n2088# 0.013101f
C32 drain_right.n16 a_n1180_n2088# 0.013872f
C33 drain_right.n17 a_n1180_n2088# 0.030966f
C34 drain_right.n18 a_n1180_n2088# 0.030966f
C35 drain_right.n19 a_n1180_n2088# 0.013872f
C36 drain_right.n20 a_n1180_n2088# 0.013101f
C37 drain_right.n21 a_n1180_n2088# 0.02438f
C38 drain_right.n22 a_n1180_n2088# 0.02438f
C39 drain_right.n23 a_n1180_n2088# 0.013101f
C40 drain_right.n24 a_n1180_n2088# 0.013872f
C41 drain_right.n25 a_n1180_n2088# 0.030966f
C42 drain_right.n26 a_n1180_n2088# 0.067035f
C43 drain_right.n27 a_n1180_n2088# 0.013872f
C44 drain_right.n28 a_n1180_n2088# 0.013101f
C45 drain_right.n29 a_n1180_n2088# 0.056354f
C46 drain_right.n30 a_n1180_n2088# 0.054823f
C47 drain_right.t0 a_n1180_n2088# 0.115596f
C48 drain_right.t4 a_n1180_n2088# 0.115596f
C49 drain_right.n31 a_n1180_n2088# 0.964341f
C50 drain_right.n32 a_n1180_n2088# 0.98745f
C51 drain_right.t5 a_n1180_n2088# 0.115596f
C52 drain_right.t1 a_n1180_n2088# 0.115596f
C53 drain_right.n33 a_n1180_n2088# 0.966186f
C54 drain_right.n34 a_n1180_n2088# 0.034269f
C55 drain_right.n35 a_n1180_n2088# 0.02438f
C56 drain_right.n36 a_n1180_n2088# 0.013101f
C57 drain_right.n37 a_n1180_n2088# 0.030966f
C58 drain_right.n38 a_n1180_n2088# 0.013872f
C59 drain_right.n39 a_n1180_n2088# 0.02438f
C60 drain_right.n40 a_n1180_n2088# 0.013101f
C61 drain_right.n41 a_n1180_n2088# 0.030966f
C62 drain_right.n42 a_n1180_n2088# 0.013872f
C63 drain_right.n43 a_n1180_n2088# 0.10433f
C64 drain_right.t3 a_n1180_n2088# 0.05047f
C65 drain_right.n44 a_n1180_n2088# 0.023224f
C66 drain_right.n45 a_n1180_n2088# 0.018291f
C67 drain_right.n46 a_n1180_n2088# 0.013101f
C68 drain_right.n47 a_n1180_n2088# 0.580104f
C69 drain_right.n48 a_n1180_n2088# 0.02438f
C70 drain_right.n49 a_n1180_n2088# 0.013101f
C71 drain_right.n50 a_n1180_n2088# 0.013872f
C72 drain_right.n51 a_n1180_n2088# 0.030966f
C73 drain_right.n52 a_n1180_n2088# 0.030966f
C74 drain_right.n53 a_n1180_n2088# 0.013872f
C75 drain_right.n54 a_n1180_n2088# 0.013101f
C76 drain_right.n55 a_n1180_n2088# 0.02438f
C77 drain_right.n56 a_n1180_n2088# 0.02438f
C78 drain_right.n57 a_n1180_n2088# 0.013101f
C79 drain_right.n58 a_n1180_n2088# 0.013872f
C80 drain_right.n59 a_n1180_n2088# 0.030966f
C81 drain_right.n60 a_n1180_n2088# 0.067035f
C82 drain_right.n61 a_n1180_n2088# 0.013872f
C83 drain_right.n62 a_n1180_n2088# 0.013101f
C84 drain_right.n63 a_n1180_n2088# 0.056354f
C85 drain_right.n64 a_n1180_n2088# 0.054343f
C86 drain_right.n65 a_n1180_n2088# 0.571145f
C87 minus.t4 a_n1180_n2088# 0.14821f
C88 minus.n0 a_n1180_n2088# 0.077797f
C89 minus.t2 a_n1180_n2088# 0.14821f
C90 minus.t0 a_n1180_n2088# 0.143763f
C91 minus.n1 a_n1180_n2088# 0.067718f
C92 minus.n2 a_n1180_n2088# 0.077748f
C93 minus.n3 a_n1180_n2088# 0.868584f
C94 minus.t3 a_n1180_n2088# 0.14821f
C95 minus.n4 a_n1180_n2088# 0.077797f
C96 minus.t5 a_n1180_n2088# 0.143763f
C97 minus.n5 a_n1180_n2088# 0.067718f
C98 minus.t1 a_n1180_n2088# 0.14821f
C99 minus.n6 a_n1180_n2088# 0.077748f
C100 minus.n7 a_n1180_n2088# 0.26085f
C101 minus.n8 a_n1180_n2088# 1.02158f
C102 source.n0 a_n1180_n2088# 0.037767f
C103 source.n1 a_n1180_n2088# 0.026869f
C104 source.n2 a_n1180_n2088# 0.014438f
C105 source.n3 a_n1180_n2088# 0.034127f
C106 source.n4 a_n1180_n2088# 0.015288f
C107 source.n5 a_n1180_n2088# 0.026869f
C108 source.n6 a_n1180_n2088# 0.014438f
C109 source.n7 a_n1180_n2088# 0.034127f
C110 source.n8 a_n1180_n2088# 0.015288f
C111 source.n9 a_n1180_n2088# 0.114981f
C112 source.t7 a_n1180_n2088# 0.055622f
C113 source.n10 a_n1180_n2088# 0.025595f
C114 source.n11 a_n1180_n2088# 0.020158f
C115 source.n12 a_n1180_n2088# 0.014438f
C116 source.n13 a_n1180_n2088# 0.639325f
C117 source.n14 a_n1180_n2088# 0.026869f
C118 source.n15 a_n1180_n2088# 0.014438f
C119 source.n16 a_n1180_n2088# 0.015288f
C120 source.n17 a_n1180_n2088# 0.034127f
C121 source.n18 a_n1180_n2088# 0.034127f
C122 source.n19 a_n1180_n2088# 0.015288f
C123 source.n20 a_n1180_n2088# 0.014438f
C124 source.n21 a_n1180_n2088# 0.026869f
C125 source.n22 a_n1180_n2088# 0.026869f
C126 source.n23 a_n1180_n2088# 0.014438f
C127 source.n24 a_n1180_n2088# 0.015288f
C128 source.n25 a_n1180_n2088# 0.034127f
C129 source.n26 a_n1180_n2088# 0.073879f
C130 source.n27 a_n1180_n2088# 0.015288f
C131 source.n28 a_n1180_n2088# 0.014438f
C132 source.n29 a_n1180_n2088# 0.062107f
C133 source.n30 a_n1180_n2088# 0.041338f
C134 source.n31 a_n1180_n2088# 0.644424f
C135 source.t9 a_n1180_n2088# 0.127397f
C136 source.t11 a_n1180_n2088# 0.127397f
C137 source.n32 a_n1180_n2088# 0.992176f
C138 source.n33 a_n1180_n2088# 0.357483f
C139 source.n34 a_n1180_n2088# 0.037767f
C140 source.n35 a_n1180_n2088# 0.026869f
C141 source.n36 a_n1180_n2088# 0.014438f
C142 source.n37 a_n1180_n2088# 0.034127f
C143 source.n38 a_n1180_n2088# 0.015288f
C144 source.n39 a_n1180_n2088# 0.026869f
C145 source.n40 a_n1180_n2088# 0.014438f
C146 source.n41 a_n1180_n2088# 0.034127f
C147 source.n42 a_n1180_n2088# 0.015288f
C148 source.n43 a_n1180_n2088# 0.114981f
C149 source.t4 a_n1180_n2088# 0.055622f
C150 source.n44 a_n1180_n2088# 0.025595f
C151 source.n45 a_n1180_n2088# 0.020158f
C152 source.n46 a_n1180_n2088# 0.014438f
C153 source.n47 a_n1180_n2088# 0.639325f
C154 source.n48 a_n1180_n2088# 0.026869f
C155 source.n49 a_n1180_n2088# 0.014438f
C156 source.n50 a_n1180_n2088# 0.015288f
C157 source.n51 a_n1180_n2088# 0.034127f
C158 source.n52 a_n1180_n2088# 0.034127f
C159 source.n53 a_n1180_n2088# 0.015288f
C160 source.n54 a_n1180_n2088# 0.014438f
C161 source.n55 a_n1180_n2088# 0.026869f
C162 source.n56 a_n1180_n2088# 0.026869f
C163 source.n57 a_n1180_n2088# 0.014438f
C164 source.n58 a_n1180_n2088# 0.015288f
C165 source.n59 a_n1180_n2088# 0.034127f
C166 source.n60 a_n1180_n2088# 0.073879f
C167 source.n61 a_n1180_n2088# 0.015288f
C168 source.n62 a_n1180_n2088# 0.014438f
C169 source.n63 a_n1180_n2088# 0.062107f
C170 source.n64 a_n1180_n2088# 0.041338f
C171 source.n65 a_n1180_n2088# 0.128559f
C172 source.t5 a_n1180_n2088# 0.127397f
C173 source.t0 a_n1180_n2088# 0.127397f
C174 source.n66 a_n1180_n2088# 0.992176f
C175 source.n67 a_n1180_n2088# 1.26148f
C176 source.t10 a_n1180_n2088# 0.127397f
C177 source.t8 a_n1180_n2088# 0.127397f
C178 source.n68 a_n1180_n2088# 0.992169f
C179 source.n69 a_n1180_n2088# 1.26149f
C180 source.n70 a_n1180_n2088# 0.037767f
C181 source.n71 a_n1180_n2088# 0.026869f
C182 source.n72 a_n1180_n2088# 0.014438f
C183 source.n73 a_n1180_n2088# 0.034127f
C184 source.n74 a_n1180_n2088# 0.015288f
C185 source.n75 a_n1180_n2088# 0.026869f
C186 source.n76 a_n1180_n2088# 0.014438f
C187 source.n77 a_n1180_n2088# 0.034127f
C188 source.n78 a_n1180_n2088# 0.015288f
C189 source.n79 a_n1180_n2088# 0.114981f
C190 source.t6 a_n1180_n2088# 0.055622f
C191 source.n80 a_n1180_n2088# 0.025595f
C192 source.n81 a_n1180_n2088# 0.020158f
C193 source.n82 a_n1180_n2088# 0.014438f
C194 source.n83 a_n1180_n2088# 0.639325f
C195 source.n84 a_n1180_n2088# 0.026869f
C196 source.n85 a_n1180_n2088# 0.014438f
C197 source.n86 a_n1180_n2088# 0.015288f
C198 source.n87 a_n1180_n2088# 0.034127f
C199 source.n88 a_n1180_n2088# 0.034127f
C200 source.n89 a_n1180_n2088# 0.015288f
C201 source.n90 a_n1180_n2088# 0.014438f
C202 source.n91 a_n1180_n2088# 0.026869f
C203 source.n92 a_n1180_n2088# 0.026869f
C204 source.n93 a_n1180_n2088# 0.014438f
C205 source.n94 a_n1180_n2088# 0.015288f
C206 source.n95 a_n1180_n2088# 0.034127f
C207 source.n96 a_n1180_n2088# 0.073879f
C208 source.n97 a_n1180_n2088# 0.015288f
C209 source.n98 a_n1180_n2088# 0.014438f
C210 source.n99 a_n1180_n2088# 0.062107f
C211 source.n100 a_n1180_n2088# 0.041338f
C212 source.n101 a_n1180_n2088# 0.128559f
C213 source.t1 a_n1180_n2088# 0.127397f
C214 source.t3 a_n1180_n2088# 0.127397f
C215 source.n102 a_n1180_n2088# 0.992169f
C216 source.n103 a_n1180_n2088# 0.35749f
C217 source.n104 a_n1180_n2088# 0.037767f
C218 source.n105 a_n1180_n2088# 0.026869f
C219 source.n106 a_n1180_n2088# 0.014438f
C220 source.n107 a_n1180_n2088# 0.034127f
C221 source.n108 a_n1180_n2088# 0.015288f
C222 source.n109 a_n1180_n2088# 0.026869f
C223 source.n110 a_n1180_n2088# 0.014438f
C224 source.n111 a_n1180_n2088# 0.034127f
C225 source.n112 a_n1180_n2088# 0.015288f
C226 source.n113 a_n1180_n2088# 0.114981f
C227 source.t2 a_n1180_n2088# 0.055622f
C228 source.n114 a_n1180_n2088# 0.025595f
C229 source.n115 a_n1180_n2088# 0.020158f
C230 source.n116 a_n1180_n2088# 0.014438f
C231 source.n117 a_n1180_n2088# 0.639325f
C232 source.n118 a_n1180_n2088# 0.026869f
C233 source.n119 a_n1180_n2088# 0.014438f
C234 source.n120 a_n1180_n2088# 0.015288f
C235 source.n121 a_n1180_n2088# 0.034127f
C236 source.n122 a_n1180_n2088# 0.034127f
C237 source.n123 a_n1180_n2088# 0.015288f
C238 source.n124 a_n1180_n2088# 0.014438f
C239 source.n125 a_n1180_n2088# 0.026869f
C240 source.n126 a_n1180_n2088# 0.026869f
C241 source.n127 a_n1180_n2088# 0.014438f
C242 source.n128 a_n1180_n2088# 0.015288f
C243 source.n129 a_n1180_n2088# 0.034127f
C244 source.n130 a_n1180_n2088# 0.073879f
C245 source.n131 a_n1180_n2088# 0.015288f
C246 source.n132 a_n1180_n2088# 0.014438f
C247 source.n133 a_n1180_n2088# 0.062107f
C248 source.n134 a_n1180_n2088# 0.041338f
C249 source.n135 a_n1180_n2088# 0.255603f
C250 source.n136 a_n1180_n2088# 1.09763f
C251 drain_left.n0 a_n1180_n2088# 0.033884f
C252 drain_left.n1 a_n1180_n2088# 0.024107f
C253 drain_left.n2 a_n1180_n2088# 0.012954f
C254 drain_left.n3 a_n1180_n2088# 0.030618f
C255 drain_left.n4 a_n1180_n2088# 0.013716f
C256 drain_left.n5 a_n1180_n2088# 0.024107f
C257 drain_left.n6 a_n1180_n2088# 0.012954f
C258 drain_left.n7 a_n1180_n2088# 0.030618f
C259 drain_left.n8 a_n1180_n2088# 0.013716f
C260 drain_left.n9 a_n1180_n2088# 0.103159f
C261 drain_left.t1 a_n1180_n2088# 0.049903f
C262 drain_left.n10 a_n1180_n2088# 0.022964f
C263 drain_left.n11 a_n1180_n2088# 0.018086f
C264 drain_left.n12 a_n1180_n2088# 0.012954f
C265 drain_left.n13 a_n1180_n2088# 0.573592f
C266 drain_left.n14 a_n1180_n2088# 0.024107f
C267 drain_left.n15 a_n1180_n2088# 0.012954f
C268 drain_left.n16 a_n1180_n2088# 0.013716f
C269 drain_left.n17 a_n1180_n2088# 0.030618f
C270 drain_left.n18 a_n1180_n2088# 0.030618f
C271 drain_left.n19 a_n1180_n2088# 0.013716f
C272 drain_left.n20 a_n1180_n2088# 0.012954f
C273 drain_left.n21 a_n1180_n2088# 0.024107f
C274 drain_left.n22 a_n1180_n2088# 0.024107f
C275 drain_left.n23 a_n1180_n2088# 0.012954f
C276 drain_left.n24 a_n1180_n2088# 0.013716f
C277 drain_left.n25 a_n1180_n2088# 0.030618f
C278 drain_left.n26 a_n1180_n2088# 0.066283f
C279 drain_left.n27 a_n1180_n2088# 0.013716f
C280 drain_left.n28 a_n1180_n2088# 0.012954f
C281 drain_left.n29 a_n1180_n2088# 0.055721f
C282 drain_left.n30 a_n1180_n2088# 0.054207f
C283 drain_left.t5 a_n1180_n2088# 0.114298f
C284 drain_left.t0 a_n1180_n2088# 0.114298f
C285 drain_left.n31 a_n1180_n2088# 0.953515f
C286 drain_left.n32 a_n1180_n2088# 1.02587f
C287 drain_left.n33 a_n1180_n2088# 0.033884f
C288 drain_left.n34 a_n1180_n2088# 0.024107f
C289 drain_left.n35 a_n1180_n2088# 0.012954f
C290 drain_left.n36 a_n1180_n2088# 0.030618f
C291 drain_left.n37 a_n1180_n2088# 0.013716f
C292 drain_left.n38 a_n1180_n2088# 0.024107f
C293 drain_left.n39 a_n1180_n2088# 0.012954f
C294 drain_left.n40 a_n1180_n2088# 0.030618f
C295 drain_left.n41 a_n1180_n2088# 0.013716f
C296 drain_left.n42 a_n1180_n2088# 0.103159f
C297 drain_left.t4 a_n1180_n2088# 0.049903f
C298 drain_left.n43 a_n1180_n2088# 0.022964f
C299 drain_left.n44 a_n1180_n2088# 0.018086f
C300 drain_left.n45 a_n1180_n2088# 0.012954f
C301 drain_left.n46 a_n1180_n2088# 0.573592f
C302 drain_left.n47 a_n1180_n2088# 0.024107f
C303 drain_left.n48 a_n1180_n2088# 0.012954f
C304 drain_left.n49 a_n1180_n2088# 0.013716f
C305 drain_left.n50 a_n1180_n2088# 0.030618f
C306 drain_left.n51 a_n1180_n2088# 0.030618f
C307 drain_left.n52 a_n1180_n2088# 0.013716f
C308 drain_left.n53 a_n1180_n2088# 0.012954f
C309 drain_left.n54 a_n1180_n2088# 0.024107f
C310 drain_left.n55 a_n1180_n2088# 0.024107f
C311 drain_left.n56 a_n1180_n2088# 0.012954f
C312 drain_left.n57 a_n1180_n2088# 0.013716f
C313 drain_left.n58 a_n1180_n2088# 0.030618f
C314 drain_left.n59 a_n1180_n2088# 0.066283f
C315 drain_left.n60 a_n1180_n2088# 0.013716f
C316 drain_left.n61 a_n1180_n2088# 0.012954f
C317 drain_left.n62 a_n1180_n2088# 0.055721f
C318 drain_left.n63 a_n1180_n2088# 0.054596f
C319 drain_left.t3 a_n1180_n2088# 0.114298f
C320 drain_left.t2 a_n1180_n2088# 0.114298f
C321 drain_left.n64 a_n1180_n2088# 0.953248f
C322 drain_left.n65 a_n1180_n2088# 0.55671f
C323 plus.t2 a_n1180_n2088# 0.151148f
C324 plus.n0 a_n1180_n2088# 0.079339f
C325 plus.t0 a_n1180_n2088# 0.146613f
C326 plus.n1 a_n1180_n2088# 0.06906f
C327 plus.t4 a_n1180_n2088# 0.151148f
C328 plus.n2 a_n1180_n2088# 0.079289f
C329 plus.n3 a_n1180_n2088# 0.335651f
C330 plus.t5 a_n1180_n2088# 0.151148f
C331 plus.n4 a_n1180_n2088# 0.079339f
C332 plus.t1 a_n1180_n2088# 0.151148f
C333 plus.t3 a_n1180_n2088# 0.146613f
C334 plus.n5 a_n1180_n2088# 0.06906f
C335 plus.n6 a_n1180_n2088# 0.079289f
C336 plus.n7 a_n1180_n2088# 0.80581f
.ends

