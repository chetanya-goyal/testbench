* NGSPICE file created from diffpair313.ext - technology: sky130A

.subckt diffpair313 minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t7 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X1 drain_right.t7 minus.t0 source.t7 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X3 a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X4 drain_left.t1 plus.t1 source.t14 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X5 a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X6 source.t5 minus.t1 drain_right.t6 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X7 a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X8 drain_right.t5 minus.t2 source.t0 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X9 drain_left.t4 plus.t2 source.t13 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X10 source.t4 minus.t3 drain_right.t4 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X11 source.t2 minus.t4 drain_right.t3 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X12 drain_right.t2 minus.t5 source.t1 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X13 source.t3 minus.t6 drain_right.t1 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X14 drain_left.t5 plus.t3 source.t12 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X15 source.t11 plus.t4 drain_left.t3 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X16 drain_left.t0 plus.t5 source.t10 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X17 source.t9 plus.t6 drain_left.t2 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X18 drain_right.t0 minus.t7 source.t6 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X19 source.t8 plus.t7 drain_left.t6 a_n1846_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
R0 plus.n2 plus.t6 250.457
R1 plus.n10 plus.t2 250.457
R2 plus.n6 plus.t3 229.855
R3 plus.n4 plus.t4 229.855
R4 plus.n3 plus.t5 229.855
R5 plus.n14 plus.t7 229.855
R6 plus.n12 plus.t1 229.855
R7 plus.n11 plus.t0 229.855
R8 plus.n5 plus.n0 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n13 plus.n8 161.3
R11 plus.n15 plus.n14 161.3
R12 plus.n4 plus.n1 80.6037
R13 plus.n12 plus.n9 80.6037
R14 plus.n4 plus.n3 48.2005
R15 plus.n12 plus.n11 48.2005
R16 plus.n5 plus.n4 41.6278
R17 plus.n13 plus.n12 41.6278
R18 plus.n2 plus.n1 31.6158
R19 plus.n10 plus.n9 31.6158
R20 plus plus.n15 27.874
R21 plus.n3 plus.n2 17.6494
R22 plus.n11 plus.n10 17.6494
R23 plus plus.n7 10.0232
R24 plus.n6 plus.n5 6.57323
R25 plus.n14 plus.n13 6.57323
R26 plus.n1 plus.n0 0.285035
R27 plus.n9 plus.n8 0.285035
R28 plus.n7 plus.n0 0.189894
R29 plus.n15 plus.n8 0.189894
R30 drain_left.n5 drain_left.n3 68.165
R31 drain_left.n2 drain_left.n1 67.6224
R32 drain_left.n2 drain_left.n0 67.6224
R33 drain_left.n5 drain_left.n4 67.1907
R34 drain_left drain_left.n2 26.2311
R35 drain_left drain_left.n5 6.62735
R36 drain_left.n1 drain_left.t7 3.3005
R37 drain_left.n1 drain_left.t4 3.3005
R38 drain_left.n0 drain_left.t6 3.3005
R39 drain_left.n0 drain_left.t1 3.3005
R40 drain_left.n4 drain_left.t3 3.3005
R41 drain_left.n4 drain_left.t5 3.3005
R42 drain_left.n3 drain_left.t2 3.3005
R43 drain_left.n3 drain_left.t0 3.3005
R44 source.n258 source.n232 289.615
R45 source.n224 source.n198 289.615
R46 source.n192 source.n166 289.615
R47 source.n158 source.n132 289.615
R48 source.n26 source.n0 289.615
R49 source.n60 source.n34 289.615
R50 source.n92 source.n66 289.615
R51 source.n126 source.n100 289.615
R52 source.n243 source.n242 185
R53 source.n240 source.n239 185
R54 source.n249 source.n248 185
R55 source.n251 source.n250 185
R56 source.n236 source.n235 185
R57 source.n257 source.n256 185
R58 source.n259 source.n258 185
R59 source.n209 source.n208 185
R60 source.n206 source.n205 185
R61 source.n215 source.n214 185
R62 source.n217 source.n216 185
R63 source.n202 source.n201 185
R64 source.n223 source.n222 185
R65 source.n225 source.n224 185
R66 source.n177 source.n176 185
R67 source.n174 source.n173 185
R68 source.n183 source.n182 185
R69 source.n185 source.n184 185
R70 source.n170 source.n169 185
R71 source.n191 source.n190 185
R72 source.n193 source.n192 185
R73 source.n143 source.n142 185
R74 source.n140 source.n139 185
R75 source.n149 source.n148 185
R76 source.n151 source.n150 185
R77 source.n136 source.n135 185
R78 source.n157 source.n156 185
R79 source.n159 source.n158 185
R80 source.n27 source.n26 185
R81 source.n25 source.n24 185
R82 source.n4 source.n3 185
R83 source.n19 source.n18 185
R84 source.n17 source.n16 185
R85 source.n8 source.n7 185
R86 source.n11 source.n10 185
R87 source.n61 source.n60 185
R88 source.n59 source.n58 185
R89 source.n38 source.n37 185
R90 source.n53 source.n52 185
R91 source.n51 source.n50 185
R92 source.n42 source.n41 185
R93 source.n45 source.n44 185
R94 source.n93 source.n92 185
R95 source.n91 source.n90 185
R96 source.n70 source.n69 185
R97 source.n85 source.n84 185
R98 source.n83 source.n82 185
R99 source.n74 source.n73 185
R100 source.n77 source.n76 185
R101 source.n127 source.n126 185
R102 source.n125 source.n124 185
R103 source.n104 source.n103 185
R104 source.n119 source.n118 185
R105 source.n117 source.n116 185
R106 source.n108 source.n107 185
R107 source.n111 source.n110 185
R108 source.t6 source.n241 147.661
R109 source.t2 source.n207 147.661
R110 source.t13 source.n175 147.661
R111 source.t8 source.n141 147.661
R112 source.t12 source.n9 147.661
R113 source.t9 source.n43 147.661
R114 source.t1 source.n75 147.661
R115 source.t3 source.n109 147.661
R116 source.n242 source.n239 104.615
R117 source.n249 source.n239 104.615
R118 source.n250 source.n249 104.615
R119 source.n250 source.n235 104.615
R120 source.n257 source.n235 104.615
R121 source.n258 source.n257 104.615
R122 source.n208 source.n205 104.615
R123 source.n215 source.n205 104.615
R124 source.n216 source.n215 104.615
R125 source.n216 source.n201 104.615
R126 source.n223 source.n201 104.615
R127 source.n224 source.n223 104.615
R128 source.n176 source.n173 104.615
R129 source.n183 source.n173 104.615
R130 source.n184 source.n183 104.615
R131 source.n184 source.n169 104.615
R132 source.n191 source.n169 104.615
R133 source.n192 source.n191 104.615
R134 source.n142 source.n139 104.615
R135 source.n149 source.n139 104.615
R136 source.n150 source.n149 104.615
R137 source.n150 source.n135 104.615
R138 source.n157 source.n135 104.615
R139 source.n158 source.n157 104.615
R140 source.n26 source.n25 104.615
R141 source.n25 source.n3 104.615
R142 source.n18 source.n3 104.615
R143 source.n18 source.n17 104.615
R144 source.n17 source.n7 104.615
R145 source.n10 source.n7 104.615
R146 source.n60 source.n59 104.615
R147 source.n59 source.n37 104.615
R148 source.n52 source.n37 104.615
R149 source.n52 source.n51 104.615
R150 source.n51 source.n41 104.615
R151 source.n44 source.n41 104.615
R152 source.n92 source.n91 104.615
R153 source.n91 source.n69 104.615
R154 source.n84 source.n69 104.615
R155 source.n84 source.n83 104.615
R156 source.n83 source.n73 104.615
R157 source.n76 source.n73 104.615
R158 source.n126 source.n125 104.615
R159 source.n125 source.n103 104.615
R160 source.n118 source.n103 104.615
R161 source.n118 source.n117 104.615
R162 source.n117 source.n107 104.615
R163 source.n110 source.n107 104.615
R164 source.n242 source.t6 52.3082
R165 source.n208 source.t2 52.3082
R166 source.n176 source.t13 52.3082
R167 source.n142 source.t8 52.3082
R168 source.n10 source.t12 52.3082
R169 source.n44 source.t9 52.3082
R170 source.n76 source.t1 52.3082
R171 source.n110 source.t3 52.3082
R172 source.n33 source.n32 50.512
R173 source.n99 source.n98 50.512
R174 source.n231 source.n230 50.5119
R175 source.n165 source.n164 50.5119
R176 source.n263 source.n262 32.1853
R177 source.n229 source.n228 32.1853
R178 source.n197 source.n196 32.1853
R179 source.n163 source.n162 32.1853
R180 source.n31 source.n30 32.1853
R181 source.n65 source.n64 32.1853
R182 source.n97 source.n96 32.1853
R183 source.n131 source.n130 32.1853
R184 source.n163 source.n131 17.7164
R185 source.n243 source.n241 15.6674
R186 source.n209 source.n207 15.6674
R187 source.n177 source.n175 15.6674
R188 source.n143 source.n141 15.6674
R189 source.n11 source.n9 15.6674
R190 source.n45 source.n43 15.6674
R191 source.n77 source.n75 15.6674
R192 source.n111 source.n109 15.6674
R193 source.n244 source.n240 12.8005
R194 source.n210 source.n206 12.8005
R195 source.n178 source.n174 12.8005
R196 source.n144 source.n140 12.8005
R197 source.n12 source.n8 12.8005
R198 source.n46 source.n42 12.8005
R199 source.n78 source.n74 12.8005
R200 source.n112 source.n108 12.8005
R201 source.n248 source.n247 12.0247
R202 source.n214 source.n213 12.0247
R203 source.n182 source.n181 12.0247
R204 source.n148 source.n147 12.0247
R205 source.n16 source.n15 12.0247
R206 source.n50 source.n49 12.0247
R207 source.n82 source.n81 12.0247
R208 source.n116 source.n115 12.0247
R209 source.n264 source.n31 11.9664
R210 source.n251 source.n238 11.249
R211 source.n217 source.n204 11.249
R212 source.n185 source.n172 11.249
R213 source.n151 source.n138 11.249
R214 source.n19 source.n6 11.249
R215 source.n53 source.n40 11.249
R216 source.n85 source.n72 11.249
R217 source.n119 source.n106 11.249
R218 source.n252 source.n236 10.4732
R219 source.n218 source.n202 10.4732
R220 source.n186 source.n170 10.4732
R221 source.n152 source.n136 10.4732
R222 source.n20 source.n4 10.4732
R223 source.n54 source.n38 10.4732
R224 source.n86 source.n70 10.4732
R225 source.n120 source.n104 10.4732
R226 source.n256 source.n255 9.69747
R227 source.n222 source.n221 9.69747
R228 source.n190 source.n189 9.69747
R229 source.n156 source.n155 9.69747
R230 source.n24 source.n23 9.69747
R231 source.n58 source.n57 9.69747
R232 source.n90 source.n89 9.69747
R233 source.n124 source.n123 9.69747
R234 source.n262 source.n261 9.45567
R235 source.n228 source.n227 9.45567
R236 source.n196 source.n195 9.45567
R237 source.n162 source.n161 9.45567
R238 source.n30 source.n29 9.45567
R239 source.n64 source.n63 9.45567
R240 source.n96 source.n95 9.45567
R241 source.n130 source.n129 9.45567
R242 source.n261 source.n260 9.3005
R243 source.n234 source.n233 9.3005
R244 source.n255 source.n254 9.3005
R245 source.n253 source.n252 9.3005
R246 source.n238 source.n237 9.3005
R247 source.n247 source.n246 9.3005
R248 source.n245 source.n244 9.3005
R249 source.n227 source.n226 9.3005
R250 source.n200 source.n199 9.3005
R251 source.n221 source.n220 9.3005
R252 source.n219 source.n218 9.3005
R253 source.n204 source.n203 9.3005
R254 source.n213 source.n212 9.3005
R255 source.n211 source.n210 9.3005
R256 source.n195 source.n194 9.3005
R257 source.n168 source.n167 9.3005
R258 source.n189 source.n188 9.3005
R259 source.n187 source.n186 9.3005
R260 source.n172 source.n171 9.3005
R261 source.n181 source.n180 9.3005
R262 source.n179 source.n178 9.3005
R263 source.n161 source.n160 9.3005
R264 source.n134 source.n133 9.3005
R265 source.n155 source.n154 9.3005
R266 source.n153 source.n152 9.3005
R267 source.n138 source.n137 9.3005
R268 source.n147 source.n146 9.3005
R269 source.n145 source.n144 9.3005
R270 source.n29 source.n28 9.3005
R271 source.n2 source.n1 9.3005
R272 source.n23 source.n22 9.3005
R273 source.n21 source.n20 9.3005
R274 source.n6 source.n5 9.3005
R275 source.n15 source.n14 9.3005
R276 source.n13 source.n12 9.3005
R277 source.n63 source.n62 9.3005
R278 source.n36 source.n35 9.3005
R279 source.n57 source.n56 9.3005
R280 source.n55 source.n54 9.3005
R281 source.n40 source.n39 9.3005
R282 source.n49 source.n48 9.3005
R283 source.n47 source.n46 9.3005
R284 source.n95 source.n94 9.3005
R285 source.n68 source.n67 9.3005
R286 source.n89 source.n88 9.3005
R287 source.n87 source.n86 9.3005
R288 source.n72 source.n71 9.3005
R289 source.n81 source.n80 9.3005
R290 source.n79 source.n78 9.3005
R291 source.n129 source.n128 9.3005
R292 source.n102 source.n101 9.3005
R293 source.n123 source.n122 9.3005
R294 source.n121 source.n120 9.3005
R295 source.n106 source.n105 9.3005
R296 source.n115 source.n114 9.3005
R297 source.n113 source.n112 9.3005
R298 source.n259 source.n234 8.92171
R299 source.n225 source.n200 8.92171
R300 source.n193 source.n168 8.92171
R301 source.n159 source.n134 8.92171
R302 source.n27 source.n2 8.92171
R303 source.n61 source.n36 8.92171
R304 source.n93 source.n68 8.92171
R305 source.n127 source.n102 8.92171
R306 source.n260 source.n232 8.14595
R307 source.n226 source.n198 8.14595
R308 source.n194 source.n166 8.14595
R309 source.n160 source.n132 8.14595
R310 source.n28 source.n0 8.14595
R311 source.n62 source.n34 8.14595
R312 source.n94 source.n66 8.14595
R313 source.n128 source.n100 8.14595
R314 source.n262 source.n232 5.81868
R315 source.n228 source.n198 5.81868
R316 source.n196 source.n166 5.81868
R317 source.n162 source.n132 5.81868
R318 source.n30 source.n0 5.81868
R319 source.n64 source.n34 5.81868
R320 source.n96 source.n66 5.81868
R321 source.n130 source.n100 5.81868
R322 source.n264 source.n263 5.7505
R323 source.n260 source.n259 5.04292
R324 source.n226 source.n225 5.04292
R325 source.n194 source.n193 5.04292
R326 source.n160 source.n159 5.04292
R327 source.n28 source.n27 5.04292
R328 source.n62 source.n61 5.04292
R329 source.n94 source.n93 5.04292
R330 source.n128 source.n127 5.04292
R331 source.n245 source.n241 4.38594
R332 source.n211 source.n207 4.38594
R333 source.n179 source.n175 4.38594
R334 source.n145 source.n141 4.38594
R335 source.n13 source.n9 4.38594
R336 source.n47 source.n43 4.38594
R337 source.n79 source.n75 4.38594
R338 source.n113 source.n109 4.38594
R339 source.n256 source.n234 4.26717
R340 source.n222 source.n200 4.26717
R341 source.n190 source.n168 4.26717
R342 source.n156 source.n134 4.26717
R343 source.n24 source.n2 4.26717
R344 source.n58 source.n36 4.26717
R345 source.n90 source.n68 4.26717
R346 source.n124 source.n102 4.26717
R347 source.n255 source.n236 3.49141
R348 source.n221 source.n202 3.49141
R349 source.n189 source.n170 3.49141
R350 source.n155 source.n136 3.49141
R351 source.n23 source.n4 3.49141
R352 source.n57 source.n38 3.49141
R353 source.n89 source.n70 3.49141
R354 source.n123 source.n104 3.49141
R355 source.n230 source.t7 3.3005
R356 source.n230 source.t5 3.3005
R357 source.n164 source.t14 3.3005
R358 source.n164 source.t15 3.3005
R359 source.n32 source.t10 3.3005
R360 source.n32 source.t11 3.3005
R361 source.n98 source.t0 3.3005
R362 source.n98 source.t4 3.3005
R363 source.n252 source.n251 2.71565
R364 source.n218 source.n217 2.71565
R365 source.n186 source.n185 2.71565
R366 source.n152 source.n151 2.71565
R367 source.n20 source.n19 2.71565
R368 source.n54 source.n53 2.71565
R369 source.n86 source.n85 2.71565
R370 source.n120 source.n119 2.71565
R371 source.n248 source.n238 1.93989
R372 source.n214 source.n204 1.93989
R373 source.n182 source.n172 1.93989
R374 source.n148 source.n138 1.93989
R375 source.n16 source.n6 1.93989
R376 source.n50 source.n40 1.93989
R377 source.n82 source.n72 1.93989
R378 source.n116 source.n106 1.93989
R379 source.n247 source.n240 1.16414
R380 source.n213 source.n206 1.16414
R381 source.n181 source.n174 1.16414
R382 source.n147 source.n140 1.16414
R383 source.n15 source.n8 1.16414
R384 source.n49 source.n42 1.16414
R385 source.n81 source.n74 1.16414
R386 source.n115 source.n108 1.16414
R387 source.n131 source.n99 0.974638
R388 source.n99 source.n97 0.974638
R389 source.n65 source.n33 0.974638
R390 source.n33 source.n31 0.974638
R391 source.n165 source.n163 0.974638
R392 source.n197 source.n165 0.974638
R393 source.n231 source.n229 0.974638
R394 source.n263 source.n231 0.974638
R395 source.n97 source.n65 0.470328
R396 source.n229 source.n197 0.470328
R397 source.n244 source.n243 0.388379
R398 source.n210 source.n209 0.388379
R399 source.n178 source.n177 0.388379
R400 source.n144 source.n143 0.388379
R401 source.n12 source.n11 0.388379
R402 source.n46 source.n45 0.388379
R403 source.n78 source.n77 0.388379
R404 source.n112 source.n111 0.388379
R405 source source.n264 0.188
R406 source.n246 source.n245 0.155672
R407 source.n246 source.n237 0.155672
R408 source.n253 source.n237 0.155672
R409 source.n254 source.n253 0.155672
R410 source.n254 source.n233 0.155672
R411 source.n261 source.n233 0.155672
R412 source.n212 source.n211 0.155672
R413 source.n212 source.n203 0.155672
R414 source.n219 source.n203 0.155672
R415 source.n220 source.n219 0.155672
R416 source.n220 source.n199 0.155672
R417 source.n227 source.n199 0.155672
R418 source.n180 source.n179 0.155672
R419 source.n180 source.n171 0.155672
R420 source.n187 source.n171 0.155672
R421 source.n188 source.n187 0.155672
R422 source.n188 source.n167 0.155672
R423 source.n195 source.n167 0.155672
R424 source.n146 source.n145 0.155672
R425 source.n146 source.n137 0.155672
R426 source.n153 source.n137 0.155672
R427 source.n154 source.n153 0.155672
R428 source.n154 source.n133 0.155672
R429 source.n161 source.n133 0.155672
R430 source.n29 source.n1 0.155672
R431 source.n22 source.n1 0.155672
R432 source.n22 source.n21 0.155672
R433 source.n21 source.n5 0.155672
R434 source.n14 source.n5 0.155672
R435 source.n14 source.n13 0.155672
R436 source.n63 source.n35 0.155672
R437 source.n56 source.n35 0.155672
R438 source.n56 source.n55 0.155672
R439 source.n55 source.n39 0.155672
R440 source.n48 source.n39 0.155672
R441 source.n48 source.n47 0.155672
R442 source.n95 source.n67 0.155672
R443 source.n88 source.n67 0.155672
R444 source.n88 source.n87 0.155672
R445 source.n87 source.n71 0.155672
R446 source.n80 source.n71 0.155672
R447 source.n80 source.n79 0.155672
R448 source.n129 source.n101 0.155672
R449 source.n122 source.n101 0.155672
R450 source.n122 source.n121 0.155672
R451 source.n121 source.n105 0.155672
R452 source.n114 source.n105 0.155672
R453 source.n114 source.n113 0.155672
R454 minus.n2 minus.t5 250.457
R455 minus.n10 minus.t4 250.457
R456 minus.n1 minus.t3 229.855
R457 minus.n4 minus.t2 229.855
R458 minus.n6 minus.t6 229.855
R459 minus.n9 minus.t0 229.855
R460 minus.n12 minus.t1 229.855
R461 minus.n14 minus.t7 229.855
R462 minus.n7 minus.n6 161.3
R463 minus.n5 minus.n0 161.3
R464 minus.n15 minus.n14 161.3
R465 minus.n13 minus.n8 161.3
R466 minus.n4 minus.n3 80.6037
R467 minus.n12 minus.n11 80.6037
R468 minus.n4 minus.n1 48.2005
R469 minus.n12 minus.n9 48.2005
R470 minus.n5 minus.n4 41.6278
R471 minus.n13 minus.n12 41.6278
R472 minus.n16 minus.n7 31.7202
R473 minus.n3 minus.n2 31.6158
R474 minus.n11 minus.n10 31.6158
R475 minus.n2 minus.n1 17.6494
R476 minus.n10 minus.n9 17.6494
R477 minus.n16 minus.n15 6.65202
R478 minus.n6 minus.n5 6.57323
R479 minus.n14 minus.n13 6.57323
R480 minus.n3 minus.n0 0.285035
R481 minus.n11 minus.n8 0.285035
R482 minus.n7 minus.n0 0.189894
R483 minus.n15 minus.n8 0.189894
R484 minus minus.n16 0.188
R485 drain_right.n5 drain_right.n3 68.1648
R486 drain_right.n2 drain_right.n1 67.6224
R487 drain_right.n2 drain_right.n0 67.6224
R488 drain_right.n5 drain_right.n4 67.1908
R489 drain_right drain_right.n2 25.6779
R490 drain_right drain_right.n5 6.62735
R491 drain_right.n1 drain_right.t6 3.3005
R492 drain_right.n1 drain_right.t0 3.3005
R493 drain_right.n0 drain_right.t3 3.3005
R494 drain_right.n0 drain_right.t7 3.3005
R495 drain_right.n3 drain_right.t4 3.3005
R496 drain_right.n3 drain_right.t2 3.3005
R497 drain_right.n4 drain_right.t1 3.3005
R498 drain_right.n4 drain_right.t5 3.3005
C0 drain_left source 6.43793f
C1 drain_right drain_left 0.873724f
C2 drain_left minus 0.17159f
C3 drain_right source 6.44032f
C4 drain_left plus 3.32869f
C5 minus source 3.249f
C6 drain_right minus 3.14944f
C7 source plus 3.26302f
C8 drain_right plus 0.333957f
C9 minus plus 4.33214f
C10 drain_right a_n1846_n2088# 4.5566f
C11 drain_left a_n1846_n2088# 4.83325f
C12 source a_n1846_n2088# 5.481861f
C13 minus a_n1846_n2088# 6.667921f
C14 plus a_n1846_n2088# 8.00836f
C15 drain_right.t3 a_n1846_n2088# 0.12249f
C16 drain_right.t7 a_n1846_n2088# 0.12249f
C17 drain_right.n0 a_n1846_n2088# 1.02373f
C18 drain_right.t6 a_n1846_n2088# 0.12249f
C19 drain_right.t0 a_n1846_n2088# 0.12249f
C20 drain_right.n1 a_n1846_n2088# 1.02373f
C21 drain_right.n2 a_n1846_n2088# 1.57853f
C22 drain_right.t4 a_n1846_n2088# 0.12249f
C23 drain_right.t2 a_n1846_n2088# 0.12249f
C24 drain_right.n3 a_n1846_n2088# 1.02703f
C25 drain_right.t1 a_n1846_n2088# 0.12249f
C26 drain_right.t5 a_n1846_n2088# 0.12249f
C27 drain_right.n4 a_n1846_n2088# 1.02157f
C28 drain_right.n5 a_n1846_n2088# 0.980317f
C29 minus.n0 a_n1846_n2088# 0.056715f
C30 minus.t3 a_n1846_n2088# 0.591761f
C31 minus.n1 a_n1846_n2088# 0.282125f
C32 minus.t2 a_n1846_n2088# 0.591761f
C33 minus.t5 a_n1846_n2088# 0.614253f
C34 minus.n2 a_n1846_n2088# 0.254485f
C35 minus.n3 a_n1846_n2088# 0.243262f
C36 minus.n4 a_n1846_n2088# 0.281433f
C37 minus.n5 a_n1846_n2088# 0.009645f
C38 minus.t6 a_n1846_n2088# 0.591761f
C39 minus.n6 a_n1846_n2088# 0.265499f
C40 minus.n7 a_n1846_n2088# 1.22022f
C41 minus.n8 a_n1846_n2088# 0.056715f
C42 minus.t0 a_n1846_n2088# 0.591761f
C43 minus.n9 a_n1846_n2088# 0.282125f
C44 minus.t4 a_n1846_n2088# 0.614253f
C45 minus.n10 a_n1846_n2088# 0.254485f
C46 minus.n11 a_n1846_n2088# 0.243262f
C47 minus.t1 a_n1846_n2088# 0.591761f
C48 minus.n12 a_n1846_n2088# 0.281433f
C49 minus.n13 a_n1846_n2088# 0.009645f
C50 minus.t7 a_n1846_n2088# 0.591761f
C51 minus.n14 a_n1846_n2088# 0.265499f
C52 minus.n15 a_n1846_n2088# 0.292991f
C53 minus.n16 a_n1846_n2088# 1.49348f
C54 source.n0 a_n1846_n2088# 0.03017f
C55 source.n1 a_n1846_n2088# 0.021464f
C56 source.n2 a_n1846_n2088# 0.011534f
C57 source.n3 a_n1846_n2088# 0.027262f
C58 source.n4 a_n1846_n2088# 0.012212f
C59 source.n5 a_n1846_n2088# 0.021464f
C60 source.n6 a_n1846_n2088# 0.011534f
C61 source.n7 a_n1846_n2088# 0.027262f
C62 source.n8 a_n1846_n2088# 0.012212f
C63 source.n9 a_n1846_n2088# 0.091851f
C64 source.t12 a_n1846_n2088# 0.044433f
C65 source.n10 a_n1846_n2088# 0.020446f
C66 source.n11 a_n1846_n2088# 0.016103f
C67 source.n12 a_n1846_n2088# 0.011534f
C68 source.n13 a_n1846_n2088# 0.510716f
C69 source.n14 a_n1846_n2088# 0.021464f
C70 source.n15 a_n1846_n2088# 0.011534f
C71 source.n16 a_n1846_n2088# 0.012212f
C72 source.n17 a_n1846_n2088# 0.027262f
C73 source.n18 a_n1846_n2088# 0.027262f
C74 source.n19 a_n1846_n2088# 0.012212f
C75 source.n20 a_n1846_n2088# 0.011534f
C76 source.n21 a_n1846_n2088# 0.021464f
C77 source.n22 a_n1846_n2088# 0.021464f
C78 source.n23 a_n1846_n2088# 0.011534f
C79 source.n24 a_n1846_n2088# 0.012212f
C80 source.n25 a_n1846_n2088# 0.027262f
C81 source.n26 a_n1846_n2088# 0.059017f
C82 source.n27 a_n1846_n2088# 0.012212f
C83 source.n28 a_n1846_n2088# 0.011534f
C84 source.n29 a_n1846_n2088# 0.049613f
C85 source.n30 a_n1846_n2088# 0.033023f
C86 source.n31 a_n1846_n2088# 0.570899f
C87 source.t10 a_n1846_n2088# 0.101769f
C88 source.t11 a_n1846_n2088# 0.101769f
C89 source.n32 a_n1846_n2088# 0.792587f
C90 source.n33 a_n1846_n2088# 0.335951f
C91 source.n34 a_n1846_n2088# 0.03017f
C92 source.n35 a_n1846_n2088# 0.021464f
C93 source.n36 a_n1846_n2088# 0.011534f
C94 source.n37 a_n1846_n2088# 0.027262f
C95 source.n38 a_n1846_n2088# 0.012212f
C96 source.n39 a_n1846_n2088# 0.021464f
C97 source.n40 a_n1846_n2088# 0.011534f
C98 source.n41 a_n1846_n2088# 0.027262f
C99 source.n42 a_n1846_n2088# 0.012212f
C100 source.n43 a_n1846_n2088# 0.091851f
C101 source.t9 a_n1846_n2088# 0.044433f
C102 source.n44 a_n1846_n2088# 0.020446f
C103 source.n45 a_n1846_n2088# 0.016103f
C104 source.n46 a_n1846_n2088# 0.011534f
C105 source.n47 a_n1846_n2088# 0.510716f
C106 source.n48 a_n1846_n2088# 0.021464f
C107 source.n49 a_n1846_n2088# 0.011534f
C108 source.n50 a_n1846_n2088# 0.012212f
C109 source.n51 a_n1846_n2088# 0.027262f
C110 source.n52 a_n1846_n2088# 0.027262f
C111 source.n53 a_n1846_n2088# 0.012212f
C112 source.n54 a_n1846_n2088# 0.011534f
C113 source.n55 a_n1846_n2088# 0.021464f
C114 source.n56 a_n1846_n2088# 0.021464f
C115 source.n57 a_n1846_n2088# 0.011534f
C116 source.n58 a_n1846_n2088# 0.012212f
C117 source.n59 a_n1846_n2088# 0.027262f
C118 source.n60 a_n1846_n2088# 0.059017f
C119 source.n61 a_n1846_n2088# 0.012212f
C120 source.n62 a_n1846_n2088# 0.011534f
C121 source.n63 a_n1846_n2088# 0.049613f
C122 source.n64 a_n1846_n2088# 0.033023f
C123 source.n65 a_n1846_n2088# 0.118199f
C124 source.n66 a_n1846_n2088# 0.03017f
C125 source.n67 a_n1846_n2088# 0.021464f
C126 source.n68 a_n1846_n2088# 0.011534f
C127 source.n69 a_n1846_n2088# 0.027262f
C128 source.n70 a_n1846_n2088# 0.012212f
C129 source.n71 a_n1846_n2088# 0.021464f
C130 source.n72 a_n1846_n2088# 0.011534f
C131 source.n73 a_n1846_n2088# 0.027262f
C132 source.n74 a_n1846_n2088# 0.012212f
C133 source.n75 a_n1846_n2088# 0.091851f
C134 source.t1 a_n1846_n2088# 0.044433f
C135 source.n76 a_n1846_n2088# 0.020446f
C136 source.n77 a_n1846_n2088# 0.016103f
C137 source.n78 a_n1846_n2088# 0.011534f
C138 source.n79 a_n1846_n2088# 0.510716f
C139 source.n80 a_n1846_n2088# 0.021464f
C140 source.n81 a_n1846_n2088# 0.011534f
C141 source.n82 a_n1846_n2088# 0.012212f
C142 source.n83 a_n1846_n2088# 0.027262f
C143 source.n84 a_n1846_n2088# 0.027262f
C144 source.n85 a_n1846_n2088# 0.012212f
C145 source.n86 a_n1846_n2088# 0.011534f
C146 source.n87 a_n1846_n2088# 0.021464f
C147 source.n88 a_n1846_n2088# 0.021464f
C148 source.n89 a_n1846_n2088# 0.011534f
C149 source.n90 a_n1846_n2088# 0.012212f
C150 source.n91 a_n1846_n2088# 0.027262f
C151 source.n92 a_n1846_n2088# 0.059017f
C152 source.n93 a_n1846_n2088# 0.012212f
C153 source.n94 a_n1846_n2088# 0.011534f
C154 source.n95 a_n1846_n2088# 0.049613f
C155 source.n96 a_n1846_n2088# 0.033023f
C156 source.n97 a_n1846_n2088# 0.118199f
C157 source.t0 a_n1846_n2088# 0.101769f
C158 source.t4 a_n1846_n2088# 0.101769f
C159 source.n98 a_n1846_n2088# 0.792587f
C160 source.n99 a_n1846_n2088# 0.335951f
C161 source.n100 a_n1846_n2088# 0.03017f
C162 source.n101 a_n1846_n2088# 0.021464f
C163 source.n102 a_n1846_n2088# 0.011534f
C164 source.n103 a_n1846_n2088# 0.027262f
C165 source.n104 a_n1846_n2088# 0.012212f
C166 source.n105 a_n1846_n2088# 0.021464f
C167 source.n106 a_n1846_n2088# 0.011534f
C168 source.n107 a_n1846_n2088# 0.027262f
C169 source.n108 a_n1846_n2088# 0.012212f
C170 source.n109 a_n1846_n2088# 0.091851f
C171 source.t3 a_n1846_n2088# 0.044433f
C172 source.n110 a_n1846_n2088# 0.020446f
C173 source.n111 a_n1846_n2088# 0.016103f
C174 source.n112 a_n1846_n2088# 0.011534f
C175 source.n113 a_n1846_n2088# 0.510716f
C176 source.n114 a_n1846_n2088# 0.021464f
C177 source.n115 a_n1846_n2088# 0.011534f
C178 source.n116 a_n1846_n2088# 0.012212f
C179 source.n117 a_n1846_n2088# 0.027262f
C180 source.n118 a_n1846_n2088# 0.027262f
C181 source.n119 a_n1846_n2088# 0.012212f
C182 source.n120 a_n1846_n2088# 0.011534f
C183 source.n121 a_n1846_n2088# 0.021464f
C184 source.n122 a_n1846_n2088# 0.021464f
C185 source.n123 a_n1846_n2088# 0.011534f
C186 source.n124 a_n1846_n2088# 0.012212f
C187 source.n125 a_n1846_n2088# 0.027262f
C188 source.n126 a_n1846_n2088# 0.059017f
C189 source.n127 a_n1846_n2088# 0.012212f
C190 source.n128 a_n1846_n2088# 0.011534f
C191 source.n129 a_n1846_n2088# 0.049613f
C192 source.n130 a_n1846_n2088# 0.033023f
C193 source.n131 a_n1846_n2088# 0.855851f
C194 source.n132 a_n1846_n2088# 0.03017f
C195 source.n133 a_n1846_n2088# 0.021464f
C196 source.n134 a_n1846_n2088# 0.011534f
C197 source.n135 a_n1846_n2088# 0.027262f
C198 source.n136 a_n1846_n2088# 0.012212f
C199 source.n137 a_n1846_n2088# 0.021464f
C200 source.n138 a_n1846_n2088# 0.011534f
C201 source.n139 a_n1846_n2088# 0.027262f
C202 source.n140 a_n1846_n2088# 0.012212f
C203 source.n141 a_n1846_n2088# 0.091851f
C204 source.t8 a_n1846_n2088# 0.044433f
C205 source.n142 a_n1846_n2088# 0.020446f
C206 source.n143 a_n1846_n2088# 0.016103f
C207 source.n144 a_n1846_n2088# 0.011534f
C208 source.n145 a_n1846_n2088# 0.510716f
C209 source.n146 a_n1846_n2088# 0.021464f
C210 source.n147 a_n1846_n2088# 0.011534f
C211 source.n148 a_n1846_n2088# 0.012212f
C212 source.n149 a_n1846_n2088# 0.027262f
C213 source.n150 a_n1846_n2088# 0.027262f
C214 source.n151 a_n1846_n2088# 0.012212f
C215 source.n152 a_n1846_n2088# 0.011534f
C216 source.n153 a_n1846_n2088# 0.021464f
C217 source.n154 a_n1846_n2088# 0.021464f
C218 source.n155 a_n1846_n2088# 0.011534f
C219 source.n156 a_n1846_n2088# 0.012212f
C220 source.n157 a_n1846_n2088# 0.027262f
C221 source.n158 a_n1846_n2088# 0.059017f
C222 source.n159 a_n1846_n2088# 0.012212f
C223 source.n160 a_n1846_n2088# 0.011534f
C224 source.n161 a_n1846_n2088# 0.049613f
C225 source.n162 a_n1846_n2088# 0.033023f
C226 source.n163 a_n1846_n2088# 0.855851f
C227 source.t14 a_n1846_n2088# 0.101769f
C228 source.t15 a_n1846_n2088# 0.101769f
C229 source.n164 a_n1846_n2088# 0.792581f
C230 source.n165 a_n1846_n2088# 0.335957f
C231 source.n166 a_n1846_n2088# 0.03017f
C232 source.n167 a_n1846_n2088# 0.021464f
C233 source.n168 a_n1846_n2088# 0.011534f
C234 source.n169 a_n1846_n2088# 0.027262f
C235 source.n170 a_n1846_n2088# 0.012212f
C236 source.n171 a_n1846_n2088# 0.021464f
C237 source.n172 a_n1846_n2088# 0.011534f
C238 source.n173 a_n1846_n2088# 0.027262f
C239 source.n174 a_n1846_n2088# 0.012212f
C240 source.n175 a_n1846_n2088# 0.091851f
C241 source.t13 a_n1846_n2088# 0.044433f
C242 source.n176 a_n1846_n2088# 0.020446f
C243 source.n177 a_n1846_n2088# 0.016103f
C244 source.n178 a_n1846_n2088# 0.011534f
C245 source.n179 a_n1846_n2088# 0.510716f
C246 source.n180 a_n1846_n2088# 0.021464f
C247 source.n181 a_n1846_n2088# 0.011534f
C248 source.n182 a_n1846_n2088# 0.012212f
C249 source.n183 a_n1846_n2088# 0.027262f
C250 source.n184 a_n1846_n2088# 0.027262f
C251 source.n185 a_n1846_n2088# 0.012212f
C252 source.n186 a_n1846_n2088# 0.011534f
C253 source.n187 a_n1846_n2088# 0.021464f
C254 source.n188 a_n1846_n2088# 0.021464f
C255 source.n189 a_n1846_n2088# 0.011534f
C256 source.n190 a_n1846_n2088# 0.012212f
C257 source.n191 a_n1846_n2088# 0.027262f
C258 source.n192 a_n1846_n2088# 0.059017f
C259 source.n193 a_n1846_n2088# 0.012212f
C260 source.n194 a_n1846_n2088# 0.011534f
C261 source.n195 a_n1846_n2088# 0.049613f
C262 source.n196 a_n1846_n2088# 0.033023f
C263 source.n197 a_n1846_n2088# 0.118199f
C264 source.n198 a_n1846_n2088# 0.03017f
C265 source.n199 a_n1846_n2088# 0.021464f
C266 source.n200 a_n1846_n2088# 0.011534f
C267 source.n201 a_n1846_n2088# 0.027262f
C268 source.n202 a_n1846_n2088# 0.012212f
C269 source.n203 a_n1846_n2088# 0.021464f
C270 source.n204 a_n1846_n2088# 0.011534f
C271 source.n205 a_n1846_n2088# 0.027262f
C272 source.n206 a_n1846_n2088# 0.012212f
C273 source.n207 a_n1846_n2088# 0.091851f
C274 source.t2 a_n1846_n2088# 0.044433f
C275 source.n208 a_n1846_n2088# 0.020446f
C276 source.n209 a_n1846_n2088# 0.016103f
C277 source.n210 a_n1846_n2088# 0.011534f
C278 source.n211 a_n1846_n2088# 0.510716f
C279 source.n212 a_n1846_n2088# 0.021464f
C280 source.n213 a_n1846_n2088# 0.011534f
C281 source.n214 a_n1846_n2088# 0.012212f
C282 source.n215 a_n1846_n2088# 0.027262f
C283 source.n216 a_n1846_n2088# 0.027262f
C284 source.n217 a_n1846_n2088# 0.012212f
C285 source.n218 a_n1846_n2088# 0.011534f
C286 source.n219 a_n1846_n2088# 0.021464f
C287 source.n220 a_n1846_n2088# 0.021464f
C288 source.n221 a_n1846_n2088# 0.011534f
C289 source.n222 a_n1846_n2088# 0.012212f
C290 source.n223 a_n1846_n2088# 0.027262f
C291 source.n224 a_n1846_n2088# 0.059017f
C292 source.n225 a_n1846_n2088# 0.012212f
C293 source.n226 a_n1846_n2088# 0.011534f
C294 source.n227 a_n1846_n2088# 0.049613f
C295 source.n228 a_n1846_n2088# 0.033023f
C296 source.n229 a_n1846_n2088# 0.118199f
C297 source.t7 a_n1846_n2088# 0.101769f
C298 source.t5 a_n1846_n2088# 0.101769f
C299 source.n230 a_n1846_n2088# 0.792581f
C300 source.n231 a_n1846_n2088# 0.335957f
C301 source.n232 a_n1846_n2088# 0.03017f
C302 source.n233 a_n1846_n2088# 0.021464f
C303 source.n234 a_n1846_n2088# 0.011534f
C304 source.n235 a_n1846_n2088# 0.027262f
C305 source.n236 a_n1846_n2088# 0.012212f
C306 source.n237 a_n1846_n2088# 0.021464f
C307 source.n238 a_n1846_n2088# 0.011534f
C308 source.n239 a_n1846_n2088# 0.027262f
C309 source.n240 a_n1846_n2088# 0.012212f
C310 source.n241 a_n1846_n2088# 0.091851f
C311 source.t6 a_n1846_n2088# 0.044433f
C312 source.n242 a_n1846_n2088# 0.020446f
C313 source.n243 a_n1846_n2088# 0.016103f
C314 source.n244 a_n1846_n2088# 0.011534f
C315 source.n245 a_n1846_n2088# 0.510716f
C316 source.n246 a_n1846_n2088# 0.021464f
C317 source.n247 a_n1846_n2088# 0.011534f
C318 source.n248 a_n1846_n2088# 0.012212f
C319 source.n249 a_n1846_n2088# 0.027262f
C320 source.n250 a_n1846_n2088# 0.027262f
C321 source.n251 a_n1846_n2088# 0.012212f
C322 source.n252 a_n1846_n2088# 0.011534f
C323 source.n253 a_n1846_n2088# 0.021464f
C324 source.n254 a_n1846_n2088# 0.021464f
C325 source.n255 a_n1846_n2088# 0.011534f
C326 source.n256 a_n1846_n2088# 0.012212f
C327 source.n257 a_n1846_n2088# 0.027262f
C328 source.n258 a_n1846_n2088# 0.059017f
C329 source.n259 a_n1846_n2088# 0.012212f
C330 source.n260 a_n1846_n2088# 0.011534f
C331 source.n261 a_n1846_n2088# 0.049613f
C332 source.n262 a_n1846_n2088# 0.033023f
C333 source.n263 a_n1846_n2088# 0.262857f
C334 source.n264 a_n1846_n2088# 0.893214f
C335 drain_left.t6 a_n1846_n2088# 0.123753f
C336 drain_left.t1 a_n1846_n2088# 0.123753f
C337 drain_left.n0 a_n1846_n2088# 1.03428f
C338 drain_left.t7 a_n1846_n2088# 0.123753f
C339 drain_left.t4 a_n1846_n2088# 0.123753f
C340 drain_left.n1 a_n1846_n2088# 1.03428f
C341 drain_left.n2 a_n1846_n2088# 1.64779f
C342 drain_left.t2 a_n1846_n2088# 0.123753f
C343 drain_left.t0 a_n1846_n2088# 0.123753f
C344 drain_left.n3 a_n1846_n2088# 1.03762f
C345 drain_left.t3 a_n1846_n2088# 0.123753f
C346 drain_left.t5 a_n1846_n2088# 0.123753f
C347 drain_left.n4 a_n1846_n2088# 1.0321f
C348 drain_left.n5 a_n1846_n2088# 0.990419f
C349 plus.n0 a_n1846_n2088# 0.058797f
C350 plus.t3 a_n1846_n2088# 0.613483f
C351 plus.t4 a_n1846_n2088# 0.613483f
C352 plus.n1 a_n1846_n2088# 0.252192f
C353 plus.t5 a_n1846_n2088# 0.613483f
C354 plus.t6 a_n1846_n2088# 0.636801f
C355 plus.n2 a_n1846_n2088# 0.263827f
C356 plus.n3 a_n1846_n2088# 0.292482f
C357 plus.n4 a_n1846_n2088# 0.291764f
C358 plus.n5 a_n1846_n2088# 0.009999f
C359 plus.n6 a_n1846_n2088# 0.275245f
C360 plus.n7 a_n1846_n2088# 0.393955f
C361 plus.n8 a_n1846_n2088# 0.058797f
C362 plus.t7 a_n1846_n2088# 0.613483f
C363 plus.n9 a_n1846_n2088# 0.252192f
C364 plus.t1 a_n1846_n2088# 0.613483f
C365 plus.t2 a_n1846_n2088# 0.636801f
C366 plus.n10 a_n1846_n2088# 0.263827f
C367 plus.t0 a_n1846_n2088# 0.613483f
C368 plus.n11 a_n1846_n2088# 0.292482f
C369 plus.n12 a_n1846_n2088# 0.291764f
C370 plus.n13 a_n1846_n2088# 0.009999f
C371 plus.n14 a_n1846_n2088# 0.275245f
C372 plus.n15 a_n1846_n2088# 1.14412f
.ends

