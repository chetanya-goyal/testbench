* NGSPICE file created from diffpair521.ext - technology: sky130A

.subckt diffpair521 minus drain_right drain_left source plus
X0 source.t7 plus.t0 drain_left.t3 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X1 drain_left.t2 plus.t1 source.t6 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X2 source.t0 minus.t0 drain_right.t3 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X3 source.t5 plus.t2 drain_left.t1 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X4 drain_right.t2 minus.t1 source.t1 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X5 source.t2 minus.t2 drain_right.t1 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X6 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X7 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X8 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X9 drain_right.t0 minus.t3 source.t3 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X10 drain_left.t0 plus.t3 source.t4 a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X11 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
R0 plus.n0 plus.t2 822.548
R1 plus.n1 plus.t1 822.548
R2 plus.n0 plus.t3 822.524
R3 plus.n1 plus.t0 822.524
R4 plus plus.n1 99.0155
R5 plus plus.n0 83.5586
R6 drain_left drain_left.n0 91.9499
R7 drain_left drain_left.n1 67.2479
R8 drain_left.n0 drain_left.t3 1.3205
R9 drain_left.n0 drain_left.t2 1.3205
R10 drain_left.n1 drain_left.t1 1.3205
R11 drain_left.n1 drain_left.t0 1.3205
R12 source.n1 source.t5 45.521
R13 source.n2 source.t3 45.521
R14 source.n3 source.t0 45.521
R15 source.n7 source.t1 45.5208
R16 source.n6 source.t2 45.5208
R17 source.n5 source.t6 45.5208
R18 source.n4 source.t7 45.5208
R19 source.n0 source.t4 45.5208
R20 source.n4 source.n3 24.276
R21 source.n8 source.n0 18.6553
R22 source.n8 source.n7 5.62119
R23 source.n3 source.n2 0.716017
R24 source.n1 source.n0 0.716017
R25 source.n5 source.n4 0.716017
R26 source.n7 source.n6 0.716017
R27 source.n2 source.n1 0.470328
R28 source.n6 source.n5 0.470328
R29 source source.n8 0.188
R30 minus.n0 minus.t3 822.548
R31 minus.n1 minus.t2 822.548
R32 minus.n0 minus.t0 822.524
R33 minus.n1 minus.t1 822.524
R34 minus.n2 minus.n0 106.27
R35 minus.n2 minus.n1 76.7783
R36 minus minus.n2 0.188
R37 drain_right drain_right.n0 91.3967
R38 drain_right drain_right.n1 67.2479
R39 drain_right.n0 drain_right.t1 1.3205
R40 drain_right.n0 drain_right.t2 1.3205
R41 drain_right.n1 drain_right.t3 1.3205
R42 drain_right.n1 drain_right.t0 1.3205
C0 drain_left source 9.46804f
C1 drain_left minus 0.170454f
C2 source drain_right 9.467791f
C3 minus drain_right 3.31192f
C4 source minus 2.72935f
C5 plus drain_left 3.42537f
C6 plus drain_right 0.266739f
C7 plus source 2.74339f
C8 plus minus 5.21392f
C9 drain_left drain_right 0.522435f
C10 drain_right a_n1214_n3888# 7.33525f
C11 drain_left a_n1214_n3888# 7.53766f
C12 source a_n1214_n3888# 10.384101f
C13 minus a_n1214_n3888# 4.785806f
C14 plus a_n1214_n3888# 8.753481f
C15 drain_right.t1 a_n1214_n3888# 0.347818f
C16 drain_right.t2 a_n1214_n3888# 0.347818f
C17 drain_right.n0 a_n1214_n3888# 3.63914f
C18 drain_right.t3 a_n1214_n3888# 0.347818f
C19 drain_right.t0 a_n1214_n3888# 0.347818f
C20 drain_right.n1 a_n1214_n3888# 3.20443f
C21 minus.t3 a_n1214_n3888# 1.1697f
C22 minus.t0 a_n1214_n3888# 1.16968f
C23 minus.n0 a_n1214_n3888# 1.55032f
C24 minus.t2 a_n1214_n3888# 1.1697f
C25 minus.t1 a_n1214_n3888# 1.16968f
C26 minus.n1 a_n1214_n3888# 0.916116f
C27 minus.n2 a_n1214_n3888# 4.01912f
C28 source.t4 a_n1214_n3888# 2.23335f
C29 source.n0 a_n1214_n3888# 1.04951f
C30 source.t5 a_n1214_n3888# 2.23336f
C31 source.n1 a_n1214_n3888# 0.290568f
C32 source.t3 a_n1214_n3888# 2.23336f
C33 source.n2 a_n1214_n3888# 0.290568f
C34 source.t0 a_n1214_n3888# 2.23336f
C35 source.n3 a_n1214_n3888# 1.33265f
C36 source.t7 a_n1214_n3888# 2.23335f
C37 source.n4 a_n1214_n3888# 1.33266f
C38 source.t6 a_n1214_n3888# 2.23335f
C39 source.n5 a_n1214_n3888# 0.290571f
C40 source.t2 a_n1214_n3888# 2.23335f
C41 source.n6 a_n1214_n3888# 0.290571f
C42 source.t1 a_n1214_n3888# 2.23335f
C43 source.n7 a_n1214_n3888# 0.392901f
C44 source.n8 a_n1214_n3888# 1.23486f
C45 drain_left.t3 a_n1214_n3888# 0.34742f
C46 drain_left.t2 a_n1214_n3888# 0.34742f
C47 drain_left.n0 a_n1214_n3888# 3.66176f
C48 drain_left.t1 a_n1214_n3888# 0.34742f
C49 drain_left.t0 a_n1214_n3888# 0.34742f
C50 drain_left.n1 a_n1214_n3888# 3.20076f
C51 plus.t3 a_n1214_n3888# 1.19182f
C52 plus.t2 a_n1214_n3888# 1.19184f
C53 plus.n0 a_n1214_n3888# 1.01982f
C54 plus.t0 a_n1214_n3888# 1.19182f
C55 plus.t1 a_n1214_n3888# 1.19184f
C56 plus.n1 a_n1214_n3888# 1.37918f
.ends

