* NGSPICE file created from diffpair248.ext - technology: sky130A

.subckt diffpair248 minus drain_right drain_left source plus
X0 source.t37 plus.t0 drain_left.t9 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X1 drain_left.t2 plus.t1 source.t36 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X2 source.t8 minus.t0 drain_right.t19 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X3 source.t1 minus.t1 drain_right.t18 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X4 drain_left.t1 plus.t2 source.t35 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X5 drain_left.t0 plus.t3 source.t34 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 drain_right.t17 minus.t2 source.t4 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 drain_right.t16 minus.t3 source.t11 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X9 drain_right.t15 minus.t4 source.t13 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X10 source.t33 plus.t4 drain_left.t12 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X11 source.t14 minus.t5 drain_right.t14 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X12 source.t9 minus.t6 drain_right.t13 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X13 source.t38 minus.t7 drain_right.t12 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X14 a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X15 drain_right.t11 minus.t8 source.t39 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X16 drain_right.t10 minus.t9 source.t3 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X17 drain_right.t9 minus.t10 source.t0 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 source.t32 plus.t5 drain_left.t14 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X19 source.t2 minus.t11 drain_right.t8 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X20 drain_right.t7 minus.t12 source.t16 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X21 drain_right.t6 minus.t13 source.t10 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 drain_left.t7 plus.t6 source.t31 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X23 source.t30 plus.t7 drain_left.t6 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X24 drain_right.t5 minus.t14 source.t6 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X25 drain_right.t4 minus.t15 source.t12 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X26 source.t15 minus.t16 drain_right.t3 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X27 a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X28 source.t5 minus.t17 drain_right.t2 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X29 source.t29 plus.t8 drain_left.t18 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X30 drain_left.t17 plus.t9 source.t28 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X31 source.t7 minus.t18 drain_right.t1 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X32 a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X33 drain_left.t16 plus.t10 source.t27 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X34 source.t26 plus.t11 drain_left.t8 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X35 source.t25 plus.t12 drain_left.t19 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X36 source.t17 minus.t19 drain_right.t0 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X37 drain_left.t10 plus.t13 source.t24 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X38 source.t23 plus.t14 drain_left.t11 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X39 drain_left.t4 plus.t15 source.t22 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X40 drain_left.t5 plus.t16 source.t21 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X41 source.t20 plus.t17 drain_left.t3 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X42 drain_left.t13 plus.t18 source.t19 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X43 source.t18 plus.t19 drain_left.t15 a_n2146_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
R0 plus.n6 plus.t7 1234.94
R1 plus.n27 plus.t10 1234.94
R2 plus.n36 plus.t2 1234.94
R3 plus.n56 plus.t5 1234.94
R4 plus.n5 plus.t16 1172.87
R5 plus.n9 plus.t12 1172.87
R6 plus.n3 plus.t9 1172.87
R7 plus.n15 plus.t19 1172.87
R8 plus.n17 plus.t15 1172.87
R9 plus.n18 plus.t11 1172.87
R10 plus.n24 plus.t6 1172.87
R11 plus.n26 plus.t14 1172.87
R12 plus.n35 plus.t4 1172.87
R13 plus.n39 plus.t13 1172.87
R14 plus.n33 plus.t0 1172.87
R15 plus.n45 plus.t3 1172.87
R16 plus.n47 plus.t8 1172.87
R17 plus.n32 plus.t18 1172.87
R18 plus.n53 plus.t17 1172.87
R19 plus.n55 plus.t1 1172.87
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 69.3793
R47 plus.n19 plus.n18 69.3793
R48 plus.n48 plus.n32 69.3793
R49 plus.n44 plus.n33 69.3793
R50 plus.n9 plus.n8 54.7732
R51 plus.n25 plus.n24 54.7732
R52 plus.n54 plus.n53 54.7732
R53 plus.n39 plus.n38 54.7732
R54 plus.n16 plus.n15 47.4702
R55 plus.n17 plus.n16 47.4702
R56 plus.n47 plus.n46 47.4702
R57 plus.n46 plus.n45 47.4702
R58 plus.n8 plus.n5 40.1672
R59 plus.n26 plus.n25 40.1672
R60 plus.n55 plus.n54 40.1672
R61 plus.n38 plus.n35 40.1672
R62 plus.n6 plus.n5 32.8641
R63 plus.n27 plus.n26 32.8641
R64 plus.n56 plus.n55 32.8641
R65 plus.n36 plus.n35 32.8641
R66 plus plus.n57 28.9195
R67 plus.n15 plus.n14 25.5611
R68 plus.n19 plus.n17 25.5611
R69 plus.n48 plus.n47 25.5611
R70 plus.n45 plus.n44 25.5611
R71 plus.n10 plus.n9 18.2581
R72 plus.n24 plus.n23 18.2581
R73 plus.n53 plus.n52 18.2581
R74 plus.n40 plus.n39 18.2581
R75 plus plus.n28 9.93232
R76 plus.n11 plus.n3 3.65202
R77 plus.n18 plus.n1 3.65202
R78 plus.n32 plus.n30 3.65202
R79 plus.n41 plus.n33 3.65202
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 drain_left.n10 drain_left.n8 67.7512
R99 drain_left.n6 drain_left.n4 67.751
R100 drain_left.n2 drain_left.n0 67.751
R101 drain_left.n14 drain_left.n13 67.1908
R102 drain_left.n12 drain_left.n11 67.1908
R103 drain_left.n10 drain_left.n9 67.1908
R104 drain_left.n16 drain_left.n15 67.1907
R105 drain_left.n7 drain_left.n3 67.1907
R106 drain_left.n6 drain_left.n5 67.1907
R107 drain_left.n2 drain_left.n1 67.1907
R108 drain_left drain_left.n7 27.3044
R109 drain_left drain_left.n16 6.21356
R110 drain_left.n3 drain_left.t18 5.0005
R111 drain_left.n3 drain_left.t0 5.0005
R112 drain_left.n4 drain_left.t12 5.0005
R113 drain_left.n4 drain_left.t1 5.0005
R114 drain_left.n5 drain_left.t9 5.0005
R115 drain_left.n5 drain_left.t10 5.0005
R116 drain_left.n1 drain_left.t3 5.0005
R117 drain_left.n1 drain_left.t13 5.0005
R118 drain_left.n0 drain_left.t14 5.0005
R119 drain_left.n0 drain_left.t2 5.0005
R120 drain_left.n15 drain_left.t11 5.0005
R121 drain_left.n15 drain_left.t16 5.0005
R122 drain_left.n13 drain_left.t8 5.0005
R123 drain_left.n13 drain_left.t7 5.0005
R124 drain_left.n11 drain_left.t15 5.0005
R125 drain_left.n11 drain_left.t4 5.0005
R126 drain_left.n9 drain_left.t19 5.0005
R127 drain_left.n9 drain_left.t17 5.0005
R128 drain_left.n8 drain_left.t6 5.0005
R129 drain_left.n8 drain_left.t5 5.0005
R130 drain_left.n12 drain_left.n10 0.560845
R131 drain_left.n14 drain_left.n12 0.560845
R132 drain_left.n16 drain_left.n14 0.560845
R133 drain_left.n7 drain_left.n6 0.505499
R134 drain_left.n7 drain_left.n2 0.505499
R135 source.n9 source.t30 55.512
R136 source.n10 source.t39 55.512
R137 source.n19 source.t17 55.512
R138 source.n0 source.t27 55.5119
R139 source.n39 source.t13 55.5119
R140 source.n30 source.t15 55.5119
R141 source.n29 source.t35 55.5119
R142 source.n20 source.t32 55.5119
R143 source.n2 source.n1 50.512
R144 source.n4 source.n3 50.512
R145 source.n6 source.n5 50.512
R146 source.n8 source.n7 50.512
R147 source.n12 source.n11 50.512
R148 source.n14 source.n13 50.512
R149 source.n16 source.n15 50.512
R150 source.n18 source.n17 50.512
R151 source.n38 source.n37 50.5119
R152 source.n36 source.n35 50.5119
R153 source.n34 source.n33 50.5119
R154 source.n32 source.n31 50.5119
R155 source.n28 source.n27 50.5119
R156 source.n26 source.n25 50.5119
R157 source.n24 source.n23 50.5119
R158 source.n22 source.n21 50.5119
R159 source.n20 source.n19 17.3026
R160 source.n40 source.n0 11.7595
R161 source.n40 source.n39 5.5436
R162 source.n37 source.t16 5.0005
R163 source.n37 source.t1 5.0005
R164 source.n35 source.t11 5.0005
R165 source.n35 source.t9 5.0005
R166 source.n33 source.t0 5.0005
R167 source.n33 source.t8 5.0005
R168 source.n31 source.t4 5.0005
R169 source.n31 source.t14 5.0005
R170 source.n27 source.t24 5.0005
R171 source.n27 source.t33 5.0005
R172 source.n25 source.t34 5.0005
R173 source.n25 source.t37 5.0005
R174 source.n23 source.t19 5.0005
R175 source.n23 source.t29 5.0005
R176 source.n21 source.t36 5.0005
R177 source.n21 source.t20 5.0005
R178 source.n1 source.t31 5.0005
R179 source.n1 source.t23 5.0005
R180 source.n3 source.t22 5.0005
R181 source.n3 source.t26 5.0005
R182 source.n5 source.t28 5.0005
R183 source.n5 source.t18 5.0005
R184 source.n7 source.t21 5.0005
R185 source.n7 source.t25 5.0005
R186 source.n11 source.t6 5.0005
R187 source.n11 source.t38 5.0005
R188 source.n13 source.t3 5.0005
R189 source.n13 source.t2 5.0005
R190 source.n15 source.t12 5.0005
R191 source.n15 source.t7 5.0005
R192 source.n17 source.t10 5.0005
R193 source.n17 source.t5 5.0005
R194 source.n19 source.n18 0.560845
R195 source.n18 source.n16 0.560845
R196 source.n16 source.n14 0.560845
R197 source.n14 source.n12 0.560845
R198 source.n12 source.n10 0.560845
R199 source.n9 source.n8 0.560845
R200 source.n8 source.n6 0.560845
R201 source.n6 source.n4 0.560845
R202 source.n4 source.n2 0.560845
R203 source.n2 source.n0 0.560845
R204 source.n22 source.n20 0.560845
R205 source.n24 source.n22 0.560845
R206 source.n26 source.n24 0.560845
R207 source.n28 source.n26 0.560845
R208 source.n29 source.n28 0.560845
R209 source.n32 source.n30 0.560845
R210 source.n34 source.n32 0.560845
R211 source.n36 source.n34 0.560845
R212 source.n38 source.n36 0.560845
R213 source.n39 source.n38 0.560845
R214 source.n10 source.n9 0.470328
R215 source.n30 source.n29 0.470328
R216 source source.n40 0.188
R217 minus.n27 minus.t19 1234.94
R218 minus.n7 minus.t8 1234.94
R219 minus.n56 minus.t4 1234.94
R220 minus.n35 minus.t16 1234.94
R221 minus.n26 minus.t13 1172.87
R222 minus.n24 minus.t17 1172.87
R223 minus.n3 minus.t15 1172.87
R224 minus.n18 minus.t18 1172.87
R225 minus.n16 minus.t9 1172.87
R226 minus.n4 minus.t11 1172.87
R227 minus.n10 minus.t14 1172.87
R228 minus.n6 minus.t7 1172.87
R229 minus.n55 minus.t1 1172.87
R230 minus.n53 minus.t12 1172.87
R231 minus.n47 minus.t6 1172.87
R232 minus.n46 minus.t3 1172.87
R233 minus.n44 minus.t0 1172.87
R234 minus.n32 minus.t10 1172.87
R235 minus.n38 minus.t5 1172.87
R236 minus.n34 minus.t2 1172.87
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 69.3793
R264 minus.n15 minus.n4 69.3793
R265 minus.n43 minus.n32 69.3793
R266 minus.n48 minus.n47 69.3793
R267 minus.n25 minus.n24 54.7732
R268 minus.n10 minus.n9 54.7732
R269 minus.n38 minus.n37 54.7732
R270 minus.n54 minus.n53 54.7732
R271 minus.n18 minus.n17 47.4702
R272 minus.n17 minus.n16 47.4702
R273 minus.n45 minus.n44 47.4702
R274 minus.n46 minus.n45 47.4702
R275 minus.n26 minus.n25 40.1672
R276 minus.n9 minus.n6 40.1672
R277 minus.n37 minus.n34 40.1672
R278 minus.n55 minus.n54 40.1672
R279 minus.n27 minus.n26 32.8641
R280 minus.n7 minus.n6 32.8641
R281 minus.n35 minus.n34 32.8641
R282 minus.n56 minus.n55 32.8641
R283 minus.n58 minus.n28 32.7657
R284 minus.n19 minus.n18 25.5611
R285 minus.n16 minus.n15 25.5611
R286 minus.n44 minus.n43 25.5611
R287 minus.n48 minus.n46 25.5611
R288 minus.n24 minus.n23 18.2581
R289 minus.n11 minus.n10 18.2581
R290 minus.n39 minus.n38 18.2581
R291 minus.n53 minus.n52 18.2581
R292 minus.n58 minus.n57 6.56111
R293 minus.n3 minus.n1 3.65202
R294 minus.n12 minus.n4 3.65202
R295 minus.n40 minus.n32 3.65202
R296 minus.n47 minus.n30 3.65202
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 67.751
R317 drain_right.n6 drain_right.n4 67.751
R318 drain_right.n2 drain_right.n0 67.751
R319 drain_right.n10 drain_right.n9 67.1908
R320 drain_right.n12 drain_right.n11 67.1908
R321 drain_right.n14 drain_right.n13 67.1908
R322 drain_right.n16 drain_right.n15 67.1908
R323 drain_right.n7 drain_right.n3 67.1907
R324 drain_right.n6 drain_right.n5 67.1907
R325 drain_right.n2 drain_right.n1 67.1907
R326 drain_right drain_right.n7 26.7511
R327 drain_right drain_right.n16 6.21356
R328 drain_right.n3 drain_right.t19 5.0005
R329 drain_right.n3 drain_right.t16 5.0005
R330 drain_right.n4 drain_right.t18 5.0005
R331 drain_right.n4 drain_right.t15 5.0005
R332 drain_right.n5 drain_right.t13 5.0005
R333 drain_right.n5 drain_right.t7 5.0005
R334 drain_right.n1 drain_right.t14 5.0005
R335 drain_right.n1 drain_right.t9 5.0005
R336 drain_right.n0 drain_right.t3 5.0005
R337 drain_right.n0 drain_right.t17 5.0005
R338 drain_right.n8 drain_right.t12 5.0005
R339 drain_right.n8 drain_right.t11 5.0005
R340 drain_right.n9 drain_right.t8 5.0005
R341 drain_right.n9 drain_right.t5 5.0005
R342 drain_right.n11 drain_right.t1 5.0005
R343 drain_right.n11 drain_right.t10 5.0005
R344 drain_right.n13 drain_right.t2 5.0005
R345 drain_right.n13 drain_right.t4 5.0005
R346 drain_right.n15 drain_right.t0 5.0005
R347 drain_right.n15 drain_right.t6 5.0005
R348 drain_right.n16 drain_right.n14 0.560845
R349 drain_right.n14 drain_right.n12 0.560845
R350 drain_right.n12 drain_right.n10 0.560845
R351 drain_right.n7 drain_right.n6 0.505499
R352 drain_right.n7 drain_right.n2 0.505499
C0 drain_left plus 2.6279f
C1 drain_left minus 0.171338f
C2 plus minus 4.70176f
C3 drain_left source 20.8286f
C4 plus source 2.32014f
C5 minus source 2.30612f
C6 drain_left drain_right 1.13563f
C7 drain_right plus 0.364841f
C8 drain_right minus 2.41721f
C9 drain_right source 20.8291f
C10 drain_right a_n2146_n2088# 5.28349f
C11 drain_left a_n2146_n2088# 5.60129f
C12 source a_n2146_n2088# 5.540656f
C13 minus a_n2146_n2088# 7.442463f
C14 plus a_n2146_n2088# 9.19155f
C15 drain_right.t3 a_n2146_n2088# 0.202053f
C16 drain_right.t17 a_n2146_n2088# 0.202053f
C17 drain_right.n0 a_n2146_n2088# 1.2524f
C18 drain_right.t14 a_n2146_n2088# 0.202053f
C19 drain_right.t9 a_n2146_n2088# 0.202053f
C20 drain_right.n1 a_n2146_n2088# 1.24958f
C21 drain_right.n2 a_n2146_n2088# 0.66447f
C22 drain_right.t19 a_n2146_n2088# 0.202053f
C23 drain_right.t16 a_n2146_n2088# 0.202053f
C24 drain_right.n3 a_n2146_n2088# 1.24958f
C25 drain_right.t18 a_n2146_n2088# 0.202053f
C26 drain_right.t15 a_n2146_n2088# 0.202053f
C27 drain_right.n4 a_n2146_n2088# 1.2524f
C28 drain_right.t13 a_n2146_n2088# 0.202053f
C29 drain_right.t7 a_n2146_n2088# 0.202053f
C30 drain_right.n5 a_n2146_n2088# 1.24958f
C31 drain_right.n6 a_n2146_n2088# 0.66447f
C32 drain_right.n7 a_n2146_n2088# 1.32369f
C33 drain_right.t12 a_n2146_n2088# 0.202053f
C34 drain_right.t11 a_n2146_n2088# 0.202053f
C35 drain_right.n8 a_n2146_n2088# 1.2524f
C36 drain_right.t8 a_n2146_n2088# 0.202053f
C37 drain_right.t5 a_n2146_n2088# 0.202053f
C38 drain_right.n9 a_n2146_n2088# 1.24958f
C39 drain_right.n10 a_n2146_n2088# 0.668189f
C40 drain_right.t1 a_n2146_n2088# 0.202053f
C41 drain_right.t10 a_n2146_n2088# 0.202053f
C42 drain_right.n11 a_n2146_n2088# 1.24958f
C43 drain_right.n12 a_n2146_n2088# 0.329839f
C44 drain_right.t2 a_n2146_n2088# 0.202053f
C45 drain_right.t4 a_n2146_n2088# 0.202053f
C46 drain_right.n13 a_n2146_n2088# 1.24958f
C47 drain_right.n14 a_n2146_n2088# 0.329839f
C48 drain_right.t0 a_n2146_n2088# 0.202053f
C49 drain_right.t6 a_n2146_n2088# 0.202053f
C50 drain_right.n15 a_n2146_n2088# 1.24958f
C51 drain_right.n16 a_n2146_n2088# 0.564719f
C52 minus.n0 a_n2146_n2088# 0.051598f
C53 minus.t19 a_n2146_n2088# 0.135884f
C54 minus.t13 a_n2146_n2088# 0.132311f
C55 minus.t17 a_n2146_n2088# 0.132311f
C56 minus.n1 a_n2146_n2088# 0.017912f
C57 minus.n2 a_n2146_n2088# 0.051598f
C58 minus.t15 a_n2146_n2088# 0.132311f
C59 minus.n3 a_n2146_n2088# 0.068686f
C60 minus.t18 a_n2146_n2088# 0.132311f
C61 minus.t9 a_n2146_n2088# 0.132311f
C62 minus.t11 a_n2146_n2088# 0.132311f
C63 minus.n4 a_n2146_n2088# 0.068686f
C64 minus.n5 a_n2146_n2088# 0.051598f
C65 minus.t14 a_n2146_n2088# 0.132311f
C66 minus.t7 a_n2146_n2088# 0.132311f
C67 minus.n6 a_n2146_n2088# 0.068686f
C68 minus.t8 a_n2146_n2088# 0.135884f
C69 minus.n7 a_n2146_n2088# 0.089467f
C70 minus.n8 a_n2146_n2088# 0.119023f
C71 minus.n9 a_n2146_n2088# 0.021889f
C72 minus.n10 a_n2146_n2088# 0.068686f
C73 minus.n11 a_n2146_n2088# 0.021093f
C74 minus.n12 a_n2146_n2088# 0.017912f
C75 minus.n13 a_n2146_n2088# 0.051598f
C76 minus.n14 a_n2146_n2088# 0.051598f
C77 minus.n15 a_n2146_n2088# 0.021889f
C78 minus.n16 a_n2146_n2088# 0.068686f
C79 minus.n17 a_n2146_n2088# 0.021889f
C80 minus.n18 a_n2146_n2088# 0.068686f
C81 minus.n19 a_n2146_n2088# 0.021889f
C82 minus.n20 a_n2146_n2088# 0.051598f
C83 minus.n21 a_n2146_n2088# 0.051598f
C84 minus.n22 a_n2146_n2088# 0.051598f
C85 minus.n23 a_n2146_n2088# 0.021093f
C86 minus.n24 a_n2146_n2088# 0.068686f
C87 minus.n25 a_n2146_n2088# 0.021889f
C88 minus.n26 a_n2146_n2088# 0.068686f
C89 minus.n27 a_n2146_n2088# 0.089388f
C90 minus.n28 a_n2146_n2088# 1.55804f
C91 minus.n29 a_n2146_n2088# 0.051598f
C92 minus.t1 a_n2146_n2088# 0.132311f
C93 minus.t12 a_n2146_n2088# 0.132311f
C94 minus.n30 a_n2146_n2088# 0.017912f
C95 minus.n31 a_n2146_n2088# 0.051598f
C96 minus.t3 a_n2146_n2088# 0.132311f
C97 minus.t0 a_n2146_n2088# 0.132311f
C98 minus.t10 a_n2146_n2088# 0.132311f
C99 minus.n32 a_n2146_n2088# 0.068686f
C100 minus.n33 a_n2146_n2088# 0.051598f
C101 minus.t5 a_n2146_n2088# 0.132311f
C102 minus.t2 a_n2146_n2088# 0.132311f
C103 minus.n34 a_n2146_n2088# 0.068686f
C104 minus.t16 a_n2146_n2088# 0.135884f
C105 minus.n35 a_n2146_n2088# 0.089467f
C106 minus.n36 a_n2146_n2088# 0.119023f
C107 minus.n37 a_n2146_n2088# 0.021889f
C108 minus.n38 a_n2146_n2088# 0.068686f
C109 minus.n39 a_n2146_n2088# 0.021093f
C110 minus.n40 a_n2146_n2088# 0.017912f
C111 minus.n41 a_n2146_n2088# 0.051598f
C112 minus.n42 a_n2146_n2088# 0.051598f
C113 minus.n43 a_n2146_n2088# 0.021889f
C114 minus.n44 a_n2146_n2088# 0.068686f
C115 minus.n45 a_n2146_n2088# 0.021889f
C116 minus.n46 a_n2146_n2088# 0.068686f
C117 minus.t6 a_n2146_n2088# 0.132311f
C118 minus.n47 a_n2146_n2088# 0.068686f
C119 minus.n48 a_n2146_n2088# 0.021889f
C120 minus.n49 a_n2146_n2088# 0.051598f
C121 minus.n50 a_n2146_n2088# 0.051598f
C122 minus.n51 a_n2146_n2088# 0.051598f
C123 minus.n52 a_n2146_n2088# 0.021093f
C124 minus.n53 a_n2146_n2088# 0.068686f
C125 minus.n54 a_n2146_n2088# 0.021889f
C126 minus.n55 a_n2146_n2088# 0.068686f
C127 minus.t4 a_n2146_n2088# 0.135884f
C128 minus.n56 a_n2146_n2088# 0.089388f
C129 minus.n57 a_n2146_n2088# 0.344742f
C130 minus.n58 a_n2146_n2088# 1.9076f
C131 source.t27 a_n2146_n2088# 1.30918f
C132 source.n0 a_n2146_n2088# 0.963131f
C133 source.t31 a_n2146_n2088# 0.186391f
C134 source.t23 a_n2146_n2088# 0.186391f
C135 source.n1 a_n2146_n2088# 1.08482f
C136 source.n2 a_n2146_n2088# 0.336908f
C137 source.t22 a_n2146_n2088# 0.186391f
C138 source.t26 a_n2146_n2088# 0.186391f
C139 source.n3 a_n2146_n2088# 1.08482f
C140 source.n4 a_n2146_n2088# 0.336908f
C141 source.t28 a_n2146_n2088# 0.186391f
C142 source.t18 a_n2146_n2088# 0.186391f
C143 source.n5 a_n2146_n2088# 1.08482f
C144 source.n6 a_n2146_n2088# 0.336908f
C145 source.t21 a_n2146_n2088# 0.186391f
C146 source.t25 a_n2146_n2088# 0.186391f
C147 source.n7 a_n2146_n2088# 1.08482f
C148 source.n8 a_n2146_n2088# 0.336908f
C149 source.t30 a_n2146_n2088# 1.30918f
C150 source.n9 a_n2146_n2088# 0.440483f
C151 source.t39 a_n2146_n2088# 1.30918f
C152 source.n10 a_n2146_n2088# 0.440483f
C153 source.t6 a_n2146_n2088# 0.186391f
C154 source.t38 a_n2146_n2088# 0.186391f
C155 source.n11 a_n2146_n2088# 1.08482f
C156 source.n12 a_n2146_n2088# 0.336908f
C157 source.t3 a_n2146_n2088# 0.186391f
C158 source.t2 a_n2146_n2088# 0.186391f
C159 source.n13 a_n2146_n2088# 1.08482f
C160 source.n14 a_n2146_n2088# 0.336908f
C161 source.t12 a_n2146_n2088# 0.186391f
C162 source.t7 a_n2146_n2088# 0.186391f
C163 source.n15 a_n2146_n2088# 1.08482f
C164 source.n16 a_n2146_n2088# 0.336908f
C165 source.t10 a_n2146_n2088# 0.186391f
C166 source.t5 a_n2146_n2088# 0.186391f
C167 source.n17 a_n2146_n2088# 1.08482f
C168 source.n18 a_n2146_n2088# 0.336908f
C169 source.t17 a_n2146_n2088# 1.30918f
C170 source.n19 a_n2146_n2088# 1.29756f
C171 source.t32 a_n2146_n2088# 1.30918f
C172 source.n20 a_n2146_n2088# 1.29757f
C173 source.t36 a_n2146_n2088# 0.186391f
C174 source.t20 a_n2146_n2088# 0.186391f
C175 source.n21 a_n2146_n2088# 1.08482f
C176 source.n22 a_n2146_n2088# 0.336915f
C177 source.t19 a_n2146_n2088# 0.186391f
C178 source.t29 a_n2146_n2088# 0.186391f
C179 source.n23 a_n2146_n2088# 1.08482f
C180 source.n24 a_n2146_n2088# 0.336915f
C181 source.t34 a_n2146_n2088# 0.186391f
C182 source.t37 a_n2146_n2088# 0.186391f
C183 source.n25 a_n2146_n2088# 1.08482f
C184 source.n26 a_n2146_n2088# 0.336915f
C185 source.t24 a_n2146_n2088# 0.186391f
C186 source.t33 a_n2146_n2088# 0.186391f
C187 source.n27 a_n2146_n2088# 1.08482f
C188 source.n28 a_n2146_n2088# 0.336915f
C189 source.t35 a_n2146_n2088# 1.30918f
C190 source.n29 a_n2146_n2088# 0.440489f
C191 source.t15 a_n2146_n2088# 1.30918f
C192 source.n30 a_n2146_n2088# 0.440489f
C193 source.t4 a_n2146_n2088# 0.186391f
C194 source.t14 a_n2146_n2088# 0.186391f
C195 source.n31 a_n2146_n2088# 1.08482f
C196 source.n32 a_n2146_n2088# 0.336915f
C197 source.t0 a_n2146_n2088# 0.186391f
C198 source.t8 a_n2146_n2088# 0.186391f
C199 source.n33 a_n2146_n2088# 1.08482f
C200 source.n34 a_n2146_n2088# 0.336915f
C201 source.t11 a_n2146_n2088# 0.186391f
C202 source.t9 a_n2146_n2088# 0.186391f
C203 source.n35 a_n2146_n2088# 1.08482f
C204 source.n36 a_n2146_n2088# 0.336915f
C205 source.t16 a_n2146_n2088# 0.186391f
C206 source.t1 a_n2146_n2088# 0.186391f
C207 source.n37 a_n2146_n2088# 1.08482f
C208 source.n38 a_n2146_n2088# 0.336915f
C209 source.t13 a_n2146_n2088# 1.30918f
C210 source.n39 a_n2146_n2088# 0.588104f
C211 source.n40 a_n2146_n2088# 1.06235f
C212 drain_left.t14 a_n2146_n2088# 0.202833f
C213 drain_left.t2 a_n2146_n2088# 0.202833f
C214 drain_left.n0 a_n2146_n2088# 1.25723f
C215 drain_left.t3 a_n2146_n2088# 0.202833f
C216 drain_left.t13 a_n2146_n2088# 0.202833f
C217 drain_left.n1 a_n2146_n2088# 1.2544f
C218 drain_left.n2 a_n2146_n2088# 0.667035f
C219 drain_left.t18 a_n2146_n2088# 0.202833f
C220 drain_left.t0 a_n2146_n2088# 0.202833f
C221 drain_left.n3 a_n2146_n2088# 1.2544f
C222 drain_left.t12 a_n2146_n2088# 0.202833f
C223 drain_left.t1 a_n2146_n2088# 0.202833f
C224 drain_left.n4 a_n2146_n2088# 1.25723f
C225 drain_left.t9 a_n2146_n2088# 0.202833f
C226 drain_left.t10 a_n2146_n2088# 0.202833f
C227 drain_left.n5 a_n2146_n2088# 1.2544f
C228 drain_left.n6 a_n2146_n2088# 0.667035f
C229 drain_left.n7 a_n2146_n2088# 1.38582f
C230 drain_left.t6 a_n2146_n2088# 0.202833f
C231 drain_left.t5 a_n2146_n2088# 0.202833f
C232 drain_left.n8 a_n2146_n2088# 1.25724f
C233 drain_left.t19 a_n2146_n2088# 0.202833f
C234 drain_left.t17 a_n2146_n2088# 0.202833f
C235 drain_left.n9 a_n2146_n2088# 1.25441f
C236 drain_left.n10 a_n2146_n2088# 0.670763f
C237 drain_left.t15 a_n2146_n2088# 0.202833f
C238 drain_left.t4 a_n2146_n2088# 0.202833f
C239 drain_left.n11 a_n2146_n2088# 1.25441f
C240 drain_left.n12 a_n2146_n2088# 0.331112f
C241 drain_left.t8 a_n2146_n2088# 0.202833f
C242 drain_left.t7 a_n2146_n2088# 0.202833f
C243 drain_left.n13 a_n2146_n2088# 1.25441f
C244 drain_left.n14 a_n2146_n2088# 0.331112f
C245 drain_left.t11 a_n2146_n2088# 0.202833f
C246 drain_left.t16 a_n2146_n2088# 0.202833f
C247 drain_left.n15 a_n2146_n2088# 1.2544f
C248 drain_left.n16 a_n2146_n2088# 0.566904f
C249 plus.n0 a_n2146_n2088# 0.053288f
C250 plus.t14 a_n2146_n2088# 0.136643f
C251 plus.t6 a_n2146_n2088# 0.136643f
C252 plus.n1 a_n2146_n2088# 0.018499f
C253 plus.n2 a_n2146_n2088# 0.053288f
C254 plus.t15 a_n2146_n2088# 0.136643f
C255 plus.t19 a_n2146_n2088# 0.136643f
C256 plus.t9 a_n2146_n2088# 0.136643f
C257 plus.n3 a_n2146_n2088# 0.070935f
C258 plus.n4 a_n2146_n2088# 0.053288f
C259 plus.t12 a_n2146_n2088# 0.136643f
C260 plus.t16 a_n2146_n2088# 0.136643f
C261 plus.n5 a_n2146_n2088# 0.070935f
C262 plus.t7 a_n2146_n2088# 0.140333f
C263 plus.n6 a_n2146_n2088# 0.092397f
C264 plus.n7 a_n2146_n2088# 0.12292f
C265 plus.n8 a_n2146_n2088# 0.022605f
C266 plus.n9 a_n2146_n2088# 0.070935f
C267 plus.n10 a_n2146_n2088# 0.021784f
C268 plus.n11 a_n2146_n2088# 0.018499f
C269 plus.n12 a_n2146_n2088# 0.053288f
C270 plus.n13 a_n2146_n2088# 0.053288f
C271 plus.n14 a_n2146_n2088# 0.022605f
C272 plus.n15 a_n2146_n2088# 0.070935f
C273 plus.n16 a_n2146_n2088# 0.022605f
C274 plus.n17 a_n2146_n2088# 0.070935f
C275 plus.t11 a_n2146_n2088# 0.136643f
C276 plus.n18 a_n2146_n2088# 0.070935f
C277 plus.n19 a_n2146_n2088# 0.022605f
C278 plus.n20 a_n2146_n2088# 0.053288f
C279 plus.n21 a_n2146_n2088# 0.053288f
C280 plus.n22 a_n2146_n2088# 0.053288f
C281 plus.n23 a_n2146_n2088# 0.021784f
C282 plus.n24 a_n2146_n2088# 0.070935f
C283 plus.n25 a_n2146_n2088# 0.022605f
C284 plus.n26 a_n2146_n2088# 0.070935f
C285 plus.t10 a_n2146_n2088# 0.140333f
C286 plus.n27 a_n2146_n2088# 0.092315f
C287 plus.n28 a_n2146_n2088# 0.464603f
C288 plus.n29 a_n2146_n2088# 0.053288f
C289 plus.t5 a_n2146_n2088# 0.140333f
C290 plus.t1 a_n2146_n2088# 0.136643f
C291 plus.t17 a_n2146_n2088# 0.136643f
C292 plus.n30 a_n2146_n2088# 0.018499f
C293 plus.n31 a_n2146_n2088# 0.053288f
C294 plus.t18 a_n2146_n2088# 0.136643f
C295 plus.n32 a_n2146_n2088# 0.070935f
C296 plus.t8 a_n2146_n2088# 0.136643f
C297 plus.t3 a_n2146_n2088# 0.136643f
C298 plus.t0 a_n2146_n2088# 0.136643f
C299 plus.n33 a_n2146_n2088# 0.070935f
C300 plus.n34 a_n2146_n2088# 0.053288f
C301 plus.t13 a_n2146_n2088# 0.136643f
C302 plus.t4 a_n2146_n2088# 0.136643f
C303 plus.n35 a_n2146_n2088# 0.070935f
C304 plus.t2 a_n2146_n2088# 0.140333f
C305 plus.n36 a_n2146_n2088# 0.092397f
C306 plus.n37 a_n2146_n2088# 0.12292f
C307 plus.n38 a_n2146_n2088# 0.022605f
C308 plus.n39 a_n2146_n2088# 0.070935f
C309 plus.n40 a_n2146_n2088# 0.021784f
C310 plus.n41 a_n2146_n2088# 0.018499f
C311 plus.n42 a_n2146_n2088# 0.053288f
C312 plus.n43 a_n2146_n2088# 0.053288f
C313 plus.n44 a_n2146_n2088# 0.022605f
C314 plus.n45 a_n2146_n2088# 0.070935f
C315 plus.n46 a_n2146_n2088# 0.022605f
C316 plus.n47 a_n2146_n2088# 0.070935f
C317 plus.n48 a_n2146_n2088# 0.022605f
C318 plus.n49 a_n2146_n2088# 0.053288f
C319 plus.n50 a_n2146_n2088# 0.053288f
C320 plus.n51 a_n2146_n2088# 0.053288f
C321 plus.n52 a_n2146_n2088# 0.021784f
C322 plus.n53 a_n2146_n2088# 0.070935f
C323 plus.n54 a_n2146_n2088# 0.022605f
C324 plus.n55 a_n2146_n2088# 0.070935f
C325 plus.n56 a_n2146_n2088# 0.092315f
C326 plus.n57 a_n2146_n2088# 1.45455f
.ends

