* NGSPICE file created from diffpair487.ext - technology: sky130A

.subckt diffpair487 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t5 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X1 drain_right.t15 minus.t1 source.t30 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X2 drain_right.t7 minus.t2 source.t29 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X3 source.t28 minus.t3 drain_right.t10 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X4 source.t7 plus.t0 drain_left.t15 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X5 drain_left.t14 plus.t1 source.t9 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X6 a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X7 a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X8 drain_left.t13 plus.t2 source.t11 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X9 source.t6 plus.t3 drain_left.t12 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X10 source.t27 minus.t4 drain_right.t13 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X11 drain_right.t4 minus.t5 source.t26 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X12 drain_right.t1 minus.t6 source.t25 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X13 source.t8 plus.t4 drain_left.t11 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X14 a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X15 source.t24 minus.t7 drain_right.t3 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X16 source.t23 minus.t8 drain_right.t6 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X17 drain_left.t10 plus.t5 source.t2 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X18 source.t1 plus.t6 drain_left.t9 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X19 drain_right.t9 minus.t9 source.t22 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X20 drain_right.t12 minus.t10 source.t21 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X21 drain_left.t8 plus.t7 source.t3 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X22 source.t20 minus.t11 drain_right.t0 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X23 drain_left.t7 plus.t8 source.t5 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X24 source.t19 minus.t12 drain_right.t14 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X25 drain_right.t2 minus.t13 source.t18 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X26 drain_left.t6 plus.t9 source.t10 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X27 source.t12 plus.t10 drain_left.t5 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X28 source.t0 plus.t11 drain_left.t4 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X29 drain_right.t8 minus.t14 source.t17 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X30 drain_left.t3 plus.t12 source.t14 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X31 drain_left.t2 plus.t13 source.t4 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X32 source.t13 plus.t14 drain_left.t1 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X33 a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X34 source.t15 plus.t15 drain_left.t0 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X35 source.t16 minus.t15 drain_right.t11 a_n1886_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
R0 minus.n21 minus.t11 2659.03
R1 minus.n5 minus.t5 2659.03
R2 minus.n44 minus.t2 2659.03
R3 minus.n28 minus.t3 2659.03
R4 minus.n20 minus.t10 2618.87
R5 minus.n1 minus.t12 2618.87
R6 minus.n14 minus.t6 2618.87
R7 minus.n12 minus.t7 2618.87
R8 minus.n3 minus.t9 2618.87
R9 minus.n6 minus.t4 2618.87
R10 minus.n43 minus.t0 2618.87
R11 minus.n24 minus.t14 2618.87
R12 minus.n37 minus.t8 2618.87
R13 minus.n35 minus.t1 2618.87
R14 minus.n26 minus.t15 2618.87
R15 minus.n29 minus.t13 2618.87
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 69.3793
R39 minus.n11 minus.n3 69.3793
R40 minus.n34 minus.n26 69.3793
R41 minus.n38 minus.n24 69.3793
R42 minus.n21 minus.n20 54.7732
R43 minus.n6 minus.n5 54.7732
R44 minus.n29 minus.n28 54.7732
R45 minus.n44 minus.n43 54.7732
R46 minus.n14 minus.n13 47.4702
R47 minus.n13 minus.n12 47.4702
R48 minus.n36 minus.n35 47.4702
R49 minus.n37 minus.n36 47.4702
R50 minus.n46 minus.n22 38.5422
R51 minus.n15 minus.n14 25.5611
R52 minus.n12 minus.n11 25.5611
R53 minus.n35 minus.n34 25.5611
R54 minus.n38 minus.n37 25.5611
R55 minus.n20 minus.n19 18.2581
R56 minus.n7 minus.n6 18.2581
R57 minus.n30 minus.n29 18.2581
R58 minus.n43 minus.n42 18.2581
R59 minus.n46 minus.n45 6.50429
R60 minus.n18 minus.n1 3.65202
R61 minus.n8 minus.n3 3.65202
R62 minus.n31 minus.n26 3.65202
R63 minus.n41 minus.n24 3.65202
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 drain_right.n9 drain_right.n7 61.44
R80 drain_right.n5 drain_right.n3 61.4399
R81 drain_right.n2 drain_right.n0 61.4399
R82 drain_right.n9 drain_right.n8 60.8798
R83 drain_right.n11 drain_right.n10 60.8798
R84 drain_right.n13 drain_right.n12 60.8798
R85 drain_right.n5 drain_right.n4 60.8796
R86 drain_right.n2 drain_right.n1 60.8796
R87 drain_right drain_right.n6 32.7288
R88 drain_right drain_right.n13 6.21356
R89 drain_right.n3 drain_right.t5 2.0005
R90 drain_right.n3 drain_right.t7 2.0005
R91 drain_right.n4 drain_right.t6 2.0005
R92 drain_right.n4 drain_right.t8 2.0005
R93 drain_right.n1 drain_right.t11 2.0005
R94 drain_right.n1 drain_right.t15 2.0005
R95 drain_right.n0 drain_right.t10 2.0005
R96 drain_right.n0 drain_right.t2 2.0005
R97 drain_right.n7 drain_right.t13 2.0005
R98 drain_right.n7 drain_right.t4 2.0005
R99 drain_right.n8 drain_right.t3 2.0005
R100 drain_right.n8 drain_right.t9 2.0005
R101 drain_right.n10 drain_right.t14 2.0005
R102 drain_right.n10 drain_right.t1 2.0005
R103 drain_right.n12 drain_right.t0 2.0005
R104 drain_right.n12 drain_right.t12 2.0005
R105 drain_right.n13 drain_right.n11 0.560845
R106 drain_right.n11 drain_right.n9 0.560845
R107 drain_right.n6 drain_right.n5 0.225326
R108 drain_right.n6 drain_right.n2 0.225326
R109 source.n7 source.t1 46.201
R110 source.n8 source.t26 46.201
R111 source.n15 source.t20 46.201
R112 source.n31 source.t29 46.2008
R113 source.n24 source.t28 46.2008
R114 source.n23 source.t3 46.2008
R115 source.n16 source.t6 46.2008
R116 source.n0 source.t2 46.2008
R117 source.n2 source.n1 44.201
R118 source.n4 source.n3 44.201
R119 source.n6 source.n5 44.201
R120 source.n10 source.n9 44.201
R121 source.n12 source.n11 44.201
R122 source.n14 source.n13 44.201
R123 source.n30 source.n29 44.2008
R124 source.n28 source.n27 44.2008
R125 source.n26 source.n25 44.2008
R126 source.n22 source.n21 44.2008
R127 source.n20 source.n19 44.2008
R128 source.n18 source.n17 44.2008
R129 source.n16 source.n15 24.1208
R130 source.n32 source.n0 18.5777
R131 source.n32 source.n31 5.5436
R132 source.n29 source.t17 2.0005
R133 source.n29 source.t31 2.0005
R134 source.n27 source.t30 2.0005
R135 source.n27 source.t23 2.0005
R136 source.n25 source.t18 2.0005
R137 source.n25 source.t16 2.0005
R138 source.n21 source.t9 2.0005
R139 source.n21 source.t13 2.0005
R140 source.n19 source.t10 2.0005
R141 source.n19 source.t8 2.0005
R142 source.n17 source.t11 2.0005
R143 source.n17 source.t7 2.0005
R144 source.n1 source.t14 2.0005
R145 source.n1 source.t12 2.0005
R146 source.n3 source.t5 2.0005
R147 source.n3 source.t15 2.0005
R148 source.n5 source.t4 2.0005
R149 source.n5 source.t0 2.0005
R150 source.n9 source.t22 2.0005
R151 source.n9 source.t27 2.0005
R152 source.n11 source.t25 2.0005
R153 source.n11 source.t24 2.0005
R154 source.n13 source.t21 2.0005
R155 source.n13 source.t19 2.0005
R156 source.n15 source.n14 0.560845
R157 source.n14 source.n12 0.560845
R158 source.n12 source.n10 0.560845
R159 source.n10 source.n8 0.560845
R160 source.n7 source.n6 0.560845
R161 source.n6 source.n4 0.560845
R162 source.n4 source.n2 0.560845
R163 source.n2 source.n0 0.560845
R164 source.n18 source.n16 0.560845
R165 source.n20 source.n18 0.560845
R166 source.n22 source.n20 0.560845
R167 source.n23 source.n22 0.560845
R168 source.n26 source.n24 0.560845
R169 source.n28 source.n26 0.560845
R170 source.n30 source.n28 0.560845
R171 source.n31 source.n30 0.560845
R172 source.n8 source.n7 0.470328
R173 source.n24 source.n23 0.470328
R174 source source.n32 0.188
R175 plus.n5 plus.t6 2659.03
R176 plus.n21 plus.t5 2659.03
R177 plus.n28 plus.t7 2659.03
R178 plus.n44 plus.t3 2659.03
R179 plus.n6 plus.t13 2618.87
R180 plus.n3 plus.t11 2618.87
R181 plus.n12 plus.t8 2618.87
R182 plus.n14 plus.t15 2618.87
R183 plus.n1 plus.t12 2618.87
R184 plus.n20 plus.t10 2618.87
R185 plus.n29 plus.t14 2618.87
R186 plus.n26 plus.t1 2618.87
R187 plus.n35 plus.t4 2618.87
R188 plus.n37 plus.t9 2618.87
R189 plus.n24 plus.t0 2618.87
R190 plus.n43 plus.t2 2618.87
R191 plus.n5 plus.n4 161.489
R192 plus.n28 plus.n27 161.489
R193 plus.n7 plus.n4 161.3
R194 plus.n9 plus.n8 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n13 plus.n2 161.3
R197 plus.n16 plus.n15 161.3
R198 plus.n18 plus.n17 161.3
R199 plus.n19 plus.n0 161.3
R200 plus.n22 plus.n21 161.3
R201 plus.n30 plus.n27 161.3
R202 plus.n32 plus.n31 161.3
R203 plus.n34 plus.n33 161.3
R204 plus.n36 plus.n25 161.3
R205 plus.n39 plus.n38 161.3
R206 plus.n41 plus.n40 161.3
R207 plus.n42 plus.n23 161.3
R208 plus.n45 plus.n44 161.3
R209 plus.n8 plus.n7 73.0308
R210 plus.n19 plus.n18 73.0308
R211 plus.n42 plus.n41 73.0308
R212 plus.n31 plus.n30 73.0308
R213 plus.n11 plus.n3 69.3793
R214 plus.n15 plus.n1 69.3793
R215 plus.n38 plus.n24 69.3793
R216 plus.n34 plus.n26 69.3793
R217 plus.n6 plus.n5 54.7732
R218 plus.n21 plus.n20 54.7732
R219 plus.n44 plus.n43 54.7732
R220 plus.n29 plus.n28 54.7732
R221 plus.n13 plus.n12 47.4702
R222 plus.n14 plus.n13 47.4702
R223 plus.n37 plus.n36 47.4702
R224 plus.n36 plus.n35 47.4702
R225 plus plus.n45 31.2869
R226 plus.n12 plus.n11 25.5611
R227 plus.n15 plus.n14 25.5611
R228 plus.n38 plus.n37 25.5611
R229 plus.n35 plus.n34 25.5611
R230 plus.n7 plus.n6 18.2581
R231 plus.n20 plus.n19 18.2581
R232 plus.n43 plus.n42 18.2581
R233 plus.n30 plus.n29 18.2581
R234 plus plus.n22 13.2846
R235 plus.n8 plus.n3 3.65202
R236 plus.n18 plus.n1 3.65202
R237 plus.n41 plus.n24 3.65202
R238 plus.n31 plus.n26 3.65202
R239 plus.n9 plus.n4 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n2 0.189894
R242 plus.n16 plus.n2 0.189894
R243 plus.n17 plus.n16 0.189894
R244 plus.n17 plus.n0 0.189894
R245 plus.n22 plus.n0 0.189894
R246 plus.n45 plus.n23 0.189894
R247 plus.n40 plus.n23 0.189894
R248 plus.n40 plus.n39 0.189894
R249 plus.n39 plus.n25 0.189894
R250 plus.n33 plus.n25 0.189894
R251 plus.n33 plus.n32 0.189894
R252 plus.n32 plus.n27 0.189894
R253 drain_left.n9 drain_left.n7 61.4402
R254 drain_left.n5 drain_left.n3 61.4399
R255 drain_left.n2 drain_left.n0 61.4399
R256 drain_left.n11 drain_left.n10 60.8798
R257 drain_left.n9 drain_left.n8 60.8798
R258 drain_left.n13 drain_left.n12 60.8796
R259 drain_left.n5 drain_left.n4 60.8796
R260 drain_left.n2 drain_left.n1 60.8796
R261 drain_left drain_left.n6 33.282
R262 drain_left drain_left.n13 6.21356
R263 drain_left.n3 drain_left.t1 2.0005
R264 drain_left.n3 drain_left.t8 2.0005
R265 drain_left.n4 drain_left.t11 2.0005
R266 drain_left.n4 drain_left.t14 2.0005
R267 drain_left.n1 drain_left.t15 2.0005
R268 drain_left.n1 drain_left.t6 2.0005
R269 drain_left.n0 drain_left.t12 2.0005
R270 drain_left.n0 drain_left.t13 2.0005
R271 drain_left.n12 drain_left.t5 2.0005
R272 drain_left.n12 drain_left.t10 2.0005
R273 drain_left.n10 drain_left.t0 2.0005
R274 drain_left.n10 drain_left.t3 2.0005
R275 drain_left.n8 drain_left.t4 2.0005
R276 drain_left.n8 drain_left.t7 2.0005
R277 drain_left.n7 drain_left.t9 2.0005
R278 drain_left.n7 drain_left.t2 2.0005
R279 drain_left.n11 drain_left.n9 0.560845
R280 drain_left.n13 drain_left.n11 0.560845
R281 drain_left.n6 drain_left.n5 0.225326
R282 drain_left.n6 drain_left.n2 0.225326
C0 plus source 3.67449f
C1 minus source 3.66045f
C2 drain_right plus 0.337321f
C3 drain_left source 38.209f
C4 drain_right minus 4.29854f
C5 drain_right drain_left 0.96779f
C6 plus minus 6.04791f
C7 plus drain_left 4.48213f
C8 drain_left minus 0.170952f
C9 drain_right source 38.2094f
C10 drain_right a_n1886_n3888# 6.65322f
C11 drain_left a_n1886_n3888# 6.93547f
C12 source a_n1886_n3888# 10.405945f
C13 minus a_n1886_n3888# 7.168919f
C14 plus a_n1886_n3888# 9.540549f
C15 drain_left.t12 a_n1886_n3888# 0.507323f
C16 drain_left.t13 a_n1886_n3888# 0.507323f
C17 drain_left.n0 a_n1886_n3888# 3.37463f
C18 drain_left.t15 a_n1886_n3888# 0.507323f
C19 drain_left.t6 a_n1886_n3888# 0.507323f
C20 drain_left.n1 a_n1886_n3888# 3.37148f
C21 drain_left.n2 a_n1886_n3888# 0.647351f
C22 drain_left.t1 a_n1886_n3888# 0.507323f
C23 drain_left.t8 a_n1886_n3888# 0.507323f
C24 drain_left.n3 a_n1886_n3888# 3.37463f
C25 drain_left.t11 a_n1886_n3888# 0.507323f
C26 drain_left.t14 a_n1886_n3888# 0.507323f
C27 drain_left.n4 a_n1886_n3888# 3.37148f
C28 drain_left.n5 a_n1886_n3888# 0.647351f
C29 drain_left.n6 a_n1886_n3888# 1.59793f
C30 drain_left.t9 a_n1886_n3888# 0.507323f
C31 drain_left.t2 a_n1886_n3888# 0.507323f
C32 drain_left.n7 a_n1886_n3888# 3.37463f
C33 drain_left.t4 a_n1886_n3888# 0.507323f
C34 drain_left.t7 a_n1886_n3888# 0.507323f
C35 drain_left.n8 a_n1886_n3888# 3.37148f
C36 drain_left.n9 a_n1886_n3888# 0.674972f
C37 drain_left.t0 a_n1886_n3888# 0.507323f
C38 drain_left.t3 a_n1886_n3888# 0.507323f
C39 drain_left.n10 a_n1886_n3888# 3.37148f
C40 drain_left.n11 a_n1886_n3888# 0.333369f
C41 drain_left.t5 a_n1886_n3888# 0.507323f
C42 drain_left.t10 a_n1886_n3888# 0.507323f
C43 drain_left.n12 a_n1886_n3888# 3.37147f
C44 drain_left.n13 a_n1886_n3888# 0.569279f
C45 plus.n0 a_n1886_n3888# 0.055153f
C46 plus.t10 a_n1886_n3888# 0.350087f
C47 plus.t12 a_n1886_n3888# 0.350087f
C48 plus.n1 a_n1886_n3888# 0.142971f
C49 plus.n2 a_n1886_n3888# 0.055153f
C50 plus.t15 a_n1886_n3888# 0.350087f
C51 plus.t8 a_n1886_n3888# 0.350087f
C52 plus.t11 a_n1886_n3888# 0.350087f
C53 plus.n3 a_n1886_n3888# 0.142971f
C54 plus.n4 a_n1886_n3888# 0.117034f
C55 plus.t13 a_n1886_n3888# 0.350087f
C56 plus.t6 a_n1886_n3888# 0.352208f
C57 plus.n5 a_n1886_n3888# 0.161769f
C58 plus.n6 a_n1886_n3888# 0.142971f
C59 plus.n7 a_n1886_n3888# 0.022546f
C60 plus.n8 a_n1886_n3888# 0.019146f
C61 plus.n9 a_n1886_n3888# 0.055153f
C62 plus.n10 a_n1886_n3888# 0.055153f
C63 plus.n11 a_n1886_n3888# 0.023397f
C64 plus.n12 a_n1886_n3888# 0.142971f
C65 plus.n13 a_n1886_n3888# 0.023397f
C66 plus.n14 a_n1886_n3888# 0.142971f
C67 plus.n15 a_n1886_n3888# 0.023397f
C68 plus.n16 a_n1886_n3888# 0.055153f
C69 plus.n17 a_n1886_n3888# 0.055153f
C70 plus.n18 a_n1886_n3888# 0.019146f
C71 plus.n19 a_n1886_n3888# 0.022546f
C72 plus.n20 a_n1886_n3888# 0.142971f
C73 plus.t5 a_n1886_n3888# 0.352208f
C74 plus.n21 a_n1886_n3888# 0.161697f
C75 plus.n22 a_n1886_n3888# 0.697513f
C76 plus.n23 a_n1886_n3888# 0.055153f
C77 plus.t3 a_n1886_n3888# 0.352208f
C78 plus.t2 a_n1886_n3888# 0.350087f
C79 plus.t0 a_n1886_n3888# 0.350087f
C80 plus.n24 a_n1886_n3888# 0.142971f
C81 plus.n25 a_n1886_n3888# 0.055153f
C82 plus.t9 a_n1886_n3888# 0.350087f
C83 plus.t4 a_n1886_n3888# 0.350087f
C84 plus.t1 a_n1886_n3888# 0.350087f
C85 plus.n26 a_n1886_n3888# 0.142971f
C86 plus.n27 a_n1886_n3888# 0.117034f
C87 plus.t14 a_n1886_n3888# 0.350087f
C88 plus.t7 a_n1886_n3888# 0.352208f
C89 plus.n28 a_n1886_n3888# 0.161769f
C90 plus.n29 a_n1886_n3888# 0.142971f
C91 plus.n30 a_n1886_n3888# 0.022546f
C92 plus.n31 a_n1886_n3888# 0.019146f
C93 plus.n32 a_n1886_n3888# 0.055153f
C94 plus.n33 a_n1886_n3888# 0.055153f
C95 plus.n34 a_n1886_n3888# 0.023397f
C96 plus.n35 a_n1886_n3888# 0.142971f
C97 plus.n36 a_n1886_n3888# 0.023397f
C98 plus.n37 a_n1886_n3888# 0.142971f
C99 plus.n38 a_n1886_n3888# 0.023397f
C100 plus.n39 a_n1886_n3888# 0.055153f
C101 plus.n40 a_n1886_n3888# 0.055153f
C102 plus.n41 a_n1886_n3888# 0.019146f
C103 plus.n42 a_n1886_n3888# 0.022546f
C104 plus.n43 a_n1886_n3888# 0.142971f
C105 plus.n44 a_n1886_n3888# 0.161697f
C106 plus.n45 a_n1886_n3888# 1.76798f
C107 source.t2 a_n1886_n3888# 3.39333f
C108 source.n0 a_n1886_n3888# 1.51063f
C109 source.t14 a_n1886_n3888# 0.426164f
C110 source.t12 a_n1886_n3888# 0.426164f
C111 source.n1 a_n1886_n3888# 2.7605f
C112 source.n2 a_n1886_n3888# 0.319419f
C113 source.t5 a_n1886_n3888# 0.426164f
C114 source.t15 a_n1886_n3888# 0.426164f
C115 source.n3 a_n1886_n3888# 2.7605f
C116 source.n4 a_n1886_n3888# 0.319419f
C117 source.t4 a_n1886_n3888# 0.426164f
C118 source.t0 a_n1886_n3888# 0.426164f
C119 source.n5 a_n1886_n3888# 2.7605f
C120 source.n6 a_n1886_n3888# 0.319419f
C121 source.t1 a_n1886_n3888# 3.39333f
C122 source.n7 a_n1886_n3888# 0.446757f
C123 source.t26 a_n1886_n3888# 3.39333f
C124 source.n8 a_n1886_n3888# 0.446757f
C125 source.t22 a_n1886_n3888# 0.426164f
C126 source.t27 a_n1886_n3888# 0.426164f
C127 source.n9 a_n1886_n3888# 2.7605f
C128 source.n10 a_n1886_n3888# 0.319419f
C129 source.t25 a_n1886_n3888# 0.426164f
C130 source.t24 a_n1886_n3888# 0.426164f
C131 source.n11 a_n1886_n3888# 2.7605f
C132 source.n12 a_n1886_n3888# 0.319419f
C133 source.t21 a_n1886_n3888# 0.426164f
C134 source.t19 a_n1886_n3888# 0.426164f
C135 source.n13 a_n1886_n3888# 2.7605f
C136 source.n14 a_n1886_n3888# 0.319419f
C137 source.t20 a_n1886_n3888# 3.39333f
C138 source.n15 a_n1886_n3888# 1.90565f
C139 source.t6 a_n1886_n3888# 3.39333f
C140 source.n16 a_n1886_n3888# 1.90565f
C141 source.t11 a_n1886_n3888# 0.426164f
C142 source.t7 a_n1886_n3888# 0.426164f
C143 source.n17 a_n1886_n3888# 2.76049f
C144 source.n18 a_n1886_n3888# 0.319422f
C145 source.t10 a_n1886_n3888# 0.426164f
C146 source.t8 a_n1886_n3888# 0.426164f
C147 source.n19 a_n1886_n3888# 2.76049f
C148 source.n20 a_n1886_n3888# 0.319422f
C149 source.t9 a_n1886_n3888# 0.426164f
C150 source.t13 a_n1886_n3888# 0.426164f
C151 source.n21 a_n1886_n3888# 2.76049f
C152 source.n22 a_n1886_n3888# 0.319422f
C153 source.t3 a_n1886_n3888# 3.39333f
C154 source.n23 a_n1886_n3888# 0.446761f
C155 source.t28 a_n1886_n3888# 3.39333f
C156 source.n24 a_n1886_n3888# 0.446761f
C157 source.t18 a_n1886_n3888# 0.426164f
C158 source.t16 a_n1886_n3888# 0.426164f
C159 source.n25 a_n1886_n3888# 2.76049f
C160 source.n26 a_n1886_n3888# 0.319422f
C161 source.t30 a_n1886_n3888# 0.426164f
C162 source.t23 a_n1886_n3888# 0.426164f
C163 source.n27 a_n1886_n3888# 2.76049f
C164 source.n28 a_n1886_n3888# 0.319422f
C165 source.t17 a_n1886_n3888# 0.426164f
C166 source.t31 a_n1886_n3888# 0.426164f
C167 source.n29 a_n1886_n3888# 2.76049f
C168 source.n30 a_n1886_n3888# 0.319422f
C169 source.t29 a_n1886_n3888# 3.39333f
C170 source.n31 a_n1886_n3888# 0.581763f
C171 source.n32 a_n1886_n3888# 1.73579f
C172 drain_right.t10 a_n1886_n3888# 0.506257f
C173 drain_right.t2 a_n1886_n3888# 0.506257f
C174 drain_right.n0 a_n1886_n3888# 3.36753f
C175 drain_right.t11 a_n1886_n3888# 0.506257f
C176 drain_right.t15 a_n1886_n3888# 0.506257f
C177 drain_right.n1 a_n1886_n3888# 3.3644f
C178 drain_right.n2 a_n1886_n3888# 0.64599f
C179 drain_right.t5 a_n1886_n3888# 0.506257f
C180 drain_right.t7 a_n1886_n3888# 0.506257f
C181 drain_right.n3 a_n1886_n3888# 3.36753f
C182 drain_right.t6 a_n1886_n3888# 0.506257f
C183 drain_right.t8 a_n1886_n3888# 0.506257f
C184 drain_right.n4 a_n1886_n3888# 3.3644f
C185 drain_right.n5 a_n1886_n3888# 0.64599f
C186 drain_right.n6 a_n1886_n3888# 1.53595f
C187 drain_right.t13 a_n1886_n3888# 0.506257f
C188 drain_right.t4 a_n1886_n3888# 0.506257f
C189 drain_right.n7 a_n1886_n3888# 3.36753f
C190 drain_right.t3 a_n1886_n3888# 0.506257f
C191 drain_right.t9 a_n1886_n3888# 0.506257f
C192 drain_right.n8 a_n1886_n3888# 3.3644f
C193 drain_right.n9 a_n1886_n3888# 0.673564f
C194 drain_right.t14 a_n1886_n3888# 0.506257f
C195 drain_right.t1 a_n1886_n3888# 0.506257f
C196 drain_right.n10 a_n1886_n3888# 3.3644f
C197 drain_right.n11 a_n1886_n3888# 0.332669f
C198 drain_right.t0 a_n1886_n3888# 0.506257f
C199 drain_right.t12 a_n1886_n3888# 0.506257f
C200 drain_right.n12 a_n1886_n3888# 3.3644f
C201 drain_right.n13 a_n1886_n3888# 0.568072f
C202 minus.n0 a_n1886_n3888# 0.053952f
C203 minus.t11 a_n1886_n3888# 0.344541f
C204 minus.t10 a_n1886_n3888# 0.342466f
C205 minus.t12 a_n1886_n3888# 0.342466f
C206 minus.n1 a_n1886_n3888# 0.139859f
C207 minus.n2 a_n1886_n3888# 0.053952f
C208 minus.t6 a_n1886_n3888# 0.342466f
C209 minus.t7 a_n1886_n3888# 0.342466f
C210 minus.t9 a_n1886_n3888# 0.342466f
C211 minus.n3 a_n1886_n3888# 0.139859f
C212 minus.n4 a_n1886_n3888# 0.114486f
C213 minus.t4 a_n1886_n3888# 0.342466f
C214 minus.t5 a_n1886_n3888# 0.344541f
C215 minus.n5 a_n1886_n3888# 0.158248f
C216 minus.n6 a_n1886_n3888# 0.139859f
C217 minus.n7 a_n1886_n3888# 0.022056f
C218 minus.n8 a_n1886_n3888# 0.018729f
C219 minus.n9 a_n1886_n3888# 0.053952f
C220 minus.n10 a_n1886_n3888# 0.053952f
C221 minus.n11 a_n1886_n3888# 0.022887f
C222 minus.n12 a_n1886_n3888# 0.139859f
C223 minus.n13 a_n1886_n3888# 0.022887f
C224 minus.n14 a_n1886_n3888# 0.139859f
C225 minus.n15 a_n1886_n3888# 0.022887f
C226 minus.n16 a_n1886_n3888# 0.053952f
C227 minus.n17 a_n1886_n3888# 0.053952f
C228 minus.n18 a_n1886_n3888# 0.018729f
C229 minus.n19 a_n1886_n3888# 0.022056f
C230 minus.n20 a_n1886_n3888# 0.139859f
C231 minus.n21 a_n1886_n3888# 0.158177f
C232 minus.n22 a_n1886_n3888# 2.10111f
C233 minus.n23 a_n1886_n3888# 0.053952f
C234 minus.t0 a_n1886_n3888# 0.342466f
C235 minus.t14 a_n1886_n3888# 0.342466f
C236 minus.n24 a_n1886_n3888# 0.139859f
C237 minus.n25 a_n1886_n3888# 0.053952f
C238 minus.t8 a_n1886_n3888# 0.342466f
C239 minus.t1 a_n1886_n3888# 0.342466f
C240 minus.t15 a_n1886_n3888# 0.342466f
C241 minus.n26 a_n1886_n3888# 0.139859f
C242 minus.n27 a_n1886_n3888# 0.114486f
C243 minus.t13 a_n1886_n3888# 0.342466f
C244 minus.t3 a_n1886_n3888# 0.344541f
C245 minus.n28 a_n1886_n3888# 0.158248f
C246 minus.n29 a_n1886_n3888# 0.139859f
C247 minus.n30 a_n1886_n3888# 0.022056f
C248 minus.n31 a_n1886_n3888# 0.018729f
C249 minus.n32 a_n1886_n3888# 0.053952f
C250 minus.n33 a_n1886_n3888# 0.053952f
C251 minus.n34 a_n1886_n3888# 0.022887f
C252 minus.n35 a_n1886_n3888# 0.139859f
C253 minus.n36 a_n1886_n3888# 0.022887f
C254 minus.n37 a_n1886_n3888# 0.139859f
C255 minus.n38 a_n1886_n3888# 0.022887f
C256 minus.n39 a_n1886_n3888# 0.053952f
C257 minus.n40 a_n1886_n3888# 0.053952f
C258 minus.n41 a_n1886_n3888# 0.018729f
C259 minus.n42 a_n1886_n3888# 0.022056f
C260 minus.n43 a_n1886_n3888# 0.139859f
C261 minus.t2 a_n1886_n3888# 0.344541f
C262 minus.n44 a_n1886_n3888# 0.158177f
C263 minus.n45 a_n1886_n3888# 0.35327f
C264 minus.n46 a_n1886_n3888# 2.53441f
.ends

