* NGSPICE file created from diffpair87.ext - technology: sky130A

.subckt diffpair87 minus drain_right drain_left source plus
X0 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X5 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X6 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X7 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X8 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X9 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X10 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X12 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X14 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X18 a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X19 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X20 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X21 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X22 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X24 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X25 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X26 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X27 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X28 source minus drain_right a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X29 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X30 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X31 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X32 drain_right minus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X33 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X34 drain_left plus source a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X35 source plus drain_left a_n1886_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
.ends

