* NGSPICE file created from diffpair234.ext - technology: sky130A

.subckt diffpair234 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t12 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X1 drain_left.t9 plus.t0 source.t1 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X2 a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X3 drain_right.t8 minus.t1 source.t19 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X4 a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X5 drain_right.t7 minus.t2 source.t18 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X6 drain_left.t8 plus.t1 source.t7 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X7 drain_left.t7 plus.t2 source.t9 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X8 a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X9 drain_right.t6 minus.t3 source.t17 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X10 source.t16 minus.t4 drain_right.t5 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X11 source.t13 minus.t5 drain_right.t4 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X12 source.t14 minus.t6 drain_right.t3 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X13 drain_right.t2 minus.t7 source.t11 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X14 source.t4 plus.t3 drain_left.t6 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X15 source.t15 minus.t8 drain_right.t1 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X16 source.t8 plus.t4 drain_left.t5 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X17 drain_right.t0 minus.t9 source.t10 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X18 source.t5 plus.t5 drain_left.t4 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 drain_left.t3 plus.t6 source.t3 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X20 a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X21 drain_left.t2 plus.t7 source.t6 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X22 source.t0 plus.t8 drain_left.t1 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X23 drain_left.t0 plus.t9 source.t2 a_n2072_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
R0 minus.n3 minus.t7 162.675
R1 minus.n13 minus.t1 162.675
R2 minus.n9 minus.n8 161.3
R3 minus.n7 minus.n0 161.3
R4 minus.n19 minus.n18 161.3
R5 minus.n17 minus.n10 161.3
R6 minus.n2 minus.t5 139.48
R7 minus.n1 minus.t3 139.48
R8 minus.n6 minus.t8 139.48
R9 minus.n8 minus.t9 139.48
R10 minus.n12 minus.t4 139.48
R11 minus.n11 minus.t2 139.48
R12 minus.n16 minus.t6 139.48
R13 minus.n18 minus.t0 139.48
R14 minus.n6 minus.n5 80.6037
R15 minus.n4 minus.n1 80.6037
R16 minus.n16 minus.n15 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n7 minus.n6 32.1338
R23 minus.n17 minus.n16 32.1338
R24 minus.n4 minus.n3 31.8629
R25 minus.n14 minus.n13 31.8629
R26 minus.n20 minus.n9 30.3282
R27 minus.n3 minus.n2 16.2333
R28 minus.n13 minus.n12 16.2333
R29 minus.n8 minus.n7 16.0672
R30 minus.n18 minus.n17 16.0672
R31 minus.n20 minus.n19 6.67664
R32 minus.n5 minus.n4 0.380177
R33 minus.n15 minus.n14 0.380177
R34 minus.n5 minus.n0 0.285035
R35 minus.n15 minus.n10 0.285035
R36 minus.n9 minus.n0 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 source.n0 source.t6 69.6943
R40 source.n5 source.t11 69.6943
R41 source.n19 source.t12 69.6942
R42 source.n14 source.t7 69.6942
R43 source.n2 source.n1 63.0943
R44 source.n4 source.n3 63.0943
R45 source.n7 source.n6 63.0943
R46 source.n9 source.n8 63.0943
R47 source.n18 source.n17 63.0942
R48 source.n16 source.n15 63.0942
R49 source.n13 source.n12 63.0942
R50 source.n11 source.n10 63.0942
R51 source.n11 source.n9 16.4178
R52 source.n20 source.n0 9.69368
R53 source.n17 source.t18 6.6005
R54 source.n17 source.t14 6.6005
R55 source.n15 source.t19 6.6005
R56 source.n15 source.t16 6.6005
R57 source.n12 source.t9 6.6005
R58 source.n12 source.t4 6.6005
R59 source.n10 source.t1 6.6005
R60 source.n10 source.t8 6.6005
R61 source.n1 source.t3 6.6005
R62 source.n1 source.t5 6.6005
R63 source.n3 source.t2 6.6005
R64 source.n3 source.t0 6.6005
R65 source.n6 source.t17 6.6005
R66 source.n6 source.t13 6.6005
R67 source.n8 source.t10 6.6005
R68 source.n8 source.t15 6.6005
R69 source.n20 source.n19 5.7505
R70 source.n9 source.n7 0.974638
R71 source.n7 source.n5 0.974638
R72 source.n4 source.n2 0.974638
R73 source.n2 source.n0 0.974638
R74 source.n13 source.n11 0.974638
R75 source.n14 source.n13 0.974638
R76 source.n18 source.n16 0.974638
R77 source.n19 source.n18 0.974638
R78 source.n5 source.n4 0.957397
R79 source.n16 source.n14 0.957397
R80 source source.n20 0.188
R81 drain_right.n1 drain_right.t8 87.3471
R82 drain_right.n7 drain_right.t0 86.3731
R83 drain_right.n6 drain_right.n4 80.7472
R84 drain_right.n3 drain_right.n2 80.4483
R85 drain_right.n6 drain_right.n5 79.7731
R86 drain_right.n1 drain_right.n0 79.773
R87 drain_right drain_right.n3 24.1358
R88 drain_right.n2 drain_right.t3 6.6005
R89 drain_right.n2 drain_right.t9 6.6005
R90 drain_right.n0 drain_right.t5 6.6005
R91 drain_right.n0 drain_right.t7 6.6005
R92 drain_right.n4 drain_right.t4 6.6005
R93 drain_right.n4 drain_right.t2 6.6005
R94 drain_right.n5 drain_right.t1 6.6005
R95 drain_right.n5 drain_right.t6 6.6005
R96 drain_right drain_right.n7 6.14028
R97 drain_right.n7 drain_right.n6 0.974638
R98 drain_right.n3 drain_right.n1 0.188688
R99 plus.n3 plus.t9 162.675
R100 plus.n13 plus.t1 162.675
R101 plus.n7 plus.n0 161.3
R102 plus.n9 plus.n8 161.3
R103 plus.n17 plus.n10 161.3
R104 plus.n19 plus.n18 161.3
R105 plus.n8 plus.t7 139.48
R106 plus.n6 plus.t5 139.48
R107 plus.n5 plus.t6 139.48
R108 plus.n4 plus.t8 139.48
R109 plus.n18 plus.t0 139.48
R110 plus.n16 plus.t4 139.48
R111 plus.n15 plus.t2 139.48
R112 plus.n14 plus.t3 139.48
R113 plus.n5 plus.n2 80.6037
R114 plus.n6 plus.n1 80.6037
R115 plus.n15 plus.n12 80.6037
R116 plus.n16 plus.n11 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n7 plus.n6 32.1338
R122 plus.n17 plus.n16 32.1338
R123 plus.n3 plus.n2 31.8629
R124 plus.n13 plus.n12 31.8629
R125 plus plus.n19 27.6183
R126 plus.n4 plus.n3 16.2333
R127 plus.n14 plus.n13 16.2333
R128 plus.n8 plus.n7 16.0672
R129 plus.n18 plus.n17 16.0672
R130 plus plus.n9 8.91148
R131 plus.n2 plus.n1 0.380177
R132 plus.n12 plus.n11 0.380177
R133 plus.n1 plus.n0 0.285035
R134 plus.n11 plus.n10 0.285035
R135 plus.n9 plus.n0 0.189894
R136 plus.n19 plus.n10 0.189894
R137 drain_left.n5 drain_left.t0 87.3472
R138 drain_left.n1 drain_left.t9 87.3471
R139 drain_left.n3 drain_left.n2 80.4483
R140 drain_left.n7 drain_left.n6 79.7731
R141 drain_left.n5 drain_left.n4 79.7731
R142 drain_left.n1 drain_left.n0 79.773
R143 drain_left drain_left.n3 24.689
R144 drain_left drain_left.n7 6.62735
R145 drain_left.n2 drain_left.t6 6.6005
R146 drain_left.n2 drain_left.t8 6.6005
R147 drain_left.n0 drain_left.t5 6.6005
R148 drain_left.n0 drain_left.t7 6.6005
R149 drain_left.n6 drain_left.t4 6.6005
R150 drain_left.n6 drain_left.t2 6.6005
R151 drain_left.n4 drain_left.t1 6.6005
R152 drain_left.n4 drain_left.t3 6.6005
R153 drain_left.n7 drain_left.n5 0.974638
R154 drain_left.n3 drain_left.n1 0.188688
C0 drain_right plus 0.364576f
C1 drain_left drain_right 1.03121f
C2 minus source 2.47786f
C3 plus minus 4.06428f
C4 plus source 2.49197f
C5 drain_left minus 0.177583f
C6 drain_right minus 2.12886f
C7 drain_left source 5.41115f
C8 drain_right source 5.41097f
C9 drain_left plus 2.33099f
C10 drain_right a_n2072_n1488# 4.51396f
C11 drain_left a_n2072_n1488# 4.83873f
C12 source a_n2072_n1488# 3.08638f
C13 minus a_n2072_n1488# 7.381784f
C14 plus a_n2072_n1488# 8.612939f
C15 drain_left.t9 a_n2072_n1488# 0.535561f
C16 drain_left.t5 a_n2072_n1488# 0.057476f
C17 drain_left.t7 a_n2072_n1488# 0.057476f
C18 drain_left.n0 a_n2072_n1488# 0.414509f
C19 drain_left.n1 a_n2072_n1488# 0.603498f
C20 drain_left.t6 a_n2072_n1488# 0.057476f
C21 drain_left.t8 a_n2072_n1488# 0.057476f
C22 drain_left.n2 a_n2072_n1488# 0.417309f
C23 drain_left.n3 a_n2072_n1488# 1.1459f
C24 drain_left.t0 a_n2072_n1488# 0.535563f
C25 drain_left.t1 a_n2072_n1488# 0.057476f
C26 drain_left.t3 a_n2072_n1488# 0.057476f
C27 drain_left.n4 a_n2072_n1488# 0.414511f
C28 drain_left.n5 a_n2072_n1488# 0.661906f
C29 drain_left.t4 a_n2072_n1488# 0.057476f
C30 drain_left.t2 a_n2072_n1488# 0.057476f
C31 drain_left.n6 a_n2072_n1488# 0.414511f
C32 drain_left.n7 a_n2072_n1488# 0.563668f
C33 plus.n0 a_n2072_n1488# 0.059815f
C34 plus.t7 a_n2072_n1488# 0.322605f
C35 plus.t5 a_n2072_n1488# 0.322605f
C36 plus.n1 a_n2072_n1488# 0.074664f
C37 plus.t6 a_n2072_n1488# 0.322605f
C38 plus.n2 a_n2072_n1488# 0.275086f
C39 plus.t8 a_n2072_n1488# 0.322605f
C40 plus.t9 a_n2072_n1488# 0.349292f
C41 plus.n3 a_n2072_n1488# 0.165554f
C42 plus.n4 a_n2072_n1488# 0.196475f
C43 plus.n5 a_n2072_n1488# 0.197559f
C44 plus.n6 a_n2072_n1488# 0.194519f
C45 plus.n7 a_n2072_n1488# 0.010172f
C46 plus.n8 a_n2072_n1488# 0.181307f
C47 plus.n9 a_n2072_n1488# 0.354347f
C48 plus.n10 a_n2072_n1488# 0.059815f
C49 plus.t0 a_n2072_n1488# 0.322605f
C50 plus.n11 a_n2072_n1488# 0.074664f
C51 plus.t4 a_n2072_n1488# 0.322605f
C52 plus.n12 a_n2072_n1488# 0.275086f
C53 plus.t2 a_n2072_n1488# 0.322605f
C54 plus.t1 a_n2072_n1488# 0.349292f
C55 plus.n13 a_n2072_n1488# 0.165554f
C56 plus.t3 a_n2072_n1488# 0.322605f
C57 plus.n14 a_n2072_n1488# 0.196475f
C58 plus.n15 a_n2072_n1488# 0.197559f
C59 plus.n16 a_n2072_n1488# 0.194519f
C60 plus.n17 a_n2072_n1488# 0.010172f
C61 plus.n18 a_n2072_n1488# 0.181307f
C62 plus.n19 a_n2072_n1488# 1.12389f
C63 drain_right.t8 a_n2072_n1488# 0.528156f
C64 drain_right.t5 a_n2072_n1488# 0.056681f
C65 drain_right.t7 a_n2072_n1488# 0.056681f
C66 drain_right.n0 a_n2072_n1488# 0.408778f
C67 drain_right.n1 a_n2072_n1488# 0.595153f
C68 drain_right.t3 a_n2072_n1488# 0.056681f
C69 drain_right.t9 a_n2072_n1488# 0.056681f
C70 drain_right.n2 a_n2072_n1488# 0.411539f
C71 drain_right.n3 a_n2072_n1488# 1.0828f
C72 drain_right.t4 a_n2072_n1488# 0.056681f
C73 drain_right.t2 a_n2072_n1488# 0.056681f
C74 drain_right.n4 a_n2072_n1488# 0.413016f
C75 drain_right.t1 a_n2072_n1488# 0.056681f
C76 drain_right.t6 a_n2072_n1488# 0.056681f
C77 drain_right.n5 a_n2072_n1488# 0.40878f
C78 drain_right.n6 a_n2072_n1488# 0.688359f
C79 drain_right.t0 a_n2072_n1488# 0.524647f
C80 drain_right.n7 a_n2072_n1488# 0.539527f
C81 source.t6 a_n2072_n1488# 0.591854f
C82 source.n0 a_n2072_n1488# 0.880788f
C83 source.t3 a_n2072_n1488# 0.071275f
C84 source.t5 a_n2072_n1488# 0.071275f
C85 source.n1 a_n2072_n1488# 0.451924f
C86 source.n2 a_n2072_n1488# 0.450647f
C87 source.t2 a_n2072_n1488# 0.071275f
C88 source.t0 a_n2072_n1488# 0.071275f
C89 source.n3 a_n2072_n1488# 0.451924f
C90 source.n4 a_n2072_n1488# 0.448977f
C91 source.t11 a_n2072_n1488# 0.591854f
C92 source.n5 a_n2072_n1488# 0.503433f
C93 source.t17 a_n2072_n1488# 0.071275f
C94 source.t13 a_n2072_n1488# 0.071275f
C95 source.n6 a_n2072_n1488# 0.451924f
C96 source.n7 a_n2072_n1488# 0.450647f
C97 source.t10 a_n2072_n1488# 0.071275f
C98 source.t15 a_n2072_n1488# 0.071275f
C99 source.n8 a_n2072_n1488# 0.451924f
C100 source.n9 a_n2072_n1488# 1.2443f
C101 source.t1 a_n2072_n1488# 0.071275f
C102 source.t8 a_n2072_n1488# 0.071275f
C103 source.n10 a_n2072_n1488# 0.451921f
C104 source.n11 a_n2072_n1488# 1.24431f
C105 source.t9 a_n2072_n1488# 0.071275f
C106 source.t4 a_n2072_n1488# 0.071275f
C107 source.n12 a_n2072_n1488# 0.451921f
C108 source.n13 a_n2072_n1488# 0.45065f
C109 source.t7 a_n2072_n1488# 0.591851f
C110 source.n14 a_n2072_n1488# 0.503436f
C111 source.t19 a_n2072_n1488# 0.071275f
C112 source.t16 a_n2072_n1488# 0.071275f
C113 source.n15 a_n2072_n1488# 0.451921f
C114 source.n16 a_n2072_n1488# 0.44898f
C115 source.t18 a_n2072_n1488# 0.071275f
C116 source.t14 a_n2072_n1488# 0.071275f
C117 source.n17 a_n2072_n1488# 0.451921f
C118 source.n18 a_n2072_n1488# 0.45065f
C119 source.t12 a_n2072_n1488# 0.591851f
C120 source.n19 a_n2072_n1488# 0.658874f
C121 source.n20 a_n2072_n1488# 0.890504f
C122 minus.n0 a_n2072_n1488# 0.057882f
C123 minus.t3 a_n2072_n1488# 0.312176f
C124 minus.n1 a_n2072_n1488# 0.191173f
C125 minus.t8 a_n2072_n1488# 0.312176f
C126 minus.t7 a_n2072_n1488# 0.338f
C127 minus.t5 a_n2072_n1488# 0.312176f
C128 minus.n2 a_n2072_n1488# 0.190123f
C129 minus.n3 a_n2072_n1488# 0.160202f
C130 minus.n4 a_n2072_n1488# 0.266193f
C131 minus.n5 a_n2072_n1488# 0.072251f
C132 minus.n6 a_n2072_n1488# 0.188231f
C133 minus.n7 a_n2072_n1488# 0.009843f
C134 minus.t9 a_n2072_n1488# 0.312176f
C135 minus.n8 a_n2072_n1488# 0.175446f
C136 minus.n9 a_n2072_n1488# 1.15658f
C137 minus.n10 a_n2072_n1488# 0.057882f
C138 minus.t2 a_n2072_n1488# 0.312176f
C139 minus.n11 a_n2072_n1488# 0.191173f
C140 minus.t1 a_n2072_n1488# 0.338f
C141 minus.t4 a_n2072_n1488# 0.312176f
C142 minus.n12 a_n2072_n1488# 0.190123f
C143 minus.n13 a_n2072_n1488# 0.160202f
C144 minus.n14 a_n2072_n1488# 0.266193f
C145 minus.n15 a_n2072_n1488# 0.072251f
C146 minus.t6 a_n2072_n1488# 0.312176f
C147 minus.n16 a_n2072_n1488# 0.188231f
C148 minus.n17 a_n2072_n1488# 0.009843f
C149 minus.t0 a_n2072_n1488# 0.312176f
C150 minus.n18 a_n2072_n1488# 0.175446f
C151 minus.n19 a_n2072_n1488# 0.301494f
C152 minus.n20 a_n2072_n1488# 1.41735f
.ends

