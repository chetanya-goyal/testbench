* NGSPICE file created from diffpair609.ext - technology: sky130A

.subckt diffpair609 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t29 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t28 plus.t1 drain_left.t22 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X3 drain_right.t23 minus.t0 source.t17 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X4 drain_left.t21 plus.t2 source.t40 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X5 source.t39 plus.t3 drain_left.t20 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t38 plus.t4 drain_left.t19 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X7 source.t14 minus.t1 drain_right.t22 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 source.t19 minus.t2 drain_right.t21 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X9 source.t23 plus.t5 drain_left.t18 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 drain_right.t20 minus.t3 source.t3 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X11 source.t37 plus.t6 drain_left.t17 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X12 drain_left.t16 plus.t7 source.t32 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X13 source.t31 plus.t8 drain_left.t15 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X14 source.t8 minus.t4 drain_right.t19 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 drain_right.t18 minus.t5 source.t4 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X16 source.t7 minus.t6 drain_right.t17 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X17 drain_right.t16 minus.t7 source.t21 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X18 drain_left.t14 plus.t9 source.t30 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 drain_right.t15 minus.t8 source.t20 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X20 source.t10 minus.t9 drain_right.t14 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X21 drain_left.t13 plus.t10 source.t41 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X22 drain_left.t12 plus.t11 source.t27 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 drain_left.t11 plus.t12 source.t22 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X24 source.t26 plus.t13 drain_left.t10 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X25 source.t9 minus.t10 drain_right.t13 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X26 drain_right.t12 minus.t11 source.t46 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X27 a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X28 source.t47 minus.t12 drain_right.t11 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X29 drain_left.t9 plus.t14 source.t25 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X30 source.t42 plus.t15 drain_left.t8 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X31 source.t44 plus.t16 drain_left.t7 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X32 drain_right.t10 minus.t13 source.t5 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X33 drain_left.t6 plus.t17 source.t43 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X34 drain_right.t9 minus.t14 source.t18 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X35 drain_right.t8 minus.t15 source.t1 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X36 a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X37 source.t12 minus.t16 drain_right.t7 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X38 source.t16 minus.t17 drain_right.t6 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X39 drain_left.t5 plus.t18 source.t45 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X40 drain_right.t5 minus.t18 source.t6 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X41 source.t11 minus.t19 drain_right.t4 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X42 drain_right.t3 minus.t20 source.t15 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X43 source.t0 minus.t21 drain_right.t2 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X44 source.t24 plus.t19 drain_left.t4 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X45 a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X46 source.t2 minus.t22 drain_right.t1 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X47 drain_right.t0 minus.t23 source.t13 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X48 drain_left.t3 plus.t20 source.t36 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X49 source.t35 plus.t21 drain_left.t2 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X50 source.t34 plus.t22 drain_left.t1 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X51 drain_left.t0 plus.t23 source.t33 a_n2874_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
R0 plus.n11 plus.t8 1068.92
R1 plus.n45 plus.t0 1068.92
R2 plus.n32 plus.t2 1042.57
R3 plus.n30 plus.t3 1042.57
R4 plus.n29 plus.t17 1042.57
R5 plus.n3 plus.t5 1042.57
R6 plus.n23 plus.t20 1042.57
R7 plus.n22 plus.t13 1042.57
R8 plus.n6 plus.t23 1042.57
R9 plus.n17 plus.t19 1042.57
R10 plus.n15 plus.t10 1042.57
R11 plus.n9 plus.t21 1042.57
R12 plus.n10 plus.t18 1042.57
R13 plus.n66 plus.t22 1042.57
R14 plus.n64 plus.t9 1042.57
R15 plus.n63 plus.t15 1042.57
R16 plus.n37 plus.t14 1042.57
R17 plus.n57 plus.t4 1042.57
R18 plus.n56 plus.t11 1042.57
R19 plus.n40 plus.t16 1042.57
R20 plus.n51 plus.t7 1042.57
R21 plus.n49 plus.t6 1042.57
R22 plus.n43 plus.t12 1042.57
R23 plus.n44 plus.t1 1042.57
R24 plus.n12 plus.n9 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n15 plus.n8 161.3
R27 plus.n16 plus.n7 161.3
R28 plus.n18 plus.n17 161.3
R29 plus.n19 plus.n6 161.3
R30 plus.n21 plus.n20 161.3
R31 plus.n22 plus.n5 161.3
R32 plus.n23 plus.n4 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n26 plus.n3 161.3
R35 plus.n28 plus.n27 161.3
R36 plus.n29 plus.n2 161.3
R37 plus.n30 plus.n1 161.3
R38 plus.n31 plus.n0 161.3
R39 plus.n33 plus.n32 161.3
R40 plus.n46 plus.n43 161.3
R41 plus.n48 plus.n47 161.3
R42 plus.n49 plus.n42 161.3
R43 plus.n50 plus.n41 161.3
R44 plus.n52 plus.n51 161.3
R45 plus.n53 plus.n40 161.3
R46 plus.n55 plus.n54 161.3
R47 plus.n56 plus.n39 161.3
R48 plus.n57 plus.n38 161.3
R49 plus.n59 plus.n58 161.3
R50 plus.n60 plus.n37 161.3
R51 plus.n62 plus.n61 161.3
R52 plus.n63 plus.n36 161.3
R53 plus.n64 plus.n35 161.3
R54 plus.n65 plus.n34 161.3
R55 plus.n67 plus.n66 161.3
R56 plus.n30 plus.n29 48.2005
R57 plus.n23 plus.n22 48.2005
R58 plus.n17 plus.n6 48.2005
R59 plus.n10 plus.n9 48.2005
R60 plus.n64 plus.n63 48.2005
R61 plus.n57 plus.n56 48.2005
R62 plus.n51 plus.n40 48.2005
R63 plus.n44 plus.n43 48.2005
R64 plus.n24 plus.n3 47.4702
R65 plus.n16 plus.n15 47.4702
R66 plus.n58 plus.n37 47.4702
R67 plus.n50 plus.n49 47.4702
R68 plus.n32 plus.n31 46.0096
R69 plus.n66 plus.n65 46.0096
R70 plus.n12 plus.n11 45.0871
R71 plus.n46 plus.n45 45.0871
R72 plus plus.n67 36.946
R73 plus.n28 plus.n3 25.5611
R74 plus.n15 plus.n14 25.5611
R75 plus.n62 plus.n37 25.5611
R76 plus.n49 plus.n48 25.5611
R77 plus.n21 plus.n6 24.1005
R78 plus.n22 plus.n21 24.1005
R79 plus.n56 plus.n55 24.1005
R80 plus.n55 plus.n40 24.1005
R81 plus.n29 plus.n28 22.6399
R82 plus.n14 plus.n9 22.6399
R83 plus.n63 plus.n62 22.6399
R84 plus.n48 plus.n43 22.6399
R85 plus plus.n33 15.2013
R86 plus.n11 plus.n10 14.1472
R87 plus.n45 plus.n44 14.1472
R88 plus.n31 plus.n30 2.19141
R89 plus.n65 plus.n64 2.19141
R90 plus.n24 plus.n23 0.730803
R91 plus.n17 plus.n16 0.730803
R92 plus.n58 plus.n57 0.730803
R93 plus.n51 plus.n50 0.730803
R94 plus.n13 plus.n12 0.189894
R95 plus.n13 plus.n8 0.189894
R96 plus.n8 plus.n7 0.189894
R97 plus.n18 plus.n7 0.189894
R98 plus.n19 plus.n18 0.189894
R99 plus.n20 plus.n19 0.189894
R100 plus.n20 plus.n5 0.189894
R101 plus.n5 plus.n4 0.189894
R102 plus.n25 plus.n4 0.189894
R103 plus.n26 plus.n25 0.189894
R104 plus.n27 plus.n26 0.189894
R105 plus.n27 plus.n2 0.189894
R106 plus.n2 plus.n1 0.189894
R107 plus.n1 plus.n0 0.189894
R108 plus.n33 plus.n0 0.189894
R109 plus.n67 plus.n34 0.189894
R110 plus.n35 plus.n34 0.189894
R111 plus.n36 plus.n35 0.189894
R112 plus.n61 plus.n36 0.189894
R113 plus.n61 plus.n60 0.189894
R114 plus.n60 plus.n59 0.189894
R115 plus.n59 plus.n38 0.189894
R116 plus.n39 plus.n38 0.189894
R117 plus.n54 plus.n39 0.189894
R118 plus.n54 plus.n53 0.189894
R119 plus.n53 plus.n52 0.189894
R120 plus.n52 plus.n41 0.189894
R121 plus.n42 plus.n41 0.189894
R122 plus.n47 plus.n42 0.189894
R123 plus.n47 plus.n46 0.189894
R124 source.n0 source.t40 44.1297
R125 source.n11 source.t31 44.1296
R126 source.n12 source.t18 44.1296
R127 source.n23 source.t2 44.1296
R128 source.n47 source.t3 44.1295
R129 source.n36 source.t7 44.1295
R130 source.n35 source.t29 44.1295
R131 source.n24 source.t34 44.1295
R132 source.n2 source.n1 43.1397
R133 source.n4 source.n3 43.1397
R134 source.n6 source.n5 43.1397
R135 source.n8 source.n7 43.1397
R136 source.n10 source.n9 43.1397
R137 source.n14 source.n13 43.1397
R138 source.n16 source.n15 43.1397
R139 source.n18 source.n17 43.1397
R140 source.n20 source.n19 43.1397
R141 source.n22 source.n21 43.1397
R142 source.n46 source.n45 43.1396
R143 source.n44 source.n43 43.1396
R144 source.n42 source.n41 43.1396
R145 source.n40 source.n39 43.1396
R146 source.n38 source.n37 43.1396
R147 source.n34 source.n33 43.1396
R148 source.n32 source.n31 43.1396
R149 source.n30 source.n29 43.1396
R150 source.n28 source.n27 43.1396
R151 source.n26 source.n25 43.1396
R152 source.n24 source.n23 28.0638
R153 source.n48 source.n0 22.4432
R154 source.n48 source.n47 5.62119
R155 source.n45 source.t13 0.9905
R156 source.n45 source.t12 0.9905
R157 source.n43 source.t46 0.9905
R158 source.n43 source.t19 0.9905
R159 source.n41 source.t15 0.9905
R160 source.n41 source.t11 0.9905
R161 source.n39 source.t5 0.9905
R162 source.n39 source.t10 0.9905
R163 source.n37 source.t4 0.9905
R164 source.n37 source.t16 0.9905
R165 source.n33 source.t22 0.9905
R166 source.n33 source.t28 0.9905
R167 source.n31 source.t32 0.9905
R168 source.n31 source.t37 0.9905
R169 source.n29 source.t27 0.9905
R170 source.n29 source.t44 0.9905
R171 source.n27 source.t25 0.9905
R172 source.n27 source.t38 0.9905
R173 source.n25 source.t30 0.9905
R174 source.n25 source.t42 0.9905
R175 source.n1 source.t43 0.9905
R176 source.n1 source.t39 0.9905
R177 source.n3 source.t36 0.9905
R178 source.n3 source.t23 0.9905
R179 source.n5 source.t33 0.9905
R180 source.n5 source.t26 0.9905
R181 source.n7 source.t41 0.9905
R182 source.n7 source.t24 0.9905
R183 source.n9 source.t45 0.9905
R184 source.n9 source.t35 0.9905
R185 source.n13 source.t20 0.9905
R186 source.n13 source.t14 0.9905
R187 source.n15 source.t21 0.9905
R188 source.n15 source.t0 0.9905
R189 source.n17 source.t17 0.9905
R190 source.n17 source.t9 0.9905
R191 source.n19 source.t6 0.9905
R192 source.n19 source.t47 0.9905
R193 source.n21 source.t1 0.9905
R194 source.n21 source.t8 0.9905
R195 source.n23 source.n22 0.716017
R196 source.n22 source.n20 0.716017
R197 source.n20 source.n18 0.716017
R198 source.n18 source.n16 0.716017
R199 source.n16 source.n14 0.716017
R200 source.n14 source.n12 0.716017
R201 source.n11 source.n10 0.716017
R202 source.n10 source.n8 0.716017
R203 source.n8 source.n6 0.716017
R204 source.n6 source.n4 0.716017
R205 source.n4 source.n2 0.716017
R206 source.n2 source.n0 0.716017
R207 source.n26 source.n24 0.716017
R208 source.n28 source.n26 0.716017
R209 source.n30 source.n28 0.716017
R210 source.n32 source.n30 0.716017
R211 source.n34 source.n32 0.716017
R212 source.n35 source.n34 0.716017
R213 source.n38 source.n36 0.716017
R214 source.n40 source.n38 0.716017
R215 source.n42 source.n40 0.716017
R216 source.n44 source.n42 0.716017
R217 source.n46 source.n44 0.716017
R218 source.n47 source.n46 0.716017
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 60.534
R223 drain_left.n7 drain_left.n5 60.5339
R224 drain_left.n2 drain_left.n0 60.5339
R225 drain_left.n21 drain_left.n20 59.8185
R226 drain_left.n19 drain_left.n18 59.8185
R227 drain_left.n17 drain_left.n16 59.8185
R228 drain_left.n15 drain_left.n14 59.8185
R229 drain_left.n13 drain_left.n12 59.8185
R230 drain_left.n7 drain_left.n6 59.8184
R231 drain_left.n9 drain_left.n8 59.8184
R232 drain_left.n4 drain_left.n3 59.8184
R233 drain_left.n2 drain_left.n1 59.8184
R234 drain_left drain_left.n10 40.2251
R235 drain_left drain_left.n21 6.36873
R236 drain_left.n5 drain_left.t22 0.9905
R237 drain_left.n5 drain_left.t23 0.9905
R238 drain_left.n6 drain_left.t17 0.9905
R239 drain_left.n6 drain_left.t11 0.9905
R240 drain_left.n8 drain_left.t7 0.9905
R241 drain_left.n8 drain_left.t16 0.9905
R242 drain_left.n3 drain_left.t19 0.9905
R243 drain_left.n3 drain_left.t12 0.9905
R244 drain_left.n1 drain_left.t8 0.9905
R245 drain_left.n1 drain_left.t9 0.9905
R246 drain_left.n0 drain_left.t1 0.9905
R247 drain_left.n0 drain_left.t14 0.9905
R248 drain_left.n20 drain_left.t20 0.9905
R249 drain_left.n20 drain_left.t21 0.9905
R250 drain_left.n18 drain_left.t18 0.9905
R251 drain_left.n18 drain_left.t6 0.9905
R252 drain_left.n16 drain_left.t10 0.9905
R253 drain_left.n16 drain_left.t3 0.9905
R254 drain_left.n14 drain_left.t4 0.9905
R255 drain_left.n14 drain_left.t0 0.9905
R256 drain_left.n12 drain_left.t2 0.9905
R257 drain_left.n12 drain_left.t13 0.9905
R258 drain_left.n11 drain_left.t15 0.9905
R259 drain_left.n11 drain_left.t5 0.9905
R260 drain_left.n9 drain_left.n7 0.716017
R261 drain_left.n4 drain_left.n2 0.716017
R262 drain_left.n15 drain_left.n13 0.716017
R263 drain_left.n17 drain_left.n15 0.716017
R264 drain_left.n19 drain_left.n17 0.716017
R265 drain_left.n21 drain_left.n19 0.716017
R266 drain_left.n10 drain_left.n9 0.302913
R267 drain_left.n10 drain_left.n4 0.302913
R268 minus.n9 minus.t14 1068.92
R269 minus.n43 minus.t6 1068.92
R270 minus.n8 minus.t1 1042.57
R271 minus.n7 minus.t8 1042.57
R272 minus.n13 minus.t21 1042.57
R273 minus.n5 minus.t7 1042.57
R274 minus.n18 minus.t10 1042.57
R275 minus.n20 minus.t0 1042.57
R276 minus.n3 minus.t12 1042.57
R277 minus.n25 minus.t18 1042.57
R278 minus.n1 minus.t4 1042.57
R279 minus.n30 minus.t15 1042.57
R280 minus.n32 minus.t22 1042.57
R281 minus.n42 minus.t5 1042.57
R282 minus.n41 minus.t17 1042.57
R283 minus.n47 minus.t13 1042.57
R284 minus.n39 minus.t9 1042.57
R285 minus.n52 minus.t20 1042.57
R286 minus.n54 minus.t19 1042.57
R287 minus.n37 minus.t11 1042.57
R288 minus.n59 minus.t2 1042.57
R289 minus.n35 minus.t23 1042.57
R290 minus.n64 minus.t16 1042.57
R291 minus.n66 minus.t3 1042.57
R292 minus.n33 minus.n32 161.3
R293 minus.n31 minus.n0 161.3
R294 minus.n30 minus.n29 161.3
R295 minus.n28 minus.n1 161.3
R296 minus.n27 minus.n26 161.3
R297 minus.n25 minus.n2 161.3
R298 minus.n24 minus.n23 161.3
R299 minus.n22 minus.n3 161.3
R300 minus.n21 minus.n20 161.3
R301 minus.n19 minus.n4 161.3
R302 minus.n18 minus.n17 161.3
R303 minus.n16 minus.n5 161.3
R304 minus.n15 minus.n14 161.3
R305 minus.n13 minus.n6 161.3
R306 minus.n12 minus.n11 161.3
R307 minus.n10 minus.n7 161.3
R308 minus.n67 minus.n66 161.3
R309 minus.n65 minus.n34 161.3
R310 minus.n64 minus.n63 161.3
R311 minus.n62 minus.n35 161.3
R312 minus.n61 minus.n60 161.3
R313 minus.n59 minus.n36 161.3
R314 minus.n58 minus.n57 161.3
R315 minus.n56 minus.n37 161.3
R316 minus.n55 minus.n54 161.3
R317 minus.n53 minus.n38 161.3
R318 minus.n52 minus.n51 161.3
R319 minus.n50 minus.n39 161.3
R320 minus.n49 minus.n48 161.3
R321 minus.n47 minus.n40 161.3
R322 minus.n46 minus.n45 161.3
R323 minus.n44 minus.n41 161.3
R324 minus.n8 minus.n7 48.2005
R325 minus.n18 minus.n5 48.2005
R326 minus.n20 minus.n3 48.2005
R327 minus.n30 minus.n1 48.2005
R328 minus.n42 minus.n41 48.2005
R329 minus.n52 minus.n39 48.2005
R330 minus.n54 minus.n37 48.2005
R331 minus.n64 minus.n35 48.2005
R332 minus.n14 minus.n13 47.4702
R333 minus.n25 minus.n24 47.4702
R334 minus.n48 minus.n47 47.4702
R335 minus.n59 minus.n58 47.4702
R336 minus.n68 minus.n33 46.0952
R337 minus.n32 minus.n31 46.0096
R338 minus.n66 minus.n65 46.0096
R339 minus.n10 minus.n9 45.0871
R340 minus.n44 minus.n43 45.0871
R341 minus.n13 minus.n12 25.5611
R342 minus.n26 minus.n25 25.5611
R343 minus.n47 minus.n46 25.5611
R344 minus.n60 minus.n59 25.5611
R345 minus.n20 minus.n19 24.1005
R346 minus.n19 minus.n18 24.1005
R347 minus.n53 minus.n52 24.1005
R348 minus.n54 minus.n53 24.1005
R349 minus.n12 minus.n7 22.6399
R350 minus.n26 minus.n1 22.6399
R351 minus.n46 minus.n41 22.6399
R352 minus.n60 minus.n35 22.6399
R353 minus.n9 minus.n8 14.1472
R354 minus.n43 minus.n42 14.1472
R355 minus.n68 minus.n67 6.52702
R356 minus.n31 minus.n30 2.19141
R357 minus.n65 minus.n64 2.19141
R358 minus.n14 minus.n5 0.730803
R359 minus.n24 minus.n3 0.730803
R360 minus.n48 minus.n39 0.730803
R361 minus.n58 minus.n37 0.730803
R362 minus.n33 minus.n0 0.189894
R363 minus.n29 minus.n0 0.189894
R364 minus.n29 minus.n28 0.189894
R365 minus.n28 minus.n27 0.189894
R366 minus.n27 minus.n2 0.189894
R367 minus.n23 minus.n2 0.189894
R368 minus.n23 minus.n22 0.189894
R369 minus.n22 minus.n21 0.189894
R370 minus.n21 minus.n4 0.189894
R371 minus.n17 minus.n4 0.189894
R372 minus.n17 minus.n16 0.189894
R373 minus.n16 minus.n15 0.189894
R374 minus.n15 minus.n6 0.189894
R375 minus.n11 minus.n6 0.189894
R376 minus.n11 minus.n10 0.189894
R377 minus.n45 minus.n44 0.189894
R378 minus.n45 minus.n40 0.189894
R379 minus.n49 minus.n40 0.189894
R380 minus.n50 minus.n49 0.189894
R381 minus.n51 minus.n50 0.189894
R382 minus.n51 minus.n38 0.189894
R383 minus.n55 minus.n38 0.189894
R384 minus.n56 minus.n55 0.189894
R385 minus.n57 minus.n56 0.189894
R386 minus.n57 minus.n36 0.189894
R387 minus.n61 minus.n36 0.189894
R388 minus.n62 minus.n61 0.189894
R389 minus.n63 minus.n62 0.189894
R390 minus.n63 minus.n34 0.189894
R391 minus.n67 minus.n34 0.189894
R392 minus minus.n68 0.188
R393 drain_right.n13 drain_right.n11 60.534
R394 drain_right.n7 drain_right.n5 60.5339
R395 drain_right.n2 drain_right.n0 60.5339
R396 drain_right.n13 drain_right.n12 59.8185
R397 drain_right.n15 drain_right.n14 59.8185
R398 drain_right.n17 drain_right.n16 59.8185
R399 drain_right.n19 drain_right.n18 59.8185
R400 drain_right.n21 drain_right.n20 59.8185
R401 drain_right.n7 drain_right.n6 59.8184
R402 drain_right.n9 drain_right.n8 59.8184
R403 drain_right.n4 drain_right.n3 59.8184
R404 drain_right.n2 drain_right.n1 59.8184
R405 drain_right drain_right.n10 39.6719
R406 drain_right drain_right.n21 6.36873
R407 drain_right.n5 drain_right.t7 0.9905
R408 drain_right.n5 drain_right.t20 0.9905
R409 drain_right.n6 drain_right.t21 0.9905
R410 drain_right.n6 drain_right.t0 0.9905
R411 drain_right.n8 drain_right.t4 0.9905
R412 drain_right.n8 drain_right.t12 0.9905
R413 drain_right.n3 drain_right.t14 0.9905
R414 drain_right.n3 drain_right.t3 0.9905
R415 drain_right.n1 drain_right.t6 0.9905
R416 drain_right.n1 drain_right.t10 0.9905
R417 drain_right.n0 drain_right.t17 0.9905
R418 drain_right.n0 drain_right.t18 0.9905
R419 drain_right.n11 drain_right.t22 0.9905
R420 drain_right.n11 drain_right.t9 0.9905
R421 drain_right.n12 drain_right.t2 0.9905
R422 drain_right.n12 drain_right.t15 0.9905
R423 drain_right.n14 drain_right.t13 0.9905
R424 drain_right.n14 drain_right.t16 0.9905
R425 drain_right.n16 drain_right.t11 0.9905
R426 drain_right.n16 drain_right.t23 0.9905
R427 drain_right.n18 drain_right.t19 0.9905
R428 drain_right.n18 drain_right.t5 0.9905
R429 drain_right.n20 drain_right.t1 0.9905
R430 drain_right.n20 drain_right.t8 0.9905
R431 drain_right.n9 drain_right.n7 0.716017
R432 drain_right.n4 drain_right.n2 0.716017
R433 drain_right.n21 drain_right.n19 0.716017
R434 drain_right.n19 drain_right.n17 0.716017
R435 drain_right.n17 drain_right.n15 0.716017
R436 drain_right.n15 drain_right.n13 0.716017
R437 drain_right.n10 drain_right.n9 0.302913
R438 drain_right.n10 drain_right.n4 0.302913
C0 minus source 19.4783f
C1 source drain_left 53.7813f
C2 plus drain_right 0.443411f
C3 plus minus 8.223009f
C4 minus drain_right 19.734098f
C5 plus drain_left 20.0205f
C6 plus source 19.4924f
C7 drain_left drain_right 1.55979f
C8 source drain_right 53.782898f
C9 minus drain_left 0.173624f
C10 drain_right a_n2874_n4888# 9.03784f
C11 drain_left a_n2874_n4888# 9.4458f
C12 source a_n2874_n4888# 13.652222f
C13 minus a_n2874_n4888# 12.059871f
C14 plus a_n2874_n4888# 14.46159f
C15 drain_right.t17 a_n2874_n4888# 0.465898f
C16 drain_right.t18 a_n2874_n4888# 0.465898f
C17 drain_right.n0 a_n2874_n4888# 4.26403f
C18 drain_right.t6 a_n2874_n4888# 0.465898f
C19 drain_right.t10 a_n2874_n4888# 0.465898f
C20 drain_right.n1 a_n2874_n4888# 4.25934f
C21 drain_right.n2 a_n2874_n4888# 0.77656f
C22 drain_right.t14 a_n2874_n4888# 0.465898f
C23 drain_right.t3 a_n2874_n4888# 0.465898f
C24 drain_right.n3 a_n2874_n4888# 4.25934f
C25 drain_right.n4 a_n2874_n4888# 0.347707f
C26 drain_right.t7 a_n2874_n4888# 0.465898f
C27 drain_right.t20 a_n2874_n4888# 0.465898f
C28 drain_right.n5 a_n2874_n4888# 4.26403f
C29 drain_right.t21 a_n2874_n4888# 0.465898f
C30 drain_right.t0 a_n2874_n4888# 0.465898f
C31 drain_right.n6 a_n2874_n4888# 4.25934f
C32 drain_right.n7 a_n2874_n4888# 0.77656f
C33 drain_right.t4 a_n2874_n4888# 0.465898f
C34 drain_right.t12 a_n2874_n4888# 0.465898f
C35 drain_right.n8 a_n2874_n4888# 4.25934f
C36 drain_right.n9 a_n2874_n4888# 0.347707f
C37 drain_right.n10 a_n2874_n4888# 2.29134f
C38 drain_right.t22 a_n2874_n4888# 0.465898f
C39 drain_right.t9 a_n2874_n4888# 0.465898f
C40 drain_right.n11 a_n2874_n4888# 4.26403f
C41 drain_right.t2 a_n2874_n4888# 0.465898f
C42 drain_right.t15 a_n2874_n4888# 0.465898f
C43 drain_right.n12 a_n2874_n4888# 4.25934f
C44 drain_right.n13 a_n2874_n4888# 0.776572f
C45 drain_right.t13 a_n2874_n4888# 0.465898f
C46 drain_right.t16 a_n2874_n4888# 0.465898f
C47 drain_right.n14 a_n2874_n4888# 4.25934f
C48 drain_right.n15 a_n2874_n4888# 0.384693f
C49 drain_right.t11 a_n2874_n4888# 0.465898f
C50 drain_right.t23 a_n2874_n4888# 0.465898f
C51 drain_right.n16 a_n2874_n4888# 4.25934f
C52 drain_right.n17 a_n2874_n4888# 0.384693f
C53 drain_right.t19 a_n2874_n4888# 0.465898f
C54 drain_right.t5 a_n2874_n4888# 0.465898f
C55 drain_right.n18 a_n2874_n4888# 4.25934f
C56 drain_right.n19 a_n2874_n4888# 0.384693f
C57 drain_right.t1 a_n2874_n4888# 0.465898f
C58 drain_right.t8 a_n2874_n4888# 0.465898f
C59 drain_right.n20 a_n2874_n4888# 4.25934f
C60 drain_right.n21 a_n2874_n4888# 0.637955f
C61 minus.n0 a_n2874_n4888# 0.043355f
C62 minus.t4 a_n2874_n4888# 1.22775f
C63 minus.n1 a_n2874_n4888# 0.465352f
C64 minus.t15 a_n2874_n4888# 1.22775f
C65 minus.n2 a_n2874_n4888# 0.043355f
C66 minus.t12 a_n2874_n4888# 1.22775f
C67 minus.n3 a_n2874_n4888# 0.461343f
C68 minus.n4 a_n2874_n4888# 0.043355f
C69 minus.t7 a_n2874_n4888# 1.22775f
C70 minus.n5 a_n2874_n4888# 0.461343f
C71 minus.t10 a_n2874_n4888# 1.22775f
C72 minus.n6 a_n2874_n4888# 0.043355f
C73 minus.t8 a_n2874_n4888# 1.22775f
C74 minus.n7 a_n2874_n4888# 0.465352f
C75 minus.t14 a_n2874_n4888# 1.23913f
C76 minus.t1 a_n2874_n4888# 1.22775f
C77 minus.n8 a_n2874_n4888# 0.470482f
C78 minus.n9 a_n2874_n4888# 0.451258f
C79 minus.n10 a_n2874_n4888# 0.176037f
C80 minus.n11 a_n2874_n4888# 0.043355f
C81 minus.n12 a_n2874_n4888# 0.009838f
C82 minus.t21 a_n2874_n4888# 1.22775f
C83 minus.n13 a_n2874_n4888# 0.465753f
C84 minus.n14 a_n2874_n4888# 0.009838f
C85 minus.n15 a_n2874_n4888# 0.043355f
C86 minus.n16 a_n2874_n4888# 0.043355f
C87 minus.n17 a_n2874_n4888# 0.043355f
C88 minus.n18 a_n2874_n4888# 0.46562f
C89 minus.n19 a_n2874_n4888# 0.009838f
C90 minus.t0 a_n2874_n4888# 1.22775f
C91 minus.n20 a_n2874_n4888# 0.46562f
C92 minus.n21 a_n2874_n4888# 0.043355f
C93 minus.n22 a_n2874_n4888# 0.043355f
C94 minus.n23 a_n2874_n4888# 0.043355f
C95 minus.n24 a_n2874_n4888# 0.009838f
C96 minus.t18 a_n2874_n4888# 1.22775f
C97 minus.n25 a_n2874_n4888# 0.465753f
C98 minus.n26 a_n2874_n4888# 0.009838f
C99 minus.n27 a_n2874_n4888# 0.043355f
C100 minus.n28 a_n2874_n4888# 0.043355f
C101 minus.n29 a_n2874_n4888# 0.043355f
C102 minus.n30 a_n2874_n4888# 0.46161f
C103 minus.n31 a_n2874_n4888# 0.009838f
C104 minus.t22 a_n2874_n4888# 1.22775f
C105 minus.n32 a_n2874_n4888# 0.460808f
C106 minus.n33 a_n2874_n4888# 2.19758f
C107 minus.n34 a_n2874_n4888# 0.043355f
C108 minus.t23 a_n2874_n4888# 1.22775f
C109 minus.n35 a_n2874_n4888# 0.465352f
C110 minus.n36 a_n2874_n4888# 0.043355f
C111 minus.t11 a_n2874_n4888# 1.22775f
C112 minus.n37 a_n2874_n4888# 0.461343f
C113 minus.n38 a_n2874_n4888# 0.043355f
C114 minus.t9 a_n2874_n4888# 1.22775f
C115 minus.n39 a_n2874_n4888# 0.461343f
C116 minus.n40 a_n2874_n4888# 0.043355f
C117 minus.t17 a_n2874_n4888# 1.22775f
C118 minus.n41 a_n2874_n4888# 0.465352f
C119 minus.t6 a_n2874_n4888# 1.23913f
C120 minus.t5 a_n2874_n4888# 1.22775f
C121 minus.n42 a_n2874_n4888# 0.470482f
C122 minus.n43 a_n2874_n4888# 0.451258f
C123 minus.n44 a_n2874_n4888# 0.176037f
C124 minus.n45 a_n2874_n4888# 0.043355f
C125 minus.n46 a_n2874_n4888# 0.009838f
C126 minus.t13 a_n2874_n4888# 1.22775f
C127 minus.n47 a_n2874_n4888# 0.465753f
C128 minus.n48 a_n2874_n4888# 0.009838f
C129 minus.n49 a_n2874_n4888# 0.043355f
C130 minus.n50 a_n2874_n4888# 0.043355f
C131 minus.n51 a_n2874_n4888# 0.043355f
C132 minus.t20 a_n2874_n4888# 1.22775f
C133 minus.n52 a_n2874_n4888# 0.46562f
C134 minus.n53 a_n2874_n4888# 0.009838f
C135 minus.t19 a_n2874_n4888# 1.22775f
C136 minus.n54 a_n2874_n4888# 0.46562f
C137 minus.n55 a_n2874_n4888# 0.043355f
C138 minus.n56 a_n2874_n4888# 0.043355f
C139 minus.n57 a_n2874_n4888# 0.043355f
C140 minus.n58 a_n2874_n4888# 0.009838f
C141 minus.t2 a_n2874_n4888# 1.22775f
C142 minus.n59 a_n2874_n4888# 0.465753f
C143 minus.n60 a_n2874_n4888# 0.009838f
C144 minus.n61 a_n2874_n4888# 0.043355f
C145 minus.n62 a_n2874_n4888# 0.043355f
C146 minus.n63 a_n2874_n4888# 0.043355f
C147 minus.t16 a_n2874_n4888# 1.22775f
C148 minus.n64 a_n2874_n4888# 0.46161f
C149 minus.n65 a_n2874_n4888# 0.009838f
C150 minus.t3 a_n2874_n4888# 1.22775f
C151 minus.n66 a_n2874_n4888# 0.460808f
C152 minus.n67 a_n2874_n4888# 0.286196f
C153 minus.n68 a_n2874_n4888# 2.59428f
C154 drain_left.t1 a_n2874_n4888# 0.467067f
C155 drain_left.t14 a_n2874_n4888# 0.467067f
C156 drain_left.n0 a_n2874_n4888# 4.27473f
C157 drain_left.t8 a_n2874_n4888# 0.467067f
C158 drain_left.t9 a_n2874_n4888# 0.467067f
C159 drain_left.n1 a_n2874_n4888# 4.27003f
C160 drain_left.n2 a_n2874_n4888# 0.778508f
C161 drain_left.t19 a_n2874_n4888# 0.467067f
C162 drain_left.t12 a_n2874_n4888# 0.467067f
C163 drain_left.n3 a_n2874_n4888# 4.27003f
C164 drain_left.n4 a_n2874_n4888# 0.348579f
C165 drain_left.t22 a_n2874_n4888# 0.467067f
C166 drain_left.t23 a_n2874_n4888# 0.467067f
C167 drain_left.n5 a_n2874_n4888# 4.27473f
C168 drain_left.t17 a_n2874_n4888# 0.467067f
C169 drain_left.t11 a_n2874_n4888# 0.467067f
C170 drain_left.n6 a_n2874_n4888# 4.27003f
C171 drain_left.n7 a_n2874_n4888# 0.778508f
C172 drain_left.t7 a_n2874_n4888# 0.467067f
C173 drain_left.t16 a_n2874_n4888# 0.467067f
C174 drain_left.n8 a_n2874_n4888# 4.27003f
C175 drain_left.n9 a_n2874_n4888# 0.348579f
C176 drain_left.n10 a_n2874_n4888# 2.35772f
C177 drain_left.t15 a_n2874_n4888# 0.467067f
C178 drain_left.t5 a_n2874_n4888# 0.467067f
C179 drain_left.n11 a_n2874_n4888# 4.27472f
C180 drain_left.t2 a_n2874_n4888# 0.467067f
C181 drain_left.t13 a_n2874_n4888# 0.467067f
C182 drain_left.n12 a_n2874_n4888# 4.27002f
C183 drain_left.n13 a_n2874_n4888# 0.77852f
C184 drain_left.t4 a_n2874_n4888# 0.467067f
C185 drain_left.t0 a_n2874_n4888# 0.467067f
C186 drain_left.n14 a_n2874_n4888# 4.27002f
C187 drain_left.n15 a_n2874_n4888# 0.385658f
C188 drain_left.t10 a_n2874_n4888# 0.467067f
C189 drain_left.t3 a_n2874_n4888# 0.467067f
C190 drain_left.n16 a_n2874_n4888# 4.27002f
C191 drain_left.n17 a_n2874_n4888# 0.385658f
C192 drain_left.t18 a_n2874_n4888# 0.467067f
C193 drain_left.t6 a_n2874_n4888# 0.467067f
C194 drain_left.n18 a_n2874_n4888# 4.27002f
C195 drain_left.n19 a_n2874_n4888# 0.385658f
C196 drain_left.t20 a_n2874_n4888# 0.467067f
C197 drain_left.t21 a_n2874_n4888# 0.467067f
C198 drain_left.n20 a_n2874_n4888# 4.27002f
C199 drain_left.n21 a_n2874_n4888# 0.639556f
C200 source.t40 a_n2874_n4888# 4.68055f
C201 source.n0 a_n2874_n4888# 2.01349f
C202 source.t43 a_n2874_n4888# 0.409555f
C203 source.t39 a_n2874_n4888# 0.409555f
C204 source.n1 a_n2874_n4888# 3.6616f
C205 source.n2 a_n2874_n4888# 0.385588f
C206 source.t36 a_n2874_n4888# 0.409555f
C207 source.t23 a_n2874_n4888# 0.409555f
C208 source.n3 a_n2874_n4888# 3.6616f
C209 source.n4 a_n2874_n4888# 0.385588f
C210 source.t33 a_n2874_n4888# 0.409555f
C211 source.t26 a_n2874_n4888# 0.409555f
C212 source.n5 a_n2874_n4888# 3.6616f
C213 source.n6 a_n2874_n4888# 0.385588f
C214 source.t41 a_n2874_n4888# 0.409555f
C215 source.t24 a_n2874_n4888# 0.409555f
C216 source.n7 a_n2874_n4888# 3.6616f
C217 source.n8 a_n2874_n4888# 0.385588f
C218 source.t45 a_n2874_n4888# 0.409555f
C219 source.t35 a_n2874_n4888# 0.409555f
C220 source.n9 a_n2874_n4888# 3.6616f
C221 source.n10 a_n2874_n4888# 0.385588f
C222 source.t31 a_n2874_n4888# 4.68056f
C223 source.n11 a_n2874_n4888# 0.463078f
C224 source.t18 a_n2874_n4888# 4.68056f
C225 source.n12 a_n2874_n4888# 0.463078f
C226 source.t20 a_n2874_n4888# 0.409555f
C227 source.t14 a_n2874_n4888# 0.409555f
C228 source.n13 a_n2874_n4888# 3.6616f
C229 source.n14 a_n2874_n4888# 0.385588f
C230 source.t21 a_n2874_n4888# 0.409555f
C231 source.t0 a_n2874_n4888# 0.409555f
C232 source.n15 a_n2874_n4888# 3.6616f
C233 source.n16 a_n2874_n4888# 0.385588f
C234 source.t17 a_n2874_n4888# 0.409555f
C235 source.t9 a_n2874_n4888# 0.409555f
C236 source.n17 a_n2874_n4888# 3.6616f
C237 source.n18 a_n2874_n4888# 0.385588f
C238 source.t6 a_n2874_n4888# 0.409555f
C239 source.t47 a_n2874_n4888# 0.409555f
C240 source.n19 a_n2874_n4888# 3.6616f
C241 source.n20 a_n2874_n4888# 0.385588f
C242 source.t1 a_n2874_n4888# 0.409555f
C243 source.t8 a_n2874_n4888# 0.409555f
C244 source.n21 a_n2874_n4888# 3.6616f
C245 source.n22 a_n2874_n4888# 0.385588f
C246 source.t2 a_n2874_n4888# 4.68056f
C247 source.n23 a_n2874_n4888# 2.47881f
C248 source.t34 a_n2874_n4888# 4.68053f
C249 source.n24 a_n2874_n4888# 2.47883f
C250 source.t30 a_n2874_n4888# 0.409555f
C251 source.t42 a_n2874_n4888# 0.409555f
C252 source.n25 a_n2874_n4888# 3.6616f
C253 source.n26 a_n2874_n4888# 0.385581f
C254 source.t25 a_n2874_n4888# 0.409555f
C255 source.t38 a_n2874_n4888# 0.409555f
C256 source.n27 a_n2874_n4888# 3.6616f
C257 source.n28 a_n2874_n4888# 0.385581f
C258 source.t27 a_n2874_n4888# 0.409555f
C259 source.t44 a_n2874_n4888# 0.409555f
C260 source.n29 a_n2874_n4888# 3.6616f
C261 source.n30 a_n2874_n4888# 0.385581f
C262 source.t32 a_n2874_n4888# 0.409555f
C263 source.t37 a_n2874_n4888# 0.409555f
C264 source.n31 a_n2874_n4888# 3.6616f
C265 source.n32 a_n2874_n4888# 0.385581f
C266 source.t22 a_n2874_n4888# 0.409555f
C267 source.t28 a_n2874_n4888# 0.409555f
C268 source.n33 a_n2874_n4888# 3.6616f
C269 source.n34 a_n2874_n4888# 0.385581f
C270 source.t29 a_n2874_n4888# 4.68053f
C271 source.n35 a_n2874_n4888# 0.463104f
C272 source.t7 a_n2874_n4888# 4.68053f
C273 source.n36 a_n2874_n4888# 0.463104f
C274 source.t4 a_n2874_n4888# 0.409555f
C275 source.t16 a_n2874_n4888# 0.409555f
C276 source.n37 a_n2874_n4888# 3.6616f
C277 source.n38 a_n2874_n4888# 0.385581f
C278 source.t5 a_n2874_n4888# 0.409555f
C279 source.t10 a_n2874_n4888# 0.409555f
C280 source.n39 a_n2874_n4888# 3.6616f
C281 source.n40 a_n2874_n4888# 0.385581f
C282 source.t15 a_n2874_n4888# 0.409555f
C283 source.t11 a_n2874_n4888# 0.409555f
C284 source.n41 a_n2874_n4888# 3.6616f
C285 source.n42 a_n2874_n4888# 0.385581f
C286 source.t46 a_n2874_n4888# 0.409555f
C287 source.t19 a_n2874_n4888# 0.409555f
C288 source.n43 a_n2874_n4888# 3.6616f
C289 source.n44 a_n2874_n4888# 0.385581f
C290 source.t13 a_n2874_n4888# 0.409555f
C291 source.t12 a_n2874_n4888# 0.409555f
C292 source.n45 a_n2874_n4888# 3.6616f
C293 source.n46 a_n2874_n4888# 0.385581f
C294 source.t3 a_n2874_n4888# 4.68053f
C295 source.n47 a_n2874_n4888# 0.620827f
C296 source.n48 a_n2874_n4888# 2.34177f
C297 plus.n0 a_n2874_n4888# 0.04371f
C298 plus.t2 a_n2874_n4888# 1.23781f
C299 plus.t3 a_n2874_n4888# 1.23781f
C300 plus.n1 a_n2874_n4888# 0.04371f
C301 plus.t17 a_n2874_n4888# 1.23781f
C302 plus.n2 a_n2874_n4888# 0.04371f
C303 plus.t5 a_n2874_n4888# 1.23781f
C304 plus.n3 a_n2874_n4888# 0.46957f
C305 plus.n4 a_n2874_n4888# 0.04371f
C306 plus.t20 a_n2874_n4888# 1.23781f
C307 plus.t13 a_n2874_n4888# 1.23781f
C308 plus.n5 a_n2874_n4888# 0.04371f
C309 plus.t23 a_n2874_n4888# 1.23781f
C310 plus.n6 a_n2874_n4888# 0.469435f
C311 plus.n7 a_n2874_n4888# 0.04371f
C312 plus.t19 a_n2874_n4888# 1.23781f
C313 plus.t10 a_n2874_n4888# 1.23781f
C314 plus.n8 a_n2874_n4888# 0.04371f
C315 plus.t21 a_n2874_n4888# 1.23781f
C316 plus.n9 a_n2874_n4888# 0.469165f
C317 plus.t18 a_n2874_n4888# 1.23781f
C318 plus.n10 a_n2874_n4888# 0.474337f
C319 plus.t8 a_n2874_n4888# 1.24928f
C320 plus.n11 a_n2874_n4888# 0.454956f
C321 plus.n12 a_n2874_n4888# 0.17748f
C322 plus.n13 a_n2874_n4888# 0.04371f
C323 plus.n14 a_n2874_n4888# 0.009919f
C324 plus.n15 a_n2874_n4888# 0.46957f
C325 plus.n16 a_n2874_n4888# 0.009919f
C326 plus.n17 a_n2874_n4888# 0.465123f
C327 plus.n18 a_n2874_n4888# 0.04371f
C328 plus.n19 a_n2874_n4888# 0.04371f
C329 plus.n20 a_n2874_n4888# 0.04371f
C330 plus.n21 a_n2874_n4888# 0.009919f
C331 plus.n22 a_n2874_n4888# 0.469435f
C332 plus.n23 a_n2874_n4888# 0.465123f
C333 plus.n24 a_n2874_n4888# 0.009919f
C334 plus.n25 a_n2874_n4888# 0.04371f
C335 plus.n26 a_n2874_n4888# 0.04371f
C336 plus.n27 a_n2874_n4888# 0.04371f
C337 plus.n28 a_n2874_n4888# 0.009919f
C338 plus.n29 a_n2874_n4888# 0.469165f
C339 plus.n30 a_n2874_n4888# 0.465392f
C340 plus.n31 a_n2874_n4888# 0.009919f
C341 plus.n32 a_n2874_n4888# 0.464584f
C342 plus.n33 a_n2874_n4888# 0.666418f
C343 plus.n34 a_n2874_n4888# 0.04371f
C344 plus.t22 a_n2874_n4888# 1.23781f
C345 plus.n35 a_n2874_n4888# 0.04371f
C346 plus.t9 a_n2874_n4888# 1.23781f
C347 plus.n36 a_n2874_n4888# 0.04371f
C348 plus.t15 a_n2874_n4888# 1.23781f
C349 plus.t14 a_n2874_n4888# 1.23781f
C350 plus.n37 a_n2874_n4888# 0.46957f
C351 plus.n38 a_n2874_n4888# 0.04371f
C352 plus.t4 a_n2874_n4888# 1.23781f
C353 plus.n39 a_n2874_n4888# 0.04371f
C354 plus.t11 a_n2874_n4888# 1.23781f
C355 plus.t16 a_n2874_n4888# 1.23781f
C356 plus.n40 a_n2874_n4888# 0.469435f
C357 plus.n41 a_n2874_n4888# 0.04371f
C358 plus.t7 a_n2874_n4888# 1.23781f
C359 plus.n42 a_n2874_n4888# 0.04371f
C360 plus.t6 a_n2874_n4888# 1.23781f
C361 plus.t12 a_n2874_n4888# 1.23781f
C362 plus.n43 a_n2874_n4888# 0.469165f
C363 plus.t0 a_n2874_n4888# 1.24928f
C364 plus.t1 a_n2874_n4888# 1.23781f
C365 plus.n44 a_n2874_n4888# 0.474337f
C366 plus.n45 a_n2874_n4888# 0.454956f
C367 plus.n46 a_n2874_n4888# 0.17748f
C368 plus.n47 a_n2874_n4888# 0.04371f
C369 plus.n48 a_n2874_n4888# 0.009919f
C370 plus.n49 a_n2874_n4888# 0.46957f
C371 plus.n50 a_n2874_n4888# 0.009919f
C372 plus.n51 a_n2874_n4888# 0.465123f
C373 plus.n52 a_n2874_n4888# 0.04371f
C374 plus.n53 a_n2874_n4888# 0.04371f
C375 plus.n54 a_n2874_n4888# 0.04371f
C376 plus.n55 a_n2874_n4888# 0.009919f
C377 plus.n56 a_n2874_n4888# 0.469435f
C378 plus.n57 a_n2874_n4888# 0.465123f
C379 plus.n58 a_n2874_n4888# 0.009919f
C380 plus.n59 a_n2874_n4888# 0.04371f
C381 plus.n60 a_n2874_n4888# 0.04371f
C382 plus.n61 a_n2874_n4888# 0.04371f
C383 plus.n62 a_n2874_n4888# 0.009919f
C384 plus.n63 a_n2874_n4888# 0.469165f
C385 plus.n64 a_n2874_n4888# 0.465392f
C386 plus.n65 a_n2874_n4888# 0.009919f
C387 plus.n66 a_n2874_n4888# 0.464584f
C388 plus.n67 a_n2874_n4888# 1.77986f
.ends

