* NGSPICE file created from diffpair495.ext - technology: sky130A

.subckt diffpair495 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t19 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t10 plus.t1 source.t20 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X2 drain_left.t9 plus.t2 source.t23 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X3 drain_right.t11 minus.t0 source.t1 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X4 source.t13 plus.t3 drain_left.t8 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 drain_left.t7 plus.t4 source.t15 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 source.t7 minus.t1 drain_right.t10 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X7 source.t9 minus.t2 drain_right.t9 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 source.t5 minus.t3 drain_right.t8 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 source.t6 minus.t4 drain_right.t7 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X10 drain_left.t6 plus.t5 source.t17 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X11 source.t22 plus.t6 drain_left.t5 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X12 drain_right.t6 minus.t5 source.t10 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X13 drain_right.t5 minus.t6 source.t4 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X14 a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X15 drain_right.t4 minus.t7 source.t8 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X16 drain_right.t3 minus.t8 source.t11 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X17 drain_right.t2 minus.t9 source.t0 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X18 a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X19 source.t2 minus.t10 drain_right.t1 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X20 a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X21 source.t14 plus.t7 drain_left.t4 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X22 drain_left.t3 plus.t8 source.t16 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X23 source.t3 minus.t11 drain_right.t0 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X24 source.t12 plus.t9 drain_left.t2 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X25 source.t21 plus.t10 drain_left.t1 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X26 a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X27 source.t18 plus.t11 drain_left.t0 a_n1458_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n2 plus.t6 2011.62
R1 plus.n11 plus.t5 2011.62
R2 plus.n15 plus.t2 2011.62
R3 plus.n24 plus.t10 2011.62
R4 plus.n3 plus.t4 1964.15
R5 plus.n1 plus.t11 1964.15
R6 plus.n8 plus.t8 1964.15
R7 plus.n10 plus.t7 1964.15
R8 plus.n16 plus.t3 1964.15
R9 plus.n14 plus.t1 1964.15
R10 plus.n21 plus.t9 1964.15
R11 plus.n23 plus.t0 1964.15
R12 plus.n5 plus.n2 161.489
R13 plus.n18 plus.n15 161.489
R14 plus.n5 plus.n4 161.3
R15 plus.n7 plus.n6 161.3
R16 plus.n9 plus.n0 161.3
R17 plus.n12 plus.n11 161.3
R18 plus.n18 plus.n17 161.3
R19 plus.n20 plus.n19 161.3
R20 plus.n22 plus.n13 161.3
R21 plus.n25 plus.n24 161.3
R22 plus.n4 plus.n3 43.0884
R23 plus.n10 plus.n9 43.0884
R24 plus.n23 plus.n22 43.0884
R25 plus.n17 plus.n16 43.0884
R26 plus.n7 plus.n1 38.7066
R27 plus.n8 plus.n7 38.7066
R28 plus.n21 plus.n20 38.7066
R29 plus.n20 plus.n14 38.7066
R30 plus.n4 plus.n1 34.3247
R31 plus.n9 plus.n8 34.3247
R32 plus.n22 plus.n21 34.3247
R33 plus.n17 plus.n14 34.3247
R34 plus.n3 plus.n2 29.9429
R35 plus.n11 plus.n10 29.9429
R36 plus.n24 plus.n23 29.9429
R37 plus.n16 plus.n15 29.9429
R38 plus plus.n25 29.6164
R39 plus plus.n12 13.2353
R40 plus.n6 plus.n5 0.189894
R41 plus.n6 plus.n0 0.189894
R42 plus.n12 plus.n0 0.189894
R43 plus.n25 plus.n13 0.189894
R44 plus.n19 plus.n13 0.189894
R45 plus.n19 plus.n18 0.189894
R46 source.n5 source.t22 45.521
R47 source.n6 source.t11 45.521
R48 source.n11 source.t7 45.521
R49 source.n23 source.t8 45.5208
R50 source.n18 source.t6 45.5208
R51 source.n17 source.t23 45.5208
R52 source.n12 source.t21 45.5208
R53 source.n0 source.t17 45.5208
R54 source.n2 source.n1 44.201
R55 source.n4 source.n3 44.201
R56 source.n8 source.n7 44.201
R57 source.n10 source.n9 44.201
R58 source.n22 source.n21 44.2008
R59 source.n20 source.n19 44.2008
R60 source.n16 source.n15 44.2008
R61 source.n14 source.n13 44.2008
R62 source.n12 source.n11 24.0173
R63 source.n24 source.n0 18.526
R64 source.n24 source.n23 5.49188
R65 source.n21 source.t10 1.3205
R66 source.n21 source.t2 1.3205
R67 source.n19 source.t4 1.3205
R68 source.n19 source.t9 1.3205
R69 source.n15 source.t20 1.3205
R70 source.n15 source.t13 1.3205
R71 source.n13 source.t19 1.3205
R72 source.n13 source.t12 1.3205
R73 source.n1 source.t16 1.3205
R74 source.n1 source.t14 1.3205
R75 source.n3 source.t15 1.3205
R76 source.n3 source.t18 1.3205
R77 source.n7 source.t1 1.3205
R78 source.n7 source.t5 1.3205
R79 source.n9 source.t0 1.3205
R80 source.n9 source.t3 1.3205
R81 source.n6 source.n5 0.470328
R82 source.n18 source.n17 0.470328
R83 source.n11 source.n10 0.457397
R84 source.n10 source.n8 0.457397
R85 source.n8 source.n6 0.457397
R86 source.n5 source.n4 0.457397
R87 source.n4 source.n2 0.457397
R88 source.n2 source.n0 0.457397
R89 source.n14 source.n12 0.457397
R90 source.n16 source.n14 0.457397
R91 source.n17 source.n16 0.457397
R92 source.n20 source.n18 0.457397
R93 source.n22 source.n20 0.457397
R94 source.n23 source.n22 0.457397
R95 source source.n24 0.188
R96 drain_left.n6 drain_left.n4 61.3367
R97 drain_left.n3 drain_left.n2 61.2811
R98 drain_left.n3 drain_left.n0 61.2811
R99 drain_left.n6 drain_left.n5 60.8798
R100 drain_left.n8 drain_left.n7 60.8796
R101 drain_left.n3 drain_left.n1 60.8796
R102 drain_left drain_left.n3 31.9243
R103 drain_left drain_left.n8 6.11011
R104 drain_left.n1 drain_left.t2 1.3205
R105 drain_left.n1 drain_left.t10 1.3205
R106 drain_left.n2 drain_left.t8 1.3205
R107 drain_left.n2 drain_left.t9 1.3205
R108 drain_left.n0 drain_left.t1 1.3205
R109 drain_left.n0 drain_left.t11 1.3205
R110 drain_left.n7 drain_left.t4 1.3205
R111 drain_left.n7 drain_left.t6 1.3205
R112 drain_left.n5 drain_left.t0 1.3205
R113 drain_left.n5 drain_left.t3 1.3205
R114 drain_left.n4 drain_left.t5 1.3205
R115 drain_left.n4 drain_left.t7 1.3205
R116 drain_left.n8 drain_left.n6 0.457397
R117 minus.n11 minus.t1 2011.62
R118 minus.n2 minus.t8 2011.62
R119 minus.n24 minus.t7 2011.62
R120 minus.n15 minus.t4 2011.62
R121 minus.n10 minus.t9 1964.15
R122 minus.n8 minus.t11 1964.15
R123 minus.n1 minus.t0 1964.15
R124 minus.n3 minus.t3 1964.15
R125 minus.n23 minus.t10 1964.15
R126 minus.n21 minus.t5 1964.15
R127 minus.n14 minus.t2 1964.15
R128 minus.n16 minus.t6 1964.15
R129 minus.n5 minus.n2 161.489
R130 minus.n18 minus.n15 161.489
R131 minus.n12 minus.n11 161.3
R132 minus.n9 minus.n0 161.3
R133 minus.n7 minus.n6 161.3
R134 minus.n5 minus.n4 161.3
R135 minus.n25 minus.n24 161.3
R136 minus.n22 minus.n13 161.3
R137 minus.n20 minus.n19 161.3
R138 minus.n18 minus.n17 161.3
R139 minus.n10 minus.n9 43.0884
R140 minus.n4 minus.n3 43.0884
R141 minus.n17 minus.n16 43.0884
R142 minus.n23 minus.n22 43.0884
R143 minus.n8 minus.n7 38.7066
R144 minus.n7 minus.n1 38.7066
R145 minus.n20 minus.n14 38.7066
R146 minus.n21 minus.n20 38.7066
R147 minus.n26 minus.n12 36.8717
R148 minus.n9 minus.n8 34.3247
R149 minus.n4 minus.n1 34.3247
R150 minus.n17 minus.n14 34.3247
R151 minus.n22 minus.n21 34.3247
R152 minus.n11 minus.n10 29.9429
R153 minus.n3 minus.n2 29.9429
R154 minus.n16 minus.n15 29.9429
R155 minus.n24 minus.n23 29.9429
R156 minus.n26 minus.n25 6.45505
R157 minus.n12 minus.n0 0.189894
R158 minus.n6 minus.n0 0.189894
R159 minus.n6 minus.n5 0.189894
R160 minus.n19 minus.n18 0.189894
R161 minus.n19 minus.n13 0.189894
R162 minus.n25 minus.n13 0.189894
R163 minus minus.n26 0.188
R164 drain_right.n6 drain_right.n4 61.3365
R165 drain_right.n3 drain_right.n2 61.2811
R166 drain_right.n3 drain_right.n0 61.2811
R167 drain_right.n6 drain_right.n5 60.8798
R168 drain_right.n8 drain_right.n7 60.8798
R169 drain_right.n3 drain_right.n1 60.8796
R170 drain_right drain_right.n3 31.3711
R171 drain_right drain_right.n8 6.11011
R172 drain_right.n1 drain_right.t9 1.3205
R173 drain_right.n1 drain_right.t6 1.3205
R174 drain_right.n2 drain_right.t1 1.3205
R175 drain_right.n2 drain_right.t4 1.3205
R176 drain_right.n0 drain_right.t7 1.3205
R177 drain_right.n0 drain_right.t5 1.3205
R178 drain_right.n4 drain_right.t8 1.3205
R179 drain_right.n4 drain_right.t3 1.3205
R180 drain_right.n5 drain_right.t0 1.3205
R181 drain_right.n5 drain_right.t11 1.3205
R182 drain_right.n7 drain_right.t10 1.3205
R183 drain_right.n7 drain_right.t2 1.3205
R184 drain_right.n8 drain_right.n6 0.457397
C0 plus minus 5.52833f
C1 plus drain_left 4.44241f
C2 drain_left minus 0.17046f
C3 source drain_right 34.6502f
C4 plus drain_right 0.292203f
C5 drain_right minus 4.30353f
C6 drain_left drain_right 0.711832f
C7 plus source 3.73288f
C8 source minus 3.71884f
C9 source drain_left 34.6511f
C10 drain_right a_n1458_n3888# 7.1143f
C11 drain_left a_n1458_n3888# 7.3525f
C12 source a_n1458_n3888# 10.065277f
C13 minus a_n1458_n3888# 5.835226f
C14 plus a_n1458_n3888# 8.11596f
C15 drain_right.t7 a_n1458_n3888# 0.455935f
C16 drain_right.t5 a_n1458_n3888# 0.455935f
C17 drain_right.n0 a_n1458_n3888# 4.123991f
C18 drain_right.t9 a_n1458_n3888# 0.455935f
C19 drain_right.t6 a_n1458_n3888# 0.455935f
C20 drain_right.n1 a_n1458_n3888# 4.12112f
C21 drain_right.t1 a_n1458_n3888# 0.455935f
C22 drain_right.t4 a_n1458_n3888# 0.455935f
C23 drain_right.n2 a_n1458_n3888# 4.123991f
C24 drain_right.n3 a_n1458_n3888# 3.162f
C25 drain_right.t8 a_n1458_n3888# 0.455935f
C26 drain_right.t3 a_n1458_n3888# 0.455935f
C27 drain_right.n4 a_n1458_n3888# 4.12441f
C28 drain_right.t0 a_n1458_n3888# 0.455935f
C29 drain_right.t11 a_n1458_n3888# 0.455935f
C30 drain_right.n5 a_n1458_n3888# 4.12112f
C31 drain_right.n6 a_n1458_n3888# 0.868798f
C32 drain_right.t10 a_n1458_n3888# 0.455935f
C33 drain_right.t2 a_n1458_n3888# 0.455935f
C34 drain_right.n7 a_n1458_n3888# 4.12112f
C35 drain_right.n8 a_n1458_n3888# 0.743092f
C36 minus.n0 a_n1458_n3888# 0.055941f
C37 minus.t1 a_n1458_n3888# 0.477901f
C38 minus.t9 a_n1458_n3888# 0.473454f
C39 minus.t11 a_n1458_n3888# 0.473454f
C40 minus.t0 a_n1458_n3888# 0.473454f
C41 minus.n1 a_n1458_n3888# 0.187605f
C42 minus.t8 a_n1458_n3888# 0.477901f
C43 minus.n2 a_n1458_n3888# 0.203692f
C44 minus.t3 a_n1458_n3888# 0.473454f
C45 minus.n3 a_n1458_n3888# 0.187605f
C46 minus.n4 a_n1458_n3888# 0.019592f
C47 minus.n5 a_n1458_n3888# 0.123874f
C48 minus.n6 a_n1458_n3888# 0.055941f
C49 minus.n7 a_n1458_n3888# 0.019592f
C50 minus.n8 a_n1458_n3888# 0.187605f
C51 minus.n9 a_n1458_n3888# 0.019592f
C52 minus.n10 a_n1458_n3888# 0.187605f
C53 minus.n11 a_n1458_n3888# 0.203612f
C54 minus.n12 a_n1458_n3888# 2.03308f
C55 minus.n13 a_n1458_n3888# 0.055941f
C56 minus.t10 a_n1458_n3888# 0.473454f
C57 minus.t5 a_n1458_n3888# 0.473454f
C58 minus.t2 a_n1458_n3888# 0.473454f
C59 minus.n14 a_n1458_n3888# 0.187605f
C60 minus.t4 a_n1458_n3888# 0.477901f
C61 minus.n15 a_n1458_n3888# 0.203692f
C62 minus.t6 a_n1458_n3888# 0.473454f
C63 minus.n16 a_n1458_n3888# 0.187605f
C64 minus.n17 a_n1458_n3888# 0.019592f
C65 minus.n18 a_n1458_n3888# 0.123874f
C66 minus.n19 a_n1458_n3888# 0.055941f
C67 minus.n20 a_n1458_n3888# 0.019592f
C68 minus.n21 a_n1458_n3888# 0.187605f
C69 minus.n22 a_n1458_n3888# 0.019592f
C70 minus.n23 a_n1458_n3888# 0.187605f
C71 minus.t7 a_n1458_n3888# 0.477901f
C72 minus.n24 a_n1458_n3888# 0.203612f
C73 minus.n25 a_n1458_n3888# 0.35979f
C74 minus.n26 a_n1458_n3888# 2.46665f
C75 drain_left.t1 a_n1458_n3888# 0.455347f
C76 drain_left.t11 a_n1458_n3888# 0.455347f
C77 drain_left.n0 a_n1458_n3888# 4.11868f
C78 drain_left.t2 a_n1458_n3888# 0.455347f
C79 drain_left.t10 a_n1458_n3888# 0.455347f
C80 drain_left.n1 a_n1458_n3888# 4.1158f
C81 drain_left.t8 a_n1458_n3888# 0.455347f
C82 drain_left.t9 a_n1458_n3888# 0.455347f
C83 drain_left.n2 a_n1458_n3888# 4.11868f
C84 drain_left.n3 a_n1458_n3888# 3.23841f
C85 drain_left.t5 a_n1458_n3888# 0.455347f
C86 drain_left.t7 a_n1458_n3888# 0.455347f
C87 drain_left.n4 a_n1458_n3888# 4.11911f
C88 drain_left.t0 a_n1458_n3888# 0.455347f
C89 drain_left.t3 a_n1458_n3888# 0.455347f
C90 drain_left.n5 a_n1458_n3888# 4.11581f
C91 drain_left.n6 a_n1458_n3888# 0.867664f
C92 drain_left.t4 a_n1458_n3888# 0.455347f
C93 drain_left.t6 a_n1458_n3888# 0.455347f
C94 drain_left.n7 a_n1458_n3888# 4.11579f
C95 drain_left.n8 a_n1458_n3888# 0.742149f
C96 source.t17 a_n1458_n3888# 3.97537f
C97 source.n0 a_n1458_n3888# 1.8279f
C98 source.t16 a_n1458_n3888# 0.354734f
C99 source.t14 a_n1458_n3888# 0.354734f
C100 source.n1 a_n1458_n3888# 3.11604f
C101 source.n2 a_n1458_n3888# 0.382899f
C102 source.t15 a_n1458_n3888# 0.354734f
C103 source.t18 a_n1458_n3888# 0.354734f
C104 source.n3 a_n1458_n3888# 3.11604f
C105 source.n4 a_n1458_n3888# 0.382899f
C106 source.t22 a_n1458_n3888# 3.97537f
C107 source.n5 a_n1458_n3888# 0.492272f
C108 source.t11 a_n1458_n3888# 3.97537f
C109 source.n6 a_n1458_n3888# 0.492272f
C110 source.t1 a_n1458_n3888# 0.354734f
C111 source.t5 a_n1458_n3888# 0.354734f
C112 source.n7 a_n1458_n3888# 3.11604f
C113 source.n8 a_n1458_n3888# 0.382899f
C114 source.t0 a_n1458_n3888# 0.354734f
C115 source.t3 a_n1458_n3888# 0.354734f
C116 source.n9 a_n1458_n3888# 3.11604f
C117 source.n10 a_n1458_n3888# 0.382899f
C118 source.t7 a_n1458_n3888# 3.97537f
C119 source.n11 a_n1458_n3888# 2.32224f
C120 source.t21 a_n1458_n3888# 3.97537f
C121 source.n12 a_n1458_n3888# 2.32225f
C122 source.t19 a_n1458_n3888# 0.354734f
C123 source.t12 a_n1458_n3888# 0.354734f
C124 source.n13 a_n1458_n3888# 3.11604f
C125 source.n14 a_n1458_n3888# 0.382903f
C126 source.t20 a_n1458_n3888# 0.354734f
C127 source.t13 a_n1458_n3888# 0.354734f
C128 source.n15 a_n1458_n3888# 3.11604f
C129 source.n16 a_n1458_n3888# 0.382903f
C130 source.t23 a_n1458_n3888# 3.97537f
C131 source.n17 a_n1458_n3888# 0.492277f
C132 source.t6 a_n1458_n3888# 3.97537f
C133 source.n18 a_n1458_n3888# 0.492277f
C134 source.t4 a_n1458_n3888# 0.354734f
C135 source.t9 a_n1458_n3888# 0.354734f
C136 source.n19 a_n1458_n3888# 3.11604f
C137 source.n20 a_n1458_n3888# 0.382903f
C138 source.t10 a_n1458_n3888# 0.354734f
C139 source.t2 a_n1458_n3888# 0.354734f
C140 source.n21 a_n1458_n3888# 3.11604f
C141 source.n22 a_n1458_n3888# 0.382903f
C142 source.t8 a_n1458_n3888# 3.97537f
C143 source.n23 a_n1458_n3888# 0.654549f
C144 source.n24 a_n1458_n3888# 2.18333f
C145 plus.n0 a_n1458_n3888# 0.056832f
C146 plus.t7 a_n1458_n3888# 0.480992f
C147 plus.t8 a_n1458_n3888# 0.480992f
C148 plus.t11 a_n1458_n3888# 0.480992f
C149 plus.n1 a_n1458_n3888# 0.190592f
C150 plus.t6 a_n1458_n3888# 0.48551f
C151 plus.n2 a_n1458_n3888# 0.206934f
C152 plus.t4 a_n1458_n3888# 0.480992f
C153 plus.n3 a_n1458_n3888# 0.190592f
C154 plus.n4 a_n1458_n3888# 0.019904f
C155 plus.n5 a_n1458_n3888# 0.125846f
C156 plus.n6 a_n1458_n3888# 0.056832f
C157 plus.n7 a_n1458_n3888# 0.019904f
C158 plus.n8 a_n1458_n3888# 0.190592f
C159 plus.n9 a_n1458_n3888# 0.019904f
C160 plus.n10 a_n1458_n3888# 0.190592f
C161 plus.t5 a_n1458_n3888# 0.48551f
C162 plus.n11 a_n1458_n3888# 0.206853f
C163 plus.n12 a_n1458_n3888# 0.712146f
C164 plus.n13 a_n1458_n3888# 0.056832f
C165 plus.t10 a_n1458_n3888# 0.48551f
C166 plus.t0 a_n1458_n3888# 0.480992f
C167 plus.t9 a_n1458_n3888# 0.480992f
C168 plus.t1 a_n1458_n3888# 0.480992f
C169 plus.n14 a_n1458_n3888# 0.190592f
C170 plus.t2 a_n1458_n3888# 0.48551f
C171 plus.n15 a_n1458_n3888# 0.206934f
C172 plus.t3 a_n1458_n3888# 0.480992f
C173 plus.n16 a_n1458_n3888# 0.190592f
C174 plus.n17 a_n1458_n3888# 0.019904f
C175 plus.n18 a_n1458_n3888# 0.125846f
C176 plus.n19 a_n1458_n3888# 0.056832f
C177 plus.n20 a_n1458_n3888# 0.019904f
C178 plus.n21 a_n1458_n3888# 0.190592f
C179 plus.n22 a_n1458_n3888# 0.019904f
C180 plus.n23 a_n1458_n3888# 0.190592f
C181 plus.n24 a_n1458_n3888# 0.206853f
C182 plus.n25 a_n1458_n3888# 1.69143f
.ends

