* NGSPICE file created from diffpair521.ext - technology: sky130A

.subckt diffpair521 minus drain_right drain_left source plus
X0 source plus drain_left a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X1 drain_left plus source a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X2 source minus drain_right a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X3 source plus drain_left a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X4 drain_right minus source a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X5 source minus drain_right a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X6 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X7 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X8 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X9 drain_right minus source a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X10 drain_left plus source a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X11 a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# a_n1214_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
.ends

