* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X1 source.t19 plus.t0 drain_left.t1 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X2 drain_right.t9 minus.t0 source.t2 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X3 drain_right.t8 minus.t1 source.t3 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X4 source.t6 minus.t2 drain_right.t7 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 drain_left.t2 plus.t1 source.t18 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X6 source.t8 minus.t3 drain_right.t6 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X7 drain_right.t5 minus.t4 source.t0 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 drain_left.t0 plus.t2 source.t17 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X9 source.t16 plus.t3 drain_left.t5 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X10 source.t9 minus.t5 drain_right.t4 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 drain_left.t6 plus.t4 source.t15 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X12 drain_left.t7 plus.t5 source.t14 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 drain_right.t3 minus.t6 source.t1 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X14 source.t13 plus.t6 drain_left.t8 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 drain_left.t3 plus.t7 source.t12 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X16 a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X17 drain_right.t2 minus.t7 source.t5 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X18 a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X19 source.t11 plus.t8 drain_left.t4 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X20 source.t7 minus.t8 drain_right.t1 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 drain_right.t0 minus.t9 source.t4 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X22 a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X23 drain_left.t9 plus.t9 source.t10 a_n1832_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n6 plus.n1 161.3
R1 plus.n7 plus.n0 161.3
R2 plus.n9 plus.n8 161.3
R3 plus.n16 plus.n11 161.3
R4 plus.n17 plus.n10 161.3
R5 plus.n19 plus.n18 161.3
R6 plus.n3 plus.t7 131.839
R7 plus.n13 plus.t2 131.839
R8 plus.n8 plus.t1 105.638
R9 plus.n6 plus.t3 105.638
R10 plus.n5 plus.t5 105.638
R11 plus.n4 plus.t6 105.638
R12 plus.n18 plus.t4 105.638
R13 plus.n16 plus.t8 105.638
R14 plus.n15 plus.t9 105.638
R15 plus.n14 plus.t0 105.638
R16 plus.n5 plus.n2 80.6037
R17 plus.n15 plus.n12 80.6037
R18 plus.n6 plus.n5 48.2005
R19 plus.n5 plus.n4 48.2005
R20 plus.n16 plus.n15 48.2005
R21 plus.n15 plus.n14 48.2005
R22 plus.n8 plus.n7 45.2793
R23 plus.n18 plus.n17 45.2793
R24 plus.n3 plus.n2 45.1669
R25 plus.n13 plus.n12 45.1669
R26 plus plus.n19 25.8759
R27 plus.n4 plus.n3 14.3992
R28 plus.n14 plus.n13 14.3992
R29 plus plus.n9 8.07815
R30 plus.n7 plus.n6 2.92171
R31 plus.n17 plus.n16 2.92171
R32 plus.n2 plus.n1 0.285035
R33 plus.n12 plus.n11 0.285035
R34 plus.n1 plus.n0 0.189894
R35 plus.n9 plus.n0 0.189894
R36 plus.n19 plus.n10 0.189894
R37 plus.n11 plus.n10 0.189894
R38 drain_left.n5 drain_left.t3 260.735
R39 drain_left.n1 drain_left.t6 260.733
R40 drain_left.n3 drain_left.n2 240.678
R41 drain_left.n7 drain_left.n6 240.132
R42 drain_left.n5 drain_left.n4 240.132
R43 drain_left.n1 drain_left.n0 240.131
R44 drain_left drain_left.n3 22.4411
R45 drain_left.n2 drain_left.t1 19.8005
R46 drain_left.n2 drain_left.t0 19.8005
R47 drain_left.n0 drain_left.t4 19.8005
R48 drain_left.n0 drain_left.t9 19.8005
R49 drain_left.n6 drain_left.t5 19.8005
R50 drain_left.n6 drain_left.t2 19.8005
R51 drain_left.n4 drain_left.t8 19.8005
R52 drain_left.n4 drain_left.t7 19.8005
R53 drain_left drain_left.n7 6.45494
R54 drain_left.n7 drain_left.n5 0.802224
R55 drain_left.n3 drain_left.n1 0.145585
R56 source.n0 source.t18 243.255
R57 source.n5 source.t1 243.255
R58 source.n19 source.t5 243.254
R59 source.n14 source.t17 243.254
R60 source.n2 source.n1 223.454
R61 source.n4 source.n3 223.454
R62 source.n7 source.n6 223.454
R63 source.n9 source.n8 223.454
R64 source.n18 source.n17 223.453
R65 source.n16 source.n15 223.453
R66 source.n13 source.n12 223.453
R67 source.n11 source.n10 223.453
R68 source.n17 source.t3 19.8005
R69 source.n17 source.t7 19.8005
R70 source.n15 source.t4 19.8005
R71 source.n15 source.t6 19.8005
R72 source.n12 source.t10 19.8005
R73 source.n12 source.t19 19.8005
R74 source.n10 source.t15 19.8005
R75 source.n10 source.t11 19.8005
R76 source.n1 source.t14 19.8005
R77 source.n1 source.t16 19.8005
R78 source.n3 source.t12 19.8005
R79 source.n3 source.t13 19.8005
R80 source.n6 source.t0 19.8005
R81 source.n6 source.t9 19.8005
R82 source.n8 source.t2 19.8005
R83 source.n8 source.t8 19.8005
R84 source.n11 source.n9 14.5578
R85 source.n20 source.n0 8.09232
R86 source.n20 source.n19 5.66429
R87 source.n5 source.n4 0.87119
R88 source.n16 source.n14 0.87119
R89 source.n9 source.n7 0.802224
R90 source.n7 source.n5 0.802224
R91 source.n4 source.n2 0.802224
R92 source.n2 source.n0 0.802224
R93 source.n13 source.n11 0.802224
R94 source.n14 source.n13 0.802224
R95 source.n18 source.n16 0.802224
R96 source.n19 source.n18 0.802224
R97 source source.n20 0.188
R98 minus.n9 minus.n8 161.3
R99 minus.n7 minus.n0 161.3
R100 minus.n6 minus.n5 161.3
R101 minus.n19 minus.n18 161.3
R102 minus.n17 minus.n10 161.3
R103 minus.n16 minus.n15 161.3
R104 minus.n3 minus.t6 131.839
R105 minus.n13 minus.t9 131.839
R106 minus.n2 minus.t5 105.638
R107 minus.n1 minus.t4 105.638
R108 minus.n6 minus.t3 105.638
R109 minus.n8 minus.t0 105.638
R110 minus.n12 minus.t2 105.638
R111 minus.n11 minus.t1 105.638
R112 minus.n16 minus.t8 105.638
R113 minus.n18 minus.t7 105.638
R114 minus.n4 minus.n1 80.6037
R115 minus.n14 minus.n11 80.6037
R116 minus.n2 minus.n1 48.2005
R117 minus.n6 minus.n1 48.2005
R118 minus.n12 minus.n11 48.2005
R119 minus.n16 minus.n11 48.2005
R120 minus.n8 minus.n7 45.2793
R121 minus.n18 minus.n17 45.2793
R122 minus.n4 minus.n3 45.1669
R123 minus.n14 minus.n13 45.1669
R124 minus.n20 minus.n9 27.8282
R125 minus.n3 minus.n2 14.3992
R126 minus.n13 minus.n12 14.3992
R127 minus.n20 minus.n19 6.60088
R128 minus.n7 minus.n6 2.92171
R129 minus.n17 minus.n16 2.92171
R130 minus.n5 minus.n4 0.285035
R131 minus.n15 minus.n14 0.285035
R132 minus.n9 minus.n0 0.189894
R133 minus.n5 minus.n0 0.189894
R134 minus.n15 minus.n10 0.189894
R135 minus.n19 minus.n10 0.189894
R136 minus minus.n20 0.188
R137 drain_right.n1 drain_right.t0 260.733
R138 drain_right.n7 drain_right.t9 259.933
R139 drain_right.n6 drain_right.n4 240.935
R140 drain_right.n3 drain_right.n2 240.678
R141 drain_right.n6 drain_right.n5 240.132
R142 drain_right.n1 drain_right.n0 240.131
R143 drain_right drain_right.n3 21.8878
R144 drain_right.n2 drain_right.t1 19.8005
R145 drain_right.n2 drain_right.t2 19.8005
R146 drain_right.n0 drain_right.t7 19.8005
R147 drain_right.n0 drain_right.t8 19.8005
R148 drain_right.n4 drain_right.t4 19.8005
R149 drain_right.n4 drain_right.t3 19.8005
R150 drain_right.n5 drain_right.t6 19.8005
R151 drain_right.n5 drain_right.t5 19.8005
R152 drain_right drain_right.n7 6.05408
R153 drain_right.n7 drain_right.n6 0.802224
R154 drain_right.n3 drain_right.n1 0.145585
C0 drain_left drain_right 0.906277f
C1 minus source 1.29358f
C2 plus minus 3.40204f
C3 plus source 1.30749f
C4 drain_left minus 0.179981f
C5 drain_right minus 0.903434f
C6 drain_left source 3.52913f
C7 drain_right source 3.52894f
C8 drain_left plus 1.08085f
C9 drain_right plus 0.342246f
C10 drain_right a_n1832_n1088# 3.44356f
C11 drain_left a_n1832_n1088# 3.686267f
C12 source a_n1832_n1088# 2.164418f
C13 minus a_n1832_n1088# 6.237153f
C14 plus a_n1832_n1088# 6.862583f
C15 drain_right.t0 a_n1832_n1088# 0.096346f
C16 drain_right.t7 a_n1832_n1088# 0.015476f
C17 drain_right.t8 a_n1832_n1088# 0.015476f
C18 drain_right.n0 a_n1832_n1088# 0.060135f
C19 drain_right.n1 a_n1832_n1088# 0.401259f
C20 drain_right.t1 a_n1832_n1088# 0.015476f
C21 drain_right.t2 a_n1832_n1088# 0.015476f
C22 drain_right.n2 a_n1832_n1088# 0.060658f
C23 drain_right.n3 a_n1832_n1088# 0.729251f
C24 drain_right.t4 a_n1832_n1088# 0.015476f
C25 drain_right.t3 a_n1832_n1088# 0.015476f
C26 drain_right.n4 a_n1832_n1088# 0.060953f
C27 drain_right.t6 a_n1832_n1088# 0.015476f
C28 drain_right.t5 a_n1832_n1088# 0.015476f
C29 drain_right.n5 a_n1832_n1088# 0.060135f
C30 drain_right.n6 a_n1832_n1088# 0.483344f
C31 drain_right.t9 a_n1832_n1088# 0.095725f
C32 drain_right.n7 a_n1832_n1088# 0.377917f
C33 minus.n0 a_n1832_n1088# 0.02947f
C34 minus.t4 a_n1832_n1088# 0.059959f
C35 minus.n1 a_n1832_n1088# 0.067718f
C36 minus.t3 a_n1832_n1088# 0.059959f
C37 minus.t6 a_n1832_n1088# 0.072074f
C38 minus.t5 a_n1832_n1088# 0.059959f
C39 minus.n2 a_n1832_n1088# 0.067223f
C40 minus.n3 a_n1832_n1088# 0.050279f
C41 minus.n4 a_n1832_n1088# 0.142442f
C42 minus.n5 a_n1832_n1088# 0.039324f
C43 minus.n6 a_n1832_n1088# 0.061394f
C44 minus.n7 a_n1832_n1088# 0.006687f
C45 minus.t0 a_n1832_n1088# 0.059959f
C46 minus.n8 a_n1832_n1088# 0.060667f
C47 minus.n9 a_n1832_n1088# 0.675584f
C48 minus.n10 a_n1832_n1088# 0.02947f
C49 minus.t1 a_n1832_n1088# 0.059959f
C50 minus.n11 a_n1832_n1088# 0.067718f
C51 minus.t9 a_n1832_n1088# 0.072074f
C52 minus.t2 a_n1832_n1088# 0.059959f
C53 minus.n12 a_n1832_n1088# 0.067223f
C54 minus.n13 a_n1832_n1088# 0.050279f
C55 minus.n14 a_n1832_n1088# 0.142442f
C56 minus.n15 a_n1832_n1088# 0.039324f
C57 minus.t8 a_n1832_n1088# 0.059959f
C58 minus.n16 a_n1832_n1088# 0.061394f
C59 minus.n17 a_n1832_n1088# 0.006687f
C60 minus.t7 a_n1832_n1088# 0.059959f
C61 minus.n18 a_n1832_n1088# 0.060667f
C62 minus.n19 a_n1832_n1088# 0.199638f
C63 minus.n20 a_n1832_n1088# 0.831192f
C64 source.t18 a_n1832_n1088# 0.116658f
C65 source.n0 a_n1832_n1088# 0.540416f
C66 source.t14 a_n1832_n1088# 0.02096f
C67 source.t16 a_n1832_n1088# 0.02096f
C68 source.n1 a_n1832_n1088# 0.067975f
C69 source.n2 a_n1832_n1088# 0.299936f
C70 source.t12 a_n1832_n1088# 0.02096f
C71 source.t13 a_n1832_n1088# 0.02096f
C72 source.n3 a_n1832_n1088# 0.067975f
C73 source.n4 a_n1832_n1088# 0.30583f
C74 source.t1 a_n1832_n1088# 0.116658f
C75 source.n5 a_n1832_n1088# 0.314309f
C76 source.t0 a_n1832_n1088# 0.02096f
C77 source.t9 a_n1832_n1088# 0.02096f
C78 source.n6 a_n1832_n1088# 0.067975f
C79 source.n7 a_n1832_n1088# 0.299936f
C80 source.t2 a_n1832_n1088# 0.02096f
C81 source.t8 a_n1832_n1088# 0.02096f
C82 source.n8 a_n1832_n1088# 0.067975f
C83 source.n9 a_n1832_n1088# 0.817689f
C84 source.t15 a_n1832_n1088# 0.02096f
C85 source.t11 a_n1832_n1088# 0.02096f
C86 source.n10 a_n1832_n1088# 0.067975f
C87 source.n11 a_n1832_n1088# 0.817689f
C88 source.t10 a_n1832_n1088# 0.02096f
C89 source.t19 a_n1832_n1088# 0.02096f
C90 source.n12 a_n1832_n1088# 0.067975f
C91 source.n13 a_n1832_n1088# 0.299936f
C92 source.t17 a_n1832_n1088# 0.116658f
C93 source.n14 a_n1832_n1088# 0.31431f
C94 source.t4 a_n1832_n1088# 0.02096f
C95 source.t6 a_n1832_n1088# 0.02096f
C96 source.n15 a_n1832_n1088# 0.067975f
C97 source.n16 a_n1832_n1088# 0.30583f
C98 source.t3 a_n1832_n1088# 0.02096f
C99 source.t7 a_n1832_n1088# 0.02096f
C100 source.n17 a_n1832_n1088# 0.067975f
C101 source.n18 a_n1832_n1088# 0.299936f
C102 source.t5 a_n1832_n1088# 0.116658f
C103 source.n19 a_n1832_n1088# 0.44729f
C104 source.n20 a_n1832_n1088# 0.546459f
C105 drain_left.t6 a_n1832_n1088# 0.094282f
C106 drain_left.t4 a_n1832_n1088# 0.015144f
C107 drain_left.t9 a_n1832_n1088# 0.015144f
C108 drain_left.n0 a_n1832_n1088# 0.058847f
C109 drain_left.n1 a_n1832_n1088# 0.392664f
C110 drain_left.t1 a_n1832_n1088# 0.015144f
C111 drain_left.t0 a_n1832_n1088# 0.015144f
C112 drain_left.n2 a_n1832_n1088# 0.059359f
C113 drain_left.n3 a_n1832_n1088# 0.750679f
C114 drain_left.t3 a_n1832_n1088# 0.094282f
C115 drain_left.t8 a_n1832_n1088# 0.015144f
C116 drain_left.t7 a_n1832_n1088# 0.015144f
C117 drain_left.n4 a_n1832_n1088# 0.058847f
C118 drain_left.n5 a_n1832_n1088# 0.430151f
C119 drain_left.t5 a_n1832_n1088# 0.015144f
C120 drain_left.t2 a_n1832_n1088# 0.015144f
C121 drain_left.n6 a_n1832_n1088# 0.058847f
C122 drain_left.n7 a_n1832_n1088# 0.40015f
C123 plus.n0 a_n1832_n1088# 0.029996f
C124 plus.t1 a_n1832_n1088# 0.061029f
C125 plus.t3 a_n1832_n1088# 0.061029f
C126 plus.n1 a_n1832_n1088# 0.040026f
C127 plus.t5 a_n1832_n1088# 0.061029f
C128 plus.n2 a_n1832_n1088# 0.144983f
C129 plus.t6 a_n1832_n1088# 0.061029f
C130 plus.t7 a_n1832_n1088# 0.07336f
C131 plus.n3 a_n1832_n1088# 0.051176f
C132 plus.n4 a_n1832_n1088# 0.068423f
C133 plus.n5 a_n1832_n1088# 0.068926f
C134 plus.n6 a_n1832_n1088# 0.062489f
C135 plus.n7 a_n1832_n1088# 0.006807f
C136 plus.n8 a_n1832_n1088# 0.06175f
C137 plus.n9 a_n1832_n1088# 0.21313f
C138 plus.n10 a_n1832_n1088# 0.029996f
C139 plus.t4 a_n1832_n1088# 0.061029f
C140 plus.n11 a_n1832_n1088# 0.040026f
C141 plus.t8 a_n1832_n1088# 0.061029f
C142 plus.n12 a_n1832_n1088# 0.144983f
C143 plus.t9 a_n1832_n1088# 0.061029f
C144 plus.t2 a_n1832_n1088# 0.07336f
C145 plus.n13 a_n1832_n1088# 0.051176f
C146 plus.t0 a_n1832_n1088# 0.061029f
C147 plus.n14 a_n1832_n1088# 0.068423f
C148 plus.n15 a_n1832_n1088# 0.068926f
C149 plus.n16 a_n1832_n1088# 0.062489f
C150 plus.n17 a_n1832_n1088# 0.006807f
C151 plus.n18 a_n1832_n1088# 0.06175f
C152 plus.n19 a_n1832_n1088# 0.667104f
.ends

