* NGSPICE file created from diffpair273.ext - technology: sky130A

.subckt diffpair273 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t13 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t15 plus.t0 drain_left.t7 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 source.t0 plus.t1 drain_left.t6 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X3 source.t1 plus.t2 drain_left.t5 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X4 drain_right.t6 minus.t1 source.t12 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X5 drain_right.t5 minus.t2 source.t7 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X6 a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X7 drain_left.t4 plus.t3 source.t6 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X8 drain_left.t3 plus.t4 source.t5 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X9 drain_left.t2 plus.t5 source.t2 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 source.t10 minus.t3 drain_right.t4 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X11 drain_right.t3 minus.t4 source.t8 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X12 source.t11 minus.t5 drain_right.t2 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X13 source.t9 minus.t6 drain_right.t1 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X14 source.t4 plus.t6 drain_left.t1 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X15 a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X16 source.t14 minus.t7 drain_right.t0 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X17 a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X18 drain_left.t0 plus.t7 source.t3 a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X19 a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# a_n1346_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
R0 minus.n7 minus.t3 614.915
R1 minus.n2 minus.t4 614.915
R2 minus.n16 minus.t1 614.915
R3 minus.n11 minus.t6 614.915
R4 minus.n6 minus.t0 586.433
R5 minus.n1 minus.t7 586.433
R6 minus.n15 minus.t5 586.433
R7 minus.n10 minus.t2 586.433
R8 minus.n3 minus.n2 161.489
R9 minus.n12 minus.n11 161.489
R10 minus.n8 minus.n7 161.3
R11 minus.n5 minus.n0 161.3
R12 minus.n4 minus.n3 161.3
R13 minus.n17 minus.n16 161.3
R14 minus.n14 minus.n9 161.3
R15 minus.n13 minus.n12 161.3
R16 minus.n5 minus.n4 73.0308
R17 minus.n14 minus.n13 73.0308
R18 minus.n7 minus.n6 63.5369
R19 minus.n2 minus.n1 63.5369
R20 minus.n11 minus.n10 63.5369
R21 minus.n16 minus.n15 63.5369
R22 minus.n18 minus.n8 29.6369
R23 minus.n6 minus.n5 9.49444
R24 minus.n4 minus.n1 9.49444
R25 minus.n13 minus.n10 9.49444
R26 minus.n15 minus.n14 9.49444
R27 minus.n18 minus.n17 6.46262
R28 minus.n8 minus.n0 0.189894
R29 minus.n3 minus.n0 0.189894
R30 minus.n12 minus.n9 0.189894
R31 minus.n17 minus.n9 0.189894
R32 minus minus.n18 0.188
R33 source.n258 source.n232 289.615
R34 source.n224 source.n198 289.615
R35 source.n192 source.n166 289.615
R36 source.n158 source.n132 289.615
R37 source.n26 source.n0 289.615
R38 source.n60 source.n34 289.615
R39 source.n92 source.n66 289.615
R40 source.n126 source.n100 289.615
R41 source.n243 source.n242 185
R42 source.n240 source.n239 185
R43 source.n249 source.n248 185
R44 source.n251 source.n250 185
R45 source.n236 source.n235 185
R46 source.n257 source.n256 185
R47 source.n259 source.n258 185
R48 source.n209 source.n208 185
R49 source.n206 source.n205 185
R50 source.n215 source.n214 185
R51 source.n217 source.n216 185
R52 source.n202 source.n201 185
R53 source.n223 source.n222 185
R54 source.n225 source.n224 185
R55 source.n177 source.n176 185
R56 source.n174 source.n173 185
R57 source.n183 source.n182 185
R58 source.n185 source.n184 185
R59 source.n170 source.n169 185
R60 source.n191 source.n190 185
R61 source.n193 source.n192 185
R62 source.n143 source.n142 185
R63 source.n140 source.n139 185
R64 source.n149 source.n148 185
R65 source.n151 source.n150 185
R66 source.n136 source.n135 185
R67 source.n157 source.n156 185
R68 source.n159 source.n158 185
R69 source.n27 source.n26 185
R70 source.n25 source.n24 185
R71 source.n4 source.n3 185
R72 source.n19 source.n18 185
R73 source.n17 source.n16 185
R74 source.n8 source.n7 185
R75 source.n11 source.n10 185
R76 source.n61 source.n60 185
R77 source.n59 source.n58 185
R78 source.n38 source.n37 185
R79 source.n53 source.n52 185
R80 source.n51 source.n50 185
R81 source.n42 source.n41 185
R82 source.n45 source.n44 185
R83 source.n93 source.n92 185
R84 source.n91 source.n90 185
R85 source.n70 source.n69 185
R86 source.n85 source.n84 185
R87 source.n83 source.n82 185
R88 source.n74 source.n73 185
R89 source.n77 source.n76 185
R90 source.n127 source.n126 185
R91 source.n125 source.n124 185
R92 source.n104 source.n103 185
R93 source.n119 source.n118 185
R94 source.n117 source.n116 185
R95 source.n108 source.n107 185
R96 source.n111 source.n110 185
R97 source.t12 source.n241 147.661
R98 source.t9 source.n207 147.661
R99 source.t5 source.n175 147.661
R100 source.t1 source.n141 147.661
R101 source.t3 source.n9 147.661
R102 source.t0 source.n43 147.661
R103 source.t8 source.n75 147.661
R104 source.t10 source.n109 147.661
R105 source.n242 source.n239 104.615
R106 source.n249 source.n239 104.615
R107 source.n250 source.n249 104.615
R108 source.n250 source.n235 104.615
R109 source.n257 source.n235 104.615
R110 source.n258 source.n257 104.615
R111 source.n208 source.n205 104.615
R112 source.n215 source.n205 104.615
R113 source.n216 source.n215 104.615
R114 source.n216 source.n201 104.615
R115 source.n223 source.n201 104.615
R116 source.n224 source.n223 104.615
R117 source.n176 source.n173 104.615
R118 source.n183 source.n173 104.615
R119 source.n184 source.n183 104.615
R120 source.n184 source.n169 104.615
R121 source.n191 source.n169 104.615
R122 source.n192 source.n191 104.615
R123 source.n142 source.n139 104.615
R124 source.n149 source.n139 104.615
R125 source.n150 source.n149 104.615
R126 source.n150 source.n135 104.615
R127 source.n157 source.n135 104.615
R128 source.n158 source.n157 104.615
R129 source.n26 source.n25 104.615
R130 source.n25 source.n3 104.615
R131 source.n18 source.n3 104.615
R132 source.n18 source.n17 104.615
R133 source.n17 source.n7 104.615
R134 source.n10 source.n7 104.615
R135 source.n60 source.n59 104.615
R136 source.n59 source.n37 104.615
R137 source.n52 source.n37 104.615
R138 source.n52 source.n51 104.615
R139 source.n51 source.n41 104.615
R140 source.n44 source.n41 104.615
R141 source.n92 source.n91 104.615
R142 source.n91 source.n69 104.615
R143 source.n84 source.n69 104.615
R144 source.n84 source.n83 104.615
R145 source.n83 source.n73 104.615
R146 source.n76 source.n73 104.615
R147 source.n126 source.n125 104.615
R148 source.n125 source.n103 104.615
R149 source.n118 source.n103 104.615
R150 source.n118 source.n117 104.615
R151 source.n117 source.n107 104.615
R152 source.n110 source.n107 104.615
R153 source.n242 source.t12 52.3082
R154 source.n208 source.t9 52.3082
R155 source.n176 source.t5 52.3082
R156 source.n142 source.t1 52.3082
R157 source.n10 source.t3 52.3082
R158 source.n44 source.t0 52.3082
R159 source.n76 source.t8 52.3082
R160 source.n110 source.t10 52.3082
R161 source.n33 source.n32 50.512
R162 source.n99 source.n98 50.512
R163 source.n231 source.n230 50.5119
R164 source.n165 source.n164 50.5119
R165 source.n263 source.n262 32.1853
R166 source.n229 source.n228 32.1853
R167 source.n197 source.n196 32.1853
R168 source.n163 source.n162 32.1853
R169 source.n31 source.n30 32.1853
R170 source.n65 source.n64 32.1853
R171 source.n97 source.n96 32.1853
R172 source.n131 source.n130 32.1853
R173 source.n163 source.n131 17.2854
R174 source.n243 source.n241 15.6674
R175 source.n209 source.n207 15.6674
R176 source.n177 source.n175 15.6674
R177 source.n143 source.n141 15.6674
R178 source.n11 source.n9 15.6674
R179 source.n45 source.n43 15.6674
R180 source.n77 source.n75 15.6674
R181 source.n111 source.n109 15.6674
R182 source.n244 source.n240 12.8005
R183 source.n210 source.n206 12.8005
R184 source.n178 source.n174 12.8005
R185 source.n144 source.n140 12.8005
R186 source.n12 source.n8 12.8005
R187 source.n46 source.n42 12.8005
R188 source.n78 source.n74 12.8005
R189 source.n112 source.n108 12.8005
R190 source.n248 source.n247 12.0247
R191 source.n214 source.n213 12.0247
R192 source.n182 source.n181 12.0247
R193 source.n148 source.n147 12.0247
R194 source.n16 source.n15 12.0247
R195 source.n50 source.n49 12.0247
R196 source.n82 source.n81 12.0247
R197 source.n116 source.n115 12.0247
R198 source.n264 source.n31 11.7509
R199 source.n251 source.n238 11.249
R200 source.n217 source.n204 11.249
R201 source.n185 source.n172 11.249
R202 source.n151 source.n138 11.249
R203 source.n19 source.n6 11.249
R204 source.n53 source.n40 11.249
R205 source.n85 source.n72 11.249
R206 source.n119 source.n106 11.249
R207 source.n252 source.n236 10.4732
R208 source.n218 source.n202 10.4732
R209 source.n186 source.n170 10.4732
R210 source.n152 source.n136 10.4732
R211 source.n20 source.n4 10.4732
R212 source.n54 source.n38 10.4732
R213 source.n86 source.n70 10.4732
R214 source.n120 source.n104 10.4732
R215 source.n256 source.n255 9.69747
R216 source.n222 source.n221 9.69747
R217 source.n190 source.n189 9.69747
R218 source.n156 source.n155 9.69747
R219 source.n24 source.n23 9.69747
R220 source.n58 source.n57 9.69747
R221 source.n90 source.n89 9.69747
R222 source.n124 source.n123 9.69747
R223 source.n262 source.n261 9.45567
R224 source.n228 source.n227 9.45567
R225 source.n196 source.n195 9.45567
R226 source.n162 source.n161 9.45567
R227 source.n30 source.n29 9.45567
R228 source.n64 source.n63 9.45567
R229 source.n96 source.n95 9.45567
R230 source.n130 source.n129 9.45567
R231 source.n261 source.n260 9.3005
R232 source.n234 source.n233 9.3005
R233 source.n255 source.n254 9.3005
R234 source.n253 source.n252 9.3005
R235 source.n238 source.n237 9.3005
R236 source.n247 source.n246 9.3005
R237 source.n245 source.n244 9.3005
R238 source.n227 source.n226 9.3005
R239 source.n200 source.n199 9.3005
R240 source.n221 source.n220 9.3005
R241 source.n219 source.n218 9.3005
R242 source.n204 source.n203 9.3005
R243 source.n213 source.n212 9.3005
R244 source.n211 source.n210 9.3005
R245 source.n195 source.n194 9.3005
R246 source.n168 source.n167 9.3005
R247 source.n189 source.n188 9.3005
R248 source.n187 source.n186 9.3005
R249 source.n172 source.n171 9.3005
R250 source.n181 source.n180 9.3005
R251 source.n179 source.n178 9.3005
R252 source.n161 source.n160 9.3005
R253 source.n134 source.n133 9.3005
R254 source.n155 source.n154 9.3005
R255 source.n153 source.n152 9.3005
R256 source.n138 source.n137 9.3005
R257 source.n147 source.n146 9.3005
R258 source.n145 source.n144 9.3005
R259 source.n29 source.n28 9.3005
R260 source.n2 source.n1 9.3005
R261 source.n23 source.n22 9.3005
R262 source.n21 source.n20 9.3005
R263 source.n6 source.n5 9.3005
R264 source.n15 source.n14 9.3005
R265 source.n13 source.n12 9.3005
R266 source.n63 source.n62 9.3005
R267 source.n36 source.n35 9.3005
R268 source.n57 source.n56 9.3005
R269 source.n55 source.n54 9.3005
R270 source.n40 source.n39 9.3005
R271 source.n49 source.n48 9.3005
R272 source.n47 source.n46 9.3005
R273 source.n95 source.n94 9.3005
R274 source.n68 source.n67 9.3005
R275 source.n89 source.n88 9.3005
R276 source.n87 source.n86 9.3005
R277 source.n72 source.n71 9.3005
R278 source.n81 source.n80 9.3005
R279 source.n79 source.n78 9.3005
R280 source.n129 source.n128 9.3005
R281 source.n102 source.n101 9.3005
R282 source.n123 source.n122 9.3005
R283 source.n121 source.n120 9.3005
R284 source.n106 source.n105 9.3005
R285 source.n115 source.n114 9.3005
R286 source.n113 source.n112 9.3005
R287 source.n259 source.n234 8.92171
R288 source.n225 source.n200 8.92171
R289 source.n193 source.n168 8.92171
R290 source.n159 source.n134 8.92171
R291 source.n27 source.n2 8.92171
R292 source.n61 source.n36 8.92171
R293 source.n93 source.n68 8.92171
R294 source.n127 source.n102 8.92171
R295 source.n260 source.n232 8.14595
R296 source.n226 source.n198 8.14595
R297 source.n194 source.n166 8.14595
R298 source.n160 source.n132 8.14595
R299 source.n28 source.n0 8.14595
R300 source.n62 source.n34 8.14595
R301 source.n94 source.n66 8.14595
R302 source.n128 source.n100 8.14595
R303 source.n262 source.n232 5.81868
R304 source.n228 source.n198 5.81868
R305 source.n196 source.n166 5.81868
R306 source.n162 source.n132 5.81868
R307 source.n30 source.n0 5.81868
R308 source.n64 source.n34 5.81868
R309 source.n96 source.n66 5.81868
R310 source.n130 source.n100 5.81868
R311 source.n264 source.n263 5.53498
R312 source.n260 source.n259 5.04292
R313 source.n226 source.n225 5.04292
R314 source.n194 source.n193 5.04292
R315 source.n160 source.n159 5.04292
R316 source.n28 source.n27 5.04292
R317 source.n62 source.n61 5.04292
R318 source.n94 source.n93 5.04292
R319 source.n128 source.n127 5.04292
R320 source.n245 source.n241 4.38594
R321 source.n211 source.n207 4.38594
R322 source.n179 source.n175 4.38594
R323 source.n145 source.n141 4.38594
R324 source.n13 source.n9 4.38594
R325 source.n47 source.n43 4.38594
R326 source.n79 source.n75 4.38594
R327 source.n113 source.n109 4.38594
R328 source.n256 source.n234 4.26717
R329 source.n222 source.n200 4.26717
R330 source.n190 source.n168 4.26717
R331 source.n156 source.n134 4.26717
R332 source.n24 source.n2 4.26717
R333 source.n58 source.n36 4.26717
R334 source.n90 source.n68 4.26717
R335 source.n124 source.n102 4.26717
R336 source.n255 source.n236 3.49141
R337 source.n221 source.n202 3.49141
R338 source.n189 source.n170 3.49141
R339 source.n155 source.n136 3.49141
R340 source.n23 source.n4 3.49141
R341 source.n57 source.n38 3.49141
R342 source.n89 source.n70 3.49141
R343 source.n123 source.n104 3.49141
R344 source.n230 source.t7 3.3005
R345 source.n230 source.t11 3.3005
R346 source.n164 source.t2 3.3005
R347 source.n164 source.t15 3.3005
R348 source.n32 source.t6 3.3005
R349 source.n32 source.t4 3.3005
R350 source.n98 source.t13 3.3005
R351 source.n98 source.t14 3.3005
R352 source.n252 source.n251 2.71565
R353 source.n218 source.n217 2.71565
R354 source.n186 source.n185 2.71565
R355 source.n152 source.n151 2.71565
R356 source.n20 source.n19 2.71565
R357 source.n54 source.n53 2.71565
R358 source.n86 source.n85 2.71565
R359 source.n120 source.n119 2.71565
R360 source.n248 source.n238 1.93989
R361 source.n214 source.n204 1.93989
R362 source.n182 source.n172 1.93989
R363 source.n148 source.n138 1.93989
R364 source.n16 source.n6 1.93989
R365 source.n50 source.n40 1.93989
R366 source.n82 source.n72 1.93989
R367 source.n116 source.n106 1.93989
R368 source.n247 source.n240 1.16414
R369 source.n213 source.n206 1.16414
R370 source.n181 source.n174 1.16414
R371 source.n147 source.n140 1.16414
R372 source.n15 source.n8 1.16414
R373 source.n49 source.n42 1.16414
R374 source.n81 source.n74 1.16414
R375 source.n115 source.n108 1.16414
R376 source.n131 source.n99 0.543603
R377 source.n99 source.n97 0.543603
R378 source.n65 source.n33 0.543603
R379 source.n33 source.n31 0.543603
R380 source.n165 source.n163 0.543603
R381 source.n197 source.n165 0.543603
R382 source.n231 source.n229 0.543603
R383 source.n263 source.n231 0.543603
R384 source.n97 source.n65 0.470328
R385 source.n229 source.n197 0.470328
R386 source.n244 source.n243 0.388379
R387 source.n210 source.n209 0.388379
R388 source.n178 source.n177 0.388379
R389 source.n144 source.n143 0.388379
R390 source.n12 source.n11 0.388379
R391 source.n46 source.n45 0.388379
R392 source.n78 source.n77 0.388379
R393 source.n112 source.n111 0.388379
R394 source source.n264 0.188
R395 source.n246 source.n245 0.155672
R396 source.n246 source.n237 0.155672
R397 source.n253 source.n237 0.155672
R398 source.n254 source.n253 0.155672
R399 source.n254 source.n233 0.155672
R400 source.n261 source.n233 0.155672
R401 source.n212 source.n211 0.155672
R402 source.n212 source.n203 0.155672
R403 source.n219 source.n203 0.155672
R404 source.n220 source.n219 0.155672
R405 source.n220 source.n199 0.155672
R406 source.n227 source.n199 0.155672
R407 source.n180 source.n179 0.155672
R408 source.n180 source.n171 0.155672
R409 source.n187 source.n171 0.155672
R410 source.n188 source.n187 0.155672
R411 source.n188 source.n167 0.155672
R412 source.n195 source.n167 0.155672
R413 source.n146 source.n145 0.155672
R414 source.n146 source.n137 0.155672
R415 source.n153 source.n137 0.155672
R416 source.n154 source.n153 0.155672
R417 source.n154 source.n133 0.155672
R418 source.n161 source.n133 0.155672
R419 source.n29 source.n1 0.155672
R420 source.n22 source.n1 0.155672
R421 source.n22 source.n21 0.155672
R422 source.n21 source.n5 0.155672
R423 source.n14 source.n5 0.155672
R424 source.n14 source.n13 0.155672
R425 source.n63 source.n35 0.155672
R426 source.n56 source.n35 0.155672
R427 source.n56 source.n55 0.155672
R428 source.n55 source.n39 0.155672
R429 source.n48 source.n39 0.155672
R430 source.n48 source.n47 0.155672
R431 source.n95 source.n67 0.155672
R432 source.n88 source.n67 0.155672
R433 source.n88 source.n87 0.155672
R434 source.n87 source.n71 0.155672
R435 source.n80 source.n71 0.155672
R436 source.n80 source.n79 0.155672
R437 source.n129 source.n101 0.155672
R438 source.n122 source.n101 0.155672
R439 source.n122 source.n121 0.155672
R440 source.n121 source.n105 0.155672
R441 source.n114 source.n105 0.155672
R442 source.n114 source.n113 0.155672
R443 drain_right.n5 drain_right.n3 67.7338
R444 drain_right.n2 drain_right.n1 67.4069
R445 drain_right.n2 drain_right.n0 67.4069
R446 drain_right.n5 drain_right.n4 67.1908
R447 drain_right drain_right.n2 24.1693
R448 drain_right drain_right.n5 6.19632
R449 drain_right.n1 drain_right.t2 3.3005
R450 drain_right.n1 drain_right.t6 3.3005
R451 drain_right.n0 drain_right.t1 3.3005
R452 drain_right.n0 drain_right.t5 3.3005
R453 drain_right.n3 drain_right.t0 3.3005
R454 drain_right.n3 drain_right.t3 3.3005
R455 drain_right.n4 drain_right.t4 3.3005
R456 drain_right.n4 drain_right.t7 3.3005
R457 plus.n2 plus.t1 614.915
R458 plus.n7 plus.t7 614.915
R459 plus.n11 plus.t4 614.915
R460 plus.n16 plus.t2 614.915
R461 plus.n1 plus.t3 586.433
R462 plus.n6 plus.t6 586.433
R463 plus.n10 plus.t0 586.433
R464 plus.n15 plus.t5 586.433
R465 plus.n3 plus.n2 161.489
R466 plus.n12 plus.n11 161.489
R467 plus.n4 plus.n3 161.3
R468 plus.n5 plus.n0 161.3
R469 plus.n8 plus.n7 161.3
R470 plus.n13 plus.n12 161.3
R471 plus.n14 plus.n9 161.3
R472 plus.n17 plus.n16 161.3
R473 plus.n5 plus.n4 73.0308
R474 plus.n14 plus.n13 73.0308
R475 plus.n2 plus.n1 63.5369
R476 plus.n7 plus.n6 63.5369
R477 plus.n16 plus.n15 63.5369
R478 plus.n11 plus.n10 63.5369
R479 plus plus.n17 25.7907
R480 plus plus.n8 9.83383
R481 plus.n4 plus.n1 9.49444
R482 plus.n6 plus.n5 9.49444
R483 plus.n15 plus.n14 9.49444
R484 plus.n13 plus.n10 9.49444
R485 plus.n3 plus.n0 0.189894
R486 plus.n8 plus.n0 0.189894
R487 plus.n17 plus.n9 0.189894
R488 plus.n12 plus.n9 0.189894
R489 drain_left.n5 drain_left.n3 67.7339
R490 drain_left.n2 drain_left.n1 67.4069
R491 drain_left.n2 drain_left.n0 67.4069
R492 drain_left.n5 drain_left.n4 67.1907
R493 drain_left drain_left.n2 24.7225
R494 drain_left drain_left.n5 6.19632
R495 drain_left.n1 drain_left.t7 3.3005
R496 drain_left.n1 drain_left.t3 3.3005
R497 drain_left.n0 drain_left.t5 3.3005
R498 drain_left.n0 drain_left.t2 3.3005
R499 drain_left.n4 drain_left.t1 3.3005
R500 drain_left.n4 drain_left.t0 3.3005
R501 drain_left.n3 drain_left.t6 3.3005
R502 drain_left.n3 drain_left.t4 3.3005
C0 source plus 1.73406f
C1 source drain_right 9.19398f
C2 minus drain_left 0.170671f
C3 plus minus 3.72105f
C4 minus drain_right 1.85677f
C5 plus drain_left 1.98397f
C6 drain_right drain_left 0.630082f
C7 plus drain_right 0.280736f
C8 source minus 1.72004f
C9 source drain_left 9.19478f
C10 drain_right a_n1346_n2088# 4.02517f
C11 drain_left a_n1346_n2088# 4.19594f
C12 source a_n1346_n2088# 5.138415f
C13 minus a_n1346_n2088# 4.708669f
C14 plus a_n1346_n2088# 5.415934f
C15 drain_left.t5 a_n1346_n2088# 0.124838f
C16 drain_left.t2 a_n1346_n2088# 0.124838f
C17 drain_left.n0 a_n1346_n2088# 1.04209f
C18 drain_left.t7 a_n1346_n2088# 0.124838f
C19 drain_left.t3 a_n1346_n2088# 0.124838f
C20 drain_left.n1 a_n1346_n2088# 1.04209f
C21 drain_left.n2 a_n1346_n2088# 1.39354f
C22 drain_left.t6 a_n1346_n2088# 0.124838f
C23 drain_left.t4 a_n1346_n2088# 0.124838f
C24 drain_left.n3 a_n1346_n2088# 1.04369f
C25 drain_left.t1 a_n1346_n2088# 0.124838f
C26 drain_left.t0 a_n1346_n2088# 0.124838f
C27 drain_left.n4 a_n1346_n2088# 1.04115f
C28 drain_left.n5 a_n1346_n2088# 0.838925f
C29 plus.n0 a_n1346_n2088# 0.028203f
C30 plus.t6 a_n1346_n2088# 0.144638f
C31 plus.t3 a_n1346_n2088# 0.144638f
C32 plus.n1 a_n1346_n2088# 0.066391f
C33 plus.t1 a_n1346_n2088# 0.147709f
C34 plus.n2 a_n1346_n2088# 0.074886f
C35 plus.n3 a_n1346_n2088# 0.059672f
C36 plus.n4 a_n1346_n2088# 0.010486f
C37 plus.n5 a_n1346_n2088# 0.010486f
C38 plus.n6 a_n1346_n2088# 0.066391f
C39 plus.t7 a_n1346_n2088# 0.147709f
C40 plus.n7 a_n1346_n2088# 0.074849f
C41 plus.n8 a_n1346_n2088# 0.239073f
C42 plus.n9 a_n1346_n2088# 0.028203f
C43 plus.t2 a_n1346_n2088# 0.147709f
C44 plus.t5 a_n1346_n2088# 0.144638f
C45 plus.t0 a_n1346_n2088# 0.144638f
C46 plus.n10 a_n1346_n2088# 0.066391f
C47 plus.t4 a_n1346_n2088# 0.147709f
C48 plus.n11 a_n1346_n2088# 0.074886f
C49 plus.n12 a_n1346_n2088# 0.059672f
C50 plus.n13 a_n1346_n2088# 0.010486f
C51 plus.n14 a_n1346_n2088# 0.010486f
C52 plus.n15 a_n1346_n2088# 0.066391f
C53 plus.n16 a_n1346_n2088# 0.074849f
C54 plus.n17 a_n1346_n2088# 0.648686f
C55 drain_right.t1 a_n1346_n2088# 0.126252f
C56 drain_right.t5 a_n1346_n2088# 0.126252f
C57 drain_right.n0 a_n1346_n2088# 1.05389f
C58 drain_right.t2 a_n1346_n2088# 0.126252f
C59 drain_right.t6 a_n1346_n2088# 0.126252f
C60 drain_right.n1 a_n1346_n2088# 1.05389f
C61 drain_right.n2 a_n1346_n2088# 1.3548f
C62 drain_right.t0 a_n1346_n2088# 0.126252f
C63 drain_right.t3 a_n1346_n2088# 0.126252f
C64 drain_right.n3 a_n1346_n2088# 1.05551f
C65 drain_right.t4 a_n1346_n2088# 0.126252f
C66 drain_right.t7 a_n1346_n2088# 0.126252f
C67 drain_right.n4 a_n1346_n2088# 1.05295f
C68 drain_right.n5 a_n1346_n2088# 0.848424f
C69 source.n0 a_n1346_n2088# 0.02968f
C70 source.n1 a_n1346_n2088# 0.021115f
C71 source.n2 a_n1346_n2088# 0.011347f
C72 source.n3 a_n1346_n2088# 0.026819f
C73 source.n4 a_n1346_n2088# 0.012014f
C74 source.n5 a_n1346_n2088# 0.021115f
C75 source.n6 a_n1346_n2088# 0.011347f
C76 source.n7 a_n1346_n2088# 0.026819f
C77 source.n8 a_n1346_n2088# 0.012014f
C78 source.n9 a_n1346_n2088# 0.090359f
C79 source.t3 a_n1346_n2088# 0.043711f
C80 source.n10 a_n1346_n2088# 0.020114f
C81 source.n11 a_n1346_n2088# 0.015842f
C82 source.n12 a_n1346_n2088# 0.011347f
C83 source.n13 a_n1346_n2088# 0.502421f
C84 source.n14 a_n1346_n2088# 0.021115f
C85 source.n15 a_n1346_n2088# 0.011347f
C86 source.n16 a_n1346_n2088# 0.012014f
C87 source.n17 a_n1346_n2088# 0.026819f
C88 source.n18 a_n1346_n2088# 0.026819f
C89 source.n19 a_n1346_n2088# 0.012014f
C90 source.n20 a_n1346_n2088# 0.011347f
C91 source.n21 a_n1346_n2088# 0.021115f
C92 source.n22 a_n1346_n2088# 0.021115f
C93 source.n23 a_n1346_n2088# 0.011347f
C94 source.n24 a_n1346_n2088# 0.012014f
C95 source.n25 a_n1346_n2088# 0.026819f
C96 source.n26 a_n1346_n2088# 0.058059f
C97 source.n27 a_n1346_n2088# 0.012014f
C98 source.n28 a_n1346_n2088# 0.011347f
C99 source.n29 a_n1346_n2088# 0.048807f
C100 source.n30 a_n1346_n2088# 0.032486f
C101 source.n31 a_n1346_n2088# 0.511458f
C102 source.t6 a_n1346_n2088# 0.100116f
C103 source.t4 a_n1346_n2088# 0.100116f
C104 source.n32 a_n1346_n2088# 0.779714f
C105 source.n33 a_n1346_n2088# 0.271841f
C106 source.n34 a_n1346_n2088# 0.02968f
C107 source.n35 a_n1346_n2088# 0.021115f
C108 source.n36 a_n1346_n2088# 0.011347f
C109 source.n37 a_n1346_n2088# 0.026819f
C110 source.n38 a_n1346_n2088# 0.012014f
C111 source.n39 a_n1346_n2088# 0.021115f
C112 source.n40 a_n1346_n2088# 0.011347f
C113 source.n41 a_n1346_n2088# 0.026819f
C114 source.n42 a_n1346_n2088# 0.012014f
C115 source.n43 a_n1346_n2088# 0.090359f
C116 source.t0 a_n1346_n2088# 0.043711f
C117 source.n44 a_n1346_n2088# 0.020114f
C118 source.n45 a_n1346_n2088# 0.015842f
C119 source.n46 a_n1346_n2088# 0.011347f
C120 source.n47 a_n1346_n2088# 0.502421f
C121 source.n48 a_n1346_n2088# 0.021115f
C122 source.n49 a_n1346_n2088# 0.011347f
C123 source.n50 a_n1346_n2088# 0.012014f
C124 source.n51 a_n1346_n2088# 0.026819f
C125 source.n52 a_n1346_n2088# 0.026819f
C126 source.n53 a_n1346_n2088# 0.012014f
C127 source.n54 a_n1346_n2088# 0.011347f
C128 source.n55 a_n1346_n2088# 0.021115f
C129 source.n56 a_n1346_n2088# 0.021115f
C130 source.n57 a_n1346_n2088# 0.011347f
C131 source.n58 a_n1346_n2088# 0.012014f
C132 source.n59 a_n1346_n2088# 0.026819f
C133 source.n60 a_n1346_n2088# 0.058059f
C134 source.n61 a_n1346_n2088# 0.012014f
C135 source.n62 a_n1346_n2088# 0.011347f
C136 source.n63 a_n1346_n2088# 0.048807f
C137 source.n64 a_n1346_n2088# 0.032486f
C138 source.n65 a_n1346_n2088# 0.086953f
C139 source.n66 a_n1346_n2088# 0.02968f
C140 source.n67 a_n1346_n2088# 0.021115f
C141 source.n68 a_n1346_n2088# 0.011347f
C142 source.n69 a_n1346_n2088# 0.026819f
C143 source.n70 a_n1346_n2088# 0.012014f
C144 source.n71 a_n1346_n2088# 0.021115f
C145 source.n72 a_n1346_n2088# 0.011347f
C146 source.n73 a_n1346_n2088# 0.026819f
C147 source.n74 a_n1346_n2088# 0.012014f
C148 source.n75 a_n1346_n2088# 0.090359f
C149 source.t8 a_n1346_n2088# 0.043711f
C150 source.n76 a_n1346_n2088# 0.020114f
C151 source.n77 a_n1346_n2088# 0.015842f
C152 source.n78 a_n1346_n2088# 0.011347f
C153 source.n79 a_n1346_n2088# 0.502421f
C154 source.n80 a_n1346_n2088# 0.021115f
C155 source.n81 a_n1346_n2088# 0.011347f
C156 source.n82 a_n1346_n2088# 0.012014f
C157 source.n83 a_n1346_n2088# 0.026819f
C158 source.n84 a_n1346_n2088# 0.026819f
C159 source.n85 a_n1346_n2088# 0.012014f
C160 source.n86 a_n1346_n2088# 0.011347f
C161 source.n87 a_n1346_n2088# 0.021115f
C162 source.n88 a_n1346_n2088# 0.021115f
C163 source.n89 a_n1346_n2088# 0.011347f
C164 source.n90 a_n1346_n2088# 0.012014f
C165 source.n91 a_n1346_n2088# 0.026819f
C166 source.n92 a_n1346_n2088# 0.058059f
C167 source.n93 a_n1346_n2088# 0.012014f
C168 source.n94 a_n1346_n2088# 0.011347f
C169 source.n95 a_n1346_n2088# 0.048807f
C170 source.n96 a_n1346_n2088# 0.032486f
C171 source.n97 a_n1346_n2088# 0.086953f
C172 source.t13 a_n1346_n2088# 0.100116f
C173 source.t14 a_n1346_n2088# 0.100116f
C174 source.n98 a_n1346_n2088# 0.779714f
C175 source.n99 a_n1346_n2088# 0.271841f
C176 source.n100 a_n1346_n2088# 0.02968f
C177 source.n101 a_n1346_n2088# 0.021115f
C178 source.n102 a_n1346_n2088# 0.011347f
C179 source.n103 a_n1346_n2088# 0.026819f
C180 source.n104 a_n1346_n2088# 0.012014f
C181 source.n105 a_n1346_n2088# 0.021115f
C182 source.n106 a_n1346_n2088# 0.011347f
C183 source.n107 a_n1346_n2088# 0.026819f
C184 source.n108 a_n1346_n2088# 0.012014f
C185 source.n109 a_n1346_n2088# 0.090359f
C186 source.t10 a_n1346_n2088# 0.043711f
C187 source.n110 a_n1346_n2088# 0.020114f
C188 source.n111 a_n1346_n2088# 0.015842f
C189 source.n112 a_n1346_n2088# 0.011347f
C190 source.n113 a_n1346_n2088# 0.502421f
C191 source.n114 a_n1346_n2088# 0.021115f
C192 source.n115 a_n1346_n2088# 0.011347f
C193 source.n116 a_n1346_n2088# 0.012014f
C194 source.n117 a_n1346_n2088# 0.026819f
C195 source.n118 a_n1346_n2088# 0.026819f
C196 source.n119 a_n1346_n2088# 0.012014f
C197 source.n120 a_n1346_n2088# 0.011347f
C198 source.n121 a_n1346_n2088# 0.021115f
C199 source.n122 a_n1346_n2088# 0.021115f
C200 source.n123 a_n1346_n2088# 0.011347f
C201 source.n124 a_n1346_n2088# 0.012014f
C202 source.n125 a_n1346_n2088# 0.026819f
C203 source.n126 a_n1346_n2088# 0.058059f
C204 source.n127 a_n1346_n2088# 0.012014f
C205 source.n128 a_n1346_n2088# 0.011347f
C206 source.n129 a_n1346_n2088# 0.048807f
C207 source.n130 a_n1346_n2088# 0.032486f
C208 source.n131 a_n1346_n2088# 0.783297f
C209 source.n132 a_n1346_n2088# 0.02968f
C210 source.n133 a_n1346_n2088# 0.021115f
C211 source.n134 a_n1346_n2088# 0.011347f
C212 source.n135 a_n1346_n2088# 0.026819f
C213 source.n136 a_n1346_n2088# 0.012014f
C214 source.n137 a_n1346_n2088# 0.021115f
C215 source.n138 a_n1346_n2088# 0.011347f
C216 source.n139 a_n1346_n2088# 0.026819f
C217 source.n140 a_n1346_n2088# 0.012014f
C218 source.n141 a_n1346_n2088# 0.090359f
C219 source.t1 a_n1346_n2088# 0.043711f
C220 source.n142 a_n1346_n2088# 0.020114f
C221 source.n143 a_n1346_n2088# 0.015842f
C222 source.n144 a_n1346_n2088# 0.011347f
C223 source.n145 a_n1346_n2088# 0.502421f
C224 source.n146 a_n1346_n2088# 0.021115f
C225 source.n147 a_n1346_n2088# 0.011347f
C226 source.n148 a_n1346_n2088# 0.012014f
C227 source.n149 a_n1346_n2088# 0.026819f
C228 source.n150 a_n1346_n2088# 0.026819f
C229 source.n151 a_n1346_n2088# 0.012014f
C230 source.n152 a_n1346_n2088# 0.011347f
C231 source.n153 a_n1346_n2088# 0.021115f
C232 source.n154 a_n1346_n2088# 0.021115f
C233 source.n155 a_n1346_n2088# 0.011347f
C234 source.n156 a_n1346_n2088# 0.012014f
C235 source.n157 a_n1346_n2088# 0.026819f
C236 source.n158 a_n1346_n2088# 0.058059f
C237 source.n159 a_n1346_n2088# 0.012014f
C238 source.n160 a_n1346_n2088# 0.011347f
C239 source.n161 a_n1346_n2088# 0.048807f
C240 source.n162 a_n1346_n2088# 0.032486f
C241 source.n163 a_n1346_n2088# 0.783297f
C242 source.t2 a_n1346_n2088# 0.100116f
C243 source.t15 a_n1346_n2088# 0.100116f
C244 source.n164 a_n1346_n2088# 0.779709f
C245 source.n165 a_n1346_n2088# 0.271846f
C246 source.n166 a_n1346_n2088# 0.02968f
C247 source.n167 a_n1346_n2088# 0.021115f
C248 source.n168 a_n1346_n2088# 0.011347f
C249 source.n169 a_n1346_n2088# 0.026819f
C250 source.n170 a_n1346_n2088# 0.012014f
C251 source.n171 a_n1346_n2088# 0.021115f
C252 source.n172 a_n1346_n2088# 0.011347f
C253 source.n173 a_n1346_n2088# 0.026819f
C254 source.n174 a_n1346_n2088# 0.012014f
C255 source.n175 a_n1346_n2088# 0.090359f
C256 source.t5 a_n1346_n2088# 0.043711f
C257 source.n176 a_n1346_n2088# 0.020114f
C258 source.n177 a_n1346_n2088# 0.015842f
C259 source.n178 a_n1346_n2088# 0.011347f
C260 source.n179 a_n1346_n2088# 0.502421f
C261 source.n180 a_n1346_n2088# 0.021115f
C262 source.n181 a_n1346_n2088# 0.011347f
C263 source.n182 a_n1346_n2088# 0.012014f
C264 source.n183 a_n1346_n2088# 0.026819f
C265 source.n184 a_n1346_n2088# 0.026819f
C266 source.n185 a_n1346_n2088# 0.012014f
C267 source.n186 a_n1346_n2088# 0.011347f
C268 source.n187 a_n1346_n2088# 0.021115f
C269 source.n188 a_n1346_n2088# 0.021115f
C270 source.n189 a_n1346_n2088# 0.011347f
C271 source.n190 a_n1346_n2088# 0.012014f
C272 source.n191 a_n1346_n2088# 0.026819f
C273 source.n192 a_n1346_n2088# 0.058059f
C274 source.n193 a_n1346_n2088# 0.012014f
C275 source.n194 a_n1346_n2088# 0.011347f
C276 source.n195 a_n1346_n2088# 0.048807f
C277 source.n196 a_n1346_n2088# 0.032486f
C278 source.n197 a_n1346_n2088# 0.086953f
C279 source.n198 a_n1346_n2088# 0.02968f
C280 source.n199 a_n1346_n2088# 0.021115f
C281 source.n200 a_n1346_n2088# 0.011347f
C282 source.n201 a_n1346_n2088# 0.026819f
C283 source.n202 a_n1346_n2088# 0.012014f
C284 source.n203 a_n1346_n2088# 0.021115f
C285 source.n204 a_n1346_n2088# 0.011347f
C286 source.n205 a_n1346_n2088# 0.026819f
C287 source.n206 a_n1346_n2088# 0.012014f
C288 source.n207 a_n1346_n2088# 0.090359f
C289 source.t9 a_n1346_n2088# 0.043711f
C290 source.n208 a_n1346_n2088# 0.020114f
C291 source.n209 a_n1346_n2088# 0.015842f
C292 source.n210 a_n1346_n2088# 0.011347f
C293 source.n211 a_n1346_n2088# 0.502421f
C294 source.n212 a_n1346_n2088# 0.021115f
C295 source.n213 a_n1346_n2088# 0.011347f
C296 source.n214 a_n1346_n2088# 0.012014f
C297 source.n215 a_n1346_n2088# 0.026819f
C298 source.n216 a_n1346_n2088# 0.026819f
C299 source.n217 a_n1346_n2088# 0.012014f
C300 source.n218 a_n1346_n2088# 0.011347f
C301 source.n219 a_n1346_n2088# 0.021115f
C302 source.n220 a_n1346_n2088# 0.021115f
C303 source.n221 a_n1346_n2088# 0.011347f
C304 source.n222 a_n1346_n2088# 0.012014f
C305 source.n223 a_n1346_n2088# 0.026819f
C306 source.n224 a_n1346_n2088# 0.058059f
C307 source.n225 a_n1346_n2088# 0.012014f
C308 source.n226 a_n1346_n2088# 0.011347f
C309 source.n227 a_n1346_n2088# 0.048807f
C310 source.n228 a_n1346_n2088# 0.032486f
C311 source.n229 a_n1346_n2088# 0.086953f
C312 source.t7 a_n1346_n2088# 0.100116f
C313 source.t11 a_n1346_n2088# 0.100116f
C314 source.n230 a_n1346_n2088# 0.779709f
C315 source.n231 a_n1346_n2088# 0.271846f
C316 source.n232 a_n1346_n2088# 0.02968f
C317 source.n233 a_n1346_n2088# 0.021115f
C318 source.n234 a_n1346_n2088# 0.011347f
C319 source.n235 a_n1346_n2088# 0.026819f
C320 source.n236 a_n1346_n2088# 0.012014f
C321 source.n237 a_n1346_n2088# 0.021115f
C322 source.n238 a_n1346_n2088# 0.011347f
C323 source.n239 a_n1346_n2088# 0.026819f
C324 source.n240 a_n1346_n2088# 0.012014f
C325 source.n241 a_n1346_n2088# 0.090359f
C326 source.t12 a_n1346_n2088# 0.043711f
C327 source.n242 a_n1346_n2088# 0.020114f
C328 source.n243 a_n1346_n2088# 0.015842f
C329 source.n244 a_n1346_n2088# 0.011347f
C330 source.n245 a_n1346_n2088# 0.502421f
C331 source.n246 a_n1346_n2088# 0.021115f
C332 source.n247 a_n1346_n2088# 0.011347f
C333 source.n248 a_n1346_n2088# 0.012014f
C334 source.n249 a_n1346_n2088# 0.026819f
C335 source.n250 a_n1346_n2088# 0.026819f
C336 source.n251 a_n1346_n2088# 0.012014f
C337 source.n252 a_n1346_n2088# 0.011347f
C338 source.n253 a_n1346_n2088# 0.021115f
C339 source.n254 a_n1346_n2088# 0.021115f
C340 source.n255 a_n1346_n2088# 0.011347f
C341 source.n256 a_n1346_n2088# 0.012014f
C342 source.n257 a_n1346_n2088# 0.026819f
C343 source.n258 a_n1346_n2088# 0.058059f
C344 source.n259 a_n1346_n2088# 0.012014f
C345 source.n260 a_n1346_n2088# 0.011347f
C346 source.n261 a_n1346_n2088# 0.048807f
C347 source.n262 a_n1346_n2088# 0.032486f
C348 source.n263 a_n1346_n2088# 0.206149f
C349 source.n264 a_n1346_n2088# 0.864006f
C350 minus.n0 a_n1346_n2088# 0.027775f
C351 minus.t3 a_n1346_n2088# 0.145467f
C352 minus.t0 a_n1346_n2088# 0.142442f
C353 minus.t7 a_n1346_n2088# 0.142442f
C354 minus.n1 a_n1346_n2088# 0.065383f
C355 minus.t4 a_n1346_n2088# 0.145467f
C356 minus.n2 a_n1346_n2088# 0.073749f
C357 minus.n3 a_n1346_n2088# 0.058766f
C358 minus.n4 a_n1346_n2088# 0.010327f
C359 minus.n5 a_n1346_n2088# 0.010327f
C360 minus.n6 a_n1346_n2088# 0.065383f
C361 minus.n7 a_n1346_n2088# 0.073713f
C362 minus.n8 a_n1346_n2088# 0.706639f
C363 minus.n9 a_n1346_n2088# 0.027775f
C364 minus.t5 a_n1346_n2088# 0.142442f
C365 minus.t2 a_n1346_n2088# 0.142442f
C366 minus.n10 a_n1346_n2088# 0.065383f
C367 minus.t6 a_n1346_n2088# 0.145467f
C368 minus.n11 a_n1346_n2088# 0.073749f
C369 minus.n12 a_n1346_n2088# 0.058766f
C370 minus.n13 a_n1346_n2088# 0.010327f
C371 minus.n14 a_n1346_n2088# 0.010327f
C372 minus.n15 a_n1346_n2088# 0.065383f
C373 minus.t1 a_n1346_n2088# 0.145467f
C374 minus.n16 a_n1346_n2088# 0.073713f
C375 minus.n17 a_n1346_n2088# 0.179133f
C376 minus.n18 a_n1346_n2088# 0.873506f
.ends

