* NGSPICE file created from diffpair670.ext - technology: sky130A

.subckt diffpair670 minus drain_right drain_left source plus
X0 drain_right minus source a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.3
X1 a_n968_n5892# a_n968_n5892# a_n968_n5892# a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X2 drain_left plus source a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.3
X3 a_n968_n5892# a_n968_n5892# a_n968_n5892# a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X4 drain_right minus source a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.3
X5 drain_left plus source a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.3
X6 a_n968_n5892# a_n968_n5892# a_n968_n5892# a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X7 a_n968_n5892# a_n968_n5892# a_n968_n5892# a_n968_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
.ends

