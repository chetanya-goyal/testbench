* NGSPICE file created from diffpair276.ext - technology: sky130A

.subckt diffpair276 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t20 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X1 drain_right.t12 minus.t1 source.t18 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 source.t14 minus.t2 drain_right.t11 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X3 drain_right.t10 minus.t3 source.t15 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X4 source.t7 plus.t0 drain_left.t13 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X5 drain_left.t12 plus.t1 source.t11 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X6 source.t5 plus.t2 drain_left.t11 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 source.t6 plus.t3 drain_left.t10 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X8 drain_right.t9 minus.t4 source.t16 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X9 source.t23 minus.t5 drain_right.t8 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 source.t24 minus.t6 drain_right.t7 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X11 a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X12 a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X13 source.t21 minus.t7 drain_right.t6 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 drain_left.t9 plus.t4 source.t10 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X15 source.t0 plus.t5 drain_left.t8 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X16 drain_left.t7 plus.t6 source.t13 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X17 drain_left.t6 plus.t7 source.t3 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X18 source.t27 minus.t8 drain_right.t5 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X19 drain_right.t4 minus.t9 source.t22 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X20 source.t1 plus.t8 drain_left.t5 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X21 a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X22 drain_right.t3 minus.t10 source.t26 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X23 drain_right.t2 minus.t11 source.t17 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X24 drain_left.t4 plus.t9 source.t2 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X25 drain_right.t1 minus.t12 source.t25 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X26 drain_left.t3 plus.t10 source.t4 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X27 drain_left.t2 plus.t11 source.t8 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X28 a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X29 source.t19 minus.t13 drain_right.t0 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X30 drain_left.t1 plus.t12 source.t12 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X31 source.t9 plus.t13 drain_left.t0 a_n1724_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n15 minus.t4 643.398
R1 minus.n3 minus.t9 643.398
R2 minus.n32 minus.t0 643.398
R3 minus.n20 minus.t11 643.398
R4 minus.n1 minus.t8 586.433
R5 minus.n14 minus.t2 586.433
R6 minus.n12 minus.t12 586.433
R7 minus.n6 minus.t3 586.433
R8 minus.n4 minus.t13 586.433
R9 minus.n18 minus.t5 586.433
R10 minus.n31 minus.t7 586.433
R11 minus.n29 minus.t1 586.433
R12 minus.n23 minus.t10 586.433
R13 minus.n21 minus.t6 586.433
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n15 minus.n14 35.055
R41 minus.n4 minus.n3 35.055
R42 minus.n21 minus.n20 35.055
R43 minus.n32 minus.n31 35.055
R44 minus.n34 minus.n16 31.1425
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 source.n146 source.n120 289.615
R62 source.n108 source.n82 289.615
R63 source.n26 source.n0 289.615
R64 source.n64 source.n38 289.615
R65 source.n131 source.n130 185
R66 source.n128 source.n127 185
R67 source.n137 source.n136 185
R68 source.n139 source.n138 185
R69 source.n124 source.n123 185
R70 source.n145 source.n144 185
R71 source.n147 source.n146 185
R72 source.n93 source.n92 185
R73 source.n90 source.n89 185
R74 source.n99 source.n98 185
R75 source.n101 source.n100 185
R76 source.n86 source.n85 185
R77 source.n107 source.n106 185
R78 source.n109 source.n108 185
R79 source.n27 source.n26 185
R80 source.n25 source.n24 185
R81 source.n4 source.n3 185
R82 source.n19 source.n18 185
R83 source.n17 source.n16 185
R84 source.n8 source.n7 185
R85 source.n11 source.n10 185
R86 source.n65 source.n64 185
R87 source.n63 source.n62 185
R88 source.n42 source.n41 185
R89 source.n57 source.n56 185
R90 source.n55 source.n54 185
R91 source.n46 source.n45 185
R92 source.n49 source.n48 185
R93 source.t20 source.n129 147.661
R94 source.t13 source.n91 147.661
R95 source.t12 source.n9 147.661
R96 source.t22 source.n47 147.661
R97 source.n130 source.n127 104.615
R98 source.n137 source.n127 104.615
R99 source.n138 source.n137 104.615
R100 source.n138 source.n123 104.615
R101 source.n145 source.n123 104.615
R102 source.n146 source.n145 104.615
R103 source.n92 source.n89 104.615
R104 source.n99 source.n89 104.615
R105 source.n100 source.n99 104.615
R106 source.n100 source.n85 104.615
R107 source.n107 source.n85 104.615
R108 source.n108 source.n107 104.615
R109 source.n26 source.n25 104.615
R110 source.n25 source.n3 104.615
R111 source.n18 source.n3 104.615
R112 source.n18 source.n17 104.615
R113 source.n17 source.n7 104.615
R114 source.n10 source.n7 104.615
R115 source.n64 source.n63 104.615
R116 source.n63 source.n41 104.615
R117 source.n56 source.n41 104.615
R118 source.n56 source.n55 104.615
R119 source.n55 source.n45 104.615
R120 source.n48 source.n45 104.615
R121 source.n130 source.t20 52.3082
R122 source.n92 source.t13 52.3082
R123 source.n10 source.t12 52.3082
R124 source.n48 source.t22 52.3082
R125 source.n33 source.n32 50.512
R126 source.n35 source.n34 50.512
R127 source.n37 source.n36 50.512
R128 source.n71 source.n70 50.512
R129 source.n73 source.n72 50.512
R130 source.n75 source.n74 50.512
R131 source.n119 source.n118 50.5119
R132 source.n117 source.n116 50.5119
R133 source.n115 source.n114 50.5119
R134 source.n81 source.n80 50.5119
R135 source.n79 source.n78 50.5119
R136 source.n77 source.n76 50.5119
R137 source.n151 source.n150 32.1853
R138 source.n113 source.n112 32.1853
R139 source.n31 source.n30 32.1853
R140 source.n69 source.n68 32.1853
R141 source.n77 source.n75 17.8285
R142 source.n131 source.n129 15.6674
R143 source.n93 source.n91 15.6674
R144 source.n11 source.n9 15.6674
R145 source.n49 source.n47 15.6674
R146 source.n132 source.n128 12.8005
R147 source.n94 source.n90 12.8005
R148 source.n12 source.n8 12.8005
R149 source.n50 source.n46 12.8005
R150 source.n136 source.n135 12.0247
R151 source.n98 source.n97 12.0247
R152 source.n16 source.n15 12.0247
R153 source.n54 source.n53 12.0247
R154 source.n152 source.n31 11.7509
R155 source.n139 source.n126 11.249
R156 source.n101 source.n88 11.249
R157 source.n19 source.n6 11.249
R158 source.n57 source.n44 11.249
R159 source.n140 source.n124 10.4732
R160 source.n102 source.n86 10.4732
R161 source.n20 source.n4 10.4732
R162 source.n58 source.n42 10.4732
R163 source.n144 source.n143 9.69747
R164 source.n106 source.n105 9.69747
R165 source.n24 source.n23 9.69747
R166 source.n62 source.n61 9.69747
R167 source.n150 source.n149 9.45567
R168 source.n112 source.n111 9.45567
R169 source.n30 source.n29 9.45567
R170 source.n68 source.n67 9.45567
R171 source.n149 source.n148 9.3005
R172 source.n122 source.n121 9.3005
R173 source.n143 source.n142 9.3005
R174 source.n141 source.n140 9.3005
R175 source.n126 source.n125 9.3005
R176 source.n135 source.n134 9.3005
R177 source.n133 source.n132 9.3005
R178 source.n111 source.n110 9.3005
R179 source.n84 source.n83 9.3005
R180 source.n105 source.n104 9.3005
R181 source.n103 source.n102 9.3005
R182 source.n88 source.n87 9.3005
R183 source.n97 source.n96 9.3005
R184 source.n95 source.n94 9.3005
R185 source.n29 source.n28 9.3005
R186 source.n2 source.n1 9.3005
R187 source.n23 source.n22 9.3005
R188 source.n21 source.n20 9.3005
R189 source.n6 source.n5 9.3005
R190 source.n15 source.n14 9.3005
R191 source.n13 source.n12 9.3005
R192 source.n67 source.n66 9.3005
R193 source.n40 source.n39 9.3005
R194 source.n61 source.n60 9.3005
R195 source.n59 source.n58 9.3005
R196 source.n44 source.n43 9.3005
R197 source.n53 source.n52 9.3005
R198 source.n51 source.n50 9.3005
R199 source.n147 source.n122 8.92171
R200 source.n109 source.n84 8.92171
R201 source.n27 source.n2 8.92171
R202 source.n65 source.n40 8.92171
R203 source.n148 source.n120 8.14595
R204 source.n110 source.n82 8.14595
R205 source.n28 source.n0 8.14595
R206 source.n66 source.n38 8.14595
R207 source.n150 source.n120 5.81868
R208 source.n112 source.n82 5.81868
R209 source.n30 source.n0 5.81868
R210 source.n68 source.n38 5.81868
R211 source.n152 source.n151 5.53498
R212 source.n148 source.n147 5.04292
R213 source.n110 source.n109 5.04292
R214 source.n28 source.n27 5.04292
R215 source.n66 source.n65 5.04292
R216 source.n133 source.n129 4.38594
R217 source.n95 source.n91 4.38594
R218 source.n13 source.n9 4.38594
R219 source.n51 source.n47 4.38594
R220 source.n144 source.n122 4.26717
R221 source.n106 source.n84 4.26717
R222 source.n24 source.n2 4.26717
R223 source.n62 source.n40 4.26717
R224 source.n143 source.n124 3.49141
R225 source.n105 source.n86 3.49141
R226 source.n23 source.n4 3.49141
R227 source.n61 source.n42 3.49141
R228 source.n118 source.t18 3.3005
R229 source.n118 source.t21 3.3005
R230 source.n116 source.t26 3.3005
R231 source.n116 source.t23 3.3005
R232 source.n114 source.t17 3.3005
R233 source.n114 source.t24 3.3005
R234 source.n80 source.t3 3.3005
R235 source.n80 source.t7 3.3005
R236 source.n78 source.t4 3.3005
R237 source.n78 source.t5 3.3005
R238 source.n76 source.t8 3.3005
R239 source.n76 source.t6 3.3005
R240 source.n32 source.t10 3.3005
R241 source.n32 source.t1 3.3005
R242 source.n34 source.t2 3.3005
R243 source.n34 source.t9 3.3005
R244 source.n36 source.t11 3.3005
R245 source.n36 source.t0 3.3005
R246 source.n70 source.t15 3.3005
R247 source.n70 source.t19 3.3005
R248 source.n72 source.t25 3.3005
R249 source.n72 source.t27 3.3005
R250 source.n74 source.t16 3.3005
R251 source.n74 source.t14 3.3005
R252 source.n140 source.n139 2.71565
R253 source.n102 source.n101 2.71565
R254 source.n20 source.n19 2.71565
R255 source.n58 source.n57 2.71565
R256 source.n136 source.n126 1.93989
R257 source.n98 source.n88 1.93989
R258 source.n16 source.n6 1.93989
R259 source.n54 source.n44 1.93989
R260 source.n135 source.n128 1.16414
R261 source.n97 source.n90 1.16414
R262 source.n15 source.n8 1.16414
R263 source.n53 source.n46 1.16414
R264 source.n69 source.n37 0.741879
R265 source.n115 source.n113 0.741879
R266 source.n75 source.n73 0.543603
R267 source.n73 source.n71 0.543603
R268 source.n71 source.n69 0.543603
R269 source.n37 source.n35 0.543603
R270 source.n35 source.n33 0.543603
R271 source.n33 source.n31 0.543603
R272 source.n79 source.n77 0.543603
R273 source.n81 source.n79 0.543603
R274 source.n113 source.n81 0.543603
R275 source.n117 source.n115 0.543603
R276 source.n119 source.n117 0.543603
R277 source.n151 source.n119 0.543603
R278 source.n132 source.n131 0.388379
R279 source.n94 source.n93 0.388379
R280 source.n12 source.n11 0.388379
R281 source.n50 source.n49 0.388379
R282 source source.n152 0.188
R283 source.n134 source.n133 0.155672
R284 source.n134 source.n125 0.155672
R285 source.n141 source.n125 0.155672
R286 source.n142 source.n141 0.155672
R287 source.n142 source.n121 0.155672
R288 source.n149 source.n121 0.155672
R289 source.n96 source.n95 0.155672
R290 source.n96 source.n87 0.155672
R291 source.n103 source.n87 0.155672
R292 source.n104 source.n103 0.155672
R293 source.n104 source.n83 0.155672
R294 source.n111 source.n83 0.155672
R295 source.n29 source.n1 0.155672
R296 source.n22 source.n1 0.155672
R297 source.n22 source.n21 0.155672
R298 source.n21 source.n5 0.155672
R299 source.n14 source.n5 0.155672
R300 source.n14 source.n13 0.155672
R301 source.n67 source.n39 0.155672
R302 source.n60 source.n39 0.155672
R303 source.n60 source.n59 0.155672
R304 source.n59 source.n43 0.155672
R305 source.n52 source.n43 0.155672
R306 source.n52 source.n51 0.155672
R307 drain_right.n26 drain_right.n0 289.615
R308 drain_right.n68 drain_right.n42 289.615
R309 drain_right.n11 drain_right.n10 185
R310 drain_right.n8 drain_right.n7 185
R311 drain_right.n17 drain_right.n16 185
R312 drain_right.n19 drain_right.n18 185
R313 drain_right.n4 drain_right.n3 185
R314 drain_right.n25 drain_right.n24 185
R315 drain_right.n27 drain_right.n26 185
R316 drain_right.n69 drain_right.n68 185
R317 drain_right.n67 drain_right.n66 185
R318 drain_right.n46 drain_right.n45 185
R319 drain_right.n61 drain_right.n60 185
R320 drain_right.n59 drain_right.n58 185
R321 drain_right.n50 drain_right.n49 185
R322 drain_right.n53 drain_right.n52 185
R323 drain_right.t2 drain_right.n9 147.661
R324 drain_right.t9 drain_right.n51 147.661
R325 drain_right.n10 drain_right.n7 104.615
R326 drain_right.n17 drain_right.n7 104.615
R327 drain_right.n18 drain_right.n17 104.615
R328 drain_right.n18 drain_right.n3 104.615
R329 drain_right.n25 drain_right.n3 104.615
R330 drain_right.n26 drain_right.n25 104.615
R331 drain_right.n68 drain_right.n67 104.615
R332 drain_right.n67 drain_right.n45 104.615
R333 drain_right.n60 drain_right.n45 104.615
R334 drain_right.n60 drain_right.n59 104.615
R335 drain_right.n59 drain_right.n49 104.615
R336 drain_right.n52 drain_right.n49 104.615
R337 drain_right.n35 drain_right.n33 67.7338
R338 drain_right.n39 drain_right.n37 67.7338
R339 drain_right.n39 drain_right.n38 67.1908
R340 drain_right.n41 drain_right.n40 67.1908
R341 drain_right.n35 drain_right.n34 67.1907
R342 drain_right.n32 drain_right.n31 67.1907
R343 drain_right.n10 drain_right.t2 52.3082
R344 drain_right.n52 drain_right.t9 52.3082
R345 drain_right.n32 drain_right.n30 49.4072
R346 drain_right.n73 drain_right.n72 48.8641
R347 drain_right drain_right.n36 25.3912
R348 drain_right.n11 drain_right.n9 15.6674
R349 drain_right.n53 drain_right.n51 15.6674
R350 drain_right.n12 drain_right.n8 12.8005
R351 drain_right.n54 drain_right.n50 12.8005
R352 drain_right.n16 drain_right.n15 12.0247
R353 drain_right.n58 drain_right.n57 12.0247
R354 drain_right.n19 drain_right.n6 11.249
R355 drain_right.n61 drain_right.n48 11.249
R356 drain_right.n20 drain_right.n4 10.4732
R357 drain_right.n62 drain_right.n46 10.4732
R358 drain_right.n24 drain_right.n23 9.69747
R359 drain_right.n66 drain_right.n65 9.69747
R360 drain_right.n30 drain_right.n29 9.45567
R361 drain_right.n72 drain_right.n71 9.45567
R362 drain_right.n29 drain_right.n28 9.3005
R363 drain_right.n2 drain_right.n1 9.3005
R364 drain_right.n23 drain_right.n22 9.3005
R365 drain_right.n21 drain_right.n20 9.3005
R366 drain_right.n6 drain_right.n5 9.3005
R367 drain_right.n15 drain_right.n14 9.3005
R368 drain_right.n13 drain_right.n12 9.3005
R369 drain_right.n71 drain_right.n70 9.3005
R370 drain_right.n44 drain_right.n43 9.3005
R371 drain_right.n65 drain_right.n64 9.3005
R372 drain_right.n63 drain_right.n62 9.3005
R373 drain_right.n48 drain_right.n47 9.3005
R374 drain_right.n57 drain_right.n56 9.3005
R375 drain_right.n55 drain_right.n54 9.3005
R376 drain_right.n27 drain_right.n2 8.92171
R377 drain_right.n69 drain_right.n44 8.92171
R378 drain_right.n28 drain_right.n0 8.14595
R379 drain_right.n70 drain_right.n42 8.14595
R380 drain_right drain_right.n73 5.92477
R381 drain_right.n30 drain_right.n0 5.81868
R382 drain_right.n72 drain_right.n42 5.81868
R383 drain_right.n28 drain_right.n27 5.04292
R384 drain_right.n70 drain_right.n69 5.04292
R385 drain_right.n13 drain_right.n9 4.38594
R386 drain_right.n55 drain_right.n51 4.38594
R387 drain_right.n24 drain_right.n2 4.26717
R388 drain_right.n66 drain_right.n44 4.26717
R389 drain_right.n23 drain_right.n4 3.49141
R390 drain_right.n65 drain_right.n46 3.49141
R391 drain_right.n33 drain_right.t6 3.3005
R392 drain_right.n33 drain_right.t13 3.3005
R393 drain_right.n34 drain_right.t8 3.3005
R394 drain_right.n34 drain_right.t12 3.3005
R395 drain_right.n31 drain_right.t7 3.3005
R396 drain_right.n31 drain_right.t3 3.3005
R397 drain_right.n37 drain_right.t0 3.3005
R398 drain_right.n37 drain_right.t4 3.3005
R399 drain_right.n38 drain_right.t5 3.3005
R400 drain_right.n38 drain_right.t10 3.3005
R401 drain_right.n40 drain_right.t11 3.3005
R402 drain_right.n40 drain_right.t1 3.3005
R403 drain_right.n20 drain_right.n19 2.71565
R404 drain_right.n62 drain_right.n61 2.71565
R405 drain_right.n16 drain_right.n6 1.93989
R406 drain_right.n58 drain_right.n48 1.93989
R407 drain_right.n15 drain_right.n8 1.16414
R408 drain_right.n57 drain_right.n50 1.16414
R409 drain_right.n73 drain_right.n41 0.543603
R410 drain_right.n41 drain_right.n39 0.543603
R411 drain_right.n12 drain_right.n11 0.388379
R412 drain_right.n54 drain_right.n53 0.388379
R413 drain_right.n36 drain_right.n32 0.352482
R414 drain_right.n14 drain_right.n13 0.155672
R415 drain_right.n14 drain_right.n5 0.155672
R416 drain_right.n21 drain_right.n5 0.155672
R417 drain_right.n22 drain_right.n21 0.155672
R418 drain_right.n22 drain_right.n1 0.155672
R419 drain_right.n29 drain_right.n1 0.155672
R420 drain_right.n71 drain_right.n43 0.155672
R421 drain_right.n64 drain_right.n43 0.155672
R422 drain_right.n64 drain_right.n63 0.155672
R423 drain_right.n63 drain_right.n47 0.155672
R424 drain_right.n56 drain_right.n47 0.155672
R425 drain_right.n56 drain_right.n55 0.155672
R426 drain_right.n36 drain_right.n35 0.0809298
R427 plus.n3 plus.t1 643.398
R428 plus.n15 plus.t12 643.398
R429 plus.n20 plus.t6 643.398
R430 plus.n32 plus.t11 643.398
R431 plus.n1 plus.t13 586.433
R432 plus.n4 plus.t5 586.433
R433 plus.n6 plus.t9 586.433
R434 plus.n12 plus.t4 586.433
R435 plus.n14 plus.t8 586.433
R436 plus.n18 plus.t2 586.433
R437 plus.n21 plus.t0 586.433
R438 plus.n23 plus.t7 586.433
R439 plus.n29 plus.t10 586.433
R440 plus.n31 plus.t3 586.433
R441 plus.n3 plus.n2 161.489
R442 plus.n20 plus.n19 161.489
R443 plus.n5 plus.n2 161.3
R444 plus.n8 plus.n7 161.3
R445 plus.n9 plus.n1 161.3
R446 plus.n11 plus.n10 161.3
R447 plus.n13 plus.n0 161.3
R448 plus.n16 plus.n15 161.3
R449 plus.n22 plus.n19 161.3
R450 plus.n25 plus.n24 161.3
R451 plus.n26 plus.n18 161.3
R452 plus.n28 plus.n27 161.3
R453 plus.n30 plus.n17 161.3
R454 plus.n33 plus.n32 161.3
R455 plus.n7 plus.n1 73.0308
R456 plus.n11 plus.n1 73.0308
R457 plus.n28 plus.n18 73.0308
R458 plus.n24 plus.n18 73.0308
R459 plus.n6 plus.n5 54.0429
R460 plus.n13 plus.n12 54.0429
R461 plus.n30 plus.n29 54.0429
R462 plus.n23 plus.n22 54.0429
R463 plus.n5 plus.n4 37.9763
R464 plus.n14 plus.n13 37.9763
R465 plus.n31 plus.n30 37.9763
R466 plus.n22 plus.n21 37.9763
R467 plus.n4 plus.n3 35.055
R468 plus.n15 plus.n14 35.055
R469 plus.n32 plus.n31 35.055
R470 plus.n21 plus.n20 35.055
R471 plus plus.n33 27.2964
R472 plus.n7 plus.n6 18.9884
R473 plus.n12 plus.n11 18.9884
R474 plus.n29 plus.n28 18.9884
R475 plus.n24 plus.n23 18.9884
R476 plus plus.n16 9.9077
R477 plus.n8 plus.n2 0.189894
R478 plus.n9 plus.n8 0.189894
R479 plus.n10 plus.n9 0.189894
R480 plus.n10 plus.n0 0.189894
R481 plus.n16 plus.n0 0.189894
R482 plus.n33 plus.n17 0.189894
R483 plus.n27 plus.n17 0.189894
R484 plus.n27 plus.n26 0.189894
R485 plus.n26 plus.n25 0.189894
R486 plus.n25 plus.n19 0.189894
R487 drain_left.n26 drain_left.n0 289.615
R488 drain_left.n63 drain_left.n37 289.615
R489 drain_left.n11 drain_left.n10 185
R490 drain_left.n8 drain_left.n7 185
R491 drain_left.n17 drain_left.n16 185
R492 drain_left.n19 drain_left.n18 185
R493 drain_left.n4 drain_left.n3 185
R494 drain_left.n25 drain_left.n24 185
R495 drain_left.n27 drain_left.n26 185
R496 drain_left.n64 drain_left.n63 185
R497 drain_left.n62 drain_left.n61 185
R498 drain_left.n41 drain_left.n40 185
R499 drain_left.n56 drain_left.n55 185
R500 drain_left.n54 drain_left.n53 185
R501 drain_left.n45 drain_left.n44 185
R502 drain_left.n48 drain_left.n47 185
R503 drain_left.t2 drain_left.n9 147.661
R504 drain_left.t12 drain_left.n46 147.661
R505 drain_left.n10 drain_left.n7 104.615
R506 drain_left.n17 drain_left.n7 104.615
R507 drain_left.n18 drain_left.n17 104.615
R508 drain_left.n18 drain_left.n3 104.615
R509 drain_left.n25 drain_left.n3 104.615
R510 drain_left.n26 drain_left.n25 104.615
R511 drain_left.n63 drain_left.n62 104.615
R512 drain_left.n62 drain_left.n40 104.615
R513 drain_left.n55 drain_left.n40 104.615
R514 drain_left.n55 drain_left.n54 104.615
R515 drain_left.n54 drain_left.n44 104.615
R516 drain_left.n47 drain_left.n44 104.615
R517 drain_left.n35 drain_left.n33 67.7338
R518 drain_left.n71 drain_left.n70 67.1908
R519 drain_left.n69 drain_left.n68 67.1908
R520 drain_left.n73 drain_left.n72 67.1907
R521 drain_left.n35 drain_left.n34 67.1907
R522 drain_left.n32 drain_left.n31 67.1907
R523 drain_left.n10 drain_left.t2 52.3082
R524 drain_left.n47 drain_left.t12 52.3082
R525 drain_left.n32 drain_left.n30 49.4072
R526 drain_left.n69 drain_left.n67 49.4072
R527 drain_left drain_left.n36 25.9445
R528 drain_left.n11 drain_left.n9 15.6674
R529 drain_left.n48 drain_left.n46 15.6674
R530 drain_left.n12 drain_left.n8 12.8005
R531 drain_left.n49 drain_left.n45 12.8005
R532 drain_left.n16 drain_left.n15 12.0247
R533 drain_left.n53 drain_left.n52 12.0247
R534 drain_left.n19 drain_left.n6 11.249
R535 drain_left.n56 drain_left.n43 11.249
R536 drain_left.n20 drain_left.n4 10.4732
R537 drain_left.n57 drain_left.n41 10.4732
R538 drain_left.n24 drain_left.n23 9.69747
R539 drain_left.n61 drain_left.n60 9.69747
R540 drain_left.n30 drain_left.n29 9.45567
R541 drain_left.n67 drain_left.n66 9.45567
R542 drain_left.n29 drain_left.n28 9.3005
R543 drain_left.n2 drain_left.n1 9.3005
R544 drain_left.n23 drain_left.n22 9.3005
R545 drain_left.n21 drain_left.n20 9.3005
R546 drain_left.n6 drain_left.n5 9.3005
R547 drain_left.n15 drain_left.n14 9.3005
R548 drain_left.n13 drain_left.n12 9.3005
R549 drain_left.n66 drain_left.n65 9.3005
R550 drain_left.n39 drain_left.n38 9.3005
R551 drain_left.n60 drain_left.n59 9.3005
R552 drain_left.n58 drain_left.n57 9.3005
R553 drain_left.n43 drain_left.n42 9.3005
R554 drain_left.n52 drain_left.n51 9.3005
R555 drain_left.n50 drain_left.n49 9.3005
R556 drain_left.n27 drain_left.n2 8.92171
R557 drain_left.n64 drain_left.n39 8.92171
R558 drain_left.n28 drain_left.n0 8.14595
R559 drain_left.n65 drain_left.n37 8.14595
R560 drain_left drain_left.n73 6.19632
R561 drain_left.n30 drain_left.n0 5.81868
R562 drain_left.n67 drain_left.n37 5.81868
R563 drain_left.n28 drain_left.n27 5.04292
R564 drain_left.n65 drain_left.n64 5.04292
R565 drain_left.n13 drain_left.n9 4.38594
R566 drain_left.n50 drain_left.n46 4.38594
R567 drain_left.n24 drain_left.n2 4.26717
R568 drain_left.n61 drain_left.n39 4.26717
R569 drain_left.n23 drain_left.n4 3.49141
R570 drain_left.n60 drain_left.n41 3.49141
R571 drain_left.n33 drain_left.t13 3.3005
R572 drain_left.n33 drain_left.t7 3.3005
R573 drain_left.n34 drain_left.t11 3.3005
R574 drain_left.n34 drain_left.t6 3.3005
R575 drain_left.n31 drain_left.t10 3.3005
R576 drain_left.n31 drain_left.t3 3.3005
R577 drain_left.n72 drain_left.t5 3.3005
R578 drain_left.n72 drain_left.t1 3.3005
R579 drain_left.n70 drain_left.t0 3.3005
R580 drain_left.n70 drain_left.t9 3.3005
R581 drain_left.n68 drain_left.t8 3.3005
R582 drain_left.n68 drain_left.t4 3.3005
R583 drain_left.n20 drain_left.n19 2.71565
R584 drain_left.n57 drain_left.n56 2.71565
R585 drain_left.n16 drain_left.n6 1.93989
R586 drain_left.n53 drain_left.n43 1.93989
R587 drain_left.n15 drain_left.n8 1.16414
R588 drain_left.n52 drain_left.n45 1.16414
R589 drain_left.n71 drain_left.n69 0.543603
R590 drain_left.n73 drain_left.n71 0.543603
R591 drain_left.n12 drain_left.n11 0.388379
R592 drain_left.n49 drain_left.n48 0.388379
R593 drain_left.n36 drain_left.n32 0.352482
R594 drain_left.n14 drain_left.n13 0.155672
R595 drain_left.n14 drain_left.n5 0.155672
R596 drain_left.n21 drain_left.n5 0.155672
R597 drain_left.n22 drain_left.n21 0.155672
R598 drain_left.n22 drain_left.n1 0.155672
R599 drain_left.n29 drain_left.n1 0.155672
R600 drain_left.n66 drain_left.n38 0.155672
R601 drain_left.n59 drain_left.n38 0.155672
R602 drain_left.n59 drain_left.n58 0.155672
R603 drain_left.n58 drain_left.n42 0.155672
R604 drain_left.n51 drain_left.n42 0.155672
R605 drain_left.n51 drain_left.n50 0.155672
R606 drain_left.n36 drain_left.n35 0.0809298
C0 drain_left drain_right 0.881295f
C1 source drain_right 15.325701f
C2 plus minus 4.18806f
C3 minus drain_right 2.87378f
C4 plus drain_right 0.32231f
C5 drain_left source 15.3313f
C6 drain_left minus 0.171678f
C7 source minus 2.84488f
C8 drain_left plus 3.03901f
C9 source plus 2.85922f
C10 drain_right a_n1724_n2088# 5.49462f
C11 drain_left a_n1724_n2088# 5.7671f
C12 source a_n1724_n2088# 3.994913f
C13 minus a_n1724_n2088# 6.231949f
C14 plus a_n1724_n2088# 7.82006f
C15 drain_left.n0 a_n1724_n2088# 0.042639f
C16 drain_left.n1 a_n1724_n2088# 0.030335f
C17 drain_left.n2 a_n1724_n2088# 0.016301f
C18 drain_left.n3 a_n1724_n2088# 0.038529f
C19 drain_left.n4 a_n1724_n2088# 0.01726f
C20 drain_left.n5 a_n1724_n2088# 0.030335f
C21 drain_left.n6 a_n1724_n2088# 0.016301f
C22 drain_left.n7 a_n1724_n2088# 0.038529f
C23 drain_left.n8 a_n1724_n2088# 0.01726f
C24 drain_left.n9 a_n1724_n2088# 0.129814f
C25 drain_left.t2 a_n1724_n2088# 0.062798f
C26 drain_left.n10 a_n1724_n2088# 0.028897f
C27 drain_left.n11 a_n1724_n2088# 0.022759f
C28 drain_left.n12 a_n1724_n2088# 0.016301f
C29 drain_left.n13 a_n1724_n2088# 0.721798f
C30 drain_left.n14 a_n1724_n2088# 0.030335f
C31 drain_left.n15 a_n1724_n2088# 0.016301f
C32 drain_left.n16 a_n1724_n2088# 0.01726f
C33 drain_left.n17 a_n1724_n2088# 0.038529f
C34 drain_left.n18 a_n1724_n2088# 0.038529f
C35 drain_left.n19 a_n1724_n2088# 0.01726f
C36 drain_left.n20 a_n1724_n2088# 0.016301f
C37 drain_left.n21 a_n1724_n2088# 0.030335f
C38 drain_left.n22 a_n1724_n2088# 0.030335f
C39 drain_left.n23 a_n1724_n2088# 0.016301f
C40 drain_left.n24 a_n1724_n2088# 0.01726f
C41 drain_left.n25 a_n1724_n2088# 0.038529f
C42 drain_left.n26 a_n1724_n2088# 0.083409f
C43 drain_left.n27 a_n1724_n2088# 0.01726f
C44 drain_left.n28 a_n1724_n2088# 0.016301f
C45 drain_left.n29 a_n1724_n2088# 0.070119f
C46 drain_left.n30 a_n1724_n2088# 0.068842f
C47 drain_left.t10 a_n1724_n2088# 0.143831f
C48 drain_left.t3 a_n1724_n2088# 0.143831f
C49 drain_left.n31 a_n1724_n2088# 1.19955f
C50 drain_left.n32 a_n1724_n2088# 0.445975f
C51 drain_left.t13 a_n1724_n2088# 0.143831f
C52 drain_left.t7 a_n1724_n2088# 0.143831f
C53 drain_left.n33 a_n1724_n2088# 1.20248f
C54 drain_left.t11 a_n1724_n2088# 0.143831f
C55 drain_left.t6 a_n1724_n2088# 0.143831f
C56 drain_left.n34 a_n1724_n2088# 1.19955f
C57 drain_left.n35 a_n1724_n2088# 0.677584f
C58 drain_left.n36 a_n1724_n2088# 1.04826f
C59 drain_left.n37 a_n1724_n2088# 0.042639f
C60 drain_left.n38 a_n1724_n2088# 0.030335f
C61 drain_left.n39 a_n1724_n2088# 0.016301f
C62 drain_left.n40 a_n1724_n2088# 0.038529f
C63 drain_left.n41 a_n1724_n2088# 0.01726f
C64 drain_left.n42 a_n1724_n2088# 0.030335f
C65 drain_left.n43 a_n1724_n2088# 0.016301f
C66 drain_left.n44 a_n1724_n2088# 0.038529f
C67 drain_left.n45 a_n1724_n2088# 0.01726f
C68 drain_left.n46 a_n1724_n2088# 0.129814f
C69 drain_left.t12 a_n1724_n2088# 0.062798f
C70 drain_left.n47 a_n1724_n2088# 0.028897f
C71 drain_left.n48 a_n1724_n2088# 0.022759f
C72 drain_left.n49 a_n1724_n2088# 0.016301f
C73 drain_left.n50 a_n1724_n2088# 0.721798f
C74 drain_left.n51 a_n1724_n2088# 0.030335f
C75 drain_left.n52 a_n1724_n2088# 0.016301f
C76 drain_left.n53 a_n1724_n2088# 0.01726f
C77 drain_left.n54 a_n1724_n2088# 0.038529f
C78 drain_left.n55 a_n1724_n2088# 0.038529f
C79 drain_left.n56 a_n1724_n2088# 0.01726f
C80 drain_left.n57 a_n1724_n2088# 0.016301f
C81 drain_left.n58 a_n1724_n2088# 0.030335f
C82 drain_left.n59 a_n1724_n2088# 0.030335f
C83 drain_left.n60 a_n1724_n2088# 0.016301f
C84 drain_left.n61 a_n1724_n2088# 0.01726f
C85 drain_left.n62 a_n1724_n2088# 0.038529f
C86 drain_left.n63 a_n1724_n2088# 0.083409f
C87 drain_left.n64 a_n1724_n2088# 0.01726f
C88 drain_left.n65 a_n1724_n2088# 0.016301f
C89 drain_left.n66 a_n1724_n2088# 0.070119f
C90 drain_left.n67 a_n1724_n2088# 0.068842f
C91 drain_left.t8 a_n1724_n2088# 0.143831f
C92 drain_left.t4 a_n1724_n2088# 0.143831f
C93 drain_left.n68 a_n1724_n2088# 1.19956f
C94 drain_left.n69 a_n1724_n2088# 0.462653f
C95 drain_left.t0 a_n1724_n2088# 0.143831f
C96 drain_left.t9 a_n1724_n2088# 0.143831f
C97 drain_left.n70 a_n1724_n2088# 1.19956f
C98 drain_left.n71 a_n1724_n2088# 0.35238f
C99 drain_left.t5 a_n1724_n2088# 0.143831f
C100 drain_left.t1 a_n1724_n2088# 0.143831f
C101 drain_left.n72 a_n1724_n2088# 1.19955f
C102 drain_left.n73 a_n1724_n2088# 0.604884f
C103 plus.n0 a_n1724_n2088# 0.052973f
C104 plus.t8 a_n1724_n2088# 0.271672f
C105 plus.t4 a_n1724_n2088# 0.271672f
C106 plus.t13 a_n1724_n2088# 0.271672f
C107 plus.n1 a_n1724_n2088# 0.142275f
C108 plus.n2 a_n1724_n2088# 0.124804f
C109 plus.t9 a_n1724_n2088# 0.271672f
C110 plus.t5 a_n1724_n2088# 0.271672f
C111 plus.t1 a_n1724_n2088# 0.283262f
C112 plus.n3 a_n1724_n2088# 0.14122f
C113 plus.n4 a_n1724_n2088# 0.124702f
C114 plus.n5 a_n1724_n2088# 0.021819f
C115 plus.n6 a_n1724_n2088# 0.124702f
C116 plus.n7 a_n1724_n2088# 0.021819f
C117 plus.n8 a_n1724_n2088# 0.052973f
C118 plus.n9 a_n1724_n2088# 0.052973f
C119 plus.n10 a_n1724_n2088# 0.052973f
C120 plus.n11 a_n1724_n2088# 0.021819f
C121 plus.n12 a_n1724_n2088# 0.124702f
C122 plus.n13 a_n1724_n2088# 0.021819f
C123 plus.n14 a_n1724_n2088# 0.124702f
C124 plus.t12 a_n1724_n2088# 0.283262f
C125 plus.n15 a_n1724_n2088# 0.141136f
C126 plus.n16 a_n1724_n2088# 0.458664f
C127 plus.n17 a_n1724_n2088# 0.052973f
C128 plus.t11 a_n1724_n2088# 0.283262f
C129 plus.t3 a_n1724_n2088# 0.271672f
C130 plus.t10 a_n1724_n2088# 0.271672f
C131 plus.t2 a_n1724_n2088# 0.271672f
C132 plus.n18 a_n1724_n2088# 0.142275f
C133 plus.n19 a_n1724_n2088# 0.124804f
C134 plus.t7 a_n1724_n2088# 0.271672f
C135 plus.t0 a_n1724_n2088# 0.271672f
C136 plus.t6 a_n1724_n2088# 0.283262f
C137 plus.n20 a_n1724_n2088# 0.14122f
C138 plus.n21 a_n1724_n2088# 0.124702f
C139 plus.n22 a_n1724_n2088# 0.021819f
C140 plus.n23 a_n1724_n2088# 0.124702f
C141 plus.n24 a_n1724_n2088# 0.021819f
C142 plus.n25 a_n1724_n2088# 0.052973f
C143 plus.n26 a_n1724_n2088# 0.052973f
C144 plus.n27 a_n1724_n2088# 0.052973f
C145 plus.n28 a_n1724_n2088# 0.021819f
C146 plus.n29 a_n1724_n2088# 0.124702f
C147 plus.n30 a_n1724_n2088# 0.021819f
C148 plus.n31 a_n1724_n2088# 0.124702f
C149 plus.n32 a_n1724_n2088# 0.141136f
C150 plus.n33 a_n1724_n2088# 1.32815f
C151 drain_right.n0 a_n1724_n2088# 0.042683f
C152 drain_right.n1 a_n1724_n2088# 0.030366f
C153 drain_right.n2 a_n1724_n2088# 0.016318f
C154 drain_right.n3 a_n1724_n2088# 0.038569f
C155 drain_right.n4 a_n1724_n2088# 0.017277f
C156 drain_right.n5 a_n1724_n2088# 0.030366f
C157 drain_right.n6 a_n1724_n2088# 0.016318f
C158 drain_right.n7 a_n1724_n2088# 0.038569f
C159 drain_right.n8 a_n1724_n2088# 0.017277f
C160 drain_right.n9 a_n1724_n2088# 0.129947f
C161 drain_right.t2 a_n1724_n2088# 0.062862f
C162 drain_right.n10 a_n1724_n2088# 0.028927f
C163 drain_right.n11 a_n1724_n2088# 0.022782f
C164 drain_right.n12 a_n1724_n2088# 0.016318f
C165 drain_right.n13 a_n1724_n2088# 0.722539f
C166 drain_right.n14 a_n1724_n2088# 0.030366f
C167 drain_right.n15 a_n1724_n2088# 0.016318f
C168 drain_right.n16 a_n1724_n2088# 0.017277f
C169 drain_right.n17 a_n1724_n2088# 0.038569f
C170 drain_right.n18 a_n1724_n2088# 0.038569f
C171 drain_right.n19 a_n1724_n2088# 0.017277f
C172 drain_right.n20 a_n1724_n2088# 0.016318f
C173 drain_right.n21 a_n1724_n2088# 0.030366f
C174 drain_right.n22 a_n1724_n2088# 0.030366f
C175 drain_right.n23 a_n1724_n2088# 0.016318f
C176 drain_right.n24 a_n1724_n2088# 0.017277f
C177 drain_right.n25 a_n1724_n2088# 0.038569f
C178 drain_right.n26 a_n1724_n2088# 0.083495f
C179 drain_right.n27 a_n1724_n2088# 0.017277f
C180 drain_right.n28 a_n1724_n2088# 0.016318f
C181 drain_right.n29 a_n1724_n2088# 0.07019f
C182 drain_right.n30 a_n1724_n2088# 0.068913f
C183 drain_right.t7 a_n1724_n2088# 0.143979f
C184 drain_right.t3 a_n1724_n2088# 0.143979f
C185 drain_right.n31 a_n1724_n2088# 1.20078f
C186 drain_right.n32 a_n1724_n2088# 0.446433f
C187 drain_right.t6 a_n1724_n2088# 0.143979f
C188 drain_right.t13 a_n1724_n2088# 0.143979f
C189 drain_right.n33 a_n1724_n2088# 1.20371f
C190 drain_right.t8 a_n1724_n2088# 0.143979f
C191 drain_right.t12 a_n1724_n2088# 0.143979f
C192 drain_right.n34 a_n1724_n2088# 1.20078f
C193 drain_right.n35 a_n1724_n2088# 0.67828f
C194 drain_right.n36 a_n1724_n2088# 0.987578f
C195 drain_right.t0 a_n1724_n2088# 0.143979f
C196 drain_right.t4 a_n1724_n2088# 0.143979f
C197 drain_right.n37 a_n1724_n2088# 1.20371f
C198 drain_right.t5 a_n1724_n2088# 0.143979f
C199 drain_right.t10 a_n1724_n2088# 0.143979f
C200 drain_right.n38 a_n1724_n2088# 1.20079f
C201 drain_right.n39 a_n1724_n2088# 0.714793f
C202 drain_right.t11 a_n1724_n2088# 0.143979f
C203 drain_right.t1 a_n1724_n2088# 0.143979f
C204 drain_right.n40 a_n1724_n2088# 1.20079f
C205 drain_right.n41 a_n1724_n2088# 0.352741f
C206 drain_right.n42 a_n1724_n2088# 0.042683f
C207 drain_right.n43 a_n1724_n2088# 0.030366f
C208 drain_right.n44 a_n1724_n2088# 0.016318f
C209 drain_right.n45 a_n1724_n2088# 0.038569f
C210 drain_right.n46 a_n1724_n2088# 0.017277f
C211 drain_right.n47 a_n1724_n2088# 0.030366f
C212 drain_right.n48 a_n1724_n2088# 0.016318f
C213 drain_right.n49 a_n1724_n2088# 0.038569f
C214 drain_right.n50 a_n1724_n2088# 0.017277f
C215 drain_right.n51 a_n1724_n2088# 0.129947f
C216 drain_right.t9 a_n1724_n2088# 0.062862f
C217 drain_right.n52 a_n1724_n2088# 0.028927f
C218 drain_right.n53 a_n1724_n2088# 0.022782f
C219 drain_right.n54 a_n1724_n2088# 0.016318f
C220 drain_right.n55 a_n1724_n2088# 0.722539f
C221 drain_right.n56 a_n1724_n2088# 0.030366f
C222 drain_right.n57 a_n1724_n2088# 0.016318f
C223 drain_right.n58 a_n1724_n2088# 0.017277f
C224 drain_right.n59 a_n1724_n2088# 0.038569f
C225 drain_right.n60 a_n1724_n2088# 0.038569f
C226 drain_right.n61 a_n1724_n2088# 0.017277f
C227 drain_right.n62 a_n1724_n2088# 0.016318f
C228 drain_right.n63 a_n1724_n2088# 0.030366f
C229 drain_right.n64 a_n1724_n2088# 0.030366f
C230 drain_right.n65 a_n1724_n2088# 0.016318f
C231 drain_right.n66 a_n1724_n2088# 0.017277f
C232 drain_right.n67 a_n1724_n2088# 0.038569f
C233 drain_right.n68 a_n1724_n2088# 0.083495f
C234 drain_right.n69 a_n1724_n2088# 0.017277f
C235 drain_right.n70 a_n1724_n2088# 0.016318f
C236 drain_right.n71 a_n1724_n2088# 0.07019f
C237 drain_right.n72 a_n1724_n2088# 0.067686f
C238 drain_right.n73 a_n1724_n2088# 0.364945f
C239 source.n0 a_n1724_n2088# 0.046311f
C240 source.n1 a_n1724_n2088# 0.032948f
C241 source.n2 a_n1724_n2088# 0.017705f
C242 source.n3 a_n1724_n2088# 0.041848f
C243 source.n4 a_n1724_n2088# 0.018746f
C244 source.n5 a_n1724_n2088# 0.032948f
C245 source.n6 a_n1724_n2088# 0.017705f
C246 source.n7 a_n1724_n2088# 0.041848f
C247 source.n8 a_n1724_n2088# 0.018746f
C248 source.n9 a_n1724_n2088# 0.140994f
C249 source.t12 a_n1724_n2088# 0.068206f
C250 source.n10 a_n1724_n2088# 0.031386f
C251 source.n11 a_n1724_n2088# 0.024719f
C252 source.n12 a_n1724_n2088# 0.017705f
C253 source.n13 a_n1724_n2088# 0.783963f
C254 source.n14 a_n1724_n2088# 0.032948f
C255 source.n15 a_n1724_n2088# 0.017705f
C256 source.n16 a_n1724_n2088# 0.018746f
C257 source.n17 a_n1724_n2088# 0.041848f
C258 source.n18 a_n1724_n2088# 0.041848f
C259 source.n19 a_n1724_n2088# 0.018746f
C260 source.n20 a_n1724_n2088# 0.017705f
C261 source.n21 a_n1724_n2088# 0.032948f
C262 source.n22 a_n1724_n2088# 0.032948f
C263 source.n23 a_n1724_n2088# 0.017705f
C264 source.n24 a_n1724_n2088# 0.018746f
C265 source.n25 a_n1724_n2088# 0.041848f
C266 source.n26 a_n1724_n2088# 0.090593f
C267 source.n27 a_n1724_n2088# 0.018746f
C268 source.n28 a_n1724_n2088# 0.017705f
C269 source.n29 a_n1724_n2088# 0.076158f
C270 source.n30 a_n1724_n2088# 0.05069f
C271 source.n31 a_n1724_n2088# 0.798064f
C272 source.t10 a_n1724_n2088# 0.156218f
C273 source.t1 a_n1724_n2088# 0.156218f
C274 source.n32 a_n1724_n2088# 1.21664f
C275 source.n33 a_n1724_n2088# 0.424172f
C276 source.t2 a_n1724_n2088# 0.156218f
C277 source.t9 a_n1724_n2088# 0.156218f
C278 source.n34 a_n1724_n2088# 1.21664f
C279 source.n35 a_n1724_n2088# 0.424172f
C280 source.t11 a_n1724_n2088# 0.156218f
C281 source.t0 a_n1724_n2088# 0.156218f
C282 source.n36 a_n1724_n2088# 1.21664f
C283 source.n37 a_n1724_n2088# 0.445223f
C284 source.n38 a_n1724_n2088# 0.046311f
C285 source.n39 a_n1724_n2088# 0.032948f
C286 source.n40 a_n1724_n2088# 0.017705f
C287 source.n41 a_n1724_n2088# 0.041848f
C288 source.n42 a_n1724_n2088# 0.018746f
C289 source.n43 a_n1724_n2088# 0.032948f
C290 source.n44 a_n1724_n2088# 0.017705f
C291 source.n45 a_n1724_n2088# 0.041848f
C292 source.n46 a_n1724_n2088# 0.018746f
C293 source.n47 a_n1724_n2088# 0.140994f
C294 source.t22 a_n1724_n2088# 0.068206f
C295 source.n48 a_n1724_n2088# 0.031386f
C296 source.n49 a_n1724_n2088# 0.024719f
C297 source.n50 a_n1724_n2088# 0.017705f
C298 source.n51 a_n1724_n2088# 0.783963f
C299 source.n52 a_n1724_n2088# 0.032948f
C300 source.n53 a_n1724_n2088# 0.017705f
C301 source.n54 a_n1724_n2088# 0.018746f
C302 source.n55 a_n1724_n2088# 0.041848f
C303 source.n56 a_n1724_n2088# 0.041848f
C304 source.n57 a_n1724_n2088# 0.018746f
C305 source.n58 a_n1724_n2088# 0.017705f
C306 source.n59 a_n1724_n2088# 0.032948f
C307 source.n60 a_n1724_n2088# 0.032948f
C308 source.n61 a_n1724_n2088# 0.017705f
C309 source.n62 a_n1724_n2088# 0.018746f
C310 source.n63 a_n1724_n2088# 0.041848f
C311 source.n64 a_n1724_n2088# 0.090593f
C312 source.n65 a_n1724_n2088# 0.018746f
C313 source.n66 a_n1724_n2088# 0.017705f
C314 source.n67 a_n1724_n2088# 0.076158f
C315 source.n68 a_n1724_n2088# 0.05069f
C316 source.n69 a_n1724_n2088# 0.164508f
C317 source.t15 a_n1724_n2088# 0.156218f
C318 source.t19 a_n1724_n2088# 0.156218f
C319 source.n70 a_n1724_n2088# 1.21664f
C320 source.n71 a_n1724_n2088# 0.424172f
C321 source.t25 a_n1724_n2088# 0.156218f
C322 source.t27 a_n1724_n2088# 0.156218f
C323 source.n72 a_n1724_n2088# 1.21664f
C324 source.n73 a_n1724_n2088# 0.424172f
C325 source.t16 a_n1724_n2088# 0.156218f
C326 source.t14 a_n1724_n2088# 0.156218f
C327 source.n74 a_n1724_n2088# 1.21664f
C328 source.n75 a_n1724_n2088# 1.56061f
C329 source.t8 a_n1724_n2088# 0.156218f
C330 source.t6 a_n1724_n2088# 0.156218f
C331 source.n76 a_n1724_n2088# 1.21663f
C332 source.n77 a_n1724_n2088# 1.56062f
C333 source.t4 a_n1724_n2088# 0.156218f
C334 source.t5 a_n1724_n2088# 0.156218f
C335 source.n78 a_n1724_n2088# 1.21663f
C336 source.n79 a_n1724_n2088# 0.424181f
C337 source.t3 a_n1724_n2088# 0.156218f
C338 source.t7 a_n1724_n2088# 0.156218f
C339 source.n80 a_n1724_n2088# 1.21663f
C340 source.n81 a_n1724_n2088# 0.424181f
C341 source.n82 a_n1724_n2088# 0.046311f
C342 source.n83 a_n1724_n2088# 0.032948f
C343 source.n84 a_n1724_n2088# 0.017705f
C344 source.n85 a_n1724_n2088# 0.041848f
C345 source.n86 a_n1724_n2088# 0.018746f
C346 source.n87 a_n1724_n2088# 0.032948f
C347 source.n88 a_n1724_n2088# 0.017705f
C348 source.n89 a_n1724_n2088# 0.041848f
C349 source.n90 a_n1724_n2088# 0.018746f
C350 source.n91 a_n1724_n2088# 0.140994f
C351 source.t13 a_n1724_n2088# 0.068206f
C352 source.n92 a_n1724_n2088# 0.031386f
C353 source.n93 a_n1724_n2088# 0.024719f
C354 source.n94 a_n1724_n2088# 0.017705f
C355 source.n95 a_n1724_n2088# 0.783963f
C356 source.n96 a_n1724_n2088# 0.032948f
C357 source.n97 a_n1724_n2088# 0.017705f
C358 source.n98 a_n1724_n2088# 0.018746f
C359 source.n99 a_n1724_n2088# 0.041848f
C360 source.n100 a_n1724_n2088# 0.041848f
C361 source.n101 a_n1724_n2088# 0.018746f
C362 source.n102 a_n1724_n2088# 0.017705f
C363 source.n103 a_n1724_n2088# 0.032948f
C364 source.n104 a_n1724_n2088# 0.032948f
C365 source.n105 a_n1724_n2088# 0.017705f
C366 source.n106 a_n1724_n2088# 0.018746f
C367 source.n107 a_n1724_n2088# 0.041848f
C368 source.n108 a_n1724_n2088# 0.090593f
C369 source.n109 a_n1724_n2088# 0.018746f
C370 source.n110 a_n1724_n2088# 0.017705f
C371 source.n111 a_n1724_n2088# 0.076158f
C372 source.n112 a_n1724_n2088# 0.05069f
C373 source.n113 a_n1724_n2088# 0.164508f
C374 source.t17 a_n1724_n2088# 0.156218f
C375 source.t24 a_n1724_n2088# 0.156218f
C376 source.n114 a_n1724_n2088# 1.21663f
C377 source.n115 a_n1724_n2088# 0.445231f
C378 source.t26 a_n1724_n2088# 0.156218f
C379 source.t23 a_n1724_n2088# 0.156218f
C380 source.n116 a_n1724_n2088# 1.21663f
C381 source.n117 a_n1724_n2088# 0.424181f
C382 source.t18 a_n1724_n2088# 0.156218f
C383 source.t21 a_n1724_n2088# 0.156218f
C384 source.n118 a_n1724_n2088# 1.21663f
C385 source.n119 a_n1724_n2088# 0.424181f
C386 source.n120 a_n1724_n2088# 0.046311f
C387 source.n121 a_n1724_n2088# 0.032948f
C388 source.n122 a_n1724_n2088# 0.017705f
C389 source.n123 a_n1724_n2088# 0.041848f
C390 source.n124 a_n1724_n2088# 0.018746f
C391 source.n125 a_n1724_n2088# 0.032948f
C392 source.n126 a_n1724_n2088# 0.017705f
C393 source.n127 a_n1724_n2088# 0.041848f
C394 source.n128 a_n1724_n2088# 0.018746f
C395 source.n129 a_n1724_n2088# 0.140994f
C396 source.t20 a_n1724_n2088# 0.068206f
C397 source.n130 a_n1724_n2088# 0.031386f
C398 source.n131 a_n1724_n2088# 0.024719f
C399 source.n132 a_n1724_n2088# 0.017705f
C400 source.n133 a_n1724_n2088# 0.783963f
C401 source.n134 a_n1724_n2088# 0.032948f
C402 source.n135 a_n1724_n2088# 0.017705f
C403 source.n136 a_n1724_n2088# 0.018746f
C404 source.n137 a_n1724_n2088# 0.041848f
C405 source.n138 a_n1724_n2088# 0.041848f
C406 source.n139 a_n1724_n2088# 0.018746f
C407 source.n140 a_n1724_n2088# 0.017705f
C408 source.n141 a_n1724_n2088# 0.032948f
C409 source.n142 a_n1724_n2088# 0.032948f
C410 source.n143 a_n1724_n2088# 0.017705f
C411 source.n144 a_n1724_n2088# 0.018746f
C412 source.n145 a_n1724_n2088# 0.041848f
C413 source.n146 a_n1724_n2088# 0.090593f
C414 source.n147 a_n1724_n2088# 0.018746f
C415 source.n148 a_n1724_n2088# 0.017705f
C416 source.n149 a_n1724_n2088# 0.076158f
C417 source.n150 a_n1724_n2088# 0.05069f
C418 source.n151 a_n1724_n2088# 0.321669f
C419 source.n152 a_n1724_n2088# 1.34817f
C420 minus.n0 a_n1724_n2088# 0.051379f
C421 minus.t4 a_n1724_n2088# 0.274739f
C422 minus.t2 a_n1724_n2088# 0.263498f
C423 minus.t12 a_n1724_n2088# 0.263498f
C424 minus.t8 a_n1724_n2088# 0.263498f
C425 minus.n1 a_n1724_n2088# 0.137994f
C426 minus.n2 a_n1724_n2088# 0.121049f
C427 minus.t3 a_n1724_n2088# 0.263498f
C428 minus.t13 a_n1724_n2088# 0.263498f
C429 minus.t9 a_n1724_n2088# 0.274739f
C430 minus.n3 a_n1724_n2088# 0.136971f
C431 minus.n4 a_n1724_n2088# 0.12095f
C432 minus.n5 a_n1724_n2088# 0.021162f
C433 minus.n6 a_n1724_n2088# 0.12095f
C434 minus.n7 a_n1724_n2088# 0.021162f
C435 minus.n8 a_n1724_n2088# 0.051379f
C436 minus.n9 a_n1724_n2088# 0.051379f
C437 minus.n10 a_n1724_n2088# 0.051379f
C438 minus.n11 a_n1724_n2088# 0.021162f
C439 minus.n12 a_n1724_n2088# 0.12095f
C440 minus.n13 a_n1724_n2088# 0.021162f
C441 minus.n14 a_n1724_n2088# 0.12095f
C442 minus.n15 a_n1724_n2088# 0.136889f
C443 minus.n16 a_n1724_n2088# 1.4255f
C444 minus.n17 a_n1724_n2088# 0.051379f
C445 minus.t7 a_n1724_n2088# 0.263498f
C446 minus.t1 a_n1724_n2088# 0.263498f
C447 minus.t5 a_n1724_n2088# 0.263498f
C448 minus.n18 a_n1724_n2088# 0.137994f
C449 minus.n19 a_n1724_n2088# 0.121049f
C450 minus.t10 a_n1724_n2088# 0.263498f
C451 minus.t6 a_n1724_n2088# 0.263498f
C452 minus.t11 a_n1724_n2088# 0.274739f
C453 minus.n20 a_n1724_n2088# 0.136971f
C454 minus.n21 a_n1724_n2088# 0.12095f
C455 minus.n22 a_n1724_n2088# 0.021162f
C456 minus.n23 a_n1724_n2088# 0.12095f
C457 minus.n24 a_n1724_n2088# 0.021162f
C458 minus.n25 a_n1724_n2088# 0.051379f
C459 minus.n26 a_n1724_n2088# 0.051379f
C460 minus.n27 a_n1724_n2088# 0.051379f
C461 minus.n28 a_n1724_n2088# 0.021162f
C462 minus.n29 a_n1724_n2088# 0.12095f
C463 minus.n30 a_n1724_n2088# 0.021162f
C464 minus.n31 a_n1724_n2088# 0.12095f
C465 minus.t0 a_n1724_n2088# 0.274739f
C466 minus.n32 a_n1724_n2088# 0.136889f
C467 minus.n33 a_n1724_n2088# 0.340311f
C468 minus.n34 a_n1724_n2088# 1.75279f
.ends

