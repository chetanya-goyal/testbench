* NGSPICE file created from diffpair334.ext - technology: sky130A

.subckt diffpair334 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t19 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X2 drain_right.t8 minus.t1 source.t12 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X3 drain_right.t7 minus.t2 source.t13 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 source.t16 minus.t3 drain_right.t6 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 source.t18 minus.t4 drain_right.t5 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X6 source.t4 plus.t0 drain_left.t9 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X7 drain_right.t4 minus.t5 source.t14 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X8 a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X9 source.t10 minus.t6 drain_right.t3 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X10 a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X11 drain_left.t8 plus.t1 source.t7 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X12 source.t3 plus.t2 drain_left.t7 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X13 drain_right.t2 minus.t7 source.t15 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X14 drain_right.t1 minus.t8 source.t17 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X15 drain_left.t6 plus.t3 source.t6 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X16 drain_left.t5 plus.t4 source.t8 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X17 drain_left.t4 plus.t5 source.t0 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X18 drain_left.t3 plus.t6 source.t1 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X19 source.t2 plus.t7 drain_left.t2 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X20 source.t5 plus.t8 drain_left.t1 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X21 source.t11 minus.t9 drain_right.t0 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X22 a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X23 drain_left.t0 plus.t9 source.t9 a_n1352_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n8 minus.t8 1286.43
R1 minus.n2 minus.t7 1286.43
R2 minus.n18 minus.t5 1286.43
R3 minus.n12 minus.t1 1286.43
R4 minus.n7 minus.t9 1241.15
R5 minus.n5 minus.t2 1241.15
R6 minus.n1 minus.t6 1241.15
R7 minus.n17 minus.t3 1241.15
R8 minus.n15 minus.t0 1241.15
R9 minus.n11 minus.t4 1241.15
R10 minus.n3 minus.n2 161.489
R11 minus.n13 minus.n12 161.489
R12 minus.n9 minus.n8 161.3
R13 minus.n6 minus.n0 161.3
R14 minus.n4 minus.n3 161.3
R15 minus.n19 minus.n18 161.3
R16 minus.n16 minus.n10 161.3
R17 minus.n14 minus.n13 161.3
R18 minus.n7 minus.n6 40.8975
R19 minus.n4 minus.n1 40.8975
R20 minus.n14 minus.n11 40.8975
R21 minus.n17 minus.n16 40.8975
R22 minus.n6 minus.n5 36.5157
R23 minus.n5 minus.n4 36.5157
R24 minus.n15 minus.n14 36.5157
R25 minus.n16 minus.n15 36.5157
R26 minus.n8 minus.n7 32.1338
R27 minus.n2 minus.n1 32.1338
R28 minus.n12 minus.n11 32.1338
R29 minus.n18 minus.n17 32.1338
R30 minus.n20 minus.n9 31.9191
R31 minus.n20 minus.n19 6.44936
R32 minus.n9 minus.n0 0.189894
R33 minus.n3 minus.n0 0.189894
R34 minus.n13 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n5 source.t15 51.0588
R38 source.n19 source.t14 51.0586
R39 source.n14 source.t8 51.0586
R40 source.n0 source.t1 51.0586
R41 source.n2 source.n1 48.8588
R42 source.n4 source.n3 48.8588
R43 source.n7 source.n6 48.8588
R44 source.n9 source.n8 48.8588
R45 source.n18 source.n17 48.8586
R46 source.n16 source.n15 48.8586
R47 source.n13 source.n12 48.8586
R48 source.n11 source.n10 48.8586
R49 source.n11 source.n9 19.9288
R50 source.n20 source.n0 13.9805
R51 source.n20 source.n19 5.49188
R52 source.n17 source.t19 2.2005
R53 source.n17 source.t16 2.2005
R54 source.n15 source.t12 2.2005
R55 source.n15 source.t18 2.2005
R56 source.n12 source.t0 2.2005
R57 source.n12 source.t5 2.2005
R58 source.n10 source.t6 2.2005
R59 source.n10 source.t3 2.2005
R60 source.n1 source.t9 2.2005
R61 source.n1 source.t2 2.2005
R62 source.n3 source.t7 2.2005
R63 source.n3 source.t4 2.2005
R64 source.n6 source.t13 2.2005
R65 source.n6 source.t10 2.2005
R66 source.n8 source.t17 2.2005
R67 source.n8 source.t11 2.2005
R68 source.n5 source.n4 0.698776
R69 source.n16 source.n14 0.698776
R70 source.n9 source.n7 0.457397
R71 source.n7 source.n5 0.457397
R72 source.n4 source.n2 0.457397
R73 source.n2 source.n0 0.457397
R74 source.n13 source.n11 0.457397
R75 source.n14 source.n13 0.457397
R76 source.n18 source.n16 0.457397
R77 source.n19 source.n18 0.457397
R78 source source.n20 0.188
R79 drain_right.n1 drain_right.t8 68.1942
R80 drain_right.n7 drain_right.t1 67.7376
R81 drain_right.n6 drain_right.n4 65.9943
R82 drain_right.n3 drain_right.n2 65.8247
R83 drain_right.n6 drain_right.n5 65.5376
R84 drain_right.n1 drain_right.n0 65.5373
R85 drain_right drain_right.n3 26.4829
R86 drain_right drain_right.n7 5.88166
R87 drain_right.n2 drain_right.t6 2.2005
R88 drain_right.n2 drain_right.t4 2.2005
R89 drain_right.n0 drain_right.t5 2.2005
R90 drain_right.n0 drain_right.t9 2.2005
R91 drain_right.n4 drain_right.t3 2.2005
R92 drain_right.n4 drain_right.t2 2.2005
R93 drain_right.n5 drain_right.t0 2.2005
R94 drain_right.n5 drain_right.t7 2.2005
R95 drain_right.n7 drain_right.n6 0.457397
R96 drain_right.n3 drain_right.n1 0.0593781
R97 plus.n2 plus.t1 1286.43
R98 plus.n8 plus.t6 1286.43
R99 plus.n12 plus.t4 1286.43
R100 plus.n18 plus.t3 1286.43
R101 plus.n1 plus.t0 1241.15
R102 plus.n5 plus.t9 1241.15
R103 plus.n7 plus.t7 1241.15
R104 plus.n11 plus.t8 1241.15
R105 plus.n15 plus.t5 1241.15
R106 plus.n17 plus.t2 1241.15
R107 plus.n3 plus.n2 161.489
R108 plus.n13 plus.n12 161.489
R109 plus.n4 plus.n3 161.3
R110 plus.n6 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n14 plus.n13 161.3
R113 plus.n16 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n4 plus.n1 40.8975
R116 plus.n7 plus.n6 40.8975
R117 plus.n17 plus.n16 40.8975
R118 plus.n14 plus.n11 40.8975
R119 plus.n5 plus.n4 36.5157
R120 plus.n6 plus.n5 36.5157
R121 plus.n16 plus.n15 36.5157
R122 plus.n15 plus.n14 36.5157
R123 plus.n2 plus.n1 32.1338
R124 plus.n8 plus.n7 32.1338
R125 plus.n18 plus.n17 32.1338
R126 plus.n12 plus.n11 32.1338
R127 plus plus.n19 26.9365
R128 plus plus.n9 10.9569
R129 plus.n3 plus.n0 0.189894
R130 plus.n9 plus.n0 0.189894
R131 plus.n19 plus.n10 0.189894
R132 plus.n13 plus.n10 0.189894
R133 drain_left.n5 drain_left.t8 68.1945
R134 drain_left.n1 drain_left.t6 68.1942
R135 drain_left.n3 drain_left.n2 65.8247
R136 drain_left.n5 drain_left.n4 65.5376
R137 drain_left.n7 drain_left.n6 65.5374
R138 drain_left.n1 drain_left.n0 65.5373
R139 drain_left drain_left.n3 27.0362
R140 drain_left drain_left.n7 6.11011
R141 drain_left.n2 drain_left.t1 2.2005
R142 drain_left.n2 drain_left.t5 2.2005
R143 drain_left.n0 drain_left.t7 2.2005
R144 drain_left.n0 drain_left.t4 2.2005
R145 drain_left.n6 drain_left.t2 2.2005
R146 drain_left.n6 drain_left.t3 2.2005
R147 drain_left.n4 drain_left.t9 2.2005
R148 drain_left.n4 drain_left.t0 2.2005
R149 drain_left.n7 drain_left.n5 0.457397
R150 drain_left.n3 drain_left.n1 0.0593781
C0 plus source 2.08254f
C1 drain_left minus 0.170748f
C2 drain_right minus 2.40031f
C3 drain_left source 19.2113f
C4 drain_right source 19.2015f
C5 drain_left plus 2.52601f
C6 drain_right plus 0.283112f
C7 drain_left drain_right 0.661658f
C8 minus source 2.06798f
C9 plus minus 4.285f
C10 drain_right a_n1352_n2688# 6.10943f
C11 drain_left a_n1352_n2688# 6.32328f
C12 source a_n1352_n2688# 4.932425f
C13 minus a_n1352_n2688# 5.01069f
C14 plus a_n1352_n2688# 6.86367f
C15 drain_left.t6 a_n1352_n2688# 2.61604f
C16 drain_left.t7 a_n1352_n2688# 0.23472f
C17 drain_left.t4 a_n1352_n2688# 0.23472f
C18 drain_left.n0 a_n1352_n2688# 2.05302f
C19 drain_left.n1 a_n1352_n2688# 0.735568f
C20 drain_left.t1 a_n1352_n2688# 0.23472f
C21 drain_left.t5 a_n1352_n2688# 0.23472f
C22 drain_left.n2 a_n1352_n2688# 2.05459f
C23 drain_left.n3 a_n1352_n2688# 1.56761f
C24 drain_left.t8 a_n1352_n2688# 2.61604f
C25 drain_left.t9 a_n1352_n2688# 0.23472f
C26 drain_left.t0 a_n1352_n2688# 0.23472f
C27 drain_left.n4 a_n1352_n2688# 2.05302f
C28 drain_left.n5 a_n1352_n2688# 0.764891f
C29 drain_left.t2 a_n1352_n2688# 0.23472f
C30 drain_left.t3 a_n1352_n2688# 0.23472f
C31 drain_left.n6 a_n1352_n2688# 2.05301f
C32 drain_left.n7 a_n1352_n2688# 0.631638f
C33 plus.n0 a_n1352_n2688# 0.058586f
C34 plus.t7 a_n1352_n2688# 0.298816f
C35 plus.t9 a_n1352_n2688# 0.298816f
C36 plus.t0 a_n1352_n2688# 0.298816f
C37 plus.n1 a_n1352_n2688# 0.1308f
C38 plus.t1 a_n1352_n2688# 0.303432f
C39 plus.n2 a_n1352_n2688# 0.147146f
C40 plus.n3 a_n1352_n2688# 0.128648f
C41 plus.n4 a_n1352_n2688# 0.020518f
C42 plus.n5 a_n1352_n2688# 0.1308f
C43 plus.n6 a_n1352_n2688# 0.020518f
C44 plus.n7 a_n1352_n2688# 0.1308f
C45 plus.t6 a_n1352_n2688# 0.303432f
C46 plus.n8 a_n1352_n2688# 0.147063f
C47 plus.n9 a_n1352_n2688# 0.568278f
C48 plus.n10 a_n1352_n2688# 0.058586f
C49 plus.t3 a_n1352_n2688# 0.303432f
C50 plus.t2 a_n1352_n2688# 0.298816f
C51 plus.t5 a_n1352_n2688# 0.298816f
C52 plus.t8 a_n1352_n2688# 0.298816f
C53 plus.n11 a_n1352_n2688# 0.1308f
C54 plus.t4 a_n1352_n2688# 0.303432f
C55 plus.n12 a_n1352_n2688# 0.147146f
C56 plus.n13 a_n1352_n2688# 0.128648f
C57 plus.n14 a_n1352_n2688# 0.020518f
C58 plus.n15 a_n1352_n2688# 0.1308f
C59 plus.n16 a_n1352_n2688# 0.020518f
C60 plus.n17 a_n1352_n2688# 0.1308f
C61 plus.n18 a_n1352_n2688# 0.147063f
C62 plus.n19 a_n1352_n2688# 1.46993f
C63 drain_right.t8 a_n1352_n2688# 2.61957f
C64 drain_right.t5 a_n1352_n2688# 0.235037f
C65 drain_right.t9 a_n1352_n2688# 0.235037f
C66 drain_right.n0 a_n1352_n2688# 2.05579f
C67 drain_right.n1 a_n1352_n2688# 0.73656f
C68 drain_right.t6 a_n1352_n2688# 0.235037f
C69 drain_right.t4 a_n1352_n2688# 0.235037f
C70 drain_right.n2 a_n1352_n2688# 2.05736f
C71 drain_right.n3 a_n1352_n2688# 1.50108f
C72 drain_right.t3 a_n1352_n2688# 0.235037f
C73 drain_right.t2 a_n1352_n2688# 0.235037f
C74 drain_right.n4 a_n1352_n2688# 2.05838f
C75 drain_right.t0 a_n1352_n2688# 0.235037f
C76 drain_right.t7 a_n1352_n2688# 0.235037f
C77 drain_right.n5 a_n1352_n2688# 2.05579f
C78 drain_right.n6 a_n1352_n2688# 0.734757f
C79 drain_right.t1 a_n1352_n2688# 2.61685f
C80 drain_right.n7 a_n1352_n2688# 0.675233f
C81 source.t1 a_n1352_n2688# 2.62587f
C82 source.n0 a_n1352_n2688# 1.49384f
C83 source.t9 a_n1352_n2688# 0.24625f
C84 source.t2 a_n1352_n2688# 0.24625f
C85 source.n1 a_n1352_n2688# 2.06144f
C86 source.n2 a_n1352_n2688# 0.424652f
C87 source.t7 a_n1352_n2688# 0.24625f
C88 source.t4 a_n1352_n2688# 0.24625f
C89 source.n3 a_n1352_n2688# 2.06144f
C90 source.n4 a_n1352_n2688# 0.451582f
C91 source.t15 a_n1352_n2688# 2.62588f
C92 source.n5 a_n1352_n2688# 0.558732f
C93 source.t13 a_n1352_n2688# 0.24625f
C94 source.t10 a_n1352_n2688# 0.24625f
C95 source.n6 a_n1352_n2688# 2.06144f
C96 source.n7 a_n1352_n2688# 0.424652f
C97 source.t17 a_n1352_n2688# 0.24625f
C98 source.t11 a_n1352_n2688# 0.24625f
C99 source.n8 a_n1352_n2688# 2.06144f
C100 source.n9 a_n1352_n2688# 1.93762f
C101 source.t6 a_n1352_n2688# 0.24625f
C102 source.t3 a_n1352_n2688# 0.24625f
C103 source.n10 a_n1352_n2688# 2.06143f
C104 source.n11 a_n1352_n2688# 1.93763f
C105 source.t0 a_n1352_n2688# 0.24625f
C106 source.t5 a_n1352_n2688# 0.24625f
C107 source.n12 a_n1352_n2688# 2.06143f
C108 source.n13 a_n1352_n2688# 0.424658f
C109 source.t8 a_n1352_n2688# 2.62587f
C110 source.n14 a_n1352_n2688# 0.558739f
C111 source.t12 a_n1352_n2688# 0.24625f
C112 source.t18 a_n1352_n2688# 0.24625f
C113 source.n15 a_n1352_n2688# 2.06143f
C114 source.n16 a_n1352_n2688# 0.451588f
C115 source.t19 a_n1352_n2688# 0.24625f
C116 source.t16 a_n1352_n2688# 0.24625f
C117 source.n17 a_n1352_n2688# 2.06143f
C118 source.n18 a_n1352_n2688# 0.424658f
C119 source.t14 a_n1352_n2688# 2.62587f
C120 source.n19 a_n1352_n2688# 0.720995f
C121 source.n20 a_n1352_n2688# 1.7974f
C122 minus.n0 a_n1352_n2688# 0.057166f
C123 minus.t8 a_n1352_n2688# 0.296081f
C124 minus.t9 a_n1352_n2688# 0.291577f
C125 minus.t2 a_n1352_n2688# 0.291577f
C126 minus.t6 a_n1352_n2688# 0.291577f
C127 minus.n1 a_n1352_n2688# 0.127632f
C128 minus.t7 a_n1352_n2688# 0.296081f
C129 minus.n2 a_n1352_n2688# 0.143581f
C130 minus.n3 a_n1352_n2688# 0.125531f
C131 minus.n4 a_n1352_n2688# 0.020021f
C132 minus.n5 a_n1352_n2688# 0.127632f
C133 minus.n6 a_n1352_n2688# 0.020021f
C134 minus.n7 a_n1352_n2688# 0.127632f
C135 minus.n8 a_n1352_n2688# 0.143501f
C136 minus.n9 a_n1352_n2688# 1.64802f
C137 minus.n10 a_n1352_n2688# 0.057166f
C138 minus.t3 a_n1352_n2688# 0.291577f
C139 minus.t0 a_n1352_n2688# 0.291577f
C140 minus.t4 a_n1352_n2688# 0.291577f
C141 minus.n11 a_n1352_n2688# 0.127632f
C142 minus.t1 a_n1352_n2688# 0.296081f
C143 minus.n12 a_n1352_n2688# 0.143581f
C144 minus.n13 a_n1352_n2688# 0.125531f
C145 minus.n14 a_n1352_n2688# 0.020021f
C146 minus.n15 a_n1352_n2688# 0.127632f
C147 minus.n16 a_n1352_n2688# 0.020021f
C148 minus.n17 a_n1352_n2688# 0.127632f
C149 minus.t5 a_n1352_n2688# 0.296081f
C150 minus.n18 a_n1352_n2688# 0.143501f
C151 minus.n19 a_n1352_n2688# 0.366903f
C152 minus.n20 a_n1352_n2688# 2.02832f
.ends

