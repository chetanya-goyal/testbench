* NGSPICE file created from diffpair412.ext - technology: sky130A

.subckt diffpair412 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t8 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X1 drain_right.t4 minus.t1 source.t10 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X2 drain_right.t3 minus.t2 source.t6 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X3 source.t0 plus.t0 drain_left.t5 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X4 source.t7 minus.t3 drain_right.t2 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X5 source.t11 minus.t4 drain_right.t1 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
X6 a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.2
X7 drain_left.t4 plus.t1 source.t2 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X8 a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X9 a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X10 drain_right.t0 minus.t5 source.t9 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X11 drain_left.t3 plus.t2 source.t5 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.2
X12 drain_left.t2 plus.t3 source.t4 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X13 a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.2
X14 drain_left.t1 plus.t4 source.t1 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.2
X15 source.t3 plus.t5 drain_left.t0 a_n1140_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.2
R0 minus.n2 minus.t0 1643.55
R1 minus.n0 minus.t5 1643.55
R2 minus.n6 minus.t1 1643.55
R3 minus.n4 minus.t2 1643.55
R4 minus.n1 minus.t4 1602.65
R5 minus.n5 minus.t3 1602.65
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 33.3774
R15 minus.n8 minus.n7 6.438
R16 minus minus.n8 0.188
R17 source.n266 source.n206 289.615
R18 source.n198 source.n138 289.615
R19 source.n60 source.n0 289.615
R20 source.n128 source.n68 289.615
R21 source.n226 source.n225 185
R22 source.n231 source.n230 185
R23 source.n233 source.n232 185
R24 source.n222 source.n221 185
R25 source.n239 source.n238 185
R26 source.n241 source.n240 185
R27 source.n218 source.n217 185
R28 source.n248 source.n247 185
R29 source.n249 source.n216 185
R30 source.n251 source.n250 185
R31 source.n214 source.n213 185
R32 source.n257 source.n256 185
R33 source.n259 source.n258 185
R34 source.n210 source.n209 185
R35 source.n265 source.n264 185
R36 source.n267 source.n266 185
R37 source.n158 source.n157 185
R38 source.n163 source.n162 185
R39 source.n165 source.n164 185
R40 source.n154 source.n153 185
R41 source.n171 source.n170 185
R42 source.n173 source.n172 185
R43 source.n150 source.n149 185
R44 source.n180 source.n179 185
R45 source.n181 source.n148 185
R46 source.n183 source.n182 185
R47 source.n146 source.n145 185
R48 source.n189 source.n188 185
R49 source.n191 source.n190 185
R50 source.n142 source.n141 185
R51 source.n197 source.n196 185
R52 source.n199 source.n198 185
R53 source.n61 source.n60 185
R54 source.n59 source.n58 185
R55 source.n4 source.n3 185
R56 source.n53 source.n52 185
R57 source.n51 source.n50 185
R58 source.n8 source.n7 185
R59 source.n45 source.n44 185
R60 source.n43 source.n10 185
R61 source.n42 source.n41 185
R62 source.n13 source.n11 185
R63 source.n36 source.n35 185
R64 source.n34 source.n33 185
R65 source.n17 source.n16 185
R66 source.n28 source.n27 185
R67 source.n26 source.n25 185
R68 source.n21 source.n20 185
R69 source.n129 source.n128 185
R70 source.n127 source.n126 185
R71 source.n72 source.n71 185
R72 source.n121 source.n120 185
R73 source.n119 source.n118 185
R74 source.n76 source.n75 185
R75 source.n113 source.n112 185
R76 source.n111 source.n78 185
R77 source.n110 source.n109 185
R78 source.n81 source.n79 185
R79 source.n104 source.n103 185
R80 source.n102 source.n101 185
R81 source.n85 source.n84 185
R82 source.n96 source.n95 185
R83 source.n94 source.n93 185
R84 source.n89 source.n88 185
R85 source.n227 source.t10 149.524
R86 source.n159 source.t4 149.524
R87 source.n22 source.t1 149.524
R88 source.n90 source.t9 149.524
R89 source.n231 source.n225 104.615
R90 source.n232 source.n231 104.615
R91 source.n232 source.n221 104.615
R92 source.n239 source.n221 104.615
R93 source.n240 source.n239 104.615
R94 source.n240 source.n217 104.615
R95 source.n248 source.n217 104.615
R96 source.n249 source.n248 104.615
R97 source.n250 source.n249 104.615
R98 source.n250 source.n213 104.615
R99 source.n257 source.n213 104.615
R100 source.n258 source.n257 104.615
R101 source.n258 source.n209 104.615
R102 source.n265 source.n209 104.615
R103 source.n266 source.n265 104.615
R104 source.n163 source.n157 104.615
R105 source.n164 source.n163 104.615
R106 source.n164 source.n153 104.615
R107 source.n171 source.n153 104.615
R108 source.n172 source.n171 104.615
R109 source.n172 source.n149 104.615
R110 source.n180 source.n149 104.615
R111 source.n181 source.n180 104.615
R112 source.n182 source.n181 104.615
R113 source.n182 source.n145 104.615
R114 source.n189 source.n145 104.615
R115 source.n190 source.n189 104.615
R116 source.n190 source.n141 104.615
R117 source.n197 source.n141 104.615
R118 source.n198 source.n197 104.615
R119 source.n60 source.n59 104.615
R120 source.n59 source.n3 104.615
R121 source.n52 source.n3 104.615
R122 source.n52 source.n51 104.615
R123 source.n51 source.n7 104.615
R124 source.n44 source.n7 104.615
R125 source.n44 source.n43 104.615
R126 source.n43 source.n42 104.615
R127 source.n42 source.n11 104.615
R128 source.n35 source.n11 104.615
R129 source.n35 source.n34 104.615
R130 source.n34 source.n16 104.615
R131 source.n27 source.n16 104.615
R132 source.n27 source.n26 104.615
R133 source.n26 source.n20 104.615
R134 source.n128 source.n127 104.615
R135 source.n127 source.n71 104.615
R136 source.n120 source.n71 104.615
R137 source.n120 source.n119 104.615
R138 source.n119 source.n75 104.615
R139 source.n112 source.n75 104.615
R140 source.n112 source.n111 104.615
R141 source.n111 source.n110 104.615
R142 source.n110 source.n79 104.615
R143 source.n103 source.n79 104.615
R144 source.n103 source.n102 104.615
R145 source.n102 source.n84 104.615
R146 source.n95 source.n84 104.615
R147 source.n95 source.n94 104.615
R148 source.n94 source.n88 104.615
R149 source.t10 source.n225 52.3082
R150 source.t4 source.n157 52.3082
R151 source.t1 source.n20 52.3082
R152 source.t9 source.n88 52.3082
R153 source.n67 source.n66 42.8739
R154 source.n135 source.n134 42.8739
R155 source.n205 source.n204 42.8737
R156 source.n137 source.n136 42.8737
R157 source.n271 source.n270 29.8581
R158 source.n203 source.n202 29.8581
R159 source.n65 source.n64 29.8581
R160 source.n133 source.n132 29.8581
R161 source.n137 source.n135 22.2015
R162 source.n272 source.n65 16.2532
R163 source.n251 source.n216 13.1884
R164 source.n183 source.n148 13.1884
R165 source.n45 source.n10 13.1884
R166 source.n113 source.n78 13.1884
R167 source.n247 source.n246 12.8005
R168 source.n252 source.n214 12.8005
R169 source.n179 source.n178 12.8005
R170 source.n184 source.n146 12.8005
R171 source.n46 source.n8 12.8005
R172 source.n41 source.n12 12.8005
R173 source.n114 source.n76 12.8005
R174 source.n109 source.n80 12.8005
R175 source.n245 source.n218 12.0247
R176 source.n256 source.n255 12.0247
R177 source.n177 source.n150 12.0247
R178 source.n188 source.n187 12.0247
R179 source.n50 source.n49 12.0247
R180 source.n40 source.n13 12.0247
R181 source.n118 source.n117 12.0247
R182 source.n108 source.n81 12.0247
R183 source.n242 source.n241 11.249
R184 source.n259 source.n212 11.249
R185 source.n174 source.n173 11.249
R186 source.n191 source.n144 11.249
R187 source.n53 source.n6 11.249
R188 source.n37 source.n36 11.249
R189 source.n121 source.n74 11.249
R190 source.n105 source.n104 11.249
R191 source.n238 source.n220 10.4732
R192 source.n260 source.n210 10.4732
R193 source.n170 source.n152 10.4732
R194 source.n192 source.n142 10.4732
R195 source.n54 source.n4 10.4732
R196 source.n33 source.n15 10.4732
R197 source.n122 source.n72 10.4732
R198 source.n101 source.n83 10.4732
R199 source.n227 source.n226 10.2747
R200 source.n159 source.n158 10.2747
R201 source.n22 source.n21 10.2747
R202 source.n90 source.n89 10.2747
R203 source.n237 source.n222 9.69747
R204 source.n264 source.n263 9.69747
R205 source.n169 source.n154 9.69747
R206 source.n196 source.n195 9.69747
R207 source.n58 source.n57 9.69747
R208 source.n32 source.n17 9.69747
R209 source.n126 source.n125 9.69747
R210 source.n100 source.n85 9.69747
R211 source.n270 source.n269 9.45567
R212 source.n202 source.n201 9.45567
R213 source.n64 source.n63 9.45567
R214 source.n132 source.n131 9.45567
R215 source.n269 source.n268 9.3005
R216 source.n208 source.n207 9.3005
R217 source.n263 source.n262 9.3005
R218 source.n261 source.n260 9.3005
R219 source.n212 source.n211 9.3005
R220 source.n255 source.n254 9.3005
R221 source.n253 source.n252 9.3005
R222 source.n229 source.n228 9.3005
R223 source.n224 source.n223 9.3005
R224 source.n235 source.n234 9.3005
R225 source.n237 source.n236 9.3005
R226 source.n220 source.n219 9.3005
R227 source.n243 source.n242 9.3005
R228 source.n245 source.n244 9.3005
R229 source.n246 source.n215 9.3005
R230 source.n201 source.n200 9.3005
R231 source.n140 source.n139 9.3005
R232 source.n195 source.n194 9.3005
R233 source.n193 source.n192 9.3005
R234 source.n144 source.n143 9.3005
R235 source.n187 source.n186 9.3005
R236 source.n185 source.n184 9.3005
R237 source.n161 source.n160 9.3005
R238 source.n156 source.n155 9.3005
R239 source.n167 source.n166 9.3005
R240 source.n169 source.n168 9.3005
R241 source.n152 source.n151 9.3005
R242 source.n175 source.n174 9.3005
R243 source.n177 source.n176 9.3005
R244 source.n178 source.n147 9.3005
R245 source.n24 source.n23 9.3005
R246 source.n19 source.n18 9.3005
R247 source.n30 source.n29 9.3005
R248 source.n32 source.n31 9.3005
R249 source.n15 source.n14 9.3005
R250 source.n38 source.n37 9.3005
R251 source.n40 source.n39 9.3005
R252 source.n12 source.n9 9.3005
R253 source.n63 source.n62 9.3005
R254 source.n2 source.n1 9.3005
R255 source.n57 source.n56 9.3005
R256 source.n55 source.n54 9.3005
R257 source.n6 source.n5 9.3005
R258 source.n49 source.n48 9.3005
R259 source.n47 source.n46 9.3005
R260 source.n92 source.n91 9.3005
R261 source.n87 source.n86 9.3005
R262 source.n98 source.n97 9.3005
R263 source.n100 source.n99 9.3005
R264 source.n83 source.n82 9.3005
R265 source.n106 source.n105 9.3005
R266 source.n108 source.n107 9.3005
R267 source.n80 source.n77 9.3005
R268 source.n131 source.n130 9.3005
R269 source.n70 source.n69 9.3005
R270 source.n125 source.n124 9.3005
R271 source.n123 source.n122 9.3005
R272 source.n74 source.n73 9.3005
R273 source.n117 source.n116 9.3005
R274 source.n115 source.n114 9.3005
R275 source.n234 source.n233 8.92171
R276 source.n267 source.n208 8.92171
R277 source.n166 source.n165 8.92171
R278 source.n199 source.n140 8.92171
R279 source.n61 source.n2 8.92171
R280 source.n29 source.n28 8.92171
R281 source.n129 source.n70 8.92171
R282 source.n97 source.n96 8.92171
R283 source.n230 source.n224 8.14595
R284 source.n268 source.n206 8.14595
R285 source.n162 source.n156 8.14595
R286 source.n200 source.n138 8.14595
R287 source.n62 source.n0 8.14595
R288 source.n25 source.n19 8.14595
R289 source.n130 source.n68 8.14595
R290 source.n93 source.n87 8.14595
R291 source.n229 source.n226 7.3702
R292 source.n161 source.n158 7.3702
R293 source.n24 source.n21 7.3702
R294 source.n92 source.n89 7.3702
R295 source.n230 source.n229 5.81868
R296 source.n270 source.n206 5.81868
R297 source.n162 source.n161 5.81868
R298 source.n202 source.n138 5.81868
R299 source.n64 source.n0 5.81868
R300 source.n25 source.n24 5.81868
R301 source.n132 source.n68 5.81868
R302 source.n93 source.n92 5.81868
R303 source.n272 source.n271 5.49188
R304 source.n233 source.n224 5.04292
R305 source.n268 source.n267 5.04292
R306 source.n165 source.n156 5.04292
R307 source.n200 source.n199 5.04292
R308 source.n62 source.n61 5.04292
R309 source.n28 source.n19 5.04292
R310 source.n130 source.n129 5.04292
R311 source.n96 source.n87 5.04292
R312 source.n234 source.n222 4.26717
R313 source.n264 source.n208 4.26717
R314 source.n166 source.n154 4.26717
R315 source.n196 source.n140 4.26717
R316 source.n58 source.n2 4.26717
R317 source.n29 source.n17 4.26717
R318 source.n126 source.n70 4.26717
R319 source.n97 source.n85 4.26717
R320 source.n238 source.n237 3.49141
R321 source.n263 source.n210 3.49141
R322 source.n170 source.n169 3.49141
R323 source.n195 source.n142 3.49141
R324 source.n57 source.n4 3.49141
R325 source.n33 source.n32 3.49141
R326 source.n125 source.n72 3.49141
R327 source.n101 source.n100 3.49141
R328 source.n228 source.n227 2.84303
R329 source.n160 source.n159 2.84303
R330 source.n23 source.n22 2.84303
R331 source.n91 source.n90 2.84303
R332 source.n241 source.n220 2.71565
R333 source.n260 source.n259 2.71565
R334 source.n173 source.n152 2.71565
R335 source.n192 source.n191 2.71565
R336 source.n54 source.n53 2.71565
R337 source.n36 source.n15 2.71565
R338 source.n122 source.n121 2.71565
R339 source.n104 source.n83 2.71565
R340 source.n242 source.n218 1.93989
R341 source.n256 source.n212 1.93989
R342 source.n174 source.n150 1.93989
R343 source.n188 source.n144 1.93989
R344 source.n50 source.n6 1.93989
R345 source.n37 source.n13 1.93989
R346 source.n118 source.n74 1.93989
R347 source.n105 source.n81 1.93989
R348 source.n204 source.t6 1.6505
R349 source.n204 source.t7 1.6505
R350 source.n136 source.t5 1.6505
R351 source.n136 source.t3 1.6505
R352 source.n66 source.t2 1.6505
R353 source.n66 source.t0 1.6505
R354 source.n134 source.t8 1.6505
R355 source.n134 source.t11 1.6505
R356 source.n247 source.n245 1.16414
R357 source.n255 source.n214 1.16414
R358 source.n179 source.n177 1.16414
R359 source.n187 source.n146 1.16414
R360 source.n49 source.n8 1.16414
R361 source.n41 source.n40 1.16414
R362 source.n117 source.n76 1.16414
R363 source.n109 source.n108 1.16414
R364 source.n133 source.n67 0.698776
R365 source.n205 source.n203 0.698776
R366 source.n135 source.n133 0.457397
R367 source.n67 source.n65 0.457397
R368 source.n203 source.n137 0.457397
R369 source.n271 source.n205 0.457397
R370 source.n246 source.n216 0.388379
R371 source.n252 source.n251 0.388379
R372 source.n178 source.n148 0.388379
R373 source.n184 source.n183 0.388379
R374 source.n46 source.n45 0.388379
R375 source.n12 source.n10 0.388379
R376 source.n114 source.n113 0.388379
R377 source.n80 source.n78 0.388379
R378 source source.n272 0.188
R379 source.n228 source.n223 0.155672
R380 source.n235 source.n223 0.155672
R381 source.n236 source.n235 0.155672
R382 source.n236 source.n219 0.155672
R383 source.n243 source.n219 0.155672
R384 source.n244 source.n243 0.155672
R385 source.n244 source.n215 0.155672
R386 source.n253 source.n215 0.155672
R387 source.n254 source.n253 0.155672
R388 source.n254 source.n211 0.155672
R389 source.n261 source.n211 0.155672
R390 source.n262 source.n261 0.155672
R391 source.n262 source.n207 0.155672
R392 source.n269 source.n207 0.155672
R393 source.n160 source.n155 0.155672
R394 source.n167 source.n155 0.155672
R395 source.n168 source.n167 0.155672
R396 source.n168 source.n151 0.155672
R397 source.n175 source.n151 0.155672
R398 source.n176 source.n175 0.155672
R399 source.n176 source.n147 0.155672
R400 source.n185 source.n147 0.155672
R401 source.n186 source.n185 0.155672
R402 source.n186 source.n143 0.155672
R403 source.n193 source.n143 0.155672
R404 source.n194 source.n193 0.155672
R405 source.n194 source.n139 0.155672
R406 source.n201 source.n139 0.155672
R407 source.n63 source.n1 0.155672
R408 source.n56 source.n1 0.155672
R409 source.n56 source.n55 0.155672
R410 source.n55 source.n5 0.155672
R411 source.n48 source.n5 0.155672
R412 source.n48 source.n47 0.155672
R413 source.n47 source.n9 0.155672
R414 source.n39 source.n9 0.155672
R415 source.n39 source.n38 0.155672
R416 source.n38 source.n14 0.155672
R417 source.n31 source.n14 0.155672
R418 source.n31 source.n30 0.155672
R419 source.n30 source.n18 0.155672
R420 source.n23 source.n18 0.155672
R421 source.n131 source.n69 0.155672
R422 source.n124 source.n69 0.155672
R423 source.n124 source.n123 0.155672
R424 source.n123 source.n73 0.155672
R425 source.n116 source.n73 0.155672
R426 source.n116 source.n115 0.155672
R427 source.n115 source.n77 0.155672
R428 source.n107 source.n77 0.155672
R429 source.n107 source.n106 0.155672
R430 source.n106 source.n82 0.155672
R431 source.n99 source.n82 0.155672
R432 source.n99 source.n98 0.155672
R433 source.n98 source.n86 0.155672
R434 source.n91 source.n86 0.155672
R435 drain_right.n60 drain_right.n0 289.615
R436 drain_right.n128 drain_right.n68 289.615
R437 drain_right.n20 drain_right.n19 185
R438 drain_right.n25 drain_right.n24 185
R439 drain_right.n27 drain_right.n26 185
R440 drain_right.n16 drain_right.n15 185
R441 drain_right.n33 drain_right.n32 185
R442 drain_right.n35 drain_right.n34 185
R443 drain_right.n12 drain_right.n11 185
R444 drain_right.n42 drain_right.n41 185
R445 drain_right.n43 drain_right.n10 185
R446 drain_right.n45 drain_right.n44 185
R447 drain_right.n8 drain_right.n7 185
R448 drain_right.n51 drain_right.n50 185
R449 drain_right.n53 drain_right.n52 185
R450 drain_right.n4 drain_right.n3 185
R451 drain_right.n59 drain_right.n58 185
R452 drain_right.n61 drain_right.n60 185
R453 drain_right.n129 drain_right.n128 185
R454 drain_right.n127 drain_right.n126 185
R455 drain_right.n72 drain_right.n71 185
R456 drain_right.n121 drain_right.n120 185
R457 drain_right.n119 drain_right.n118 185
R458 drain_right.n76 drain_right.n75 185
R459 drain_right.n113 drain_right.n112 185
R460 drain_right.n111 drain_right.n78 185
R461 drain_right.n110 drain_right.n109 185
R462 drain_right.n81 drain_right.n79 185
R463 drain_right.n104 drain_right.n103 185
R464 drain_right.n102 drain_right.n101 185
R465 drain_right.n85 drain_right.n84 185
R466 drain_right.n96 drain_right.n95 185
R467 drain_right.n94 drain_right.n93 185
R468 drain_right.n89 drain_right.n88 185
R469 drain_right.n21 drain_right.t3 149.524
R470 drain_right.n90 drain_right.t5 149.524
R471 drain_right.n25 drain_right.n19 104.615
R472 drain_right.n26 drain_right.n25 104.615
R473 drain_right.n26 drain_right.n15 104.615
R474 drain_right.n33 drain_right.n15 104.615
R475 drain_right.n34 drain_right.n33 104.615
R476 drain_right.n34 drain_right.n11 104.615
R477 drain_right.n42 drain_right.n11 104.615
R478 drain_right.n43 drain_right.n42 104.615
R479 drain_right.n44 drain_right.n43 104.615
R480 drain_right.n44 drain_right.n7 104.615
R481 drain_right.n51 drain_right.n7 104.615
R482 drain_right.n52 drain_right.n51 104.615
R483 drain_right.n52 drain_right.n3 104.615
R484 drain_right.n59 drain_right.n3 104.615
R485 drain_right.n60 drain_right.n59 104.615
R486 drain_right.n128 drain_right.n127 104.615
R487 drain_right.n127 drain_right.n71 104.615
R488 drain_right.n120 drain_right.n71 104.615
R489 drain_right.n120 drain_right.n119 104.615
R490 drain_right.n119 drain_right.n75 104.615
R491 drain_right.n112 drain_right.n75 104.615
R492 drain_right.n112 drain_right.n111 104.615
R493 drain_right.n111 drain_right.n110 104.615
R494 drain_right.n110 drain_right.n79 104.615
R495 drain_right.n103 drain_right.n79 104.615
R496 drain_right.n103 drain_right.n102 104.615
R497 drain_right.n102 drain_right.n84 104.615
R498 drain_right.n95 drain_right.n84 104.615
R499 drain_right.n95 drain_right.n94 104.615
R500 drain_right.n94 drain_right.n88 104.615
R501 drain_right.n133 drain_right.n67 60.0094
R502 drain_right.n66 drain_right.n65 59.6114
R503 drain_right.t3 drain_right.n19 52.3082
R504 drain_right.t5 drain_right.n88 52.3082
R505 drain_right.n66 drain_right.n64 46.8242
R506 drain_right.n133 drain_right.n132 46.5369
R507 drain_right drain_right.n66 28.0703
R508 drain_right.n45 drain_right.n10 13.1884
R509 drain_right.n113 drain_right.n78 13.1884
R510 drain_right.n41 drain_right.n40 12.8005
R511 drain_right.n46 drain_right.n8 12.8005
R512 drain_right.n114 drain_right.n76 12.8005
R513 drain_right.n109 drain_right.n80 12.8005
R514 drain_right.n39 drain_right.n12 12.0247
R515 drain_right.n50 drain_right.n49 12.0247
R516 drain_right.n118 drain_right.n117 12.0247
R517 drain_right.n108 drain_right.n81 12.0247
R518 drain_right.n36 drain_right.n35 11.249
R519 drain_right.n53 drain_right.n6 11.249
R520 drain_right.n121 drain_right.n74 11.249
R521 drain_right.n105 drain_right.n104 11.249
R522 drain_right.n32 drain_right.n14 10.4732
R523 drain_right.n54 drain_right.n4 10.4732
R524 drain_right.n122 drain_right.n72 10.4732
R525 drain_right.n101 drain_right.n83 10.4732
R526 drain_right.n21 drain_right.n20 10.2747
R527 drain_right.n90 drain_right.n89 10.2747
R528 drain_right.n31 drain_right.n16 9.69747
R529 drain_right.n58 drain_right.n57 9.69747
R530 drain_right.n126 drain_right.n125 9.69747
R531 drain_right.n100 drain_right.n85 9.69747
R532 drain_right.n64 drain_right.n63 9.45567
R533 drain_right.n132 drain_right.n131 9.45567
R534 drain_right.n63 drain_right.n62 9.3005
R535 drain_right.n2 drain_right.n1 9.3005
R536 drain_right.n57 drain_right.n56 9.3005
R537 drain_right.n55 drain_right.n54 9.3005
R538 drain_right.n6 drain_right.n5 9.3005
R539 drain_right.n49 drain_right.n48 9.3005
R540 drain_right.n47 drain_right.n46 9.3005
R541 drain_right.n23 drain_right.n22 9.3005
R542 drain_right.n18 drain_right.n17 9.3005
R543 drain_right.n29 drain_right.n28 9.3005
R544 drain_right.n31 drain_right.n30 9.3005
R545 drain_right.n14 drain_right.n13 9.3005
R546 drain_right.n37 drain_right.n36 9.3005
R547 drain_right.n39 drain_right.n38 9.3005
R548 drain_right.n40 drain_right.n9 9.3005
R549 drain_right.n92 drain_right.n91 9.3005
R550 drain_right.n87 drain_right.n86 9.3005
R551 drain_right.n98 drain_right.n97 9.3005
R552 drain_right.n100 drain_right.n99 9.3005
R553 drain_right.n83 drain_right.n82 9.3005
R554 drain_right.n106 drain_right.n105 9.3005
R555 drain_right.n108 drain_right.n107 9.3005
R556 drain_right.n80 drain_right.n77 9.3005
R557 drain_right.n131 drain_right.n130 9.3005
R558 drain_right.n70 drain_right.n69 9.3005
R559 drain_right.n125 drain_right.n124 9.3005
R560 drain_right.n123 drain_right.n122 9.3005
R561 drain_right.n74 drain_right.n73 9.3005
R562 drain_right.n117 drain_right.n116 9.3005
R563 drain_right.n115 drain_right.n114 9.3005
R564 drain_right.n28 drain_right.n27 8.92171
R565 drain_right.n61 drain_right.n2 8.92171
R566 drain_right.n129 drain_right.n70 8.92171
R567 drain_right.n97 drain_right.n96 8.92171
R568 drain_right.n24 drain_right.n18 8.14595
R569 drain_right.n62 drain_right.n0 8.14595
R570 drain_right.n130 drain_right.n68 8.14595
R571 drain_right.n93 drain_right.n87 8.14595
R572 drain_right.n23 drain_right.n20 7.3702
R573 drain_right.n92 drain_right.n89 7.3702
R574 drain_right drain_right.n133 5.88166
R575 drain_right.n24 drain_right.n23 5.81868
R576 drain_right.n64 drain_right.n0 5.81868
R577 drain_right.n132 drain_right.n68 5.81868
R578 drain_right.n93 drain_right.n92 5.81868
R579 drain_right.n27 drain_right.n18 5.04292
R580 drain_right.n62 drain_right.n61 5.04292
R581 drain_right.n130 drain_right.n129 5.04292
R582 drain_right.n96 drain_right.n87 5.04292
R583 drain_right.n28 drain_right.n16 4.26717
R584 drain_right.n58 drain_right.n2 4.26717
R585 drain_right.n126 drain_right.n70 4.26717
R586 drain_right.n97 drain_right.n85 4.26717
R587 drain_right.n32 drain_right.n31 3.49141
R588 drain_right.n57 drain_right.n4 3.49141
R589 drain_right.n125 drain_right.n72 3.49141
R590 drain_right.n101 drain_right.n100 3.49141
R591 drain_right.n22 drain_right.n21 2.84303
R592 drain_right.n91 drain_right.n90 2.84303
R593 drain_right.n35 drain_right.n14 2.71565
R594 drain_right.n54 drain_right.n53 2.71565
R595 drain_right.n122 drain_right.n121 2.71565
R596 drain_right.n104 drain_right.n83 2.71565
R597 drain_right.n36 drain_right.n12 1.93989
R598 drain_right.n50 drain_right.n6 1.93989
R599 drain_right.n118 drain_right.n74 1.93989
R600 drain_right.n105 drain_right.n81 1.93989
R601 drain_right.n65 drain_right.t2 1.6505
R602 drain_right.n65 drain_right.t4 1.6505
R603 drain_right.n67 drain_right.t1 1.6505
R604 drain_right.n67 drain_right.t0 1.6505
R605 drain_right.n41 drain_right.n39 1.16414
R606 drain_right.n49 drain_right.n8 1.16414
R607 drain_right.n117 drain_right.n76 1.16414
R608 drain_right.n109 drain_right.n108 1.16414
R609 drain_right.n40 drain_right.n10 0.388379
R610 drain_right.n46 drain_right.n45 0.388379
R611 drain_right.n114 drain_right.n113 0.388379
R612 drain_right.n80 drain_right.n78 0.388379
R613 drain_right.n22 drain_right.n17 0.155672
R614 drain_right.n29 drain_right.n17 0.155672
R615 drain_right.n30 drain_right.n29 0.155672
R616 drain_right.n30 drain_right.n13 0.155672
R617 drain_right.n37 drain_right.n13 0.155672
R618 drain_right.n38 drain_right.n37 0.155672
R619 drain_right.n38 drain_right.n9 0.155672
R620 drain_right.n47 drain_right.n9 0.155672
R621 drain_right.n48 drain_right.n47 0.155672
R622 drain_right.n48 drain_right.n5 0.155672
R623 drain_right.n55 drain_right.n5 0.155672
R624 drain_right.n56 drain_right.n55 0.155672
R625 drain_right.n56 drain_right.n1 0.155672
R626 drain_right.n63 drain_right.n1 0.155672
R627 drain_right.n131 drain_right.n69 0.155672
R628 drain_right.n124 drain_right.n69 0.155672
R629 drain_right.n124 drain_right.n123 0.155672
R630 drain_right.n123 drain_right.n73 0.155672
R631 drain_right.n116 drain_right.n73 0.155672
R632 drain_right.n116 drain_right.n115 0.155672
R633 drain_right.n115 drain_right.n77 0.155672
R634 drain_right.n107 drain_right.n77 0.155672
R635 drain_right.n107 drain_right.n106 0.155672
R636 drain_right.n106 drain_right.n82 0.155672
R637 drain_right.n99 drain_right.n82 0.155672
R638 drain_right.n99 drain_right.n98 0.155672
R639 drain_right.n98 drain_right.n86 0.155672
R640 drain_right.n91 drain_right.n86 0.155672
R641 plus.n0 plus.t1 1643.55
R642 plus.n2 plus.t4 1643.55
R643 plus.n4 plus.t3 1643.55
R644 plus.n6 plus.t2 1643.55
R645 plus.n1 plus.t0 1602.65
R646 plus.n5 plus.t5 1602.65
R647 plus.n3 plus.n0 161.489
R648 plus.n7 plus.n4 161.489
R649 plus.n3 plus.n2 161.3
R650 plus.n7 plus.n6 161.3
R651 plus.n1 plus.n0 36.5157
R652 plus.n2 plus.n1 36.5157
R653 plus.n6 plus.n5 36.5157
R654 plus.n5 plus.n4 36.5157
R655 plus plus.n7 27.2585
R656 plus plus.n3 12.0819
R657 drain_left.n60 drain_left.n0 289.615
R658 drain_left.n127 drain_left.n67 289.615
R659 drain_left.n20 drain_left.n19 185
R660 drain_left.n25 drain_left.n24 185
R661 drain_left.n27 drain_left.n26 185
R662 drain_left.n16 drain_left.n15 185
R663 drain_left.n33 drain_left.n32 185
R664 drain_left.n35 drain_left.n34 185
R665 drain_left.n12 drain_left.n11 185
R666 drain_left.n42 drain_left.n41 185
R667 drain_left.n43 drain_left.n10 185
R668 drain_left.n45 drain_left.n44 185
R669 drain_left.n8 drain_left.n7 185
R670 drain_left.n51 drain_left.n50 185
R671 drain_left.n53 drain_left.n52 185
R672 drain_left.n4 drain_left.n3 185
R673 drain_left.n59 drain_left.n58 185
R674 drain_left.n61 drain_left.n60 185
R675 drain_left.n128 drain_left.n127 185
R676 drain_left.n126 drain_left.n125 185
R677 drain_left.n71 drain_left.n70 185
R678 drain_left.n120 drain_left.n119 185
R679 drain_left.n118 drain_left.n117 185
R680 drain_left.n75 drain_left.n74 185
R681 drain_left.n112 drain_left.n111 185
R682 drain_left.n110 drain_left.n77 185
R683 drain_left.n109 drain_left.n108 185
R684 drain_left.n80 drain_left.n78 185
R685 drain_left.n103 drain_left.n102 185
R686 drain_left.n101 drain_left.n100 185
R687 drain_left.n84 drain_left.n83 185
R688 drain_left.n95 drain_left.n94 185
R689 drain_left.n93 drain_left.n92 185
R690 drain_left.n88 drain_left.n87 185
R691 drain_left.n21 drain_left.t3 149.524
R692 drain_left.n89 drain_left.t4 149.524
R693 drain_left.n25 drain_left.n19 104.615
R694 drain_left.n26 drain_left.n25 104.615
R695 drain_left.n26 drain_left.n15 104.615
R696 drain_left.n33 drain_left.n15 104.615
R697 drain_left.n34 drain_left.n33 104.615
R698 drain_left.n34 drain_left.n11 104.615
R699 drain_left.n42 drain_left.n11 104.615
R700 drain_left.n43 drain_left.n42 104.615
R701 drain_left.n44 drain_left.n43 104.615
R702 drain_left.n44 drain_left.n7 104.615
R703 drain_left.n51 drain_left.n7 104.615
R704 drain_left.n52 drain_left.n51 104.615
R705 drain_left.n52 drain_left.n3 104.615
R706 drain_left.n59 drain_left.n3 104.615
R707 drain_left.n60 drain_left.n59 104.615
R708 drain_left.n127 drain_left.n126 104.615
R709 drain_left.n126 drain_left.n70 104.615
R710 drain_left.n119 drain_left.n70 104.615
R711 drain_left.n119 drain_left.n118 104.615
R712 drain_left.n118 drain_left.n74 104.615
R713 drain_left.n111 drain_left.n74 104.615
R714 drain_left.n111 drain_left.n110 104.615
R715 drain_left.n110 drain_left.n109 104.615
R716 drain_left.n109 drain_left.n78 104.615
R717 drain_left.n102 drain_left.n78 104.615
R718 drain_left.n102 drain_left.n101 104.615
R719 drain_left.n101 drain_left.n83 104.615
R720 drain_left.n94 drain_left.n83 104.615
R721 drain_left.n94 drain_left.n93 104.615
R722 drain_left.n93 drain_left.n87 104.615
R723 drain_left.n66 drain_left.n65 59.6114
R724 drain_left.n133 drain_left.n132 59.5525
R725 drain_left.t3 drain_left.n19 52.3082
R726 drain_left.t4 drain_left.n87 52.3082
R727 drain_left.n133 drain_left.n131 46.9938
R728 drain_left.n66 drain_left.n64 46.8242
R729 drain_left drain_left.n66 28.6235
R730 drain_left.n45 drain_left.n10 13.1884
R731 drain_left.n112 drain_left.n77 13.1884
R732 drain_left.n41 drain_left.n40 12.8005
R733 drain_left.n46 drain_left.n8 12.8005
R734 drain_left.n113 drain_left.n75 12.8005
R735 drain_left.n108 drain_left.n79 12.8005
R736 drain_left.n39 drain_left.n12 12.0247
R737 drain_left.n50 drain_left.n49 12.0247
R738 drain_left.n117 drain_left.n116 12.0247
R739 drain_left.n107 drain_left.n80 12.0247
R740 drain_left.n36 drain_left.n35 11.249
R741 drain_left.n53 drain_left.n6 11.249
R742 drain_left.n120 drain_left.n73 11.249
R743 drain_left.n104 drain_left.n103 11.249
R744 drain_left.n32 drain_left.n14 10.4732
R745 drain_left.n54 drain_left.n4 10.4732
R746 drain_left.n121 drain_left.n71 10.4732
R747 drain_left.n100 drain_left.n82 10.4732
R748 drain_left.n21 drain_left.n20 10.2747
R749 drain_left.n89 drain_left.n88 10.2747
R750 drain_left.n31 drain_left.n16 9.69747
R751 drain_left.n58 drain_left.n57 9.69747
R752 drain_left.n125 drain_left.n124 9.69747
R753 drain_left.n99 drain_left.n84 9.69747
R754 drain_left.n64 drain_left.n63 9.45567
R755 drain_left.n131 drain_left.n130 9.45567
R756 drain_left.n63 drain_left.n62 9.3005
R757 drain_left.n2 drain_left.n1 9.3005
R758 drain_left.n57 drain_left.n56 9.3005
R759 drain_left.n55 drain_left.n54 9.3005
R760 drain_left.n6 drain_left.n5 9.3005
R761 drain_left.n49 drain_left.n48 9.3005
R762 drain_left.n47 drain_left.n46 9.3005
R763 drain_left.n23 drain_left.n22 9.3005
R764 drain_left.n18 drain_left.n17 9.3005
R765 drain_left.n29 drain_left.n28 9.3005
R766 drain_left.n31 drain_left.n30 9.3005
R767 drain_left.n14 drain_left.n13 9.3005
R768 drain_left.n37 drain_left.n36 9.3005
R769 drain_left.n39 drain_left.n38 9.3005
R770 drain_left.n40 drain_left.n9 9.3005
R771 drain_left.n91 drain_left.n90 9.3005
R772 drain_left.n86 drain_left.n85 9.3005
R773 drain_left.n97 drain_left.n96 9.3005
R774 drain_left.n99 drain_left.n98 9.3005
R775 drain_left.n82 drain_left.n81 9.3005
R776 drain_left.n105 drain_left.n104 9.3005
R777 drain_left.n107 drain_left.n106 9.3005
R778 drain_left.n79 drain_left.n76 9.3005
R779 drain_left.n130 drain_left.n129 9.3005
R780 drain_left.n69 drain_left.n68 9.3005
R781 drain_left.n124 drain_left.n123 9.3005
R782 drain_left.n122 drain_left.n121 9.3005
R783 drain_left.n73 drain_left.n72 9.3005
R784 drain_left.n116 drain_left.n115 9.3005
R785 drain_left.n114 drain_left.n113 9.3005
R786 drain_left.n28 drain_left.n27 8.92171
R787 drain_left.n61 drain_left.n2 8.92171
R788 drain_left.n128 drain_left.n69 8.92171
R789 drain_left.n96 drain_left.n95 8.92171
R790 drain_left.n24 drain_left.n18 8.14595
R791 drain_left.n62 drain_left.n0 8.14595
R792 drain_left.n129 drain_left.n67 8.14595
R793 drain_left.n92 drain_left.n86 8.14595
R794 drain_left.n23 drain_left.n20 7.3702
R795 drain_left.n91 drain_left.n88 7.3702
R796 drain_left drain_left.n133 6.11011
R797 drain_left.n24 drain_left.n23 5.81868
R798 drain_left.n64 drain_left.n0 5.81868
R799 drain_left.n131 drain_left.n67 5.81868
R800 drain_left.n92 drain_left.n91 5.81868
R801 drain_left.n27 drain_left.n18 5.04292
R802 drain_left.n62 drain_left.n61 5.04292
R803 drain_left.n129 drain_left.n128 5.04292
R804 drain_left.n95 drain_left.n86 5.04292
R805 drain_left.n28 drain_left.n16 4.26717
R806 drain_left.n58 drain_left.n2 4.26717
R807 drain_left.n125 drain_left.n69 4.26717
R808 drain_left.n96 drain_left.n84 4.26717
R809 drain_left.n32 drain_left.n31 3.49141
R810 drain_left.n57 drain_left.n4 3.49141
R811 drain_left.n124 drain_left.n71 3.49141
R812 drain_left.n100 drain_left.n99 3.49141
R813 drain_left.n22 drain_left.n21 2.84303
R814 drain_left.n90 drain_left.n89 2.84303
R815 drain_left.n35 drain_left.n14 2.71565
R816 drain_left.n54 drain_left.n53 2.71565
R817 drain_left.n121 drain_left.n120 2.71565
R818 drain_left.n103 drain_left.n82 2.71565
R819 drain_left.n36 drain_left.n12 1.93989
R820 drain_left.n50 drain_left.n6 1.93989
R821 drain_left.n117 drain_left.n73 1.93989
R822 drain_left.n104 drain_left.n80 1.93989
R823 drain_left.n65 drain_left.t0 1.6505
R824 drain_left.n65 drain_left.t2 1.6505
R825 drain_left.n132 drain_left.t5 1.6505
R826 drain_left.n132 drain_left.t1 1.6505
R827 drain_left.n41 drain_left.n39 1.16414
R828 drain_left.n49 drain_left.n8 1.16414
R829 drain_left.n116 drain_left.n75 1.16414
R830 drain_left.n108 drain_left.n107 1.16414
R831 drain_left.n40 drain_left.n10 0.388379
R832 drain_left.n46 drain_left.n45 0.388379
R833 drain_left.n113 drain_left.n112 0.388379
R834 drain_left.n79 drain_left.n77 0.388379
R835 drain_left.n22 drain_left.n17 0.155672
R836 drain_left.n29 drain_left.n17 0.155672
R837 drain_left.n30 drain_left.n29 0.155672
R838 drain_left.n30 drain_left.n13 0.155672
R839 drain_left.n37 drain_left.n13 0.155672
R840 drain_left.n38 drain_left.n37 0.155672
R841 drain_left.n38 drain_left.n9 0.155672
R842 drain_left.n47 drain_left.n9 0.155672
R843 drain_left.n48 drain_left.n47 0.155672
R844 drain_left.n48 drain_left.n5 0.155672
R845 drain_left.n55 drain_left.n5 0.155672
R846 drain_left.n56 drain_left.n55 0.155672
R847 drain_left.n56 drain_left.n1 0.155672
R848 drain_left.n63 drain_left.n1 0.155672
R849 drain_left.n130 drain_left.n68 0.155672
R850 drain_left.n123 drain_left.n68 0.155672
R851 drain_left.n123 drain_left.n122 0.155672
R852 drain_left.n122 drain_left.n72 0.155672
R853 drain_left.n115 drain_left.n72 0.155672
R854 drain_left.n115 drain_left.n114 0.155672
R855 drain_left.n114 drain_left.n76 0.155672
R856 drain_left.n106 drain_left.n76 0.155672
R857 drain_left.n106 drain_left.n105 0.155672
R858 drain_left.n105 drain_left.n81 0.155672
R859 drain_left.n98 drain_left.n81 0.155672
R860 drain_left.n98 drain_left.n97 0.155672
R861 drain_left.n97 drain_left.n85 0.155672
R862 drain_left.n90 drain_left.n85 0.155672
C0 plus drain_right 0.261274f
C1 plus source 1.66161f
C2 minus drain_left 0.170484f
C3 drain_left drain_right 0.535026f
C4 drain_left source 16.404099f
C5 plus drain_left 2.27627f
C6 minus drain_right 2.1734f
C7 minus source 1.64687f
C8 plus minus 4.57614f
C9 source drain_right 16.391098f
C10 drain_right a_n1140_n3288# 6.52569f
C11 drain_left a_n1140_n3288# 6.70626f
C12 source a_n1140_n3288# 5.992964f
C13 minus a_n1140_n3288# 4.365132f
C14 plus a_n1140_n3288# 6.09021f
C15 drain_left.n0 a_n1140_n3288# 0.040612f
C16 drain_left.n1 a_n1140_n3288# 0.030659f
C17 drain_left.n2 a_n1140_n3288# 0.016475f
C18 drain_left.n3 a_n1140_n3288# 0.03894f
C19 drain_left.n4 a_n1140_n3288# 0.017444f
C20 drain_left.n5 a_n1140_n3288# 0.030659f
C21 drain_left.n6 a_n1140_n3288# 0.016475f
C22 drain_left.n7 a_n1140_n3288# 0.03894f
C23 drain_left.n8 a_n1140_n3288# 0.017444f
C24 drain_left.n9 a_n1140_n3288# 0.030659f
C25 drain_left.n10 a_n1140_n3288# 0.016959f
C26 drain_left.n11 a_n1140_n3288# 0.03894f
C27 drain_left.n12 a_n1140_n3288# 0.017444f
C28 drain_left.n13 a_n1140_n3288# 0.030659f
C29 drain_left.n14 a_n1140_n3288# 0.016475f
C30 drain_left.n15 a_n1140_n3288# 0.03894f
C31 drain_left.n16 a_n1140_n3288# 0.017444f
C32 drain_left.n17 a_n1140_n3288# 0.030659f
C33 drain_left.n18 a_n1140_n3288# 0.016475f
C34 drain_left.n19 a_n1140_n3288# 0.029205f
C35 drain_left.n20 a_n1140_n3288# 0.027528f
C36 drain_left.t3 a_n1140_n3288# 0.065768f
C37 drain_left.n21 a_n1140_n3288# 0.221048f
C38 drain_left.n22 a_n1140_n3288# 1.54669f
C39 drain_left.n23 a_n1140_n3288# 0.016475f
C40 drain_left.n24 a_n1140_n3288# 0.017444f
C41 drain_left.n25 a_n1140_n3288# 0.03894f
C42 drain_left.n26 a_n1140_n3288# 0.03894f
C43 drain_left.n27 a_n1140_n3288# 0.017444f
C44 drain_left.n28 a_n1140_n3288# 0.016475f
C45 drain_left.n29 a_n1140_n3288# 0.030659f
C46 drain_left.n30 a_n1140_n3288# 0.030659f
C47 drain_left.n31 a_n1140_n3288# 0.016475f
C48 drain_left.n32 a_n1140_n3288# 0.017444f
C49 drain_left.n33 a_n1140_n3288# 0.03894f
C50 drain_left.n34 a_n1140_n3288# 0.03894f
C51 drain_left.n35 a_n1140_n3288# 0.017444f
C52 drain_left.n36 a_n1140_n3288# 0.016475f
C53 drain_left.n37 a_n1140_n3288# 0.030659f
C54 drain_left.n38 a_n1140_n3288# 0.030659f
C55 drain_left.n39 a_n1140_n3288# 0.016475f
C56 drain_left.n40 a_n1140_n3288# 0.016475f
C57 drain_left.n41 a_n1140_n3288# 0.017444f
C58 drain_left.n42 a_n1140_n3288# 0.03894f
C59 drain_left.n43 a_n1140_n3288# 0.03894f
C60 drain_left.n44 a_n1140_n3288# 0.03894f
C61 drain_left.n45 a_n1140_n3288# 0.016959f
C62 drain_left.n46 a_n1140_n3288# 0.016475f
C63 drain_left.n47 a_n1140_n3288# 0.030659f
C64 drain_left.n48 a_n1140_n3288# 0.030659f
C65 drain_left.n49 a_n1140_n3288# 0.016475f
C66 drain_left.n50 a_n1140_n3288# 0.017444f
C67 drain_left.n51 a_n1140_n3288# 0.03894f
C68 drain_left.n52 a_n1140_n3288# 0.03894f
C69 drain_left.n53 a_n1140_n3288# 0.017444f
C70 drain_left.n54 a_n1140_n3288# 0.016475f
C71 drain_left.n55 a_n1140_n3288# 0.030659f
C72 drain_left.n56 a_n1140_n3288# 0.030659f
C73 drain_left.n57 a_n1140_n3288# 0.016475f
C74 drain_left.n58 a_n1140_n3288# 0.017444f
C75 drain_left.n59 a_n1140_n3288# 0.03894f
C76 drain_left.n60 a_n1140_n3288# 0.07991f
C77 drain_left.n61 a_n1140_n3288# 0.017444f
C78 drain_left.n62 a_n1140_n3288# 0.016475f
C79 drain_left.n63 a_n1140_n3288# 0.065841f
C80 drain_left.n64 a_n1140_n3288# 0.065849f
C81 drain_left.t0 a_n1140_n3288# 0.290732f
C82 drain_left.t2 a_n1140_n3288# 0.290732f
C83 drain_left.n65 a_n1140_n3288# 2.58739f
C84 drain_left.n66 a_n1140_n3288# 1.68114f
C85 drain_left.n67 a_n1140_n3288# 0.040612f
C86 drain_left.n68 a_n1140_n3288# 0.030659f
C87 drain_left.n69 a_n1140_n3288# 0.016475f
C88 drain_left.n70 a_n1140_n3288# 0.03894f
C89 drain_left.n71 a_n1140_n3288# 0.017444f
C90 drain_left.n72 a_n1140_n3288# 0.030659f
C91 drain_left.n73 a_n1140_n3288# 0.016475f
C92 drain_left.n74 a_n1140_n3288# 0.03894f
C93 drain_left.n75 a_n1140_n3288# 0.017444f
C94 drain_left.n76 a_n1140_n3288# 0.030659f
C95 drain_left.n77 a_n1140_n3288# 0.016959f
C96 drain_left.n78 a_n1140_n3288# 0.03894f
C97 drain_left.n79 a_n1140_n3288# 0.016475f
C98 drain_left.n80 a_n1140_n3288# 0.017444f
C99 drain_left.n81 a_n1140_n3288# 0.030659f
C100 drain_left.n82 a_n1140_n3288# 0.016475f
C101 drain_left.n83 a_n1140_n3288# 0.03894f
C102 drain_left.n84 a_n1140_n3288# 0.017444f
C103 drain_left.n85 a_n1140_n3288# 0.030659f
C104 drain_left.n86 a_n1140_n3288# 0.016475f
C105 drain_left.n87 a_n1140_n3288# 0.029205f
C106 drain_left.n88 a_n1140_n3288# 0.027528f
C107 drain_left.t4 a_n1140_n3288# 0.065768f
C108 drain_left.n89 a_n1140_n3288# 0.221048f
C109 drain_left.n90 a_n1140_n3288# 1.54669f
C110 drain_left.n91 a_n1140_n3288# 0.016475f
C111 drain_left.n92 a_n1140_n3288# 0.017444f
C112 drain_left.n93 a_n1140_n3288# 0.03894f
C113 drain_left.n94 a_n1140_n3288# 0.03894f
C114 drain_left.n95 a_n1140_n3288# 0.017444f
C115 drain_left.n96 a_n1140_n3288# 0.016475f
C116 drain_left.n97 a_n1140_n3288# 0.030659f
C117 drain_left.n98 a_n1140_n3288# 0.030659f
C118 drain_left.n99 a_n1140_n3288# 0.016475f
C119 drain_left.n100 a_n1140_n3288# 0.017444f
C120 drain_left.n101 a_n1140_n3288# 0.03894f
C121 drain_left.n102 a_n1140_n3288# 0.03894f
C122 drain_left.n103 a_n1140_n3288# 0.017444f
C123 drain_left.n104 a_n1140_n3288# 0.016475f
C124 drain_left.n105 a_n1140_n3288# 0.030659f
C125 drain_left.n106 a_n1140_n3288# 0.030659f
C126 drain_left.n107 a_n1140_n3288# 0.016475f
C127 drain_left.n108 a_n1140_n3288# 0.017444f
C128 drain_left.n109 a_n1140_n3288# 0.03894f
C129 drain_left.n110 a_n1140_n3288# 0.03894f
C130 drain_left.n111 a_n1140_n3288# 0.03894f
C131 drain_left.n112 a_n1140_n3288# 0.016959f
C132 drain_left.n113 a_n1140_n3288# 0.016475f
C133 drain_left.n114 a_n1140_n3288# 0.030659f
C134 drain_left.n115 a_n1140_n3288# 0.030659f
C135 drain_left.n116 a_n1140_n3288# 0.016475f
C136 drain_left.n117 a_n1140_n3288# 0.017444f
C137 drain_left.n118 a_n1140_n3288# 0.03894f
C138 drain_left.n119 a_n1140_n3288# 0.03894f
C139 drain_left.n120 a_n1140_n3288# 0.017444f
C140 drain_left.n121 a_n1140_n3288# 0.016475f
C141 drain_left.n122 a_n1140_n3288# 0.030659f
C142 drain_left.n123 a_n1140_n3288# 0.030659f
C143 drain_left.n124 a_n1140_n3288# 0.016475f
C144 drain_left.n125 a_n1140_n3288# 0.017444f
C145 drain_left.n126 a_n1140_n3288# 0.03894f
C146 drain_left.n127 a_n1140_n3288# 0.07991f
C147 drain_left.n128 a_n1140_n3288# 0.017444f
C148 drain_left.n129 a_n1140_n3288# 0.016475f
C149 drain_left.n130 a_n1140_n3288# 0.065841f
C150 drain_left.n131 a_n1140_n3288# 0.0663f
C151 drain_left.t5 a_n1140_n3288# 0.290732f
C152 drain_left.t1 a_n1140_n3288# 0.290732f
C153 drain_left.n132 a_n1140_n3288# 2.58706f
C154 drain_left.n133 a_n1140_n3288# 0.698808f
C155 plus.t1 a_n1140_n3288# 0.349665f
C156 plus.n0 a_n1140_n3288# 0.156337f
C157 plus.t0 a_n1140_n3288# 0.346134f
C158 plus.n1 a_n1140_n3288# 0.142554f
C159 plus.t4 a_n1140_n3288# 0.349665f
C160 plus.n2 a_n1140_n3288# 0.156268f
C161 plus.n3 a_n1140_n3288# 0.622601f
C162 plus.t3 a_n1140_n3288# 0.349665f
C163 plus.n4 a_n1140_n3288# 0.156337f
C164 plus.t2 a_n1140_n3288# 0.349665f
C165 plus.t5 a_n1140_n3288# 0.346134f
C166 plus.n5 a_n1140_n3288# 0.142554f
C167 plus.n6 a_n1140_n3288# 0.156268f
C168 plus.n7 a_n1140_n3288# 1.39043f
C169 drain_right.n0 a_n1140_n3288# 0.040655f
C170 drain_right.n1 a_n1140_n3288# 0.030692f
C171 drain_right.n2 a_n1140_n3288# 0.016493f
C172 drain_right.n3 a_n1140_n3288# 0.038982f
C173 drain_right.n4 a_n1140_n3288# 0.017463f
C174 drain_right.n5 a_n1140_n3288# 0.030692f
C175 drain_right.n6 a_n1140_n3288# 0.016493f
C176 drain_right.n7 a_n1140_n3288# 0.038982f
C177 drain_right.n8 a_n1140_n3288# 0.017463f
C178 drain_right.n9 a_n1140_n3288# 0.030692f
C179 drain_right.n10 a_n1140_n3288# 0.016978f
C180 drain_right.n11 a_n1140_n3288# 0.038982f
C181 drain_right.n12 a_n1140_n3288# 0.017463f
C182 drain_right.n13 a_n1140_n3288# 0.030692f
C183 drain_right.n14 a_n1140_n3288# 0.016493f
C184 drain_right.n15 a_n1140_n3288# 0.038982f
C185 drain_right.n16 a_n1140_n3288# 0.017463f
C186 drain_right.n17 a_n1140_n3288# 0.030692f
C187 drain_right.n18 a_n1140_n3288# 0.016493f
C188 drain_right.n19 a_n1140_n3288# 0.029237f
C189 drain_right.n20 a_n1140_n3288# 0.027557f
C190 drain_right.t3 a_n1140_n3288# 0.065838f
C191 drain_right.n21 a_n1140_n3288# 0.221285f
C192 drain_right.n22 a_n1140_n3288# 1.54835f
C193 drain_right.n23 a_n1140_n3288# 0.016493f
C194 drain_right.n24 a_n1140_n3288# 0.017463f
C195 drain_right.n25 a_n1140_n3288# 0.038982f
C196 drain_right.n26 a_n1140_n3288# 0.038982f
C197 drain_right.n27 a_n1140_n3288# 0.017463f
C198 drain_right.n28 a_n1140_n3288# 0.016493f
C199 drain_right.n29 a_n1140_n3288# 0.030692f
C200 drain_right.n30 a_n1140_n3288# 0.030692f
C201 drain_right.n31 a_n1140_n3288# 0.016493f
C202 drain_right.n32 a_n1140_n3288# 0.017463f
C203 drain_right.n33 a_n1140_n3288# 0.038982f
C204 drain_right.n34 a_n1140_n3288# 0.038982f
C205 drain_right.n35 a_n1140_n3288# 0.017463f
C206 drain_right.n36 a_n1140_n3288# 0.016493f
C207 drain_right.n37 a_n1140_n3288# 0.030692f
C208 drain_right.n38 a_n1140_n3288# 0.030692f
C209 drain_right.n39 a_n1140_n3288# 0.016493f
C210 drain_right.n40 a_n1140_n3288# 0.016493f
C211 drain_right.n41 a_n1140_n3288# 0.017463f
C212 drain_right.n42 a_n1140_n3288# 0.038982f
C213 drain_right.n43 a_n1140_n3288# 0.038982f
C214 drain_right.n44 a_n1140_n3288# 0.038982f
C215 drain_right.n45 a_n1140_n3288# 0.016978f
C216 drain_right.n46 a_n1140_n3288# 0.016493f
C217 drain_right.n47 a_n1140_n3288# 0.030692f
C218 drain_right.n48 a_n1140_n3288# 0.030692f
C219 drain_right.n49 a_n1140_n3288# 0.016493f
C220 drain_right.n50 a_n1140_n3288# 0.017463f
C221 drain_right.n51 a_n1140_n3288# 0.038982f
C222 drain_right.n52 a_n1140_n3288# 0.038982f
C223 drain_right.n53 a_n1140_n3288# 0.017463f
C224 drain_right.n54 a_n1140_n3288# 0.016493f
C225 drain_right.n55 a_n1140_n3288# 0.030692f
C226 drain_right.n56 a_n1140_n3288# 0.030692f
C227 drain_right.n57 a_n1140_n3288# 0.016493f
C228 drain_right.n58 a_n1140_n3288# 0.017463f
C229 drain_right.n59 a_n1140_n3288# 0.038982f
C230 drain_right.n60 a_n1140_n3288# 0.079996f
C231 drain_right.n61 a_n1140_n3288# 0.017463f
C232 drain_right.n62 a_n1140_n3288# 0.016493f
C233 drain_right.n63 a_n1140_n3288# 0.065911f
C234 drain_right.n64 a_n1140_n3288# 0.065919f
C235 drain_right.t2 a_n1140_n3288# 0.291044f
C236 drain_right.t4 a_n1140_n3288# 0.291044f
C237 drain_right.n65 a_n1140_n3288# 2.59017f
C238 drain_right.n66 a_n1140_n3288# 1.61843f
C239 drain_right.t1 a_n1140_n3288# 0.291044f
C240 drain_right.t0 a_n1140_n3288# 0.291044f
C241 drain_right.n67 a_n1140_n3288# 2.59258f
C242 drain_right.n68 a_n1140_n3288# 0.040655f
C243 drain_right.n69 a_n1140_n3288# 0.030692f
C244 drain_right.n70 a_n1140_n3288# 0.016493f
C245 drain_right.n71 a_n1140_n3288# 0.038982f
C246 drain_right.n72 a_n1140_n3288# 0.017463f
C247 drain_right.n73 a_n1140_n3288# 0.030692f
C248 drain_right.n74 a_n1140_n3288# 0.016493f
C249 drain_right.n75 a_n1140_n3288# 0.038982f
C250 drain_right.n76 a_n1140_n3288# 0.017463f
C251 drain_right.n77 a_n1140_n3288# 0.030692f
C252 drain_right.n78 a_n1140_n3288# 0.016978f
C253 drain_right.n79 a_n1140_n3288# 0.038982f
C254 drain_right.n80 a_n1140_n3288# 0.016493f
C255 drain_right.n81 a_n1140_n3288# 0.017463f
C256 drain_right.n82 a_n1140_n3288# 0.030692f
C257 drain_right.n83 a_n1140_n3288# 0.016493f
C258 drain_right.n84 a_n1140_n3288# 0.038982f
C259 drain_right.n85 a_n1140_n3288# 0.017463f
C260 drain_right.n86 a_n1140_n3288# 0.030692f
C261 drain_right.n87 a_n1140_n3288# 0.016493f
C262 drain_right.n88 a_n1140_n3288# 0.029237f
C263 drain_right.n89 a_n1140_n3288# 0.027557f
C264 drain_right.t5 a_n1140_n3288# 0.065838f
C265 drain_right.n90 a_n1140_n3288# 0.221285f
C266 drain_right.n91 a_n1140_n3288# 1.54835f
C267 drain_right.n92 a_n1140_n3288# 0.016493f
C268 drain_right.n93 a_n1140_n3288# 0.017463f
C269 drain_right.n94 a_n1140_n3288# 0.038982f
C270 drain_right.n95 a_n1140_n3288# 0.038982f
C271 drain_right.n96 a_n1140_n3288# 0.017463f
C272 drain_right.n97 a_n1140_n3288# 0.016493f
C273 drain_right.n98 a_n1140_n3288# 0.030692f
C274 drain_right.n99 a_n1140_n3288# 0.030692f
C275 drain_right.n100 a_n1140_n3288# 0.016493f
C276 drain_right.n101 a_n1140_n3288# 0.017463f
C277 drain_right.n102 a_n1140_n3288# 0.038982f
C278 drain_right.n103 a_n1140_n3288# 0.038982f
C279 drain_right.n104 a_n1140_n3288# 0.017463f
C280 drain_right.n105 a_n1140_n3288# 0.016493f
C281 drain_right.n106 a_n1140_n3288# 0.030692f
C282 drain_right.n107 a_n1140_n3288# 0.030692f
C283 drain_right.n108 a_n1140_n3288# 0.016493f
C284 drain_right.n109 a_n1140_n3288# 0.017463f
C285 drain_right.n110 a_n1140_n3288# 0.038982f
C286 drain_right.n111 a_n1140_n3288# 0.038982f
C287 drain_right.n112 a_n1140_n3288# 0.038982f
C288 drain_right.n113 a_n1140_n3288# 0.016978f
C289 drain_right.n114 a_n1140_n3288# 0.016493f
C290 drain_right.n115 a_n1140_n3288# 0.030692f
C291 drain_right.n116 a_n1140_n3288# 0.030692f
C292 drain_right.n117 a_n1140_n3288# 0.016493f
C293 drain_right.n118 a_n1140_n3288# 0.017463f
C294 drain_right.n119 a_n1140_n3288# 0.038982f
C295 drain_right.n120 a_n1140_n3288# 0.038982f
C296 drain_right.n121 a_n1140_n3288# 0.017463f
C297 drain_right.n122 a_n1140_n3288# 0.016493f
C298 drain_right.n123 a_n1140_n3288# 0.030692f
C299 drain_right.n124 a_n1140_n3288# 0.030692f
C300 drain_right.n125 a_n1140_n3288# 0.016493f
C301 drain_right.n126 a_n1140_n3288# 0.017463f
C302 drain_right.n127 a_n1140_n3288# 0.038982f
C303 drain_right.n128 a_n1140_n3288# 0.079996f
C304 drain_right.n129 a_n1140_n3288# 0.017463f
C305 drain_right.n130 a_n1140_n3288# 0.016493f
C306 drain_right.n131 a_n1140_n3288# 0.065911f
C307 drain_right.n132 a_n1140_n3288# 0.065385f
C308 drain_right.n133 a_n1140_n3288# 0.708435f
C309 source.n0 a_n1140_n3288# 0.037798f
C310 source.n1 a_n1140_n3288# 0.028535f
C311 source.n2 a_n1140_n3288# 0.015333f
C312 source.n3 a_n1140_n3288# 0.036243f
C313 source.n4 a_n1140_n3288# 0.016235f
C314 source.n5 a_n1140_n3288# 0.028535f
C315 source.n6 a_n1140_n3288# 0.015333f
C316 source.n7 a_n1140_n3288# 0.036243f
C317 source.n8 a_n1140_n3288# 0.016235f
C318 source.n9 a_n1140_n3288# 0.028535f
C319 source.n10 a_n1140_n3288# 0.015784f
C320 source.n11 a_n1140_n3288# 0.036243f
C321 source.n12 a_n1140_n3288# 0.015333f
C322 source.n13 a_n1140_n3288# 0.016235f
C323 source.n14 a_n1140_n3288# 0.028535f
C324 source.n15 a_n1140_n3288# 0.015333f
C325 source.n16 a_n1140_n3288# 0.036243f
C326 source.n17 a_n1140_n3288# 0.016235f
C327 source.n18 a_n1140_n3288# 0.028535f
C328 source.n19 a_n1140_n3288# 0.015333f
C329 source.n20 a_n1140_n3288# 0.027182f
C330 source.n21 a_n1140_n3288# 0.025621f
C331 source.t1 a_n1140_n3288# 0.061211f
C332 source.n22 a_n1140_n3288# 0.205734f
C333 source.n23 a_n1140_n3288# 1.43954f
C334 source.n24 a_n1140_n3288# 0.015333f
C335 source.n25 a_n1140_n3288# 0.016235f
C336 source.n26 a_n1140_n3288# 0.036243f
C337 source.n27 a_n1140_n3288# 0.036243f
C338 source.n28 a_n1140_n3288# 0.016235f
C339 source.n29 a_n1140_n3288# 0.015333f
C340 source.n30 a_n1140_n3288# 0.028535f
C341 source.n31 a_n1140_n3288# 0.028535f
C342 source.n32 a_n1140_n3288# 0.015333f
C343 source.n33 a_n1140_n3288# 0.016235f
C344 source.n34 a_n1140_n3288# 0.036243f
C345 source.n35 a_n1140_n3288# 0.036243f
C346 source.n36 a_n1140_n3288# 0.016235f
C347 source.n37 a_n1140_n3288# 0.015333f
C348 source.n38 a_n1140_n3288# 0.028535f
C349 source.n39 a_n1140_n3288# 0.028535f
C350 source.n40 a_n1140_n3288# 0.015333f
C351 source.n41 a_n1140_n3288# 0.016235f
C352 source.n42 a_n1140_n3288# 0.036243f
C353 source.n43 a_n1140_n3288# 0.036243f
C354 source.n44 a_n1140_n3288# 0.036243f
C355 source.n45 a_n1140_n3288# 0.015784f
C356 source.n46 a_n1140_n3288# 0.015333f
C357 source.n47 a_n1140_n3288# 0.028535f
C358 source.n48 a_n1140_n3288# 0.028535f
C359 source.n49 a_n1140_n3288# 0.015333f
C360 source.n50 a_n1140_n3288# 0.016235f
C361 source.n51 a_n1140_n3288# 0.036243f
C362 source.n52 a_n1140_n3288# 0.036243f
C363 source.n53 a_n1140_n3288# 0.016235f
C364 source.n54 a_n1140_n3288# 0.015333f
C365 source.n55 a_n1140_n3288# 0.028535f
C366 source.n56 a_n1140_n3288# 0.028535f
C367 source.n57 a_n1140_n3288# 0.015333f
C368 source.n58 a_n1140_n3288# 0.016235f
C369 source.n59 a_n1140_n3288# 0.036243f
C370 source.n60 a_n1140_n3288# 0.074374f
C371 source.n61 a_n1140_n3288# 0.016235f
C372 source.n62 a_n1140_n3288# 0.015333f
C373 source.n63 a_n1140_n3288# 0.061279f
C374 source.n64 a_n1140_n3288# 0.041046f
C375 source.n65 a_n1140_n3288# 1.13538f
C376 source.t2 a_n1140_n3288# 0.27059f
C377 source.t0 a_n1140_n3288# 0.27059f
C378 source.n66 a_n1140_n3288# 2.3168f
C379 source.n67 a_n1140_n3288# 0.397947f
C380 source.n68 a_n1140_n3288# 0.037798f
C381 source.n69 a_n1140_n3288# 0.028535f
C382 source.n70 a_n1140_n3288# 0.015333f
C383 source.n71 a_n1140_n3288# 0.036243f
C384 source.n72 a_n1140_n3288# 0.016235f
C385 source.n73 a_n1140_n3288# 0.028535f
C386 source.n74 a_n1140_n3288# 0.015333f
C387 source.n75 a_n1140_n3288# 0.036243f
C388 source.n76 a_n1140_n3288# 0.016235f
C389 source.n77 a_n1140_n3288# 0.028535f
C390 source.n78 a_n1140_n3288# 0.015784f
C391 source.n79 a_n1140_n3288# 0.036243f
C392 source.n80 a_n1140_n3288# 0.015333f
C393 source.n81 a_n1140_n3288# 0.016235f
C394 source.n82 a_n1140_n3288# 0.028535f
C395 source.n83 a_n1140_n3288# 0.015333f
C396 source.n84 a_n1140_n3288# 0.036243f
C397 source.n85 a_n1140_n3288# 0.016235f
C398 source.n86 a_n1140_n3288# 0.028535f
C399 source.n87 a_n1140_n3288# 0.015333f
C400 source.n88 a_n1140_n3288# 0.027182f
C401 source.n89 a_n1140_n3288# 0.025621f
C402 source.t9 a_n1140_n3288# 0.061211f
C403 source.n90 a_n1140_n3288# 0.205734f
C404 source.n91 a_n1140_n3288# 1.43954f
C405 source.n92 a_n1140_n3288# 0.015333f
C406 source.n93 a_n1140_n3288# 0.016235f
C407 source.n94 a_n1140_n3288# 0.036243f
C408 source.n95 a_n1140_n3288# 0.036243f
C409 source.n96 a_n1140_n3288# 0.016235f
C410 source.n97 a_n1140_n3288# 0.015333f
C411 source.n98 a_n1140_n3288# 0.028535f
C412 source.n99 a_n1140_n3288# 0.028535f
C413 source.n100 a_n1140_n3288# 0.015333f
C414 source.n101 a_n1140_n3288# 0.016235f
C415 source.n102 a_n1140_n3288# 0.036243f
C416 source.n103 a_n1140_n3288# 0.036243f
C417 source.n104 a_n1140_n3288# 0.016235f
C418 source.n105 a_n1140_n3288# 0.015333f
C419 source.n106 a_n1140_n3288# 0.028535f
C420 source.n107 a_n1140_n3288# 0.028535f
C421 source.n108 a_n1140_n3288# 0.015333f
C422 source.n109 a_n1140_n3288# 0.016235f
C423 source.n110 a_n1140_n3288# 0.036243f
C424 source.n111 a_n1140_n3288# 0.036243f
C425 source.n112 a_n1140_n3288# 0.036243f
C426 source.n113 a_n1140_n3288# 0.015784f
C427 source.n114 a_n1140_n3288# 0.015333f
C428 source.n115 a_n1140_n3288# 0.028535f
C429 source.n116 a_n1140_n3288# 0.028535f
C430 source.n117 a_n1140_n3288# 0.015333f
C431 source.n118 a_n1140_n3288# 0.016235f
C432 source.n119 a_n1140_n3288# 0.036243f
C433 source.n120 a_n1140_n3288# 0.036243f
C434 source.n121 a_n1140_n3288# 0.016235f
C435 source.n122 a_n1140_n3288# 0.015333f
C436 source.n123 a_n1140_n3288# 0.028535f
C437 source.n124 a_n1140_n3288# 0.028535f
C438 source.n125 a_n1140_n3288# 0.015333f
C439 source.n126 a_n1140_n3288# 0.016235f
C440 source.n127 a_n1140_n3288# 0.036243f
C441 source.n128 a_n1140_n3288# 0.074374f
C442 source.n129 a_n1140_n3288# 0.016235f
C443 source.n130 a_n1140_n3288# 0.015333f
C444 source.n131 a_n1140_n3288# 0.061279f
C445 source.n132 a_n1140_n3288# 0.041046f
C446 source.n133 a_n1140_n3288# 0.127949f
C447 source.t8 a_n1140_n3288# 0.27059f
C448 source.t11 a_n1140_n3288# 0.27059f
C449 source.n134 a_n1140_n3288# 2.3168f
C450 source.n135 a_n1140_n3288# 1.89323f
C451 source.t5 a_n1140_n3288# 0.27059f
C452 source.t3 a_n1140_n3288# 0.27059f
C453 source.n136 a_n1140_n3288# 2.31678f
C454 source.n137 a_n1140_n3288# 1.89324f
C455 source.n138 a_n1140_n3288# 0.037798f
C456 source.n139 a_n1140_n3288# 0.028535f
C457 source.n140 a_n1140_n3288# 0.015333f
C458 source.n141 a_n1140_n3288# 0.036243f
C459 source.n142 a_n1140_n3288# 0.016235f
C460 source.n143 a_n1140_n3288# 0.028535f
C461 source.n144 a_n1140_n3288# 0.015333f
C462 source.n145 a_n1140_n3288# 0.036243f
C463 source.n146 a_n1140_n3288# 0.016235f
C464 source.n147 a_n1140_n3288# 0.028535f
C465 source.n148 a_n1140_n3288# 0.015784f
C466 source.n149 a_n1140_n3288# 0.036243f
C467 source.n150 a_n1140_n3288# 0.016235f
C468 source.n151 a_n1140_n3288# 0.028535f
C469 source.n152 a_n1140_n3288# 0.015333f
C470 source.n153 a_n1140_n3288# 0.036243f
C471 source.n154 a_n1140_n3288# 0.016235f
C472 source.n155 a_n1140_n3288# 0.028535f
C473 source.n156 a_n1140_n3288# 0.015333f
C474 source.n157 a_n1140_n3288# 0.027182f
C475 source.n158 a_n1140_n3288# 0.025621f
C476 source.t4 a_n1140_n3288# 0.061211f
C477 source.n159 a_n1140_n3288# 0.205734f
C478 source.n160 a_n1140_n3288# 1.43954f
C479 source.n161 a_n1140_n3288# 0.015333f
C480 source.n162 a_n1140_n3288# 0.016235f
C481 source.n163 a_n1140_n3288# 0.036243f
C482 source.n164 a_n1140_n3288# 0.036243f
C483 source.n165 a_n1140_n3288# 0.016235f
C484 source.n166 a_n1140_n3288# 0.015333f
C485 source.n167 a_n1140_n3288# 0.028535f
C486 source.n168 a_n1140_n3288# 0.028535f
C487 source.n169 a_n1140_n3288# 0.015333f
C488 source.n170 a_n1140_n3288# 0.016235f
C489 source.n171 a_n1140_n3288# 0.036243f
C490 source.n172 a_n1140_n3288# 0.036243f
C491 source.n173 a_n1140_n3288# 0.016235f
C492 source.n174 a_n1140_n3288# 0.015333f
C493 source.n175 a_n1140_n3288# 0.028535f
C494 source.n176 a_n1140_n3288# 0.028535f
C495 source.n177 a_n1140_n3288# 0.015333f
C496 source.n178 a_n1140_n3288# 0.015333f
C497 source.n179 a_n1140_n3288# 0.016235f
C498 source.n180 a_n1140_n3288# 0.036243f
C499 source.n181 a_n1140_n3288# 0.036243f
C500 source.n182 a_n1140_n3288# 0.036243f
C501 source.n183 a_n1140_n3288# 0.015784f
C502 source.n184 a_n1140_n3288# 0.015333f
C503 source.n185 a_n1140_n3288# 0.028535f
C504 source.n186 a_n1140_n3288# 0.028535f
C505 source.n187 a_n1140_n3288# 0.015333f
C506 source.n188 a_n1140_n3288# 0.016235f
C507 source.n189 a_n1140_n3288# 0.036243f
C508 source.n190 a_n1140_n3288# 0.036243f
C509 source.n191 a_n1140_n3288# 0.016235f
C510 source.n192 a_n1140_n3288# 0.015333f
C511 source.n193 a_n1140_n3288# 0.028535f
C512 source.n194 a_n1140_n3288# 0.028535f
C513 source.n195 a_n1140_n3288# 0.015333f
C514 source.n196 a_n1140_n3288# 0.016235f
C515 source.n197 a_n1140_n3288# 0.036243f
C516 source.n198 a_n1140_n3288# 0.074374f
C517 source.n199 a_n1140_n3288# 0.016235f
C518 source.n200 a_n1140_n3288# 0.015333f
C519 source.n201 a_n1140_n3288# 0.061279f
C520 source.n202 a_n1140_n3288# 0.041046f
C521 source.n203 a_n1140_n3288# 0.127949f
C522 source.t6 a_n1140_n3288# 0.27059f
C523 source.t7 a_n1140_n3288# 0.27059f
C524 source.n204 a_n1140_n3288# 2.31678f
C525 source.n205 a_n1140_n3288# 0.397961f
C526 source.n206 a_n1140_n3288# 0.037798f
C527 source.n207 a_n1140_n3288# 0.028535f
C528 source.n208 a_n1140_n3288# 0.015333f
C529 source.n209 a_n1140_n3288# 0.036243f
C530 source.n210 a_n1140_n3288# 0.016235f
C531 source.n211 a_n1140_n3288# 0.028535f
C532 source.n212 a_n1140_n3288# 0.015333f
C533 source.n213 a_n1140_n3288# 0.036243f
C534 source.n214 a_n1140_n3288# 0.016235f
C535 source.n215 a_n1140_n3288# 0.028535f
C536 source.n216 a_n1140_n3288# 0.015784f
C537 source.n217 a_n1140_n3288# 0.036243f
C538 source.n218 a_n1140_n3288# 0.016235f
C539 source.n219 a_n1140_n3288# 0.028535f
C540 source.n220 a_n1140_n3288# 0.015333f
C541 source.n221 a_n1140_n3288# 0.036243f
C542 source.n222 a_n1140_n3288# 0.016235f
C543 source.n223 a_n1140_n3288# 0.028535f
C544 source.n224 a_n1140_n3288# 0.015333f
C545 source.n225 a_n1140_n3288# 0.027182f
C546 source.n226 a_n1140_n3288# 0.025621f
C547 source.t10 a_n1140_n3288# 0.061211f
C548 source.n227 a_n1140_n3288# 0.205734f
C549 source.n228 a_n1140_n3288# 1.43954f
C550 source.n229 a_n1140_n3288# 0.015333f
C551 source.n230 a_n1140_n3288# 0.016235f
C552 source.n231 a_n1140_n3288# 0.036243f
C553 source.n232 a_n1140_n3288# 0.036243f
C554 source.n233 a_n1140_n3288# 0.016235f
C555 source.n234 a_n1140_n3288# 0.015333f
C556 source.n235 a_n1140_n3288# 0.028535f
C557 source.n236 a_n1140_n3288# 0.028535f
C558 source.n237 a_n1140_n3288# 0.015333f
C559 source.n238 a_n1140_n3288# 0.016235f
C560 source.n239 a_n1140_n3288# 0.036243f
C561 source.n240 a_n1140_n3288# 0.036243f
C562 source.n241 a_n1140_n3288# 0.016235f
C563 source.n242 a_n1140_n3288# 0.015333f
C564 source.n243 a_n1140_n3288# 0.028535f
C565 source.n244 a_n1140_n3288# 0.028535f
C566 source.n245 a_n1140_n3288# 0.015333f
C567 source.n246 a_n1140_n3288# 0.015333f
C568 source.n247 a_n1140_n3288# 0.016235f
C569 source.n248 a_n1140_n3288# 0.036243f
C570 source.n249 a_n1140_n3288# 0.036243f
C571 source.n250 a_n1140_n3288# 0.036243f
C572 source.n251 a_n1140_n3288# 0.015784f
C573 source.n252 a_n1140_n3288# 0.015333f
C574 source.n253 a_n1140_n3288# 0.028535f
C575 source.n254 a_n1140_n3288# 0.028535f
C576 source.n255 a_n1140_n3288# 0.015333f
C577 source.n256 a_n1140_n3288# 0.016235f
C578 source.n257 a_n1140_n3288# 0.036243f
C579 source.n258 a_n1140_n3288# 0.036243f
C580 source.n259 a_n1140_n3288# 0.016235f
C581 source.n260 a_n1140_n3288# 0.015333f
C582 source.n261 a_n1140_n3288# 0.028535f
C583 source.n262 a_n1140_n3288# 0.028535f
C584 source.n263 a_n1140_n3288# 0.015333f
C585 source.n264 a_n1140_n3288# 0.016235f
C586 source.n265 a_n1140_n3288# 0.036243f
C587 source.n266 a_n1140_n3288# 0.074374f
C588 source.n267 a_n1140_n3288# 0.016235f
C589 source.n268 a_n1140_n3288# 0.015333f
C590 source.n269 a_n1140_n3288# 0.061279f
C591 source.n270 a_n1140_n3288# 0.041046f
C592 source.n271 a_n1140_n3288# 0.26167f
C593 source.n272 a_n1140_n3288# 1.78569f
C594 minus.t5 a_n1140_n3288# 0.339519f
C595 minus.n0 a_n1140_n3288# 0.151801f
C596 minus.t0 a_n1140_n3288# 0.339519f
C597 minus.t4 a_n1140_n3288# 0.33609f
C598 minus.n1 a_n1140_n3288# 0.138417f
C599 minus.n2 a_n1140_n3288# 0.151733f
C600 minus.n3 a_n1140_n3288# 1.59435f
C601 minus.t2 a_n1140_n3288# 0.339519f
C602 minus.n4 a_n1140_n3288# 0.151801f
C603 minus.t3 a_n1140_n3288# 0.33609f
C604 minus.n5 a_n1140_n3288# 0.138417f
C605 minus.t1 a_n1140_n3288# 0.339519f
C606 minus.n6 a_n1140_n3288# 0.151733f
C607 minus.n7 a_n1140_n3288# 0.37416f
C608 minus.n8 a_n1140_n3288# 1.88479f
.ends

