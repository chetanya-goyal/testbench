* NGSPICE file created from diffpair501.ext - technology: sky130A

.subckt diffpair501 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t6 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X1 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X2 source.t2 plus.t0 drain_left.t3 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X3 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X4 drain_left.t2 plus.t1 source.t0 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X5 drain_left.t1 plus.t2 source.t1 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X6 source.t4 minus.t1 drain_right.t2 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X7 source.t7 minus.t2 drain_right.t1 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X9 source.t3 plus.t3 drain_left.t0 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X10 drain_right.t0 minus.t3 source.t5 a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X11 a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# a_n1064_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
R0 minus.n0 minus.t1 1613.68
R1 minus.n0 minus.t0 1613.68
R2 minus.n1 minus.t3 1613.68
R3 minus.n1 minus.t2 1613.68
R4 minus.n2 minus.n0 196.709
R5 minus.n2 minus.n1 167.77
R6 minus minus.n2 0.188
R7 source.n1 source.t3 45.521
R8 source.n2 source.t6 45.521
R9 source.n3 source.t4 45.521
R10 source.n7 source.t5 45.5208
R11 source.n6 source.t7 45.5208
R12 source.n5 source.t1 45.5208
R13 source.n4 source.t2 45.5208
R14 source.n0 source.t0 45.5208
R15 source.n4 source.n3 24.0756
R16 source.n8 source.n0 18.5627
R17 source.n8 source.n7 5.51343
R18 source.n3 source.n2 0.5005
R19 source.n1 source.n0 0.5005
R20 source.n5 source.n4 0.5005
R21 source.n7 source.n6 0.5005
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 90.9808
R26 drain_right drain_right.n1 67.0323
R27 drain_right.n0 drain_right.t1 1.3205
R28 drain_right.n0 drain_right.t0 1.3205
R29 drain_right.n1 drain_right.t2 1.3205
R30 drain_right.n1 drain_right.t3 1.3205
R31 plus.n0 plus.t3 1613.68
R32 plus.n0 plus.t1 1613.68
R33 plus.n1 plus.t2 1613.68
R34 plus.n1 plus.t0 1613.68
R35 plus plus.n1 189.454
R36 plus plus.n0 174.55
R37 drain_left drain_left.n0 91.534
R38 drain_left drain_left.n1 67.0323
R39 drain_left.n0 drain_left.t3 1.3205
R40 drain_left.n0 drain_left.t1 1.3205
R41 drain_left.n1 drain_left.t0 1.3205
R42 drain_left.n1 drain_left.t2 1.3205
C0 drain_left drain_right 0.467153f
C1 drain_left source 12.5092f
C2 drain_left minus 0.171285f
C3 source drain_right 12.507401f
C4 minus drain_right 2.32761f
C5 source minus 1.63459f
C6 plus drain_left 2.42544f
C7 plus drain_right 0.251889f
C8 plus source 1.64863f
C9 plus minus 5.02981f
C10 drain_right a_n1064_n3892# 7.85614f
C11 drain_left a_n1064_n3892# 8.05177f
C12 source a_n1064_n3892# 9.643491f
C13 minus a_n1064_n3892# 4.254276f
C14 plus a_n1064_n3892# 8.0915f
C15 drain_left.t3 a_n1064_n3892# 0.404358f
C16 drain_left.t1 a_n1064_n3892# 0.404358f
C17 drain_left.n0 a_n1064_n3892# 4.25704f
C18 drain_left.t0 a_n1064_n3892# 0.404358f
C19 drain_left.t2 a_n1064_n3892# 0.404358f
C20 drain_left.n1 a_n1064_n3892# 3.71775f
C21 plus.t3 a_n1064_n3892# 0.561577f
C22 plus.t1 a_n1064_n3892# 0.561577f
C23 plus.n0 a_n1064_n3892# 0.494551f
C24 plus.t0 a_n1064_n3892# 0.561577f
C25 plus.t2 a_n1064_n3892# 0.561577f
C26 plus.n1 a_n1064_n3892# 0.662748f
C27 drain_right.t1 a_n1064_n3892# 0.405274f
C28 drain_right.t0 a_n1064_n3892# 0.405274f
C29 drain_right.n0 a_n1064_n3892# 4.23551f
C30 drain_right.t2 a_n1064_n3892# 0.405274f
C31 drain_right.t3 a_n1064_n3892# 0.405274f
C32 drain_right.n1 a_n1064_n3892# 3.72617f
C33 source.t0 a_n1064_n3892# 2.30109f
C34 source.n0 a_n1064_n3892# 1.06294f
C35 source.t3 a_n1064_n3892# 2.30109f
C36 source.n1 a_n1064_n3892# 0.28735f
C37 source.t6 a_n1064_n3892# 2.30109f
C38 source.n2 a_n1064_n3892# 0.28735f
C39 source.t4 a_n1064_n3892# 2.30109f
C40 source.n3 a_n1064_n3892# 1.3501f
C41 source.t2 a_n1064_n3892# 2.30109f
C42 source.n4 a_n1064_n3892# 1.35011f
C43 source.t1 a_n1064_n3892# 2.30109f
C44 source.n5 a_n1064_n3892# 0.287353f
C45 source.t7 a_n1064_n3892# 2.30109f
C46 source.n6 a_n1064_n3892# 0.287353f
C47 source.t5 a_n1064_n3892# 2.30109f
C48 source.n7 a_n1064_n3892# 0.383213f
C49 source.n8 a_n1064_n3892# 1.26638f
C50 minus.t1 a_n1064_n3892# 0.546146f
C51 minus.t0 a_n1064_n3892# 0.546146f
C52 minus.n0 a_n1064_n3892# 0.747107f
C53 minus.t2 a_n1064_n3892# 0.546146f
C54 minus.t3 a_n1064_n3892# 0.546146f
C55 minus.n1 a_n1064_n3892# 0.444573f
C56 minus.n2 a_n1064_n3892# 3.89018f
.ends

