* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X1 drain_right.t0 minus.t1 source.t1 a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X2 drain_left.t1 plus.t0 source.t3 a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X3 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X4 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5 drain_left.t0 plus.t1 source.t0 a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X6 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
R0 minus.n0 minus.t0 579.333
R1 minus.n0 minus.t1 561.333
R2 minus minus.n0 0.188
R3 source.n0 source.t3 253.454
R4 source.n1 source.t2 253.454
R5 source.n3 source.t1 253.453
R6 source.n2 source.t0 253.453
R7 source.n2 source.n1 14.0902
R8 source.n4 source.n0 7.98679
R9 source.n4 source.n3 5.5436
R10 source.n1 source.n0 0.7505
R11 source.n3 source.n2 0.7505
R12 source source.n4 0.188
R13 drain_right drain_right.t0 289.413
R14 drain_right drain_right.t1 276.065
R15 plus plus.t1 577.381
R16 plus plus.t0 562.811
R17 drain_left drain_left.t0 289.966
R18 drain_left drain_left.t1 276.346
C0 drain_left minus 0.178817f
C1 source plus 0.36424f
C2 drain_right source 1.665f
C3 drain_left plus 0.395415f
C4 drain_right drain_left 0.423967f
C5 minus plus 2.34042f
C6 drain_right minus 0.306873f
C7 drain_right plus 0.251385f
C8 source drain_left 1.66516f
C9 source minus 0.350323f
C10 drain_right a_n976_n1092# 1.57271f
C11 drain_left a_n976_n1092# 1.66964f
C12 source a_n976_n1092# 1.67047f
C13 minus a_n976_n1092# 2.755354f
C14 plus a_n976_n1092# 4.77335f
C15 plus.t0 a_n976_n1092# 0.039087f
C16 plus.t1 a_n976_n1092# 0.068471f
C17 minus.t0 a_n976_n1092# 0.068862f
C18 minus.t1 a_n976_n1092# 0.036454f
C19 minus.n0 a_n976_n1092# 2.16384f
.ends

