* NGSPICE file created from diffpair437.ext - technology: sky130A

.subckt diffpair437 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t13 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X1 source.t30 minus.t1 drain_right.t11 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X2 drain_left.t15 plus.t0 source.t1 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X3 source.t29 minus.t2 drain_right.t3 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X4 drain_right.t10 minus.t3 source.t28 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X5 a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.3
X6 drain_left.t14 plus.t1 source.t3 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X7 source.t6 plus.t2 drain_left.t13 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X8 drain_left.t12 plus.t3 source.t9 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X9 a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X10 drain_right.t8 minus.t4 source.t27 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X11 source.t26 minus.t5 drain_right.t14 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X12 source.t25 minus.t6 drain_right.t15 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X13 source.t0 plus.t4 drain_left.t11 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X14 source.t10 plus.t5 drain_left.t10 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X15 drain_left.t9 plus.t6 source.t5 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X16 source.t24 minus.t7 drain_right.t9 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X17 source.t11 plus.t7 drain_left.t8 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X18 source.t14 plus.t8 drain_left.t7 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X19 drain_right.t12 minus.t8 source.t23 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X20 a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X21 drain_left.t6 plus.t9 source.t2 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X22 a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X23 drain_right.t4 minus.t9 source.t22 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X24 drain_right.t7 minus.t10 source.t21 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X25 source.t13 plus.t10 drain_left.t5 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X26 drain_right.t0 minus.t11 source.t20 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X27 source.t4 plus.t11 drain_left.t4 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X28 drain_right.t1 minus.t12 source.t19 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X29 drain_right.t5 minus.t13 source.t18 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X30 drain_left.t3 plus.t12 source.t7 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X31 drain_left.t2 plus.t13 source.t15 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X32 source.t17 minus.t14 drain_right.t2 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X33 source.t16 minus.t15 drain_right.t6 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X34 source.t8 plus.t14 drain_left.t1 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X35 drain_left.t0 plus.t15 source.t12 a_n1850_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
R0 minus.n21 minus.t15 1098.38
R1 minus.n5 minus.t8 1098.38
R2 minus.n44 minus.t11 1098.38
R3 minus.n28 minus.t1 1098.38
R4 minus.n20 minus.t4 1068.43
R5 minus.n1 minus.t2 1068.43
R6 minus.n14 minus.t13 1068.43
R7 minus.n12 minus.t7 1068.43
R8 minus.n3 minus.t3 1068.43
R9 minus.n6 minus.t14 1068.43
R10 minus.n43 minus.t5 1068.43
R11 minus.n24 minus.t12 1068.43
R12 minus.n37 minus.t6 1068.43
R13 minus.n35 minus.t9 1068.43
R14 minus.n26 minus.t0 1068.43
R15 minus.n29 minus.t10 1068.43
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 64.9975
R39 minus.n11 minus.n3 64.9975
R40 minus.n34 minus.n26 64.9975
R41 minus.n38 minus.n24 64.9975
R42 minus.n21 minus.n20 62.0763
R43 minus.n6 minus.n5 62.0763
R44 minus.n29 minus.n28 62.0763
R45 minus.n44 minus.n43 62.0763
R46 minus.n14 minus.n13 46.0096
R47 minus.n13 minus.n12 46.0096
R48 minus.n36 minus.n35 46.0096
R49 minus.n37 minus.n36 46.0096
R50 minus.n46 minus.n22 36.0952
R51 minus.n15 minus.n14 27.0217
R52 minus.n12 minus.n11 27.0217
R53 minus.n35 minus.n34 27.0217
R54 minus.n38 minus.n37 27.0217
R55 minus.n20 minus.n19 10.955
R56 minus.n7 minus.n6 10.955
R57 minus.n30 minus.n29 10.955
R58 minus.n43 minus.n42 10.955
R59 minus.n18 minus.n1 8.03383
R60 minus.n8 minus.n3 8.03383
R61 minus.n31 minus.n26 8.03383
R62 minus.n41 minus.n24 8.03383
R63 minus.n46 minus.n45 6.46641
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 drain_right.n5 drain_right.n3 60.0956
R80 drain_right.n2 drain_right.n0 60.0956
R81 drain_right.n9 drain_right.n7 60.0956
R82 drain_right.n9 drain_right.n8 59.5527
R83 drain_right.n11 drain_right.n10 59.5527
R84 drain_right.n13 drain_right.n12 59.5527
R85 drain_right.n5 drain_right.n4 59.5525
R86 drain_right.n2 drain_right.n1 59.5525
R87 drain_right drain_right.n6 30.344
R88 drain_right drain_right.n13 6.19632
R89 drain_right.n3 drain_right.t14 1.6505
R90 drain_right.n3 drain_right.t0 1.6505
R91 drain_right.n4 drain_right.t15 1.6505
R92 drain_right.n4 drain_right.t1 1.6505
R93 drain_right.n1 drain_right.t13 1.6505
R94 drain_right.n1 drain_right.t4 1.6505
R95 drain_right.n0 drain_right.t11 1.6505
R96 drain_right.n0 drain_right.t7 1.6505
R97 drain_right.n7 drain_right.t2 1.6505
R98 drain_right.n7 drain_right.t12 1.6505
R99 drain_right.n8 drain_right.t9 1.6505
R100 drain_right.n8 drain_right.t10 1.6505
R101 drain_right.n10 drain_right.t3 1.6505
R102 drain_right.n10 drain_right.t5 1.6505
R103 drain_right.n12 drain_right.t6 1.6505
R104 drain_right.n12 drain_right.t8 1.6505
R105 drain_right.n13 drain_right.n11 0.543603
R106 drain_right.n11 drain_right.n9 0.543603
R107 drain_right.n6 drain_right.n5 0.216706
R108 drain_right.n6 drain_right.n2 0.216706
R109 source.n546 source.n486 289.615
R110 source.n474 source.n414 289.615
R111 source.n408 source.n348 289.615
R112 source.n336 source.n276 289.615
R113 source.n60 source.n0 289.615
R114 source.n132 source.n72 289.615
R115 source.n198 source.n138 289.615
R116 source.n270 source.n210 289.615
R117 source.n506 source.n505 185
R118 source.n511 source.n510 185
R119 source.n513 source.n512 185
R120 source.n502 source.n501 185
R121 source.n519 source.n518 185
R122 source.n521 source.n520 185
R123 source.n498 source.n497 185
R124 source.n528 source.n527 185
R125 source.n529 source.n496 185
R126 source.n531 source.n530 185
R127 source.n494 source.n493 185
R128 source.n537 source.n536 185
R129 source.n539 source.n538 185
R130 source.n490 source.n489 185
R131 source.n545 source.n544 185
R132 source.n547 source.n546 185
R133 source.n434 source.n433 185
R134 source.n439 source.n438 185
R135 source.n441 source.n440 185
R136 source.n430 source.n429 185
R137 source.n447 source.n446 185
R138 source.n449 source.n448 185
R139 source.n426 source.n425 185
R140 source.n456 source.n455 185
R141 source.n457 source.n424 185
R142 source.n459 source.n458 185
R143 source.n422 source.n421 185
R144 source.n465 source.n464 185
R145 source.n467 source.n466 185
R146 source.n418 source.n417 185
R147 source.n473 source.n472 185
R148 source.n475 source.n474 185
R149 source.n368 source.n367 185
R150 source.n373 source.n372 185
R151 source.n375 source.n374 185
R152 source.n364 source.n363 185
R153 source.n381 source.n380 185
R154 source.n383 source.n382 185
R155 source.n360 source.n359 185
R156 source.n390 source.n389 185
R157 source.n391 source.n358 185
R158 source.n393 source.n392 185
R159 source.n356 source.n355 185
R160 source.n399 source.n398 185
R161 source.n401 source.n400 185
R162 source.n352 source.n351 185
R163 source.n407 source.n406 185
R164 source.n409 source.n408 185
R165 source.n296 source.n295 185
R166 source.n301 source.n300 185
R167 source.n303 source.n302 185
R168 source.n292 source.n291 185
R169 source.n309 source.n308 185
R170 source.n311 source.n310 185
R171 source.n288 source.n287 185
R172 source.n318 source.n317 185
R173 source.n319 source.n286 185
R174 source.n321 source.n320 185
R175 source.n284 source.n283 185
R176 source.n327 source.n326 185
R177 source.n329 source.n328 185
R178 source.n280 source.n279 185
R179 source.n335 source.n334 185
R180 source.n337 source.n336 185
R181 source.n61 source.n60 185
R182 source.n59 source.n58 185
R183 source.n4 source.n3 185
R184 source.n53 source.n52 185
R185 source.n51 source.n50 185
R186 source.n8 source.n7 185
R187 source.n45 source.n44 185
R188 source.n43 source.n10 185
R189 source.n42 source.n41 185
R190 source.n13 source.n11 185
R191 source.n36 source.n35 185
R192 source.n34 source.n33 185
R193 source.n17 source.n16 185
R194 source.n28 source.n27 185
R195 source.n26 source.n25 185
R196 source.n21 source.n20 185
R197 source.n133 source.n132 185
R198 source.n131 source.n130 185
R199 source.n76 source.n75 185
R200 source.n125 source.n124 185
R201 source.n123 source.n122 185
R202 source.n80 source.n79 185
R203 source.n117 source.n116 185
R204 source.n115 source.n82 185
R205 source.n114 source.n113 185
R206 source.n85 source.n83 185
R207 source.n108 source.n107 185
R208 source.n106 source.n105 185
R209 source.n89 source.n88 185
R210 source.n100 source.n99 185
R211 source.n98 source.n97 185
R212 source.n93 source.n92 185
R213 source.n199 source.n198 185
R214 source.n197 source.n196 185
R215 source.n142 source.n141 185
R216 source.n191 source.n190 185
R217 source.n189 source.n188 185
R218 source.n146 source.n145 185
R219 source.n183 source.n182 185
R220 source.n181 source.n148 185
R221 source.n180 source.n179 185
R222 source.n151 source.n149 185
R223 source.n174 source.n173 185
R224 source.n172 source.n171 185
R225 source.n155 source.n154 185
R226 source.n166 source.n165 185
R227 source.n164 source.n163 185
R228 source.n159 source.n158 185
R229 source.n271 source.n270 185
R230 source.n269 source.n268 185
R231 source.n214 source.n213 185
R232 source.n263 source.n262 185
R233 source.n261 source.n260 185
R234 source.n218 source.n217 185
R235 source.n255 source.n254 185
R236 source.n253 source.n220 185
R237 source.n252 source.n251 185
R238 source.n223 source.n221 185
R239 source.n246 source.n245 185
R240 source.n244 source.n243 185
R241 source.n227 source.n226 185
R242 source.n238 source.n237 185
R243 source.n236 source.n235 185
R244 source.n231 source.n230 185
R245 source.n507 source.t20 149.524
R246 source.n435 source.t30 149.524
R247 source.n369 source.t7 149.524
R248 source.n297 source.t4 149.524
R249 source.n22 source.t1 149.524
R250 source.n94 source.t6 149.524
R251 source.n160 source.t23 149.524
R252 source.n232 source.t16 149.524
R253 source.n511 source.n505 104.615
R254 source.n512 source.n511 104.615
R255 source.n512 source.n501 104.615
R256 source.n519 source.n501 104.615
R257 source.n520 source.n519 104.615
R258 source.n520 source.n497 104.615
R259 source.n528 source.n497 104.615
R260 source.n529 source.n528 104.615
R261 source.n530 source.n529 104.615
R262 source.n530 source.n493 104.615
R263 source.n537 source.n493 104.615
R264 source.n538 source.n537 104.615
R265 source.n538 source.n489 104.615
R266 source.n545 source.n489 104.615
R267 source.n546 source.n545 104.615
R268 source.n439 source.n433 104.615
R269 source.n440 source.n439 104.615
R270 source.n440 source.n429 104.615
R271 source.n447 source.n429 104.615
R272 source.n448 source.n447 104.615
R273 source.n448 source.n425 104.615
R274 source.n456 source.n425 104.615
R275 source.n457 source.n456 104.615
R276 source.n458 source.n457 104.615
R277 source.n458 source.n421 104.615
R278 source.n465 source.n421 104.615
R279 source.n466 source.n465 104.615
R280 source.n466 source.n417 104.615
R281 source.n473 source.n417 104.615
R282 source.n474 source.n473 104.615
R283 source.n373 source.n367 104.615
R284 source.n374 source.n373 104.615
R285 source.n374 source.n363 104.615
R286 source.n381 source.n363 104.615
R287 source.n382 source.n381 104.615
R288 source.n382 source.n359 104.615
R289 source.n390 source.n359 104.615
R290 source.n391 source.n390 104.615
R291 source.n392 source.n391 104.615
R292 source.n392 source.n355 104.615
R293 source.n399 source.n355 104.615
R294 source.n400 source.n399 104.615
R295 source.n400 source.n351 104.615
R296 source.n407 source.n351 104.615
R297 source.n408 source.n407 104.615
R298 source.n301 source.n295 104.615
R299 source.n302 source.n301 104.615
R300 source.n302 source.n291 104.615
R301 source.n309 source.n291 104.615
R302 source.n310 source.n309 104.615
R303 source.n310 source.n287 104.615
R304 source.n318 source.n287 104.615
R305 source.n319 source.n318 104.615
R306 source.n320 source.n319 104.615
R307 source.n320 source.n283 104.615
R308 source.n327 source.n283 104.615
R309 source.n328 source.n327 104.615
R310 source.n328 source.n279 104.615
R311 source.n335 source.n279 104.615
R312 source.n336 source.n335 104.615
R313 source.n60 source.n59 104.615
R314 source.n59 source.n3 104.615
R315 source.n52 source.n3 104.615
R316 source.n52 source.n51 104.615
R317 source.n51 source.n7 104.615
R318 source.n44 source.n7 104.615
R319 source.n44 source.n43 104.615
R320 source.n43 source.n42 104.615
R321 source.n42 source.n11 104.615
R322 source.n35 source.n11 104.615
R323 source.n35 source.n34 104.615
R324 source.n34 source.n16 104.615
R325 source.n27 source.n16 104.615
R326 source.n27 source.n26 104.615
R327 source.n26 source.n20 104.615
R328 source.n132 source.n131 104.615
R329 source.n131 source.n75 104.615
R330 source.n124 source.n75 104.615
R331 source.n124 source.n123 104.615
R332 source.n123 source.n79 104.615
R333 source.n116 source.n79 104.615
R334 source.n116 source.n115 104.615
R335 source.n115 source.n114 104.615
R336 source.n114 source.n83 104.615
R337 source.n107 source.n83 104.615
R338 source.n107 source.n106 104.615
R339 source.n106 source.n88 104.615
R340 source.n99 source.n88 104.615
R341 source.n99 source.n98 104.615
R342 source.n98 source.n92 104.615
R343 source.n198 source.n197 104.615
R344 source.n197 source.n141 104.615
R345 source.n190 source.n141 104.615
R346 source.n190 source.n189 104.615
R347 source.n189 source.n145 104.615
R348 source.n182 source.n145 104.615
R349 source.n182 source.n181 104.615
R350 source.n181 source.n180 104.615
R351 source.n180 source.n149 104.615
R352 source.n173 source.n149 104.615
R353 source.n173 source.n172 104.615
R354 source.n172 source.n154 104.615
R355 source.n165 source.n154 104.615
R356 source.n165 source.n164 104.615
R357 source.n164 source.n158 104.615
R358 source.n270 source.n269 104.615
R359 source.n269 source.n213 104.615
R360 source.n262 source.n213 104.615
R361 source.n262 source.n261 104.615
R362 source.n261 source.n217 104.615
R363 source.n254 source.n217 104.615
R364 source.n254 source.n253 104.615
R365 source.n253 source.n252 104.615
R366 source.n252 source.n221 104.615
R367 source.n245 source.n221 104.615
R368 source.n245 source.n244 104.615
R369 source.n244 source.n226 104.615
R370 source.n237 source.n226 104.615
R371 source.n237 source.n236 104.615
R372 source.n236 source.n230 104.615
R373 source.t20 source.n505 52.3082
R374 source.t30 source.n433 52.3082
R375 source.t7 source.n367 52.3082
R376 source.t4 source.n295 52.3082
R377 source.t1 source.n20 52.3082
R378 source.t6 source.n92 52.3082
R379 source.t23 source.n158 52.3082
R380 source.t16 source.n230 52.3082
R381 source.n67 source.n66 42.8739
R382 source.n69 source.n68 42.8739
R383 source.n71 source.n70 42.8739
R384 source.n205 source.n204 42.8739
R385 source.n207 source.n206 42.8739
R386 source.n209 source.n208 42.8739
R387 source.n485 source.n484 42.8737
R388 source.n483 source.n482 42.8737
R389 source.n481 source.n480 42.8737
R390 source.n347 source.n346 42.8737
R391 source.n345 source.n344 42.8737
R392 source.n343 source.n342 42.8737
R393 source.n551 source.n550 29.8581
R394 source.n479 source.n478 29.8581
R395 source.n413 source.n412 29.8581
R396 source.n341 source.n340 29.8581
R397 source.n65 source.n64 29.8581
R398 source.n137 source.n136 29.8581
R399 source.n203 source.n202 29.8581
R400 source.n275 source.n274 29.8581
R401 source.n341 source.n275 21.8308
R402 source.n552 source.n65 16.2963
R403 source.n531 source.n496 13.1884
R404 source.n459 source.n424 13.1884
R405 source.n393 source.n358 13.1884
R406 source.n321 source.n286 13.1884
R407 source.n45 source.n10 13.1884
R408 source.n117 source.n82 13.1884
R409 source.n183 source.n148 13.1884
R410 source.n255 source.n220 13.1884
R411 source.n527 source.n526 12.8005
R412 source.n532 source.n494 12.8005
R413 source.n455 source.n454 12.8005
R414 source.n460 source.n422 12.8005
R415 source.n389 source.n388 12.8005
R416 source.n394 source.n356 12.8005
R417 source.n317 source.n316 12.8005
R418 source.n322 source.n284 12.8005
R419 source.n46 source.n8 12.8005
R420 source.n41 source.n12 12.8005
R421 source.n118 source.n80 12.8005
R422 source.n113 source.n84 12.8005
R423 source.n184 source.n146 12.8005
R424 source.n179 source.n150 12.8005
R425 source.n256 source.n218 12.8005
R426 source.n251 source.n222 12.8005
R427 source.n525 source.n498 12.0247
R428 source.n536 source.n535 12.0247
R429 source.n453 source.n426 12.0247
R430 source.n464 source.n463 12.0247
R431 source.n387 source.n360 12.0247
R432 source.n398 source.n397 12.0247
R433 source.n315 source.n288 12.0247
R434 source.n326 source.n325 12.0247
R435 source.n50 source.n49 12.0247
R436 source.n40 source.n13 12.0247
R437 source.n122 source.n121 12.0247
R438 source.n112 source.n85 12.0247
R439 source.n188 source.n187 12.0247
R440 source.n178 source.n151 12.0247
R441 source.n260 source.n259 12.0247
R442 source.n250 source.n223 12.0247
R443 source.n522 source.n521 11.249
R444 source.n539 source.n492 11.249
R445 source.n450 source.n449 11.249
R446 source.n467 source.n420 11.249
R447 source.n384 source.n383 11.249
R448 source.n401 source.n354 11.249
R449 source.n312 source.n311 11.249
R450 source.n329 source.n282 11.249
R451 source.n53 source.n6 11.249
R452 source.n37 source.n36 11.249
R453 source.n125 source.n78 11.249
R454 source.n109 source.n108 11.249
R455 source.n191 source.n144 11.249
R456 source.n175 source.n174 11.249
R457 source.n263 source.n216 11.249
R458 source.n247 source.n246 11.249
R459 source.n518 source.n500 10.4732
R460 source.n540 source.n490 10.4732
R461 source.n446 source.n428 10.4732
R462 source.n468 source.n418 10.4732
R463 source.n380 source.n362 10.4732
R464 source.n402 source.n352 10.4732
R465 source.n308 source.n290 10.4732
R466 source.n330 source.n280 10.4732
R467 source.n54 source.n4 10.4732
R468 source.n33 source.n15 10.4732
R469 source.n126 source.n76 10.4732
R470 source.n105 source.n87 10.4732
R471 source.n192 source.n142 10.4732
R472 source.n171 source.n153 10.4732
R473 source.n264 source.n214 10.4732
R474 source.n243 source.n225 10.4732
R475 source.n507 source.n506 10.2747
R476 source.n435 source.n434 10.2747
R477 source.n369 source.n368 10.2747
R478 source.n297 source.n296 10.2747
R479 source.n22 source.n21 10.2747
R480 source.n94 source.n93 10.2747
R481 source.n160 source.n159 10.2747
R482 source.n232 source.n231 10.2747
R483 source.n517 source.n502 9.69747
R484 source.n544 source.n543 9.69747
R485 source.n445 source.n430 9.69747
R486 source.n472 source.n471 9.69747
R487 source.n379 source.n364 9.69747
R488 source.n406 source.n405 9.69747
R489 source.n307 source.n292 9.69747
R490 source.n334 source.n333 9.69747
R491 source.n58 source.n57 9.69747
R492 source.n32 source.n17 9.69747
R493 source.n130 source.n129 9.69747
R494 source.n104 source.n89 9.69747
R495 source.n196 source.n195 9.69747
R496 source.n170 source.n155 9.69747
R497 source.n268 source.n267 9.69747
R498 source.n242 source.n227 9.69747
R499 source.n550 source.n549 9.45567
R500 source.n478 source.n477 9.45567
R501 source.n412 source.n411 9.45567
R502 source.n340 source.n339 9.45567
R503 source.n64 source.n63 9.45567
R504 source.n136 source.n135 9.45567
R505 source.n202 source.n201 9.45567
R506 source.n274 source.n273 9.45567
R507 source.n549 source.n548 9.3005
R508 source.n488 source.n487 9.3005
R509 source.n543 source.n542 9.3005
R510 source.n541 source.n540 9.3005
R511 source.n492 source.n491 9.3005
R512 source.n535 source.n534 9.3005
R513 source.n533 source.n532 9.3005
R514 source.n509 source.n508 9.3005
R515 source.n504 source.n503 9.3005
R516 source.n515 source.n514 9.3005
R517 source.n517 source.n516 9.3005
R518 source.n500 source.n499 9.3005
R519 source.n523 source.n522 9.3005
R520 source.n525 source.n524 9.3005
R521 source.n526 source.n495 9.3005
R522 source.n477 source.n476 9.3005
R523 source.n416 source.n415 9.3005
R524 source.n471 source.n470 9.3005
R525 source.n469 source.n468 9.3005
R526 source.n420 source.n419 9.3005
R527 source.n463 source.n462 9.3005
R528 source.n461 source.n460 9.3005
R529 source.n437 source.n436 9.3005
R530 source.n432 source.n431 9.3005
R531 source.n443 source.n442 9.3005
R532 source.n445 source.n444 9.3005
R533 source.n428 source.n427 9.3005
R534 source.n451 source.n450 9.3005
R535 source.n453 source.n452 9.3005
R536 source.n454 source.n423 9.3005
R537 source.n411 source.n410 9.3005
R538 source.n350 source.n349 9.3005
R539 source.n405 source.n404 9.3005
R540 source.n403 source.n402 9.3005
R541 source.n354 source.n353 9.3005
R542 source.n397 source.n396 9.3005
R543 source.n395 source.n394 9.3005
R544 source.n371 source.n370 9.3005
R545 source.n366 source.n365 9.3005
R546 source.n377 source.n376 9.3005
R547 source.n379 source.n378 9.3005
R548 source.n362 source.n361 9.3005
R549 source.n385 source.n384 9.3005
R550 source.n387 source.n386 9.3005
R551 source.n388 source.n357 9.3005
R552 source.n339 source.n338 9.3005
R553 source.n278 source.n277 9.3005
R554 source.n333 source.n332 9.3005
R555 source.n331 source.n330 9.3005
R556 source.n282 source.n281 9.3005
R557 source.n325 source.n324 9.3005
R558 source.n323 source.n322 9.3005
R559 source.n299 source.n298 9.3005
R560 source.n294 source.n293 9.3005
R561 source.n305 source.n304 9.3005
R562 source.n307 source.n306 9.3005
R563 source.n290 source.n289 9.3005
R564 source.n313 source.n312 9.3005
R565 source.n315 source.n314 9.3005
R566 source.n316 source.n285 9.3005
R567 source.n24 source.n23 9.3005
R568 source.n19 source.n18 9.3005
R569 source.n30 source.n29 9.3005
R570 source.n32 source.n31 9.3005
R571 source.n15 source.n14 9.3005
R572 source.n38 source.n37 9.3005
R573 source.n40 source.n39 9.3005
R574 source.n12 source.n9 9.3005
R575 source.n63 source.n62 9.3005
R576 source.n2 source.n1 9.3005
R577 source.n57 source.n56 9.3005
R578 source.n55 source.n54 9.3005
R579 source.n6 source.n5 9.3005
R580 source.n49 source.n48 9.3005
R581 source.n47 source.n46 9.3005
R582 source.n96 source.n95 9.3005
R583 source.n91 source.n90 9.3005
R584 source.n102 source.n101 9.3005
R585 source.n104 source.n103 9.3005
R586 source.n87 source.n86 9.3005
R587 source.n110 source.n109 9.3005
R588 source.n112 source.n111 9.3005
R589 source.n84 source.n81 9.3005
R590 source.n135 source.n134 9.3005
R591 source.n74 source.n73 9.3005
R592 source.n129 source.n128 9.3005
R593 source.n127 source.n126 9.3005
R594 source.n78 source.n77 9.3005
R595 source.n121 source.n120 9.3005
R596 source.n119 source.n118 9.3005
R597 source.n162 source.n161 9.3005
R598 source.n157 source.n156 9.3005
R599 source.n168 source.n167 9.3005
R600 source.n170 source.n169 9.3005
R601 source.n153 source.n152 9.3005
R602 source.n176 source.n175 9.3005
R603 source.n178 source.n177 9.3005
R604 source.n150 source.n147 9.3005
R605 source.n201 source.n200 9.3005
R606 source.n140 source.n139 9.3005
R607 source.n195 source.n194 9.3005
R608 source.n193 source.n192 9.3005
R609 source.n144 source.n143 9.3005
R610 source.n187 source.n186 9.3005
R611 source.n185 source.n184 9.3005
R612 source.n234 source.n233 9.3005
R613 source.n229 source.n228 9.3005
R614 source.n240 source.n239 9.3005
R615 source.n242 source.n241 9.3005
R616 source.n225 source.n224 9.3005
R617 source.n248 source.n247 9.3005
R618 source.n250 source.n249 9.3005
R619 source.n222 source.n219 9.3005
R620 source.n273 source.n272 9.3005
R621 source.n212 source.n211 9.3005
R622 source.n267 source.n266 9.3005
R623 source.n265 source.n264 9.3005
R624 source.n216 source.n215 9.3005
R625 source.n259 source.n258 9.3005
R626 source.n257 source.n256 9.3005
R627 source.n514 source.n513 8.92171
R628 source.n547 source.n488 8.92171
R629 source.n442 source.n441 8.92171
R630 source.n475 source.n416 8.92171
R631 source.n376 source.n375 8.92171
R632 source.n409 source.n350 8.92171
R633 source.n304 source.n303 8.92171
R634 source.n337 source.n278 8.92171
R635 source.n61 source.n2 8.92171
R636 source.n29 source.n28 8.92171
R637 source.n133 source.n74 8.92171
R638 source.n101 source.n100 8.92171
R639 source.n199 source.n140 8.92171
R640 source.n167 source.n166 8.92171
R641 source.n271 source.n212 8.92171
R642 source.n239 source.n238 8.92171
R643 source.n510 source.n504 8.14595
R644 source.n548 source.n486 8.14595
R645 source.n438 source.n432 8.14595
R646 source.n476 source.n414 8.14595
R647 source.n372 source.n366 8.14595
R648 source.n410 source.n348 8.14595
R649 source.n300 source.n294 8.14595
R650 source.n338 source.n276 8.14595
R651 source.n62 source.n0 8.14595
R652 source.n25 source.n19 8.14595
R653 source.n134 source.n72 8.14595
R654 source.n97 source.n91 8.14595
R655 source.n200 source.n138 8.14595
R656 source.n163 source.n157 8.14595
R657 source.n272 source.n210 8.14595
R658 source.n235 source.n229 8.14595
R659 source.n509 source.n506 7.3702
R660 source.n437 source.n434 7.3702
R661 source.n371 source.n368 7.3702
R662 source.n299 source.n296 7.3702
R663 source.n24 source.n21 7.3702
R664 source.n96 source.n93 7.3702
R665 source.n162 source.n159 7.3702
R666 source.n234 source.n231 7.3702
R667 source.n510 source.n509 5.81868
R668 source.n550 source.n486 5.81868
R669 source.n438 source.n437 5.81868
R670 source.n478 source.n414 5.81868
R671 source.n372 source.n371 5.81868
R672 source.n412 source.n348 5.81868
R673 source.n300 source.n299 5.81868
R674 source.n340 source.n276 5.81868
R675 source.n64 source.n0 5.81868
R676 source.n25 source.n24 5.81868
R677 source.n136 source.n72 5.81868
R678 source.n97 source.n96 5.81868
R679 source.n202 source.n138 5.81868
R680 source.n163 source.n162 5.81868
R681 source.n274 source.n210 5.81868
R682 source.n235 source.n234 5.81868
R683 source.n552 source.n551 5.53498
R684 source.n513 source.n504 5.04292
R685 source.n548 source.n547 5.04292
R686 source.n441 source.n432 5.04292
R687 source.n476 source.n475 5.04292
R688 source.n375 source.n366 5.04292
R689 source.n410 source.n409 5.04292
R690 source.n303 source.n294 5.04292
R691 source.n338 source.n337 5.04292
R692 source.n62 source.n61 5.04292
R693 source.n28 source.n19 5.04292
R694 source.n134 source.n133 5.04292
R695 source.n100 source.n91 5.04292
R696 source.n200 source.n199 5.04292
R697 source.n166 source.n157 5.04292
R698 source.n272 source.n271 5.04292
R699 source.n238 source.n229 5.04292
R700 source.n514 source.n502 4.26717
R701 source.n544 source.n488 4.26717
R702 source.n442 source.n430 4.26717
R703 source.n472 source.n416 4.26717
R704 source.n376 source.n364 4.26717
R705 source.n406 source.n350 4.26717
R706 source.n304 source.n292 4.26717
R707 source.n334 source.n278 4.26717
R708 source.n58 source.n2 4.26717
R709 source.n29 source.n17 4.26717
R710 source.n130 source.n74 4.26717
R711 source.n101 source.n89 4.26717
R712 source.n196 source.n140 4.26717
R713 source.n167 source.n155 4.26717
R714 source.n268 source.n212 4.26717
R715 source.n239 source.n227 4.26717
R716 source.n518 source.n517 3.49141
R717 source.n543 source.n490 3.49141
R718 source.n446 source.n445 3.49141
R719 source.n471 source.n418 3.49141
R720 source.n380 source.n379 3.49141
R721 source.n405 source.n352 3.49141
R722 source.n308 source.n307 3.49141
R723 source.n333 source.n280 3.49141
R724 source.n57 source.n4 3.49141
R725 source.n33 source.n32 3.49141
R726 source.n129 source.n76 3.49141
R727 source.n105 source.n104 3.49141
R728 source.n195 source.n142 3.49141
R729 source.n171 source.n170 3.49141
R730 source.n267 source.n214 3.49141
R731 source.n243 source.n242 3.49141
R732 source.n508 source.n507 2.84303
R733 source.n436 source.n435 2.84303
R734 source.n370 source.n369 2.84303
R735 source.n298 source.n297 2.84303
R736 source.n23 source.n22 2.84303
R737 source.n95 source.n94 2.84303
R738 source.n161 source.n160 2.84303
R739 source.n233 source.n232 2.84303
R740 source.n521 source.n500 2.71565
R741 source.n540 source.n539 2.71565
R742 source.n449 source.n428 2.71565
R743 source.n468 source.n467 2.71565
R744 source.n383 source.n362 2.71565
R745 source.n402 source.n401 2.71565
R746 source.n311 source.n290 2.71565
R747 source.n330 source.n329 2.71565
R748 source.n54 source.n53 2.71565
R749 source.n36 source.n15 2.71565
R750 source.n126 source.n125 2.71565
R751 source.n108 source.n87 2.71565
R752 source.n192 source.n191 2.71565
R753 source.n174 source.n153 2.71565
R754 source.n264 source.n263 2.71565
R755 source.n246 source.n225 2.71565
R756 source.n522 source.n498 1.93989
R757 source.n536 source.n492 1.93989
R758 source.n450 source.n426 1.93989
R759 source.n464 source.n420 1.93989
R760 source.n384 source.n360 1.93989
R761 source.n398 source.n354 1.93989
R762 source.n312 source.n288 1.93989
R763 source.n326 source.n282 1.93989
R764 source.n50 source.n6 1.93989
R765 source.n37 source.n13 1.93989
R766 source.n122 source.n78 1.93989
R767 source.n109 source.n85 1.93989
R768 source.n188 source.n144 1.93989
R769 source.n175 source.n151 1.93989
R770 source.n260 source.n216 1.93989
R771 source.n247 source.n223 1.93989
R772 source.n484 source.t19 1.6505
R773 source.n484 source.t26 1.6505
R774 source.n482 source.t22 1.6505
R775 source.n482 source.t25 1.6505
R776 source.n480 source.t21 1.6505
R777 source.n480 source.t31 1.6505
R778 source.n346 source.t15 1.6505
R779 source.n346 source.t10 1.6505
R780 source.n344 source.t3 1.6505
R781 source.n344 source.t11 1.6505
R782 source.n342 source.t9 1.6505
R783 source.n342 source.t14 1.6505
R784 source.n66 source.t2 1.6505
R785 source.n66 source.t8 1.6505
R786 source.n68 source.t12 1.6505
R787 source.n68 source.t0 1.6505
R788 source.n70 source.t5 1.6505
R789 source.n70 source.t13 1.6505
R790 source.n204 source.t28 1.6505
R791 source.n204 source.t17 1.6505
R792 source.n206 source.t18 1.6505
R793 source.n206 source.t24 1.6505
R794 source.n208 source.t27 1.6505
R795 source.n208 source.t29 1.6505
R796 source.n527 source.n525 1.16414
R797 source.n535 source.n494 1.16414
R798 source.n455 source.n453 1.16414
R799 source.n463 source.n422 1.16414
R800 source.n389 source.n387 1.16414
R801 source.n397 source.n356 1.16414
R802 source.n317 source.n315 1.16414
R803 source.n325 source.n284 1.16414
R804 source.n49 source.n8 1.16414
R805 source.n41 source.n40 1.16414
R806 source.n121 source.n80 1.16414
R807 source.n113 source.n112 1.16414
R808 source.n187 source.n146 1.16414
R809 source.n179 source.n178 1.16414
R810 source.n259 source.n218 1.16414
R811 source.n251 source.n250 1.16414
R812 source.n275 source.n209 0.543603
R813 source.n209 source.n207 0.543603
R814 source.n207 source.n205 0.543603
R815 source.n205 source.n203 0.543603
R816 source.n137 source.n71 0.543603
R817 source.n71 source.n69 0.543603
R818 source.n69 source.n67 0.543603
R819 source.n67 source.n65 0.543603
R820 source.n343 source.n341 0.543603
R821 source.n345 source.n343 0.543603
R822 source.n347 source.n345 0.543603
R823 source.n413 source.n347 0.543603
R824 source.n481 source.n479 0.543603
R825 source.n483 source.n481 0.543603
R826 source.n485 source.n483 0.543603
R827 source.n551 source.n485 0.543603
R828 source.n203 source.n137 0.470328
R829 source.n479 source.n413 0.470328
R830 source.n526 source.n496 0.388379
R831 source.n532 source.n531 0.388379
R832 source.n454 source.n424 0.388379
R833 source.n460 source.n459 0.388379
R834 source.n388 source.n358 0.388379
R835 source.n394 source.n393 0.388379
R836 source.n316 source.n286 0.388379
R837 source.n322 source.n321 0.388379
R838 source.n46 source.n45 0.388379
R839 source.n12 source.n10 0.388379
R840 source.n118 source.n117 0.388379
R841 source.n84 source.n82 0.388379
R842 source.n184 source.n183 0.388379
R843 source.n150 source.n148 0.388379
R844 source.n256 source.n255 0.388379
R845 source.n222 source.n220 0.388379
R846 source source.n552 0.188
R847 source.n508 source.n503 0.155672
R848 source.n515 source.n503 0.155672
R849 source.n516 source.n515 0.155672
R850 source.n516 source.n499 0.155672
R851 source.n523 source.n499 0.155672
R852 source.n524 source.n523 0.155672
R853 source.n524 source.n495 0.155672
R854 source.n533 source.n495 0.155672
R855 source.n534 source.n533 0.155672
R856 source.n534 source.n491 0.155672
R857 source.n541 source.n491 0.155672
R858 source.n542 source.n541 0.155672
R859 source.n542 source.n487 0.155672
R860 source.n549 source.n487 0.155672
R861 source.n436 source.n431 0.155672
R862 source.n443 source.n431 0.155672
R863 source.n444 source.n443 0.155672
R864 source.n444 source.n427 0.155672
R865 source.n451 source.n427 0.155672
R866 source.n452 source.n451 0.155672
R867 source.n452 source.n423 0.155672
R868 source.n461 source.n423 0.155672
R869 source.n462 source.n461 0.155672
R870 source.n462 source.n419 0.155672
R871 source.n469 source.n419 0.155672
R872 source.n470 source.n469 0.155672
R873 source.n470 source.n415 0.155672
R874 source.n477 source.n415 0.155672
R875 source.n370 source.n365 0.155672
R876 source.n377 source.n365 0.155672
R877 source.n378 source.n377 0.155672
R878 source.n378 source.n361 0.155672
R879 source.n385 source.n361 0.155672
R880 source.n386 source.n385 0.155672
R881 source.n386 source.n357 0.155672
R882 source.n395 source.n357 0.155672
R883 source.n396 source.n395 0.155672
R884 source.n396 source.n353 0.155672
R885 source.n403 source.n353 0.155672
R886 source.n404 source.n403 0.155672
R887 source.n404 source.n349 0.155672
R888 source.n411 source.n349 0.155672
R889 source.n298 source.n293 0.155672
R890 source.n305 source.n293 0.155672
R891 source.n306 source.n305 0.155672
R892 source.n306 source.n289 0.155672
R893 source.n313 source.n289 0.155672
R894 source.n314 source.n313 0.155672
R895 source.n314 source.n285 0.155672
R896 source.n323 source.n285 0.155672
R897 source.n324 source.n323 0.155672
R898 source.n324 source.n281 0.155672
R899 source.n331 source.n281 0.155672
R900 source.n332 source.n331 0.155672
R901 source.n332 source.n277 0.155672
R902 source.n339 source.n277 0.155672
R903 source.n63 source.n1 0.155672
R904 source.n56 source.n1 0.155672
R905 source.n56 source.n55 0.155672
R906 source.n55 source.n5 0.155672
R907 source.n48 source.n5 0.155672
R908 source.n48 source.n47 0.155672
R909 source.n47 source.n9 0.155672
R910 source.n39 source.n9 0.155672
R911 source.n39 source.n38 0.155672
R912 source.n38 source.n14 0.155672
R913 source.n31 source.n14 0.155672
R914 source.n31 source.n30 0.155672
R915 source.n30 source.n18 0.155672
R916 source.n23 source.n18 0.155672
R917 source.n135 source.n73 0.155672
R918 source.n128 source.n73 0.155672
R919 source.n128 source.n127 0.155672
R920 source.n127 source.n77 0.155672
R921 source.n120 source.n77 0.155672
R922 source.n120 source.n119 0.155672
R923 source.n119 source.n81 0.155672
R924 source.n111 source.n81 0.155672
R925 source.n111 source.n110 0.155672
R926 source.n110 source.n86 0.155672
R927 source.n103 source.n86 0.155672
R928 source.n103 source.n102 0.155672
R929 source.n102 source.n90 0.155672
R930 source.n95 source.n90 0.155672
R931 source.n201 source.n139 0.155672
R932 source.n194 source.n139 0.155672
R933 source.n194 source.n193 0.155672
R934 source.n193 source.n143 0.155672
R935 source.n186 source.n143 0.155672
R936 source.n186 source.n185 0.155672
R937 source.n185 source.n147 0.155672
R938 source.n177 source.n147 0.155672
R939 source.n177 source.n176 0.155672
R940 source.n176 source.n152 0.155672
R941 source.n169 source.n152 0.155672
R942 source.n169 source.n168 0.155672
R943 source.n168 source.n156 0.155672
R944 source.n161 source.n156 0.155672
R945 source.n273 source.n211 0.155672
R946 source.n266 source.n211 0.155672
R947 source.n266 source.n265 0.155672
R948 source.n265 source.n215 0.155672
R949 source.n258 source.n215 0.155672
R950 source.n258 source.n257 0.155672
R951 source.n257 source.n219 0.155672
R952 source.n249 source.n219 0.155672
R953 source.n249 source.n248 0.155672
R954 source.n248 source.n224 0.155672
R955 source.n241 source.n224 0.155672
R956 source.n241 source.n240 0.155672
R957 source.n240 source.n228 0.155672
R958 source.n233 source.n228 0.155672
R959 plus.n5 plus.t2 1098.38
R960 plus.n21 plus.t0 1098.38
R961 plus.n28 plus.t12 1098.38
R962 plus.n44 plus.t11 1098.38
R963 plus.n6 plus.t6 1068.43
R964 plus.n3 plus.t10 1068.43
R965 plus.n12 plus.t15 1068.43
R966 plus.n14 plus.t4 1068.43
R967 plus.n1 plus.t9 1068.43
R968 plus.n20 plus.t14 1068.43
R969 plus.n29 plus.t5 1068.43
R970 plus.n26 plus.t13 1068.43
R971 plus.n35 plus.t7 1068.43
R972 plus.n37 plus.t1 1068.43
R973 plus.n24 plus.t8 1068.43
R974 plus.n43 plus.t3 1068.43
R975 plus.n5 plus.n4 161.489
R976 plus.n28 plus.n27 161.489
R977 plus.n7 plus.n4 161.3
R978 plus.n9 plus.n8 161.3
R979 plus.n11 plus.n10 161.3
R980 plus.n13 plus.n2 161.3
R981 plus.n16 plus.n15 161.3
R982 plus.n18 plus.n17 161.3
R983 plus.n19 plus.n0 161.3
R984 plus.n22 plus.n21 161.3
R985 plus.n30 plus.n27 161.3
R986 plus.n32 plus.n31 161.3
R987 plus.n34 plus.n33 161.3
R988 plus.n36 plus.n25 161.3
R989 plus.n39 plus.n38 161.3
R990 plus.n41 plus.n40 161.3
R991 plus.n42 plus.n23 161.3
R992 plus.n45 plus.n44 161.3
R993 plus.n8 plus.n7 73.0308
R994 plus.n19 plus.n18 73.0308
R995 plus.n42 plus.n41 73.0308
R996 plus.n31 plus.n30 73.0308
R997 plus.n11 plus.n3 64.9975
R998 plus.n15 plus.n1 64.9975
R999 plus.n38 plus.n24 64.9975
R1000 plus.n34 plus.n26 64.9975
R1001 plus.n6 plus.n5 62.0763
R1002 plus.n21 plus.n20 62.0763
R1003 plus.n44 plus.n43 62.0763
R1004 plus.n29 plus.n28 62.0763
R1005 plus.n13 plus.n12 46.0096
R1006 plus.n14 plus.n13 46.0096
R1007 plus.n37 plus.n36 46.0096
R1008 plus.n36 plus.n35 46.0096
R1009 plus plus.n45 29.9763
R1010 plus.n12 plus.n11 27.0217
R1011 plus.n15 plus.n14 27.0217
R1012 plus.n38 plus.n37 27.0217
R1013 plus.n35 plus.n34 27.0217
R1014 plus plus.n22 12.1103
R1015 plus.n7 plus.n6 10.955
R1016 plus.n20 plus.n19 10.955
R1017 plus.n43 plus.n42 10.955
R1018 plus.n30 plus.n29 10.955
R1019 plus.n8 plus.n3 8.03383
R1020 plus.n18 plus.n1 8.03383
R1021 plus.n41 plus.n24 8.03383
R1022 plus.n31 plus.n26 8.03383
R1023 plus.n9 plus.n4 0.189894
R1024 plus.n10 plus.n9 0.189894
R1025 plus.n10 plus.n2 0.189894
R1026 plus.n16 plus.n2 0.189894
R1027 plus.n17 plus.n16 0.189894
R1028 plus.n17 plus.n0 0.189894
R1029 plus.n22 plus.n0 0.189894
R1030 plus.n45 plus.n23 0.189894
R1031 plus.n40 plus.n23 0.189894
R1032 plus.n40 plus.n39 0.189894
R1033 plus.n39 plus.n25 0.189894
R1034 plus.n33 plus.n25 0.189894
R1035 plus.n33 plus.n32 0.189894
R1036 plus.n32 plus.n27 0.189894
R1037 drain_left.n9 drain_left.n7 60.0958
R1038 drain_left.n5 drain_left.n3 60.0956
R1039 drain_left.n2 drain_left.n0 60.0956
R1040 drain_left.n11 drain_left.n10 59.5527
R1041 drain_left.n9 drain_left.n8 59.5527
R1042 drain_left.n5 drain_left.n4 59.5525
R1043 drain_left.n2 drain_left.n1 59.5525
R1044 drain_left.n13 drain_left.n12 59.5525
R1045 drain_left drain_left.n6 30.8972
R1046 drain_left drain_left.n13 6.19632
R1047 drain_left.n3 drain_left.t10 1.6505
R1048 drain_left.n3 drain_left.t3 1.6505
R1049 drain_left.n4 drain_left.t8 1.6505
R1050 drain_left.n4 drain_left.t2 1.6505
R1051 drain_left.n1 drain_left.t7 1.6505
R1052 drain_left.n1 drain_left.t14 1.6505
R1053 drain_left.n0 drain_left.t4 1.6505
R1054 drain_left.n0 drain_left.t12 1.6505
R1055 drain_left.n12 drain_left.t1 1.6505
R1056 drain_left.n12 drain_left.t15 1.6505
R1057 drain_left.n10 drain_left.t11 1.6505
R1058 drain_left.n10 drain_left.t6 1.6505
R1059 drain_left.n8 drain_left.t5 1.6505
R1060 drain_left.n8 drain_left.t0 1.6505
R1061 drain_left.n7 drain_left.t13 1.6505
R1062 drain_left.n7 drain_left.t9 1.6505
R1063 drain_left.n11 drain_left.n9 0.543603
R1064 drain_left.n13 drain_left.n11 0.543603
R1065 drain_left.n6 drain_left.n5 0.216706
R1066 drain_left.n6 drain_left.n2 0.216706
C0 drain_right plus 0.334364f
C1 drain_right minus 5.89809f
C2 plus source 5.60855f
C3 source minus 5.59451f
C4 drain_right source 30.4984f
C5 plus drain_left 6.0778f
C6 minus drain_left 0.171647f
C7 drain_right drain_left 0.948737f
C8 source drain_left 30.498098f
C9 plus minus 5.46309f
C10 drain_right a_n1850_n3288# 6.57855f
C11 drain_left a_n1850_n3288# 6.86706f
C12 source a_n1850_n3288# 8.717459f
C13 minus a_n1850_n3288# 7.231881f
C14 plus a_n1850_n3288# 9.22191f
C15 drain_left.t4 a_n1850_n3288# 0.322196f
C16 drain_left.t12 a_n1850_n3288# 0.322196f
C17 drain_left.n0 a_n1850_n3288# 2.87082f
C18 drain_left.t7 a_n1850_n3288# 0.322196f
C19 drain_left.t14 a_n1850_n3288# 0.322196f
C20 drain_left.n1 a_n1850_n3288# 2.86704f
C21 drain_left.n2 a_n1850_n3288# 0.78591f
C22 drain_left.t10 a_n1850_n3288# 0.322196f
C23 drain_left.t3 a_n1850_n3288# 0.322196f
C24 drain_left.n3 a_n1850_n3288# 2.87082f
C25 drain_left.t8 a_n1850_n3288# 0.322196f
C26 drain_left.t2 a_n1850_n3288# 0.322196f
C27 drain_left.n4 a_n1850_n3288# 2.86704f
C28 drain_left.n5 a_n1850_n3288# 0.78591f
C29 drain_left.n6 a_n1850_n3288# 1.66541f
C30 drain_left.t13 a_n1850_n3288# 0.322196f
C31 drain_left.t9 a_n1850_n3288# 0.322196f
C32 drain_left.n7 a_n1850_n3288# 2.87083f
C33 drain_left.t5 a_n1850_n3288# 0.322196f
C34 drain_left.t0 a_n1850_n3288# 0.322196f
C35 drain_left.n8 a_n1850_n3288# 2.86705f
C36 drain_left.n9 a_n1850_n3288# 0.818033f
C37 drain_left.t11 a_n1850_n3288# 0.322196f
C38 drain_left.t6 a_n1850_n3288# 0.322196f
C39 drain_left.n10 a_n1850_n3288# 2.86705f
C40 drain_left.n11 a_n1850_n3288# 0.404061f
C41 drain_left.t1 a_n1850_n3288# 0.322196f
C42 drain_left.t15 a_n1850_n3288# 0.322196f
C43 drain_left.n12 a_n1850_n3288# 2.86704f
C44 drain_left.n13 a_n1850_n3288# 0.686884f
C45 plus.n0 a_n1850_n3288# 0.051541f
C46 plus.t14 a_n1850_n3288# 0.524327f
C47 plus.t9 a_n1850_n3288# 0.524327f
C48 plus.n1 a_n1850_n3288# 0.207998f
C49 plus.n2 a_n1850_n3288# 0.051541f
C50 plus.t4 a_n1850_n3288# 0.524327f
C51 plus.t15 a_n1850_n3288# 0.524327f
C52 plus.t10 a_n1850_n3288# 0.524327f
C53 plus.n3 a_n1850_n3288# 0.207998f
C54 plus.n4 a_n1850_n3288# 0.109688f
C55 plus.t6 a_n1850_n3288# 0.524327f
C56 plus.t2 a_n1850_n3288# 0.530002f
C57 plus.n5 a_n1850_n3288# 0.223779f
C58 plus.n6 a_n1850_n3288# 0.207998f
C59 plus.n7 a_n1850_n3288# 0.019481f
C60 plus.n8 a_n1850_n3288# 0.018846f
C61 plus.n9 a_n1850_n3288# 0.051541f
C62 plus.n10 a_n1850_n3288# 0.051541f
C63 plus.n11 a_n1850_n3288# 0.021229f
C64 plus.n12 a_n1850_n3288# 0.207998f
C65 plus.n13 a_n1850_n3288# 0.021229f
C66 plus.n14 a_n1850_n3288# 0.207998f
C67 plus.n15 a_n1850_n3288# 0.021229f
C68 plus.n16 a_n1850_n3288# 0.051541f
C69 plus.n17 a_n1850_n3288# 0.051541f
C70 plus.n18 a_n1850_n3288# 0.018846f
C71 plus.n19 a_n1850_n3288# 0.019481f
C72 plus.n20 a_n1850_n3288# 0.207998f
C73 plus.t0 a_n1850_n3288# 0.530002f
C74 plus.n21 a_n1850_n3288# 0.223711f
C75 plus.n22 a_n1850_n3288# 0.572526f
C76 plus.n23 a_n1850_n3288# 0.051541f
C77 plus.t11 a_n1850_n3288# 0.530002f
C78 plus.t3 a_n1850_n3288# 0.524327f
C79 plus.t8 a_n1850_n3288# 0.524327f
C80 plus.n24 a_n1850_n3288# 0.207998f
C81 plus.n25 a_n1850_n3288# 0.051541f
C82 plus.t1 a_n1850_n3288# 0.524327f
C83 plus.t7 a_n1850_n3288# 0.524327f
C84 plus.t13 a_n1850_n3288# 0.524327f
C85 plus.n26 a_n1850_n3288# 0.207998f
C86 plus.n27 a_n1850_n3288# 0.109688f
C87 plus.t5 a_n1850_n3288# 0.524327f
C88 plus.t12 a_n1850_n3288# 0.530002f
C89 plus.n28 a_n1850_n3288# 0.223779f
C90 plus.n29 a_n1850_n3288# 0.207998f
C91 plus.n30 a_n1850_n3288# 0.019481f
C92 plus.n31 a_n1850_n3288# 0.018846f
C93 plus.n32 a_n1850_n3288# 0.051541f
C94 plus.n33 a_n1850_n3288# 0.051541f
C95 plus.n34 a_n1850_n3288# 0.021229f
C96 plus.n35 a_n1850_n3288# 0.207998f
C97 plus.n36 a_n1850_n3288# 0.021229f
C98 plus.n37 a_n1850_n3288# 0.207998f
C99 plus.n38 a_n1850_n3288# 0.021229f
C100 plus.n39 a_n1850_n3288# 0.051541f
C101 plus.n40 a_n1850_n3288# 0.051541f
C102 plus.n41 a_n1850_n3288# 0.018846f
C103 plus.n42 a_n1850_n3288# 0.019481f
C104 plus.n43 a_n1850_n3288# 0.207998f
C105 plus.n44 a_n1850_n3288# 0.223711f
C106 plus.n45 a_n1850_n3288# 1.53201f
C107 source.n0 a_n1850_n3288# 0.037637f
C108 source.n1 a_n1850_n3288# 0.028413f
C109 source.n2 a_n1850_n3288# 0.015268f
C110 source.n3 a_n1850_n3288# 0.036088f
C111 source.n4 a_n1850_n3288# 0.016166f
C112 source.n5 a_n1850_n3288# 0.028413f
C113 source.n6 a_n1850_n3288# 0.015268f
C114 source.n7 a_n1850_n3288# 0.036088f
C115 source.n8 a_n1850_n3288# 0.016166f
C116 source.n9 a_n1850_n3288# 0.028413f
C117 source.n10 a_n1850_n3288# 0.015717f
C118 source.n11 a_n1850_n3288# 0.036088f
C119 source.n12 a_n1850_n3288# 0.015268f
C120 source.n13 a_n1850_n3288# 0.016166f
C121 source.n14 a_n1850_n3288# 0.028413f
C122 source.n15 a_n1850_n3288# 0.015268f
C123 source.n16 a_n1850_n3288# 0.036088f
C124 source.n17 a_n1850_n3288# 0.016166f
C125 source.n18 a_n1850_n3288# 0.028413f
C126 source.n19 a_n1850_n3288# 0.015268f
C127 source.n20 a_n1850_n3288# 0.027066f
C128 source.n21 a_n1850_n3288# 0.025511f
C129 source.t1 a_n1850_n3288# 0.06095f
C130 source.n22 a_n1850_n3288# 0.204856f
C131 source.n23 a_n1850_n3288# 1.4334f
C132 source.n24 a_n1850_n3288# 0.015268f
C133 source.n25 a_n1850_n3288# 0.016166f
C134 source.n26 a_n1850_n3288# 0.036088f
C135 source.n27 a_n1850_n3288# 0.036088f
C136 source.n28 a_n1850_n3288# 0.016166f
C137 source.n29 a_n1850_n3288# 0.015268f
C138 source.n30 a_n1850_n3288# 0.028413f
C139 source.n31 a_n1850_n3288# 0.028413f
C140 source.n32 a_n1850_n3288# 0.015268f
C141 source.n33 a_n1850_n3288# 0.016166f
C142 source.n34 a_n1850_n3288# 0.036088f
C143 source.n35 a_n1850_n3288# 0.036088f
C144 source.n36 a_n1850_n3288# 0.016166f
C145 source.n37 a_n1850_n3288# 0.015268f
C146 source.n38 a_n1850_n3288# 0.028413f
C147 source.n39 a_n1850_n3288# 0.028413f
C148 source.n40 a_n1850_n3288# 0.015268f
C149 source.n41 a_n1850_n3288# 0.016166f
C150 source.n42 a_n1850_n3288# 0.036088f
C151 source.n43 a_n1850_n3288# 0.036088f
C152 source.n44 a_n1850_n3288# 0.036088f
C153 source.n45 a_n1850_n3288# 0.015717f
C154 source.n46 a_n1850_n3288# 0.015268f
C155 source.n47 a_n1850_n3288# 0.028413f
C156 source.n48 a_n1850_n3288# 0.028413f
C157 source.n49 a_n1850_n3288# 0.015268f
C158 source.n50 a_n1850_n3288# 0.016166f
C159 source.n51 a_n1850_n3288# 0.036088f
C160 source.n52 a_n1850_n3288# 0.036088f
C161 source.n53 a_n1850_n3288# 0.016166f
C162 source.n54 a_n1850_n3288# 0.015268f
C163 source.n55 a_n1850_n3288# 0.028413f
C164 source.n56 a_n1850_n3288# 0.028413f
C165 source.n57 a_n1850_n3288# 0.015268f
C166 source.n58 a_n1850_n3288# 0.016166f
C167 source.n59 a_n1850_n3288# 0.036088f
C168 source.n60 a_n1850_n3288# 0.074057f
C169 source.n61 a_n1850_n3288# 0.016166f
C170 source.n62 a_n1850_n3288# 0.015268f
C171 source.n63 a_n1850_n3288# 0.061018f
C172 source.n64 a_n1850_n3288# 0.040871f
C173 source.n65 a_n1850_n3288# 1.14349f
C174 source.t2 a_n1850_n3288# 0.269436f
C175 source.t8 a_n1850_n3288# 0.269436f
C176 source.n66 a_n1850_n3288# 2.30692f
C177 source.n67 a_n1850_n3288# 0.389935f
C178 source.t12 a_n1850_n3288# 0.269436f
C179 source.t0 a_n1850_n3288# 0.269436f
C180 source.n68 a_n1850_n3288# 2.30692f
C181 source.n69 a_n1850_n3288# 0.389935f
C182 source.t5 a_n1850_n3288# 0.269436f
C183 source.t13 a_n1850_n3288# 0.269436f
C184 source.n70 a_n1850_n3288# 2.30692f
C185 source.n71 a_n1850_n3288# 0.389935f
C186 source.n72 a_n1850_n3288# 0.037637f
C187 source.n73 a_n1850_n3288# 0.028413f
C188 source.n74 a_n1850_n3288# 0.015268f
C189 source.n75 a_n1850_n3288# 0.036088f
C190 source.n76 a_n1850_n3288# 0.016166f
C191 source.n77 a_n1850_n3288# 0.028413f
C192 source.n78 a_n1850_n3288# 0.015268f
C193 source.n79 a_n1850_n3288# 0.036088f
C194 source.n80 a_n1850_n3288# 0.016166f
C195 source.n81 a_n1850_n3288# 0.028413f
C196 source.n82 a_n1850_n3288# 0.015717f
C197 source.n83 a_n1850_n3288# 0.036088f
C198 source.n84 a_n1850_n3288# 0.015268f
C199 source.n85 a_n1850_n3288# 0.016166f
C200 source.n86 a_n1850_n3288# 0.028413f
C201 source.n87 a_n1850_n3288# 0.015268f
C202 source.n88 a_n1850_n3288# 0.036088f
C203 source.n89 a_n1850_n3288# 0.016166f
C204 source.n90 a_n1850_n3288# 0.028413f
C205 source.n91 a_n1850_n3288# 0.015268f
C206 source.n92 a_n1850_n3288# 0.027066f
C207 source.n93 a_n1850_n3288# 0.025511f
C208 source.t6 a_n1850_n3288# 0.06095f
C209 source.n94 a_n1850_n3288# 0.204856f
C210 source.n95 a_n1850_n3288# 1.4334f
C211 source.n96 a_n1850_n3288# 0.015268f
C212 source.n97 a_n1850_n3288# 0.016166f
C213 source.n98 a_n1850_n3288# 0.036088f
C214 source.n99 a_n1850_n3288# 0.036088f
C215 source.n100 a_n1850_n3288# 0.016166f
C216 source.n101 a_n1850_n3288# 0.015268f
C217 source.n102 a_n1850_n3288# 0.028413f
C218 source.n103 a_n1850_n3288# 0.028413f
C219 source.n104 a_n1850_n3288# 0.015268f
C220 source.n105 a_n1850_n3288# 0.016166f
C221 source.n106 a_n1850_n3288# 0.036088f
C222 source.n107 a_n1850_n3288# 0.036088f
C223 source.n108 a_n1850_n3288# 0.016166f
C224 source.n109 a_n1850_n3288# 0.015268f
C225 source.n110 a_n1850_n3288# 0.028413f
C226 source.n111 a_n1850_n3288# 0.028413f
C227 source.n112 a_n1850_n3288# 0.015268f
C228 source.n113 a_n1850_n3288# 0.016166f
C229 source.n114 a_n1850_n3288# 0.036088f
C230 source.n115 a_n1850_n3288# 0.036088f
C231 source.n116 a_n1850_n3288# 0.036088f
C232 source.n117 a_n1850_n3288# 0.015717f
C233 source.n118 a_n1850_n3288# 0.015268f
C234 source.n119 a_n1850_n3288# 0.028413f
C235 source.n120 a_n1850_n3288# 0.028413f
C236 source.n121 a_n1850_n3288# 0.015268f
C237 source.n122 a_n1850_n3288# 0.016166f
C238 source.n123 a_n1850_n3288# 0.036088f
C239 source.n124 a_n1850_n3288# 0.036088f
C240 source.n125 a_n1850_n3288# 0.016166f
C241 source.n126 a_n1850_n3288# 0.015268f
C242 source.n127 a_n1850_n3288# 0.028413f
C243 source.n128 a_n1850_n3288# 0.028413f
C244 source.n129 a_n1850_n3288# 0.015268f
C245 source.n130 a_n1850_n3288# 0.016166f
C246 source.n131 a_n1850_n3288# 0.036088f
C247 source.n132 a_n1850_n3288# 0.074057f
C248 source.n133 a_n1850_n3288# 0.016166f
C249 source.n134 a_n1850_n3288# 0.015268f
C250 source.n135 a_n1850_n3288# 0.061018f
C251 source.n136 a_n1850_n3288# 0.040871f
C252 source.n137 a_n1850_n3288# 0.114381f
C253 source.n138 a_n1850_n3288# 0.037637f
C254 source.n139 a_n1850_n3288# 0.028413f
C255 source.n140 a_n1850_n3288# 0.015268f
C256 source.n141 a_n1850_n3288# 0.036088f
C257 source.n142 a_n1850_n3288# 0.016166f
C258 source.n143 a_n1850_n3288# 0.028413f
C259 source.n144 a_n1850_n3288# 0.015268f
C260 source.n145 a_n1850_n3288# 0.036088f
C261 source.n146 a_n1850_n3288# 0.016166f
C262 source.n147 a_n1850_n3288# 0.028413f
C263 source.n148 a_n1850_n3288# 0.015717f
C264 source.n149 a_n1850_n3288# 0.036088f
C265 source.n150 a_n1850_n3288# 0.015268f
C266 source.n151 a_n1850_n3288# 0.016166f
C267 source.n152 a_n1850_n3288# 0.028413f
C268 source.n153 a_n1850_n3288# 0.015268f
C269 source.n154 a_n1850_n3288# 0.036088f
C270 source.n155 a_n1850_n3288# 0.016166f
C271 source.n156 a_n1850_n3288# 0.028413f
C272 source.n157 a_n1850_n3288# 0.015268f
C273 source.n158 a_n1850_n3288# 0.027066f
C274 source.n159 a_n1850_n3288# 0.025511f
C275 source.t23 a_n1850_n3288# 0.06095f
C276 source.n160 a_n1850_n3288# 0.204856f
C277 source.n161 a_n1850_n3288# 1.4334f
C278 source.n162 a_n1850_n3288# 0.015268f
C279 source.n163 a_n1850_n3288# 0.016166f
C280 source.n164 a_n1850_n3288# 0.036088f
C281 source.n165 a_n1850_n3288# 0.036088f
C282 source.n166 a_n1850_n3288# 0.016166f
C283 source.n167 a_n1850_n3288# 0.015268f
C284 source.n168 a_n1850_n3288# 0.028413f
C285 source.n169 a_n1850_n3288# 0.028413f
C286 source.n170 a_n1850_n3288# 0.015268f
C287 source.n171 a_n1850_n3288# 0.016166f
C288 source.n172 a_n1850_n3288# 0.036088f
C289 source.n173 a_n1850_n3288# 0.036088f
C290 source.n174 a_n1850_n3288# 0.016166f
C291 source.n175 a_n1850_n3288# 0.015268f
C292 source.n176 a_n1850_n3288# 0.028413f
C293 source.n177 a_n1850_n3288# 0.028413f
C294 source.n178 a_n1850_n3288# 0.015268f
C295 source.n179 a_n1850_n3288# 0.016166f
C296 source.n180 a_n1850_n3288# 0.036088f
C297 source.n181 a_n1850_n3288# 0.036088f
C298 source.n182 a_n1850_n3288# 0.036088f
C299 source.n183 a_n1850_n3288# 0.015717f
C300 source.n184 a_n1850_n3288# 0.015268f
C301 source.n185 a_n1850_n3288# 0.028413f
C302 source.n186 a_n1850_n3288# 0.028413f
C303 source.n187 a_n1850_n3288# 0.015268f
C304 source.n188 a_n1850_n3288# 0.016166f
C305 source.n189 a_n1850_n3288# 0.036088f
C306 source.n190 a_n1850_n3288# 0.036088f
C307 source.n191 a_n1850_n3288# 0.016166f
C308 source.n192 a_n1850_n3288# 0.015268f
C309 source.n193 a_n1850_n3288# 0.028413f
C310 source.n194 a_n1850_n3288# 0.028413f
C311 source.n195 a_n1850_n3288# 0.015268f
C312 source.n196 a_n1850_n3288# 0.016166f
C313 source.n197 a_n1850_n3288# 0.036088f
C314 source.n198 a_n1850_n3288# 0.074057f
C315 source.n199 a_n1850_n3288# 0.016166f
C316 source.n200 a_n1850_n3288# 0.015268f
C317 source.n201 a_n1850_n3288# 0.061018f
C318 source.n202 a_n1850_n3288# 0.040871f
C319 source.n203 a_n1850_n3288# 0.114381f
C320 source.t28 a_n1850_n3288# 0.269436f
C321 source.t17 a_n1850_n3288# 0.269436f
C322 source.n204 a_n1850_n3288# 2.30692f
C323 source.n205 a_n1850_n3288# 0.389935f
C324 source.t18 a_n1850_n3288# 0.269436f
C325 source.t24 a_n1850_n3288# 0.269436f
C326 source.n206 a_n1850_n3288# 2.30692f
C327 source.n207 a_n1850_n3288# 0.389935f
C328 source.t27 a_n1850_n3288# 0.269436f
C329 source.t29 a_n1850_n3288# 0.269436f
C330 source.n208 a_n1850_n3288# 2.30692f
C331 source.n209 a_n1850_n3288# 0.389935f
C332 source.n210 a_n1850_n3288# 0.037637f
C333 source.n211 a_n1850_n3288# 0.028413f
C334 source.n212 a_n1850_n3288# 0.015268f
C335 source.n213 a_n1850_n3288# 0.036088f
C336 source.n214 a_n1850_n3288# 0.016166f
C337 source.n215 a_n1850_n3288# 0.028413f
C338 source.n216 a_n1850_n3288# 0.015268f
C339 source.n217 a_n1850_n3288# 0.036088f
C340 source.n218 a_n1850_n3288# 0.016166f
C341 source.n219 a_n1850_n3288# 0.028413f
C342 source.n220 a_n1850_n3288# 0.015717f
C343 source.n221 a_n1850_n3288# 0.036088f
C344 source.n222 a_n1850_n3288# 0.015268f
C345 source.n223 a_n1850_n3288# 0.016166f
C346 source.n224 a_n1850_n3288# 0.028413f
C347 source.n225 a_n1850_n3288# 0.015268f
C348 source.n226 a_n1850_n3288# 0.036088f
C349 source.n227 a_n1850_n3288# 0.016166f
C350 source.n228 a_n1850_n3288# 0.028413f
C351 source.n229 a_n1850_n3288# 0.015268f
C352 source.n230 a_n1850_n3288# 0.027066f
C353 source.n231 a_n1850_n3288# 0.025511f
C354 source.t16 a_n1850_n3288# 0.06095f
C355 source.n232 a_n1850_n3288# 0.204856f
C356 source.n233 a_n1850_n3288# 1.4334f
C357 source.n234 a_n1850_n3288# 0.015268f
C358 source.n235 a_n1850_n3288# 0.016166f
C359 source.n236 a_n1850_n3288# 0.036088f
C360 source.n237 a_n1850_n3288# 0.036088f
C361 source.n238 a_n1850_n3288# 0.016166f
C362 source.n239 a_n1850_n3288# 0.015268f
C363 source.n240 a_n1850_n3288# 0.028413f
C364 source.n241 a_n1850_n3288# 0.028413f
C365 source.n242 a_n1850_n3288# 0.015268f
C366 source.n243 a_n1850_n3288# 0.016166f
C367 source.n244 a_n1850_n3288# 0.036088f
C368 source.n245 a_n1850_n3288# 0.036088f
C369 source.n246 a_n1850_n3288# 0.016166f
C370 source.n247 a_n1850_n3288# 0.015268f
C371 source.n248 a_n1850_n3288# 0.028413f
C372 source.n249 a_n1850_n3288# 0.028413f
C373 source.n250 a_n1850_n3288# 0.015268f
C374 source.n251 a_n1850_n3288# 0.016166f
C375 source.n252 a_n1850_n3288# 0.036088f
C376 source.n253 a_n1850_n3288# 0.036088f
C377 source.n254 a_n1850_n3288# 0.036088f
C378 source.n255 a_n1850_n3288# 0.015717f
C379 source.n256 a_n1850_n3288# 0.015268f
C380 source.n257 a_n1850_n3288# 0.028413f
C381 source.n258 a_n1850_n3288# 0.028413f
C382 source.n259 a_n1850_n3288# 0.015268f
C383 source.n260 a_n1850_n3288# 0.016166f
C384 source.n261 a_n1850_n3288# 0.036088f
C385 source.n262 a_n1850_n3288# 0.036088f
C386 source.n263 a_n1850_n3288# 0.016166f
C387 source.n264 a_n1850_n3288# 0.015268f
C388 source.n265 a_n1850_n3288# 0.028413f
C389 source.n266 a_n1850_n3288# 0.028413f
C390 source.n267 a_n1850_n3288# 0.015268f
C391 source.n268 a_n1850_n3288# 0.016166f
C392 source.n269 a_n1850_n3288# 0.036088f
C393 source.n270 a_n1850_n3288# 0.074057f
C394 source.n271 a_n1850_n3288# 0.016166f
C395 source.n272 a_n1850_n3288# 0.015268f
C396 source.n273 a_n1850_n3288# 0.061018f
C397 source.n274 a_n1850_n3288# 0.040871f
C398 source.n275 a_n1850_n3288# 1.59026f
C399 source.n276 a_n1850_n3288# 0.037637f
C400 source.n277 a_n1850_n3288# 0.028413f
C401 source.n278 a_n1850_n3288# 0.015268f
C402 source.n279 a_n1850_n3288# 0.036088f
C403 source.n280 a_n1850_n3288# 0.016166f
C404 source.n281 a_n1850_n3288# 0.028413f
C405 source.n282 a_n1850_n3288# 0.015268f
C406 source.n283 a_n1850_n3288# 0.036088f
C407 source.n284 a_n1850_n3288# 0.016166f
C408 source.n285 a_n1850_n3288# 0.028413f
C409 source.n286 a_n1850_n3288# 0.015717f
C410 source.n287 a_n1850_n3288# 0.036088f
C411 source.n288 a_n1850_n3288# 0.016166f
C412 source.n289 a_n1850_n3288# 0.028413f
C413 source.n290 a_n1850_n3288# 0.015268f
C414 source.n291 a_n1850_n3288# 0.036088f
C415 source.n292 a_n1850_n3288# 0.016166f
C416 source.n293 a_n1850_n3288# 0.028413f
C417 source.n294 a_n1850_n3288# 0.015268f
C418 source.n295 a_n1850_n3288# 0.027066f
C419 source.n296 a_n1850_n3288# 0.025511f
C420 source.t4 a_n1850_n3288# 0.06095f
C421 source.n297 a_n1850_n3288# 0.204856f
C422 source.n298 a_n1850_n3288# 1.4334f
C423 source.n299 a_n1850_n3288# 0.015268f
C424 source.n300 a_n1850_n3288# 0.016166f
C425 source.n301 a_n1850_n3288# 0.036088f
C426 source.n302 a_n1850_n3288# 0.036088f
C427 source.n303 a_n1850_n3288# 0.016166f
C428 source.n304 a_n1850_n3288# 0.015268f
C429 source.n305 a_n1850_n3288# 0.028413f
C430 source.n306 a_n1850_n3288# 0.028413f
C431 source.n307 a_n1850_n3288# 0.015268f
C432 source.n308 a_n1850_n3288# 0.016166f
C433 source.n309 a_n1850_n3288# 0.036088f
C434 source.n310 a_n1850_n3288# 0.036088f
C435 source.n311 a_n1850_n3288# 0.016166f
C436 source.n312 a_n1850_n3288# 0.015268f
C437 source.n313 a_n1850_n3288# 0.028413f
C438 source.n314 a_n1850_n3288# 0.028413f
C439 source.n315 a_n1850_n3288# 0.015268f
C440 source.n316 a_n1850_n3288# 0.015268f
C441 source.n317 a_n1850_n3288# 0.016166f
C442 source.n318 a_n1850_n3288# 0.036088f
C443 source.n319 a_n1850_n3288# 0.036088f
C444 source.n320 a_n1850_n3288# 0.036088f
C445 source.n321 a_n1850_n3288# 0.015717f
C446 source.n322 a_n1850_n3288# 0.015268f
C447 source.n323 a_n1850_n3288# 0.028413f
C448 source.n324 a_n1850_n3288# 0.028413f
C449 source.n325 a_n1850_n3288# 0.015268f
C450 source.n326 a_n1850_n3288# 0.016166f
C451 source.n327 a_n1850_n3288# 0.036088f
C452 source.n328 a_n1850_n3288# 0.036088f
C453 source.n329 a_n1850_n3288# 0.016166f
C454 source.n330 a_n1850_n3288# 0.015268f
C455 source.n331 a_n1850_n3288# 0.028413f
C456 source.n332 a_n1850_n3288# 0.028413f
C457 source.n333 a_n1850_n3288# 0.015268f
C458 source.n334 a_n1850_n3288# 0.016166f
C459 source.n335 a_n1850_n3288# 0.036088f
C460 source.n336 a_n1850_n3288# 0.074057f
C461 source.n337 a_n1850_n3288# 0.016166f
C462 source.n338 a_n1850_n3288# 0.015268f
C463 source.n339 a_n1850_n3288# 0.061018f
C464 source.n340 a_n1850_n3288# 0.040871f
C465 source.n341 a_n1850_n3288# 1.59026f
C466 source.t9 a_n1850_n3288# 0.269436f
C467 source.t14 a_n1850_n3288# 0.269436f
C468 source.n342 a_n1850_n3288# 2.3069f
C469 source.n343 a_n1850_n3288# 0.389949f
C470 source.t3 a_n1850_n3288# 0.269436f
C471 source.t11 a_n1850_n3288# 0.269436f
C472 source.n344 a_n1850_n3288# 2.3069f
C473 source.n345 a_n1850_n3288# 0.389949f
C474 source.t15 a_n1850_n3288# 0.269436f
C475 source.t10 a_n1850_n3288# 0.269436f
C476 source.n346 a_n1850_n3288# 2.3069f
C477 source.n347 a_n1850_n3288# 0.389949f
C478 source.n348 a_n1850_n3288# 0.037637f
C479 source.n349 a_n1850_n3288# 0.028413f
C480 source.n350 a_n1850_n3288# 0.015268f
C481 source.n351 a_n1850_n3288# 0.036088f
C482 source.n352 a_n1850_n3288# 0.016166f
C483 source.n353 a_n1850_n3288# 0.028413f
C484 source.n354 a_n1850_n3288# 0.015268f
C485 source.n355 a_n1850_n3288# 0.036088f
C486 source.n356 a_n1850_n3288# 0.016166f
C487 source.n357 a_n1850_n3288# 0.028413f
C488 source.n358 a_n1850_n3288# 0.015717f
C489 source.n359 a_n1850_n3288# 0.036088f
C490 source.n360 a_n1850_n3288# 0.016166f
C491 source.n361 a_n1850_n3288# 0.028413f
C492 source.n362 a_n1850_n3288# 0.015268f
C493 source.n363 a_n1850_n3288# 0.036088f
C494 source.n364 a_n1850_n3288# 0.016166f
C495 source.n365 a_n1850_n3288# 0.028413f
C496 source.n366 a_n1850_n3288# 0.015268f
C497 source.n367 a_n1850_n3288# 0.027066f
C498 source.n368 a_n1850_n3288# 0.025511f
C499 source.t7 a_n1850_n3288# 0.06095f
C500 source.n369 a_n1850_n3288# 0.204856f
C501 source.n370 a_n1850_n3288# 1.4334f
C502 source.n371 a_n1850_n3288# 0.015268f
C503 source.n372 a_n1850_n3288# 0.016166f
C504 source.n373 a_n1850_n3288# 0.036088f
C505 source.n374 a_n1850_n3288# 0.036088f
C506 source.n375 a_n1850_n3288# 0.016166f
C507 source.n376 a_n1850_n3288# 0.015268f
C508 source.n377 a_n1850_n3288# 0.028413f
C509 source.n378 a_n1850_n3288# 0.028413f
C510 source.n379 a_n1850_n3288# 0.015268f
C511 source.n380 a_n1850_n3288# 0.016166f
C512 source.n381 a_n1850_n3288# 0.036088f
C513 source.n382 a_n1850_n3288# 0.036088f
C514 source.n383 a_n1850_n3288# 0.016166f
C515 source.n384 a_n1850_n3288# 0.015268f
C516 source.n385 a_n1850_n3288# 0.028413f
C517 source.n386 a_n1850_n3288# 0.028413f
C518 source.n387 a_n1850_n3288# 0.015268f
C519 source.n388 a_n1850_n3288# 0.015268f
C520 source.n389 a_n1850_n3288# 0.016166f
C521 source.n390 a_n1850_n3288# 0.036088f
C522 source.n391 a_n1850_n3288# 0.036088f
C523 source.n392 a_n1850_n3288# 0.036088f
C524 source.n393 a_n1850_n3288# 0.015717f
C525 source.n394 a_n1850_n3288# 0.015268f
C526 source.n395 a_n1850_n3288# 0.028413f
C527 source.n396 a_n1850_n3288# 0.028413f
C528 source.n397 a_n1850_n3288# 0.015268f
C529 source.n398 a_n1850_n3288# 0.016166f
C530 source.n399 a_n1850_n3288# 0.036088f
C531 source.n400 a_n1850_n3288# 0.036088f
C532 source.n401 a_n1850_n3288# 0.016166f
C533 source.n402 a_n1850_n3288# 0.015268f
C534 source.n403 a_n1850_n3288# 0.028413f
C535 source.n404 a_n1850_n3288# 0.028413f
C536 source.n405 a_n1850_n3288# 0.015268f
C537 source.n406 a_n1850_n3288# 0.016166f
C538 source.n407 a_n1850_n3288# 0.036088f
C539 source.n408 a_n1850_n3288# 0.074057f
C540 source.n409 a_n1850_n3288# 0.016166f
C541 source.n410 a_n1850_n3288# 0.015268f
C542 source.n411 a_n1850_n3288# 0.061018f
C543 source.n412 a_n1850_n3288# 0.040871f
C544 source.n413 a_n1850_n3288# 0.114381f
C545 source.n414 a_n1850_n3288# 0.037637f
C546 source.n415 a_n1850_n3288# 0.028413f
C547 source.n416 a_n1850_n3288# 0.015268f
C548 source.n417 a_n1850_n3288# 0.036088f
C549 source.n418 a_n1850_n3288# 0.016166f
C550 source.n419 a_n1850_n3288# 0.028413f
C551 source.n420 a_n1850_n3288# 0.015268f
C552 source.n421 a_n1850_n3288# 0.036088f
C553 source.n422 a_n1850_n3288# 0.016166f
C554 source.n423 a_n1850_n3288# 0.028413f
C555 source.n424 a_n1850_n3288# 0.015717f
C556 source.n425 a_n1850_n3288# 0.036088f
C557 source.n426 a_n1850_n3288# 0.016166f
C558 source.n427 a_n1850_n3288# 0.028413f
C559 source.n428 a_n1850_n3288# 0.015268f
C560 source.n429 a_n1850_n3288# 0.036088f
C561 source.n430 a_n1850_n3288# 0.016166f
C562 source.n431 a_n1850_n3288# 0.028413f
C563 source.n432 a_n1850_n3288# 0.015268f
C564 source.n433 a_n1850_n3288# 0.027066f
C565 source.n434 a_n1850_n3288# 0.025511f
C566 source.t30 a_n1850_n3288# 0.06095f
C567 source.n435 a_n1850_n3288# 0.204856f
C568 source.n436 a_n1850_n3288# 1.4334f
C569 source.n437 a_n1850_n3288# 0.015268f
C570 source.n438 a_n1850_n3288# 0.016166f
C571 source.n439 a_n1850_n3288# 0.036088f
C572 source.n440 a_n1850_n3288# 0.036088f
C573 source.n441 a_n1850_n3288# 0.016166f
C574 source.n442 a_n1850_n3288# 0.015268f
C575 source.n443 a_n1850_n3288# 0.028413f
C576 source.n444 a_n1850_n3288# 0.028413f
C577 source.n445 a_n1850_n3288# 0.015268f
C578 source.n446 a_n1850_n3288# 0.016166f
C579 source.n447 a_n1850_n3288# 0.036088f
C580 source.n448 a_n1850_n3288# 0.036088f
C581 source.n449 a_n1850_n3288# 0.016166f
C582 source.n450 a_n1850_n3288# 0.015268f
C583 source.n451 a_n1850_n3288# 0.028413f
C584 source.n452 a_n1850_n3288# 0.028413f
C585 source.n453 a_n1850_n3288# 0.015268f
C586 source.n454 a_n1850_n3288# 0.015268f
C587 source.n455 a_n1850_n3288# 0.016166f
C588 source.n456 a_n1850_n3288# 0.036088f
C589 source.n457 a_n1850_n3288# 0.036088f
C590 source.n458 a_n1850_n3288# 0.036088f
C591 source.n459 a_n1850_n3288# 0.015717f
C592 source.n460 a_n1850_n3288# 0.015268f
C593 source.n461 a_n1850_n3288# 0.028413f
C594 source.n462 a_n1850_n3288# 0.028413f
C595 source.n463 a_n1850_n3288# 0.015268f
C596 source.n464 a_n1850_n3288# 0.016166f
C597 source.n465 a_n1850_n3288# 0.036088f
C598 source.n466 a_n1850_n3288# 0.036088f
C599 source.n467 a_n1850_n3288# 0.016166f
C600 source.n468 a_n1850_n3288# 0.015268f
C601 source.n469 a_n1850_n3288# 0.028413f
C602 source.n470 a_n1850_n3288# 0.028413f
C603 source.n471 a_n1850_n3288# 0.015268f
C604 source.n472 a_n1850_n3288# 0.016166f
C605 source.n473 a_n1850_n3288# 0.036088f
C606 source.n474 a_n1850_n3288# 0.074057f
C607 source.n475 a_n1850_n3288# 0.016166f
C608 source.n476 a_n1850_n3288# 0.015268f
C609 source.n477 a_n1850_n3288# 0.061018f
C610 source.n478 a_n1850_n3288# 0.040871f
C611 source.n479 a_n1850_n3288# 0.114381f
C612 source.t21 a_n1850_n3288# 0.269436f
C613 source.t31 a_n1850_n3288# 0.269436f
C614 source.n480 a_n1850_n3288# 2.3069f
C615 source.n481 a_n1850_n3288# 0.389949f
C616 source.t22 a_n1850_n3288# 0.269436f
C617 source.t25 a_n1850_n3288# 0.269436f
C618 source.n482 a_n1850_n3288# 2.3069f
C619 source.n483 a_n1850_n3288# 0.389949f
C620 source.t19 a_n1850_n3288# 0.269436f
C621 source.t26 a_n1850_n3288# 0.269436f
C622 source.n484 a_n1850_n3288# 2.3069f
C623 source.n485 a_n1850_n3288# 0.389949f
C624 source.n486 a_n1850_n3288# 0.037637f
C625 source.n487 a_n1850_n3288# 0.028413f
C626 source.n488 a_n1850_n3288# 0.015268f
C627 source.n489 a_n1850_n3288# 0.036088f
C628 source.n490 a_n1850_n3288# 0.016166f
C629 source.n491 a_n1850_n3288# 0.028413f
C630 source.n492 a_n1850_n3288# 0.015268f
C631 source.n493 a_n1850_n3288# 0.036088f
C632 source.n494 a_n1850_n3288# 0.016166f
C633 source.n495 a_n1850_n3288# 0.028413f
C634 source.n496 a_n1850_n3288# 0.015717f
C635 source.n497 a_n1850_n3288# 0.036088f
C636 source.n498 a_n1850_n3288# 0.016166f
C637 source.n499 a_n1850_n3288# 0.028413f
C638 source.n500 a_n1850_n3288# 0.015268f
C639 source.n501 a_n1850_n3288# 0.036088f
C640 source.n502 a_n1850_n3288# 0.016166f
C641 source.n503 a_n1850_n3288# 0.028413f
C642 source.n504 a_n1850_n3288# 0.015268f
C643 source.n505 a_n1850_n3288# 0.027066f
C644 source.n506 a_n1850_n3288# 0.025511f
C645 source.t20 a_n1850_n3288# 0.06095f
C646 source.n507 a_n1850_n3288# 0.204856f
C647 source.n508 a_n1850_n3288# 1.4334f
C648 source.n509 a_n1850_n3288# 0.015268f
C649 source.n510 a_n1850_n3288# 0.016166f
C650 source.n511 a_n1850_n3288# 0.036088f
C651 source.n512 a_n1850_n3288# 0.036088f
C652 source.n513 a_n1850_n3288# 0.016166f
C653 source.n514 a_n1850_n3288# 0.015268f
C654 source.n515 a_n1850_n3288# 0.028413f
C655 source.n516 a_n1850_n3288# 0.028413f
C656 source.n517 a_n1850_n3288# 0.015268f
C657 source.n518 a_n1850_n3288# 0.016166f
C658 source.n519 a_n1850_n3288# 0.036088f
C659 source.n520 a_n1850_n3288# 0.036088f
C660 source.n521 a_n1850_n3288# 0.016166f
C661 source.n522 a_n1850_n3288# 0.015268f
C662 source.n523 a_n1850_n3288# 0.028413f
C663 source.n524 a_n1850_n3288# 0.028413f
C664 source.n525 a_n1850_n3288# 0.015268f
C665 source.n526 a_n1850_n3288# 0.015268f
C666 source.n527 a_n1850_n3288# 0.016166f
C667 source.n528 a_n1850_n3288# 0.036088f
C668 source.n529 a_n1850_n3288# 0.036088f
C669 source.n530 a_n1850_n3288# 0.036088f
C670 source.n531 a_n1850_n3288# 0.015717f
C671 source.n532 a_n1850_n3288# 0.015268f
C672 source.n533 a_n1850_n3288# 0.028413f
C673 source.n534 a_n1850_n3288# 0.028413f
C674 source.n535 a_n1850_n3288# 0.015268f
C675 source.n536 a_n1850_n3288# 0.016166f
C676 source.n537 a_n1850_n3288# 0.036088f
C677 source.n538 a_n1850_n3288# 0.036088f
C678 source.n539 a_n1850_n3288# 0.016166f
C679 source.n540 a_n1850_n3288# 0.015268f
C680 source.n541 a_n1850_n3288# 0.028413f
C681 source.n542 a_n1850_n3288# 0.028413f
C682 source.n543 a_n1850_n3288# 0.015268f
C683 source.n544 a_n1850_n3288# 0.016166f
C684 source.n545 a_n1850_n3288# 0.036088f
C685 source.n546 a_n1850_n3288# 0.074057f
C686 source.n547 a_n1850_n3288# 0.016166f
C687 source.n548 a_n1850_n3288# 0.015268f
C688 source.n549 a_n1850_n3288# 0.061018f
C689 source.n550 a_n1850_n3288# 0.040871f
C690 source.n551 a_n1850_n3288# 0.274773f
C691 source.n552 a_n1850_n3288# 1.78248f
C692 drain_right.t11 a_n1850_n3288# 0.321603f
C693 drain_right.t7 a_n1850_n3288# 0.321603f
C694 drain_right.n0 a_n1850_n3288# 2.86554f
C695 drain_right.t13 a_n1850_n3288# 0.321603f
C696 drain_right.t4 a_n1850_n3288# 0.321603f
C697 drain_right.n1 a_n1850_n3288# 2.86177f
C698 drain_right.n2 a_n1850_n3288# 0.784465f
C699 drain_right.t14 a_n1850_n3288# 0.321603f
C700 drain_right.t0 a_n1850_n3288# 0.321603f
C701 drain_right.n3 a_n1850_n3288# 2.86554f
C702 drain_right.t15 a_n1850_n3288# 0.321603f
C703 drain_right.t1 a_n1850_n3288# 0.321603f
C704 drain_right.n4 a_n1850_n3288# 2.86177f
C705 drain_right.n5 a_n1850_n3288# 0.784465f
C706 drain_right.n6 a_n1850_n3288# 1.59202f
C707 drain_right.t2 a_n1850_n3288# 0.321603f
C708 drain_right.t12 a_n1850_n3288# 0.321603f
C709 drain_right.n7 a_n1850_n3288# 2.86554f
C710 drain_right.t9 a_n1850_n3288# 0.321603f
C711 drain_right.t10 a_n1850_n3288# 0.321603f
C712 drain_right.n8 a_n1850_n3288# 2.86178f
C713 drain_right.n9 a_n1850_n3288# 0.816539f
C714 drain_right.t3 a_n1850_n3288# 0.321603f
C715 drain_right.t5 a_n1850_n3288# 0.321603f
C716 drain_right.n10 a_n1850_n3288# 2.86178f
C717 drain_right.n11 a_n1850_n3288# 0.403318f
C718 drain_right.t6 a_n1850_n3288# 0.321603f
C719 drain_right.t8 a_n1850_n3288# 0.321603f
C720 drain_right.n12 a_n1850_n3288# 2.86178f
C721 drain_right.n13 a_n1850_n3288# 0.685609f
C722 minus.n0 a_n1850_n3288# 0.050635f
C723 minus.t15 a_n1850_n3288# 0.520684f
C724 minus.t4 a_n1850_n3288# 0.515109f
C725 minus.t2 a_n1850_n3288# 0.515109f
C726 minus.n1 a_n1850_n3288# 0.204341f
C727 minus.n2 a_n1850_n3288# 0.050635f
C728 minus.t13 a_n1850_n3288# 0.515109f
C729 minus.t7 a_n1850_n3288# 0.515109f
C730 minus.t3 a_n1850_n3288# 0.515109f
C731 minus.n3 a_n1850_n3288# 0.204341f
C732 minus.n4 a_n1850_n3288# 0.107759f
C733 minus.t14 a_n1850_n3288# 0.515109f
C734 minus.t8 a_n1850_n3288# 0.520684f
C735 minus.n5 a_n1850_n3288# 0.219845f
C736 minus.n6 a_n1850_n3288# 0.204341f
C737 minus.n7 a_n1850_n3288# 0.019139f
C738 minus.n8 a_n1850_n3288# 0.018514f
C739 minus.n9 a_n1850_n3288# 0.050635f
C740 minus.n10 a_n1850_n3288# 0.050635f
C741 minus.n11 a_n1850_n3288# 0.020856f
C742 minus.n12 a_n1850_n3288# 0.204341f
C743 minus.n13 a_n1850_n3288# 0.020856f
C744 minus.n14 a_n1850_n3288# 0.204341f
C745 minus.n15 a_n1850_n3288# 0.020856f
C746 minus.n16 a_n1850_n3288# 0.050635f
C747 minus.n17 a_n1850_n3288# 0.050635f
C748 minus.n18 a_n1850_n3288# 0.018514f
C749 minus.n19 a_n1850_n3288# 0.019139f
C750 minus.n20 a_n1850_n3288# 0.204341f
C751 minus.n21 a_n1850_n3288# 0.219778f
C752 minus.n22 a_n1850_n3288# 1.78057f
C753 minus.n23 a_n1850_n3288# 0.050635f
C754 minus.t5 a_n1850_n3288# 0.515109f
C755 minus.t12 a_n1850_n3288# 0.515109f
C756 minus.n24 a_n1850_n3288# 0.204341f
C757 minus.n25 a_n1850_n3288# 0.050635f
C758 minus.t6 a_n1850_n3288# 0.515109f
C759 minus.t9 a_n1850_n3288# 0.515109f
C760 minus.t0 a_n1850_n3288# 0.515109f
C761 minus.n26 a_n1850_n3288# 0.204341f
C762 minus.n27 a_n1850_n3288# 0.107759f
C763 minus.t10 a_n1850_n3288# 0.515109f
C764 minus.t1 a_n1850_n3288# 0.520684f
C765 minus.n28 a_n1850_n3288# 0.219845f
C766 minus.n29 a_n1850_n3288# 0.204341f
C767 minus.n30 a_n1850_n3288# 0.019139f
C768 minus.n31 a_n1850_n3288# 0.018514f
C769 minus.n32 a_n1850_n3288# 0.050635f
C770 minus.n33 a_n1850_n3288# 0.050635f
C771 minus.n34 a_n1850_n3288# 0.020856f
C772 minus.n35 a_n1850_n3288# 0.204341f
C773 minus.n36 a_n1850_n3288# 0.020856f
C774 minus.n37 a_n1850_n3288# 0.204341f
C775 minus.n38 a_n1850_n3288# 0.020856f
C776 minus.n39 a_n1850_n3288# 0.050635f
C777 minus.n40 a_n1850_n3288# 0.050635f
C778 minus.n41 a_n1850_n3288# 0.018514f
C779 minus.n42 a_n1850_n3288# 0.019139f
C780 minus.n43 a_n1850_n3288# 0.204341f
C781 minus.t11 a_n1850_n3288# 0.520684f
C782 minus.n44 a_n1850_n3288# 0.219778f
C783 minus.n45 a_n1850_n3288# 0.327026f
C784 minus.n46 a_n1850_n3288# 2.16489f
.ends

