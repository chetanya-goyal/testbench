* NGSPICE file created from diffpair585.ext - technology: sky130A

.subckt diffpair585 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t21 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X1 drain_left.t10 plus.t1 source.t19 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X2 drain_left.t9 plus.t2 source.t13 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X3 drain_right.t11 minus.t0 source.t4 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X4 source.t1 minus.t1 drain_right.t10 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X5 source.t7 minus.t2 drain_right.t9 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X6 source.t9 minus.t3 drain_right.t8 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X7 source.t12 plus.t3 drain_left.t8 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X8 a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X9 a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X10 source.t17 plus.t4 drain_left.t7 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X11 drain_right.t7 minus.t4 source.t8 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X12 source.t2 minus.t5 drain_right.t6 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X13 drain_left.t6 plus.t5 source.t18 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X14 source.t5 minus.t6 drain_right.t5 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X15 source.t20 plus.t6 drain_left.t5 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X16 source.t11 plus.t7 drain_left.t4 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X17 a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X18 drain_left.t3 plus.t8 source.t10 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X19 a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X20 drain_right.t4 minus.t7 source.t6 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X21 drain_right.t3 minus.t8 source.t0 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X22 drain_right.t2 minus.t9 source.t3 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X23 drain_right.t1 minus.t10 source.t22 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X24 source.t16 plus.t9 drain_left.t2 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X25 source.t23 minus.t11 drain_right.t0 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X26 drain_left.t1 plus.t10 source.t15 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X27 source.t14 plus.t11 drain_left.t0 a_n1528_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
R0 plus.n2 plus.t4 2082.53
R1 plus.n13 plus.t10 2082.53
R2 plus.n17 plus.t2 2082.53
R3 plus.n28 plus.t11 2082.53
R4 plus.n3 plus.t1 2053.32
R5 plus.n4 plus.t7 2053.32
R6 plus.n10 plus.t0 2053.32
R7 plus.n12 plus.t6 2053.32
R8 plus.n19 plus.t9 2053.32
R9 plus.n18 plus.t8 2053.32
R10 plus.n25 plus.t3 2053.32
R11 plus.n27 plus.t5 2053.32
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 67.1884
R27 plus.n11 plus.n10 67.1884
R28 plus.n26 plus.n25 67.1884
R29 plus.n20 plus.n18 67.1884
R30 plus.n3 plus.n2 55.5035
R31 plus.n13 plus.n12 55.5035
R32 plus.n28 plus.n27 55.5035
R33 plus.n19 plus.n17 55.5035
R34 plus plus.n29 31.7566
R35 plus.n5 plus.n3 17.5278
R36 plus.n12 plus.n11 17.5278
R37 plus.n27 plus.n26 17.5278
R38 plus.n20 plus.n19 17.5278
R39 plus plus.n14 15.1103
R40 plus.n4 plus.n1 5.84292
R41 plus.n10 plus.n9 5.84292
R42 plus.n25 plus.n24 5.84292
R43 plus.n18 plus.n16 5.84292
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n0 source.t15 44.1297
R53 source.n5 source.t17 44.1296
R54 source.n6 source.t0 44.1296
R55 source.n11 source.t2 44.1296
R56 source.n23 source.t4 44.1295
R57 source.n18 source.t7 44.1295
R58 source.n17 source.t13 44.1295
R59 source.n12 source.t14 44.1295
R60 source.n2 source.n1 43.1397
R61 source.n4 source.n3 43.1397
R62 source.n8 source.n7 43.1397
R63 source.n10 source.n9 43.1397
R64 source.n22 source.n21 43.1396
R65 source.n20 source.n19 43.1396
R66 source.n16 source.n15 43.1396
R67 source.n14 source.n13 43.1396
R68 source.n12 source.n11 27.8483
R69 source.n24 source.n0 22.3354
R70 source.n24 source.n23 5.51343
R71 source.n21 source.t3 0.9905
R72 source.n21 source.t5 0.9905
R73 source.n19 source.t8 0.9905
R74 source.n19 source.t23 0.9905
R75 source.n15 source.t10 0.9905
R76 source.n15 source.t16 0.9905
R77 source.n13 source.t18 0.9905
R78 source.n13 source.t12 0.9905
R79 source.n1 source.t21 0.9905
R80 source.n1 source.t20 0.9905
R81 source.n3 source.t19 0.9905
R82 source.n3 source.t11 0.9905
R83 source.n7 source.t6 0.9905
R84 source.n7 source.t9 0.9905
R85 source.n9 source.t22 0.9905
R86 source.n9 source.t1 0.9905
R87 source.n11 source.n10 0.5005
R88 source.n10 source.n8 0.5005
R89 source.n8 source.n6 0.5005
R90 source.n5 source.n4 0.5005
R91 source.n4 source.n2 0.5005
R92 source.n2 source.n0 0.5005
R93 source.n14 source.n12 0.5005
R94 source.n16 source.n14 0.5005
R95 source.n17 source.n16 0.5005
R96 source.n20 source.n18 0.5005
R97 source.n22 source.n20 0.5005
R98 source.n23 source.n22 0.5005
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 60.3185
R103 drain_left.n3 drain_left.n2 60.2631
R104 drain_left.n3 drain_left.n0 60.2631
R105 drain_left.n8 drain_left.n7 59.8185
R106 drain_left.n6 drain_left.n5 59.8185
R107 drain_left.n3 drain_left.n1 59.8184
R108 drain_left drain_left.n3 35.9277
R109 drain_left drain_left.n8 6.15322
R110 drain_left.n1 drain_left.t8 0.9905
R111 drain_left.n1 drain_left.t3 0.9905
R112 drain_left.n2 drain_left.t2 0.9905
R113 drain_left.n2 drain_left.t9 0.9905
R114 drain_left.n0 drain_left.t0 0.9905
R115 drain_left.n0 drain_left.t6 0.9905
R116 drain_left.n7 drain_left.t5 0.9905
R117 drain_left.n7 drain_left.t1 0.9905
R118 drain_left.n5 drain_left.t4 0.9905
R119 drain_left.n5 drain_left.t11 0.9905
R120 drain_left.n4 drain_left.t7 0.9905
R121 drain_left.n4 drain_left.t10 0.9905
R122 drain_left.n8 drain_left.n6 0.5005
R123 minus.n13 minus.t5 2082.53
R124 minus.n2 minus.t8 2082.53
R125 minus.n28 minus.t0 2082.53
R126 minus.n17 minus.t2 2082.53
R127 minus.n12 minus.t10 2053.32
R128 minus.n10 minus.t1 2053.32
R129 minus.n3 minus.t7 2053.32
R130 minus.n4 minus.t3 2053.32
R131 minus.n27 minus.t6 2053.32
R132 minus.n25 minus.t9 2053.32
R133 minus.n19 minus.t11 2053.32
R134 minus.n18 minus.t4 2053.32
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 67.1884
R150 minus.n5 minus.n3 67.1884
R151 minus.n20 minus.n19 67.1884
R152 minus.n26 minus.n25 67.1884
R153 minus.n13 minus.n12 55.5035
R154 minus.n4 minus.n2 55.5035
R155 minus.n18 minus.n17 55.5035
R156 minus.n28 minus.n27 55.5035
R157 minus.n30 minus.n14 40.9058
R158 minus.n12 minus.n11 17.5278
R159 minus.n5 minus.n4 17.5278
R160 minus.n20 minus.n18 17.5278
R161 minus.n27 minus.n26 17.5278
R162 minus.n30 minus.n29 6.43611
R163 minus.n10 minus.n9 5.84292
R164 minus.n3 minus.n1 5.84292
R165 minus.n19 minus.n16 5.84292
R166 minus.n25 minus.n24 5.84292
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 60.3185
R177 drain_right.n3 drain_right.n2 60.2631
R178 drain_right.n3 drain_right.n0 60.2631
R179 drain_right.n6 drain_right.n5 59.8185
R180 drain_right.n8 drain_right.n7 59.8185
R181 drain_right.n3 drain_right.n1 59.8184
R182 drain_right drain_right.n3 35.3745
R183 drain_right drain_right.n8 6.15322
R184 drain_right.n1 drain_right.t0 0.9905
R185 drain_right.n1 drain_right.t2 0.9905
R186 drain_right.n2 drain_right.t5 0.9905
R187 drain_right.n2 drain_right.t11 0.9905
R188 drain_right.n0 drain_right.t9 0.9905
R189 drain_right.n0 drain_right.t7 0.9905
R190 drain_right.n4 drain_right.t8 0.9905
R191 drain_right.n4 drain_right.t3 0.9905
R192 drain_right.n5 drain_right.t10 0.9905
R193 drain_right.n5 drain_right.t4 0.9905
R194 drain_right.n7 drain_right.t6 0.9905
R195 drain_right.n7 drain_right.t1 0.9905
R196 drain_right.n8 drain_right.n6 0.5005
C0 minus drain_left 0.171004f
C1 plus drain_left 6.68092f
C2 minus drain_right 6.53476f
C3 plus drain_right 0.300071f
C4 source drain_left 41.122604f
C5 minus plus 6.54371f
C6 source drain_right 41.121998f
C7 source minus 5.77816f
C8 source plus 5.7922f
C9 drain_right drain_left 0.751086f
C10 drain_right a_n1528_n4888# 8.03215f
C11 drain_left a_n1528_n4888# 8.284349f
C12 source a_n1528_n4888# 12.874455f
C13 minus a_n1528_n4888# 6.461996f
C14 plus a_n1528_n4888# 9.039419f
C15 drain_right.t9 a_n1528_n4888# 0.569182f
C16 drain_right.t7 a_n1528_n4888# 0.569182f
C17 drain_right.n0 a_n1528_n4888# 5.20676f
C18 drain_right.t0 a_n1528_n4888# 0.569182f
C19 drain_right.t2 a_n1528_n4888# 0.569182f
C20 drain_right.n1 a_n1528_n4888# 5.20359f
C21 drain_right.t5 a_n1528_n4888# 0.569182f
C22 drain_right.t11 a_n1528_n4888# 0.569182f
C23 drain_right.n2 a_n1528_n4888# 5.20676f
C24 drain_right.n3 a_n1528_n4888# 3.49285f
C25 drain_right.t8 a_n1528_n4888# 0.569182f
C26 drain_right.t3 a_n1528_n4888# 0.569182f
C27 drain_right.n4 a_n1528_n4888# 5.207181f
C28 drain_right.t10 a_n1528_n4888# 0.569182f
C29 drain_right.t4 a_n1528_n4888# 0.569182f
C30 drain_right.n5 a_n1528_n4888# 5.20358f
C31 drain_right.n6 a_n1528_n4888# 0.850815f
C32 drain_right.t6 a_n1528_n4888# 0.569182f
C33 drain_right.t1 a_n1528_n4888# 0.569182f
C34 drain_right.n7 a_n1528_n4888# 5.20358f
C35 drain_right.n8 a_n1528_n4888# 0.717224f
C36 minus.n0 a_n1528_n4888# 0.054099f
C37 minus.t5 a_n1528_n4888# 0.765826f
C38 minus.t10 a_n1528_n4888# 0.761841f
C39 minus.t1 a_n1528_n4888# 0.761841f
C40 minus.n1 a_n1528_n4888# 0.019281f
C41 minus.t8 a_n1528_n4888# 0.765826f
C42 minus.n2 a_n1528_n4888# 0.300816f
C43 minus.t7 a_n1528_n4888# 0.761841f
C44 minus.n3 a_n1528_n4888# 0.285785f
C45 minus.t3 a_n1528_n4888# 0.761841f
C46 minus.n4 a_n1528_n4888# 0.285785f
C47 minus.n5 a_n1528_n4888# 0.020615f
C48 minus.n6 a_n1528_n4888# 0.113131f
C49 minus.n7 a_n1528_n4888# 0.054099f
C50 minus.n8 a_n1528_n4888# 0.054099f
C51 minus.n9 a_n1528_n4888# 0.019281f
C52 minus.n10 a_n1528_n4888# 0.285785f
C53 minus.n11 a_n1528_n4888# 0.020615f
C54 minus.n12 a_n1528_n4888# 0.285785f
C55 minus.n13 a_n1528_n4888# 0.300747f
C56 minus.n14 a_n1528_n4888# 2.30169f
C57 minus.n15 a_n1528_n4888# 0.054099f
C58 minus.t6 a_n1528_n4888# 0.761841f
C59 minus.t9 a_n1528_n4888# 0.761841f
C60 minus.n16 a_n1528_n4888# 0.019281f
C61 minus.t2 a_n1528_n4888# 0.765826f
C62 minus.n17 a_n1528_n4888# 0.300816f
C63 minus.t4 a_n1528_n4888# 0.761841f
C64 minus.n18 a_n1528_n4888# 0.285785f
C65 minus.t11 a_n1528_n4888# 0.761841f
C66 minus.n19 a_n1528_n4888# 0.285785f
C67 minus.n20 a_n1528_n4888# 0.020615f
C68 minus.n21 a_n1528_n4888# 0.113131f
C69 minus.n22 a_n1528_n4888# 0.054099f
C70 minus.n23 a_n1528_n4888# 0.054099f
C71 minus.n24 a_n1528_n4888# 0.019281f
C72 minus.n25 a_n1528_n4888# 0.285785f
C73 minus.n26 a_n1528_n4888# 0.020615f
C74 minus.n27 a_n1528_n4888# 0.285785f
C75 minus.t0 a_n1528_n4888# 0.765826f
C76 minus.n28 a_n1528_n4888# 0.300747f
C77 minus.n29 a_n1528_n4888# 0.345516f
C78 minus.n30 a_n1528_n4888# 2.75939f
C79 drain_left.t0 a_n1528_n4888# 0.569887f
C80 drain_left.t6 a_n1528_n4888# 0.569887f
C81 drain_left.n0 a_n1528_n4888# 5.21321f
C82 drain_left.t8 a_n1528_n4888# 0.569887f
C83 drain_left.t3 a_n1528_n4888# 0.569887f
C84 drain_left.n1 a_n1528_n4888# 5.21003f
C85 drain_left.t2 a_n1528_n4888# 0.569887f
C86 drain_left.t9 a_n1528_n4888# 0.569887f
C87 drain_left.n2 a_n1528_n4888# 5.21321f
C88 drain_left.n3 a_n1528_n4888# 3.57259f
C89 drain_left.t7 a_n1528_n4888# 0.569887f
C90 drain_left.t10 a_n1528_n4888# 0.569887f
C91 drain_left.n4 a_n1528_n4888# 5.21363f
C92 drain_left.t4 a_n1528_n4888# 0.569887f
C93 drain_left.t11 a_n1528_n4888# 0.569887f
C94 drain_left.n5 a_n1528_n4888# 5.21002f
C95 drain_left.n6 a_n1528_n4888# 0.851868f
C96 drain_left.t5 a_n1528_n4888# 0.569887f
C97 drain_left.t1 a_n1528_n4888# 0.569887f
C98 drain_left.n7 a_n1528_n4888# 5.21002f
C99 drain_left.n8 a_n1528_n4888# 0.718112f
C100 source.t15 a_n1528_n4888# 5.00607f
C101 source.n0 a_n1528_n4888# 2.12318f
C102 source.t21 a_n1528_n4888# 0.438039f
C103 source.t20 a_n1528_n4888# 0.438039f
C104 source.n1 a_n1528_n4888# 3.91625f
C105 source.n2 a_n1528_n4888# 0.373911f
C106 source.t19 a_n1528_n4888# 0.438039f
C107 source.t11 a_n1528_n4888# 0.438039f
C108 source.n3 a_n1528_n4888# 3.91625f
C109 source.n4 a_n1528_n4888# 0.373911f
C110 source.t17 a_n1528_n4888# 5.00609f
C111 source.n5 a_n1528_n4888# 0.476037f
C112 source.t0 a_n1528_n4888# 5.00609f
C113 source.n6 a_n1528_n4888# 0.476037f
C114 source.t6 a_n1528_n4888# 0.438039f
C115 source.t9 a_n1528_n4888# 0.438039f
C116 source.n7 a_n1528_n4888# 3.91625f
C117 source.n8 a_n1528_n4888# 0.373911f
C118 source.t22 a_n1528_n4888# 0.438039f
C119 source.t1 a_n1528_n4888# 0.438039f
C120 source.n9 a_n1528_n4888# 3.91625f
C121 source.n10 a_n1528_n4888# 0.373911f
C122 source.t2 a_n1528_n4888# 5.00609f
C123 source.n11 a_n1528_n4888# 2.61271f
C124 source.t14 a_n1528_n4888# 5.00606f
C125 source.n12 a_n1528_n4888# 2.61274f
C126 source.t18 a_n1528_n4888# 0.438039f
C127 source.t12 a_n1528_n4888# 0.438039f
C128 source.n13 a_n1528_n4888# 3.91626f
C129 source.n14 a_n1528_n4888# 0.373903f
C130 source.t10 a_n1528_n4888# 0.438039f
C131 source.t16 a_n1528_n4888# 0.438039f
C132 source.n15 a_n1528_n4888# 3.91626f
C133 source.n16 a_n1528_n4888# 0.373903f
C134 source.t13 a_n1528_n4888# 5.00606f
C135 source.n17 a_n1528_n4888# 0.476065f
C136 source.t7 a_n1528_n4888# 5.00606f
C137 source.n18 a_n1528_n4888# 0.476065f
C138 source.t8 a_n1528_n4888# 0.438039f
C139 source.t23 a_n1528_n4888# 0.438039f
C140 source.n19 a_n1528_n4888# 3.91626f
C141 source.n20 a_n1528_n4888# 0.373903f
C142 source.t3 a_n1528_n4888# 0.438039f
C143 source.t5 a_n1528_n4888# 0.438039f
C144 source.n21 a_n1528_n4888# 3.91626f
C145 source.n22 a_n1528_n4888# 0.373903f
C146 source.t4 a_n1528_n4888# 5.00606f
C147 source.n23 a_n1528_n4888# 0.62944f
C148 source.n24 a_n1528_n4888# 2.49255f
C149 plus.n0 a_n1528_n4888# 0.054994f
C150 plus.t6 a_n1528_n4888# 0.774452f
C151 plus.t0 a_n1528_n4888# 0.774452f
C152 plus.n1 a_n1528_n4888# 0.0196f
C153 plus.t4 a_n1528_n4888# 0.778504f
C154 plus.n2 a_n1528_n4888# 0.305796f
C155 plus.t1 a_n1528_n4888# 0.774452f
C156 plus.n3 a_n1528_n4888# 0.290516f
C157 plus.t7 a_n1528_n4888# 0.774452f
C158 plus.n4 a_n1528_n4888# 0.290516f
C159 plus.n5 a_n1528_n4888# 0.020956f
C160 plus.n6 a_n1528_n4888# 0.115004f
C161 plus.n7 a_n1528_n4888# 0.054994f
C162 plus.n8 a_n1528_n4888# 0.054994f
C163 plus.n9 a_n1528_n4888# 0.0196f
C164 plus.n10 a_n1528_n4888# 0.290516f
C165 plus.n11 a_n1528_n4888# 0.020956f
C166 plus.n12 a_n1528_n4888# 0.290516f
C167 plus.t10 a_n1528_n4888# 0.778504f
C168 plus.n13 a_n1528_n4888# 0.305725f
C169 plus.n14 a_n1528_n4888# 0.826959f
C170 plus.n15 a_n1528_n4888# 0.054994f
C171 plus.t11 a_n1528_n4888# 0.778504f
C172 plus.t5 a_n1528_n4888# 0.774452f
C173 plus.t3 a_n1528_n4888# 0.774452f
C174 plus.n16 a_n1528_n4888# 0.0196f
C175 plus.t2 a_n1528_n4888# 0.778504f
C176 plus.n17 a_n1528_n4888# 0.305796f
C177 plus.t8 a_n1528_n4888# 0.774452f
C178 plus.n18 a_n1528_n4888# 0.290516f
C179 plus.t9 a_n1528_n4888# 0.774452f
C180 plus.n19 a_n1528_n4888# 0.290516f
C181 plus.n20 a_n1528_n4888# 0.020956f
C182 plus.n21 a_n1528_n4888# 0.115004f
C183 plus.n22 a_n1528_n4888# 0.054994f
C184 plus.n23 a_n1528_n4888# 0.054994f
C185 plus.n24 a_n1528_n4888# 0.0196f
C186 plus.n25 a_n1528_n4888# 0.290516f
C187 plus.n26 a_n1528_n4888# 0.020956f
C188 plus.n27 a_n1528_n4888# 0.290516f
C189 plus.n28 a_n1528_n4888# 0.305725f
C190 plus.n29 a_n1528_n4888# 1.84064f
.ends

