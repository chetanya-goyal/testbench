* NGSPICE file created from diffpair637.ext - technology: sky130A

.subckt diffpair637 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t18 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X2 source.t0 minus.t0 drain_right.t15 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X3 source.t1 minus.t1 drain_right.t14 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X4 source.t17 plus.t1 drain_left.t14 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X5 drain_right.t13 minus.t2 source.t5 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X6 a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X7 source.t16 plus.t2 drain_left.t13 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X8 drain_right.t12 minus.t3 source.t9 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 drain_right.t11 minus.t4 source.t10 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 source.t25 plus.t3 drain_left.t12 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X11 drain_right.t10 minus.t5 source.t6 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 source.t11 minus.t6 drain_right.t9 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X13 source.t21 plus.t4 drain_left.t11 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X14 drain_right.t8 minus.t7 source.t15 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X15 drain_right.t7 minus.t8 source.t7 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X16 drain_right.t6 minus.t9 source.t14 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_left.t10 plus.t5 source.t30 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X18 a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X19 source.t3 minus.t10 drain_right.t5 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 drain_left.t9 plus.t6 source.t28 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X21 source.t12 minus.t11 drain_right.t4 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X22 drain_right.t3 minus.t12 source.t13 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X23 source.t27 plus.t7 drain_left.t8 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X24 drain_left.t7 plus.t8 source.t20 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X25 drain_left.t6 plus.t9 source.t31 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X26 source.t8 minus.t13 drain_right.t2 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X27 source.t23 plus.t10 drain_left.t5 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X28 drain_left.t4 plus.t11 source.t24 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X29 a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X30 drain_left.t3 plus.t12 source.t19 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X31 source.t26 plus.t13 drain_left.t2 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X32 drain_left.t1 plus.t14 source.t22 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X33 source.t2 minus.t14 drain_right.t1 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X34 source.t4 minus.t15 drain_right.t0 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X35 source.t29 plus.t15 drain_left.t0 a_n2750_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n7 plus.t15 672.628
R1 plus.n29 plus.t0 672.628
R2 plus.n20 plus.t6 651.605
R3 plus.n18 plus.t7 651.605
R4 plus.n17 plus.t8 651.605
R5 plus.n3 plus.t13 651.605
R6 plus.n11 plus.t9 651.605
R7 plus.n5 plus.t10 651.605
R8 plus.n6 plus.t14 651.605
R9 plus.n42 plus.t2 651.605
R10 plus.n40 plus.t5 651.605
R11 plus.n39 plus.t1 651.605
R12 plus.n25 plus.t11 651.605
R13 plus.n33 plus.t3 651.605
R14 plus.n27 plus.t12 651.605
R15 plus.n28 plus.t4 651.605
R16 plus.n10 plus.n9 161.3
R17 plus.n11 plus.n4 161.3
R18 plus.n13 plus.n12 161.3
R19 plus.n14 plus.n3 161.3
R20 plus.n16 plus.n15 161.3
R21 plus.n19 plus.n0 161.3
R22 plus.n21 plus.n20 161.3
R23 plus.n32 plus.n31 161.3
R24 plus.n33 plus.n26 161.3
R25 plus.n35 plus.n34 161.3
R26 plus.n36 plus.n25 161.3
R27 plus.n38 plus.n37 161.3
R28 plus.n41 plus.n22 161.3
R29 plus.n43 plus.n42 161.3
R30 plus.n8 plus.n5 80.6037
R31 plus.n17 plus.n2 80.6037
R32 plus.n18 plus.n1 80.6037
R33 plus.n30 plus.n27 80.6037
R34 plus.n39 plus.n24 80.6037
R35 plus.n40 plus.n23 80.6037
R36 plus.n18 plus.n17 48.2005
R37 plus.n6 plus.n5 48.2005
R38 plus.n40 plus.n39 48.2005
R39 plus.n28 plus.n27 48.2005
R40 plus.n17 plus.n16 43.0884
R41 plus.n10 plus.n5 43.0884
R42 plus.n39 plus.n38 43.0884
R43 plus.n32 plus.n27 43.0884
R44 plus.n19 plus.n18 40.1672
R45 plus.n41 plus.n40 40.1672
R46 plus plus.n43 36.6051
R47 plus.n8 plus.n7 31.6481
R48 plus.n30 plus.n29 31.6481
R49 plus.n12 plus.n11 24.1005
R50 plus.n12 plus.n3 24.1005
R51 plus.n34 plus.n25 24.1005
R52 plus.n34 plus.n33 24.1005
R53 plus.n7 plus.n6 17.444
R54 plus.n29 plus.n28 17.444
R55 plus plus.n21 15.33
R56 plus.n20 plus.n19 8.03383
R57 plus.n42 plus.n41 8.03383
R58 plus.n16 plus.n3 5.11262
R59 plus.n11 plus.n10 5.11262
R60 plus.n38 plus.n25 5.11262
R61 plus.n33 plus.n32 5.11262
R62 plus.n2 plus.n1 0.380177
R63 plus.n24 plus.n23 0.380177
R64 plus.n9 plus.n8 0.285035
R65 plus.n15 plus.n2 0.285035
R66 plus.n1 plus.n0 0.285035
R67 plus.n23 plus.n22 0.285035
R68 plus.n37 plus.n24 0.285035
R69 plus.n31 plus.n30 0.285035
R70 plus.n9 plus.n4 0.189894
R71 plus.n13 plus.n4 0.189894
R72 plus.n14 plus.n13 0.189894
R73 plus.n15 plus.n14 0.189894
R74 plus.n21 plus.n0 0.189894
R75 plus.n43 plus.n22 0.189894
R76 plus.n37 plus.n36 0.189894
R77 plus.n36 plus.n35 0.189894
R78 plus.n35 plus.n26 0.189894
R79 plus.n31 plus.n26 0.189894
R80 source.n0 source.t28 44.1297
R81 source.n7 source.t29 44.1296
R82 source.n8 source.t7 44.1296
R83 source.n15 source.t8 44.1296
R84 source.n31 source.t5 44.1295
R85 source.n24 source.t1 44.1295
R86 source.n23 source.t18 44.1295
R87 source.n16 source.t16 44.1295
R88 source.n2 source.n1 43.1397
R89 source.n4 source.n3 43.1397
R90 source.n6 source.n5 43.1397
R91 source.n10 source.n9 43.1397
R92 source.n12 source.n11 43.1397
R93 source.n14 source.n13 43.1397
R94 source.n30 source.n29 43.1396
R95 source.n28 source.n27 43.1396
R96 source.n26 source.n25 43.1396
R97 source.n22 source.n21 43.1396
R98 source.n20 source.n19 43.1396
R99 source.n18 source.n17 43.1396
R100 source.n16 source.n15 28.3225
R101 source.n32 source.n0 22.5725
R102 source.n32 source.n31 5.7505
R103 source.n29 source.t9 0.9905
R104 source.n29 source.t2 0.9905
R105 source.n27 source.t10 0.9905
R106 source.n27 source.t0 0.9905
R107 source.n25 source.t14 0.9905
R108 source.n25 source.t4 0.9905
R109 source.n21 source.t19 0.9905
R110 source.n21 source.t21 0.9905
R111 source.n19 source.t24 0.9905
R112 source.n19 source.t25 0.9905
R113 source.n17 source.t30 0.9905
R114 source.n17 source.t17 0.9905
R115 source.n1 source.t20 0.9905
R116 source.n1 source.t27 0.9905
R117 source.n3 source.t31 0.9905
R118 source.n3 source.t26 0.9905
R119 source.n5 source.t22 0.9905
R120 source.n5 source.t23 0.9905
R121 source.n9 source.t6 0.9905
R122 source.n9 source.t11 0.9905
R123 source.n11 source.t13 0.9905
R124 source.n11 source.t12 0.9905
R125 source.n13 source.t15 0.9905
R126 source.n13 source.t3 0.9905
R127 source.n15 source.n14 0.974638
R128 source.n14 source.n12 0.974638
R129 source.n12 source.n10 0.974638
R130 source.n10 source.n8 0.974638
R131 source.n7 source.n6 0.974638
R132 source.n6 source.n4 0.974638
R133 source.n4 source.n2 0.974638
R134 source.n2 source.n0 0.974638
R135 source.n18 source.n16 0.974638
R136 source.n20 source.n18 0.974638
R137 source.n22 source.n20 0.974638
R138 source.n23 source.n22 0.974638
R139 source.n26 source.n24 0.974638
R140 source.n28 source.n26 0.974638
R141 source.n30 source.n28 0.974638
R142 source.n31 source.n30 0.974638
R143 source.n8 source.n7 0.470328
R144 source.n24 source.n23 0.470328
R145 source source.n32 0.188
R146 drain_left.n9 drain_left.n7 60.7926
R147 drain_left.n5 drain_left.n3 60.7925
R148 drain_left.n2 drain_left.n0 60.7925
R149 drain_left.n13 drain_left.n12 59.8185
R150 drain_left.n11 drain_left.n10 59.8185
R151 drain_left.n9 drain_left.n8 59.8185
R152 drain_left.n5 drain_left.n4 59.8184
R153 drain_left.n2 drain_left.n1 59.8184
R154 drain_left drain_left.n6 39.7596
R155 drain_left drain_left.n13 6.62735
R156 drain_left.n3 drain_left.t11 0.9905
R157 drain_left.n3 drain_left.t15 0.9905
R158 drain_left.n4 drain_left.t12 0.9905
R159 drain_left.n4 drain_left.t3 0.9905
R160 drain_left.n1 drain_left.t14 0.9905
R161 drain_left.n1 drain_left.t4 0.9905
R162 drain_left.n0 drain_left.t13 0.9905
R163 drain_left.n0 drain_left.t10 0.9905
R164 drain_left.n12 drain_left.t8 0.9905
R165 drain_left.n12 drain_left.t9 0.9905
R166 drain_left.n10 drain_left.t2 0.9905
R167 drain_left.n10 drain_left.t7 0.9905
R168 drain_left.n8 drain_left.t5 0.9905
R169 drain_left.n8 drain_left.t6 0.9905
R170 drain_left.n7 drain_left.t0 0.9905
R171 drain_left.n7 drain_left.t1 0.9905
R172 drain_left.n11 drain_left.n9 0.974638
R173 drain_left.n13 drain_left.n11 0.974638
R174 drain_left.n6 drain_left.n5 0.432223
R175 drain_left.n6 drain_left.n2 0.432223
R176 minus.n5 minus.t8 672.628
R177 minus.n27 minus.t1 672.628
R178 minus.n6 minus.t6 651.605
R179 minus.n7 minus.t5 651.605
R180 minus.n3 minus.t11 651.605
R181 minus.n13 minus.t12 651.605
R182 minus.n1 minus.t10 651.605
R183 minus.n18 minus.t7 651.605
R184 minus.n20 minus.t13 651.605
R185 minus.n28 minus.t9 651.605
R186 minus.n29 minus.t15 651.605
R187 minus.n25 minus.t4 651.605
R188 minus.n35 minus.t0 651.605
R189 minus.n23 minus.t3 651.605
R190 minus.n40 minus.t14 651.605
R191 minus.n42 minus.t2 651.605
R192 minus.n21 minus.n20 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n15 minus.n14 161.3
R195 minus.n13 minus.n2 161.3
R196 minus.n12 minus.n11 161.3
R197 minus.n10 minus.n3 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n43 minus.n42 161.3
R200 minus.n41 minus.n22 161.3
R201 minus.n37 minus.n36 161.3
R202 minus.n35 minus.n24 161.3
R203 minus.n34 minus.n33 161.3
R204 minus.n32 minus.n25 161.3
R205 minus.n31 minus.n30 161.3
R206 minus.n18 minus.n17 80.6037
R207 minus.n16 minus.n1 80.6037
R208 minus.n7 minus.n4 80.6037
R209 minus.n40 minus.n39 80.6037
R210 minus.n38 minus.n23 80.6037
R211 minus.n29 minus.n26 80.6037
R212 minus.n7 minus.n6 48.2005
R213 minus.n18 minus.n1 48.2005
R214 minus.n29 minus.n28 48.2005
R215 minus.n40 minus.n23 48.2005
R216 minus.n44 minus.n21 45.7543
R217 minus.n8 minus.n7 43.0884
R218 minus.n14 minus.n1 43.0884
R219 minus.n30 minus.n29 43.0884
R220 minus.n36 minus.n23 43.0884
R221 minus.n19 minus.n18 40.1672
R222 minus.n41 minus.n40 40.1672
R223 minus.n5 minus.n4 31.6481
R224 minus.n27 minus.n26 31.6481
R225 minus.n13 minus.n12 24.1005
R226 minus.n12 minus.n3 24.1005
R227 minus.n34 minus.n25 24.1005
R228 minus.n35 minus.n34 24.1005
R229 minus.n6 minus.n5 17.444
R230 minus.n28 minus.n27 17.444
R231 minus.n20 minus.n19 8.03383
R232 minus.n42 minus.n41 8.03383
R233 minus.n44 minus.n43 6.6558
R234 minus.n8 minus.n3 5.11262
R235 minus.n14 minus.n13 5.11262
R236 minus.n30 minus.n25 5.11262
R237 minus.n36 minus.n35 5.11262
R238 minus.n17 minus.n16 0.380177
R239 minus.n39 minus.n38 0.380177
R240 minus.n17 minus.n0 0.285035
R241 minus.n16 minus.n15 0.285035
R242 minus.n9 minus.n4 0.285035
R243 minus.n31 minus.n26 0.285035
R244 minus.n38 minus.n37 0.285035
R245 minus.n39 minus.n22 0.285035
R246 minus.n21 minus.n0 0.189894
R247 minus.n15 minus.n2 0.189894
R248 minus.n11 minus.n2 0.189894
R249 minus.n11 minus.n10 0.189894
R250 minus.n10 minus.n9 0.189894
R251 minus.n32 minus.n31 0.189894
R252 minus.n33 minus.n32 0.189894
R253 minus.n33 minus.n24 0.189894
R254 minus.n37 minus.n24 0.189894
R255 minus.n43 minus.n22 0.189894
R256 minus minus.n44 0.188
R257 drain_right.n9 drain_right.n7 60.7926
R258 drain_right.n5 drain_right.n3 60.7925
R259 drain_right.n2 drain_right.n0 60.7925
R260 drain_right.n9 drain_right.n8 59.8185
R261 drain_right.n11 drain_right.n10 59.8185
R262 drain_right.n13 drain_right.n12 59.8185
R263 drain_right.n5 drain_right.n4 59.8184
R264 drain_right.n2 drain_right.n1 59.8184
R265 drain_right drain_right.n6 39.2063
R266 drain_right drain_right.n13 6.62735
R267 drain_right.n3 drain_right.t1 0.9905
R268 drain_right.n3 drain_right.t13 0.9905
R269 drain_right.n4 drain_right.t15 0.9905
R270 drain_right.n4 drain_right.t12 0.9905
R271 drain_right.n1 drain_right.t0 0.9905
R272 drain_right.n1 drain_right.t11 0.9905
R273 drain_right.n0 drain_right.t14 0.9905
R274 drain_right.n0 drain_right.t6 0.9905
R275 drain_right.n7 drain_right.t9 0.9905
R276 drain_right.n7 drain_right.t7 0.9905
R277 drain_right.n8 drain_right.t4 0.9905
R278 drain_right.n8 drain_right.t10 0.9905
R279 drain_right.n10 drain_right.t5 0.9905
R280 drain_right.n10 drain_right.t3 0.9905
R281 drain_right.n12 drain_right.t2 0.9905
R282 drain_right.n12 drain_right.t8 0.9905
R283 drain_right.n13 drain_right.n11 0.974638
R284 drain_right.n11 drain_right.n9 0.974638
R285 drain_right.n6 drain_right.n5 0.432223
R286 drain_right.n6 drain_right.n2 0.432223
C0 plus drain_right 0.430381f
C1 source drain_left 28.460701f
C2 plus source 17.7243f
C3 plus drain_left 18.1905f
C4 drain_right minus 17.917099f
C5 source minus 17.7102f
C6 minus drain_left 0.173489f
C7 plus minus 8.0575f
C8 source drain_right 28.4635f
C9 drain_right drain_left 1.44945f
C10 drain_right a_n2750_n4888# 8.37026f
C11 drain_left a_n2750_n4888# 8.75568f
C12 source a_n2750_n4888# 13.906367f
C13 minus a_n2750_n4888# 11.554412f
C14 plus a_n2750_n4888# 13.6241f
C15 drain_right.t14 a_n2750_n4888# 0.41955f
C16 drain_right.t6 a_n2750_n4888# 0.41955f
C17 drain_right.n0 a_n2750_n4888# 3.84205f
C18 drain_right.t0 a_n2750_n4888# 0.41955f
C19 drain_right.t11 a_n2750_n4888# 0.41955f
C20 drain_right.n1 a_n2750_n4888# 3.83562f
C21 drain_right.n2 a_n2750_n4888# 0.740612f
C22 drain_right.t1 a_n2750_n4888# 0.41955f
C23 drain_right.t13 a_n2750_n4888# 0.41955f
C24 drain_right.n3 a_n2750_n4888# 3.84205f
C25 drain_right.t15 a_n2750_n4888# 0.41955f
C26 drain_right.t12 a_n2750_n4888# 0.41955f
C27 drain_right.n4 a_n2750_n4888# 3.83562f
C28 drain_right.n5 a_n2750_n4888# 0.740612f
C29 drain_right.n6 a_n2750_n4888# 2.04692f
C30 drain_right.t9 a_n2750_n4888# 0.41955f
C31 drain_right.t7 a_n2750_n4888# 0.41955f
C32 drain_right.n7 a_n2750_n4888# 3.84205f
C33 drain_right.t4 a_n2750_n4888# 0.41955f
C34 drain_right.t10 a_n2750_n4888# 0.41955f
C35 drain_right.n8 a_n2750_n4888# 3.83561f
C36 drain_right.n9 a_n2750_n4888# 0.785594f
C37 drain_right.t5 a_n2750_n4888# 0.41955f
C38 drain_right.t3 a_n2750_n4888# 0.41955f
C39 drain_right.n10 a_n2750_n4888# 3.83561f
C40 drain_right.n11 a_n2750_n4888# 0.390666f
C41 drain_right.t2 a_n2750_n4888# 0.41955f
C42 drain_right.t8 a_n2750_n4888# 0.41955f
C43 drain_right.n12 a_n2750_n4888# 3.83561f
C44 drain_right.n13 a_n2750_n4888# 0.628703f
C45 minus.n0 a_n2750_n4888# 0.050824f
C46 minus.t10 a_n2750_n4888# 1.72579f
C47 minus.n1 a_n2750_n4888# 0.650931f
C48 minus.t7 a_n2750_n4888# 1.72579f
C49 minus.n2 a_n2750_n4888# 0.038088f
C50 minus.t11 a_n2750_n4888# 1.72579f
C51 minus.n3 a_n2750_n4888# 0.640057f
C52 minus.n4 a_n2750_n4888# 0.218454f
C53 minus.t8 a_n2750_n4888# 1.74589f
C54 minus.n5 a_n2750_n4888# 0.626688f
C55 minus.t6 a_n2750_n4888# 1.72579f
C56 minus.n6 a_n2750_n4888# 0.65123f
C57 minus.t5 a_n2750_n4888# 1.72579f
C58 minus.n7 a_n2750_n4888# 0.650931f
C59 minus.n8 a_n2750_n4888# 0.008643f
C60 minus.n9 a_n2750_n4888# 0.050824f
C61 minus.n10 a_n2750_n4888# 0.038088f
C62 minus.n11 a_n2750_n4888# 0.038088f
C63 minus.n12 a_n2750_n4888# 0.008643f
C64 minus.t12 a_n2750_n4888# 1.72579f
C65 minus.n13 a_n2750_n4888# 0.640057f
C66 minus.n14 a_n2750_n4888# 0.008643f
C67 minus.n15 a_n2750_n4888# 0.050824f
C68 minus.n16 a_n2750_n4888# 0.063441f
C69 minus.n17 a_n2750_n4888# 0.063441f
C70 minus.n18 a_n2750_n4888# 0.650462f
C71 minus.n19 a_n2750_n4888# 0.008643f
C72 minus.t13 a_n2750_n4888# 1.72579f
C73 minus.n20 a_n2750_n4888# 0.636652f
C74 minus.n21 a_n2750_n4888# 1.91331f
C75 minus.n22 a_n2750_n4888# 0.050824f
C76 minus.t3 a_n2750_n4888# 1.72579f
C77 minus.n23 a_n2750_n4888# 0.650931f
C78 minus.n24 a_n2750_n4888# 0.038088f
C79 minus.t4 a_n2750_n4888# 1.72579f
C80 minus.n25 a_n2750_n4888# 0.640057f
C81 minus.n26 a_n2750_n4888# 0.218454f
C82 minus.t1 a_n2750_n4888# 1.74589f
C83 minus.n27 a_n2750_n4888# 0.626688f
C84 minus.t9 a_n2750_n4888# 1.72579f
C85 minus.n28 a_n2750_n4888# 0.65123f
C86 minus.t15 a_n2750_n4888# 1.72579f
C87 minus.n29 a_n2750_n4888# 0.650931f
C88 minus.n30 a_n2750_n4888# 0.008643f
C89 minus.n31 a_n2750_n4888# 0.050824f
C90 minus.n32 a_n2750_n4888# 0.038088f
C91 minus.n33 a_n2750_n4888# 0.038088f
C92 minus.n34 a_n2750_n4888# 0.008643f
C93 minus.t0 a_n2750_n4888# 1.72579f
C94 minus.n35 a_n2750_n4888# 0.640057f
C95 minus.n36 a_n2750_n4888# 0.008643f
C96 minus.n37 a_n2750_n4888# 0.050824f
C97 minus.n38 a_n2750_n4888# 0.063441f
C98 minus.n39 a_n2750_n4888# 0.063441f
C99 minus.t14 a_n2750_n4888# 1.72579f
C100 minus.n40 a_n2750_n4888# 0.650462f
C101 minus.n41 a_n2750_n4888# 0.008643f
C102 minus.t2 a_n2750_n4888# 1.72579f
C103 minus.n42 a_n2750_n4888# 0.636652f
C104 minus.n43 a_n2750_n4888# 0.26289f
C105 minus.n44 a_n2750_n4888# 2.25871f
C106 drain_left.t13 a_n2750_n4888# 0.42132f
C107 drain_left.t10 a_n2750_n4888# 0.42132f
C108 drain_left.n0 a_n2750_n4888# 3.85826f
C109 drain_left.t14 a_n2750_n4888# 0.42132f
C110 drain_left.t4 a_n2750_n4888# 0.42132f
C111 drain_left.n1 a_n2750_n4888# 3.8518f
C112 drain_left.n2 a_n2750_n4888# 0.743736f
C113 drain_left.t11 a_n2750_n4888# 0.42132f
C114 drain_left.t15 a_n2750_n4888# 0.42132f
C115 drain_left.n3 a_n2750_n4888# 3.85826f
C116 drain_left.t12 a_n2750_n4888# 0.42132f
C117 drain_left.t3 a_n2750_n4888# 0.42132f
C118 drain_left.n4 a_n2750_n4888# 3.8518f
C119 drain_left.n5 a_n2750_n4888# 0.743736f
C120 drain_left.n6 a_n2750_n4888# 2.11035f
C121 drain_left.t0 a_n2750_n4888# 0.42132f
C122 drain_left.t1 a_n2750_n4888# 0.42132f
C123 drain_left.n7 a_n2750_n4888# 3.85825f
C124 drain_left.t5 a_n2750_n4888# 0.42132f
C125 drain_left.t6 a_n2750_n4888# 0.42132f
C126 drain_left.n8 a_n2750_n4888# 3.85179f
C127 drain_left.n9 a_n2750_n4888# 0.788907f
C128 drain_left.t2 a_n2750_n4888# 0.42132f
C129 drain_left.t7 a_n2750_n4888# 0.42132f
C130 drain_left.n10 a_n2750_n4888# 3.85179f
C131 drain_left.n11 a_n2750_n4888# 0.392314f
C132 drain_left.t8 a_n2750_n4888# 0.42132f
C133 drain_left.t9 a_n2750_n4888# 0.42132f
C134 drain_left.n12 a_n2750_n4888# 3.85179f
C135 drain_left.n13 a_n2750_n4888# 0.631355f
C136 source.t28 a_n2750_n4888# 3.98796f
C137 source.n0 a_n2750_n4888# 1.74454f
C138 source.t20 a_n2750_n4888# 0.348953f
C139 source.t27 a_n2750_n4888# 0.348953f
C140 source.n1 a_n2750_n4888# 3.11979f
C141 source.n2 a_n2750_n4888# 0.365331f
C142 source.t31 a_n2750_n4888# 0.348953f
C143 source.t26 a_n2750_n4888# 0.348953f
C144 source.n3 a_n2750_n4888# 3.11979f
C145 source.n4 a_n2750_n4888# 0.365331f
C146 source.t22 a_n2750_n4888# 0.348953f
C147 source.t23 a_n2750_n4888# 0.348953f
C148 source.n5 a_n2750_n4888# 3.11979f
C149 source.n6 a_n2750_n4888# 0.365331f
C150 source.t29 a_n2750_n4888# 3.98797f
C151 source.n7 a_n2750_n4888# 0.412955f
C152 source.t7 a_n2750_n4888# 3.98797f
C153 source.n8 a_n2750_n4888# 0.412955f
C154 source.t6 a_n2750_n4888# 0.348953f
C155 source.t11 a_n2750_n4888# 0.348953f
C156 source.n9 a_n2750_n4888# 3.11979f
C157 source.n10 a_n2750_n4888# 0.365331f
C158 source.t13 a_n2750_n4888# 0.348953f
C159 source.t12 a_n2750_n4888# 0.348953f
C160 source.n11 a_n2750_n4888# 3.11979f
C161 source.n12 a_n2750_n4888# 0.365331f
C162 source.t15 a_n2750_n4888# 0.348953f
C163 source.t3 a_n2750_n4888# 0.348953f
C164 source.n13 a_n2750_n4888# 3.11979f
C165 source.n14 a_n2750_n4888# 0.365331f
C166 source.t8 a_n2750_n4888# 3.98797f
C167 source.n15 a_n2750_n4888# 2.14881f
C168 source.t16 a_n2750_n4888# 3.98795f
C169 source.n16 a_n2750_n4888# 2.14884f
C170 source.t30 a_n2750_n4888# 0.348953f
C171 source.t17 a_n2750_n4888# 0.348953f
C172 source.n17 a_n2750_n4888# 3.11979f
C173 source.n18 a_n2750_n4888# 0.365325f
C174 source.t24 a_n2750_n4888# 0.348953f
C175 source.t25 a_n2750_n4888# 0.348953f
C176 source.n19 a_n2750_n4888# 3.11979f
C177 source.n20 a_n2750_n4888# 0.365325f
C178 source.t19 a_n2750_n4888# 0.348953f
C179 source.t21 a_n2750_n4888# 0.348953f
C180 source.n21 a_n2750_n4888# 3.11979f
C181 source.n22 a_n2750_n4888# 0.365325f
C182 source.t18 a_n2750_n4888# 3.98795f
C183 source.n23 a_n2750_n4888# 0.412977f
C184 source.t1 a_n2750_n4888# 3.98795f
C185 source.n24 a_n2750_n4888# 0.412977f
C186 source.t14 a_n2750_n4888# 0.348953f
C187 source.t4 a_n2750_n4888# 0.348953f
C188 source.n25 a_n2750_n4888# 3.11979f
C189 source.n26 a_n2750_n4888# 0.365325f
C190 source.t10 a_n2750_n4888# 0.348953f
C191 source.t0 a_n2750_n4888# 0.348953f
C192 source.n27 a_n2750_n4888# 3.11979f
C193 source.n28 a_n2750_n4888# 0.365325f
C194 source.t9 a_n2750_n4888# 0.348953f
C195 source.t2 a_n2750_n4888# 0.348953f
C196 source.n29 a_n2750_n4888# 3.11979f
C197 source.n30 a_n2750_n4888# 0.365325f
C198 source.t5 a_n2750_n4888# 3.98795f
C199 source.n31 a_n2750_n4888# 0.561781f
C200 source.n32 a_n2750_n4888# 2.00705f
C201 plus.n0 a_n2750_n4888# 0.051263f
C202 plus.t6 a_n2750_n4888# 1.7407f
C203 plus.t7 a_n2750_n4888# 1.7407f
C204 plus.n1 a_n2750_n4888# 0.063989f
C205 plus.t8 a_n2750_n4888# 1.7407f
C206 plus.n2 a_n2750_n4888# 0.063989f
C207 plus.t13 a_n2750_n4888# 1.7407f
C208 plus.n3 a_n2750_n4888# 0.645589f
C209 plus.n4 a_n2750_n4888# 0.038417f
C210 plus.t9 a_n2750_n4888# 1.7407f
C211 plus.t10 a_n2750_n4888# 1.7407f
C212 plus.n5 a_n2750_n4888# 0.656557f
C213 plus.t14 a_n2750_n4888# 1.7407f
C214 plus.n6 a_n2750_n4888# 0.656858f
C215 plus.t15 a_n2750_n4888# 1.76098f
C216 plus.n7 a_n2750_n4888# 0.632105f
C217 plus.n8 a_n2750_n4888# 0.220342f
C218 plus.n9 a_n2750_n4888# 0.051263f
C219 plus.n10 a_n2750_n4888# 0.008718f
C220 plus.n11 a_n2750_n4888# 0.645589f
C221 plus.n12 a_n2750_n4888# 0.008718f
C222 plus.n13 a_n2750_n4888# 0.038417f
C223 plus.n14 a_n2750_n4888# 0.038417f
C224 plus.n15 a_n2750_n4888# 0.051263f
C225 plus.n16 a_n2750_n4888# 0.008718f
C226 plus.n17 a_n2750_n4888# 0.656557f
C227 plus.n18 a_n2750_n4888# 0.656083f
C228 plus.n19 a_n2750_n4888# 0.008718f
C229 plus.n20 a_n2750_n4888# 0.642155f
C230 plus.n21 a_n2750_n4888# 0.597068f
C231 plus.n22 a_n2750_n4888# 0.051263f
C232 plus.t2 a_n2750_n4888# 1.7407f
C233 plus.n23 a_n2750_n4888# 0.063989f
C234 plus.t5 a_n2750_n4888# 1.7407f
C235 plus.n24 a_n2750_n4888# 0.063989f
C236 plus.t1 a_n2750_n4888# 1.7407f
C237 plus.t11 a_n2750_n4888# 1.7407f
C238 plus.n25 a_n2750_n4888# 0.645589f
C239 plus.n26 a_n2750_n4888# 0.038417f
C240 plus.t3 a_n2750_n4888# 1.7407f
C241 plus.t12 a_n2750_n4888# 1.7407f
C242 plus.n27 a_n2750_n4888# 0.656557f
C243 plus.t4 a_n2750_n4888# 1.7407f
C244 plus.n28 a_n2750_n4888# 0.656858f
C245 plus.t0 a_n2750_n4888# 1.76098f
C246 plus.n29 a_n2750_n4888# 0.632105f
C247 plus.n30 a_n2750_n4888# 0.220342f
C248 plus.n31 a_n2750_n4888# 0.051263f
C249 plus.n32 a_n2750_n4888# 0.008718f
C250 plus.n33 a_n2750_n4888# 0.645589f
C251 plus.n34 a_n2750_n4888# 0.008718f
C252 plus.n35 a_n2750_n4888# 0.038417f
C253 plus.n36 a_n2750_n4888# 0.038417f
C254 plus.n37 a_n2750_n4888# 0.051263f
C255 plus.n38 a_n2750_n4888# 0.008718f
C256 plus.n39 a_n2750_n4888# 0.656557f
C257 plus.n40 a_n2750_n4888# 0.656083f
C258 plus.n41 a_n2750_n4888# 0.008718f
C259 plus.n42 a_n2750_n4888# 0.642155f
C260 plus.n43 a_n2750_n4888# 1.5496f
.ends

