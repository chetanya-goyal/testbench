* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t4 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 source.t26 plus.t1 drain_left.t1 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X2 drain_right.t13 minus.t0 source.t6 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 source.t5 minus.t1 drain_right.t12 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X4 source.t13 minus.t2 drain_right.t11 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X5 drain_right.t10 minus.t3 source.t3 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X6 a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X7 drain_right.t9 minus.t4 source.t2 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X8 drain_left.t9 plus.t2 source.t25 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X9 drain_right.t8 minus.t5 source.t7 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X10 source.t1 minus.t6 drain_right.t7 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X11 source.t4 minus.t7 drain_right.t6 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X12 source.t24 plus.t3 drain_left.t5 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X13 drain_left.t6 plus.t4 source.t23 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X14 drain_left.t11 plus.t5 source.t22 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X15 drain_left.t10 plus.t6 source.t21 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X16 drain_left.t7 plus.t7 source.t20 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X17 drain_left.t13 plus.t8 source.t19 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X18 drain_right.t5 minus.t8 source.t10 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X19 drain_left.t8 plus.t9 source.t18 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X20 drain_right.t4 minus.t9 source.t11 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X21 drain_left.t12 plus.t10 source.t17 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X22 a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X23 a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X24 source.t16 plus.t11 drain_left.t3 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X25 source.t15 plus.t12 drain_left.t2 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X26 drain_right.t3 minus.t10 source.t12 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X27 drain_right.t2 minus.t11 source.t0 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X28 source.t8 minus.t12 drain_right.t1 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X29 source.t14 plus.t13 drain_left.t0 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X30 a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X31 source.t9 minus.t13 drain_right.t0 a_n1644_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
R0 plus.n3 plus.t2 256.776
R1 plus.n15 plus.t4 256.776
R2 plus.n20 plus.t8 256.776
R3 plus.n32 plus.t9 256.776
R4 plus.n1 plus.t0 221.72
R5 plus.n4 plus.t1 221.72
R6 plus.n6 plus.t6 221.72
R7 plus.n12 plus.t5 221.72
R8 plus.n14 plus.t13 221.72
R9 plus.n18 plus.t12 221.72
R10 plus.n21 plus.t3 221.72
R11 plus.n23 plus.t10 221.72
R12 plus.n29 plus.t7 221.72
R13 plus.n31 plus.t11 221.72
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 25.0142
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus.n7 plus.n6 11.6853
R46 plus.n12 plus.n11 11.6853
R47 plus.n29 plus.n28 11.6853
R48 plus.n24 plus.n23 11.6853
R49 plus plus.n16 7.92853
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t9 260.433
R61 drain_left.n1 drain_left.t8 260.432
R62 drain_left.n4 drain_left.n2 240.631
R63 drain_left.n11 drain_left.n10 240.132
R64 drain_left.n9 drain_left.n8 240.132
R65 drain_left.n7 drain_left.n6 240.132
R66 drain_left.n4 drain_left.n3 240.131
R67 drain_left.n1 drain_left.n0 240.131
R68 drain_left drain_left.n5 21.9087
R69 drain_left.n2 drain_left.t5 19.8005
R70 drain_left.n2 drain_left.t13 19.8005
R71 drain_left.n3 drain_left.t2 19.8005
R72 drain_left.n3 drain_left.t12 19.8005
R73 drain_left.n0 drain_left.t3 19.8005
R74 drain_left.n0 drain_left.t7 19.8005
R75 drain_left.n10 drain_left.t0 19.8005
R76 drain_left.n10 drain_left.t6 19.8005
R77 drain_left.n8 drain_left.t4 19.8005
R78 drain_left.n8 drain_left.t11 19.8005
R79 drain_left.n6 drain_left.t1 19.8005
R80 drain_left.n6 drain_left.t10 19.8005
R81 drain_left drain_left.n11 6.15322
R82 drain_left.n9 drain_left.n7 0.5005
R83 drain_left.n11 drain_left.n9 0.5005
R84 drain_left.n5 drain_left.n1 0.320154
R85 drain_left.n5 drain_left.n4 0.070154
R86 source.n0 source.t23 243.255
R87 source.n7 source.t11 243.255
R88 source.n27 source.t7 243.254
R89 source.n20 source.t19 243.254
R90 source.n2 source.n1 223.454
R91 source.n4 source.n3 223.454
R92 source.n6 source.n5 223.454
R93 source.n9 source.n8 223.454
R94 source.n11 source.n10 223.454
R95 source.n13 source.n12 223.454
R96 source.n26 source.n25 223.453
R97 source.n24 source.n23 223.453
R98 source.n22 source.n21 223.453
R99 source.n19 source.n18 223.453
R100 source.n17 source.n16 223.453
R101 source.n15 source.n14 223.453
R102 source.n25 source.t3 19.8005
R103 source.n25 source.t4 19.8005
R104 source.n23 source.t6 19.8005
R105 source.n23 source.t9 19.8005
R106 source.n21 source.t2 19.8005
R107 source.n21 source.t8 19.8005
R108 source.n18 source.t17 19.8005
R109 source.n18 source.t24 19.8005
R110 source.n16 source.t20 19.8005
R111 source.n16 source.t15 19.8005
R112 source.n14 source.t18 19.8005
R113 source.n14 source.t16 19.8005
R114 source.n1 source.t22 19.8005
R115 source.n1 source.t14 19.8005
R116 source.n3 source.t21 19.8005
R117 source.n3 source.t27 19.8005
R118 source.n5 source.t25 19.8005
R119 source.n5 source.t26 19.8005
R120 source.n8 source.t10 19.8005
R121 source.n8 source.t13 19.8005
R122 source.n10 source.t12 19.8005
R123 source.n10 source.t5 19.8005
R124 source.n12 source.t0 19.8005
R125 source.n12 source.t1 19.8005
R126 source.n15 source.n13 13.9544
R127 source.n28 source.n0 7.94146
R128 source.n28 source.n27 5.51343
R129 source.n7 source.n6 0.720328
R130 source.n22 source.n20 0.720328
R131 source.n13 source.n11 0.5005
R132 source.n11 source.n9 0.5005
R133 source.n9 source.n7 0.5005
R134 source.n6 source.n4 0.5005
R135 source.n4 source.n2 0.5005
R136 source.n2 source.n0 0.5005
R137 source.n17 source.n15 0.5005
R138 source.n19 source.n17 0.5005
R139 source.n20 source.n19 0.5005
R140 source.n24 source.n22 0.5005
R141 source.n26 source.n24 0.5005
R142 source.n27 source.n26 0.5005
R143 source source.n28 0.188
R144 minus.n15 minus.t11 256.776
R145 minus.n3 minus.t9 256.776
R146 minus.n32 minus.t5 256.776
R147 minus.n20 minus.t4 256.776
R148 minus.n1 minus.t1 221.72
R149 minus.n14 minus.t6 221.72
R150 minus.n12 minus.t10 221.72
R151 minus.n6 minus.t8 221.72
R152 minus.n4 minus.t2 221.72
R153 minus.n18 minus.t13 221.72
R154 minus.n31 minus.t7 221.72
R155 minus.n29 minus.t3 221.72
R156 minus.n23 minus.t0 221.72
R157 minus.n21 minus.t12 221.72
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 61.346
R177 minus.n6 minus.n5 61.346
R178 minus.n23 minus.n22 61.346
R179 minus.n30 minus.n29 61.346
R180 minus.n15 minus.n14 49.6611
R181 minus.n4 minus.n3 49.6611
R182 minus.n21 minus.n20 49.6611
R183 minus.n32 minus.n31 49.6611
R184 minus.n34 minus.n16 26.9664
R185 minus.n14 minus.n13 23.3702
R186 minus.n5 minus.n4 23.3702
R187 minus.n22 minus.n21 23.3702
R188 minus.n31 minus.n30 23.3702
R189 minus.n12 minus.n11 11.6853
R190 minus.n7 minus.n6 11.6853
R191 minus.n24 minus.n23 11.6853
R192 minus.n29 minus.n28 11.6853
R193 minus.n34 minus.n33 6.45126
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t9 260.432
R206 drain_right.n11 drain_right.t2 259.933
R207 drain_right.n8 drain_right.n6 240.632
R208 drain_right.n4 drain_right.n2 240.631
R209 drain_right.n8 drain_right.n7 240.132
R210 drain_right.n10 drain_right.n9 240.132
R211 drain_right.n4 drain_right.n3 240.131
R212 drain_right.n1 drain_right.n0 240.131
R213 drain_right drain_right.n5 21.3555
R214 drain_right.n2 drain_right.t6 19.8005
R215 drain_right.n2 drain_right.t8 19.8005
R216 drain_right.n3 drain_right.t0 19.8005
R217 drain_right.n3 drain_right.t10 19.8005
R218 drain_right.n0 drain_right.t1 19.8005
R219 drain_right.n0 drain_right.t13 19.8005
R220 drain_right.n6 drain_right.t11 19.8005
R221 drain_right.n6 drain_right.t4 19.8005
R222 drain_right.n7 drain_right.t12 19.8005
R223 drain_right.n7 drain_right.t5 19.8005
R224 drain_right.n9 drain_right.t7 19.8005
R225 drain_right.n9 drain_right.t3 19.8005
R226 drain_right drain_right.n11 5.90322
R227 drain_right.n11 drain_right.n10 0.5005
R228 drain_right.n10 drain_right.n8 0.5005
R229 drain_right.n5 drain_right.n1 0.320154
R230 drain_right.n5 drain_right.n4 0.070154
C0 drain_right source 4.9062f
C1 minus drain_left 0.179388f
C2 plus drain_left 0.967045f
C3 minus source 1.04276f
C4 plus source 1.05668f
C5 source drain_left 4.90817f
C6 drain_right minus 0.809026f
C7 drain_right plus 0.321841f
C8 plus minus 3.17867f
C9 drain_right drain_left 0.83657f
C10 drain_right a_n1644_n1088# 3.55559f
C11 drain_left a_n1644_n1088# 3.7877f
C12 source a_n1644_n1088# 2.128015f
C13 minus a_n1644_n1088# 5.49307f
C14 plus a_n1644_n1088# 6.183045f
C15 drain_right.t9 a_n1644_n1088# 0.123703f
C16 drain_right.t1 a_n1644_n1088# 0.019926f
C17 drain_right.t13 a_n1644_n1088# 0.019926f
C18 drain_right.n0 a_n1644_n1088# 0.077427f
C19 drain_right.n1 a_n1644_n1088# 0.479944f
C20 drain_right.t6 a_n1644_n1088# 0.019926f
C21 drain_right.t8 a_n1644_n1088# 0.019926f
C22 drain_right.n2 a_n1644_n1088# 0.077983f
C23 drain_right.t0 a_n1644_n1088# 0.019926f
C24 drain_right.t10 a_n1644_n1088# 0.019926f
C25 drain_right.n3 a_n1644_n1088# 0.077427f
C26 drain_right.n4 a_n1644_n1088# 0.498196f
C27 drain_right.n5 a_n1644_n1088# 0.572725f
C28 drain_right.t11 a_n1644_n1088# 0.019926f
C29 drain_right.t4 a_n1644_n1088# 0.019926f
C30 drain_right.n6 a_n1644_n1088# 0.077983f
C31 drain_right.t12 a_n1644_n1088# 0.019926f
C32 drain_right.t5 a_n1644_n1088# 0.019926f
C33 drain_right.n7 a_n1644_n1088# 0.077427f
C34 drain_right.n8 a_n1644_n1088# 0.524769f
C35 drain_right.t7 a_n1644_n1088# 0.019926f
C36 drain_right.t3 a_n1644_n1088# 0.019926f
C37 drain_right.n9 a_n1644_n1088# 0.077427f
C38 drain_right.n10 a_n1644_n1088# 0.257585f
C39 drain_right.t2 a_n1644_n1088# 0.123251f
C40 drain_right.n11 a_n1644_n1088# 0.443292f
C41 minus.n0 a_n1644_n1088# 0.033547f
C42 minus.t11 a_n1644_n1088# 0.029698f
C43 minus.t6 a_n1644_n1088# 0.025854f
C44 minus.t10 a_n1644_n1088# 0.025854f
C45 minus.t1 a_n1644_n1088# 0.025854f
C46 minus.n1 a_n1644_n1088# 0.03949f
C47 minus.n2 a_n1644_n1088# 0.071807f
C48 minus.t8 a_n1644_n1088# 0.025854f
C49 minus.t2 a_n1644_n1088# 0.025854f
C50 minus.t9 a_n1644_n1088# 0.029698f
C51 minus.n3 a_n1644_n1088# 0.037139f
C52 minus.n4 a_n1644_n1088# 0.028361f
C53 minus.n5 a_n1644_n1088# 0.012783f
C54 minus.n6 a_n1644_n1088# 0.028361f
C55 minus.n7 a_n1644_n1088# 0.012783f
C56 minus.n8 a_n1644_n1088# 0.033547f
C57 minus.n9 a_n1644_n1088# 0.033547f
C58 minus.n10 a_n1644_n1088# 0.033547f
C59 minus.n11 a_n1644_n1088# 0.012783f
C60 minus.n12 a_n1644_n1088# 0.028361f
C61 minus.n13 a_n1644_n1088# 0.012783f
C62 minus.n14 a_n1644_n1088# 0.028361f
C63 minus.n15 a_n1644_n1088# 0.037094f
C64 minus.n16 a_n1644_n1088# 0.722005f
C65 minus.n17 a_n1644_n1088# 0.033547f
C66 minus.t7 a_n1644_n1088# 0.025854f
C67 minus.t3 a_n1644_n1088# 0.025854f
C68 minus.t13 a_n1644_n1088# 0.025854f
C69 minus.n18 a_n1644_n1088# 0.03949f
C70 minus.n19 a_n1644_n1088# 0.071807f
C71 minus.t0 a_n1644_n1088# 0.025854f
C72 minus.t12 a_n1644_n1088# 0.025854f
C73 minus.t4 a_n1644_n1088# 0.029698f
C74 minus.n20 a_n1644_n1088# 0.037139f
C75 minus.n21 a_n1644_n1088# 0.028361f
C76 minus.n22 a_n1644_n1088# 0.012783f
C77 minus.n23 a_n1644_n1088# 0.028361f
C78 minus.n24 a_n1644_n1088# 0.012783f
C79 minus.n25 a_n1644_n1088# 0.033547f
C80 minus.n26 a_n1644_n1088# 0.033547f
C81 minus.n27 a_n1644_n1088# 0.033547f
C82 minus.n28 a_n1644_n1088# 0.012783f
C83 minus.n29 a_n1644_n1088# 0.028361f
C84 minus.n30 a_n1644_n1088# 0.012783f
C85 minus.n31 a_n1644_n1088# 0.028361f
C86 minus.t5 a_n1644_n1088# 0.029698f
C87 minus.n32 a_n1644_n1088# 0.037094f
C88 minus.n33 a_n1644_n1088# 0.215461f
C89 minus.n34 a_n1644_n1088# 0.894581f
C90 source.t23 a_n1644_n1088# 0.146305f
C91 source.n0 a_n1644_n1088# 0.619928f
C92 source.t22 a_n1644_n1088# 0.026286f
C93 source.t14 a_n1644_n1088# 0.026286f
C94 source.n1 a_n1644_n1088# 0.08525f
C95 source.n2 a_n1644_n1088# 0.31148f
C96 source.t21 a_n1644_n1088# 0.026286f
C97 source.t27 a_n1644_n1088# 0.026286f
C98 source.n3 a_n1644_n1088# 0.08525f
C99 source.n4 a_n1644_n1088# 0.31148f
C100 source.t25 a_n1644_n1088# 0.026286f
C101 source.t26 a_n1644_n1088# 0.026286f
C102 source.n5 a_n1644_n1088# 0.08525f
C103 source.n6 a_n1644_n1088# 0.335042f
C104 source.t11 a_n1644_n1088# 0.146305f
C105 source.n7 a_n1644_n1088# 0.345677f
C106 source.t10 a_n1644_n1088# 0.026286f
C107 source.t13 a_n1644_n1088# 0.026286f
C108 source.n8 a_n1644_n1088# 0.08525f
C109 source.n9 a_n1644_n1088# 0.31148f
C110 source.t12 a_n1644_n1088# 0.026286f
C111 source.t5 a_n1644_n1088# 0.026286f
C112 source.n10 a_n1644_n1088# 0.08525f
C113 source.n11 a_n1644_n1088# 0.31148f
C114 source.t0 a_n1644_n1088# 0.026286f
C115 source.t1 a_n1644_n1088# 0.026286f
C116 source.n12 a_n1644_n1088# 0.08525f
C117 source.n13 a_n1644_n1088# 0.928472f
C118 source.t18 a_n1644_n1088# 0.026286f
C119 source.t16 a_n1644_n1088# 0.026286f
C120 source.n14 a_n1644_n1088# 0.08525f
C121 source.n15 a_n1644_n1088# 0.928473f
C122 source.t20 a_n1644_n1088# 0.026286f
C123 source.t15 a_n1644_n1088# 0.026286f
C124 source.n16 a_n1644_n1088# 0.08525f
C125 source.n17 a_n1644_n1088# 0.31148f
C126 source.t17 a_n1644_n1088# 0.026286f
C127 source.t24 a_n1644_n1088# 0.026286f
C128 source.n18 a_n1644_n1088# 0.08525f
C129 source.n19 a_n1644_n1088# 0.31148f
C130 source.t19 a_n1644_n1088# 0.146305f
C131 source.n20 a_n1644_n1088# 0.345677f
C132 source.t2 a_n1644_n1088# 0.026286f
C133 source.t8 a_n1644_n1088# 0.026286f
C134 source.n21 a_n1644_n1088# 0.08525f
C135 source.n22 a_n1644_n1088# 0.335042f
C136 source.t6 a_n1644_n1088# 0.026286f
C137 source.t9 a_n1644_n1088# 0.026286f
C138 source.n23 a_n1644_n1088# 0.08525f
C139 source.n24 a_n1644_n1088# 0.31148f
C140 source.t3 a_n1644_n1088# 0.026286f
C141 source.t4 a_n1644_n1088# 0.026286f
C142 source.n25 a_n1644_n1088# 0.08525f
C143 source.n26 a_n1644_n1088# 0.31148f
C144 source.t7 a_n1644_n1088# 0.146305f
C145 source.n27 a_n1644_n1088# 0.502957f
C146 source.n28 a_n1644_n1088# 0.671805f
C147 drain_left.t8 a_n1644_n1088# 0.121262f
C148 drain_left.t3 a_n1644_n1088# 0.019533f
C149 drain_left.t7 a_n1644_n1088# 0.019533f
C150 drain_left.n0 a_n1644_n1088# 0.075899f
C151 drain_left.n1 a_n1644_n1088# 0.470473f
C152 drain_left.t5 a_n1644_n1088# 0.019533f
C153 drain_left.t13 a_n1644_n1088# 0.019533f
C154 drain_left.n2 a_n1644_n1088# 0.076444f
C155 drain_left.t2 a_n1644_n1088# 0.019533f
C156 drain_left.t12 a_n1644_n1088# 0.019533f
C157 drain_left.n3 a_n1644_n1088# 0.075899f
C158 drain_left.n4 a_n1644_n1088# 0.488365f
C159 drain_left.n5 a_n1644_n1088# 0.60926f
C160 drain_left.t9 a_n1644_n1088# 0.121262f
C161 drain_left.t1 a_n1644_n1088# 0.019533f
C162 drain_left.t10 a_n1644_n1088# 0.019533f
C163 drain_left.n6 a_n1644_n1088# 0.075899f
C164 drain_left.n7 a_n1644_n1088# 0.483044f
C165 drain_left.t4 a_n1644_n1088# 0.019533f
C166 drain_left.t11 a_n1644_n1088# 0.019533f
C167 drain_left.n8 a_n1644_n1088# 0.075899f
C168 drain_left.n9 a_n1644_n1088# 0.252502f
C169 drain_left.t0 a_n1644_n1088# 0.019533f
C170 drain_left.t6 a_n1644_n1088# 0.019533f
C171 drain_left.n10 a_n1644_n1088# 0.075899f
C172 drain_left.n11 a_n1644_n1088# 0.456531f
C173 plus.n0 a_n1644_n1088# 0.034274f
C174 plus.t13 a_n1644_n1088# 0.026414f
C175 plus.t5 a_n1644_n1088# 0.026414f
C176 plus.t0 a_n1644_n1088# 0.026414f
C177 plus.n1 a_n1644_n1088# 0.040345f
C178 plus.n2 a_n1644_n1088# 0.073362f
C179 plus.t6 a_n1644_n1088# 0.026414f
C180 plus.t1 a_n1644_n1088# 0.026414f
C181 plus.t2 a_n1644_n1088# 0.030341f
C182 plus.n3 a_n1644_n1088# 0.037943f
C183 plus.n4 a_n1644_n1088# 0.028975f
C184 plus.n5 a_n1644_n1088# 0.01306f
C185 plus.n6 a_n1644_n1088# 0.028975f
C186 plus.n7 a_n1644_n1088# 0.01306f
C187 plus.n8 a_n1644_n1088# 0.034274f
C188 plus.n9 a_n1644_n1088# 0.034274f
C189 plus.n10 a_n1644_n1088# 0.034274f
C190 plus.n11 a_n1644_n1088# 0.01306f
C191 plus.n12 a_n1644_n1088# 0.028975f
C192 plus.n13 a_n1644_n1088# 0.01306f
C193 plus.n14 a_n1644_n1088# 0.028975f
C194 plus.t4 a_n1644_n1088# 0.030341f
C195 plus.n15 a_n1644_n1088# 0.037897f
C196 plus.n16 a_n1644_n1088# 0.230824f
C197 plus.n17 a_n1644_n1088# 0.034274f
C198 plus.t9 a_n1644_n1088# 0.030341f
C199 plus.t11 a_n1644_n1088# 0.026414f
C200 plus.t7 a_n1644_n1088# 0.026414f
C201 plus.t12 a_n1644_n1088# 0.026414f
C202 plus.n18 a_n1644_n1088# 0.040345f
C203 plus.n19 a_n1644_n1088# 0.073362f
C204 plus.t10 a_n1644_n1088# 0.026414f
C205 plus.t3 a_n1644_n1088# 0.026414f
C206 plus.t8 a_n1644_n1088# 0.030341f
C207 plus.n20 a_n1644_n1088# 0.037943f
C208 plus.n21 a_n1644_n1088# 0.028975f
C209 plus.n22 a_n1644_n1088# 0.01306f
C210 plus.n23 a_n1644_n1088# 0.028975f
C211 plus.n24 a_n1644_n1088# 0.01306f
C212 plus.n25 a_n1644_n1088# 0.034274f
C213 plus.n26 a_n1644_n1088# 0.034274f
C214 plus.n27 a_n1644_n1088# 0.034274f
C215 plus.n28 a_n1644_n1088# 0.01306f
C216 plus.n29 a_n1644_n1088# 0.028975f
C217 plus.n30 a_n1644_n1088# 0.01306f
C218 plus.n31 a_n1644_n1088# 0.028975f
C219 plus.n32 a_n1644_n1088# 0.037897f
C220 plus.n33 a_n1644_n1088# 0.717125f
.ends

