* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t11 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X1 a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X2 a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X3 source.t8 minus.t0 drain_right.t9 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_left.t8 plus.t1 source.t19 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X5 drain_right.t8 minus.t1 source.t4 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X6 drain_right.t7 minus.t2 source.t1 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 drain_right.t6 minus.t3 source.t3 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 source.t14 plus.t2 drain_left.t7 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 drain_left.t6 plus.t3 source.t18 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 drain_right.t5 minus.t4 source.t5 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X11 source.t6 minus.t5 drain_right.t4 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X13 drain_left.t5 plus.t4 source.t15 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X14 drain_right.t3 minus.t6 source.t7 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X15 source.t0 minus.t7 drain_right.t2 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 source.t10 plus.t5 drain_left.t4 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 source.t13 plus.t6 drain_left.t3 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 source.t9 minus.t8 drain_right.t1 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X20 source.t12 plus.t7 drain_left.t2 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X21 drain_left.t1 plus.t8 source.t16 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X22 drain_left.t0 plus.t9 source.t17 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 drain_right.t0 minus.t9 source.t2 a_n1712_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
R0 plus.n5 plus.n4 161.3
R1 plus.n6 plus.n1 161.3
R2 plus.n8 plus.n7 161.3
R3 plus.n9 plus.n0 161.3
R4 plus.n11 plus.n10 161.3
R5 plus.n17 plus.n16 161.3
R6 plus.n18 plus.n13 161.3
R7 plus.n20 plus.n19 161.3
R8 plus.n21 plus.n12 161.3
R9 plus.n23 plus.n22 161.3
R10 plus.n2 plus.t1 147.749
R11 plus.n14 plus.t4 147.749
R12 plus.n10 plus.t8 126.766
R13 plus.n9 plus.t2 126.766
R14 plus.n1 plus.t9 126.766
R15 plus.n3 plus.t5 126.766
R16 plus.n22 plus.t0 126.766
R17 plus.n21 plus.t7 126.766
R18 plus.n13 plus.t3 126.766
R19 plus.n15 plus.t6 126.766
R20 plus.n5 plus.n2 70.4033
R21 plus.n17 plus.n14 70.4033
R22 plus.n10 plus.n9 48.2005
R23 plus.n22 plus.n21 48.2005
R24 plus.n8 plus.n1 36.5157
R25 plus.n4 plus.n1 36.5157
R26 plus.n20 plus.n13 36.5157
R27 plus.n16 plus.n13 36.5157
R28 plus plus.n23 25.3835
R29 plus.n3 plus.n2 20.9576
R30 plus.n15 plus.n14 20.9576
R31 plus.n9 plus.n8 11.6853
R32 plus.n4 plus.n3 11.6853
R33 plus.n21 plus.n20 11.6853
R34 plus.n16 plus.n15 11.6853
R35 plus plus.n11 8.04027
R36 plus.n6 plus.n5 0.189894
R37 plus.n7 plus.n6 0.189894
R38 plus.n7 plus.n0 0.189894
R39 plus.n11 plus.n0 0.189894
R40 plus.n23 plus.n12 0.189894
R41 plus.n19 plus.n12 0.189894
R42 plus.n19 plus.n18 0.189894
R43 plus.n18 plus.n17 0.189894
R44 source.n0 source.t16 243.255
R45 source.n5 source.t7 243.255
R46 source.n19 source.t2 243.254
R47 source.n14 source.t15 243.254
R48 source.n2 source.n1 223.454
R49 source.n4 source.n3 223.454
R50 source.n7 source.n6 223.454
R51 source.n9 source.n8 223.454
R52 source.n18 source.n17 223.453
R53 source.n16 source.n15 223.453
R54 source.n13 source.n12 223.453
R55 source.n11 source.n10 223.453
R56 source.n17 source.t3 19.8005
R57 source.n17 source.t6 19.8005
R58 source.n15 source.t5 19.8005
R59 source.n15 source.t0 19.8005
R60 source.n12 source.t18 19.8005
R61 source.n12 source.t13 19.8005
R62 source.n10 source.t11 19.8005
R63 source.n10 source.t12 19.8005
R64 source.n1 source.t17 19.8005
R65 source.n1 source.t14 19.8005
R66 source.n3 source.t19 19.8005
R67 source.n3 source.t10 19.8005
R68 source.n6 source.t1 19.8005
R69 source.n6 source.t8 19.8005
R70 source.n8 source.t4 19.8005
R71 source.n8 source.t9 19.8005
R72 source.n11 source.n9 14.3854
R73 source.n20 source.n0 8.04922
R74 source.n20 source.n19 5.62119
R75 source.n5 source.n4 0.828086
R76 source.n16 source.n14 0.828086
R77 source.n9 source.n7 0.716017
R78 source.n7 source.n5 0.716017
R79 source.n4 source.n2 0.716017
R80 source.n2 source.n0 0.716017
R81 source.n13 source.n11 0.716017
R82 source.n14 source.n13 0.716017
R83 source.n18 source.n16 0.716017
R84 source.n19 source.n18 0.716017
R85 source source.n20 0.188
R86 drain_left.n5 drain_left.t8 260.649
R87 drain_left.n1 drain_left.t9 260.647
R88 drain_left.n3 drain_left.n2 240.613
R89 drain_left.n7 drain_left.n6 240.132
R90 drain_left.n5 drain_left.n4 240.132
R91 drain_left.n1 drain_left.n0 240.131
R92 drain_left drain_left.n3 22.0747
R93 drain_left.n2 drain_left.t3 19.8005
R94 drain_left.n2 drain_left.t5 19.8005
R95 drain_left.n0 drain_left.t2 19.8005
R96 drain_left.n0 drain_left.t6 19.8005
R97 drain_left.n6 drain_left.t7 19.8005
R98 drain_left.n6 drain_left.t1 19.8005
R99 drain_left.n4 drain_left.t4 19.8005
R100 drain_left.n4 drain_left.t0 19.8005
R101 drain_left drain_left.n7 6.36873
R102 drain_left.n7 drain_left.n5 0.716017
R103 drain_left.n3 drain_left.n1 0.124033
R104 minus.n11 minus.n10 161.3
R105 minus.n9 minus.n0 161.3
R106 minus.n8 minus.n7 161.3
R107 minus.n6 minus.n1 161.3
R108 minus.n5 minus.n4 161.3
R109 minus.n23 minus.n22 161.3
R110 minus.n21 minus.n12 161.3
R111 minus.n20 minus.n19 161.3
R112 minus.n18 minus.n13 161.3
R113 minus.n17 minus.n16 161.3
R114 minus.n2 minus.t6 147.749
R115 minus.n14 minus.t4 147.749
R116 minus.n3 minus.t0 126.766
R117 minus.n1 minus.t2 126.766
R118 minus.n9 minus.t8 126.766
R119 minus.n10 minus.t1 126.766
R120 minus.n15 minus.t7 126.766
R121 minus.n13 minus.t3 126.766
R122 minus.n21 minus.t5 126.766
R123 minus.n22 minus.t9 126.766
R124 minus.n5 minus.n2 70.4033
R125 minus.n17 minus.n14 70.4033
R126 minus.n10 minus.n9 48.2005
R127 minus.n22 minus.n21 48.2005
R128 minus.n4 minus.n1 36.5157
R129 minus.n8 minus.n1 36.5157
R130 minus.n16 minus.n13 36.5157
R131 minus.n20 minus.n13 36.5157
R132 minus.n24 minus.n11 27.3357
R133 minus.n3 minus.n2 20.9576
R134 minus.n15 minus.n14 20.9576
R135 minus.n4 minus.n3 11.6853
R136 minus.n9 minus.n8 11.6853
R137 minus.n16 minus.n15 11.6853
R138 minus.n21 minus.n20 11.6853
R139 minus.n24 minus.n23 6.563
R140 minus.n11 minus.n0 0.189894
R141 minus.n7 minus.n0 0.189894
R142 minus.n7 minus.n6 0.189894
R143 minus.n6 minus.n5 0.189894
R144 minus.n18 minus.n17 0.189894
R145 minus.n19 minus.n18 0.189894
R146 minus.n19 minus.n12 0.189894
R147 minus.n23 minus.n12 0.189894
R148 minus minus.n24 0.188
R149 drain_right.n1 drain_right.t5 260.647
R150 drain_right.n7 drain_right.t8 259.933
R151 drain_right.n6 drain_right.n4 240.849
R152 drain_right.n3 drain_right.n2 240.613
R153 drain_right.n6 drain_right.n5 240.132
R154 drain_right.n1 drain_right.n0 240.131
R155 drain_right drain_right.n3 21.5215
R156 drain_right.n2 drain_right.t4 19.8005
R157 drain_right.n2 drain_right.t0 19.8005
R158 drain_right.n0 drain_right.t2 19.8005
R159 drain_right.n0 drain_right.t6 19.8005
R160 drain_right.n4 drain_right.t9 19.8005
R161 drain_right.n4 drain_right.t3 19.8005
R162 drain_right.n5 drain_right.t1 19.8005
R163 drain_right.n5 drain_right.t7 19.8005
R164 drain_right drain_right.n7 6.01097
R165 drain_right.n7 drain_right.n6 0.716017
R166 drain_right.n3 drain_right.n1 0.124033
C0 drain_right source 3.53729f
C1 plus minus 3.25473f
C2 minus drain_left 0.179645f
C3 plus drain_left 1.00962f
C4 minus source 1.17266f
C5 plus source 1.18657f
C6 drain_left source 3.53814f
C7 drain_right minus 0.844627f
C8 plus drain_right 0.3293f
C9 drain_right drain_left 0.843308f
C10 drain_right a_n1712_n1088# 3.337759f
C11 drain_left a_n1712_n1088# 3.566901f
C12 source a_n1712_n1088# 2.118565f
C13 minus a_n1712_n1088# 5.757642f
C14 plus a_n1712_n1088# 6.410397f
C15 drain_right.t5 a_n1712_n1088# 0.099273f
C16 drain_right.t2 a_n1712_n1088# 0.01596f
C17 drain_right.t6 a_n1712_n1088# 0.01596f
C18 drain_right.n0 a_n1712_n1088# 0.062014f
C19 drain_right.n1 a_n1712_n1088# 0.401825f
C20 drain_right.t4 a_n1712_n1088# 0.01596f
C21 drain_right.t0 a_n1712_n1088# 0.01596f
C22 drain_right.n2 a_n1712_n1088# 0.062471f
C23 drain_right.n3 a_n1712_n1088# 0.713962f
C24 drain_right.t9 a_n1712_n1088# 0.01596f
C25 drain_right.t3 a_n1712_n1088# 0.01596f
C26 drain_right.n4 a_n1712_n1088# 0.062735f
C27 drain_right.t1 a_n1712_n1088# 0.01596f
C28 drain_right.t7 a_n1712_n1088# 0.01596f
C29 drain_right.n5 a_n1712_n1088# 0.062014f
C30 drain_right.n6 a_n1712_n1088# 0.476135f
C31 drain_right.t8 a_n1712_n1088# 0.098717f
C32 drain_right.n7 a_n1712_n1088# 0.379848f
C33 minus.n0 a_n1712_n1088# 0.031388f
C34 minus.t2 a_n1712_n1088# 0.053219f
C35 minus.n1 a_n1712_n1088# 0.058647f
C36 minus.t6 a_n1712_n1088# 0.061087f
C37 minus.n2 a_n1712_n1088# 0.047719f
C38 minus.t0 a_n1712_n1088# 0.053219f
C39 minus.n3 a_n1712_n1088# 0.056905f
C40 minus.n4 a_n1712_n1088# 0.007123f
C41 minus.n5 a_n1712_n1088# 0.100129f
C42 minus.n6 a_n1712_n1088# 0.031388f
C43 minus.n7 a_n1712_n1088# 0.031388f
C44 minus.n8 a_n1712_n1088# 0.007123f
C45 minus.t8 a_n1712_n1088# 0.053219f
C46 minus.n9 a_n1712_n1088# 0.056905f
C47 minus.t1 a_n1712_n1088# 0.053219f
C48 minus.n10 a_n1712_n1088# 0.055357f
C49 minus.n11 a_n1712_n1088# 0.695938f
C50 minus.n12 a_n1712_n1088# 0.031388f
C51 minus.t3 a_n1712_n1088# 0.053219f
C52 minus.n13 a_n1712_n1088# 0.058647f
C53 minus.t4 a_n1712_n1088# 0.061087f
C54 minus.n14 a_n1712_n1088# 0.047719f
C55 minus.t7 a_n1712_n1088# 0.053219f
C56 minus.n15 a_n1712_n1088# 0.056905f
C57 minus.n16 a_n1712_n1088# 0.007123f
C58 minus.n17 a_n1712_n1088# 0.100129f
C59 minus.n18 a_n1712_n1088# 0.031388f
C60 minus.n19 a_n1712_n1088# 0.031388f
C61 minus.n20 a_n1712_n1088# 0.007123f
C62 minus.t5 a_n1712_n1088# 0.053219f
C63 minus.n21 a_n1712_n1088# 0.056905f
C64 minus.t9 a_n1712_n1088# 0.053219f
C65 minus.n22 a_n1712_n1088# 0.055357f
C66 minus.n23 a_n1712_n1088# 0.209855f
C67 minus.n24 a_n1712_n1088# 0.857524f
C68 drain_left.t9 a_n1712_n1088# 0.097082f
C69 drain_left.t2 a_n1712_n1088# 0.015607f
C70 drain_left.t6 a_n1712_n1088# 0.015607f
C71 drain_left.n0 a_n1712_n1088# 0.060645f
C72 drain_left.n1 a_n1712_n1088# 0.392955f
C73 drain_left.t3 a_n1712_n1088# 0.015607f
C74 drain_left.t5 a_n1712_n1088# 0.015607f
C75 drain_left.n2 a_n1712_n1088# 0.061092f
C76 drain_left.n3 a_n1712_n1088# 0.736412f
C77 drain_left.t8 a_n1712_n1088# 0.097082f
C78 drain_left.t4 a_n1712_n1088# 0.015607f
C79 drain_left.t0 a_n1712_n1088# 0.015607f
C80 drain_left.n4 a_n1712_n1088# 0.060645f
C81 drain_left.n5 a_n1712_n1088# 0.426922f
C82 drain_left.t7 a_n1712_n1088# 0.015607f
C83 drain_left.t1 a_n1712_n1088# 0.015607f
C84 drain_left.n6 a_n1712_n1088# 0.060645f
C85 drain_left.n7 a_n1712_n1088# 0.39887f
C86 source.t16 a_n1712_n1088# 0.119681f
C87 source.n0 a_n1712_n1088# 0.540935f
C88 source.t17 a_n1712_n1088# 0.021503f
C89 source.t14 a_n1712_n1088# 0.021503f
C90 source.n1 a_n1712_n1088# 0.069737f
C91 source.n2 a_n1712_n1088# 0.292591f
C92 source.t19 a_n1712_n1088# 0.021503f
C93 source.t10 a_n1712_n1088# 0.021503f
C94 source.n3 a_n1712_n1088# 0.069737f
C95 source.n4 a_n1712_n1088# 0.302417f
C96 source.t7 a_n1712_n1088# 0.119681f
C97 source.n5 a_n1712_n1088# 0.311117f
C98 source.t1 a_n1712_n1088# 0.021503f
C99 source.t8 a_n1712_n1088# 0.021503f
C100 source.n6 a_n1712_n1088# 0.069737f
C101 source.n7 a_n1712_n1088# 0.292591f
C102 source.t4 a_n1712_n1088# 0.021503f
C103 source.t9 a_n1712_n1088# 0.021503f
C104 source.n8 a_n1712_n1088# 0.069737f
C105 source.n9 a_n1712_n1088# 0.816203f
C106 source.t11 a_n1712_n1088# 0.021503f
C107 source.t12 a_n1712_n1088# 0.021503f
C108 source.n10 a_n1712_n1088# 0.069737f
C109 source.n11 a_n1712_n1088# 0.816204f
C110 source.t18 a_n1712_n1088# 0.021503f
C111 source.t13 a_n1712_n1088# 0.021503f
C112 source.n12 a_n1712_n1088# 0.069737f
C113 source.n13 a_n1712_n1088# 0.292591f
C114 source.t15 a_n1712_n1088# 0.119681f
C115 source.n14 a_n1712_n1088# 0.311117f
C116 source.t5 a_n1712_n1088# 0.021503f
C117 source.t0 a_n1712_n1088# 0.021503f
C118 source.n15 a_n1712_n1088# 0.069737f
C119 source.n16 a_n1712_n1088# 0.302418f
C120 source.t3 a_n1712_n1088# 0.021503f
C121 source.t6 a_n1712_n1088# 0.021503f
C122 source.n17 a_n1712_n1088# 0.069737f
C123 source.n18 a_n1712_n1088# 0.292591f
C124 source.t2 a_n1712_n1088# 0.119681f
C125 source.n19 a_n1712_n1088# 0.445367f
C126 source.n20 a_n1712_n1088# 0.557387f
C127 plus.n0 a_n1712_n1088# 0.032004f
C128 plus.t8 a_n1712_n1088# 0.054263f
C129 plus.t2 a_n1712_n1088# 0.054263f
C130 plus.t9 a_n1712_n1088# 0.054263f
C131 plus.n1 a_n1712_n1088# 0.059797f
C132 plus.t1 a_n1712_n1088# 0.062285f
C133 plus.n2 a_n1712_n1088# 0.048655f
C134 plus.t5 a_n1712_n1088# 0.054263f
C135 plus.n3 a_n1712_n1088# 0.058021f
C136 plus.n4 a_n1712_n1088# 0.007262f
C137 plus.n5 a_n1712_n1088# 0.102093f
C138 plus.n6 a_n1712_n1088# 0.032004f
C139 plus.n7 a_n1712_n1088# 0.032004f
C140 plus.n8 a_n1712_n1088# 0.007262f
C141 plus.n9 a_n1712_n1088# 0.058021f
C142 plus.n10 a_n1712_n1088# 0.056443f
C143 plus.n11 a_n1712_n1088# 0.224412f
C144 plus.n12 a_n1712_n1088# 0.032004f
C145 plus.t0 a_n1712_n1088# 0.054263f
C146 plus.t7 a_n1712_n1088# 0.054263f
C147 plus.t3 a_n1712_n1088# 0.054263f
C148 plus.n13 a_n1712_n1088# 0.059797f
C149 plus.t4 a_n1712_n1088# 0.062285f
C150 plus.n14 a_n1712_n1088# 0.048655f
C151 plus.t6 a_n1712_n1088# 0.054263f
C152 plus.n15 a_n1712_n1088# 0.058021f
C153 plus.n16 a_n1712_n1088# 0.007262f
C154 plus.n17 a_n1712_n1088# 0.102093f
C155 plus.n18 a_n1712_n1088# 0.032004f
C156 plus.n19 a_n1712_n1088# 0.032004f
C157 plus.n20 a_n1712_n1088# 0.007262f
C158 plus.n21 a_n1712_n1088# 0.058021f
C159 plus.n22 a_n1712_n1088# 0.056443f
C160 plus.n23 a_n1712_n1088# 0.689347f
.ends

