* NGSPICE file created from diffpair581.ext - technology: sky130A

.subckt diffpair581 minus drain_right drain_left source plus
X0 drain_right minus source a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X1 a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X2 source plus drain_left a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X3 a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X4 drain_left plus source a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X5 drain_left plus source a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X6 source minus drain_right a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X7 source minus drain_right a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X8 a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X9 source plus drain_left a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X10 drain_right minus source a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X11 a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# a_n1064_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
.ends

