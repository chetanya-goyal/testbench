* NGSPICE file created from diffpair177.ext - technology: sky130A

.subckt diffpair177 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t17 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X1 drain_right.t15 minus.t0 source.t13 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X2 drain_right.t14 minus.t1 source.t1 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X3 source.t8 minus.t2 drain_right.t13 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X4 drain_right.t12 minus.t3 source.t11 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X5 source.t31 plus.t1 drain_left.t14 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X6 a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.2
X7 source.t16 plus.t2 drain_left.t13 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X8 drain_left.t12 plus.t3 source.t29 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X9 source.t6 minus.t4 drain_right.t11 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X10 a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X11 drain_left.t11 plus.t4 source.t26 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X12 a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X13 source.t9 minus.t5 drain_right.t10 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X14 source.t5 minus.t6 drain_right.t9 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X15 source.t10 minus.t7 drain_right.t8 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X16 drain_left.t10 plus.t5 source.t18 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X17 drain_left.t9 plus.t6 source.t28 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X18 source.t23 plus.t7 drain_left.t8 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X19 drain_right.t7 minus.t8 source.t12 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X20 source.t24 plus.t8 drain_left.t7 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X21 a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.2
X22 source.t30 plus.t9 drain_left.t6 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X23 drain_right.t6 minus.t9 source.t3 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X24 drain_right.t5 minus.t10 source.t0 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X25 drain_right.t4 minus.t11 source.t2 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X26 drain_left.t5 plus.t10 source.t21 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X27 source.t27 plus.t11 drain_left.t4 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X28 drain_left.t3 plus.t12 source.t25 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X29 source.t4 minus.t12 drain_right.t3 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X30 source.t14 minus.t13 drain_right.t2 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X31 drain_right.t1 minus.t14 source.t7 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X32 source.t22 plus.t13 drain_left.t2 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.2
X33 drain_left.t1 plus.t14 source.t19 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.2
X34 source.t20 plus.t15 drain_left.t0 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
X35 source.t15 minus.t15 drain_right.t0 a_n1670_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.2
R0 plus.n4 plus.t7 570.003
R1 plus.n17 plus.t14 570.003
R2 plus.n23 plus.t4 570.003
R3 plus.n36 plus.t13 570.003
R4 plus.n3 plus.t3 518.15
R5 plus.n7 plus.t15 518.15
R6 plus.n9 plus.t12 518.15
R7 plus.n1 plus.t11 518.15
R8 plus.n14 plus.t6 518.15
R9 plus.n16 plus.t2 518.15
R10 plus.n22 plus.t9 518.15
R11 plus.n26 plus.t0 518.15
R12 plus.n28 plus.t8 518.15
R13 plus.n20 plus.t10 518.15
R14 plus.n33 plus.t1 518.15
R15 plus.n35 plus.t5 518.15
R16 plus.n5 plus.n4 161.489
R17 plus.n24 plus.n23 161.489
R18 plus.n6 plus.n5 161.3
R19 plus.n8 plus.n2 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n0 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n25 plus.n24 161.3
R25 plus.n27 plus.n21 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n19 161.3
R29 plus.n37 plus.n36 161.3
R30 plus.n6 plus.n3 47.4702
R31 plus.n16 plus.n15 47.4702
R32 plus.n35 plus.n34 47.4702
R33 plus.n25 plus.n22 47.4702
R34 plus.n8 plus.n7 43.0884
R35 plus.n14 plus.n13 43.0884
R36 plus.n33 plus.n32 43.0884
R37 plus.n27 plus.n26 43.0884
R38 plus.n10 plus.n9 38.7066
R39 plus.n10 plus.n1 38.7066
R40 plus.n29 plus.n20 38.7066
R41 plus.n29 plus.n28 38.7066
R42 plus.n9 plus.n8 34.3247
R43 plus.n13 plus.n1 34.3247
R44 plus.n32 plus.n20 34.3247
R45 plus.n28 plus.n27 34.3247
R46 plus.n7 plus.n6 29.9429
R47 plus.n15 plus.n14 29.9429
R48 plus.n34 plus.n33 29.9429
R49 plus.n26 plus.n25 29.9429
R50 plus plus.n37 25.8854
R51 plus.n4 plus.n3 25.5611
R52 plus.n17 plus.n16 25.5611
R53 plus.n36 plus.n35 25.5611
R54 plus.n23 plus.n22 25.5611
R55 plus plus.n18 8.70126
R56 plus.n5 plus.n2 0.189894
R57 plus.n11 plus.n2 0.189894
R58 plus.n12 plus.n11 0.189894
R59 plus.n12 plus.n0 0.189894
R60 plus.n18 plus.n0 0.189894
R61 plus.n37 plus.n19 0.189894
R62 plus.n31 plus.n19 0.189894
R63 plus.n31 plus.n30 0.189894
R64 plus.n30 plus.n21 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n0 source.t19 69.6943
R67 source.n7 source.t23 69.6943
R68 source.n8 source.t0 69.6943
R69 source.n15 source.t14 69.6943
R70 source.n31 source.t3 69.6942
R71 source.n24 source.t6 69.6942
R72 source.n23 source.t26 69.6942
R73 source.n16 source.t22 69.6942
R74 source.n2 source.n1 63.0943
R75 source.n4 source.n3 63.0943
R76 source.n6 source.n5 63.0943
R77 source.n10 source.n9 63.0943
R78 source.n12 source.n11 63.0943
R79 source.n14 source.n13 63.0943
R80 source.n30 source.n29 63.0942
R81 source.n28 source.n27 63.0942
R82 source.n26 source.n25 63.0942
R83 source.n22 source.n21 63.0942
R84 source.n20 source.n19 63.0942
R85 source.n18 source.n17 63.0942
R86 source.n16 source.n15 14.9264
R87 source.n32 source.n0 9.43506
R88 source.n29 source.t7 6.6005
R89 source.n29 source.t8 6.6005
R90 source.n27 source.t11 6.6005
R91 source.n27 source.t10 6.6005
R92 source.n25 source.t12 6.6005
R93 source.n25 source.t15 6.6005
R94 source.n21 source.t17 6.6005
R95 source.n21 source.t30 6.6005
R96 source.n19 source.t21 6.6005
R97 source.n19 source.t24 6.6005
R98 source.n17 source.t18 6.6005
R99 source.n17 source.t31 6.6005
R100 source.n1 source.t28 6.6005
R101 source.n1 source.t16 6.6005
R102 source.n3 source.t25 6.6005
R103 source.n3 source.t27 6.6005
R104 source.n5 source.t29 6.6005
R105 source.n5 source.t20 6.6005
R106 source.n9 source.t13 6.6005
R107 source.n9 source.t5 6.6005
R108 source.n11 source.t2 6.6005
R109 source.n11 source.t4 6.6005
R110 source.n13 source.t1 6.6005
R111 source.n13 source.t9 6.6005
R112 source.n32 source.n31 5.49188
R113 source.n8 source.n7 0.470328
R114 source.n24 source.n23 0.470328
R115 source.n15 source.n14 0.457397
R116 source.n14 source.n12 0.457397
R117 source.n12 source.n10 0.457397
R118 source.n10 source.n8 0.457397
R119 source.n7 source.n6 0.457397
R120 source.n6 source.n4 0.457397
R121 source.n4 source.n2 0.457397
R122 source.n2 source.n0 0.457397
R123 source.n18 source.n16 0.457397
R124 source.n20 source.n18 0.457397
R125 source.n22 source.n20 0.457397
R126 source.n23 source.n22 0.457397
R127 source.n26 source.n24 0.457397
R128 source.n28 source.n26 0.457397
R129 source.n30 source.n28 0.457397
R130 source.n31 source.n30 0.457397
R131 source source.n32 0.188
R132 drain_left.n9 drain_left.n7 80.23
R133 drain_left.n5 drain_left.n3 80.2299
R134 drain_left.n2 drain_left.n0 80.2299
R135 drain_left.n13 drain_left.n12 79.7731
R136 drain_left.n11 drain_left.n10 79.7731
R137 drain_left.n9 drain_left.n8 79.7731
R138 drain_left.n5 drain_left.n4 79.773
R139 drain_left.n2 drain_left.n1 79.773
R140 drain_left drain_left.n6 23.5187
R141 drain_left.n3 drain_left.t6 6.6005
R142 drain_left.n3 drain_left.t11 6.6005
R143 drain_left.n4 drain_left.t7 6.6005
R144 drain_left.n4 drain_left.t15 6.6005
R145 drain_left.n1 drain_left.t14 6.6005
R146 drain_left.n1 drain_left.t5 6.6005
R147 drain_left.n0 drain_left.t2 6.6005
R148 drain_left.n0 drain_left.t10 6.6005
R149 drain_left.n12 drain_left.t13 6.6005
R150 drain_left.n12 drain_left.t1 6.6005
R151 drain_left.n10 drain_left.t4 6.6005
R152 drain_left.n10 drain_left.t9 6.6005
R153 drain_left.n8 drain_left.t0 6.6005
R154 drain_left.n8 drain_left.t3 6.6005
R155 drain_left.n7 drain_left.t8 6.6005
R156 drain_left.n7 drain_left.t12 6.6005
R157 drain_left drain_left.n13 6.11011
R158 drain_left.n11 drain_left.n9 0.457397
R159 drain_left.n13 drain_left.n11 0.457397
R160 drain_left.n6 drain_left.n5 0.173602
R161 drain_left.n6 drain_left.n2 0.173602
R162 minus.n17 minus.t13 570.003
R163 minus.n4 minus.t10 570.003
R164 minus.n36 minus.t9 570.003
R165 minus.n23 minus.t4 570.003
R166 minus.n16 minus.t1 518.15
R167 minus.n14 minus.t5 518.15
R168 minus.n1 minus.t11 518.15
R169 minus.n9 minus.t12 518.15
R170 minus.n7 minus.t0 518.15
R171 minus.n3 minus.t6 518.15
R172 minus.n35 minus.t2 518.15
R173 minus.n33 minus.t14 518.15
R174 minus.n20 minus.t7 518.15
R175 minus.n28 minus.t3 518.15
R176 minus.n26 minus.t15 518.15
R177 minus.n22 minus.t8 518.15
R178 minus.n5 minus.n4 161.489
R179 minus.n24 minus.n23 161.489
R180 minus.n18 minus.n17 161.3
R181 minus.n15 minus.n0 161.3
R182 minus.n13 minus.n12 161.3
R183 minus.n11 minus.n10 161.3
R184 minus.n8 minus.n2 161.3
R185 minus.n6 minus.n5 161.3
R186 minus.n37 minus.n36 161.3
R187 minus.n34 minus.n19 161.3
R188 minus.n32 minus.n31 161.3
R189 minus.n30 minus.n29 161.3
R190 minus.n27 minus.n21 161.3
R191 minus.n25 minus.n24 161.3
R192 minus.n16 minus.n15 47.4702
R193 minus.n6 minus.n3 47.4702
R194 minus.n25 minus.n22 47.4702
R195 minus.n35 minus.n34 47.4702
R196 minus.n14 minus.n13 43.0884
R197 minus.n8 minus.n7 43.0884
R198 minus.n27 minus.n26 43.0884
R199 minus.n33 minus.n32 43.0884
R200 minus.n10 minus.n1 38.7066
R201 minus.n10 minus.n9 38.7066
R202 minus.n29 minus.n28 38.7066
R203 minus.n29 minus.n20 38.7066
R204 minus.n13 minus.n1 34.3247
R205 minus.n9 minus.n8 34.3247
R206 minus.n28 minus.n27 34.3247
R207 minus.n32 minus.n20 34.3247
R208 minus.n15 minus.n14 29.9429
R209 minus.n7 minus.n6 29.9429
R210 minus.n26 minus.n25 29.9429
R211 minus.n34 minus.n33 29.9429
R212 minus.n38 minus.n18 28.5952
R213 minus.n17 minus.n16 25.5611
R214 minus.n4 minus.n3 25.5611
R215 minus.n23 minus.n22 25.5611
R216 minus.n36 minus.n35 25.5611
R217 minus.n38 minus.n37 6.46641
R218 minus.n18 minus.n0 0.189894
R219 minus.n12 minus.n0 0.189894
R220 minus.n12 minus.n11 0.189894
R221 minus.n11 minus.n2 0.189894
R222 minus.n5 minus.n2 0.189894
R223 minus.n24 minus.n21 0.189894
R224 minus.n30 minus.n21 0.189894
R225 minus.n31 minus.n30 0.189894
R226 minus.n31 minus.n19 0.189894
R227 minus.n37 minus.n19 0.189894
R228 minus minus.n38 0.188
R229 drain_right.n9 drain_right.n7 80.23
R230 drain_right.n5 drain_right.n3 80.2299
R231 drain_right.n2 drain_right.n0 80.2299
R232 drain_right.n9 drain_right.n8 79.7731
R233 drain_right.n11 drain_right.n10 79.7731
R234 drain_right.n13 drain_right.n12 79.7731
R235 drain_right.n5 drain_right.n4 79.773
R236 drain_right.n2 drain_right.n1 79.773
R237 drain_right drain_right.n6 22.9655
R238 drain_right.n3 drain_right.t13 6.6005
R239 drain_right.n3 drain_right.t6 6.6005
R240 drain_right.n4 drain_right.t8 6.6005
R241 drain_right.n4 drain_right.t1 6.6005
R242 drain_right.n1 drain_right.t0 6.6005
R243 drain_right.n1 drain_right.t12 6.6005
R244 drain_right.n0 drain_right.t11 6.6005
R245 drain_right.n0 drain_right.t7 6.6005
R246 drain_right.n7 drain_right.t9 6.6005
R247 drain_right.n7 drain_right.t5 6.6005
R248 drain_right.n8 drain_right.t3 6.6005
R249 drain_right.n8 drain_right.t15 6.6005
R250 drain_right.n10 drain_right.t10 6.6005
R251 drain_right.n10 drain_right.t4 6.6005
R252 drain_right.n12 drain_right.t2 6.6005
R253 drain_right.n12 drain_right.t14 6.6005
R254 drain_right drain_right.n13 6.11011
R255 drain_right.n13 drain_right.n11 0.457397
R256 drain_right.n11 drain_right.n9 0.457397
R257 drain_right.n6 drain_right.n5 0.173602
R258 drain_right.n6 drain_right.n2 0.173602
C0 drain_left plus 1.6427f
C1 drain_left minus 0.175878f
C2 plus minus 3.57726f
C3 source drain_right 11.2064f
C4 drain_left drain_right 0.846053f
C5 drain_left source 11.2068f
C6 plus drain_right 0.320188f
C7 plus source 1.55247f
C8 minus drain_right 1.48171f
C9 source minus 1.53847f
C10 drain_right a_n1670_n1488# 4.21327f
C11 drain_left a_n1670_n1488# 4.45429f
C12 source a_n1670_n1488# 3.595316f
C13 minus a_n1670_n1488# 5.753903f
C14 plus a_n1670_n1488# 6.423742f
C15 drain_right.t11 a_n1670_n1488# 0.075242f
C16 drain_right.t7 a_n1670_n1488# 0.075242f
C17 drain_right.n0 a_n1670_n1488# 0.544688f
C18 drain_right.t0 a_n1670_n1488# 0.075242f
C19 drain_right.t12 a_n1670_n1488# 0.075242f
C20 drain_right.n1 a_n1670_n1488# 0.542636f
C21 drain_right.n2 a_n1670_n1488# 0.680984f
C22 drain_right.t13 a_n1670_n1488# 0.075242f
C23 drain_right.t6 a_n1670_n1488# 0.075242f
C24 drain_right.n3 a_n1670_n1488# 0.544688f
C25 drain_right.t8 a_n1670_n1488# 0.075242f
C26 drain_right.t1 a_n1670_n1488# 0.075242f
C27 drain_right.n4 a_n1670_n1488# 0.542636f
C28 drain_right.n5 a_n1670_n1488# 0.680984f
C29 drain_right.n6 a_n1670_n1488# 0.833476f
C30 drain_right.t9 a_n1670_n1488# 0.075242f
C31 drain_right.t5 a_n1670_n1488# 0.075242f
C32 drain_right.n7 a_n1670_n1488# 0.544691f
C33 drain_right.t3 a_n1670_n1488# 0.075242f
C34 drain_right.t15 a_n1670_n1488# 0.075242f
C35 drain_right.n8 a_n1670_n1488# 0.542639f
C36 drain_right.n9 a_n1670_n1488# 0.705752f
C37 drain_right.t10 a_n1670_n1488# 0.075242f
C38 drain_right.t4 a_n1670_n1488# 0.075242f
C39 drain_right.n10 a_n1670_n1488# 0.542639f
C40 drain_right.n11 a_n1670_n1488# 0.34751f
C41 drain_right.t2 a_n1670_n1488# 0.075242f
C42 drain_right.t14 a_n1670_n1488# 0.075242f
C43 drain_right.n12 a_n1670_n1488# 0.542639f
C44 drain_right.n13 a_n1670_n1488# 0.607258f
C45 minus.n0 a_n1670_n1488# 0.029091f
C46 minus.t13 a_n1670_n1488# 0.053578f
C47 minus.t1 a_n1670_n1488# 0.050546f
C48 minus.t5 a_n1670_n1488# 0.050546f
C49 minus.t11 a_n1670_n1488# 0.050546f
C50 minus.n1 a_n1670_n1488# 0.032339f
C51 minus.n2 a_n1670_n1488# 0.029091f
C52 minus.t12 a_n1670_n1488# 0.050546f
C53 minus.t0 a_n1670_n1488# 0.050546f
C54 minus.t6 a_n1670_n1488# 0.050546f
C55 minus.n3 a_n1670_n1488# 0.032339f
C56 minus.t10 a_n1670_n1488# 0.053578f
C57 minus.n4 a_n1670_n1488# 0.040525f
C58 minus.n5 a_n1670_n1488# 0.065492f
C59 minus.n6 a_n1670_n1488# 0.010188f
C60 minus.n7 a_n1670_n1488# 0.032339f
C61 minus.n8 a_n1670_n1488# 0.010188f
C62 minus.n9 a_n1670_n1488# 0.032339f
C63 minus.n10 a_n1670_n1488# 0.010188f
C64 minus.n11 a_n1670_n1488# 0.029091f
C65 minus.n12 a_n1670_n1488# 0.029091f
C66 minus.n13 a_n1670_n1488# 0.010188f
C67 minus.n14 a_n1670_n1488# 0.032339f
C68 minus.n15 a_n1670_n1488# 0.010188f
C69 minus.n16 a_n1670_n1488# 0.032339f
C70 minus.n17 a_n1670_n1488# 0.040482f
C71 minus.n18 a_n1670_n1488# 0.695603f
C72 minus.n19 a_n1670_n1488# 0.029091f
C73 minus.t2 a_n1670_n1488# 0.050546f
C74 minus.t14 a_n1670_n1488# 0.050546f
C75 minus.t7 a_n1670_n1488# 0.050546f
C76 minus.n20 a_n1670_n1488# 0.032339f
C77 minus.n21 a_n1670_n1488# 0.029091f
C78 minus.t3 a_n1670_n1488# 0.050546f
C79 minus.t15 a_n1670_n1488# 0.050546f
C80 minus.t8 a_n1670_n1488# 0.050546f
C81 minus.n22 a_n1670_n1488# 0.032339f
C82 minus.t4 a_n1670_n1488# 0.053578f
C83 minus.n23 a_n1670_n1488# 0.040525f
C84 minus.n24 a_n1670_n1488# 0.065492f
C85 minus.n25 a_n1670_n1488# 0.010188f
C86 minus.n26 a_n1670_n1488# 0.032339f
C87 minus.n27 a_n1670_n1488# 0.010188f
C88 minus.n28 a_n1670_n1488# 0.032339f
C89 minus.n29 a_n1670_n1488# 0.010188f
C90 minus.n30 a_n1670_n1488# 0.029091f
C91 minus.n31 a_n1670_n1488# 0.029091f
C92 minus.n32 a_n1670_n1488# 0.010188f
C93 minus.n33 a_n1670_n1488# 0.032339f
C94 minus.n34 a_n1670_n1488# 0.010188f
C95 minus.n35 a_n1670_n1488# 0.032339f
C96 minus.t9 a_n1670_n1488# 0.053578f
C97 minus.n36 a_n1670_n1488# 0.040482f
C98 minus.n37 a_n1670_n1488# 0.187882f
C99 minus.n38 a_n1670_n1488# 0.860876f
C100 drain_left.t2 a_n1670_n1488# 0.074417f
C101 drain_left.t10 a_n1670_n1488# 0.074417f
C102 drain_left.n0 a_n1670_n1488# 0.538716f
C103 drain_left.t14 a_n1670_n1488# 0.074417f
C104 drain_left.t5 a_n1670_n1488# 0.074417f
C105 drain_left.n1 a_n1670_n1488# 0.536687f
C106 drain_left.n2 a_n1670_n1488# 0.673518f
C107 drain_left.t6 a_n1670_n1488# 0.074417f
C108 drain_left.t11 a_n1670_n1488# 0.074417f
C109 drain_left.n3 a_n1670_n1488# 0.538716f
C110 drain_left.t7 a_n1670_n1488# 0.074417f
C111 drain_left.t15 a_n1670_n1488# 0.074417f
C112 drain_left.n4 a_n1670_n1488# 0.536687f
C113 drain_left.n5 a_n1670_n1488# 0.673518f
C114 drain_left.n6 a_n1670_n1488# 0.886663f
C115 drain_left.t8 a_n1670_n1488# 0.074417f
C116 drain_left.t12 a_n1670_n1488# 0.074417f
C117 drain_left.n7 a_n1670_n1488# 0.538719f
C118 drain_left.t0 a_n1670_n1488# 0.074417f
C119 drain_left.t3 a_n1670_n1488# 0.074417f
C120 drain_left.n8 a_n1670_n1488# 0.53669f
C121 drain_left.n9 a_n1670_n1488# 0.698014f
C122 drain_left.t4 a_n1670_n1488# 0.074417f
C123 drain_left.t9 a_n1670_n1488# 0.074417f
C124 drain_left.n10 a_n1670_n1488# 0.53669f
C125 drain_left.n11 a_n1670_n1488# 0.3437f
C126 drain_left.t13 a_n1670_n1488# 0.074417f
C127 drain_left.t1 a_n1670_n1488# 0.074417f
C128 drain_left.n12 a_n1670_n1488# 0.53669f
C129 drain_left.n13 a_n1670_n1488# 0.6006f
C130 source.t19 a_n1670_n1488# 0.597538f
C131 source.n0 a_n1670_n1488# 0.800383f
C132 source.t28 a_n1670_n1488# 0.071959f
C133 source.t16 a_n1670_n1488# 0.071959f
C134 source.n1 a_n1670_n1488# 0.456264f
C135 source.n2 a_n1670_n1488# 0.353796f
C136 source.t25 a_n1670_n1488# 0.071959f
C137 source.t27 a_n1670_n1488# 0.071959f
C138 source.n3 a_n1670_n1488# 0.456264f
C139 source.n4 a_n1670_n1488# 0.353796f
C140 source.t29 a_n1670_n1488# 0.071959f
C141 source.t20 a_n1670_n1488# 0.071959f
C142 source.n5 a_n1670_n1488# 0.456264f
C143 source.n6 a_n1670_n1488# 0.353796f
C144 source.t23 a_n1670_n1488# 0.597538f
C145 source.n7 a_n1670_n1488# 0.410039f
C146 source.t0 a_n1670_n1488# 0.597538f
C147 source.n8 a_n1670_n1488# 0.410039f
C148 source.t13 a_n1670_n1488# 0.071959f
C149 source.t5 a_n1670_n1488# 0.071959f
C150 source.n9 a_n1670_n1488# 0.456264f
C151 source.n10 a_n1670_n1488# 0.353796f
C152 source.t2 a_n1670_n1488# 0.071959f
C153 source.t4 a_n1670_n1488# 0.071959f
C154 source.n11 a_n1670_n1488# 0.456264f
C155 source.n12 a_n1670_n1488# 0.353796f
C156 source.t1 a_n1670_n1488# 0.071959f
C157 source.t9 a_n1670_n1488# 0.071959f
C158 source.n13 a_n1670_n1488# 0.456264f
C159 source.n14 a_n1670_n1488# 0.353796f
C160 source.t14 a_n1670_n1488# 0.597538f
C161 source.n15 a_n1670_n1488# 1.11478f
C162 source.t22 a_n1670_n1488# 0.597535f
C163 source.n16 a_n1670_n1488# 1.11478f
C164 source.t18 a_n1670_n1488# 0.071959f
C165 source.t31 a_n1670_n1488# 0.071959f
C166 source.n17 a_n1670_n1488# 0.456261f
C167 source.n18 a_n1670_n1488# 0.353799f
C168 source.t21 a_n1670_n1488# 0.071959f
C169 source.t24 a_n1670_n1488# 0.071959f
C170 source.n19 a_n1670_n1488# 0.456261f
C171 source.n20 a_n1670_n1488# 0.353799f
C172 source.t17 a_n1670_n1488# 0.071959f
C173 source.t30 a_n1670_n1488# 0.071959f
C174 source.n21 a_n1670_n1488# 0.456261f
C175 source.n22 a_n1670_n1488# 0.353799f
C176 source.t26 a_n1670_n1488# 0.597535f
C177 source.n23 a_n1670_n1488# 0.410042f
C178 source.t6 a_n1670_n1488# 0.597535f
C179 source.n24 a_n1670_n1488# 0.410042f
C180 source.t12 a_n1670_n1488# 0.071959f
C181 source.t15 a_n1670_n1488# 0.071959f
C182 source.n25 a_n1670_n1488# 0.456261f
C183 source.n26 a_n1670_n1488# 0.353799f
C184 source.t11 a_n1670_n1488# 0.071959f
C185 source.t10 a_n1670_n1488# 0.071959f
C186 source.n27 a_n1670_n1488# 0.456261f
C187 source.n28 a_n1670_n1488# 0.353799f
C188 source.t7 a_n1670_n1488# 0.071959f
C189 source.t8 a_n1670_n1488# 0.071959f
C190 source.n29 a_n1670_n1488# 0.456261f
C191 source.n30 a_n1670_n1488# 0.353799f
C192 source.t3 a_n1670_n1488# 0.597535f
C193 source.n31 a_n1670_n1488# 0.57463f
C194 source.n32 a_n1670_n1488# 0.876133f
C195 plus.n0 a_n1670_n1488# 0.029574f
C196 plus.t2 a_n1670_n1488# 0.051386f
C197 plus.t6 a_n1670_n1488# 0.051386f
C198 plus.t11 a_n1670_n1488# 0.051386f
C199 plus.n1 a_n1670_n1488# 0.032876f
C200 plus.n2 a_n1670_n1488# 0.029574f
C201 plus.t12 a_n1670_n1488# 0.051386f
C202 plus.t15 a_n1670_n1488# 0.051386f
C203 plus.t3 a_n1670_n1488# 0.051386f
C204 plus.n3 a_n1670_n1488# 0.032876f
C205 plus.t7 a_n1670_n1488# 0.054468f
C206 plus.n4 a_n1670_n1488# 0.041198f
C207 plus.n5 a_n1670_n1488# 0.06658f
C208 plus.n6 a_n1670_n1488# 0.010358f
C209 plus.n7 a_n1670_n1488# 0.032876f
C210 plus.n8 a_n1670_n1488# 0.010358f
C211 plus.n9 a_n1670_n1488# 0.032876f
C212 plus.n10 a_n1670_n1488# 0.010358f
C213 plus.n11 a_n1670_n1488# 0.029574f
C214 plus.n12 a_n1670_n1488# 0.029574f
C215 plus.n13 a_n1670_n1488# 0.010358f
C216 plus.n14 a_n1670_n1488# 0.032876f
C217 plus.n15 a_n1670_n1488# 0.010358f
C218 plus.n16 a_n1670_n1488# 0.032876f
C219 plus.t14 a_n1670_n1488# 0.054468f
C220 plus.n17 a_n1670_n1488# 0.041155f
C221 plus.n18 a_n1670_n1488# 0.218449f
C222 plus.n19 a_n1670_n1488# 0.029574f
C223 plus.t13 a_n1670_n1488# 0.054468f
C224 plus.t5 a_n1670_n1488# 0.051386f
C225 plus.t1 a_n1670_n1488# 0.051386f
C226 plus.t10 a_n1670_n1488# 0.051386f
C227 plus.n20 a_n1670_n1488# 0.032876f
C228 plus.n21 a_n1670_n1488# 0.029574f
C229 plus.t8 a_n1670_n1488# 0.051386f
C230 plus.t0 a_n1670_n1488# 0.051386f
C231 plus.t9 a_n1670_n1488# 0.051386f
C232 plus.n22 a_n1670_n1488# 0.032876f
C233 plus.t4 a_n1670_n1488# 0.054468f
C234 plus.n23 a_n1670_n1488# 0.041198f
C235 plus.n24 a_n1670_n1488# 0.06658f
C236 plus.n25 a_n1670_n1488# 0.010358f
C237 plus.n26 a_n1670_n1488# 0.032876f
C238 plus.n27 a_n1670_n1488# 0.010358f
C239 plus.n28 a_n1670_n1488# 0.032876f
C240 plus.n29 a_n1670_n1488# 0.010358f
C241 plus.n30 a_n1670_n1488# 0.029574f
C242 plus.n31 a_n1670_n1488# 0.029574f
C243 plus.n32 a_n1670_n1488# 0.010358f
C244 plus.n33 a_n1670_n1488# 0.032876f
C245 plus.n34 a_n1670_n1488# 0.010358f
C246 plus.n35 a_n1670_n1488# 0.032876f
C247 plus.n36 a_n1670_n1488# 0.041155f
C248 plus.n37 a_n1670_n1488# 0.665894f
.ends

