* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right minus source a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=1.425 ps=6.95 w=3 l=0.15
X1 drain_right minus source a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=1.425 ps=6.95 w=3 l=0.15
X2 drain_left plus source a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=1.425 ps=6.95 w=3 l=0.15
X3 a_n976_n1492# a_n976_n1492# a_n976_n1492# a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X4 drain_left plus source a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=1.425 ps=6.95 w=3 l=0.15
X5 a_n976_n1492# a_n976_n1492# a_n976_n1492# a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X6 a_n976_n1492# a_n976_n1492# a_n976_n1492# a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X7 a_n976_n1492# a_n976_n1492# a_n976_n1492# a_n976_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
.ends

