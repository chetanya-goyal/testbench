* NGSPICE file created from diffpair524.ext - technology: sky130A

.subckt diffpair524 minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t7 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X1 a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X2 drain_left.t4 plus.t1 source.t14 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X3 source.t17 minus.t0 drain_right.t9 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X4 drain_left.t3 plus.t2 source.t13 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X5 source.t12 plus.t3 drain_left.t8 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X6 drain_left.t9 plus.t4 source.t11 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X7 drain_right.t8 minus.t1 source.t18 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X8 source.t19 minus.t2 drain_right.t7 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X9 drain_right.t6 minus.t3 source.t1 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X10 drain_right.t5 minus.t4 source.t0 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X11 a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X12 source.t10 plus.t5 drain_left.t2 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X13 drain_right.t4 minus.t5 source.t2 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X14 drain_left.t0 plus.t6 source.t9 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X16 drain_right.t3 minus.t6 source.t4 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X17 source.t5 minus.t7 drain_right.t2 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X18 drain_right.t1 minus.t8 source.t3 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 source.t8 plus.t7 drain_left.t1 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X20 source.t16 minus.t9 drain_right.t0 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X21 drain_left.t6 plus.t8 source.t7 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X22 drain_left.t5 plus.t9 source.t6 a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X23 a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# a_n1712_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
R0 plus.n2 plus.t2 822.548
R1 plus.n14 plus.t1 822.548
R2 plus.n10 plus.t8 801.567
R3 plus.n9 plus.t5 801.567
R4 plus.n1 plus.t9 801.567
R5 plus.n3 plus.t7 801.567
R6 plus.n22 plus.t4 801.567
R7 plus.n21 plus.t3 801.567
R8 plus.n13 plus.t6 801.567
R9 plus.n15 plus.t0 801.567
R10 plus.n5 plus.n4 161.3
R11 plus.n6 plus.n1 161.3
R12 plus.n8 plus.n7 161.3
R13 plus.n9 plus.n0 161.3
R14 plus.n11 plus.n10 161.3
R15 plus.n17 plus.n16 161.3
R16 plus.n18 plus.n13 161.3
R17 plus.n20 plus.n19 161.3
R18 plus.n21 plus.n12 161.3
R19 plus.n23 plus.n22 161.3
R20 plus.n5 plus.n2 70.4033
R21 plus.n17 plus.n14 70.4033
R22 plus.n10 plus.n9 48.2005
R23 plus.n22 plus.n21 48.2005
R24 plus.n8 plus.n1 36.5157
R25 plus.n4 plus.n1 36.5157
R26 plus.n20 plus.n13 36.5157
R27 plus.n16 plus.n13 36.5157
R28 plus plus.n23 30.6865
R29 plus.n3 plus.n2 20.9576
R30 plus.n15 plus.n14 20.9576
R31 plus plus.n11 13.3433
R32 plus.n9 plus.n8 11.6853
R33 plus.n4 plus.n3 11.6853
R34 plus.n21 plus.n20 11.6853
R35 plus.n16 plus.n15 11.6853
R36 plus.n6 plus.n5 0.189894
R37 plus.n7 plus.n6 0.189894
R38 plus.n7 plus.n0 0.189894
R39 plus.n11 plus.n0 0.189894
R40 plus.n23 plus.n12 0.189894
R41 plus.n19 plus.n12 0.189894
R42 plus.n19 plus.n18 0.189894
R43 plus.n18 plus.n17 0.189894
R44 drain_left.n5 drain_left.t3 62.9153
R45 drain_left.n1 drain_left.t9 62.9151
R46 drain_left.n3 drain_left.n2 61.3609
R47 drain_left.n5 drain_left.n4 60.8798
R48 drain_left.n7 drain_left.n6 60.8796
R49 drain_left.n1 drain_left.n0 60.8796
R50 drain_left drain_left.n3 32.6807
R51 drain_left drain_left.n7 6.36873
R52 drain_left.n2 drain_left.t7 1.3205
R53 drain_left.n2 drain_left.t4 1.3205
R54 drain_left.n0 drain_left.t8 1.3205
R55 drain_left.n0 drain_left.t0 1.3205
R56 drain_left.n6 drain_left.t2 1.3205
R57 drain_left.n6 drain_left.t6 1.3205
R58 drain_left.n4 drain_left.t1 1.3205
R59 drain_left.n4 drain_left.t5 1.3205
R60 drain_left.n7 drain_left.n5 0.716017
R61 drain_left.n3 drain_left.n1 0.124033
R62 source.n5 source.t4 45.521
R63 source.n19 source.t2 45.5208
R64 source.n14 source.t14 45.5208
R65 source.n0 source.t7 45.5208
R66 source.n2 source.n1 44.201
R67 source.n4 source.n3 44.201
R68 source.n7 source.n6 44.201
R69 source.n9 source.n8 44.201
R70 source.n18 source.n17 44.2008
R71 source.n16 source.n15 44.2008
R72 source.n13 source.n12 44.2008
R73 source.n11 source.n10 44.2008
R74 source.n11 source.n9 24.9915
R75 source.n20 source.n0 18.6553
R76 source.n20 source.n19 5.62119
R77 source.n17 source.t3 1.3205
R78 source.n17 source.t5 1.3205
R79 source.n15 source.t1 1.3205
R80 source.n15 source.t19 1.3205
R81 source.n12 source.t9 1.3205
R82 source.n12 source.t15 1.3205
R83 source.n10 source.t11 1.3205
R84 source.n10 source.t12 1.3205
R85 source.n1 source.t6 1.3205
R86 source.n1 source.t10 1.3205
R87 source.n3 source.t13 1.3205
R88 source.n3 source.t8 1.3205
R89 source.n6 source.t0 1.3205
R90 source.n6 source.t17 1.3205
R91 source.n8 source.t18 1.3205
R92 source.n8 source.t16 1.3205
R93 source.n5 source.n4 0.828086
R94 source.n16 source.n14 0.828086
R95 source.n9 source.n7 0.716017
R96 source.n7 source.n5 0.716017
R97 source.n4 source.n2 0.716017
R98 source.n2 source.n0 0.716017
R99 source.n13 source.n11 0.716017
R100 source.n14 source.n13 0.716017
R101 source.n18 source.n16 0.716017
R102 source.n19 source.n18 0.716017
R103 source source.n20 0.188
R104 minus.n2 minus.t6 822.548
R105 minus.n14 minus.t3 822.548
R106 minus.n3 minus.t0 801.567
R107 minus.n1 minus.t4 801.567
R108 minus.n9 minus.t9 801.567
R109 minus.n10 minus.t1 801.567
R110 minus.n15 minus.t2 801.567
R111 minus.n13 minus.t8 801.567
R112 minus.n21 minus.t7 801.567
R113 minus.n22 minus.t5 801.567
R114 minus.n11 minus.n10 161.3
R115 minus.n9 minus.n0 161.3
R116 minus.n8 minus.n7 161.3
R117 minus.n6 minus.n1 161.3
R118 minus.n5 minus.n4 161.3
R119 minus.n23 minus.n22 161.3
R120 minus.n21 minus.n12 161.3
R121 minus.n20 minus.n19 161.3
R122 minus.n18 minus.n13 161.3
R123 minus.n17 minus.n16 161.3
R124 minus.n5 minus.n2 70.4033
R125 minus.n17 minus.n14 70.4033
R126 minus.n10 minus.n9 48.2005
R127 minus.n22 minus.n21 48.2005
R128 minus.n24 minus.n11 37.9418
R129 minus.n4 minus.n1 36.5157
R130 minus.n8 minus.n1 36.5157
R131 minus.n16 minus.n13 36.5157
R132 minus.n20 minus.n13 36.5157
R133 minus.n3 minus.n2 20.9576
R134 minus.n15 minus.n14 20.9576
R135 minus.n4 minus.n3 11.6853
R136 minus.n9 minus.n8 11.6853
R137 minus.n16 minus.n15 11.6853
R138 minus.n21 minus.n20 11.6853
R139 minus.n24 minus.n23 6.563
R140 minus.n11 minus.n0 0.189894
R141 minus.n7 minus.n0 0.189894
R142 minus.n7 minus.n6 0.189894
R143 minus.n6 minus.n5 0.189894
R144 minus.n18 minus.n17 0.189894
R145 minus.n19 minus.n18 0.189894
R146 minus.n19 minus.n12 0.189894
R147 minus.n23 minus.n12 0.189894
R148 minus minus.n24 0.188
R149 drain_right.n1 drain_right.t6 62.9151
R150 drain_right.n7 drain_right.t8 62.1998
R151 drain_right.n6 drain_right.n4 61.5952
R152 drain_right.n3 drain_right.n2 61.3609
R153 drain_right.n6 drain_right.n5 60.8798
R154 drain_right.n1 drain_right.n0 60.8796
R155 drain_right drain_right.n3 32.1275
R156 drain_right drain_right.n7 6.01097
R157 drain_right.n2 drain_right.t2 1.3205
R158 drain_right.n2 drain_right.t4 1.3205
R159 drain_right.n0 drain_right.t7 1.3205
R160 drain_right.n0 drain_right.t1 1.3205
R161 drain_right.n4 drain_right.t9 1.3205
R162 drain_right.n4 drain_right.t3 1.3205
R163 drain_right.n5 drain_right.t0 1.3205
R164 drain_right.n5 drain_right.t5 1.3205
R165 drain_right.n7 drain_right.n6 0.716017
R166 drain_right.n3 drain_right.n1 0.124033
C0 plus minus 5.83804f
C1 minus drain_left 0.171781f
C2 plus drain_left 6.98034f
C3 minus source 6.41372f
C4 plus source 6.42847f
C5 drain_left source 20.284302f
C6 drain_right minus 6.81825f
C7 plus drain_right 0.322593f
C8 drain_right drain_left 0.848261f
C9 drain_right source 20.2735f
C10 drain_right a_n1712_n3888# 7.695251f
C11 drain_left a_n1712_n3888# 7.96693f
C12 source a_n1712_n3888# 7.423024f
C13 minus a_n1712_n3888# 6.863167f
C14 plus a_n1712_n3888# 8.86243f
C15 drain_right.t6 a_n1712_n3888# 3.55994f
C16 drain_right.t7 a_n1712_n3888# 0.308202f
C17 drain_right.t1 a_n1712_n3888# 0.308202f
C18 drain_right.n0 a_n1712_n3888# 2.78579f
C19 drain_right.n1 a_n1712_n3888# 0.637918f
C20 drain_right.t2 a_n1712_n3888# 0.308202f
C21 drain_right.t4 a_n1712_n3888# 0.308202f
C22 drain_right.n2 a_n1712_n3888# 2.78833f
C23 drain_right.n3 a_n1712_n3888# 1.70088f
C24 drain_right.t9 a_n1712_n3888# 0.308202f
C25 drain_right.t3 a_n1712_n3888# 0.308202f
C26 drain_right.n4 a_n1712_n3888# 2.78977f
C27 drain_right.t0 a_n1712_n3888# 0.308202f
C28 drain_right.t5 a_n1712_n3888# 0.308202f
C29 drain_right.n5 a_n1712_n3888# 2.78579f
C30 drain_right.n6 a_n1712_n3888# 0.672205f
C31 drain_right.t8 a_n1712_n3888# 3.55592f
C32 drain_right.n7 a_n1712_n3888# 0.581792f
C33 minus.n0 a_n1712_n3888# 0.047355f
C34 minus.t4 a_n1712_n3888# 1.00927f
C35 minus.n1 a_n1712_n3888# 0.398138f
C36 minus.t6 a_n1712_n3888# 1.0193f
C37 minus.n2 a_n1712_n3888# 0.38349f
C38 minus.t0 a_n1712_n3888# 1.00927f
C39 minus.n3 a_n1712_n3888# 0.395511f
C40 minus.n4 a_n1712_n3888# 0.010746f
C41 minus.n5 a_n1712_n3888# 0.151062f
C42 minus.n6 a_n1712_n3888# 0.047355f
C43 minus.n7 a_n1712_n3888# 0.047355f
C44 minus.n8 a_n1712_n3888# 0.010746f
C45 minus.t9 a_n1712_n3888# 1.00927f
C46 minus.n9 a_n1712_n3888# 0.395511f
C47 minus.t1 a_n1712_n3888# 1.00927f
C48 minus.n10 a_n1712_n3888# 0.393175f
C49 minus.n11 a_n1712_n3888# 1.80253f
C50 minus.n12 a_n1712_n3888# 0.047355f
C51 minus.t8 a_n1712_n3888# 1.00927f
C52 minus.n13 a_n1712_n3888# 0.398138f
C53 minus.t3 a_n1712_n3888# 1.0193f
C54 minus.n14 a_n1712_n3888# 0.38349f
C55 minus.t2 a_n1712_n3888# 1.00927f
C56 minus.n15 a_n1712_n3888# 0.395511f
C57 minus.n16 a_n1712_n3888# 0.010746f
C58 minus.n17 a_n1712_n3888# 0.151062f
C59 minus.n18 a_n1712_n3888# 0.047355f
C60 minus.n19 a_n1712_n3888# 0.047355f
C61 minus.n20 a_n1712_n3888# 0.010746f
C62 minus.t7 a_n1712_n3888# 1.00927f
C63 minus.n21 a_n1712_n3888# 0.395511f
C64 minus.t5 a_n1712_n3888# 1.00927f
C65 minus.n22 a_n1712_n3888# 0.393175f
C66 minus.n23 a_n1712_n3888# 0.316603f
C67 minus.n24 a_n1712_n3888# 2.17614f
C68 source.t7 a_n1712_n3888# 3.55531f
C69 source.n0 a_n1712_n3888# 1.67073f
C70 source.t6 a_n1712_n3888# 0.317251f
C71 source.t10 a_n1712_n3888# 0.317251f
C72 source.n1 a_n1712_n3888# 2.78679f
C73 source.n2 a_n1712_n3888# 0.387047f
C74 source.t13 a_n1712_n3888# 0.317251f
C75 source.t8 a_n1712_n3888# 0.317251f
C76 source.n3 a_n1712_n3888# 2.78679f
C77 source.n4 a_n1712_n3888# 0.396712f
C78 source.t4 a_n1712_n3888# 3.55532f
C79 source.n5 a_n1712_n3888# 0.493413f
C80 source.t0 a_n1712_n3888# 0.317251f
C81 source.t17 a_n1712_n3888# 0.317251f
C82 source.n6 a_n1712_n3888# 2.78679f
C83 source.n7 a_n1712_n3888# 0.387047f
C84 source.t18 a_n1712_n3888# 0.317251f
C85 source.t16 a_n1712_n3888# 0.317251f
C86 source.n8 a_n1712_n3888# 2.78679f
C87 source.n9 a_n1712_n3888# 2.08648f
C88 source.t11 a_n1712_n3888# 0.317251f
C89 source.t12 a_n1712_n3888# 0.317251f
C90 source.n10 a_n1712_n3888# 2.78678f
C91 source.n11 a_n1712_n3888# 2.08648f
C92 source.t9 a_n1712_n3888# 0.317251f
C93 source.t15 a_n1712_n3888# 0.317251f
C94 source.n12 a_n1712_n3888# 2.78678f
C95 source.n13 a_n1712_n3888# 0.387051f
C96 source.t14 a_n1712_n3888# 3.55531f
C97 source.n14 a_n1712_n3888# 0.493417f
C98 source.t1 a_n1712_n3888# 0.317251f
C99 source.t19 a_n1712_n3888# 0.317251f
C100 source.n15 a_n1712_n3888# 2.78678f
C101 source.n16 a_n1712_n3888# 0.396716f
C102 source.t3 a_n1712_n3888# 0.317251f
C103 source.t5 a_n1712_n3888# 0.317251f
C104 source.n17 a_n1712_n3888# 2.78678f
C105 source.n18 a_n1712_n3888# 0.387051f
C106 source.t2 a_n1712_n3888# 3.55531f
C107 source.n19 a_n1712_n3888# 0.625466f
C108 source.n20 a_n1712_n3888# 1.96579f
C109 drain_left.t9 a_n1712_n3888# 3.57281f
C110 drain_left.t8 a_n1712_n3888# 0.309316f
C111 drain_left.t0 a_n1712_n3888# 0.309316f
C112 drain_left.n0 a_n1712_n3888# 2.79585f
C113 drain_left.n1 a_n1712_n3888# 0.640224f
C114 drain_left.t7 a_n1712_n3888# 0.309316f
C115 drain_left.t4 a_n1712_n3888# 0.309316f
C116 drain_left.n2 a_n1712_n3888# 2.79841f
C117 drain_left.n3 a_n1712_n3888# 1.76147f
C118 drain_left.t3 a_n1712_n3888# 3.57281f
C119 drain_left.t1 a_n1712_n3888# 0.309316f
C120 drain_left.t5 a_n1712_n3888# 0.309316f
C121 drain_left.n4 a_n1712_n3888# 2.79585f
C122 drain_left.n5 a_n1712_n3888# 0.685098f
C123 drain_left.t2 a_n1712_n3888# 0.309316f
C124 drain_left.t6 a_n1712_n3888# 0.309316f
C125 drain_left.n6 a_n1712_n3888# 2.79584f
C126 drain_left.n7 a_n1712_n3888# 0.55826f
C127 plus.n0 a_n1712_n3888# 0.048096f
C128 plus.t8 a_n1712_n3888# 1.02506f
C129 plus.t5 a_n1712_n3888# 1.02506f
C130 plus.t9 a_n1712_n3888# 1.02506f
C131 plus.n1 a_n1712_n3888# 0.404367f
C132 plus.t2 a_n1712_n3888# 1.03525f
C133 plus.n2 a_n1712_n3888# 0.38949f
C134 plus.t7 a_n1712_n3888# 1.02506f
C135 plus.n3 a_n1712_n3888# 0.401699f
C136 plus.n4 a_n1712_n3888# 0.010914f
C137 plus.n5 a_n1712_n3888# 0.153425f
C138 plus.n6 a_n1712_n3888# 0.048096f
C139 plus.n7 a_n1712_n3888# 0.048096f
C140 plus.n8 a_n1712_n3888# 0.010914f
C141 plus.n9 a_n1712_n3888# 0.401699f
C142 plus.n10 a_n1712_n3888# 0.399326f
C143 plus.n11 a_n1712_n3888# 0.614909f
C144 plus.n12 a_n1712_n3888# 0.048096f
C145 plus.t4 a_n1712_n3888# 1.02506f
C146 plus.t3 a_n1712_n3888# 1.02506f
C147 plus.t6 a_n1712_n3888# 1.02506f
C148 plus.n13 a_n1712_n3888# 0.404367f
C149 plus.t1 a_n1712_n3888# 1.03525f
C150 plus.n14 a_n1712_n3888# 0.38949f
C151 plus.t0 a_n1712_n3888# 1.02506f
C152 plus.n15 a_n1712_n3888# 0.401699f
C153 plus.n16 a_n1712_n3888# 0.010914f
C154 plus.n17 a_n1712_n3888# 0.153425f
C155 plus.n18 a_n1712_n3888# 0.048096f
C156 plus.n19 a_n1712_n3888# 0.048096f
C157 plus.n20 a_n1712_n3888# 0.010914f
C158 plus.n21 a_n1712_n3888# 0.401699f
C159 plus.n22 a_n1712_n3888# 0.399326f
C160 plus.n23 a_n1712_n3888# 1.5052f
.ends

