* NGSPICE file created from diffpair225.ext - technology: sky130A

.subckt diffpair225 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t11 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 source.t9 minus.t1 drain_right.t10 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 source.t23 plus.t0 drain_left.t11 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X3 source.t15 minus.t2 drain_right.t9 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X4 source.t5 plus.t1 drain_left.t10 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 source.t3 plus.t2 drain_left.t9 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X6 drain_right.t8 minus.t3 source.t8 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X7 source.t16 minus.t4 drain_right.t7 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X8 source.t12 minus.t5 drain_right.t6 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X9 drain_left.t8 plus.t3 source.t20 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X10 source.t21 plus.t4 drain_left.t7 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X11 a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X12 drain_right.t5 minus.t6 source.t18 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X13 drain_right.t4 minus.t7 source.t14 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X14 drain_left.t6 plus.t5 source.t7 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X15 drain_right.t3 minus.t8 source.t13 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 drain_left.t5 plus.t6 source.t1 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X17 drain_left.t4 plus.t7 source.t22 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X18 a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X19 drain_right.t2 minus.t9 source.t17 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X20 drain_left.t3 plus.t8 source.t4 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X21 drain_left.t2 plus.t9 source.t2 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X22 source.t0 plus.t10 drain_left.t1 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X24 source.t10 minus.t10 drain_right.t1 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X25 source.t19 minus.t11 drain_right.t0 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X26 a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X27 source.t6 plus.t11 drain_left.t0 a_n2158_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n5 minus.t9 182.708
R1 minus.n23 minus.t1 182.708
R2 minus.n17 minus.n16 161.3
R3 minus.n15 minus.n0 161.3
R4 minus.n14 minus.n13 161.3
R5 minus.n12 minus.n1 161.3
R6 minus.n11 minus.n10 161.3
R7 minus.n9 minus.n2 161.3
R8 minus.n8 minus.n7 161.3
R9 minus.n6 minus.n3 161.3
R10 minus.n35 minus.n34 161.3
R11 minus.n33 minus.n18 161.3
R12 minus.n32 minus.n31 161.3
R13 minus.n30 minus.n19 161.3
R14 minus.n29 minus.n28 161.3
R15 minus.n27 minus.n20 161.3
R16 minus.n26 minus.n25 161.3
R17 minus.n24 minus.n21 161.3
R18 minus.n4 minus.t2 159.405
R19 minus.n8 minus.t8 159.405
R20 minus.n10 minus.t10 159.405
R21 minus.n14 minus.t6 159.405
R22 minus.n16 minus.t11 159.405
R23 minus.n22 minus.t0 159.405
R24 minus.n26 minus.t4 159.405
R25 minus.n28 minus.t3 159.405
R26 minus.n32 minus.t5 159.405
R27 minus.n34 minus.t7 159.405
R28 minus.n6 minus.n5 44.8907
R29 minus.n24 minus.n23 44.8907
R30 minus.n16 minus.n15 32.8641
R31 minus.n34 minus.n33 32.8641
R32 minus.n36 minus.n17 30.6217
R33 minus.n4 minus.n3 28.4823
R34 minus.n14 minus.n1 28.4823
R35 minus.n22 minus.n21 28.4823
R36 minus.n32 minus.n19 28.4823
R37 minus.n10 minus.n9 24.1005
R38 minus.n9 minus.n8 24.1005
R39 minus.n27 minus.n26 24.1005
R40 minus.n28 minus.n27 24.1005
R41 minus.n8 minus.n3 19.7187
R42 minus.n10 minus.n1 19.7187
R43 minus.n26 minus.n21 19.7187
R44 minus.n28 minus.n19 19.7187
R45 minus.n5 minus.n4 18.4104
R46 minus.n23 minus.n22 18.4104
R47 minus.n15 minus.n14 15.3369
R48 minus.n33 minus.n32 15.3369
R49 minus.n36 minus.n35 6.64444
R50 minus.n17 minus.n0 0.189894
R51 minus.n13 minus.n0 0.189894
R52 minus.n13 minus.n12 0.189894
R53 minus.n12 minus.n11 0.189894
R54 minus.n11 minus.n2 0.189894
R55 minus.n7 minus.n2 0.189894
R56 minus.n7 minus.n6 0.189894
R57 minus.n25 minus.n24 0.189894
R58 minus.n25 minus.n20 0.189894
R59 minus.n29 minus.n20 0.189894
R60 minus.n30 minus.n29 0.189894
R61 minus.n31 minus.n30 0.189894
R62 minus.n31 minus.n18 0.189894
R63 minus.n35 minus.n18 0.189894
R64 minus minus.n36 0.188
R65 source.n0 source.t22 69.6943
R66 source.n5 source.t3 69.6943
R67 source.n6 source.t17 69.6943
R68 source.n11 source.t19 69.6943
R69 source.n23 source.t14 69.6942
R70 source.n18 source.t9 69.6942
R71 source.n17 source.t20 69.6942
R72 source.n12 source.t6 69.6942
R73 source.n2 source.n1 63.0943
R74 source.n4 source.n3 63.0943
R75 source.n8 source.n7 63.0943
R76 source.n10 source.n9 63.0943
R77 source.n22 source.n21 63.0942
R78 source.n20 source.n19 63.0942
R79 source.n16 source.n15 63.0942
R80 source.n14 source.n13 63.0942
R81 source.n12 source.n11 15.3575
R82 source.n24 source.n0 9.65058
R83 source.n21 source.t8 6.6005
R84 source.n21 source.t12 6.6005
R85 source.n19 source.t11 6.6005
R86 source.n19 source.t16 6.6005
R87 source.n15 source.t7 6.6005
R88 source.n15 source.t21 6.6005
R89 source.n13 source.t2 6.6005
R90 source.n13 source.t0 6.6005
R91 source.n1 source.t1 6.6005
R92 source.n1 source.t5 6.6005
R93 source.n3 source.t4 6.6005
R94 source.n3 source.t23 6.6005
R95 source.n7 source.t13 6.6005
R96 source.n7 source.t15 6.6005
R97 source.n9 source.t18 6.6005
R98 source.n9 source.t10 6.6005
R99 source.n24 source.n23 5.7074
R100 source.n11 source.n10 0.888431
R101 source.n10 source.n8 0.888431
R102 source.n8 source.n6 0.888431
R103 source.n5 source.n4 0.888431
R104 source.n4 source.n2 0.888431
R105 source.n2 source.n0 0.888431
R106 source.n14 source.n12 0.888431
R107 source.n16 source.n14 0.888431
R108 source.n17 source.n16 0.888431
R109 source.n20 source.n18 0.888431
R110 source.n22 source.n20 0.888431
R111 source.n23 source.n22 0.888431
R112 source.n6 source.n5 0.470328
R113 source.n18 source.n17 0.470328
R114 source source.n24 0.188
R115 drain_right.n6 drain_right.n4 80.661
R116 drain_right.n3 drain_right.n2 80.6056
R117 drain_right.n3 drain_right.n0 80.6056
R118 drain_right.n6 drain_right.n5 79.7731
R119 drain_right.n8 drain_right.n7 79.7731
R120 drain_right.n3 drain_right.n1 79.773
R121 drain_right drain_right.n3 24.4353
R122 drain_right.n1 drain_right.t7 6.6005
R123 drain_right.n1 drain_right.t8 6.6005
R124 drain_right.n2 drain_right.t6 6.6005
R125 drain_right.n2 drain_right.t4 6.6005
R126 drain_right.n0 drain_right.t10 6.6005
R127 drain_right.n0 drain_right.t11 6.6005
R128 drain_right.n4 drain_right.t9 6.6005
R129 drain_right.n4 drain_right.t2 6.6005
R130 drain_right.n5 drain_right.t1 6.6005
R131 drain_right.n5 drain_right.t3 6.6005
R132 drain_right.n7 drain_right.t0 6.6005
R133 drain_right.n7 drain_right.t5 6.6005
R134 drain_right drain_right.n8 6.54115
R135 drain_right.n8 drain_right.n6 0.888431
R136 plus.n5 plus.t2 182.708
R137 plus.n23 plus.t3 182.708
R138 plus.n7 plus.n6 161.3
R139 plus.n8 plus.n3 161.3
R140 plus.n10 plus.n9 161.3
R141 plus.n11 plus.n2 161.3
R142 plus.n13 plus.n12 161.3
R143 plus.n14 plus.n1 161.3
R144 plus.n15 plus.n0 161.3
R145 plus.n17 plus.n16 161.3
R146 plus.n25 plus.n24 161.3
R147 plus.n26 plus.n21 161.3
R148 plus.n28 plus.n27 161.3
R149 plus.n29 plus.n20 161.3
R150 plus.n31 plus.n30 161.3
R151 plus.n32 plus.n19 161.3
R152 plus.n33 plus.n18 161.3
R153 plus.n35 plus.n34 161.3
R154 plus.n16 plus.t7 159.405
R155 plus.n14 plus.t1 159.405
R156 plus.n2 plus.t6 159.405
R157 plus.n8 plus.t0 159.405
R158 plus.n4 plus.t8 159.405
R159 plus.n34 plus.t11 159.405
R160 plus.n32 plus.t9 159.405
R161 plus.n20 plus.t10 159.405
R162 plus.n26 plus.t5 159.405
R163 plus.n22 plus.t4 159.405
R164 plus.n6 plus.n5 44.8907
R165 plus.n24 plus.n23 44.8907
R166 plus.n16 plus.n15 32.8641
R167 plus.n34 plus.n33 32.8641
R168 plus.n14 plus.n13 28.4823
R169 plus.n7 plus.n4 28.4823
R170 plus.n32 plus.n31 28.4823
R171 plus.n25 plus.n22 28.4823
R172 plus plus.n35 27.9119
R173 plus.n9 plus.n8 24.1005
R174 plus.n9 plus.n2 24.1005
R175 plus.n27 plus.n20 24.1005
R176 plus.n27 plus.n26 24.1005
R177 plus.n13 plus.n2 19.7187
R178 plus.n8 plus.n7 19.7187
R179 plus.n31 plus.n20 19.7187
R180 plus.n26 plus.n25 19.7187
R181 plus.n5 plus.n4 18.4104
R182 plus.n23 plus.n22 18.4104
R183 plus.n15 plus.n14 15.3369
R184 plus.n33 plus.n32 15.3369
R185 plus plus.n17 8.87929
R186 plus.n6 plus.n3 0.189894
R187 plus.n10 plus.n3 0.189894
R188 plus.n11 plus.n10 0.189894
R189 plus.n12 plus.n11 0.189894
R190 plus.n12 plus.n1 0.189894
R191 plus.n1 plus.n0 0.189894
R192 plus.n17 plus.n0 0.189894
R193 plus.n35 plus.n18 0.189894
R194 plus.n19 plus.n18 0.189894
R195 plus.n30 plus.n19 0.189894
R196 plus.n30 plus.n29 0.189894
R197 plus.n29 plus.n28 0.189894
R198 plus.n28 plus.n21 0.189894
R199 plus.n24 plus.n21 0.189894
R200 drain_left.n6 drain_left.n4 80.661
R201 drain_left.n3 drain_left.n2 80.6056
R202 drain_left.n3 drain_left.n0 80.6056
R203 drain_left.n8 drain_left.n7 79.7731
R204 drain_left.n6 drain_left.n5 79.7731
R205 drain_left.n3 drain_left.n1 79.773
R206 drain_left drain_left.n3 24.9885
R207 drain_left.n1 drain_left.t1 6.6005
R208 drain_left.n1 drain_left.t6 6.6005
R209 drain_left.n2 drain_left.t7 6.6005
R210 drain_left.n2 drain_left.t8 6.6005
R211 drain_left.n0 drain_left.t0 6.6005
R212 drain_left.n0 drain_left.t2 6.6005
R213 drain_left.n7 drain_left.t10 6.6005
R214 drain_left.n7 drain_left.t4 6.6005
R215 drain_left.n5 drain_left.t11 6.6005
R216 drain_left.n5 drain_left.t5 6.6005
R217 drain_left.n4 drain_left.t9 6.6005
R218 drain_left.n4 drain_left.t3 6.6005
R219 drain_left drain_left.n8 6.54115
R220 drain_left.n8 drain_left.n6 0.888431
C0 source drain_right 5.98712f
C1 minus plus 4.17472f
C2 drain_left drain_right 1.08493f
C3 source plus 2.71727f
C4 drain_left plus 2.55651f
C5 minus source 2.70327f
C6 minus drain_left 0.176812f
C7 drain_right plus 0.372332f
C8 minus drain_right 2.34481f
C9 source drain_left 5.98508f
C10 drain_right a_n2158_n1488# 4.42299f
C11 drain_left a_n2158_n1488# 4.7632f
C12 source a_n2158_n1488# 3.805873f
C13 minus a_n2158_n1488# 7.772424f
C14 plus a_n2158_n1488# 9.05417f
C15 drain_left.t0 a_n2158_n1488# 0.063962f
C16 drain_left.t2 a_n2158_n1488# 0.063962f
C17 drain_left.n0 a_n2158_n1488# 0.465186f
C18 drain_left.t1 a_n2158_n1488# 0.063962f
C19 drain_left.t6 a_n2158_n1488# 0.063962f
C20 drain_left.n1 a_n2158_n1488# 0.46129f
C21 drain_left.t7 a_n2158_n1488# 0.063962f
C22 drain_left.t8 a_n2158_n1488# 0.063962f
C23 drain_left.n2 a_n2158_n1488# 0.465186f
C24 drain_left.n3 a_n2158_n1488# 1.96708f
C25 drain_left.t9 a_n2158_n1488# 0.063962f
C26 drain_left.t3 a_n2158_n1488# 0.063962f
C27 drain_left.n4 a_n2158_n1488# 0.465489f
C28 drain_left.t11 a_n2158_n1488# 0.063962f
C29 drain_left.t5 a_n2158_n1488# 0.063962f
C30 drain_left.n5 a_n2158_n1488# 0.461292f
C31 drain_left.n6 a_n2158_n1488# 0.747391f
C32 drain_left.t10 a_n2158_n1488# 0.063962f
C33 drain_left.t4 a_n2158_n1488# 0.063962f
C34 drain_left.n7 a_n2158_n1488# 0.461292f
C35 drain_left.n8 a_n2158_n1488# 0.609004f
C36 plus.n0 a_n2158_n1488# 0.045702f
C37 plus.t7 a_n2158_n1488# 0.287795f
C38 plus.t1 a_n2158_n1488# 0.287795f
C39 plus.n1 a_n2158_n1488# 0.045702f
C40 plus.t6 a_n2158_n1488# 0.287795f
C41 plus.n2 a_n2158_n1488# 0.167618f
C42 plus.n3 a_n2158_n1488# 0.045702f
C43 plus.t0 a_n2158_n1488# 0.287795f
C44 plus.t8 a_n2158_n1488# 0.287795f
C45 plus.n4 a_n2158_n1488# 0.17273f
C46 plus.t2 a_n2158_n1488# 0.309166f
C47 plus.n5 a_n2158_n1488# 0.150338f
C48 plus.n6 a_n2158_n1488# 0.191727f
C49 plus.n7 a_n2158_n1488# 0.010371f
C50 plus.n8 a_n2158_n1488# 0.167618f
C51 plus.n9 a_n2158_n1488# 0.010371f
C52 plus.n10 a_n2158_n1488# 0.045702f
C53 plus.n11 a_n2158_n1488# 0.045702f
C54 plus.n12 a_n2158_n1488# 0.045702f
C55 plus.n13 a_n2158_n1488# 0.010371f
C56 plus.n14 a_n2158_n1488# 0.167618f
C57 plus.n15 a_n2158_n1488# 0.010371f
C58 plus.n16 a_n2158_n1488# 0.165505f
C59 plus.n17 a_n2158_n1488# 0.357667f
C60 plus.n18 a_n2158_n1488# 0.045702f
C61 plus.t11 a_n2158_n1488# 0.287795f
C62 plus.n19 a_n2158_n1488# 0.045702f
C63 plus.t9 a_n2158_n1488# 0.287795f
C64 plus.t10 a_n2158_n1488# 0.287795f
C65 plus.n20 a_n2158_n1488# 0.167618f
C66 plus.n21 a_n2158_n1488# 0.045702f
C67 plus.t5 a_n2158_n1488# 0.287795f
C68 plus.t4 a_n2158_n1488# 0.287795f
C69 plus.n22 a_n2158_n1488# 0.17273f
C70 plus.t3 a_n2158_n1488# 0.309166f
C71 plus.n23 a_n2158_n1488# 0.150338f
C72 plus.n24 a_n2158_n1488# 0.191727f
C73 plus.n25 a_n2158_n1488# 0.010371f
C74 plus.n26 a_n2158_n1488# 0.167618f
C75 plus.n27 a_n2158_n1488# 0.010371f
C76 plus.n28 a_n2158_n1488# 0.045702f
C77 plus.n29 a_n2158_n1488# 0.045702f
C78 plus.n30 a_n2158_n1488# 0.045702f
C79 plus.n31 a_n2158_n1488# 0.010371f
C80 plus.n32 a_n2158_n1488# 0.167618f
C81 plus.n33 a_n2158_n1488# 0.010371f
C82 plus.n34 a_n2158_n1488# 0.165505f
C83 plus.n35 a_n2158_n1488# 1.16268f
C84 drain_right.t10 a_n2158_n1488# 0.062498f
C85 drain_right.t11 a_n2158_n1488# 0.062498f
C86 drain_right.n0 a_n2158_n1488# 0.454536f
C87 drain_right.t7 a_n2158_n1488# 0.062498f
C88 drain_right.t8 a_n2158_n1488# 0.062498f
C89 drain_right.n1 a_n2158_n1488# 0.45073f
C90 drain_right.t6 a_n2158_n1488# 0.062498f
C91 drain_right.t4 a_n2158_n1488# 0.062498f
C92 drain_right.n2 a_n2158_n1488# 0.454536f
C93 drain_right.n3 a_n2158_n1488# 1.87001f
C94 drain_right.t9 a_n2158_n1488# 0.062498f
C95 drain_right.t2 a_n2158_n1488# 0.062498f
C96 drain_right.n4 a_n2158_n1488# 0.454833f
C97 drain_right.t1 a_n2158_n1488# 0.062498f
C98 drain_right.t3 a_n2158_n1488# 0.062498f
C99 drain_right.n5 a_n2158_n1488# 0.450732f
C100 drain_right.n6 a_n2158_n1488# 0.730282f
C101 drain_right.t0 a_n2158_n1488# 0.062498f
C102 drain_right.t5 a_n2158_n1488# 0.062498f
C103 drain_right.n7 a_n2158_n1488# 0.450732f
C104 drain_right.n8 a_n2158_n1488# 0.595063f
C105 source.t22 a_n2158_n1488# 0.526052f
C106 source.n0 a_n2158_n1488# 0.769866f
C107 source.t1 a_n2158_n1488# 0.063351f
C108 source.t5 a_n2158_n1488# 0.063351f
C109 source.n1 a_n2158_n1488# 0.401679f
C110 source.n2 a_n2158_n1488# 0.385699f
C111 source.t4 a_n2158_n1488# 0.063351f
C112 source.t23 a_n2158_n1488# 0.063351f
C113 source.n3 a_n2158_n1488# 0.401679f
C114 source.n4 a_n2158_n1488# 0.385699f
C115 source.t3 a_n2158_n1488# 0.526052f
C116 source.n5 a_n2158_n1488# 0.398099f
C117 source.t17 a_n2158_n1488# 0.526052f
C118 source.n6 a_n2158_n1488# 0.398099f
C119 source.t13 a_n2158_n1488# 0.063351f
C120 source.t15 a_n2158_n1488# 0.063351f
C121 source.n7 a_n2158_n1488# 0.401679f
C122 source.n8 a_n2158_n1488# 0.385699f
C123 source.t18 a_n2158_n1488# 0.063351f
C124 source.t10 a_n2158_n1488# 0.063351f
C125 source.n9 a_n2158_n1488# 0.401679f
C126 source.n10 a_n2158_n1488# 0.385699f
C127 source.t19 a_n2158_n1488# 0.526052f
C128 source.n11 a_n2158_n1488# 1.05564f
C129 source.t6 a_n2158_n1488# 0.52605f
C130 source.n12 a_n2158_n1488# 1.05564f
C131 source.t2 a_n2158_n1488# 0.063351f
C132 source.t0 a_n2158_n1488# 0.063351f
C133 source.n13 a_n2158_n1488# 0.401676f
C134 source.n14 a_n2158_n1488# 0.385701f
C135 source.t7 a_n2158_n1488# 0.063351f
C136 source.t21 a_n2158_n1488# 0.063351f
C137 source.n15 a_n2158_n1488# 0.401676f
C138 source.n16 a_n2158_n1488# 0.385701f
C139 source.t20 a_n2158_n1488# 0.52605f
C140 source.n17 a_n2158_n1488# 0.398102f
C141 source.t9 a_n2158_n1488# 0.52605f
C142 source.n18 a_n2158_n1488# 0.398102f
C143 source.t11 a_n2158_n1488# 0.063351f
C144 source.t16 a_n2158_n1488# 0.063351f
C145 source.n19 a_n2158_n1488# 0.401676f
C146 source.n20 a_n2158_n1488# 0.385701f
C147 source.t8 a_n2158_n1488# 0.063351f
C148 source.t12 a_n2158_n1488# 0.063351f
C149 source.n21 a_n2158_n1488# 0.401676f
C150 source.n22 a_n2158_n1488# 0.385701f
C151 source.t14 a_n2158_n1488# 0.52605f
C152 source.n23 a_n2158_n1488# 0.572413f
C153 source.n24 a_n2158_n1488# 0.788011f
C154 minus.n0 a_n2158_n1488# 0.043833f
C155 minus.n1 a_n2158_n1488# 0.009947f
C156 minus.t6 a_n2158_n1488# 0.276021f
C157 minus.n2 a_n2158_n1488# 0.043833f
C158 minus.n3 a_n2158_n1488# 0.009947f
C159 minus.t8 a_n2158_n1488# 0.276021f
C160 minus.t9 a_n2158_n1488# 0.296518f
C161 minus.t2 a_n2158_n1488# 0.276021f
C162 minus.n4 a_n2158_n1488# 0.165664f
C163 minus.n5 a_n2158_n1488# 0.144188f
C164 minus.n6 a_n2158_n1488# 0.183883f
C165 minus.n7 a_n2158_n1488# 0.043833f
C166 minus.n8 a_n2158_n1488# 0.160761f
C167 minus.n9 a_n2158_n1488# 0.009947f
C168 minus.t10 a_n2158_n1488# 0.276021f
C169 minus.n10 a_n2158_n1488# 0.160761f
C170 minus.n11 a_n2158_n1488# 0.043833f
C171 minus.n12 a_n2158_n1488# 0.043833f
C172 minus.n13 a_n2158_n1488# 0.043833f
C173 minus.n14 a_n2158_n1488# 0.160761f
C174 minus.n15 a_n2158_n1488# 0.009947f
C175 minus.t11 a_n2158_n1488# 0.276021f
C176 minus.n16 a_n2158_n1488# 0.158734f
C177 minus.n17 a_n2158_n1488# 1.18648f
C178 minus.n18 a_n2158_n1488# 0.043833f
C179 minus.n19 a_n2158_n1488# 0.009947f
C180 minus.n20 a_n2158_n1488# 0.043833f
C181 minus.n21 a_n2158_n1488# 0.009947f
C182 minus.t1 a_n2158_n1488# 0.296518f
C183 minus.t0 a_n2158_n1488# 0.276021f
C184 minus.n22 a_n2158_n1488# 0.165664f
C185 minus.n23 a_n2158_n1488# 0.144188f
C186 minus.n24 a_n2158_n1488# 0.183883f
C187 minus.n25 a_n2158_n1488# 0.043833f
C188 minus.t4 a_n2158_n1488# 0.276021f
C189 minus.n26 a_n2158_n1488# 0.160761f
C190 minus.n27 a_n2158_n1488# 0.009947f
C191 minus.t3 a_n2158_n1488# 0.276021f
C192 minus.n28 a_n2158_n1488# 0.160761f
C193 minus.n29 a_n2158_n1488# 0.043833f
C194 minus.n30 a_n2158_n1488# 0.043833f
C195 minus.n31 a_n2158_n1488# 0.043833f
C196 minus.t5 a_n2158_n1488# 0.276021f
C197 minus.n32 a_n2158_n1488# 0.160761f
C198 minus.n33 a_n2158_n1488# 0.009947f
C199 minus.t7 a_n2158_n1488# 0.276021f
C200 minus.n34 a_n2158_n1488# 0.158734f
C201 minus.n35 a_n2158_n1488# 0.301382f
C202 minus.n36 a_n2158_n1488# 1.45504f
.ends

