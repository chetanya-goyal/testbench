* NGSPICE file created from diffpair408.ext - technology: sky130A

.subckt diffpair408 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t30 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X1 source.t37 minus.t1 drain_right.t18 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X2 a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X3 source.t2 plus.t0 drain_left.t19 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X4 a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X5 drain_left.t18 plus.t1 source.t9 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X6 source.t1 plus.t2 drain_left.t17 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X7 drain_left.t16 plus.t3 source.t5 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X8 a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X9 source.t12 plus.t4 drain_left.t15 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X10 drain_left.t14 plus.t5 source.t16 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X11 source.t21 minus.t2 drain_right.t17 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X12 source.t24 minus.t3 drain_right.t16 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 drain_left.t13 plus.t6 source.t11 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X14 source.t27 minus.t4 drain_right.t15 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X15 a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X16 drain_left.t12 plus.t7 source.t10 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 drain_right.t14 minus.t5 source.t33 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X18 drain_right.t13 minus.t6 source.t22 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 drain_right.t12 minus.t7 source.t25 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X20 source.t18 minus.t8 drain_right.t11 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X21 drain_right.t10 minus.t9 source.t31 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X22 drain_right.t9 minus.t10 source.t28 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X23 drain_right.t8 minus.t11 source.t35 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X24 source.t38 plus.t8 drain_left.t11 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X25 drain_left.t10 plus.t9 source.t39 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X26 source.t4 plus.t10 drain_left.t9 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X27 drain_right.t7 minus.t12 source.t34 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X28 drain_right.t6 minus.t13 source.t23 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X29 source.t26 minus.t14 drain_right.t5 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X30 drain_left.t8 plus.t11 source.t0 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X31 source.t20 minus.t15 drain_right.t4 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X32 source.t19 minus.t16 drain_right.t3 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X33 drain_left.t7 plus.t12 source.t3 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X34 source.t17 plus.t13 drain_left.t6 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X35 source.t15 plus.t14 drain_left.t5 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X36 source.t32 minus.t17 drain_right.t2 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X37 source.t29 minus.t18 drain_right.t1 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X38 source.t7 plus.t15 drain_left.t4 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X39 drain_left.t3 plus.t16 source.t13 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X40 drain_left.t2 plus.t17 source.t14 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X41 source.t6 plus.t18 drain_left.t1 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X42 drain_right.t0 minus.t19 source.t36 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X43 source.t8 plus.t19 drain_left.t0 a_n2146_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
R0 minus.n27 minus.t18 2198.94
R1 minus.n7 minus.t5 2198.94
R2 minus.n56 minus.t11 2198.94
R3 minus.n35 minus.t1 2198.94
R4 minus.n26 minus.t10 2136.87
R5 minus.n24 minus.t14 2136.87
R6 minus.n3 minus.t13 2136.87
R7 minus.n18 minus.t15 2136.87
R8 minus.n16 minus.t6 2136.87
R9 minus.n4 minus.t8 2136.87
R10 minus.n10 minus.t12 2136.87
R11 minus.n6 minus.t4 2136.87
R12 minus.n55 minus.t3 2136.87
R13 minus.n53 minus.t0 2136.87
R14 minus.n47 minus.t17 2136.87
R15 minus.n46 minus.t9 2136.87
R16 minus.n44 minus.t2 2136.87
R17 minus.n32 minus.t19 2136.87
R18 minus.n38 minus.t16 2136.87
R19 minus.n34 minus.t7 2136.87
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 69.3793
R47 minus.n15 minus.n4 69.3793
R48 minus.n43 minus.n32 69.3793
R49 minus.n48 minus.n47 69.3793
R50 minus.n25 minus.n24 54.7732
R51 minus.n10 minus.n9 54.7732
R52 minus.n38 minus.n37 54.7732
R53 minus.n54 minus.n53 54.7732
R54 minus.n18 minus.n17 47.4702
R55 minus.n17 minus.n16 47.4702
R56 minus.n45 minus.n44 47.4702
R57 minus.n46 minus.n45 47.4702
R58 minus.n26 minus.n25 40.1672
R59 minus.n9 minus.n6 40.1672
R60 minus.n37 minus.n34 40.1672
R61 minus.n55 minus.n54 40.1672
R62 minus.n58 minus.n28 37.3111
R63 minus.n27 minus.n26 32.8641
R64 minus.n7 minus.n6 32.8641
R65 minus.n35 minus.n34 32.8641
R66 minus.n56 minus.n55 32.8641
R67 minus.n19 minus.n18 25.5611
R68 minus.n16 minus.n15 25.5611
R69 minus.n44 minus.n43 25.5611
R70 minus.n48 minus.n46 25.5611
R71 minus.n24 minus.n23 18.2581
R72 minus.n11 minus.n10 18.2581
R73 minus.n39 minus.n38 18.2581
R74 minus.n53 minus.n52 18.2581
R75 minus.n58 minus.n57 6.56111
R76 minus.n3 minus.n1 3.65202
R77 minus.n12 minus.n4 3.65202
R78 minus.n40 minus.n32 3.65202
R79 minus.n47 minus.n30 3.65202
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 source.n9 source.t4 45.3739
R100 source.n10 source.t33 45.3739
R101 source.n19 source.t29 45.3739
R102 source.n39 source.t35 45.3737
R103 source.n30 source.t37 45.3737
R104 source.n29 source.t11 45.3737
R105 source.n20 source.t8 45.3737
R106 source.n0 source.t3 45.3737
R107 source.n2 source.n1 42.8739
R108 source.n4 source.n3 42.8739
R109 source.n6 source.n5 42.8739
R110 source.n8 source.n7 42.8739
R111 source.n12 source.n11 42.8739
R112 source.n14 source.n13 42.8739
R113 source.n16 source.n15 42.8739
R114 source.n18 source.n17 42.8739
R115 source.n38 source.n37 42.8737
R116 source.n36 source.n35 42.8737
R117 source.n34 source.n33 42.8737
R118 source.n32 source.n31 42.8737
R119 source.n28 source.n27 42.8737
R120 source.n26 source.n25 42.8737
R121 source.n24 source.n23 42.8737
R122 source.n22 source.n21 42.8737
R123 source.n20 source.n19 21.8481
R124 source.n40 source.n0 16.305
R125 source.n40 source.n39 5.5436
R126 source.n37 source.t30 2.5005
R127 source.n37 source.t24 2.5005
R128 source.n35 source.t31 2.5005
R129 source.n35 source.t32 2.5005
R130 source.n33 source.t36 2.5005
R131 source.n33 source.t21 2.5005
R132 source.n31 source.t25 2.5005
R133 source.n31 source.t19 2.5005
R134 source.n27 source.t9 2.5005
R135 source.n27 source.t38 2.5005
R136 source.n25 source.t10 2.5005
R137 source.n25 source.t12 2.5005
R138 source.n23 source.t5 2.5005
R139 source.n23 source.t2 2.5005
R140 source.n21 source.t16 2.5005
R141 source.n21 source.t1 2.5005
R142 source.n1 source.t39 2.5005
R143 source.n1 source.t7 2.5005
R144 source.n3 source.t13 2.5005
R145 source.n3 source.t17 2.5005
R146 source.n5 source.t0 2.5005
R147 source.n5 source.t6 2.5005
R148 source.n7 source.t14 2.5005
R149 source.n7 source.t15 2.5005
R150 source.n11 source.t34 2.5005
R151 source.n11 source.t27 2.5005
R152 source.n13 source.t22 2.5005
R153 source.n13 source.t18 2.5005
R154 source.n15 source.t23 2.5005
R155 source.n15 source.t20 2.5005
R156 source.n17 source.t28 2.5005
R157 source.n17 source.t26 2.5005
R158 source.n19 source.n18 0.560845
R159 source.n18 source.n16 0.560845
R160 source.n16 source.n14 0.560845
R161 source.n14 source.n12 0.560845
R162 source.n12 source.n10 0.560845
R163 source.n9 source.n8 0.560845
R164 source.n8 source.n6 0.560845
R165 source.n6 source.n4 0.560845
R166 source.n4 source.n2 0.560845
R167 source.n2 source.n0 0.560845
R168 source.n22 source.n20 0.560845
R169 source.n24 source.n22 0.560845
R170 source.n26 source.n24 0.560845
R171 source.n28 source.n26 0.560845
R172 source.n29 source.n28 0.560845
R173 source.n32 source.n30 0.560845
R174 source.n34 source.n32 0.560845
R175 source.n36 source.n34 0.560845
R176 source.n38 source.n36 0.560845
R177 source.n39 source.n38 0.560845
R178 source.n10 source.n9 0.470328
R179 source.n30 source.n29 0.470328
R180 source source.n40 0.188
R181 drain_right.n6 drain_right.n4 60.1128
R182 drain_right.n2 drain_right.n0 60.1128
R183 drain_right.n10 drain_right.n8 60.1128
R184 drain_right.n10 drain_right.n9 59.5527
R185 drain_right.n12 drain_right.n11 59.5527
R186 drain_right.n14 drain_right.n13 59.5527
R187 drain_right.n16 drain_right.n15 59.5527
R188 drain_right.n7 drain_right.n3 59.5525
R189 drain_right.n6 drain_right.n5 59.5525
R190 drain_right.n2 drain_right.n1 59.5525
R191 drain_right drain_right.n7 31.2966
R192 drain_right drain_right.n16 6.21356
R193 drain_right.n3 drain_right.t17 2.5005
R194 drain_right.n3 drain_right.t10 2.5005
R195 drain_right.n4 drain_right.t16 2.5005
R196 drain_right.n4 drain_right.t8 2.5005
R197 drain_right.n5 drain_right.t2 2.5005
R198 drain_right.n5 drain_right.t19 2.5005
R199 drain_right.n1 drain_right.t3 2.5005
R200 drain_right.n1 drain_right.t0 2.5005
R201 drain_right.n0 drain_right.t18 2.5005
R202 drain_right.n0 drain_right.t12 2.5005
R203 drain_right.n8 drain_right.t15 2.5005
R204 drain_right.n8 drain_right.t14 2.5005
R205 drain_right.n9 drain_right.t11 2.5005
R206 drain_right.n9 drain_right.t7 2.5005
R207 drain_right.n11 drain_right.t4 2.5005
R208 drain_right.n11 drain_right.t13 2.5005
R209 drain_right.n13 drain_right.t5 2.5005
R210 drain_right.n13 drain_right.t6 2.5005
R211 drain_right.n15 drain_right.t1 2.5005
R212 drain_right.n15 drain_right.t9 2.5005
R213 drain_right.n16 drain_right.n14 0.560845
R214 drain_right.n14 drain_right.n12 0.560845
R215 drain_right.n12 drain_right.n10 0.560845
R216 drain_right.n7 drain_right.n6 0.505499
R217 drain_right.n7 drain_right.n2 0.505499
R218 plus.n6 plus.t10 2198.94
R219 plus.n27 plus.t12 2198.94
R220 plus.n36 plus.t6 2198.94
R221 plus.n56 plus.t19 2198.94
R222 plus.n5 plus.t17 2136.87
R223 plus.n9 plus.t14 2136.87
R224 plus.n3 plus.t11 2136.87
R225 plus.n15 plus.t18 2136.87
R226 plus.n17 plus.t16 2136.87
R227 plus.n18 plus.t13 2136.87
R228 plus.n24 plus.t9 2136.87
R229 plus.n26 plus.t15 2136.87
R230 plus.n35 plus.t8 2136.87
R231 plus.n39 plus.t1 2136.87
R232 plus.n33 plus.t4 2136.87
R233 plus.n45 plus.t7 2136.87
R234 plus.n47 plus.t0 2136.87
R235 plus.n32 plus.t3 2136.87
R236 plus.n53 plus.t2 2136.87
R237 plus.n55 plus.t5 2136.87
R238 plus.n7 plus.n6 161.489
R239 plus.n37 plus.n36 161.489
R240 plus.n8 plus.n7 161.3
R241 plus.n10 plus.n4 161.3
R242 plus.n12 plus.n11 161.3
R243 plus.n14 plus.n13 161.3
R244 plus.n16 plus.n2 161.3
R245 plus.n20 plus.n19 161.3
R246 plus.n21 plus.n1 161.3
R247 plus.n23 plus.n22 161.3
R248 plus.n25 plus.n0 161.3
R249 plus.n28 plus.n27 161.3
R250 plus.n38 plus.n37 161.3
R251 plus.n40 plus.n34 161.3
R252 plus.n42 plus.n41 161.3
R253 plus.n44 plus.n43 161.3
R254 plus.n46 plus.n31 161.3
R255 plus.n49 plus.n48 161.3
R256 plus.n50 plus.n30 161.3
R257 plus.n52 plus.n51 161.3
R258 plus.n54 plus.n29 161.3
R259 plus.n57 plus.n56 161.3
R260 plus.n11 plus.n10 73.0308
R261 plus.n23 plus.n1 73.0308
R262 plus.n52 plus.n30 73.0308
R263 plus.n41 plus.n40 73.0308
R264 plus.n14 plus.n3 69.3793
R265 plus.n19 plus.n18 69.3793
R266 plus.n48 plus.n32 69.3793
R267 plus.n44 plus.n33 69.3793
R268 plus.n9 plus.n8 54.7732
R269 plus.n25 plus.n24 54.7732
R270 plus.n54 plus.n53 54.7732
R271 plus.n39 plus.n38 54.7732
R272 plus.n16 plus.n15 47.4702
R273 plus.n17 plus.n16 47.4702
R274 plus.n47 plus.n46 47.4702
R275 plus.n46 plus.n45 47.4702
R276 plus.n8 plus.n5 40.1672
R277 plus.n26 plus.n25 40.1672
R278 plus.n55 plus.n54 40.1672
R279 plus.n38 plus.n35 40.1672
R280 plus.n6 plus.n5 32.8641
R281 plus.n27 plus.n26 32.8641
R282 plus.n56 plus.n55 32.8641
R283 plus.n36 plus.n35 32.8641
R284 plus plus.n57 31.1922
R285 plus.n15 plus.n14 25.5611
R286 plus.n19 plus.n17 25.5611
R287 plus.n48 plus.n47 25.5611
R288 plus.n45 plus.n44 25.5611
R289 plus.n10 plus.n9 18.2581
R290 plus.n24 plus.n23 18.2581
R291 plus.n53 plus.n52 18.2581
R292 plus.n40 plus.n39 18.2581
R293 plus plus.n28 12.205
R294 plus.n11 plus.n3 3.65202
R295 plus.n18 plus.n1 3.65202
R296 plus.n32 plus.n30 3.65202
R297 plus.n41 plus.n33 3.65202
R298 plus.n7 plus.n4 0.189894
R299 plus.n12 plus.n4 0.189894
R300 plus.n13 plus.n12 0.189894
R301 plus.n13 plus.n2 0.189894
R302 plus.n20 plus.n2 0.189894
R303 plus.n21 plus.n20 0.189894
R304 plus.n22 plus.n21 0.189894
R305 plus.n22 plus.n0 0.189894
R306 plus.n28 plus.n0 0.189894
R307 plus.n57 plus.n29 0.189894
R308 plus.n51 plus.n29 0.189894
R309 plus.n51 plus.n50 0.189894
R310 plus.n50 plus.n49 0.189894
R311 plus.n49 plus.n31 0.189894
R312 plus.n43 plus.n31 0.189894
R313 plus.n43 plus.n42 0.189894
R314 plus.n42 plus.n34 0.189894
R315 plus.n37 plus.n34 0.189894
R316 drain_left.n10 drain_left.n8 60.113
R317 drain_left.n6 drain_left.n4 60.1128
R318 drain_left.n2 drain_left.n0 60.1128
R319 drain_left.n14 drain_left.n13 59.5527
R320 drain_left.n12 drain_left.n11 59.5527
R321 drain_left.n10 drain_left.n9 59.5527
R322 drain_left.n7 drain_left.n3 59.5525
R323 drain_left.n6 drain_left.n5 59.5525
R324 drain_left.n2 drain_left.n1 59.5525
R325 drain_left.n16 drain_left.n15 59.5525
R326 drain_left drain_left.n7 31.8498
R327 drain_left drain_left.n16 6.21356
R328 drain_left.n3 drain_left.t19 2.5005
R329 drain_left.n3 drain_left.t12 2.5005
R330 drain_left.n4 drain_left.t11 2.5005
R331 drain_left.n4 drain_left.t13 2.5005
R332 drain_left.n5 drain_left.t15 2.5005
R333 drain_left.n5 drain_left.t18 2.5005
R334 drain_left.n1 drain_left.t17 2.5005
R335 drain_left.n1 drain_left.t16 2.5005
R336 drain_left.n0 drain_left.t0 2.5005
R337 drain_left.n0 drain_left.t14 2.5005
R338 drain_left.n15 drain_left.t4 2.5005
R339 drain_left.n15 drain_left.t7 2.5005
R340 drain_left.n13 drain_left.t6 2.5005
R341 drain_left.n13 drain_left.t10 2.5005
R342 drain_left.n11 drain_left.t1 2.5005
R343 drain_left.n11 drain_left.t3 2.5005
R344 drain_left.n9 drain_left.t5 2.5005
R345 drain_left.n9 drain_left.t8 2.5005
R346 drain_left.n8 drain_left.t9 2.5005
R347 drain_left.n8 drain_left.t2 2.5005
R348 drain_left.n12 drain_left.n10 0.560845
R349 drain_left.n14 drain_left.n12 0.560845
R350 drain_left.n16 drain_left.n14 0.560845
R351 drain_left.n7 drain_left.n6 0.505499
R352 drain_left.n7 drain_left.n2 0.505499
C0 plus source 3.7745f
C1 minus source 3.76046f
C2 drain_left drain_right 1.13563f
C3 drain_right plus 0.364841f
C4 drain_right minus 4.22291f
C5 drain_right source 38.2587f
C6 drain_left plus 4.4336f
C7 drain_left minus 0.171338f
C8 plus minus 5.812871f
C9 drain_left source 38.258198f
C10 drain_right a_n2146_n3288# 6.44799f
C11 drain_left a_n2146_n3288# 6.76243f
C12 source a_n2146_n3288# 8.904922f
C13 minus a_n2146_n3288# 7.927526f
C14 plus a_n2146_n3288# 10.107571f
C15 drain_left.t0 a_n2146_n3288# 0.406191f
C16 drain_left.t14 a_n2146_n3288# 0.406191f
C17 drain_left.n0 a_n2146_n3288# 2.66503f
C18 drain_left.t17 a_n2146_n3288# 0.406191f
C19 drain_left.t16 a_n2146_n3288# 0.406191f
C20 drain_left.n1 a_n2146_n3288# 2.66176f
C21 drain_left.n2 a_n2146_n3288# 0.683082f
C22 drain_left.t19 a_n2146_n3288# 0.406191f
C23 drain_left.t12 a_n2146_n3288# 0.406191f
C24 drain_left.n3 a_n2146_n3288# 2.66176f
C25 drain_left.t11 a_n2146_n3288# 0.406191f
C26 drain_left.t13 a_n2146_n3288# 0.406191f
C27 drain_left.n4 a_n2146_n3288# 2.66503f
C28 drain_left.t15 a_n2146_n3288# 0.406191f
C29 drain_left.t18 a_n2146_n3288# 0.406191f
C30 drain_left.n5 a_n2146_n3288# 2.66176f
C31 drain_left.n6 a_n2146_n3288# 0.683082f
C32 drain_left.n7 a_n2146_n3288# 1.76562f
C33 drain_left.t9 a_n2146_n3288# 0.406191f
C34 drain_left.t2 a_n2146_n3288# 0.406191f
C35 drain_left.n8 a_n2146_n3288# 2.66504f
C36 drain_left.t5 a_n2146_n3288# 0.406191f
C37 drain_left.t8 a_n2146_n3288# 0.406191f
C38 drain_left.n9 a_n2146_n3288# 2.66177f
C39 drain_left.n10 a_n2146_n3288# 0.686806f
C40 drain_left.t1 a_n2146_n3288# 0.406191f
C41 drain_left.t3 a_n2146_n3288# 0.406191f
C42 drain_left.n11 a_n2146_n3288# 2.66177f
C43 drain_left.n12 a_n2146_n3288# 0.339344f
C44 drain_left.t6 a_n2146_n3288# 0.406191f
C45 drain_left.t10 a_n2146_n3288# 0.406191f
C46 drain_left.n13 a_n2146_n3288# 2.66177f
C47 drain_left.n14 a_n2146_n3288# 0.339344f
C48 drain_left.t4 a_n2146_n3288# 0.406191f
C49 drain_left.t7 a_n2146_n3288# 0.406191f
C50 drain_left.n15 a_n2146_n3288# 2.66176f
C51 drain_left.n16 a_n2146_n3288# 0.575446f
C52 plus.n0 a_n2146_n3288# 0.053392f
C53 plus.t15 a_n2146_n3288# 0.271578f
C54 plus.t9 a_n2146_n3288# 0.271578f
C55 plus.n1 a_n2146_n3288# 0.018535f
C56 plus.n2 a_n2146_n3288# 0.053392f
C57 plus.t16 a_n2146_n3288# 0.271578f
C58 plus.t18 a_n2146_n3288# 0.271578f
C59 plus.t11 a_n2146_n3288# 0.271578f
C60 plus.n3 a_n2146_n3288# 0.115963f
C61 plus.n4 a_n2146_n3288# 0.053392f
C62 plus.t14 a_n2146_n3288# 0.271578f
C63 plus.t17 a_n2146_n3288# 0.271578f
C64 plus.n5 a_n2146_n3288# 0.115963f
C65 plus.t10 a_n2146_n3288# 0.274921f
C66 plus.n6 a_n2146_n3288# 0.13782f
C67 plus.n7 a_n2146_n3288# 0.123162f
C68 plus.n8 a_n2146_n3288# 0.02265f
C69 plus.n9 a_n2146_n3288# 0.115963f
C70 plus.n10 a_n2146_n3288# 0.021827f
C71 plus.n11 a_n2146_n3288# 0.018535f
C72 plus.n12 a_n2146_n3288# 0.053392f
C73 plus.n13 a_n2146_n3288# 0.053392f
C74 plus.n14 a_n2146_n3288# 0.02265f
C75 plus.n15 a_n2146_n3288# 0.115963f
C76 plus.n16 a_n2146_n3288# 0.02265f
C77 plus.n17 a_n2146_n3288# 0.115963f
C78 plus.t13 a_n2146_n3288# 0.271578f
C79 plus.n18 a_n2146_n3288# 0.115963f
C80 plus.n19 a_n2146_n3288# 0.02265f
C81 plus.n20 a_n2146_n3288# 0.053392f
C82 plus.n21 a_n2146_n3288# 0.053392f
C83 plus.n22 a_n2146_n3288# 0.053392f
C84 plus.n23 a_n2146_n3288# 0.021827f
C85 plus.n24 a_n2146_n3288# 0.115963f
C86 plus.n25 a_n2146_n3288# 0.02265f
C87 plus.n26 a_n2146_n3288# 0.115963f
C88 plus.t12 a_n2146_n3288# 0.274921f
C89 plus.n27 a_n2146_n3288# 0.137738f
C90 plus.n28 a_n2146_n3288# 0.605165f
C91 plus.n29 a_n2146_n3288# 0.053392f
C92 plus.t19 a_n2146_n3288# 0.274921f
C93 plus.t5 a_n2146_n3288# 0.271578f
C94 plus.t2 a_n2146_n3288# 0.271578f
C95 plus.n30 a_n2146_n3288# 0.018535f
C96 plus.n31 a_n2146_n3288# 0.053392f
C97 plus.t3 a_n2146_n3288# 0.271578f
C98 plus.n32 a_n2146_n3288# 0.115963f
C99 plus.t0 a_n2146_n3288# 0.271578f
C100 plus.t7 a_n2146_n3288# 0.271578f
C101 plus.t4 a_n2146_n3288# 0.271578f
C102 plus.n33 a_n2146_n3288# 0.115963f
C103 plus.n34 a_n2146_n3288# 0.053392f
C104 plus.t1 a_n2146_n3288# 0.271578f
C105 plus.t8 a_n2146_n3288# 0.271578f
C106 plus.n35 a_n2146_n3288# 0.115963f
C107 plus.t6 a_n2146_n3288# 0.274921f
C108 plus.n36 a_n2146_n3288# 0.13782f
C109 plus.n37 a_n2146_n3288# 0.123162f
C110 plus.n38 a_n2146_n3288# 0.02265f
C111 plus.n39 a_n2146_n3288# 0.115963f
C112 plus.n40 a_n2146_n3288# 0.021827f
C113 plus.n41 a_n2146_n3288# 0.018535f
C114 plus.n42 a_n2146_n3288# 0.053392f
C115 plus.n43 a_n2146_n3288# 0.053392f
C116 plus.n44 a_n2146_n3288# 0.02265f
C117 plus.n45 a_n2146_n3288# 0.115963f
C118 plus.n46 a_n2146_n3288# 0.02265f
C119 plus.n47 a_n2146_n3288# 0.115963f
C120 plus.n48 a_n2146_n3288# 0.02265f
C121 plus.n49 a_n2146_n3288# 0.053392f
C122 plus.n50 a_n2146_n3288# 0.053392f
C123 plus.n51 a_n2146_n3288# 0.053392f
C124 plus.n52 a_n2146_n3288# 0.021827f
C125 plus.n53 a_n2146_n3288# 0.115963f
C126 plus.n54 a_n2146_n3288# 0.02265f
C127 plus.n55 a_n2146_n3288# 0.115963f
C128 plus.n56 a_n2146_n3288# 0.137738f
C129 plus.n57 a_n2146_n3288# 1.68024f
C130 drain_right.t18 a_n2146_n3288# 0.405338f
C131 drain_right.t12 a_n2146_n3288# 0.405338f
C132 drain_right.n0 a_n2146_n3288# 2.65944f
C133 drain_right.t3 a_n2146_n3288# 0.405338f
C134 drain_right.t0 a_n2146_n3288# 0.405338f
C135 drain_right.n1 a_n2146_n3288# 2.65617f
C136 drain_right.n2 a_n2146_n3288# 0.681648f
C137 drain_right.t17 a_n2146_n3288# 0.405338f
C138 drain_right.t10 a_n2146_n3288# 0.405338f
C139 drain_right.n3 a_n2146_n3288# 2.65617f
C140 drain_right.t16 a_n2146_n3288# 0.405338f
C141 drain_right.t8 a_n2146_n3288# 0.405338f
C142 drain_right.n4 a_n2146_n3288# 2.65944f
C143 drain_right.t2 a_n2146_n3288# 0.405338f
C144 drain_right.t19 a_n2146_n3288# 0.405338f
C145 drain_right.n5 a_n2146_n3288# 2.65617f
C146 drain_right.n6 a_n2146_n3288# 0.681648f
C147 drain_right.n7 a_n2146_n3288# 1.70371f
C148 drain_right.t15 a_n2146_n3288# 0.405338f
C149 drain_right.t14 a_n2146_n3288# 0.405338f
C150 drain_right.n8 a_n2146_n3288# 2.65944f
C151 drain_right.t11 a_n2146_n3288# 0.405338f
C152 drain_right.t7 a_n2146_n3288# 0.405338f
C153 drain_right.n9 a_n2146_n3288# 2.65618f
C154 drain_right.n10 a_n2146_n3288# 0.685375f
C155 drain_right.t4 a_n2146_n3288# 0.405338f
C156 drain_right.t13 a_n2146_n3288# 0.405338f
C157 drain_right.n11 a_n2146_n3288# 2.65618f
C158 drain_right.n12 a_n2146_n3288# 0.338632f
C159 drain_right.t5 a_n2146_n3288# 0.405338f
C160 drain_right.t6 a_n2146_n3288# 0.405338f
C161 drain_right.n13 a_n2146_n3288# 2.65618f
C162 drain_right.n14 a_n2146_n3288# 0.338632f
C163 drain_right.t1 a_n2146_n3288# 0.405338f
C164 drain_right.t9 a_n2146_n3288# 0.405338f
C165 drain_right.n15 a_n2146_n3288# 2.65618f
C166 drain_right.n16 a_n2146_n3288# 0.574228f
C167 source.t3 a_n2146_n3288# 2.76154f
C168 source.n0 a_n2146_n3288# 1.37716f
C169 source.t39 a_n2146_n3288# 0.356881f
C170 source.t7 a_n2146_n3288# 0.356881f
C171 source.n1 a_n2146_n3288# 2.25939f
C172 source.n2 a_n2146_n3288# 0.343642f
C173 source.t13 a_n2146_n3288# 0.356881f
C174 source.t17 a_n2146_n3288# 0.356881f
C175 source.n3 a_n2146_n3288# 2.25939f
C176 source.n4 a_n2146_n3288# 0.343642f
C177 source.t0 a_n2146_n3288# 0.356881f
C178 source.t6 a_n2146_n3288# 0.356881f
C179 source.n5 a_n2146_n3288# 2.25939f
C180 source.n6 a_n2146_n3288# 0.343642f
C181 source.t14 a_n2146_n3288# 0.356881f
C182 source.t15 a_n2146_n3288# 0.356881f
C183 source.n7 a_n2146_n3288# 2.25939f
C184 source.n8 a_n2146_n3288# 0.343642f
C185 source.t4 a_n2146_n3288# 2.76156f
C186 source.n9 a_n2146_n3288# 0.476617f
C187 source.t33 a_n2146_n3288# 2.76156f
C188 source.n10 a_n2146_n3288# 0.476617f
C189 source.t34 a_n2146_n3288# 0.356881f
C190 source.t27 a_n2146_n3288# 0.356881f
C191 source.n11 a_n2146_n3288# 2.25939f
C192 source.n12 a_n2146_n3288# 0.343642f
C193 source.t22 a_n2146_n3288# 0.356881f
C194 source.t18 a_n2146_n3288# 0.356881f
C195 source.n13 a_n2146_n3288# 2.25939f
C196 source.n14 a_n2146_n3288# 0.343642f
C197 source.t23 a_n2146_n3288# 0.356881f
C198 source.t20 a_n2146_n3288# 0.356881f
C199 source.n15 a_n2146_n3288# 2.25939f
C200 source.n16 a_n2146_n3288# 0.343642f
C201 source.t28 a_n2146_n3288# 0.356881f
C202 source.t26 a_n2146_n3288# 0.356881f
C203 source.n17 a_n2146_n3288# 2.25939f
C204 source.n18 a_n2146_n3288# 0.343642f
C205 source.t29 a_n2146_n3288# 2.76156f
C206 source.n19 a_n2146_n3288# 1.76822f
C207 source.t8 a_n2146_n3288# 2.76154f
C208 source.n20 a_n2146_n3288# 1.76823f
C209 source.t16 a_n2146_n3288# 0.356881f
C210 source.t1 a_n2146_n3288# 0.356881f
C211 source.n21 a_n2146_n3288# 2.25938f
C212 source.n22 a_n2146_n3288# 0.343655f
C213 source.t5 a_n2146_n3288# 0.356881f
C214 source.t2 a_n2146_n3288# 0.356881f
C215 source.n23 a_n2146_n3288# 2.25938f
C216 source.n24 a_n2146_n3288# 0.343655f
C217 source.t10 a_n2146_n3288# 0.356881f
C218 source.t12 a_n2146_n3288# 0.356881f
C219 source.n25 a_n2146_n3288# 2.25938f
C220 source.n26 a_n2146_n3288# 0.343655f
C221 source.t9 a_n2146_n3288# 0.356881f
C222 source.t38 a_n2146_n3288# 0.356881f
C223 source.n27 a_n2146_n3288# 2.25938f
C224 source.n28 a_n2146_n3288# 0.343655f
C225 source.t11 a_n2146_n3288# 2.76154f
C226 source.n29 a_n2146_n3288# 0.476629f
C227 source.t37 a_n2146_n3288# 2.76154f
C228 source.n30 a_n2146_n3288# 0.476629f
C229 source.t25 a_n2146_n3288# 0.356881f
C230 source.t19 a_n2146_n3288# 0.356881f
C231 source.n31 a_n2146_n3288# 2.25938f
C232 source.n32 a_n2146_n3288# 0.343655f
C233 source.t36 a_n2146_n3288# 0.356881f
C234 source.t21 a_n2146_n3288# 0.356881f
C235 source.n33 a_n2146_n3288# 2.25938f
C236 source.n34 a_n2146_n3288# 0.343655f
C237 source.t31 a_n2146_n3288# 0.356881f
C238 source.t32 a_n2146_n3288# 0.356881f
C239 source.n35 a_n2146_n3288# 2.25938f
C240 source.n36 a_n2146_n3288# 0.343655f
C241 source.t30 a_n2146_n3288# 0.356881f
C242 source.t24 a_n2146_n3288# 0.356881f
C243 source.n37 a_n2146_n3288# 2.25938f
C244 source.n38 a_n2146_n3288# 0.343655f
C245 source.t35 a_n2146_n3288# 2.76154f
C246 source.n39 a_n2146_n3288# 0.617947f
C247 source.n40 a_n2146_n3288# 1.55902f
C248 minus.n0 a_n2146_n3288# 0.052227f
C249 minus.t18 a_n2146_n3288# 0.26892f
C250 minus.t10 a_n2146_n3288# 0.26565f
C251 minus.t14 a_n2146_n3288# 0.26565f
C252 minus.n1 a_n2146_n3288# 0.01813f
C253 minus.n2 a_n2146_n3288# 0.052227f
C254 minus.t13 a_n2146_n3288# 0.26565f
C255 minus.n3 a_n2146_n3288# 0.113432f
C256 minus.t15 a_n2146_n3288# 0.26565f
C257 minus.t6 a_n2146_n3288# 0.26565f
C258 minus.t8 a_n2146_n3288# 0.26565f
C259 minus.n4 a_n2146_n3288# 0.113432f
C260 minus.n5 a_n2146_n3288# 0.052227f
C261 minus.t12 a_n2146_n3288# 0.26565f
C262 minus.t4 a_n2146_n3288# 0.26565f
C263 minus.n6 a_n2146_n3288# 0.113432f
C264 minus.t5 a_n2146_n3288# 0.26892f
C265 minus.n7 a_n2146_n3288# 0.134812f
C266 minus.n8 a_n2146_n3288# 0.120473f
C267 minus.n9 a_n2146_n3288# 0.022155f
C268 minus.n10 a_n2146_n3288# 0.113432f
C269 minus.n11 a_n2146_n3288# 0.02135f
C270 minus.n12 a_n2146_n3288# 0.01813f
C271 minus.n13 a_n2146_n3288# 0.052227f
C272 minus.n14 a_n2146_n3288# 0.052227f
C273 minus.n15 a_n2146_n3288# 0.022155f
C274 minus.n16 a_n2146_n3288# 0.113432f
C275 minus.n17 a_n2146_n3288# 0.022155f
C276 minus.n18 a_n2146_n3288# 0.113432f
C277 minus.n19 a_n2146_n3288# 0.022155f
C278 minus.n20 a_n2146_n3288# 0.052227f
C279 minus.n21 a_n2146_n3288# 0.052227f
C280 minus.n22 a_n2146_n3288# 0.052227f
C281 minus.n23 a_n2146_n3288# 0.02135f
C282 minus.n24 a_n2146_n3288# 0.113432f
C283 minus.n25 a_n2146_n3288# 0.022155f
C284 minus.n26 a_n2146_n3288# 0.113432f
C285 minus.n27 a_n2146_n3288# 0.134732f
C286 minus.n28 a_n2146_n3288# 1.9374f
C287 minus.n29 a_n2146_n3288# 0.052227f
C288 minus.t3 a_n2146_n3288# 0.26565f
C289 minus.t0 a_n2146_n3288# 0.26565f
C290 minus.n30 a_n2146_n3288# 0.01813f
C291 minus.n31 a_n2146_n3288# 0.052227f
C292 minus.t9 a_n2146_n3288# 0.26565f
C293 minus.t2 a_n2146_n3288# 0.26565f
C294 minus.t19 a_n2146_n3288# 0.26565f
C295 minus.n32 a_n2146_n3288# 0.113432f
C296 minus.n33 a_n2146_n3288# 0.052227f
C297 minus.t16 a_n2146_n3288# 0.26565f
C298 minus.t7 a_n2146_n3288# 0.26565f
C299 minus.n34 a_n2146_n3288# 0.113432f
C300 minus.t1 a_n2146_n3288# 0.26892f
C301 minus.n35 a_n2146_n3288# 0.134812f
C302 minus.n36 a_n2146_n3288# 0.120473f
C303 minus.n37 a_n2146_n3288# 0.022155f
C304 minus.n38 a_n2146_n3288# 0.113432f
C305 minus.n39 a_n2146_n3288# 0.02135f
C306 minus.n40 a_n2146_n3288# 0.01813f
C307 minus.n41 a_n2146_n3288# 0.052227f
C308 minus.n42 a_n2146_n3288# 0.052227f
C309 minus.n43 a_n2146_n3288# 0.022155f
C310 minus.n44 a_n2146_n3288# 0.113432f
C311 minus.n45 a_n2146_n3288# 0.022155f
C312 minus.n46 a_n2146_n3288# 0.113432f
C313 minus.t17 a_n2146_n3288# 0.26565f
C314 minus.n47 a_n2146_n3288# 0.113432f
C315 minus.n48 a_n2146_n3288# 0.022155f
C316 minus.n49 a_n2146_n3288# 0.052227f
C317 minus.n50 a_n2146_n3288# 0.052227f
C318 minus.n51 a_n2146_n3288# 0.052227f
C319 minus.n52 a_n2146_n3288# 0.02135f
C320 minus.n53 a_n2146_n3288# 0.113432f
C321 minus.n54 a_n2146_n3288# 0.022155f
C322 minus.n55 a_n2146_n3288# 0.113432f
C323 minus.t11 a_n2146_n3288# 0.26892f
C324 minus.n56 a_n2146_n3288# 0.134732f
C325 minus.n57 a_n2146_n3288# 0.348941f
C326 minus.n58 a_n2146_n3288# 2.34325f
.ends

