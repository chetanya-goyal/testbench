* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X2 drain_right.t9 minus.t0 source.t6 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X3 source.t0 plus.t0 drain_left.t9 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X4 drain_right.t8 minus.t1 source.t11 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t12 minus.t2 drain_right.t7 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right.t6 minus.t3 source.t14 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X7 a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X8 drain_left.t8 plus.t1 source.t16 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_left.t7 plus.t2 source.t19 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X10 source.t4 plus.t3 drain_left.t6 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X11 source.t7 minus.t4 drain_right.t5 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X12 drain_right.t4 minus.t5 source.t8 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X13 source.t18 plus.t4 drain_left.t5 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 source.t9 minus.t6 drain_right.t3 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 drain_left.t4 plus.t5 source.t5 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 drain_right.t2 minus.t7 source.t13 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X17 drain_right.t1 minus.t8 source.t15 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X18 source.t17 plus.t6 drain_left.t3 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 drain_left.t2 plus.t7 source.t1 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X20 a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X21 source.t10 minus.t9 drain_right.t0 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X22 drain_left.t1 plus.t8 source.t2 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X23 drain_left.t0 plus.t9 source.t3 a_n1832_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
R0 minus.n3 minus.t7 172.006
R1 minus.n13 minus.t3 172.006
R2 minus.n9 minus.n8 161.3
R3 minus.n7 minus.n0 161.3
R4 minus.n6 minus.n5 161.3
R5 minus.n19 minus.n18 161.3
R6 minus.n17 minus.n10 161.3
R7 minus.n16 minus.n15 161.3
R8 minus.n2 minus.t6 145.805
R9 minus.n1 minus.t5 145.805
R10 minus.n6 minus.t4 145.805
R11 minus.n8 minus.t1 145.805
R12 minus.n12 minus.t9 145.805
R13 minus.n11 minus.t8 145.805
R14 minus.n16 minus.t2 145.805
R15 minus.n18 minus.t0 145.805
R16 minus.n4 minus.n1 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n8 minus.n7 45.2793
R23 minus.n18 minus.n17 45.2793
R24 minus.n4 minus.n3 45.1669
R25 minus.n14 minus.n13 45.1669
R26 minus.n20 minus.n9 28.5857
R27 minus.n3 minus.n2 14.3992
R28 minus.n13 minus.n12 14.3992
R29 minus.n20 minus.n19 6.60088
R30 minus.n7 minus.n6 2.92171
R31 minus.n17 minus.n16 2.92171
R32 minus.n5 minus.n4 0.285035
R33 minus.n15 minus.n14 0.285035
R34 minus.n9 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n15 minus.n10 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 source.n42 source.n40 289.615
R40 source.n30 source.n28 289.615
R41 source.n2 source.n0 289.615
R42 source.n14 source.n12 289.615
R43 source.n43 source.n42 185
R44 source.n31 source.n30 185
R45 source.n3 source.n2 185
R46 source.n15 source.n14 185
R47 source.t6 source.n41 167.117
R48 source.t2 source.n29 167.117
R49 source.t19 source.n1 167.117
R50 source.t13 source.n13 167.117
R51 source.n9 source.n8 84.1169
R52 source.n11 source.n10 84.1169
R53 source.n21 source.n20 84.1169
R54 source.n23 source.n22 84.1169
R55 source.n39 source.n38 84.1168
R56 source.n37 source.n36 84.1168
R57 source.n27 source.n26 84.1168
R58 source.n25 source.n24 84.1168
R59 source.n42 source.t6 52.3082
R60 source.n30 source.t2 52.3082
R61 source.n2 source.t19 52.3082
R62 source.n14 source.t13 52.3082
R63 source.n47 source.n46 31.4096
R64 source.n35 source.n34 31.4096
R65 source.n7 source.n6 31.4096
R66 source.n19 source.n18 31.4096
R67 source.n25 source.n23 15.3154
R68 source.n38 source.t15 9.9005
R69 source.n38 source.t12 9.9005
R70 source.n36 source.t14 9.9005
R71 source.n36 source.t10 9.9005
R72 source.n26 source.t16 9.9005
R73 source.n26 source.t4 9.9005
R74 source.n24 source.t3 9.9005
R75 source.n24 source.t0 9.9005
R76 source.n8 source.t5 9.9005
R77 source.n8 source.t18 9.9005
R78 source.n10 source.t1 9.9005
R79 source.n10 source.t17 9.9005
R80 source.n20 source.t8 9.9005
R81 source.n20 source.t9 9.9005
R82 source.n22 source.t11 9.9005
R83 source.n22 source.t7 9.9005
R84 source.n43 source.n41 9.71174
R85 source.n31 source.n29 9.71174
R86 source.n3 source.n1 9.71174
R87 source.n15 source.n13 9.71174
R88 source.n46 source.n45 9.45567
R89 source.n34 source.n33 9.45567
R90 source.n6 source.n5 9.45567
R91 source.n18 source.n17 9.45567
R92 source.n45 source.n44 9.3005
R93 source.n33 source.n32 9.3005
R94 source.n5 source.n4 9.3005
R95 source.n17 source.n16 9.3005
R96 source.n48 source.n7 8.8499
R97 source.n46 source.n40 8.14595
R98 source.n34 source.n28 8.14595
R99 source.n6 source.n0 8.14595
R100 source.n18 source.n12 8.14595
R101 source.n44 source.n43 7.3702
R102 source.n32 source.n31 7.3702
R103 source.n4 source.n3 7.3702
R104 source.n16 source.n15 7.3702
R105 source.n44 source.n40 5.81868
R106 source.n32 source.n28 5.81868
R107 source.n4 source.n0 5.81868
R108 source.n16 source.n12 5.81868
R109 source.n48 source.n47 5.66429
R110 source.n45 source.n41 3.44771
R111 source.n33 source.n29 3.44771
R112 source.n5 source.n1 3.44771
R113 source.n17 source.n13 3.44771
R114 source.n19 source.n11 0.87119
R115 source.n37 source.n35 0.87119
R116 source.n23 source.n21 0.802224
R117 source.n21 source.n19 0.802224
R118 source.n11 source.n9 0.802224
R119 source.n9 source.n7 0.802224
R120 source.n27 source.n25 0.802224
R121 source.n35 source.n27 0.802224
R122 source.n39 source.n37 0.802224
R123 source.n47 source.n39 0.802224
R124 source source.n48 0.188
R125 drain_right.n2 drain_right.n0 289.615
R126 drain_right.n16 drain_right.n14 289.615
R127 drain_right.n3 drain_right.n2 185
R128 drain_right.n17 drain_right.n16 185
R129 drain_right.t6 drain_right.n1 167.117
R130 drain_right.t8 drain_right.n15 167.117
R131 drain_right.n13 drain_right.n11 101.597
R132 drain_right.n10 drain_right.n9 101.341
R133 drain_right.n13 drain_right.n12 100.796
R134 drain_right.n8 drain_right.n7 100.796
R135 drain_right.n2 drain_right.t6 52.3082
R136 drain_right.n16 drain_right.t8 52.3082
R137 drain_right.n8 drain_right.n6 48.8901
R138 drain_right.n21 drain_right.n20 48.0884
R139 drain_right drain_right.n10 22.6454
R140 drain_right.n9 drain_right.t7 9.9005
R141 drain_right.n9 drain_right.t9 9.9005
R142 drain_right.n7 drain_right.t0 9.9005
R143 drain_right.n7 drain_right.t1 9.9005
R144 drain_right.n11 drain_right.t3 9.9005
R145 drain_right.n11 drain_right.t2 9.9005
R146 drain_right.n12 drain_right.t5 9.9005
R147 drain_right.n12 drain_right.t4 9.9005
R148 drain_right.n3 drain_right.n1 9.71174
R149 drain_right.n17 drain_right.n15 9.71174
R150 drain_right.n6 drain_right.n5 9.45567
R151 drain_right.n20 drain_right.n19 9.45567
R152 drain_right.n5 drain_right.n4 9.3005
R153 drain_right.n19 drain_right.n18 9.3005
R154 drain_right.n6 drain_right.n0 8.14595
R155 drain_right.n20 drain_right.n14 8.14595
R156 drain_right.n4 drain_right.n3 7.3702
R157 drain_right.n18 drain_right.n17 7.3702
R158 drain_right drain_right.n21 6.05408
R159 drain_right.n4 drain_right.n0 5.81868
R160 drain_right.n18 drain_right.n14 5.81868
R161 drain_right.n5 drain_right.n1 3.44771
R162 drain_right.n19 drain_right.n15 3.44771
R163 drain_right.n21 drain_right.n13 0.802224
R164 drain_right.n10 drain_right.n8 0.145585
R165 plus.n3 plus.t7 172.006
R166 plus.n13 plus.t8 172.006
R167 plus.n6 plus.n1 161.3
R168 plus.n7 plus.n0 161.3
R169 plus.n9 plus.n8 161.3
R170 plus.n16 plus.n11 161.3
R171 plus.n17 plus.n10 161.3
R172 plus.n19 plus.n18 161.3
R173 plus.n8 plus.t2 145.805
R174 plus.n6 plus.t4 145.805
R175 plus.n5 plus.t5 145.805
R176 plus.n4 plus.t6 145.805
R177 plus.n18 plus.t9 145.805
R178 plus.n16 plus.t0 145.805
R179 plus.n15 plus.t1 145.805
R180 plus.n14 plus.t3 145.805
R181 plus.n5 plus.n2 80.6037
R182 plus.n15 plus.n12 80.6037
R183 plus.n6 plus.n5 48.2005
R184 plus.n5 plus.n4 48.2005
R185 plus.n16 plus.n15 48.2005
R186 plus.n15 plus.n14 48.2005
R187 plus.n8 plus.n7 45.2793
R188 plus.n18 plus.n17 45.2793
R189 plus.n3 plus.n2 45.1669
R190 plus.n13 plus.n12 45.1669
R191 plus plus.n19 26.2547
R192 plus.n4 plus.n3 14.3992
R193 plus.n14 plus.n13 14.3992
R194 plus plus.n9 8.45694
R195 plus.n7 plus.n6 2.92171
R196 plus.n17 plus.n16 2.92171
R197 plus.n2 plus.n1 0.285035
R198 plus.n12 plus.n11 0.285035
R199 plus.n1 plus.n0 0.189894
R200 plus.n9 plus.n0 0.189894
R201 plus.n19 plus.n10 0.189894
R202 plus.n11 plus.n10 0.189894
R203 drain_left.n2 drain_left.n0 289.615
R204 drain_left.n13 drain_left.n11 289.615
R205 drain_left.n3 drain_left.n2 185
R206 drain_left.n14 drain_left.n13 185
R207 drain_left.t0 drain_left.n1 167.117
R208 drain_left.t2 drain_left.n12 167.117
R209 drain_left.n10 drain_left.n9 101.341
R210 drain_left.n21 drain_left.n20 100.796
R211 drain_left.n19 drain_left.n18 100.796
R212 drain_left.n8 drain_left.n7 100.796
R213 drain_left.n2 drain_left.t0 52.3082
R214 drain_left.n13 drain_left.t2 52.3082
R215 drain_left.n8 drain_left.n6 48.8901
R216 drain_left.n19 drain_left.n17 48.8901
R217 drain_left drain_left.n10 23.1986
R218 drain_left.n9 drain_left.t6 9.9005
R219 drain_left.n9 drain_left.t1 9.9005
R220 drain_left.n7 drain_left.t9 9.9005
R221 drain_left.n7 drain_left.t8 9.9005
R222 drain_left.n20 drain_left.t5 9.9005
R223 drain_left.n20 drain_left.t7 9.9005
R224 drain_left.n18 drain_left.t3 9.9005
R225 drain_left.n18 drain_left.t4 9.9005
R226 drain_left.n3 drain_left.n1 9.71174
R227 drain_left.n14 drain_left.n12 9.71174
R228 drain_left.n6 drain_left.n5 9.45567
R229 drain_left.n17 drain_left.n16 9.45567
R230 drain_left.n5 drain_left.n4 9.3005
R231 drain_left.n16 drain_left.n15 9.3005
R232 drain_left.n6 drain_left.n0 8.14595
R233 drain_left.n17 drain_left.n11 8.14595
R234 drain_left.n4 drain_left.n3 7.3702
R235 drain_left.n15 drain_left.n14 7.3702
R236 drain_left drain_left.n21 6.45494
R237 drain_left.n4 drain_left.n0 5.81868
R238 drain_left.n15 drain_left.n11 5.81868
R239 drain_left.n5 drain_left.n1 3.44771
R240 drain_left.n16 drain_left.n12 3.44771
R241 drain_left.n21 drain_left.n19 0.802224
R242 drain_left.n10 drain_left.n8 0.145585
C0 plus minus 3.58561f
C1 drain_right minus 1.38042f
C2 source drain_left 4.60769f
C3 plus drain_right 0.340481f
C4 minus drain_left 0.178506f
C5 minus source 1.68007f
C6 plus drain_left 1.55771f
C7 plus source 1.69413f
C8 drain_right drain_left 0.906561f
C9 drain_right source 4.60684f
C10 drain_right a_n1832_n1288# 3.69474f
C11 drain_left a_n1832_n1288# 3.93986f
C12 source a_n1832_n1288# 2.584849f
C13 minus a_n1832_n1288# 6.330395f
C14 plus a_n1832_n1288# 6.885422f
C15 drain_left.n0 a_n1832_n1288# 0.027438f
C16 drain_left.n1 a_n1832_n1288# 0.06071f
C17 drain_left.t0 a_n1832_n1288# 0.045559f
C18 drain_left.n2 a_n1832_n1288# 0.047514f
C19 drain_left.n3 a_n1832_n1288# 0.015317f
C20 drain_left.n4 a_n1832_n1288# 0.010102f
C21 drain_left.n5 a_n1832_n1288# 0.133819f
C22 drain_left.n6 a_n1832_n1288# 0.044447f
C23 drain_left.t9 a_n1832_n1288# 0.029711f
C24 drain_left.t8 a_n1832_n1288# 0.029711f
C25 drain_left.n7 a_n1832_n1288# 0.186651f
C26 drain_left.n8 a_n1832_n1288# 0.287033f
C27 drain_left.t6 a_n1832_n1288# 0.029711f
C28 drain_left.t1 a_n1832_n1288# 0.029711f
C29 drain_left.n9 a_n1832_n1288# 0.187911f
C30 drain_left.n10 a_n1832_n1288# 0.778598f
C31 drain_left.n11 a_n1832_n1288# 0.027438f
C32 drain_left.n12 a_n1832_n1288# 0.06071f
C33 drain_left.t2 a_n1832_n1288# 0.045559f
C34 drain_left.n13 a_n1832_n1288# 0.047514f
C35 drain_left.n14 a_n1832_n1288# 0.015317f
C36 drain_left.n15 a_n1832_n1288# 0.010102f
C37 drain_left.n16 a_n1832_n1288# 0.133819f
C38 drain_left.n17 a_n1832_n1288# 0.044447f
C39 drain_left.t3 a_n1832_n1288# 0.029711f
C40 drain_left.t4 a_n1832_n1288# 0.029711f
C41 drain_left.n18 a_n1832_n1288# 0.186652f
C42 drain_left.n19 a_n1832_n1288# 0.323803f
C43 drain_left.t5 a_n1832_n1288# 0.029711f
C44 drain_left.t7 a_n1832_n1288# 0.029711f
C45 drain_left.n20 a_n1832_n1288# 0.186652f
C46 drain_left.n21 a_n1832_n1288# 0.404932f
C47 plus.n0 a_n1832_n1288# 0.026043f
C48 plus.t2 a_n1832_n1288# 0.096776f
C49 plus.t4 a_n1832_n1288# 0.096776f
C50 plus.n1 a_n1832_n1288# 0.03475f
C51 plus.t5 a_n1832_n1288# 0.096776f
C52 plus.n2 a_n1832_n1288# 0.125875f
C53 plus.t6 a_n1832_n1288# 0.096776f
C54 plus.t7 a_n1832_n1288# 0.107205f
C55 plus.n3 a_n1832_n1288# 0.059305f
C56 plus.n4 a_n1832_n1288# 0.074002f
C57 plus.n5 a_n1832_n1288# 0.074439f
C58 plus.n6 a_n1832_n1288# 0.068851f
C59 plus.n7 a_n1832_n1288# 0.00591f
C60 plus.n8 a_n1832_n1288# 0.068208f
C61 plus.n9 a_n1832_n1288# 0.192671f
C62 plus.n10 a_n1832_n1288# 0.026043f
C63 plus.t9 a_n1832_n1288# 0.096776f
C64 plus.n11 a_n1832_n1288# 0.03475f
C65 plus.t0 a_n1832_n1288# 0.096776f
C66 plus.n12 a_n1832_n1288# 0.125875f
C67 plus.t1 a_n1832_n1288# 0.096776f
C68 plus.t8 a_n1832_n1288# 0.107205f
C69 plus.n13 a_n1832_n1288# 0.059305f
C70 plus.t3 a_n1832_n1288# 0.096776f
C71 plus.n14 a_n1832_n1288# 0.074002f
C72 plus.n15 a_n1832_n1288# 0.074439f
C73 plus.n16 a_n1832_n1288# 0.068851f
C74 plus.n17 a_n1832_n1288# 0.00591f
C75 plus.n18 a_n1832_n1288# 0.068208f
C76 plus.n19 a_n1832_n1288# 0.597725f
C77 drain_right.n0 a_n1832_n1288# 0.027884f
C78 drain_right.n1 a_n1832_n1288# 0.061696f
C79 drain_right.t6 a_n1832_n1288# 0.0463f
C80 drain_right.n2 a_n1832_n1288# 0.048286f
C81 drain_right.n3 a_n1832_n1288# 0.015566f
C82 drain_right.n4 a_n1832_n1288# 0.010266f
C83 drain_right.n5 a_n1832_n1288# 0.135993f
C84 drain_right.n6 a_n1832_n1288# 0.045169f
C85 drain_right.t0 a_n1832_n1288# 0.030193f
C86 drain_right.t1 a_n1832_n1288# 0.030193f
C87 drain_right.n7 a_n1832_n1288# 0.189683f
C88 drain_right.n8 a_n1832_n1288# 0.291696f
C89 drain_right.t7 a_n1832_n1288# 0.030193f
C90 drain_right.t9 a_n1832_n1288# 0.030193f
C91 drain_right.n9 a_n1832_n1288# 0.190964f
C92 drain_right.n10 a_n1832_n1288# 0.753811f
C93 drain_right.t3 a_n1832_n1288# 0.030193f
C94 drain_right.t2 a_n1832_n1288# 0.030193f
C95 drain_right.n11 a_n1832_n1288# 0.191678f
C96 drain_right.t5 a_n1832_n1288# 0.030193f
C97 drain_right.t4 a_n1832_n1288# 0.030193f
C98 drain_right.n12 a_n1832_n1288# 0.189684f
C99 drain_right.n13 a_n1832_n1288# 0.495551f
C100 drain_right.n14 a_n1832_n1288# 0.027884f
C101 drain_right.n15 a_n1832_n1288# 0.061696f
C102 drain_right.t8 a_n1832_n1288# 0.0463f
C103 drain_right.n16 a_n1832_n1288# 0.048286f
C104 drain_right.n17 a_n1832_n1288# 0.015566f
C105 drain_right.n18 a_n1832_n1288# 0.010266f
C106 drain_right.n19 a_n1832_n1288# 0.135993f
C107 drain_right.n20 a_n1832_n1288# 0.043766f
C108 drain_right.n21 a_n1832_n1288# 0.257098f
C109 source.n0 a_n1832_n1288# 0.034603f
C110 source.n1 a_n1832_n1288# 0.076564f
C111 source.t19 a_n1832_n1288# 0.057457f
C112 source.n2 a_n1832_n1288# 0.059922f
C113 source.n3 a_n1832_n1288# 0.019317f
C114 source.n4 a_n1832_n1288# 0.01274f
C115 source.n5 a_n1832_n1288# 0.168766f
C116 source.n6 a_n1832_n1288# 0.037933f
C117 source.n7 a_n1832_n1288# 0.392982f
C118 source.t5 a_n1832_n1288# 0.037469f
C119 source.t18 a_n1832_n1288# 0.037469f
C120 source.n8 a_n1832_n1288# 0.200311f
C121 source.n9 a_n1832_n1288# 0.30681f
C122 source.t1 a_n1832_n1288# 0.037469f
C123 source.t17 a_n1832_n1288# 0.037469f
C124 source.n10 a_n1832_n1288# 0.200311f
C125 source.n11 a_n1832_n1288# 0.312078f
C126 source.n12 a_n1832_n1288# 0.034603f
C127 source.n13 a_n1832_n1288# 0.076564f
C128 source.t13 a_n1832_n1288# 0.057457f
C129 source.n14 a_n1832_n1288# 0.059922f
C130 source.n15 a_n1832_n1288# 0.019317f
C131 source.n16 a_n1832_n1288# 0.01274f
C132 source.n17 a_n1832_n1288# 0.168766f
C133 source.n18 a_n1832_n1288# 0.037933f
C134 source.n19 a_n1832_n1288# 0.147277f
C135 source.t8 a_n1832_n1288# 0.037469f
C136 source.t9 a_n1832_n1288# 0.037469f
C137 source.n20 a_n1832_n1288# 0.200311f
C138 source.n21 a_n1832_n1288# 0.30681f
C139 source.t11 a_n1832_n1288# 0.037469f
C140 source.t7 a_n1832_n1288# 0.037469f
C141 source.n22 a_n1832_n1288# 0.200311f
C142 source.n23 a_n1832_n1288# 0.844542f
C143 source.t3 a_n1832_n1288# 0.037469f
C144 source.t0 a_n1832_n1288# 0.037469f
C145 source.n24 a_n1832_n1288# 0.20031f
C146 source.n25 a_n1832_n1288# 0.844543f
C147 source.t16 a_n1832_n1288# 0.037469f
C148 source.t4 a_n1832_n1288# 0.037469f
C149 source.n26 a_n1832_n1288# 0.20031f
C150 source.n27 a_n1832_n1288# 0.306811f
C151 source.n28 a_n1832_n1288# 0.034603f
C152 source.n29 a_n1832_n1288# 0.076564f
C153 source.t2 a_n1832_n1288# 0.057457f
C154 source.n30 a_n1832_n1288# 0.059922f
C155 source.n31 a_n1832_n1288# 0.019317f
C156 source.n32 a_n1832_n1288# 0.01274f
C157 source.n33 a_n1832_n1288# 0.168766f
C158 source.n34 a_n1832_n1288# 0.037933f
C159 source.n35 a_n1832_n1288# 0.147277f
C160 source.t14 a_n1832_n1288# 0.037469f
C161 source.t10 a_n1832_n1288# 0.037469f
C162 source.n36 a_n1832_n1288# 0.20031f
C163 source.n37 a_n1832_n1288# 0.312079f
C164 source.t15 a_n1832_n1288# 0.037469f
C165 source.t12 a_n1832_n1288# 0.037469f
C166 source.n38 a_n1832_n1288# 0.20031f
C167 source.n39 a_n1832_n1288# 0.306811f
C168 source.n40 a_n1832_n1288# 0.034603f
C169 source.n41 a_n1832_n1288# 0.076564f
C170 source.t6 a_n1832_n1288# 0.057457f
C171 source.n42 a_n1832_n1288# 0.059922f
C172 source.n43 a_n1832_n1288# 0.019317f
C173 source.n44 a_n1832_n1288# 0.01274f
C174 source.n45 a_n1832_n1288# 0.168766f
C175 source.n46 a_n1832_n1288# 0.037933f
C176 source.n47 a_n1832_n1288# 0.266141f
C177 source.n48 a_n1832_n1288# 0.59473f
C178 minus.n0 a_n1832_n1288# 0.025667f
C179 minus.t5 a_n1832_n1288# 0.095381f
C180 minus.n1 a_n1832_n1288# 0.073366f
C181 minus.t4 a_n1832_n1288# 0.095381f
C182 minus.t7 a_n1832_n1288# 0.105659f
C183 minus.t6 a_n1832_n1288# 0.095381f
C184 minus.n2 a_n1832_n1288# 0.072935f
C185 minus.n3 a_n1832_n1288# 0.05845f
C186 minus.n4 a_n1832_n1288# 0.124061f
C187 minus.n5 a_n1832_n1288# 0.034249f
C188 minus.n6 a_n1832_n1288# 0.067858f
C189 minus.n7 a_n1832_n1288# 0.005824f
C190 minus.t1 a_n1832_n1288# 0.095381f
C191 minus.n8 a_n1832_n1288# 0.067225f
C192 minus.n9 a_n1832_n1288# 0.616752f
C193 minus.n10 a_n1832_n1288# 0.025667f
C194 minus.t8 a_n1832_n1288# 0.095381f
C195 minus.n11 a_n1832_n1288# 0.073366f
C196 minus.t3 a_n1832_n1288# 0.105659f
C197 minus.t9 a_n1832_n1288# 0.095381f
C198 minus.n12 a_n1832_n1288# 0.072935f
C199 minus.n13 a_n1832_n1288# 0.05845f
C200 minus.n14 a_n1832_n1288# 0.124061f
C201 minus.n15 a_n1832_n1288# 0.034249f
C202 minus.t2 a_n1832_n1288# 0.095381f
C203 minus.n16 a_n1832_n1288# 0.067858f
C204 minus.n17 a_n1832_n1288# 0.005824f
C205 minus.t0 a_n1832_n1288# 0.095381f
C206 minus.n18 a_n1832_n1288# 0.067225f
C207 minus.n19 a_n1832_n1288# 0.173876f
C208 minus.n20 a_n1832_n1288# 0.758884f
.ends

