* NGSPICE file created from diffpair603.ext - technology: sky130A

.subckt diffpair603 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t9 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t12 plus.t1 drain_left.t6 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 source.t1 minus.t0 drain_right.t7 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X3 source.t11 plus.t2 drain_left.t5 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X4 source.t7 plus.t3 drain_left.t4 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X5 drain_right.t6 minus.t1 source.t2 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X6 source.t3 minus.t2 drain_right.t5 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X7 a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X8 a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X9 drain_right.t4 minus.t3 source.t0 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X10 drain_left.t3 plus.t4 source.t10 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X11 drain_left.t2 plus.t5 source.t14 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X12 drain_right.t3 minus.t4 source.t15 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X13 drain_right.t2 minus.t5 source.t4 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X14 source.t6 minus.t6 drain_right.t1 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 drain_left.t1 plus.t6 source.t13 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X16 source.t5 minus.t7 drain_right.t0 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X17 a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X18 source.t8 plus.t7 drain_left.t0 a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# a_n1546_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
R0 plus.n2 plus.t3 1063.55
R1 plus.n10 plus.t0 1063.55
R2 plus.n6 plus.t4 1042.57
R3 plus.n5 plus.t7 1042.57
R4 plus.n1 plus.t6 1042.57
R5 plus.n14 plus.t2 1042.57
R6 plus.n13 plus.t5 1042.57
R7 plus.n9 plus.t1 1042.57
R8 plus.n4 plus.n3 161.3
R9 plus.n5 plus.n0 161.3
R10 plus.n7 plus.n6 161.3
R11 plus.n12 plus.n11 161.3
R12 plus.n13 plus.n8 161.3
R13 plus.n15 plus.n14 161.3
R14 plus.n3 plus.n2 70.4033
R15 plus.n11 plus.n10 70.4033
R16 plus.n6 plus.n5 48.2005
R17 plus.n14 plus.n13 48.2005
R18 plus plus.n15 31.9839
R19 plus.n4 plus.n1 24.1005
R20 plus.n5 plus.n4 24.1005
R21 plus.n13 plus.n12 24.1005
R22 plus.n12 plus.n9 24.1005
R23 plus.n2 plus.n1 20.9576
R24 plus.n10 plus.n9 20.9576
R25 plus plus.n7 15.2694
R26 plus.n3 plus.n0 0.189894
R27 plus.n7 plus.n0 0.189894
R28 plus.n15 plus.n8 0.189894
R29 plus.n11 plus.n8 0.189894
R30 source.n0 source.t10 44.1297
R31 source.n3 source.t7 44.1296
R32 source.n4 source.t4 44.1296
R33 source.n7 source.t5 44.1296
R34 source.n15 source.t15 44.1295
R35 source.n12 source.t3 44.1295
R36 source.n11 source.t9 44.1295
R37 source.n8 source.t11 44.1295
R38 source.n2 source.n1 43.1397
R39 source.n6 source.n5 43.1397
R40 source.n14 source.n13 43.1396
R41 source.n10 source.n9 43.1396
R42 source.n8 source.n7 28.0638
R43 source.n16 source.n0 22.4432
R44 source.n16 source.n15 5.62119
R45 source.n13 source.t2 0.9905
R46 source.n13 source.t6 0.9905
R47 source.n9 source.t14 0.9905
R48 source.n9 source.t12 0.9905
R49 source.n1 source.t13 0.9905
R50 source.n1 source.t8 0.9905
R51 source.n5 source.t0 0.9905
R52 source.n5 source.t1 0.9905
R53 source.n7 source.n6 0.716017
R54 source.n6 source.n4 0.716017
R55 source.n3 source.n2 0.716017
R56 source.n2 source.n0 0.716017
R57 source.n10 source.n8 0.716017
R58 source.n11 source.n10 0.716017
R59 source.n14 source.n12 0.716017
R60 source.n15 source.n14 0.716017
R61 source.n4 source.n3 0.470328
R62 source.n12 source.n11 0.470328
R63 source source.n16 0.188
R64 drain_left.n5 drain_left.n3 60.534
R65 drain_left.n2 drain_left.n1 60.1208
R66 drain_left.n2 drain_left.n0 60.1208
R67 drain_left.n5 drain_left.n4 59.8185
R68 drain_left drain_left.n2 35.932
R69 drain_left drain_left.n5 6.36873
R70 drain_left.n1 drain_left.t6 0.9905
R71 drain_left.n1 drain_left.t7 0.9905
R72 drain_left.n0 drain_left.t5 0.9905
R73 drain_left.n0 drain_left.t2 0.9905
R74 drain_left.n4 drain_left.t0 0.9905
R75 drain_left.n4 drain_left.t3 0.9905
R76 drain_left.n3 drain_left.t4 0.9905
R77 drain_left.n3 drain_left.t1 0.9905
R78 minus.n2 minus.t5 1063.55
R79 minus.n10 minus.t2 1063.55
R80 minus.n1 minus.t0 1042.57
R81 minus.n5 minus.t3 1042.57
R82 minus.n6 minus.t7 1042.57
R83 minus.n9 minus.t1 1042.57
R84 minus.n13 minus.t6 1042.57
R85 minus.n14 minus.t4 1042.57
R86 minus.n7 minus.n6 161.3
R87 minus.n5 minus.n0 161.3
R88 minus.n4 minus.n3 161.3
R89 minus.n15 minus.n14 161.3
R90 minus.n13 minus.n8 161.3
R91 minus.n12 minus.n11 161.3
R92 minus.n3 minus.n2 70.4033
R93 minus.n11 minus.n10 70.4033
R94 minus.n6 minus.n5 48.2005
R95 minus.n14 minus.n13 48.2005
R96 minus.n16 minus.n7 41.1331
R97 minus.n5 minus.n4 24.1005
R98 minus.n4 minus.n1 24.1005
R99 minus.n12 minus.n9 24.1005
R100 minus.n13 minus.n12 24.1005
R101 minus.n2 minus.n1 20.9576
R102 minus.n10 minus.n9 20.9576
R103 minus.n16 minus.n15 6.5952
R104 minus.n7 minus.n0 0.189894
R105 minus.n3 minus.n0 0.189894
R106 minus.n11 minus.n8 0.189894
R107 minus.n15 minus.n8 0.189894
R108 minus minus.n16 0.188
R109 drain_right.n5 drain_right.n3 60.534
R110 drain_right.n2 drain_right.n1 60.1208
R111 drain_right.n2 drain_right.n0 60.1208
R112 drain_right.n5 drain_right.n4 59.8185
R113 drain_right drain_right.n2 35.3788
R114 drain_right drain_right.n5 6.36873
R115 drain_right.n1 drain_right.t1 0.9905
R116 drain_right.n1 drain_right.t3 0.9905
R117 drain_right.n0 drain_right.t5 0.9905
R118 drain_right.n0 drain_right.t6 0.9905
R119 drain_right.n3 drain_right.t7 0.9905
R120 drain_right.n3 drain_right.t2 0.9905
R121 drain_right.n4 drain_right.t0 0.9905
R122 drain_right.n4 drain_right.t4 0.9905
C0 drain_right drain_left 0.727126f
C1 drain_left plus 7.551859f
C2 source drain_left 20.4899f
C3 minus drain_right 7.40383f
C4 minus plus 6.55316f
C5 source minus 6.75272f
C6 drain_right plus 0.302201f
C7 source drain_right 20.4904f
C8 source plus 6.76675f
C9 minus drain_left 0.171215f
C10 drain_right a_n1546_n4888# 7.19291f
C11 drain_left a_n1546_n4888# 7.43518f
C12 source a_n1546_n4888# 13.227349f
C13 minus a_n1546_n4888# 6.500572f
C14 plus a_n1546_n4888# 8.84733f
C15 drain_right.t5 a_n1546_n4888# 0.462948f
C16 drain_right.t6 a_n1546_n4888# 0.462948f
C17 drain_right.n0 a_n1546_n4888# 4.23417f
C18 drain_right.t1 a_n1546_n4888# 0.462948f
C19 drain_right.t3 a_n1546_n4888# 0.462948f
C20 drain_right.n1 a_n1546_n4888# 4.23417f
C21 drain_right.n2 a_n1546_n4888# 2.58271f
C22 drain_right.t7 a_n1546_n4888# 0.462948f
C23 drain_right.t2 a_n1546_n4888# 0.462948f
C24 drain_right.n3 a_n1546_n4888# 4.23703f
C25 drain_right.t0 a_n1546_n4888# 0.462948f
C26 drain_right.t4 a_n1546_n4888# 0.462948f
C27 drain_right.n4 a_n1546_n4888# 4.23237f
C28 drain_right.n5 a_n1546_n4888# 1.02331f
C29 minus.n0 a_n1546_n4888# 0.049176f
C30 minus.t0 a_n1546_n4888# 1.3926f
C31 minus.n1 a_n1546_n4888# 0.528136f
C32 minus.t5 a_n1546_n4888# 1.40292f
C33 minus.n2 a_n1546_n4888# 0.513191f
C34 minus.n3 a_n1546_n4888# 0.162003f
C35 minus.n4 a_n1546_n4888# 0.011159f
C36 minus.t3 a_n1546_n4888# 1.3926f
C37 minus.n5 a_n1546_n4888# 0.528136f
C38 minus.t7 a_n1546_n4888# 1.3926f
C39 minus.n6 a_n1546_n4888# 0.523133f
C40 minus.n7 a_n1546_n4888# 2.11486f
C41 minus.n8 a_n1546_n4888# 0.049176f
C42 minus.t1 a_n1546_n4888# 1.3926f
C43 minus.n9 a_n1546_n4888# 0.528136f
C44 minus.t2 a_n1546_n4888# 1.40292f
C45 minus.n10 a_n1546_n4888# 0.513191f
C46 minus.n11 a_n1546_n4888# 0.162003f
C47 minus.n12 a_n1546_n4888# 0.011159f
C48 minus.t6 a_n1546_n4888# 1.3926f
C49 minus.n13 a_n1546_n4888# 0.528136f
C50 minus.t4 a_n1546_n4888# 1.3926f
C51 minus.n14 a_n1546_n4888# 0.523133f
C52 minus.n15 a_n1546_n4888# 0.332476f
C53 minus.n16 a_n1546_n4888# 2.52908f
C54 drain_left.t5 a_n1546_n4888# 0.46436f
C55 drain_left.t2 a_n1546_n4888# 0.46436f
C56 drain_left.n0 a_n1546_n4888# 4.24708f
C57 drain_left.t6 a_n1546_n4888# 0.46436f
C58 drain_left.t7 a_n1546_n4888# 0.46436f
C59 drain_left.n1 a_n1546_n4888# 4.24708f
C60 drain_left.n2 a_n1546_n4888# 2.65203f
C61 drain_left.t4 a_n1546_n4888# 0.46436f
C62 drain_left.t1 a_n1546_n4888# 0.46436f
C63 drain_left.n3 a_n1546_n4888# 4.24994f
C64 drain_left.t0 a_n1546_n4888# 0.46436f
C65 drain_left.t3 a_n1546_n4888# 0.46436f
C66 drain_left.n4 a_n1546_n4888# 4.24527f
C67 drain_left.n5 a_n1546_n4888# 1.02643f
C68 source.t10 a_n1546_n4888# 3.71779f
C69 source.n0 a_n1546_n4888# 1.59932f
C70 source.t13 a_n1546_n4888# 0.325312f
C71 source.t8 a_n1546_n4888# 0.325312f
C72 source.n1 a_n1546_n4888# 2.90843f
C73 source.n2 a_n1546_n4888# 0.306275f
C74 source.t7 a_n1546_n4888# 3.7178f
C75 source.n3 a_n1546_n4888# 0.367826f
C76 source.t4 a_n1546_n4888# 3.7178f
C77 source.n4 a_n1546_n4888# 0.367826f
C78 source.t0 a_n1546_n4888# 0.325312f
C79 source.t1 a_n1546_n4888# 0.325312f
C80 source.n5 a_n1546_n4888# 2.90843f
C81 source.n6 a_n1546_n4888# 0.306275f
C82 source.t5 a_n1546_n4888# 3.7178f
C83 source.n7 a_n1546_n4888# 1.96893f
C84 source.t11 a_n1546_n4888# 3.71778f
C85 source.n8 a_n1546_n4888# 1.96895f
C86 source.t14 a_n1546_n4888# 0.325312f
C87 source.t12 a_n1546_n4888# 0.325312f
C88 source.n9 a_n1546_n4888# 2.90843f
C89 source.n10 a_n1546_n4888# 0.306269f
C90 source.t9 a_n1546_n4888# 3.71778f
C91 source.n11 a_n1546_n4888# 0.367846f
C92 source.t3 a_n1546_n4888# 3.71778f
C93 source.n12 a_n1546_n4888# 0.367846f
C94 source.t2 a_n1546_n4888# 0.325312f
C95 source.t6 a_n1546_n4888# 0.325312f
C96 source.n13 a_n1546_n4888# 2.90843f
C97 source.n14 a_n1546_n4888# 0.306269f
C98 source.t15 a_n1546_n4888# 3.71778f
C99 source.n15 a_n1546_n4888# 0.493127f
C100 source.n16 a_n1546_n4888# 1.86008f
C101 plus.n0 a_n1546_n4888# 0.049887f
C102 plus.t4 a_n1546_n4888# 1.41274f
C103 plus.t7 a_n1546_n4888# 1.41274f
C104 plus.t6 a_n1546_n4888# 1.41274f
C105 plus.n1 a_n1546_n4888# 0.535776f
C106 plus.t3 a_n1546_n4888# 1.42321f
C107 plus.n2 a_n1546_n4888# 0.520614f
C108 plus.n3 a_n1546_n4888# 0.164347f
C109 plus.n4 a_n1546_n4888# 0.01132f
C110 plus.n5 a_n1546_n4888# 0.535776f
C111 plus.n6 a_n1546_n4888# 0.530701f
C112 plus.n7 a_n1546_n4888# 0.768402f
C113 plus.n8 a_n1546_n4888# 0.049887f
C114 plus.t2 a_n1546_n4888# 1.41274f
C115 plus.t5 a_n1546_n4888# 1.41274f
C116 plus.t1 a_n1546_n4888# 1.41274f
C117 plus.n9 a_n1546_n4888# 0.535776f
C118 plus.t0 a_n1546_n4888# 1.42321f
C119 plus.n10 a_n1546_n4888# 0.520614f
C120 plus.n11 a_n1546_n4888# 0.164347f
C121 plus.n12 a_n1546_n4888# 0.01132f
C122 plus.n13 a_n1546_n4888# 0.535776f
C123 plus.n14 a_n1546_n4888# 0.530701f
C124 plus.n15 a_n1546_n4888# 1.69188f
.ends

