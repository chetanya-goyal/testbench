* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t16 plus.t0 drain_left.t9 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 source.t15 plus.t1 drain_left.t6 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t7 plus.t2 source.t14 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t0 minus.t0 drain_right.t9 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 source.t5 minus.t1 drain_right.t8 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X5 source.t13 plus.t3 drain_left.t4 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X6 drain_left.t8 plus.t4 source.t12 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X7 source.t18 minus.t2 drain_right.t7 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X8 source.t19 minus.t3 drain_right.t6 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X9 drain_right.t5 minus.t4 source.t3 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X10 drain_left.t0 plus.t5 source.t11 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X11 drain_left.t5 plus.t6 source.t10 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X13 a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X14 drain_right.t4 minus.t5 source.t2 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X15 drain_right.t3 minus.t6 source.t6 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X16 drain_right.t2 minus.t7 source.t1 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X17 drain_right.t1 minus.t8 source.t4 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X18 source.t9 plus.t7 drain_left.t2 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X19 drain_right.t0 minus.t9 source.t17 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X20 a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X21 a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X22 drain_left.t1 plus.t8 source.t8 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X23 drain_left.t3 plus.t9 source.t7 a_n1412_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
R0 plus.n2 plus.t4 378.005
R1 plus.n8 plus.t5 378.005
R2 plus.n12 plus.t9 378.005
R3 plus.n18 plus.t8 378.005
R4 plus.n1 plus.t1 318.12
R5 plus.n5 plus.t6 318.12
R6 plus.n7 plus.t0 318.12
R7 plus.n11 plus.t7 318.12
R8 plus.n15 plus.t2 318.12
R9 plus.n17 plus.t3 318.12
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus.n2 plus.n1 24.8308
R27 plus.n8 plus.n7 24.8308
R28 plus.n18 plus.n17 24.8308
R29 plus.n12 plus.n11 24.8308
R30 plus plus.n19 24.5786
R31 plus plus.n9 8.37171
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n2 drain_left.n0 289.615
R37 drain_left.n13 drain_left.n11 289.615
R38 drain_left.n3 drain_left.n2 185
R39 drain_left.n14 drain_left.n13 185
R40 drain_left.t1 drain_left.n1 167.117
R41 drain_left.t8 drain_left.n12 167.117
R42 drain_left.n10 drain_left.n9 101.115
R43 drain_left.n21 drain_left.n20 100.796
R44 drain_left.n19 drain_left.n18 100.796
R45 drain_left.n8 drain_left.n7 100.796
R46 drain_left.n2 drain_left.t1 52.3082
R47 drain_left.n13 drain_left.t8 52.3082
R48 drain_left.n8 drain_left.n6 48.5884
R49 drain_left.n19 drain_left.n17 48.5884
R50 drain_left drain_left.n10 21.9163
R51 drain_left.n9 drain_left.t2 9.9005
R52 drain_left.n9 drain_left.t3 9.9005
R53 drain_left.n7 drain_left.t4 9.9005
R54 drain_left.n7 drain_left.t7 9.9005
R55 drain_left.n20 drain_left.t9 9.9005
R56 drain_left.n20 drain_left.t0 9.9005
R57 drain_left.n18 drain_left.t6 9.9005
R58 drain_left.n18 drain_left.t5 9.9005
R59 drain_left.n3 drain_left.n1 9.71174
R60 drain_left.n14 drain_left.n12 9.71174
R61 drain_left.n6 drain_left.n5 9.45567
R62 drain_left.n17 drain_left.n16 9.45567
R63 drain_left.n5 drain_left.n4 9.3005
R64 drain_left.n16 drain_left.n15 9.3005
R65 drain_left.n6 drain_left.n0 8.14595
R66 drain_left.n17 drain_left.n11 8.14595
R67 drain_left.n4 drain_left.n3 7.3702
R68 drain_left.n15 drain_left.n14 7.3702
R69 drain_left drain_left.n21 6.15322
R70 drain_left.n4 drain_left.n0 5.81868
R71 drain_left.n15 drain_left.n11 5.81868
R72 drain_left.n5 drain_left.n1 3.44771
R73 drain_left.n16 drain_left.n12 3.44771
R74 drain_left.n21 drain_left.n19 0.5005
R75 drain_left.n10 drain_left.n8 0.070154
R76 source.n42 source.n40 289.615
R77 source.n30 source.n28 289.615
R78 source.n2 source.n0 289.615
R79 source.n14 source.n12 289.615
R80 source.n43 source.n42 185
R81 source.n31 source.n30 185
R82 source.n3 source.n2 185
R83 source.n15 source.n14 185
R84 source.t2 source.n41 167.117
R85 source.t7 source.n29 167.117
R86 source.t11 source.n1 167.117
R87 source.t4 source.n13 167.117
R88 source.n9 source.n8 84.1169
R89 source.n11 source.n10 84.1169
R90 source.n21 source.n20 84.1169
R91 source.n23 source.n22 84.1169
R92 source.n39 source.n38 84.1168
R93 source.n37 source.n36 84.1168
R94 source.n27 source.n26 84.1168
R95 source.n25 source.n24 84.1168
R96 source.n42 source.t2 52.3082
R97 source.n30 source.t7 52.3082
R98 source.n2 source.t11 52.3082
R99 source.n14 source.t4 52.3082
R100 source.n47 source.n46 31.4096
R101 source.n35 source.n34 31.4096
R102 source.n7 source.n6 31.4096
R103 source.n19 source.n18 31.4096
R104 source.n25 source.n23 14.712
R105 source.n38 source.t3 9.9005
R106 source.n38 source.t19 9.9005
R107 source.n36 source.t6 9.9005
R108 source.n36 source.t18 9.9005
R109 source.n26 source.t14 9.9005
R110 source.n26 source.t9 9.9005
R111 source.n24 source.t8 9.9005
R112 source.n24 source.t13 9.9005
R113 source.n8 source.t10 9.9005
R114 source.n8 source.t16 9.9005
R115 source.n10 source.t12 9.9005
R116 source.n10 source.t15 9.9005
R117 source.n20 source.t1 9.9005
R118 source.n20 source.t5 9.9005
R119 source.n22 source.t17 9.9005
R120 source.n22 source.t0 9.9005
R121 source.n43 source.n41 9.71174
R122 source.n31 source.n29 9.71174
R123 source.n3 source.n1 9.71174
R124 source.n15 source.n13 9.71174
R125 source.n46 source.n45 9.45567
R126 source.n34 source.n33 9.45567
R127 source.n6 source.n5 9.45567
R128 source.n18 source.n17 9.45567
R129 source.n45 source.n44 9.3005
R130 source.n33 source.n32 9.3005
R131 source.n5 source.n4 9.3005
R132 source.n17 source.n16 9.3005
R133 source.n48 source.n7 8.69904
R134 source.n46 source.n40 8.14595
R135 source.n34 source.n28 8.14595
R136 source.n6 source.n0 8.14595
R137 source.n18 source.n12 8.14595
R138 source.n44 source.n43 7.3702
R139 source.n32 source.n31 7.3702
R140 source.n4 source.n3 7.3702
R141 source.n16 source.n15 7.3702
R142 source.n44 source.n40 5.81868
R143 source.n32 source.n28 5.81868
R144 source.n4 source.n0 5.81868
R145 source.n16 source.n12 5.81868
R146 source.n48 source.n47 5.51343
R147 source.n45 source.n41 3.44771
R148 source.n33 source.n29 3.44771
R149 source.n5 source.n1 3.44771
R150 source.n17 source.n13 3.44771
R151 source.n19 source.n11 0.720328
R152 source.n37 source.n35 0.720328
R153 source.n23 source.n21 0.5005
R154 source.n21 source.n19 0.5005
R155 source.n11 source.n9 0.5005
R156 source.n9 source.n7 0.5005
R157 source.n27 source.n25 0.5005
R158 source.n35 source.n27 0.5005
R159 source.n39 source.n37 0.5005
R160 source.n47 source.n39 0.5005
R161 source source.n48 0.188
R162 minus.n8 minus.t9 378.005
R163 minus.n2 minus.t8 378.005
R164 minus.n18 minus.t5 378.005
R165 minus.n12 minus.t6 378.005
R166 minus.n7 minus.t0 318.12
R167 minus.n5 minus.t7 318.12
R168 minus.n1 minus.t1 318.12
R169 minus.n17 minus.t3 318.12
R170 minus.n15 minus.t4 318.12
R171 minus.n11 minus.t2 318.12
R172 minus.n3 minus.n2 161.489
R173 minus.n13 minus.n12 161.489
R174 minus.n9 minus.n8 161.3
R175 minus.n6 minus.n0 161.3
R176 minus.n4 minus.n3 161.3
R177 minus.n19 minus.n18 161.3
R178 minus.n16 minus.n10 161.3
R179 minus.n14 minus.n13 161.3
R180 minus.n7 minus.n6 48.2005
R181 minus.n4 minus.n1 48.2005
R182 minus.n14 minus.n11 48.2005
R183 minus.n17 minus.n16 48.2005
R184 minus.n6 minus.n5 36.5157
R185 minus.n5 minus.n4 36.5157
R186 minus.n15 minus.n14 36.5157
R187 minus.n16 minus.n15 36.5157
R188 minus.n20 minus.n9 26.9096
R189 minus.n8 minus.n7 24.8308
R190 minus.n2 minus.n1 24.8308
R191 minus.n12 minus.n11 24.8308
R192 minus.n18 minus.n17 24.8308
R193 minus.n20 minus.n19 6.51565
R194 minus.n9 minus.n0 0.189894
R195 minus.n3 minus.n0 0.189894
R196 minus.n13 minus.n10 0.189894
R197 minus.n19 minus.n10 0.189894
R198 minus minus.n20 0.188
R199 drain_right.n2 drain_right.n0 289.615
R200 drain_right.n16 drain_right.n14 289.615
R201 drain_right.n3 drain_right.n2 185
R202 drain_right.n17 drain_right.n16 185
R203 drain_right.t3 drain_right.n1 167.117
R204 drain_right.t0 drain_right.n15 167.117
R205 drain_right.n13 drain_right.n11 101.296
R206 drain_right.n10 drain_right.n9 101.115
R207 drain_right.n13 drain_right.n12 100.796
R208 drain_right.n8 drain_right.n7 100.796
R209 drain_right.n2 drain_right.t3 52.3082
R210 drain_right.n16 drain_right.t0 52.3082
R211 drain_right.n8 drain_right.n6 48.5884
R212 drain_right.n21 drain_right.n20 48.0884
R213 drain_right drain_right.n10 21.3631
R214 drain_right.n9 drain_right.t6 9.9005
R215 drain_right.n9 drain_right.t4 9.9005
R216 drain_right.n7 drain_right.t7 9.9005
R217 drain_right.n7 drain_right.t5 9.9005
R218 drain_right.n11 drain_right.t8 9.9005
R219 drain_right.n11 drain_right.t1 9.9005
R220 drain_right.n12 drain_right.t9 9.9005
R221 drain_right.n12 drain_right.t2 9.9005
R222 drain_right.n3 drain_right.n1 9.71174
R223 drain_right.n17 drain_right.n15 9.71174
R224 drain_right.n6 drain_right.n5 9.45567
R225 drain_right.n20 drain_right.n19 9.45567
R226 drain_right.n5 drain_right.n4 9.3005
R227 drain_right.n19 drain_right.n18 9.3005
R228 drain_right.n6 drain_right.n0 8.14595
R229 drain_right.n20 drain_right.n14 8.14595
R230 drain_right.n4 drain_right.n3 7.3702
R231 drain_right.n18 drain_right.n17 7.3702
R232 drain_right drain_right.n21 5.90322
R233 drain_right.n4 drain_right.n0 5.81868
R234 drain_right.n18 drain_right.n14 5.81868
R235 drain_right.n5 drain_right.n1 3.44771
R236 drain_right.n19 drain_right.n15 3.44771
R237 drain_right.n21 drain_right.n13 0.5005
R238 drain_right.n10 drain_right.n8 0.070154
C0 source drain_left 5.55091f
C1 plus drain_right 0.295235f
C2 minus drain_left 0.177288f
C3 minus source 1.00561f
C4 plus drain_left 1.04711f
C5 plus source 1.01968f
C6 drain_right drain_left 0.689799f
C7 drain_right source 5.54759f
C8 plus minus 3.06588f
C9 drain_right minus 0.913449f
C10 drain_right a_n1412_n1288# 3.49646f
C11 drain_left a_n1412_n1288# 3.7229f
C12 source a_n1412_n1288# 2.404181f
C13 minus a_n1412_n1288# 4.645155f
C14 plus a_n1412_n1288# 5.348974f
C15 drain_right.n0 a_n1412_n1288# 0.036188f
C16 drain_right.n1 a_n1412_n1288# 0.080071f
C17 drain_right.t3 a_n1412_n1288# 0.06009f
C18 drain_right.n2 a_n1412_n1288# 0.062667f
C19 drain_right.n3 a_n1412_n1288# 0.020201f
C20 drain_right.n4 a_n1412_n1288# 0.013323f
C21 drain_right.n5 a_n1412_n1288# 0.176497f
C22 drain_right.n6 a_n1412_n1288# 0.057696f
C23 drain_right.t7 a_n1412_n1288# 0.039186f
C24 drain_right.t5 a_n1412_n1288# 0.039186f
C25 drain_right.n7 a_n1412_n1288# 0.246178f
C26 drain_right.n8 a_n1412_n1288# 0.329553f
C27 drain_right.t6 a_n1412_n1288# 0.039186f
C28 drain_right.t4 a_n1412_n1288# 0.039186f
C29 drain_right.n9 a_n1412_n1288# 0.247023f
C30 drain_right.n10 a_n1412_n1288# 0.812082f
C31 drain_right.t8 a_n1412_n1288# 0.039186f
C32 drain_right.t1 a_n1412_n1288# 0.039186f
C33 drain_right.n11 a_n1412_n1288# 0.24756f
C34 drain_right.t9 a_n1412_n1288# 0.039186f
C35 drain_right.t2 a_n1412_n1288# 0.039186f
C36 drain_right.n12 a_n1412_n1288# 0.246179f
C37 drain_right.n13 a_n1412_n1288# 0.547931f
C38 drain_right.n14 a_n1412_n1288# 0.036188f
C39 drain_right.n15 a_n1412_n1288# 0.080071f
C40 drain_right.t0 a_n1412_n1288# 0.06009f
C41 drain_right.n16 a_n1412_n1288# 0.062667f
C42 drain_right.n17 a_n1412_n1288# 0.020201f
C43 drain_right.n18 a_n1412_n1288# 0.013323f
C44 drain_right.n19 a_n1412_n1288# 0.176497f
C45 drain_right.n20 a_n1412_n1288# 0.056802f
C46 drain_right.n21 a_n1412_n1288# 0.291098f
C47 minus.n0 a_n1412_n1288# 0.034088f
C48 minus.t9 a_n1412_n1288# 0.056513f
C49 minus.t0 a_n1412_n1288# 0.050154f
C50 minus.t7 a_n1412_n1288# 0.050154f
C51 minus.t1 a_n1412_n1288# 0.050154f
C52 minus.n1 a_n1412_n1288# 0.036779f
C53 minus.t8 a_n1412_n1288# 0.056513f
C54 minus.n2 a_n1412_n1288# 0.046826f
C55 minus.n3 a_n1412_n1288# 0.080102f
C56 minus.n4 a_n1412_n1288# 0.012989f
C57 minus.n5 a_n1412_n1288# 0.036779f
C58 minus.n6 a_n1412_n1288# 0.012989f
C59 minus.n7 a_n1412_n1288# 0.036779f
C60 minus.n8 a_n1412_n1288# 0.046772f
C61 minus.n9 a_n1412_n1288# 0.733122f
C62 minus.n10 a_n1412_n1288# 0.034088f
C63 minus.t3 a_n1412_n1288# 0.050154f
C64 minus.t4 a_n1412_n1288# 0.050154f
C65 minus.t2 a_n1412_n1288# 0.050154f
C66 minus.n11 a_n1412_n1288# 0.036779f
C67 minus.t6 a_n1412_n1288# 0.056513f
C68 minus.n12 a_n1412_n1288# 0.046826f
C69 minus.n13 a_n1412_n1288# 0.080102f
C70 minus.n14 a_n1412_n1288# 0.012989f
C71 minus.n15 a_n1412_n1288# 0.036779f
C72 minus.n16 a_n1412_n1288# 0.012989f
C73 minus.n17 a_n1412_n1288# 0.036779f
C74 minus.t5 a_n1412_n1288# 0.056513f
C75 minus.n18 a_n1412_n1288# 0.046772f
C76 minus.n19 a_n1412_n1288# 0.224115f
C77 minus.n20 a_n1412_n1288# 0.905193f
C78 source.n0 a_n1412_n1288# 0.044421f
C79 source.n1 a_n1412_n1288# 0.098286f
C80 source.t11 a_n1412_n1288# 0.073758f
C81 source.n2 a_n1412_n1288# 0.076922f
C82 source.n3 a_n1412_n1288# 0.024797f
C83 source.n4 a_n1412_n1288# 0.016354f
C84 source.n5 a_n1412_n1288# 0.216646f
C85 source.n6 a_n1412_n1288# 0.048695f
C86 source.n7 a_n1412_n1288# 0.451992f
C87 source.t10 a_n1412_n1288# 0.0481f
C88 source.t16 a_n1412_n1288# 0.0481f
C89 source.n8 a_n1412_n1288# 0.257141f
C90 source.n9 a_n1412_n1288# 0.334677f
C91 source.t12 a_n1412_n1288# 0.0481f
C92 source.t15 a_n1412_n1288# 0.0481f
C93 source.n10 a_n1412_n1288# 0.257141f
C94 source.n11 a_n1412_n1288# 0.356235f
C95 source.n12 a_n1412_n1288# 0.044421f
C96 source.n13 a_n1412_n1288# 0.098286f
C97 source.t4 a_n1412_n1288# 0.073758f
C98 source.n14 a_n1412_n1288# 0.076922f
C99 source.n15 a_n1412_n1288# 0.024797f
C100 source.n16 a_n1412_n1288# 0.016354f
C101 source.n17 a_n1412_n1288# 0.216646f
C102 source.n18 a_n1412_n1288# 0.048695f
C103 source.n19 a_n1412_n1288# 0.144678f
C104 source.t1 a_n1412_n1288# 0.0481f
C105 source.t5 a_n1412_n1288# 0.0481f
C106 source.n20 a_n1412_n1288# 0.257141f
C107 source.n21 a_n1412_n1288# 0.334677f
C108 source.t17 a_n1412_n1288# 0.0481f
C109 source.t0 a_n1412_n1288# 0.0481f
C110 source.n22 a_n1412_n1288# 0.257141f
C111 source.n23 a_n1412_n1288# 0.99538f
C112 source.t8 a_n1412_n1288# 0.0481f
C113 source.t13 a_n1412_n1288# 0.0481f
C114 source.n24 a_n1412_n1288# 0.25714f
C115 source.n25 a_n1412_n1288# 0.995382f
C116 source.t14 a_n1412_n1288# 0.0481f
C117 source.t9 a_n1412_n1288# 0.0481f
C118 source.n26 a_n1412_n1288# 0.25714f
C119 source.n27 a_n1412_n1288# 0.334679f
C120 source.n28 a_n1412_n1288# 0.044421f
C121 source.n29 a_n1412_n1288# 0.098286f
C122 source.t7 a_n1412_n1288# 0.073758f
C123 source.n30 a_n1412_n1288# 0.076922f
C124 source.n31 a_n1412_n1288# 0.024797f
C125 source.n32 a_n1412_n1288# 0.016354f
C126 source.n33 a_n1412_n1288# 0.216646f
C127 source.n34 a_n1412_n1288# 0.048695f
C128 source.n35 a_n1412_n1288# 0.144678f
C129 source.t6 a_n1412_n1288# 0.0481f
C130 source.t18 a_n1412_n1288# 0.0481f
C131 source.n36 a_n1412_n1288# 0.25714f
C132 source.n37 a_n1412_n1288# 0.356236f
C133 source.t3 a_n1412_n1288# 0.0481f
C134 source.t19 a_n1412_n1288# 0.0481f
C135 source.n38 a_n1412_n1288# 0.25714f
C136 source.n39 a_n1412_n1288# 0.334679f
C137 source.n40 a_n1412_n1288# 0.044421f
C138 source.n41 a_n1412_n1288# 0.098286f
C139 source.t2 a_n1412_n1288# 0.073758f
C140 source.n42 a_n1412_n1288# 0.076922f
C141 source.n43 a_n1412_n1288# 0.024797f
C142 source.n44 a_n1412_n1288# 0.016354f
C143 source.n45 a_n1412_n1288# 0.216646f
C144 source.n46 a_n1412_n1288# 0.048695f
C145 source.n47 a_n1412_n1288# 0.288578f
C146 source.n48 a_n1412_n1288# 0.750659f
C147 drain_left.n0 a_n1412_n1288# 0.036208f
C148 drain_left.n1 a_n1412_n1288# 0.080114f
C149 drain_left.t1 a_n1412_n1288# 0.060122f
C150 drain_left.n2 a_n1412_n1288# 0.062701f
C151 drain_left.n3 a_n1412_n1288# 0.020212f
C152 drain_left.n4 a_n1412_n1288# 0.01333f
C153 drain_left.n5 a_n1412_n1288# 0.176592f
C154 drain_left.n6 a_n1412_n1288# 0.057727f
C155 drain_left.t4 a_n1412_n1288# 0.039207f
C156 drain_left.t7 a_n1412_n1288# 0.039207f
C157 drain_left.n7 a_n1412_n1288# 0.246311f
C158 drain_left.n8 a_n1412_n1288# 0.329731f
C159 drain_left.t2 a_n1412_n1288# 0.039207f
C160 drain_left.t3 a_n1412_n1288# 0.039207f
C161 drain_left.n9 a_n1412_n1288# 0.247155f
C162 drain_left.n10 a_n1412_n1288# 0.86133f
C163 drain_left.n11 a_n1412_n1288# 0.036208f
C164 drain_left.n12 a_n1412_n1288# 0.080114f
C165 drain_left.t8 a_n1412_n1288# 0.060122f
C166 drain_left.n13 a_n1412_n1288# 0.062701f
C167 drain_left.n14 a_n1412_n1288# 0.020212f
C168 drain_left.n15 a_n1412_n1288# 0.01333f
C169 drain_left.n16 a_n1412_n1288# 0.176592f
C170 drain_left.n17 a_n1412_n1288# 0.057727f
C171 drain_left.t6 a_n1412_n1288# 0.039207f
C172 drain_left.t5 a_n1412_n1288# 0.039207f
C173 drain_left.n18 a_n1412_n1288# 0.246312f
C174 drain_left.n19 a_n1412_n1288# 0.355872f
C175 drain_left.t9 a_n1412_n1288# 0.039207f
C176 drain_left.t0 a_n1412_n1288# 0.039207f
C177 drain_left.n20 a_n1412_n1288# 0.246312f
C178 drain_left.n21 a_n1412_n1288# 0.474575f
C179 plus.n0 a_n1412_n1288# 0.034863f
C180 plus.t0 a_n1412_n1288# 0.051294f
C181 plus.t6 a_n1412_n1288# 0.051294f
C182 plus.t1 a_n1412_n1288# 0.051294f
C183 plus.n1 a_n1412_n1288# 0.037616f
C184 plus.t4 a_n1412_n1288# 0.057798f
C185 plus.n2 a_n1412_n1288# 0.047891f
C186 plus.n3 a_n1412_n1288# 0.081923f
C187 plus.n4 a_n1412_n1288# 0.013285f
C188 plus.n5 a_n1412_n1288# 0.037616f
C189 plus.n6 a_n1412_n1288# 0.013285f
C190 plus.n7 a_n1412_n1288# 0.037616f
C191 plus.t5 a_n1412_n1288# 0.057798f
C192 plus.n8 a_n1412_n1288# 0.047836f
C193 plus.n9 a_n1412_n1288# 0.250589f
C194 plus.n10 a_n1412_n1288# 0.034863f
C195 plus.t8 a_n1412_n1288# 0.057798f
C196 plus.t3 a_n1412_n1288# 0.051294f
C197 plus.t2 a_n1412_n1288# 0.051294f
C198 plus.t7 a_n1412_n1288# 0.051294f
C199 plus.n11 a_n1412_n1288# 0.037616f
C200 plus.t9 a_n1412_n1288# 0.057798f
C201 plus.n12 a_n1412_n1288# 0.047891f
C202 plus.n13 a_n1412_n1288# 0.081923f
C203 plus.n14 a_n1412_n1288# 0.013285f
C204 plus.n15 a_n1412_n1288# 0.037616f
C205 plus.n16 a_n1412_n1288# 0.013285f
C206 plus.n17 a_n1412_n1288# 0.037616f
C207 plus.n18 a_n1412_n1288# 0.047836f
C208 plus.n19 a_n1412_n1288# 0.719386f
.ends

