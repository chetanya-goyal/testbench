* NGSPICE file created from diffpair624.ext - technology: sky130A

.subckt diffpair624 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t8 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 drain_right.t9 minus.t0 source.t1 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X2 source.t11 plus.t1 drain_left.t8 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t18 minus.t1 drain_right.t8 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 drain_left.t7 plus.t2 source.t10 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X5 source.t4 minus.t2 drain_right.t7 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X7 a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X8 drain_right.t6 minus.t3 source.t0 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X9 a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X10 drain_left.t6 plus.t3 source.t15 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X11 drain_left.t5 plus.t4 source.t9 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X12 source.t19 minus.t4 drain_right.t5 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X13 drain_right.t4 minus.t5 source.t2 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X14 drain_right.t3 minus.t6 source.t7 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X15 a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X16 drain_right.t2 minus.t7 source.t6 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X17 source.t14 plus.t5 drain_left.t4 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X18 source.t12 plus.t6 drain_left.t3 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 drain_left.t2 plus.t7 source.t13 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X20 drain_right.t1 minus.t8 source.t3 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X21 source.t17 plus.t8 drain_left.t1 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X22 drain_left.t0 plus.t9 source.t16 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 source.t5 minus.t9 drain_right.t0 a_n1952_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n3 plus.t4 767.438
R1 plus.n17 plus.t0 767.438
R2 plus.n12 plus.t3 744.691
R3 plus.n10 plus.t5 744.691
R4 plus.n2 plus.t2 744.691
R5 plus.n4 plus.t8 744.691
R6 plus.n26 plus.t7 744.691
R7 plus.n24 plus.t6 744.691
R8 plus.n16 plus.t9 744.691
R9 plus.n18 plus.t1 744.691
R10 plus.n6 plus.n5 161.3
R11 plus.n7 plus.n2 161.3
R12 plus.n9 plus.n8 161.3
R13 plus.n10 plus.n1 161.3
R14 plus.n11 plus.n0 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n20 plus.n19 161.3
R17 plus.n21 plus.n16 161.3
R18 plus.n23 plus.n22 161.3
R19 plus.n24 plus.n15 161.3
R20 plus.n25 plus.n14 161.3
R21 plus.n27 plus.n26 161.3
R22 plus.n6 plus.n3 44.8741
R23 plus.n20 plus.n17 44.8741
R24 plus plus.n27 33.5653
R25 plus.n12 plus.n11 30.6732
R26 plus.n26 plus.n25 30.6732
R27 plus.n10 plus.n9 26.2914
R28 plus.n5 plus.n4 26.2914
R29 plus.n24 plus.n23 26.2914
R30 plus.n19 plus.n18 26.2914
R31 plus.n9 plus.n2 21.9096
R32 plus.n5 plus.n2 21.9096
R33 plus.n23 plus.n16 21.9096
R34 plus.n19 plus.n16 21.9096
R35 plus.n4 plus.n3 19.0667
R36 plus.n18 plus.n17 19.0667
R37 plus.n11 plus.n10 17.5278
R38 plus.n25 plus.n24 17.5278
R39 plus plus.n13 15.313
R40 plus.n7 plus.n6 0.189894
R41 plus.n8 plus.n7 0.189894
R42 plus.n8 plus.n1 0.189894
R43 plus.n1 plus.n0 0.189894
R44 plus.n13 plus.n0 0.189894
R45 plus.n27 plus.n14 0.189894
R46 plus.n15 plus.n14 0.189894
R47 plus.n22 plus.n15 0.189894
R48 plus.n22 plus.n21 0.189894
R49 plus.n21 plus.n20 0.189894
R50 source.n0 source.t15 44.1297
R51 source.n5 source.t3 44.1296
R52 source.n19 source.t0 44.1295
R53 source.n14 source.t8 44.1295
R54 source.n2 source.n1 43.1397
R55 source.n4 source.n3 43.1397
R56 source.n7 source.n6 43.1397
R57 source.n9 source.n8 43.1397
R58 source.n18 source.n17 43.1396
R59 source.n16 source.n15 43.1396
R60 source.n13 source.n12 43.1396
R61 source.n11 source.n10 43.1396
R62 source.n11 source.n9 29.1242
R63 source.n20 source.n0 22.5294
R64 source.n20 source.n19 5.7074
R65 source.n17 source.t1 0.9905
R66 source.n17 source.t18 0.9905
R67 source.n15 source.t2 0.9905
R68 source.n15 source.t19 0.9905
R69 source.n12 source.t16 0.9905
R70 source.n12 source.t11 0.9905
R71 source.n10 source.t13 0.9905
R72 source.n10 source.t12 0.9905
R73 source.n1 source.t10 0.9905
R74 source.n1 source.t14 0.9905
R75 source.n3 source.t9 0.9905
R76 source.n3 source.t17 0.9905
R77 source.n6 source.t6 0.9905
R78 source.n6 source.t4 0.9905
R79 source.n8 source.t7 0.9905
R80 source.n8 source.t5 0.9905
R81 source.n5 source.n4 0.914293
R82 source.n16 source.n14 0.914293
R83 source.n9 source.n7 0.888431
R84 source.n7 source.n5 0.888431
R85 source.n4 source.n2 0.888431
R86 source.n2 source.n0 0.888431
R87 source.n13 source.n11 0.888431
R88 source.n14 source.n13 0.888431
R89 source.n18 source.n16 0.888431
R90 source.n19 source.n18 0.888431
R91 source source.n20 0.188
R92 drain_left.n5 drain_left.t5 61.6963
R93 drain_left.n1 drain_left.t2 61.6962
R94 drain_left.n3 drain_left.n2 60.429
R95 drain_left.n7 drain_left.n6 59.8185
R96 drain_left.n5 drain_left.n4 59.8185
R97 drain_left.n1 drain_left.n0 59.8184
R98 drain_left drain_left.n3 37.2014
R99 drain_left drain_left.n7 6.54115
R100 drain_left.n2 drain_left.t8 0.9905
R101 drain_left.n2 drain_left.t9 0.9905
R102 drain_left.n0 drain_left.t3 0.9905
R103 drain_left.n0 drain_left.t0 0.9905
R104 drain_left.n6 drain_left.t4 0.9905
R105 drain_left.n6 drain_left.t6 0.9905
R106 drain_left.n4 drain_left.t1 0.9905
R107 drain_left.n4 drain_left.t7 0.9905
R108 drain_left.n7 drain_left.n5 0.888431
R109 drain_left.n3 drain_left.n1 0.167137
R110 minus.n3 minus.t8 767.438
R111 minus.n17 minus.t5 767.438
R112 minus.n4 minus.t2 744.691
R113 minus.n6 minus.t7 744.691
R114 minus.n10 minus.t9 744.691
R115 minus.n12 minus.t6 744.691
R116 minus.n18 minus.t4 744.691
R117 minus.n20 minus.t0 744.691
R118 minus.n24 minus.t1 744.691
R119 minus.n26 minus.t3 744.691
R120 minus.n13 minus.n12 161.3
R121 minus.n11 minus.n0 161.3
R122 minus.n10 minus.n9 161.3
R123 minus.n8 minus.n1 161.3
R124 minus.n7 minus.n6 161.3
R125 minus.n5 minus.n2 161.3
R126 minus.n27 minus.n26 161.3
R127 minus.n25 minus.n14 161.3
R128 minus.n24 minus.n23 161.3
R129 minus.n22 minus.n15 161.3
R130 minus.n21 minus.n20 161.3
R131 minus.n19 minus.n16 161.3
R132 minus.n3 minus.n2 44.8741
R133 minus.n17 minus.n16 44.8741
R134 minus.n28 minus.n13 42.7145
R135 minus.n12 minus.n11 30.6732
R136 minus.n26 minus.n25 30.6732
R137 minus.n5 minus.n4 26.2914
R138 minus.n10 minus.n1 26.2914
R139 minus.n19 minus.n18 26.2914
R140 minus.n24 minus.n15 26.2914
R141 minus.n6 minus.n5 21.9096
R142 minus.n6 minus.n1 21.9096
R143 minus.n20 minus.n19 21.9096
R144 minus.n20 minus.n15 21.9096
R145 minus.n4 minus.n3 19.0667
R146 minus.n18 minus.n17 19.0667
R147 minus.n11 minus.n10 17.5278
R148 minus.n25 minus.n24 17.5278
R149 minus.n28 minus.n27 6.63876
R150 minus.n13 minus.n0 0.189894
R151 minus.n9 minus.n0 0.189894
R152 minus.n9 minus.n8 0.189894
R153 minus.n8 minus.n7 0.189894
R154 minus.n7 minus.n2 0.189894
R155 minus.n21 minus.n16 0.189894
R156 minus.n22 minus.n21 0.189894
R157 minus.n23 minus.n22 0.189894
R158 minus.n23 minus.n14 0.189894
R159 minus.n27 minus.n14 0.189894
R160 minus minus.n28 0.188
R161 drain_right.n1 drain_right.t4 61.6962
R162 drain_right.n7 drain_right.t3 60.8084
R163 drain_right.n6 drain_right.n4 60.7064
R164 drain_right.n3 drain_right.n2 60.429
R165 drain_right.n6 drain_right.n5 59.8185
R166 drain_right.n1 drain_right.n0 59.8184
R167 drain_right drain_right.n3 36.6482
R168 drain_right drain_right.n7 6.09718
R169 drain_right.n2 drain_right.t8 0.9905
R170 drain_right.n2 drain_right.t6 0.9905
R171 drain_right.n0 drain_right.t5 0.9905
R172 drain_right.n0 drain_right.t9 0.9905
R173 drain_right.n4 drain_right.t7 0.9905
R174 drain_right.n4 drain_right.t1 0.9905
R175 drain_right.n5 drain_right.t0 0.9905
R176 drain_right.n5 drain_right.t2 0.9905
R177 drain_right.n7 drain_right.n6 0.888431
R178 drain_right.n3 drain_right.n1 0.167137
C0 drain_right plus 0.348383f
C1 drain_right drain_left 0.971685f
C2 source minus 10.4122f
C3 minus plus 7.05858f
C4 drain_left minus 0.171897f
C5 source plus 10.427f
C6 source drain_left 22.2255f
C7 drain_left plus 11.080799f
C8 drain_right minus 10.894401f
C9 source drain_right 22.2139f
C10 drain_right a_n1952_n4888# 9.14008f
C11 drain_left a_n1952_n4888# 9.4372f
C12 source a_n1952_n4888# 9.435094f
C13 minus a_n1952_n4888# 8.175349f
C14 plus a_n1952_n4888# 10.287081f
C15 drain_right.t4 a_n1952_n4888# 4.49129f
C16 drain_right.t5 a_n1952_n4888# 0.383684f
C17 drain_right.t9 a_n1952_n4888# 0.383684f
C18 drain_right.n0 a_n1952_n4888# 3.50773f
C19 drain_right.n1 a_n1952_n4888# 0.637677f
C20 drain_right.t8 a_n1952_n4888# 0.383684f
C21 drain_right.t6 a_n1952_n4888# 0.383684f
C22 drain_right.n2 a_n1952_n4888# 3.51109f
C23 drain_right.n3 a_n1952_n4888# 1.99284f
C24 drain_right.t7 a_n1952_n4888# 0.383684f
C25 drain_right.t1 a_n1952_n4888# 0.383684f
C26 drain_right.n4 a_n1952_n4888# 3.51289f
C27 drain_right.t0 a_n1952_n4888# 0.383684f
C28 drain_right.t2 a_n1952_n4888# 0.383684f
C29 drain_right.n5 a_n1952_n4888# 3.50772f
C30 drain_right.n6 a_n1952_n4888# 0.692173f
C31 drain_right.t3 a_n1952_n4888# 4.48624f
C32 drain_right.n7 a_n1952_n4888# 0.575111f
C33 minus.n0 a_n1952_n4888# 0.042424f
C34 minus.n1 a_n1952_n4888# 0.009627f
C35 minus.t9 a_n1952_n4888# 1.68195f
C36 minus.n2 a_n1952_n4888# 0.177195f
C37 minus.t8 a_n1952_n4888# 1.70054f
C38 minus.n3 a_n1952_n4888# 0.612476f
C39 minus.t2 a_n1952_n4888# 1.68195f
C40 minus.n4 a_n1952_n4888# 0.631469f
C41 minus.n5 a_n1952_n4888# 0.009627f
C42 minus.t7 a_n1952_n4888# 1.68195f
C43 minus.n6 a_n1952_n4888# 0.627194f
C44 minus.n7 a_n1952_n4888# 0.042424f
C45 minus.n8 a_n1952_n4888# 0.042424f
C46 minus.n9 a_n1952_n4888# 0.042424f
C47 minus.n10 a_n1952_n4888# 0.627194f
C48 minus.n11 a_n1952_n4888# 0.009627f
C49 minus.t6 a_n1952_n4888# 1.68195f
C50 minus.n12 a_n1952_n4888# 0.62484f
C51 minus.n13 a_n1952_n4888# 1.92974f
C52 minus.n14 a_n1952_n4888# 0.042424f
C53 minus.n15 a_n1952_n4888# 0.009627f
C54 minus.n16 a_n1952_n4888# 0.177195f
C55 minus.t5 a_n1952_n4888# 1.70054f
C56 minus.n17 a_n1952_n4888# 0.612476f
C57 minus.t4 a_n1952_n4888# 1.68195f
C58 minus.n18 a_n1952_n4888# 0.631469f
C59 minus.n19 a_n1952_n4888# 0.009627f
C60 minus.t0 a_n1952_n4888# 1.68195f
C61 minus.n20 a_n1952_n4888# 0.627194f
C62 minus.n21 a_n1952_n4888# 0.042424f
C63 minus.n22 a_n1952_n4888# 0.042424f
C64 minus.n23 a_n1952_n4888# 0.042424f
C65 minus.t1 a_n1952_n4888# 1.68195f
C66 minus.n24 a_n1952_n4888# 0.627194f
C67 minus.n25 a_n1952_n4888# 0.009627f
C68 minus.t3 a_n1952_n4888# 1.68195f
C69 minus.n26 a_n1952_n4888# 0.62484f
C70 minus.n27 a_n1952_n4888# 0.291134f
C71 minus.n28 a_n1952_n4888# 2.29669f
C72 drain_left.t2 a_n1952_n4888# 4.5055f
C73 drain_left.t3 a_n1952_n4888# 0.384898f
C74 drain_left.t0 a_n1952_n4888# 0.384898f
C75 drain_left.n0 a_n1952_n4888# 3.51883f
C76 drain_left.n1 a_n1952_n4888# 0.639695f
C77 drain_left.t8 a_n1952_n4888# 0.384898f
C78 drain_left.t9 a_n1952_n4888# 0.384898f
C79 drain_left.n2 a_n1952_n4888# 3.5222f
C80 drain_left.n3 a_n1952_n4888# 2.04977f
C81 drain_left.t5 a_n1952_n4888# 4.50552f
C82 drain_left.t1 a_n1952_n4888# 0.384898f
C83 drain_left.t7 a_n1952_n4888# 0.384898f
C84 drain_left.n4 a_n1952_n4888# 3.51882f
C85 drain_left.n5 a_n1952_n4888# 0.692896f
C86 drain_left.t4 a_n1952_n4888# 0.384898f
C87 drain_left.t6 a_n1952_n4888# 0.384898f
C88 drain_left.n6 a_n1952_n4888# 3.51882f
C89 drain_left.n7 a_n1952_n4888# 0.560279f
C90 source.t15 a_n1952_n4888# 4.47911f
C91 source.n0 a_n1952_n4888# 1.94854f
C92 source.t10 a_n1952_n4888# 0.391928f
C93 source.t14 a_n1952_n4888# 0.391928f
C94 source.n1 a_n1952_n4888# 3.50401f
C95 source.n2 a_n1952_n4888# 0.396547f
C96 source.t9 a_n1952_n4888# 0.391928f
C97 source.t17 a_n1952_n4888# 0.391928f
C98 source.n3 a_n1952_n4888# 3.50401f
C99 source.n4 a_n1952_n4888# 0.398613f
C100 source.t3 a_n1952_n4888# 4.47912f
C101 source.n5 a_n1952_n4888# 0.4924f
C102 source.t6 a_n1952_n4888# 0.391928f
C103 source.t4 a_n1952_n4888# 0.391928f
C104 source.n6 a_n1952_n4888# 3.50401f
C105 source.n7 a_n1952_n4888# 0.396547f
C106 source.t7 a_n1952_n4888# 0.391928f
C107 source.t5 a_n1952_n4888# 0.391928f
C108 source.n8 a_n1952_n4888# 3.50401f
C109 source.n9 a_n1952_n4888# 2.37684f
C110 source.t13 a_n1952_n4888# 0.391928f
C111 source.t12 a_n1952_n4888# 0.391928f
C112 source.n10 a_n1952_n4888# 3.50401f
C113 source.n11 a_n1952_n4888# 2.37683f
C114 source.t16 a_n1952_n4888# 0.391928f
C115 source.t11 a_n1952_n4888# 0.391928f
C116 source.n12 a_n1952_n4888# 3.50401f
C117 source.n13 a_n1952_n4888# 0.39654f
C118 source.t8 a_n1952_n4888# 4.47909f
C119 source.n14 a_n1952_n4888# 0.492425f
C120 source.t2 a_n1952_n4888# 0.391928f
C121 source.t19 a_n1952_n4888# 0.391928f
C122 source.n15 a_n1952_n4888# 3.50401f
C123 source.n16 a_n1952_n4888# 0.398606f
C124 source.t1 a_n1952_n4888# 0.391928f
C125 source.t18 a_n1952_n4888# 0.391928f
C126 source.n17 a_n1952_n4888# 3.50401f
C127 source.n18 a_n1952_n4888# 0.39654f
C128 source.t0 a_n1952_n4888# 4.47909f
C129 source.n19 a_n1952_n4888# 0.61871f
C130 source.n20 a_n1952_n4888# 2.24978f
C131 plus.n0 a_n1952_n4888# 0.042852f
C132 plus.t3 a_n1952_n4888# 1.69893f
C133 plus.t5 a_n1952_n4888# 1.69893f
C134 plus.n1 a_n1952_n4888# 0.042852f
C135 plus.t2 a_n1952_n4888# 1.69893f
C136 plus.n2 a_n1952_n4888# 0.633525f
C137 plus.t4 a_n1952_n4888# 1.7177f
C138 plus.n3 a_n1952_n4888# 0.618658f
C139 plus.t8 a_n1952_n4888# 1.69893f
C140 plus.n4 a_n1952_n4888# 0.637843f
C141 plus.n5 a_n1952_n4888# 0.009724f
C142 plus.n6 a_n1952_n4888# 0.178984f
C143 plus.n7 a_n1952_n4888# 0.042852f
C144 plus.n8 a_n1952_n4888# 0.042852f
C145 plus.n9 a_n1952_n4888# 0.009724f
C146 plus.n10 a_n1952_n4888# 0.633525f
C147 plus.n11 a_n1952_n4888# 0.009724f
C148 plus.n12 a_n1952_n4888# 0.631147f
C149 plus.n13 a_n1952_n4888# 0.664318f
C150 plus.n14 a_n1952_n4888# 0.042852f
C151 plus.t7 a_n1952_n4888# 1.69893f
C152 plus.n15 a_n1952_n4888# 0.042852f
C153 plus.t6 a_n1952_n4888# 1.69893f
C154 plus.t9 a_n1952_n4888# 1.69893f
C155 plus.n16 a_n1952_n4888# 0.633525f
C156 plus.t0 a_n1952_n4888# 1.7177f
C157 plus.n17 a_n1952_n4888# 0.618658f
C158 plus.t1 a_n1952_n4888# 1.69893f
C159 plus.n18 a_n1952_n4888# 0.637843f
C160 plus.n19 a_n1952_n4888# 0.009724f
C161 plus.n20 a_n1952_n4888# 0.178984f
C162 plus.n21 a_n1952_n4888# 0.042852f
C163 plus.n22 a_n1952_n4888# 0.042852f
C164 plus.n23 a_n1952_n4888# 0.009724f
C165 plus.n24 a_n1952_n4888# 0.633525f
C166 plus.n25 a_n1952_n4888# 0.009724f
C167 plus.n26 a_n1952_n4888# 0.631147f
C168 plus.n27 a_n1952_n4888# 1.54682f
.ends

