* NGSPICE file created from diffpair244.ext - technology: sky130A

.subckt diffpair244 minus drain_right drain_left source plus
X0 source.t17 plus.t0 drain_left.t5 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X1 drain_right.t9 minus.t0 source.t5 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X2 drain_left.t0 plus.t1 source.t16 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X3 a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X4 drain_left.t4 plus.t2 source.t15 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X5 source.t7 minus.t1 drain_right.t8 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 source.t14 plus.t3 drain_left.t1 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X8 a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X9 drain_right.t7 minus.t2 source.t6 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X10 a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X11 source.t0 minus.t3 drain_right.t6 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X12 drain_right.t5 minus.t4 source.t4 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X13 drain_right.t4 minus.t5 source.t1 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X14 source.t3 minus.t6 drain_right.t3 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 source.t2 minus.t7 drain_right.t2 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X16 drain_left.t6 plus.t4 source.t13 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X17 drain_right.t1 minus.t8 source.t18 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_right.t0 minus.t9 source.t19 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X19 source.t12 plus.t5 drain_left.t7 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X20 drain_left.t2 plus.t6 source.t11 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X21 drain_left.t9 plus.t7 source.t10 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 source.t9 plus.t8 drain_left.t8 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X23 drain_left.t3 plus.t9 source.t8 a_n1496_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
R0 plus.n3 plus.t4 1216.68
R1 plus.n9 plus.t9 1216.68
R2 plus.n14 plus.t1 1216.68
R3 plus.n20 plus.t2 1216.68
R4 plus.n6 plus.t6 1172.87
R5 plus.n2 plus.t8 1172.87
R6 plus.n8 plus.t5 1172.87
R7 plus.n17 plus.t7 1172.87
R8 plus.n13 plus.t3 1172.87
R9 plus.n19 plus.t0 1172.87
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 51.1217
R25 plus.n9 plus.n8 51.1217
R26 plus.n20 plus.n19 51.1217
R27 plus.n14 plus.n13 51.1217
R28 plus plus.n21 26.41
R29 plus.n2 plus.n1 21.9096
R30 plus.n8 plus.n7 21.9096
R31 plus.n19 plus.n18 21.9096
R32 plus.n13 plus.n12 21.9096
R33 plus plus.n10 9.88497
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 drain_left.n5 drain_left.t6 72.7512
R41 drain_left.n1 drain_left.t4 72.751
R42 drain_left.n3 drain_left.n2 67.5556
R43 drain_left.n5 drain_left.n4 67.1908
R44 drain_left.n7 drain_left.n6 67.1907
R45 drain_left.n1 drain_left.n0 67.1907
R46 drain_left drain_left.n3 25.2031
R47 drain_left drain_left.n7 6.21356
R48 drain_left.n2 drain_left.t1 5.0005
R49 drain_left.n2 drain_left.t0 5.0005
R50 drain_left.n0 drain_left.t5 5.0005
R51 drain_left.n0 drain_left.t9 5.0005
R52 drain_left.n6 drain_left.t7 5.0005
R53 drain_left.n6 drain_left.t3 5.0005
R54 drain_left.n4 drain_left.t8 5.0005
R55 drain_left.n4 drain_left.t2 5.0005
R56 drain_left.n7 drain_left.n5 0.560845
R57 drain_left.n3 drain_left.n1 0.0852402
R58 source.n5 source.t4 55.512
R59 source.n0 source.t8 55.5119
R60 source.n19 source.t5 55.5119
R61 source.n14 source.t16 55.5119
R62 source.n2 source.n1 50.512
R63 source.n4 source.n3 50.512
R64 source.n7 source.n6 50.512
R65 source.n9 source.n8 50.512
R66 source.n18 source.n17 50.5119
R67 source.n16 source.n15 50.5119
R68 source.n13 source.n12 50.5119
R69 source.n11 source.n10 50.5119
R70 source.n11 source.n9 17.863
R71 source.n20 source.n0 11.7595
R72 source.n20 source.n19 5.5436
R73 source.n17 source.t6 5.0005
R74 source.n17 source.t3 5.0005
R75 source.n15 source.t19 5.0005
R76 source.n15 source.t7 5.0005
R77 source.n12 source.t10 5.0005
R78 source.n12 source.t14 5.0005
R79 source.n10 source.t15 5.0005
R80 source.n10 source.t17 5.0005
R81 source.n1 source.t11 5.0005
R82 source.n1 source.t12 5.0005
R83 source.n3 source.t13 5.0005
R84 source.n3 source.t9 5.0005
R85 source.n6 source.t18 5.0005
R86 source.n6 source.t0 5.0005
R87 source.n8 source.t1 5.0005
R88 source.n8 source.t2 5.0005
R89 source.n5 source.n4 0.7505
R90 source.n16 source.n14 0.7505
R91 source.n9 source.n7 0.560845
R92 source.n7 source.n5 0.560845
R93 source.n4 source.n2 0.560845
R94 source.n2 source.n0 0.560845
R95 source.n13 source.n11 0.560845
R96 source.n14 source.n13 0.560845
R97 source.n18 source.n16 0.560845
R98 source.n19 source.n18 0.560845
R99 source source.n20 0.188
R100 minus.n9 minus.t5 1216.68
R101 minus.n3 minus.t4 1216.68
R102 minus.n20 minus.t0 1216.68
R103 minus.n14 minus.t9 1216.68
R104 minus.n6 minus.t8 1172.87
R105 minus.n8 minus.t7 1172.87
R106 minus.n2 minus.t3 1172.87
R107 minus.n17 minus.t2 1172.87
R108 minus.n19 minus.t6 1172.87
R109 minus.n13 minus.t1 1172.87
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 51.1217
R125 minus.n3 minus.n2 51.1217
R126 minus.n14 minus.n13 51.1217
R127 minus.n20 minus.n19 51.1217
R128 minus.n22 minus.n10 30.2562
R129 minus.n8 minus.n7 21.9096
R130 minus.n2 minus.n1 21.9096
R131 minus.n13 minus.n12 21.9096
R132 minus.n19 minus.n18 21.9096
R133 minus.n22 minus.n21 6.51376
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t0 72.751
R142 drain_right.n7 drain_right.t4 72.1908
R143 drain_right.n6 drain_right.n4 67.751
R144 drain_right.n3 drain_right.n2 67.5556
R145 drain_right.n6 drain_right.n5 67.1908
R146 drain_right.n1 drain_right.n0 67.1907
R147 drain_right drain_right.n3 24.6499
R148 drain_right drain_right.n7 5.93339
R149 drain_right.n2 drain_right.t3 5.0005
R150 drain_right.n2 drain_right.t9 5.0005
R151 drain_right.n0 drain_right.t8 5.0005
R152 drain_right.n0 drain_right.t7 5.0005
R153 drain_right.n4 drain_right.t6 5.0005
R154 drain_right.n4 drain_right.t5 5.0005
R155 drain_right.n5 drain_right.t2 5.0005
R156 drain_right.n5 drain_right.t1 5.0005
R157 drain_right.n7 drain_right.n6 0.560845
R158 drain_right.n3 drain_right.n1 0.0852402
C0 source plus 1.27553f
C1 plus minus 3.89236f
C2 drain_right plus 0.297565f
C3 source drain_left 11.8318f
C4 minus drain_left 0.170828f
C5 drain_right drain_left 0.734053f
C6 source minus 1.26119f
C7 drain_right source 11.8258f
C8 plus drain_left 1.59619f
C9 drain_right minus 1.45464f
C10 drain_right a_n1496_n2088# 4.64163f
C11 drain_left a_n1496_n2088# 4.85822f
C12 source a_n1496_n2088# 3.948996f
C13 minus a_n1496_n2088# 5.020319f
C14 plus a_n1496_n2088# 5.93027f
C15 drain_right.t0 a_n1496_n2088# 1.21873f
C16 drain_right.t8 a_n1496_n2088# 0.162163f
C17 drain_right.t7 a_n1496_n2088# 0.162163f
C18 drain_right.n0 a_n1496_n2088# 1.00288f
C19 drain_right.n1 a_n1496_n2088# 0.545415f
C20 drain_right.t3 a_n1496_n2088# 0.162163f
C21 drain_right.t9 a_n1496_n2088# 0.162163f
C22 drain_right.n2 a_n1496_n2088# 1.00429f
C23 drain_right.n3 a_n1496_n2088# 0.94254f
C24 drain_right.t6 a_n1496_n2088# 0.162163f
C25 drain_right.t5 a_n1496_n2088# 0.162163f
C26 drain_right.n4 a_n1496_n2088# 1.00515f
C27 drain_right.t2 a_n1496_n2088# 0.162163f
C28 drain_right.t1 a_n1496_n2088# 0.162163f
C29 drain_right.n5 a_n1496_n2088# 1.00289f
C30 drain_right.n6 a_n1496_n2088# 0.536274f
C31 drain_right.t4 a_n1496_n2088# 1.21633f
C32 drain_right.n7 a_n1496_n2088# 0.500784f
C33 minus.n0 a_n1496_n2088# 0.033226f
C34 minus.t5 a_n1496_n2088# 0.086757f
C35 minus.t7 a_n1496_n2088# 0.085201f
C36 minus.t8 a_n1496_n2088# 0.085201f
C37 minus.n1 a_n1496_n2088# 0.014095f
C38 minus.t3 a_n1496_n2088# 0.085201f
C39 minus.n2 a_n1496_n2088# 0.04423f
C40 minus.t4 a_n1496_n2088# 0.086757f
C41 minus.n3 a_n1496_n2088# 0.05579f
C42 minus.n4 a_n1496_n2088# 0.071529f
C43 minus.n5 a_n1496_n2088# 0.033226f
C44 minus.n6 a_n1496_n2088# 0.055252f
C45 minus.n7 a_n1496_n2088# 0.014095f
C46 minus.n8 a_n1496_n2088# 0.04423f
C47 minus.n9 a_n1496_n2088# 0.055745f
C48 minus.n10 a_n1496_n2088# 0.877391f
C49 minus.n11 a_n1496_n2088# 0.033226f
C50 minus.t6 a_n1496_n2088# 0.085201f
C51 minus.t2 a_n1496_n2088# 0.085201f
C52 minus.n12 a_n1496_n2088# 0.014095f
C53 minus.t9 a_n1496_n2088# 0.086757f
C54 minus.t1 a_n1496_n2088# 0.085201f
C55 minus.n13 a_n1496_n2088# 0.04423f
C56 minus.n14 a_n1496_n2088# 0.05579f
C57 minus.n15 a_n1496_n2088# 0.071529f
C58 minus.n16 a_n1496_n2088# 0.033226f
C59 minus.n17 a_n1496_n2088# 0.055252f
C60 minus.n18 a_n1496_n2088# 0.014095f
C61 minus.n19 a_n1496_n2088# 0.04423f
C62 minus.t0 a_n1496_n2088# 0.086757f
C63 minus.n20 a_n1496_n2088# 0.055745f
C64 minus.n21 a_n1496_n2088# 0.218301f
C65 minus.n22 a_n1496_n2088# 1.08142f
C66 source.t8 a_n1496_n2088# 1.23575f
C67 source.n0 a_n1496_n2088# 0.909111f
C68 source.t11 a_n1496_n2088# 0.175937f
C69 source.t12 a_n1496_n2088# 0.175937f
C70 source.n1 a_n1496_n2088# 1.02398f
C71 source.n2 a_n1496_n2088# 0.318012f
C72 source.t13 a_n1496_n2088# 0.175937f
C73 source.t9 a_n1496_n2088# 0.175937f
C74 source.n3 a_n1496_n2088# 1.02398f
C75 source.n4 a_n1496_n2088# 0.332978f
C76 source.t4 a_n1496_n2088# 1.23575f
C77 source.n5 a_n1496_n2088# 0.437887f
C78 source.t18 a_n1496_n2088# 0.175937f
C79 source.t0 a_n1496_n2088# 0.175937f
C80 source.n6 a_n1496_n2088# 1.02398f
C81 source.n7 a_n1496_n2088# 0.318012f
C82 source.t1 a_n1496_n2088# 0.175937f
C83 source.t2 a_n1496_n2088# 0.175937f
C84 source.n8 a_n1496_n2088# 1.02398f
C85 source.n9 a_n1496_n2088# 1.16409f
C86 source.t15 a_n1496_n2088# 0.175937f
C87 source.t17 a_n1496_n2088# 0.175937f
C88 source.n10 a_n1496_n2088# 1.02397f
C89 source.n11 a_n1496_n2088# 1.1641f
C90 source.t10 a_n1496_n2088# 0.175937f
C91 source.t14 a_n1496_n2088# 0.175937f
C92 source.n12 a_n1496_n2088# 1.02397f
C93 source.n13 a_n1496_n2088# 0.318018f
C94 source.t16 a_n1496_n2088# 1.23575f
C95 source.n14 a_n1496_n2088# 0.437893f
C96 source.t19 a_n1496_n2088# 0.175937f
C97 source.t7 a_n1496_n2088# 0.175937f
C98 source.n15 a_n1496_n2088# 1.02397f
C99 source.n16 a_n1496_n2088# 0.332984f
C100 source.t6 a_n1496_n2088# 0.175937f
C101 source.t3 a_n1496_n2088# 0.175937f
C102 source.n17 a_n1496_n2088# 1.02397f
C103 source.n18 a_n1496_n2088# 0.318018f
C104 source.t5 a_n1496_n2088# 1.23575f
C105 source.n19 a_n1496_n2088# 0.555118f
C106 source.n20 a_n1496_n2088# 1.00277f
C107 drain_left.t4 a_n1496_n2088# 1.20968f
C108 drain_left.t5 a_n1496_n2088# 0.160959f
C109 drain_left.t9 a_n1496_n2088# 0.160959f
C110 drain_left.n0 a_n1496_n2088# 0.995434f
C111 drain_left.n1 a_n1496_n2088# 0.541364f
C112 drain_left.t1 a_n1496_n2088# 0.160959f
C113 drain_left.t0 a_n1496_n2088# 0.160959f
C114 drain_left.n2 a_n1496_n2088# 0.996833f
C115 drain_left.n3 a_n1496_n2088# 0.98129f
C116 drain_left.t6 a_n1496_n2088# 1.20968f
C117 drain_left.t8 a_n1496_n2088# 0.160959f
C118 drain_left.t2 a_n1496_n2088# 0.160959f
C119 drain_left.n4 a_n1496_n2088# 0.995438f
C120 drain_left.n5 a_n1496_n2088# 0.569562f
C121 drain_left.t7 a_n1496_n2088# 0.160959f
C122 drain_left.t3 a_n1496_n2088# 0.160959f
C123 drain_left.n6 a_n1496_n2088# 0.995434f
C124 drain_left.n7 a_n1496_n2088# 0.449868f
C125 plus.n0 a_n1496_n2088# 0.033809f
C126 plus.t5 a_n1496_n2088# 0.086694f
C127 plus.t6 a_n1496_n2088# 0.086694f
C128 plus.n1 a_n1496_n2088# 0.014342f
C129 plus.t4 a_n1496_n2088# 0.088278f
C130 plus.t8 a_n1496_n2088# 0.086694f
C131 plus.n2 a_n1496_n2088# 0.045005f
C132 plus.n3 a_n1496_n2088# 0.056768f
C133 plus.n4 a_n1496_n2088# 0.072783f
C134 plus.n5 a_n1496_n2088# 0.033809f
C135 plus.n6 a_n1496_n2088# 0.056221f
C136 plus.n7 a_n1496_n2088# 0.014342f
C137 plus.n8 a_n1496_n2088# 0.045005f
C138 plus.t9 a_n1496_n2088# 0.088278f
C139 plus.n9 a_n1496_n2088# 0.056722f
C140 plus.n10 a_n1496_n2088# 0.290848f
C141 plus.n11 a_n1496_n2088# 0.033809f
C142 plus.t2 a_n1496_n2088# 0.088278f
C143 plus.t0 a_n1496_n2088# 0.086694f
C144 plus.t7 a_n1496_n2088# 0.086694f
C145 plus.n12 a_n1496_n2088# 0.014342f
C146 plus.t3 a_n1496_n2088# 0.086694f
C147 plus.n13 a_n1496_n2088# 0.045005f
C148 plus.t1 a_n1496_n2088# 0.088278f
C149 plus.n14 a_n1496_n2088# 0.056768f
C150 plus.n15 a_n1496_n2088# 0.072783f
C151 plus.n16 a_n1496_n2088# 0.033809f
C152 plus.n17 a_n1496_n2088# 0.056221f
C153 plus.n18 a_n1496_n2088# 0.014342f
C154 plus.n19 a_n1496_n2088# 0.045005f
C155 plus.n20 a_n1496_n2088# 0.056722f
C156 plus.n21 a_n1496_n2088# 0.807f
.ends

