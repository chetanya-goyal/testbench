* NGSPICE file created from diffpair575.ext - technology: sky130A

.subckt diffpair575 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t21 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t10 plus.t1 source.t13 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 drain_right.t11 minus.t0 source.t6 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X3 source.t20 plus.t2 drain_left.t9 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 drain_left.t8 plus.t3 source.t19 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 source.t4 minus.t1 drain_right.t10 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 source.t10 minus.t2 drain_right.t9 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X7 source.t11 minus.t3 drain_right.t8 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X8 source.t2 minus.t4 drain_right.t7 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X9 drain_right.t6 minus.t5 source.t7 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X10 drain_right.t5 minus.t6 source.t3 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 drain_left.t7 plus.t4 source.t18 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X12 source.t17 plus.t5 drain_left.t6 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X13 a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X14 drain_right.t4 minus.t7 source.t5 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X15 drain_right.t3 minus.t8 source.t8 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X16 drain_right.t2 minus.t9 source.t0 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X17 source.t9 minus.t10 drain_right.t1 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X18 a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X19 a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X20 source.t22 plus.t6 drain_left.t5 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 drain_left.t4 plus.t7 source.t16 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X22 source.t1 minus.t11 drain_right.t0 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X23 source.t12 plus.t8 drain_left.t3 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X24 source.t15 plus.t9 drain_left.t2 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X25 a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X26 source.t14 plus.t10 drain_left.t1 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X27 drain_left.t0 plus.t11 source.t23 a_n1458_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n2 plus.t5 2614.12
R1 plus.n11 plus.t4 2614.12
R2 plus.n15 plus.t0 2614.12
R3 plus.n24 plus.t9 2614.12
R4 plus.n3 plus.t3 2566.65
R5 plus.n1 plus.t10 2566.65
R6 plus.n8 plus.t7 2566.65
R7 plus.n10 plus.t6 2566.65
R8 plus.n16 plus.t2 2566.65
R9 plus.n14 plus.t1 2566.65
R10 plus.n21 plus.t8 2566.65
R11 plus.n23 plus.t11 2566.65
R12 plus.n5 plus.n2 161.489
R13 plus.n18 plus.n15 161.489
R14 plus.n5 plus.n4 161.3
R15 plus.n7 plus.n6 161.3
R16 plus.n9 plus.n0 161.3
R17 plus.n12 plus.n11 161.3
R18 plus.n18 plus.n17 161.3
R19 plus.n20 plus.n19 161.3
R20 plus.n22 plus.n13 161.3
R21 plus.n25 plus.n24 161.3
R22 plus.n4 plus.n3 43.0884
R23 plus.n10 plus.n9 43.0884
R24 plus.n23 plus.n22 43.0884
R25 plus.n17 plus.n16 43.0884
R26 plus.n7 plus.n1 38.7066
R27 plus.n8 plus.n7 38.7066
R28 plus.n21 plus.n20 38.7066
R29 plus.n20 plus.n14 38.7066
R30 plus.n4 plus.n1 34.3247
R31 plus.n9 plus.n8 34.3247
R32 plus.n22 plus.n21 34.3247
R33 plus.n17 plus.n14 34.3247
R34 plus plus.n25 31.5104
R35 plus.n3 plus.n2 29.9429
R36 plus.n11 plus.n10 29.9429
R37 plus.n24 plus.n23 29.9429
R38 plus.n16 plus.n15 29.9429
R39 plus plus.n12 15.1293
R40 plus.n6 plus.n5 0.189894
R41 plus.n6 plus.n0 0.189894
R42 plus.n12 plus.n0 0.189894
R43 plus.n25 plus.n13 0.189894
R44 plus.n19 plus.n13 0.189894
R45 plus.n19 plus.n18 0.189894
R46 source.n0 source.t18 44.1297
R47 source.n5 source.t17 44.1296
R48 source.n6 source.t8 44.1296
R49 source.n11 source.t10 44.1296
R50 source.n23 source.t5 44.1295
R51 source.n18 source.t11 44.1295
R52 source.n17 source.t21 44.1295
R53 source.n12 source.t15 44.1295
R54 source.n2 source.n1 43.1397
R55 source.n4 source.n3 43.1397
R56 source.n8 source.n7 43.1397
R57 source.n10 source.n9 43.1397
R58 source.n22 source.n21 43.1396
R59 source.n20 source.n19 43.1396
R60 source.n16 source.n15 43.1396
R61 source.n14 source.n13 43.1396
R62 source.n12 source.n11 27.8052
R63 source.n24 source.n0 22.3138
R64 source.n24 source.n23 5.49188
R65 source.n21 source.t7 0.9905
R66 source.n21 source.t9 0.9905
R67 source.n19 source.t3 0.9905
R68 source.n19 source.t4 0.9905
R69 source.n15 source.t13 0.9905
R70 source.n15 source.t20 0.9905
R71 source.n13 source.t23 0.9905
R72 source.n13 source.t12 0.9905
R73 source.n1 source.t16 0.9905
R74 source.n1 source.t22 0.9905
R75 source.n3 source.t19 0.9905
R76 source.n3 source.t14 0.9905
R77 source.n7 source.t6 0.9905
R78 source.n7 source.t2 0.9905
R79 source.n9 source.t0 0.9905
R80 source.n9 source.t1 0.9905
R81 source.n6 source.n5 0.470328
R82 source.n18 source.n17 0.470328
R83 source.n11 source.n10 0.457397
R84 source.n10 source.n8 0.457397
R85 source.n8 source.n6 0.457397
R86 source.n5 source.n4 0.457397
R87 source.n4 source.n2 0.457397
R88 source.n2 source.n0 0.457397
R89 source.n14 source.n12 0.457397
R90 source.n16 source.n14 0.457397
R91 source.n17 source.n16 0.457397
R92 source.n20 source.n18 0.457397
R93 source.n22 source.n20 0.457397
R94 source.n23 source.n22 0.457397
R95 source source.n24 0.188
R96 drain_left.n6 drain_left.n4 60.2753
R97 drain_left.n3 drain_left.n2 60.22
R98 drain_left.n3 drain_left.n0 60.22
R99 drain_left.n8 drain_left.n7 59.8185
R100 drain_left.n6 drain_left.n5 59.8185
R101 drain_left.n3 drain_left.n1 59.8184
R102 drain_left drain_left.n3 35.7122
R103 drain_left drain_left.n8 6.11011
R104 drain_left.n1 drain_left.t3 0.9905
R105 drain_left.n1 drain_left.t10 0.9905
R106 drain_left.n2 drain_left.t9 0.9905
R107 drain_left.n2 drain_left.t11 0.9905
R108 drain_left.n0 drain_left.t2 0.9905
R109 drain_left.n0 drain_left.t0 0.9905
R110 drain_left.n7 drain_left.t5 0.9905
R111 drain_left.n7 drain_left.t7 0.9905
R112 drain_left.n5 drain_left.t1 0.9905
R113 drain_left.n5 drain_left.t4 0.9905
R114 drain_left.n4 drain_left.t6 0.9905
R115 drain_left.n4 drain_left.t8 0.9905
R116 drain_left.n8 drain_left.n6 0.457397
R117 minus.n11 minus.t2 2614.12
R118 minus.n2 minus.t8 2614.12
R119 minus.n24 minus.t7 2614.12
R120 minus.n15 minus.t3 2614.12
R121 minus.n10 minus.t9 2566.65
R122 minus.n8 minus.t11 2566.65
R123 minus.n1 minus.t0 2566.65
R124 minus.n3 minus.t4 2566.65
R125 minus.n23 minus.t10 2566.65
R126 minus.n21 minus.t5 2566.65
R127 minus.n14 minus.t1 2566.65
R128 minus.n16 minus.t6 2566.65
R129 minus.n5 minus.n2 161.489
R130 minus.n18 minus.n15 161.489
R131 minus.n12 minus.n11 161.3
R132 minus.n9 minus.n0 161.3
R133 minus.n7 minus.n6 161.3
R134 minus.n5 minus.n4 161.3
R135 minus.n25 minus.n24 161.3
R136 minus.n22 minus.n13 161.3
R137 minus.n20 minus.n19 161.3
R138 minus.n18 minus.n17 161.3
R139 minus.n10 minus.n9 43.0884
R140 minus.n4 minus.n3 43.0884
R141 minus.n17 minus.n16 43.0884
R142 minus.n23 minus.n22 43.0884
R143 minus.n26 minus.n12 40.6596
R144 minus.n8 minus.n7 38.7066
R145 minus.n7 minus.n1 38.7066
R146 minus.n20 minus.n14 38.7066
R147 minus.n21 minus.n20 38.7066
R148 minus.n9 minus.n8 34.3247
R149 minus.n4 minus.n1 34.3247
R150 minus.n17 minus.n14 34.3247
R151 minus.n22 minus.n21 34.3247
R152 minus.n11 minus.n10 29.9429
R153 minus.n3 minus.n2 29.9429
R154 minus.n16 minus.n15 29.9429
R155 minus.n24 minus.n23 29.9429
R156 minus.n26 minus.n25 6.45505
R157 minus.n12 minus.n0 0.189894
R158 minus.n6 minus.n0 0.189894
R159 minus.n6 minus.n5 0.189894
R160 minus.n19 minus.n18 0.189894
R161 minus.n19 minus.n13 0.189894
R162 minus.n25 minus.n13 0.189894
R163 minus minus.n26 0.188
R164 drain_right.n6 drain_right.n4 60.2753
R165 drain_right.n3 drain_right.n2 60.22
R166 drain_right.n3 drain_right.n0 60.22
R167 drain_right.n6 drain_right.n5 59.8185
R168 drain_right.n8 drain_right.n7 59.8185
R169 drain_right.n3 drain_right.n1 59.8184
R170 drain_right drain_right.n3 35.1589
R171 drain_right drain_right.n8 6.11011
R172 drain_right.n1 drain_right.t10 0.9905
R173 drain_right.n1 drain_right.t6 0.9905
R174 drain_right.n2 drain_right.t1 0.9905
R175 drain_right.n2 drain_right.t4 0.9905
R176 drain_right.n0 drain_right.t8 0.9905
R177 drain_right.n0 drain_right.t5 0.9905
R178 drain_right.n4 drain_right.t7 0.9905
R179 drain_right.n4 drain_right.t3 0.9905
R180 drain_right.n5 drain_right.t0 0.9905
R181 drain_right.n5 drain_right.t11 0.9905
R182 drain_right.n7 drain_right.t9 0.9905
R183 drain_right.n7 drain_right.t2 0.9905
R184 drain_right.n8 drain_right.n6 0.457397
C0 plus source 4.8075f
C1 source minus 4.79346f
C2 source drain_left 45.457302f
C3 plus minus 6.45426f
C4 plus drain_left 5.73715f
C5 drain_left minus 0.17046f
C6 source drain_right 45.456398f
C7 plus drain_right 0.292203f
C8 drain_right minus 5.59827f
C9 drain_left drain_right 0.711832f
C10 drain_right a_n1458_n4888# 8.27147f
C11 drain_left a_n1458_n4888# 8.51063f
C12 source a_n1458_n4888# 12.745195f
C13 minus a_n1458_n4888# 6.172699f
C14 plus a_n1458_n4888# 8.84122f
C15 drain_right.t8 a_n1458_n4888# 0.612514f
C16 drain_right.t5 a_n1458_n4888# 0.612514f
C17 drain_right.n0 a_n1458_n4888# 5.60275f
C18 drain_right.t10 a_n1458_n4888# 0.612514f
C19 drain_right.t6 a_n1458_n4888# 0.612514f
C20 drain_right.n1 a_n1458_n4888# 5.599741f
C21 drain_right.t1 a_n1458_n4888# 0.612514f
C22 drain_right.t4 a_n1458_n4888# 0.612514f
C23 drain_right.n2 a_n1458_n4888# 5.60275f
C24 drain_right.n3 a_n1458_n4888# 3.70036f
C25 drain_right.t7 a_n1458_n4888# 0.612514f
C26 drain_right.t3 a_n1458_n4888# 0.612514f
C27 drain_right.n4 a_n1458_n4888# 5.60319f
C28 drain_right.t0 a_n1458_n4888# 0.612514f
C29 drain_right.t11 a_n1458_n4888# 0.612514f
C30 drain_right.n5 a_n1458_n4888# 5.59973f
C31 drain_right.n6 a_n1458_n4888# 0.89447f
C32 drain_right.t9 a_n1458_n4888# 0.612514f
C33 drain_right.t2 a_n1458_n4888# 0.612514f
C34 drain_right.n7 a_n1458_n4888# 5.59973f
C35 drain_right.n8 a_n1458_n4888# 0.758338f
C36 minus.n0 a_n1458_n4888# 0.056617f
C37 minus.t2 a_n1458_n4888# 0.642269f
C38 minus.t9 a_n1458_n4888# 0.637844f
C39 minus.t11 a_n1458_n4888# 0.637844f
C40 minus.t0 a_n1458_n4888# 0.637844f
C41 minus.n1 a_n1458_n4888# 0.242762f
C42 minus.t8 a_n1458_n4888# 0.642269f
C43 minus.n2 a_n1458_n4888# 0.25912f
C44 minus.t4 a_n1458_n4888# 0.637844f
C45 minus.n3 a_n1458_n4888# 0.242762f
C46 minus.n4 a_n1458_n4888# 0.019829f
C47 minus.n5 a_n1458_n4888# 0.125371f
C48 minus.n6 a_n1458_n4888# 0.056617f
C49 minus.n7 a_n1458_n4888# 0.019829f
C50 minus.n8 a_n1458_n4888# 0.242762f
C51 minus.n9 a_n1458_n4888# 0.019829f
C52 minus.n10 a_n1458_n4888# 0.242762f
C53 minus.n11 a_n1458_n4888# 0.259039f
C54 minus.n12 a_n1458_n4888# 2.38798f
C55 minus.n13 a_n1458_n4888# 0.056617f
C56 minus.t10 a_n1458_n4888# 0.637844f
C57 minus.t5 a_n1458_n4888# 0.637844f
C58 minus.t1 a_n1458_n4888# 0.637844f
C59 minus.n14 a_n1458_n4888# 0.242762f
C60 minus.t3 a_n1458_n4888# 0.642269f
C61 minus.n15 a_n1458_n4888# 0.25912f
C62 minus.t6 a_n1458_n4888# 0.637844f
C63 minus.n16 a_n1458_n4888# 0.242762f
C64 minus.n17 a_n1458_n4888# 0.019829f
C65 minus.n18 a_n1458_n4888# 0.125371f
C66 minus.n19 a_n1458_n4888# 0.056617f
C67 minus.n20 a_n1458_n4888# 0.019829f
C68 minus.n21 a_n1458_n4888# 0.242762f
C69 minus.n22 a_n1458_n4888# 0.019829f
C70 minus.n23 a_n1458_n4888# 0.242762f
C71 minus.t7 a_n1458_n4888# 0.642269f
C72 minus.n24 a_n1458_n4888# 0.259039f
C73 minus.n25 a_n1458_n4888# 0.364139f
C74 minus.n26 a_n1458_n4888# 2.86428f
C75 drain_left.t2 a_n1458_n4888# 0.611897f
C76 drain_left.t0 a_n1458_n4888# 0.611897f
C77 drain_left.n0 a_n1458_n4888# 5.59711f
C78 drain_left.t3 a_n1458_n4888# 0.611897f
C79 drain_left.t10 a_n1458_n4888# 0.611897f
C80 drain_left.n1 a_n1458_n4888# 5.5941f
C81 drain_left.t9 a_n1458_n4888# 0.611897f
C82 drain_left.t11 a_n1458_n4888# 0.611897f
C83 drain_left.n2 a_n1458_n4888# 5.59711f
C84 drain_left.n3 a_n1458_n4888# 3.77769f
C85 drain_left.t6 a_n1458_n4888# 0.611897f
C86 drain_left.t8 a_n1458_n4888# 0.611897f
C87 drain_left.n4 a_n1458_n4888# 5.59755f
C88 drain_left.t1 a_n1458_n4888# 0.611897f
C89 drain_left.t4 a_n1458_n4888# 0.611897f
C90 drain_left.n5 a_n1458_n4888# 5.59409f
C91 drain_left.n6 a_n1458_n4888# 0.893569f
C92 drain_left.t5 a_n1458_n4888# 0.611897f
C93 drain_left.t7 a_n1458_n4888# 0.611897f
C94 drain_left.n7 a_n1458_n4888# 5.59409f
C95 drain_left.n8 a_n1458_n4888# 0.757574f
C96 source.t18 a_n1458_n4888# 5.37517f
C97 source.n0 a_n1458_n4888# 2.27321f
C98 source.t16 a_n1458_n4888# 0.470335f
C99 source.t22 a_n1458_n4888# 0.470335f
C100 source.n1 a_n1458_n4888# 4.205f
C101 source.n2 a_n1458_n4888# 0.393212f
C102 source.t19 a_n1458_n4888# 0.470335f
C103 source.t14 a_n1458_n4888# 0.470335f
C104 source.n3 a_n1458_n4888# 4.205f
C105 source.n4 a_n1458_n4888# 0.393212f
C106 source.t17 a_n1458_n4888# 5.37518f
C107 source.n5 a_n1458_n4888# 0.507002f
C108 source.t8 a_n1458_n4888# 5.37518f
C109 source.n6 a_n1458_n4888# 0.507002f
C110 source.t6 a_n1458_n4888# 0.470335f
C111 source.t2 a_n1458_n4888# 0.470335f
C112 source.n7 a_n1458_n4888# 4.205f
C113 source.n8 a_n1458_n4888# 0.393212f
C114 source.t0 a_n1458_n4888# 0.470335f
C115 source.t1 a_n1458_n4888# 0.470335f
C116 source.n9 a_n1458_n4888# 4.205f
C117 source.n10 a_n1458_n4888# 0.393212f
C118 source.t10 a_n1458_n4888# 5.37518f
C119 source.n11 a_n1458_n4888# 2.79708f
C120 source.t15 a_n1458_n4888# 5.37515f
C121 source.n12 a_n1458_n4888# 2.79711f
C122 source.t23 a_n1458_n4888# 0.470335f
C123 source.t12 a_n1458_n4888# 0.470335f
C124 source.n13 a_n1458_n4888# 4.205f
C125 source.n14 a_n1458_n4888# 0.393204f
C126 source.t13 a_n1458_n4888# 0.470335f
C127 source.t20 a_n1458_n4888# 0.470335f
C128 source.n15 a_n1458_n4888# 4.205f
C129 source.n16 a_n1458_n4888# 0.393204f
C130 source.t21 a_n1458_n4888# 5.37515f
C131 source.n17 a_n1458_n4888# 0.507031f
C132 source.t11 a_n1458_n4888# 5.37515f
C133 source.n18 a_n1458_n4888# 0.507031f
C134 source.t3 a_n1458_n4888# 0.470335f
C135 source.t4 a_n1458_n4888# 0.470335f
C136 source.n19 a_n1458_n4888# 4.205f
C137 source.n20 a_n1458_n4888# 0.393204f
C138 source.t7 a_n1458_n4888# 0.470335f
C139 source.t9 a_n1458_n4888# 0.470335f
C140 source.n21 a_n1458_n4888# 4.205f
C141 source.n22 a_n1458_n4888# 0.393204f
C142 source.t5 a_n1458_n4888# 5.37515f
C143 source.n23 a_n1458_n4888# 0.668396f
C144 source.n24 a_n1458_n4888# 2.67376f
C145 plus.n0 a_n1458_n4888# 0.057341f
C146 plus.t6 a_n1458_n4888# 0.645995f
C147 plus.t7 a_n1458_n4888# 0.645995f
C148 plus.t10 a_n1458_n4888# 0.645995f
C149 plus.n1 a_n1458_n4888# 0.245864f
C150 plus.t5 a_n1458_n4888# 0.650476f
C151 plus.n2 a_n1458_n4888# 0.262431f
C152 plus.t3 a_n1458_n4888# 0.645995f
C153 plus.n3 a_n1458_n4888# 0.245864f
C154 plus.n4 a_n1458_n4888# 0.020082f
C155 plus.n5 a_n1458_n4888# 0.126973f
C156 plus.n6 a_n1458_n4888# 0.057341f
C157 plus.n7 a_n1458_n4888# 0.020082f
C158 plus.n8 a_n1458_n4888# 0.245864f
C159 plus.n9 a_n1458_n4888# 0.020082f
C160 plus.n10 a_n1458_n4888# 0.245864f
C161 plus.t4 a_n1458_n4888# 0.650476f
C162 plus.n11 a_n1458_n4888# 0.262349f
C163 plus.n12 a_n1458_n4888# 0.864744f
C164 plus.n13 a_n1458_n4888# 0.057341f
C165 plus.t9 a_n1458_n4888# 0.650476f
C166 plus.t11 a_n1458_n4888# 0.645995f
C167 plus.t8 a_n1458_n4888# 0.645995f
C168 plus.t1 a_n1458_n4888# 0.645995f
C169 plus.n14 a_n1458_n4888# 0.245864f
C170 plus.t0 a_n1458_n4888# 0.650476f
C171 plus.n15 a_n1458_n4888# 0.262431f
C172 plus.t2 a_n1458_n4888# 0.645995f
C173 plus.n16 a_n1458_n4888# 0.245864f
C174 plus.n17 a_n1458_n4888# 0.020082f
C175 plus.n18 a_n1458_n4888# 0.126973f
C176 plus.n19 a_n1458_n4888# 0.057341f
C177 plus.n20 a_n1458_n4888# 0.020082f
C178 plus.n21 a_n1458_n4888# 0.245864f
C179 plus.n22 a_n1458_n4888# 0.020082f
C180 plus.n23 a_n1458_n4888# 0.245864f
C181 plus.n24 a_n1458_n4888# 0.262349f
C182 plus.n25 a_n1458_n4888# 1.90119f
.ends

