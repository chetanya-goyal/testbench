* NGSPICE file created from diffpair274.ext - technology: sky130A

.subckt diffpair274 minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t12 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X1 drain_right.t8 minus.t1 source.t13 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 source.t5 plus.t0 drain_left.t9 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X3 a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X4 a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X5 drain_left.t8 plus.t1 source.t6 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X6 source.t0 plus.t2 drain_left.t7 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 source.t18 minus.t2 drain_right.t7 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X8 source.t11 minus.t3 drain_right.t6 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X9 drain_left.t6 plus.t3 source.t1 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X10 source.t2 plus.t4 drain_left.t5 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X11 drain_left.t4 plus.t5 source.t7 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X12 drain_left.t3 plus.t6 source.t8 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X13 source.t19 minus.t4 drain_right.t5 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X15 a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X16 drain_right.t4 minus.t5 source.t14 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X17 drain_right.t3 minus.t6 source.t15 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X18 drain_right.t2 minus.t7 source.t16 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X19 drain_left.t2 plus.t7 source.t9 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X20 drain_right.t1 minus.t8 source.t17 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X21 drain_left.t1 plus.t8 source.t4 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X22 source.t10 minus.t9 drain_right.t0 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X23 source.t3 plus.t9 drain_left.t0 a_n1472_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n9 minus.t8 624.409
R1 minus.n3 minus.t5 624.409
R2 minus.n20 minus.t0 624.409
R3 minus.n14 minus.t7 624.409
R4 minus.n6 minus.t1 586.433
R5 minus.n8 minus.t4 586.433
R6 minus.n2 minus.t9 586.433
R7 minus.n17 minus.t6 586.433
R8 minus.n19 minus.t2 586.433
R9 minus.n13 minus.t3 586.433
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 54.0429
R25 minus.n3 minus.n2 54.0429
R26 minus.n14 minus.n13 54.0429
R27 minus.n20 minus.n19 54.0429
R28 minus.n22 minus.n10 30.1388
R29 minus.n8 minus.n7 18.9884
R30 minus.n2 minus.n1 18.9884
R31 minus.n13 minus.n12 18.9884
R32 minus.n19 minus.n18 18.9884
R33 minus.n22 minus.n21 6.48724
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 source.n138 source.n112 289.615
R42 source.n102 source.n76 289.615
R43 source.n26 source.n0 289.615
R44 source.n62 source.n36 289.615
R45 source.n123 source.n122 185
R46 source.n120 source.n119 185
R47 source.n129 source.n128 185
R48 source.n131 source.n130 185
R49 source.n116 source.n115 185
R50 source.n137 source.n136 185
R51 source.n139 source.n138 185
R52 source.n87 source.n86 185
R53 source.n84 source.n83 185
R54 source.n93 source.n92 185
R55 source.n95 source.n94 185
R56 source.n80 source.n79 185
R57 source.n101 source.n100 185
R58 source.n103 source.n102 185
R59 source.n27 source.n26 185
R60 source.n25 source.n24 185
R61 source.n4 source.n3 185
R62 source.n19 source.n18 185
R63 source.n17 source.n16 185
R64 source.n8 source.n7 185
R65 source.n11 source.n10 185
R66 source.n63 source.n62 185
R67 source.n61 source.n60 185
R68 source.n40 source.n39 185
R69 source.n55 source.n54 185
R70 source.n53 source.n52 185
R71 source.n44 source.n43 185
R72 source.n47 source.n46 185
R73 source.t12 source.n121 147.661
R74 source.t7 source.n85 147.661
R75 source.t1 source.n9 147.661
R76 source.t14 source.n45 147.661
R77 source.n122 source.n119 104.615
R78 source.n129 source.n119 104.615
R79 source.n130 source.n129 104.615
R80 source.n130 source.n115 104.615
R81 source.n137 source.n115 104.615
R82 source.n138 source.n137 104.615
R83 source.n86 source.n83 104.615
R84 source.n93 source.n83 104.615
R85 source.n94 source.n93 104.615
R86 source.n94 source.n79 104.615
R87 source.n101 source.n79 104.615
R88 source.n102 source.n101 104.615
R89 source.n26 source.n25 104.615
R90 source.n25 source.n3 104.615
R91 source.n18 source.n3 104.615
R92 source.n18 source.n17 104.615
R93 source.n17 source.n7 104.615
R94 source.n10 source.n7 104.615
R95 source.n62 source.n61 104.615
R96 source.n61 source.n39 104.615
R97 source.n54 source.n39 104.615
R98 source.n54 source.n53 104.615
R99 source.n53 source.n43 104.615
R100 source.n46 source.n43 104.615
R101 source.n122 source.t12 52.3082
R102 source.n86 source.t7 52.3082
R103 source.n10 source.t1 52.3082
R104 source.n46 source.t14 52.3082
R105 source.n33 source.n32 50.512
R106 source.n35 source.n34 50.512
R107 source.n69 source.n68 50.512
R108 source.n71 source.n70 50.512
R109 source.n111 source.n110 50.5119
R110 source.n109 source.n108 50.5119
R111 source.n75 source.n74 50.5119
R112 source.n73 source.n72 50.5119
R113 source.n143 source.n142 32.1853
R114 source.n107 source.n106 32.1853
R115 source.n31 source.n30 32.1853
R116 source.n67 source.n66 32.1853
R117 source.n73 source.n71 17.8285
R118 source.n123 source.n121 15.6674
R119 source.n87 source.n85 15.6674
R120 source.n11 source.n9 15.6674
R121 source.n47 source.n45 15.6674
R122 source.n124 source.n120 12.8005
R123 source.n88 source.n84 12.8005
R124 source.n12 source.n8 12.8005
R125 source.n48 source.n44 12.8005
R126 source.n128 source.n127 12.0247
R127 source.n92 source.n91 12.0247
R128 source.n16 source.n15 12.0247
R129 source.n52 source.n51 12.0247
R130 source.n144 source.n31 11.7509
R131 source.n131 source.n118 11.249
R132 source.n95 source.n82 11.249
R133 source.n19 source.n6 11.249
R134 source.n55 source.n42 11.249
R135 source.n132 source.n116 10.4732
R136 source.n96 source.n80 10.4732
R137 source.n20 source.n4 10.4732
R138 source.n56 source.n40 10.4732
R139 source.n136 source.n135 9.69747
R140 source.n100 source.n99 9.69747
R141 source.n24 source.n23 9.69747
R142 source.n60 source.n59 9.69747
R143 source.n142 source.n141 9.45567
R144 source.n106 source.n105 9.45567
R145 source.n30 source.n29 9.45567
R146 source.n66 source.n65 9.45567
R147 source.n141 source.n140 9.3005
R148 source.n114 source.n113 9.3005
R149 source.n135 source.n134 9.3005
R150 source.n133 source.n132 9.3005
R151 source.n118 source.n117 9.3005
R152 source.n127 source.n126 9.3005
R153 source.n125 source.n124 9.3005
R154 source.n105 source.n104 9.3005
R155 source.n78 source.n77 9.3005
R156 source.n99 source.n98 9.3005
R157 source.n97 source.n96 9.3005
R158 source.n82 source.n81 9.3005
R159 source.n91 source.n90 9.3005
R160 source.n89 source.n88 9.3005
R161 source.n29 source.n28 9.3005
R162 source.n2 source.n1 9.3005
R163 source.n23 source.n22 9.3005
R164 source.n21 source.n20 9.3005
R165 source.n6 source.n5 9.3005
R166 source.n15 source.n14 9.3005
R167 source.n13 source.n12 9.3005
R168 source.n65 source.n64 9.3005
R169 source.n38 source.n37 9.3005
R170 source.n59 source.n58 9.3005
R171 source.n57 source.n56 9.3005
R172 source.n42 source.n41 9.3005
R173 source.n51 source.n50 9.3005
R174 source.n49 source.n48 9.3005
R175 source.n139 source.n114 8.92171
R176 source.n103 source.n78 8.92171
R177 source.n27 source.n2 8.92171
R178 source.n63 source.n38 8.92171
R179 source.n140 source.n112 8.14595
R180 source.n104 source.n76 8.14595
R181 source.n28 source.n0 8.14595
R182 source.n64 source.n36 8.14595
R183 source.n142 source.n112 5.81868
R184 source.n106 source.n76 5.81868
R185 source.n30 source.n0 5.81868
R186 source.n66 source.n36 5.81868
R187 source.n144 source.n143 5.53498
R188 source.n140 source.n139 5.04292
R189 source.n104 source.n103 5.04292
R190 source.n28 source.n27 5.04292
R191 source.n64 source.n63 5.04292
R192 source.n125 source.n121 4.38594
R193 source.n89 source.n85 4.38594
R194 source.n13 source.n9 4.38594
R195 source.n49 source.n45 4.38594
R196 source.n136 source.n114 4.26717
R197 source.n100 source.n78 4.26717
R198 source.n24 source.n2 4.26717
R199 source.n60 source.n38 4.26717
R200 source.n135 source.n116 3.49141
R201 source.n99 source.n80 3.49141
R202 source.n23 source.n4 3.49141
R203 source.n59 source.n40 3.49141
R204 source.n110 source.t15 3.3005
R205 source.n110 source.t18 3.3005
R206 source.n108 source.t16 3.3005
R207 source.n108 source.t11 3.3005
R208 source.n74 source.t8 3.3005
R209 source.n74 source.t5 3.3005
R210 source.n72 source.t4 3.3005
R211 source.n72 source.t0 3.3005
R212 source.n32 source.t9 3.3005
R213 source.n32 source.t3 3.3005
R214 source.n34 source.t6 3.3005
R215 source.n34 source.t2 3.3005
R216 source.n68 source.t13 3.3005
R217 source.n68 source.t10 3.3005
R218 source.n70 source.t17 3.3005
R219 source.n70 source.t19 3.3005
R220 source.n132 source.n131 2.71565
R221 source.n96 source.n95 2.71565
R222 source.n20 source.n19 2.71565
R223 source.n56 source.n55 2.71565
R224 source.n128 source.n118 1.93989
R225 source.n92 source.n82 1.93989
R226 source.n16 source.n6 1.93989
R227 source.n52 source.n42 1.93989
R228 source.n127 source.n120 1.16414
R229 source.n91 source.n84 1.16414
R230 source.n15 source.n8 1.16414
R231 source.n51 source.n44 1.16414
R232 source.n67 source.n35 0.741879
R233 source.n109 source.n107 0.741879
R234 source.n71 source.n69 0.543603
R235 source.n69 source.n67 0.543603
R236 source.n35 source.n33 0.543603
R237 source.n33 source.n31 0.543603
R238 source.n75 source.n73 0.543603
R239 source.n107 source.n75 0.543603
R240 source.n111 source.n109 0.543603
R241 source.n143 source.n111 0.543603
R242 source.n124 source.n123 0.388379
R243 source.n88 source.n87 0.388379
R244 source.n12 source.n11 0.388379
R245 source.n48 source.n47 0.388379
R246 source source.n144 0.188
R247 source.n126 source.n125 0.155672
R248 source.n126 source.n117 0.155672
R249 source.n133 source.n117 0.155672
R250 source.n134 source.n133 0.155672
R251 source.n134 source.n113 0.155672
R252 source.n141 source.n113 0.155672
R253 source.n90 source.n89 0.155672
R254 source.n90 source.n81 0.155672
R255 source.n97 source.n81 0.155672
R256 source.n98 source.n97 0.155672
R257 source.n98 source.n77 0.155672
R258 source.n105 source.n77 0.155672
R259 source.n29 source.n1 0.155672
R260 source.n22 source.n1 0.155672
R261 source.n22 source.n21 0.155672
R262 source.n21 source.n5 0.155672
R263 source.n14 source.n5 0.155672
R264 source.n14 source.n13 0.155672
R265 source.n65 source.n37 0.155672
R266 source.n58 source.n37 0.155672
R267 source.n58 source.n57 0.155672
R268 source.n57 source.n41 0.155672
R269 source.n50 source.n41 0.155672
R270 source.n50 source.n49 0.155672
R271 drain_right.n26 drain_right.n0 289.615
R272 drain_right.n64 drain_right.n38 289.615
R273 drain_right.n11 drain_right.n10 185
R274 drain_right.n8 drain_right.n7 185
R275 drain_right.n17 drain_right.n16 185
R276 drain_right.n19 drain_right.n18 185
R277 drain_right.n4 drain_right.n3 185
R278 drain_right.n25 drain_right.n24 185
R279 drain_right.n27 drain_right.n26 185
R280 drain_right.n65 drain_right.n64 185
R281 drain_right.n63 drain_right.n62 185
R282 drain_right.n42 drain_right.n41 185
R283 drain_right.n57 drain_right.n56 185
R284 drain_right.n55 drain_right.n54 185
R285 drain_right.n46 drain_right.n45 185
R286 drain_right.n49 drain_right.n48 185
R287 drain_right.t2 drain_right.n9 147.661
R288 drain_right.t1 drain_right.n47 147.661
R289 drain_right.n10 drain_right.n7 104.615
R290 drain_right.n17 drain_right.n7 104.615
R291 drain_right.n18 drain_right.n17 104.615
R292 drain_right.n18 drain_right.n3 104.615
R293 drain_right.n25 drain_right.n3 104.615
R294 drain_right.n26 drain_right.n25 104.615
R295 drain_right.n64 drain_right.n63 104.615
R296 drain_right.n63 drain_right.n41 104.615
R297 drain_right.n56 drain_right.n41 104.615
R298 drain_right.n56 drain_right.n55 104.615
R299 drain_right.n55 drain_right.n45 104.615
R300 drain_right.n48 drain_right.n45 104.615
R301 drain_right.n37 drain_right.n35 67.7338
R302 drain_right.n34 drain_right.n33 67.5426
R303 drain_right.n37 drain_right.n36 67.1908
R304 drain_right.n32 drain_right.n31 67.1907
R305 drain_right.n10 drain_right.t2 52.3082
R306 drain_right.n48 drain_right.t1 52.3082
R307 drain_right.n32 drain_right.n30 49.4072
R308 drain_right.n69 drain_right.n68 48.8641
R309 drain_right drain_right.n34 24.5766
R310 drain_right.n11 drain_right.n9 15.6674
R311 drain_right.n49 drain_right.n47 15.6674
R312 drain_right.n12 drain_right.n8 12.8005
R313 drain_right.n50 drain_right.n46 12.8005
R314 drain_right.n16 drain_right.n15 12.0247
R315 drain_right.n54 drain_right.n53 12.0247
R316 drain_right.n19 drain_right.n6 11.249
R317 drain_right.n57 drain_right.n44 11.249
R318 drain_right.n20 drain_right.n4 10.4732
R319 drain_right.n58 drain_right.n42 10.4732
R320 drain_right.n24 drain_right.n23 9.69747
R321 drain_right.n62 drain_right.n61 9.69747
R322 drain_right.n30 drain_right.n29 9.45567
R323 drain_right.n68 drain_right.n67 9.45567
R324 drain_right.n29 drain_right.n28 9.3005
R325 drain_right.n2 drain_right.n1 9.3005
R326 drain_right.n23 drain_right.n22 9.3005
R327 drain_right.n21 drain_right.n20 9.3005
R328 drain_right.n6 drain_right.n5 9.3005
R329 drain_right.n15 drain_right.n14 9.3005
R330 drain_right.n13 drain_right.n12 9.3005
R331 drain_right.n67 drain_right.n66 9.3005
R332 drain_right.n40 drain_right.n39 9.3005
R333 drain_right.n61 drain_right.n60 9.3005
R334 drain_right.n59 drain_right.n58 9.3005
R335 drain_right.n44 drain_right.n43 9.3005
R336 drain_right.n53 drain_right.n52 9.3005
R337 drain_right.n51 drain_right.n50 9.3005
R338 drain_right.n27 drain_right.n2 8.92171
R339 drain_right.n65 drain_right.n40 8.92171
R340 drain_right.n28 drain_right.n0 8.14595
R341 drain_right.n66 drain_right.n38 8.14595
R342 drain_right drain_right.n69 5.92477
R343 drain_right.n30 drain_right.n0 5.81868
R344 drain_right.n68 drain_right.n38 5.81868
R345 drain_right.n28 drain_right.n27 5.04292
R346 drain_right.n66 drain_right.n65 5.04292
R347 drain_right.n13 drain_right.n9 4.38594
R348 drain_right.n51 drain_right.n47 4.38594
R349 drain_right.n24 drain_right.n2 4.26717
R350 drain_right.n62 drain_right.n40 4.26717
R351 drain_right.n23 drain_right.n4 3.49141
R352 drain_right.n61 drain_right.n42 3.49141
R353 drain_right.n33 drain_right.t7 3.3005
R354 drain_right.n33 drain_right.t9 3.3005
R355 drain_right.n31 drain_right.t6 3.3005
R356 drain_right.n31 drain_right.t3 3.3005
R357 drain_right.n35 drain_right.t0 3.3005
R358 drain_right.n35 drain_right.t4 3.3005
R359 drain_right.n36 drain_right.t5 3.3005
R360 drain_right.n36 drain_right.t8 3.3005
R361 drain_right.n20 drain_right.n19 2.71565
R362 drain_right.n58 drain_right.n57 2.71565
R363 drain_right.n16 drain_right.n6 1.93989
R364 drain_right.n54 drain_right.n44 1.93989
R365 drain_right.n15 drain_right.n8 1.16414
R366 drain_right.n53 drain_right.n46 1.16414
R367 drain_right.n69 drain_right.n37 0.543603
R368 drain_right.n12 drain_right.n11 0.388379
R369 drain_right.n50 drain_right.n49 0.388379
R370 drain_right.n14 drain_right.n13 0.155672
R371 drain_right.n14 drain_right.n5 0.155672
R372 drain_right.n21 drain_right.n5 0.155672
R373 drain_right.n22 drain_right.n21 0.155672
R374 drain_right.n22 drain_right.n1 0.155672
R375 drain_right.n29 drain_right.n1 0.155672
R376 drain_right.n67 drain_right.n39 0.155672
R377 drain_right.n60 drain_right.n39 0.155672
R378 drain_right.n60 drain_right.n59 0.155672
R379 drain_right.n59 drain_right.n43 0.155672
R380 drain_right.n52 drain_right.n43 0.155672
R381 drain_right.n52 drain_right.n51 0.155672
R382 drain_right.n34 drain_right.n32 0.0809298
R383 plus.n3 plus.t1 624.409
R384 plus.n9 plus.t3 624.409
R385 plus.n14 plus.t5 624.409
R386 plus.n20 plus.t8 624.409
R387 plus.n6 plus.t7 586.433
R388 plus.n2 plus.t4 586.433
R389 plus.n8 plus.t9 586.433
R390 plus.n17 plus.t6 586.433
R391 plus.n13 plus.t0 586.433
R392 plus.n19 plus.t2 586.433
R393 plus.n4 plus.n3 161.489
R394 plus.n15 plus.n14 161.489
R395 plus.n4 plus.n1 161.3
R396 plus.n6 plus.n5 161.3
R397 plus.n7 plus.n0 161.3
R398 plus.n10 plus.n9 161.3
R399 plus.n15 plus.n12 161.3
R400 plus.n17 plus.n16 161.3
R401 plus.n18 plus.n11 161.3
R402 plus.n21 plus.n20 161.3
R403 plus.n6 plus.n1 73.0308
R404 plus.n7 plus.n6 73.0308
R405 plus.n18 plus.n17 73.0308
R406 plus.n17 plus.n12 73.0308
R407 plus.n3 plus.n2 54.0429
R408 plus.n9 plus.n8 54.0429
R409 plus.n20 plus.n19 54.0429
R410 plus.n14 plus.n13 54.0429
R411 plus plus.n21 26.2926
R412 plus.n2 plus.n1 18.9884
R413 plus.n8 plus.n7 18.9884
R414 plus.n19 plus.n18 18.9884
R415 plus.n13 plus.n12 18.9884
R416 plus plus.n10 9.85845
R417 plus.n5 plus.n4 0.189894
R418 plus.n5 plus.n0 0.189894
R419 plus.n10 plus.n0 0.189894
R420 plus.n21 plus.n11 0.189894
R421 plus.n16 plus.n11 0.189894
R422 plus.n16 plus.n15 0.189894
R423 drain_left.n26 drain_left.n0 289.615
R424 drain_left.n61 drain_left.n35 289.615
R425 drain_left.n11 drain_left.n10 185
R426 drain_left.n8 drain_left.n7 185
R427 drain_left.n17 drain_left.n16 185
R428 drain_left.n19 drain_left.n18 185
R429 drain_left.n4 drain_left.n3 185
R430 drain_left.n25 drain_left.n24 185
R431 drain_left.n27 drain_left.n26 185
R432 drain_left.n62 drain_left.n61 185
R433 drain_left.n60 drain_left.n59 185
R434 drain_left.n39 drain_left.n38 185
R435 drain_left.n54 drain_left.n53 185
R436 drain_left.n52 drain_left.n51 185
R437 drain_left.n43 drain_left.n42 185
R438 drain_left.n46 drain_left.n45 185
R439 drain_left.t1 drain_left.n9 147.661
R440 drain_left.t8 drain_left.n44 147.661
R441 drain_left.n10 drain_left.n7 104.615
R442 drain_left.n17 drain_left.n7 104.615
R443 drain_left.n18 drain_left.n17 104.615
R444 drain_left.n18 drain_left.n3 104.615
R445 drain_left.n25 drain_left.n3 104.615
R446 drain_left.n26 drain_left.n25 104.615
R447 drain_left.n61 drain_left.n60 104.615
R448 drain_left.n60 drain_left.n38 104.615
R449 drain_left.n53 drain_left.n38 104.615
R450 drain_left.n53 drain_left.n52 104.615
R451 drain_left.n52 drain_left.n42 104.615
R452 drain_left.n45 drain_left.n42 104.615
R453 drain_left.n34 drain_left.n33 67.5426
R454 drain_left.n67 drain_left.n66 67.1908
R455 drain_left.n69 drain_left.n68 67.1907
R456 drain_left.n32 drain_left.n31 67.1907
R457 drain_left.n10 drain_left.t1 52.3082
R458 drain_left.n45 drain_left.t8 52.3082
R459 drain_left.n32 drain_left.n30 49.4072
R460 drain_left.n67 drain_left.n65 49.4072
R461 drain_left drain_left.n34 25.1298
R462 drain_left.n11 drain_left.n9 15.6674
R463 drain_left.n46 drain_left.n44 15.6674
R464 drain_left.n12 drain_left.n8 12.8005
R465 drain_left.n47 drain_left.n43 12.8005
R466 drain_left.n16 drain_left.n15 12.0247
R467 drain_left.n51 drain_left.n50 12.0247
R468 drain_left.n19 drain_left.n6 11.249
R469 drain_left.n54 drain_left.n41 11.249
R470 drain_left.n20 drain_left.n4 10.4732
R471 drain_left.n55 drain_left.n39 10.4732
R472 drain_left.n24 drain_left.n23 9.69747
R473 drain_left.n59 drain_left.n58 9.69747
R474 drain_left.n30 drain_left.n29 9.45567
R475 drain_left.n65 drain_left.n64 9.45567
R476 drain_left.n29 drain_left.n28 9.3005
R477 drain_left.n2 drain_left.n1 9.3005
R478 drain_left.n23 drain_left.n22 9.3005
R479 drain_left.n21 drain_left.n20 9.3005
R480 drain_left.n6 drain_left.n5 9.3005
R481 drain_left.n15 drain_left.n14 9.3005
R482 drain_left.n13 drain_left.n12 9.3005
R483 drain_left.n64 drain_left.n63 9.3005
R484 drain_left.n37 drain_left.n36 9.3005
R485 drain_left.n58 drain_left.n57 9.3005
R486 drain_left.n56 drain_left.n55 9.3005
R487 drain_left.n41 drain_left.n40 9.3005
R488 drain_left.n50 drain_left.n49 9.3005
R489 drain_left.n48 drain_left.n47 9.3005
R490 drain_left.n27 drain_left.n2 8.92171
R491 drain_left.n62 drain_left.n37 8.92171
R492 drain_left.n28 drain_left.n0 8.14595
R493 drain_left.n63 drain_left.n35 8.14595
R494 drain_left drain_left.n69 6.19632
R495 drain_left.n30 drain_left.n0 5.81868
R496 drain_left.n65 drain_left.n35 5.81868
R497 drain_left.n28 drain_left.n27 5.04292
R498 drain_left.n63 drain_left.n62 5.04292
R499 drain_left.n13 drain_left.n9 4.38594
R500 drain_left.n48 drain_left.n44 4.38594
R501 drain_left.n24 drain_left.n2 4.26717
R502 drain_left.n59 drain_left.n37 4.26717
R503 drain_left.n23 drain_left.n4 3.49141
R504 drain_left.n58 drain_left.n39 3.49141
R505 drain_left.n33 drain_left.t9 3.3005
R506 drain_left.n33 drain_left.t4 3.3005
R507 drain_left.n31 drain_left.t7 3.3005
R508 drain_left.n31 drain_left.t3 3.3005
R509 drain_left.n68 drain_left.t0 3.3005
R510 drain_left.n68 drain_left.t6 3.3005
R511 drain_left.n66 drain_left.t5 3.3005
R512 drain_left.n66 drain_left.t2 3.3005
R513 drain_left.n20 drain_left.n19 2.71565
R514 drain_left.n55 drain_left.n54 2.71565
R515 drain_left.n16 drain_left.n6 1.93989
R516 drain_left.n51 drain_left.n41 1.93989
R517 drain_left.n15 drain_left.n8 1.16414
R518 drain_left.n50 drain_left.n43 1.16414
R519 drain_left.n69 drain_left.n67 0.543603
R520 drain_left.n12 drain_left.n11 0.388379
R521 drain_left.n47 drain_left.n46 0.388379
R522 drain_left.n14 drain_left.n13 0.155672
R523 drain_left.n14 drain_left.n5 0.155672
R524 drain_left.n21 drain_left.n5 0.155672
R525 drain_left.n22 drain_left.n21 0.155672
R526 drain_left.n22 drain_left.n1 0.155672
R527 drain_left.n29 drain_left.n1 0.155672
R528 drain_left.n64 drain_left.n36 0.155672
R529 drain_left.n57 drain_left.n36 0.155672
R530 drain_left.n57 drain_left.n56 0.155672
R531 drain_left.n56 drain_left.n40 0.155672
R532 drain_left.n49 drain_left.n40 0.155672
R533 drain_left.n49 drain_left.n48 0.155672
R534 drain_left.n34 drain_left.n32 0.0809298
C0 drain_left drain_right 0.722329f
C1 plus drain_right 0.295575f
C2 source drain_right 11.5935f
C3 minus drain_right 2.19651f
C4 plus drain_left 2.3355f
C5 source drain_left 11.5997f
C6 source plus 2.11543f
C7 minus drain_left 0.171269f
C8 minus plus 3.87675f
C9 source minus 2.10109f
C10 drain_right a_n1472_n2088# 5.04608f
C11 drain_left a_n1472_n2088# 5.28457f
C12 source a_n1472_n2088# 3.898896f
C13 minus a_n1472_n2088# 5.228645f
C14 plus a_n1472_n2088# 6.78415f
C15 drain_left.n0 a_n1472_n2088# 0.040983f
C16 drain_left.n1 a_n1472_n2088# 0.029157f
C17 drain_left.n2 a_n1472_n2088# 0.015668f
C18 drain_left.n3 a_n1472_n2088# 0.037033f
C19 drain_left.n4 a_n1472_n2088# 0.01659f
C20 drain_left.n5 a_n1472_n2088# 0.029157f
C21 drain_left.n6 a_n1472_n2088# 0.015668f
C22 drain_left.n7 a_n1472_n2088# 0.037033f
C23 drain_left.n8 a_n1472_n2088# 0.01659f
C24 drain_left.n9 a_n1472_n2088# 0.124773f
C25 drain_left.t1 a_n1472_n2088# 0.060359f
C26 drain_left.n10 a_n1472_n2088# 0.027775f
C27 drain_left.n11 a_n1472_n2088# 0.021875f
C28 drain_left.n12 a_n1472_n2088# 0.015668f
C29 drain_left.n13 a_n1472_n2088# 0.693771f
C30 drain_left.n14 a_n1472_n2088# 0.029157f
C31 drain_left.n15 a_n1472_n2088# 0.015668f
C32 drain_left.n16 a_n1472_n2088# 0.01659f
C33 drain_left.n17 a_n1472_n2088# 0.037033f
C34 drain_left.n18 a_n1472_n2088# 0.037033f
C35 drain_left.n19 a_n1472_n2088# 0.01659f
C36 drain_left.n20 a_n1472_n2088# 0.015668f
C37 drain_left.n21 a_n1472_n2088# 0.029157f
C38 drain_left.n22 a_n1472_n2088# 0.029157f
C39 drain_left.n23 a_n1472_n2088# 0.015668f
C40 drain_left.n24 a_n1472_n2088# 0.01659f
C41 drain_left.n25 a_n1472_n2088# 0.037033f
C42 drain_left.n26 a_n1472_n2088# 0.080171f
C43 drain_left.n27 a_n1472_n2088# 0.01659f
C44 drain_left.n28 a_n1472_n2088# 0.015668f
C45 drain_left.n29 a_n1472_n2088# 0.067396f
C46 drain_left.n30 a_n1472_n2088# 0.066169f
C47 drain_left.t7 a_n1472_n2088# 0.138246f
C48 drain_left.t3 a_n1472_n2088# 0.138246f
C49 drain_left.n31 a_n1472_n2088# 1.15297f
C50 drain_left.n32 a_n1472_n2088# 0.409629f
C51 drain_left.t9 a_n1472_n2088# 0.138246f
C52 drain_left.t4 a_n1472_n2088# 0.138246f
C53 drain_left.n33 a_n1472_n2088# 1.15472f
C54 drain_left.n34 a_n1472_n2088# 1.26548f
C55 drain_left.n35 a_n1472_n2088# 0.040983f
C56 drain_left.n36 a_n1472_n2088# 0.029157f
C57 drain_left.n37 a_n1472_n2088# 0.015668f
C58 drain_left.n38 a_n1472_n2088# 0.037033f
C59 drain_left.n39 a_n1472_n2088# 0.01659f
C60 drain_left.n40 a_n1472_n2088# 0.029157f
C61 drain_left.n41 a_n1472_n2088# 0.015668f
C62 drain_left.n42 a_n1472_n2088# 0.037033f
C63 drain_left.n43 a_n1472_n2088# 0.01659f
C64 drain_left.n44 a_n1472_n2088# 0.124773f
C65 drain_left.t8 a_n1472_n2088# 0.060359f
C66 drain_left.n45 a_n1472_n2088# 0.027775f
C67 drain_left.n46 a_n1472_n2088# 0.021875f
C68 drain_left.n47 a_n1472_n2088# 0.015668f
C69 drain_left.n48 a_n1472_n2088# 0.693771f
C70 drain_left.n49 a_n1472_n2088# 0.029157f
C71 drain_left.n50 a_n1472_n2088# 0.015668f
C72 drain_left.n51 a_n1472_n2088# 0.01659f
C73 drain_left.n52 a_n1472_n2088# 0.037033f
C74 drain_left.n53 a_n1472_n2088# 0.037033f
C75 drain_left.n54 a_n1472_n2088# 0.01659f
C76 drain_left.n55 a_n1472_n2088# 0.015668f
C77 drain_left.n56 a_n1472_n2088# 0.029157f
C78 drain_left.n57 a_n1472_n2088# 0.029157f
C79 drain_left.n58 a_n1472_n2088# 0.015668f
C80 drain_left.n59 a_n1472_n2088# 0.01659f
C81 drain_left.n60 a_n1472_n2088# 0.037033f
C82 drain_left.n61 a_n1472_n2088# 0.080171f
C83 drain_left.n62 a_n1472_n2088# 0.01659f
C84 drain_left.n63 a_n1472_n2088# 0.015668f
C85 drain_left.n64 a_n1472_n2088# 0.067396f
C86 drain_left.n65 a_n1472_n2088# 0.066169f
C87 drain_left.t5 a_n1472_n2088# 0.138246f
C88 drain_left.t2 a_n1472_n2088# 0.138246f
C89 drain_left.n66 a_n1472_n2088# 1.15298f
C90 drain_left.n67 a_n1472_n2088# 0.444688f
C91 drain_left.t0 a_n1472_n2088# 0.138246f
C92 drain_left.t6 a_n1472_n2088# 0.138246f
C93 drain_left.n68 a_n1472_n2088# 1.15297f
C94 drain_left.n69 a_n1472_n2088# 0.581396f
C95 plus.n0 a_n1472_n2088# 0.054961f
C96 plus.t9 a_n1472_n2088# 0.281867f
C97 plus.t7 a_n1472_n2088# 0.281867f
C98 plus.n1 a_n1472_n2088# 0.022637f
C99 plus.t1 a_n1472_n2088# 0.28986f
C100 plus.t4 a_n1472_n2088# 0.281867f
C101 plus.n2 a_n1472_n2088# 0.129382f
C102 plus.n3 a_n1472_n2088# 0.146137f
C103 plus.n4 a_n1472_n2088# 0.120688f
C104 plus.n5 a_n1472_n2088# 0.054961f
C105 plus.n6 a_n1472_n2088# 0.147614f
C106 plus.n7 a_n1472_n2088# 0.022637f
C107 plus.n8 a_n1472_n2088# 0.129382f
C108 plus.t3 a_n1472_n2088# 0.28986f
C109 plus.n9 a_n1472_n2088# 0.14606f
C110 plus.n10 a_n1472_n2088# 0.469232f
C111 plus.n11 a_n1472_n2088# 0.054961f
C112 plus.t8 a_n1472_n2088# 0.28986f
C113 plus.t2 a_n1472_n2088# 0.281867f
C114 plus.t6 a_n1472_n2088# 0.281867f
C115 plus.n12 a_n1472_n2088# 0.022637f
C116 plus.t0 a_n1472_n2088# 0.281867f
C117 plus.n13 a_n1472_n2088# 0.129382f
C118 plus.t5 a_n1472_n2088# 0.28986f
C119 plus.n14 a_n1472_n2088# 0.146137f
C120 plus.n15 a_n1472_n2088# 0.120688f
C121 plus.n16 a_n1472_n2088# 0.054961f
C122 plus.n17 a_n1472_n2088# 0.147614f
C123 plus.n18 a_n1472_n2088# 0.022637f
C124 plus.n19 a_n1472_n2088# 0.129382f
C125 plus.n20 a_n1472_n2088# 0.14606f
C126 plus.n21 a_n1472_n2088# 1.30183f
C127 drain_right.n0 a_n1472_n2088# 0.041025f
C128 drain_right.n1 a_n1472_n2088# 0.029187f
C129 drain_right.n2 a_n1472_n2088# 0.015684f
C130 drain_right.n3 a_n1472_n2088# 0.037071f
C131 drain_right.n4 a_n1472_n2088# 0.016606f
C132 drain_right.n5 a_n1472_n2088# 0.029187f
C133 drain_right.n6 a_n1472_n2088# 0.015684f
C134 drain_right.n7 a_n1472_n2088# 0.037071f
C135 drain_right.n8 a_n1472_n2088# 0.016606f
C136 drain_right.n9 a_n1472_n2088# 0.1249f
C137 drain_right.t2 a_n1472_n2088# 0.060421f
C138 drain_right.n10 a_n1472_n2088# 0.027803f
C139 drain_right.n11 a_n1472_n2088# 0.021897f
C140 drain_right.n12 a_n1472_n2088# 0.015684f
C141 drain_right.n13 a_n1472_n2088# 0.694478f
C142 drain_right.n14 a_n1472_n2088# 0.029187f
C143 drain_right.n15 a_n1472_n2088# 0.015684f
C144 drain_right.n16 a_n1472_n2088# 0.016606f
C145 drain_right.n17 a_n1472_n2088# 0.037071f
C146 drain_right.n18 a_n1472_n2088# 0.037071f
C147 drain_right.n19 a_n1472_n2088# 0.016606f
C148 drain_right.n20 a_n1472_n2088# 0.015684f
C149 drain_right.n21 a_n1472_n2088# 0.029187f
C150 drain_right.n22 a_n1472_n2088# 0.029187f
C151 drain_right.n23 a_n1472_n2088# 0.015684f
C152 drain_right.n24 a_n1472_n2088# 0.016606f
C153 drain_right.n25 a_n1472_n2088# 0.037071f
C154 drain_right.n26 a_n1472_n2088# 0.080252f
C155 drain_right.n27 a_n1472_n2088# 0.016606f
C156 drain_right.n28 a_n1472_n2088# 0.015684f
C157 drain_right.n29 a_n1472_n2088# 0.067465f
C158 drain_right.n30 a_n1472_n2088# 0.066237f
C159 drain_right.t6 a_n1472_n2088# 0.138387f
C160 drain_right.t3 a_n1472_n2088# 0.138387f
C161 drain_right.n31 a_n1472_n2088# 1.15415f
C162 drain_right.n32 a_n1472_n2088# 0.410047f
C163 drain_right.t7 a_n1472_n2088# 0.138387f
C164 drain_right.t9 a_n1472_n2088# 0.138387f
C165 drain_right.n33 a_n1472_n2088# 1.15589f
C166 drain_right.n34 a_n1472_n2088# 1.20715f
C167 drain_right.t0 a_n1472_n2088# 0.138387f
C168 drain_right.t4 a_n1472_n2088# 0.138387f
C169 drain_right.n35 a_n1472_n2088# 1.15696f
C170 drain_right.t5 a_n1472_n2088# 0.138387f
C171 drain_right.t8 a_n1472_n2088# 0.138387f
C172 drain_right.n36 a_n1472_n2088# 1.15415f
C173 drain_right.n37 a_n1472_n2088# 0.687032f
C174 drain_right.n38 a_n1472_n2088# 0.041025f
C175 drain_right.n39 a_n1472_n2088# 0.029187f
C176 drain_right.n40 a_n1472_n2088# 0.015684f
C177 drain_right.n41 a_n1472_n2088# 0.037071f
C178 drain_right.n42 a_n1472_n2088# 0.016606f
C179 drain_right.n43 a_n1472_n2088# 0.029187f
C180 drain_right.n44 a_n1472_n2088# 0.015684f
C181 drain_right.n45 a_n1472_n2088# 0.037071f
C182 drain_right.n46 a_n1472_n2088# 0.016606f
C183 drain_right.n47 a_n1472_n2088# 0.1249f
C184 drain_right.t1 a_n1472_n2088# 0.060421f
C185 drain_right.n48 a_n1472_n2088# 0.027803f
C186 drain_right.n49 a_n1472_n2088# 0.021897f
C187 drain_right.n50 a_n1472_n2088# 0.015684f
C188 drain_right.n51 a_n1472_n2088# 0.694478f
C189 drain_right.n52 a_n1472_n2088# 0.029187f
C190 drain_right.n53 a_n1472_n2088# 0.015684f
C191 drain_right.n54 a_n1472_n2088# 0.016606f
C192 drain_right.n55 a_n1472_n2088# 0.037071f
C193 drain_right.n56 a_n1472_n2088# 0.037071f
C194 drain_right.n57 a_n1472_n2088# 0.016606f
C195 drain_right.n58 a_n1472_n2088# 0.015684f
C196 drain_right.n59 a_n1472_n2088# 0.029187f
C197 drain_right.n60 a_n1472_n2088# 0.029187f
C198 drain_right.n61 a_n1472_n2088# 0.015684f
C199 drain_right.n62 a_n1472_n2088# 0.016606f
C200 drain_right.n63 a_n1472_n2088# 0.037071f
C201 drain_right.n64 a_n1472_n2088# 0.080252f
C202 drain_right.n65 a_n1472_n2088# 0.016606f
C203 drain_right.n66 a_n1472_n2088# 0.015684f
C204 drain_right.n67 a_n1472_n2088# 0.067465f
C205 drain_right.n68 a_n1472_n2088# 0.065057f
C206 drain_right.n69 a_n1472_n2088# 0.350772f
C207 source.n0 a_n1472_n2088# 0.044544f
C208 source.n1 a_n1472_n2088# 0.031691f
C209 source.n2 a_n1472_n2088# 0.017029f
C210 source.n3 a_n1472_n2088# 0.040251f
C211 source.n4 a_n1472_n2088# 0.018031f
C212 source.n5 a_n1472_n2088# 0.031691f
C213 source.n6 a_n1472_n2088# 0.017029f
C214 source.n7 a_n1472_n2088# 0.040251f
C215 source.n8 a_n1472_n2088# 0.018031f
C216 source.n9 a_n1472_n2088# 0.135614f
C217 source.t1 a_n1472_n2088# 0.065604f
C218 source.n10 a_n1472_n2088# 0.030188f
C219 source.n11 a_n1472_n2088# 0.023776f
C220 source.n12 a_n1472_n2088# 0.017029f
C221 source.n13 a_n1472_n2088# 0.754049f
C222 source.n14 a_n1472_n2088# 0.031691f
C223 source.n15 a_n1472_n2088# 0.017029f
C224 source.n16 a_n1472_n2088# 0.018031f
C225 source.n17 a_n1472_n2088# 0.040251f
C226 source.n18 a_n1472_n2088# 0.040251f
C227 source.n19 a_n1472_n2088# 0.018031f
C228 source.n20 a_n1472_n2088# 0.017029f
C229 source.n21 a_n1472_n2088# 0.031691f
C230 source.n22 a_n1472_n2088# 0.031691f
C231 source.n23 a_n1472_n2088# 0.017029f
C232 source.n24 a_n1472_n2088# 0.018031f
C233 source.n25 a_n1472_n2088# 0.040251f
C234 source.n26 a_n1472_n2088# 0.087136f
C235 source.n27 a_n1472_n2088# 0.018031f
C236 source.n28 a_n1472_n2088# 0.017029f
C237 source.n29 a_n1472_n2088# 0.073252f
C238 source.n30 a_n1472_n2088# 0.048756f
C239 source.n31 a_n1472_n2088# 0.767612f
C240 source.t9 a_n1472_n2088# 0.150258f
C241 source.t3 a_n1472_n2088# 0.150258f
C242 source.n32 a_n1472_n2088# 1.17022f
C243 source.n33 a_n1472_n2088# 0.407987f
C244 source.t6 a_n1472_n2088# 0.150258f
C245 source.t2 a_n1472_n2088# 0.150258f
C246 source.n34 a_n1472_n2088# 1.17022f
C247 source.n35 a_n1472_n2088# 0.428234f
C248 source.n36 a_n1472_n2088# 0.044544f
C249 source.n37 a_n1472_n2088# 0.031691f
C250 source.n38 a_n1472_n2088# 0.017029f
C251 source.n39 a_n1472_n2088# 0.040251f
C252 source.n40 a_n1472_n2088# 0.018031f
C253 source.n41 a_n1472_n2088# 0.031691f
C254 source.n42 a_n1472_n2088# 0.017029f
C255 source.n43 a_n1472_n2088# 0.040251f
C256 source.n44 a_n1472_n2088# 0.018031f
C257 source.n45 a_n1472_n2088# 0.135614f
C258 source.t14 a_n1472_n2088# 0.065604f
C259 source.n46 a_n1472_n2088# 0.030188f
C260 source.n47 a_n1472_n2088# 0.023776f
C261 source.n48 a_n1472_n2088# 0.017029f
C262 source.n49 a_n1472_n2088# 0.754049f
C263 source.n50 a_n1472_n2088# 0.031691f
C264 source.n51 a_n1472_n2088# 0.017029f
C265 source.n52 a_n1472_n2088# 0.018031f
C266 source.n53 a_n1472_n2088# 0.040251f
C267 source.n54 a_n1472_n2088# 0.040251f
C268 source.n55 a_n1472_n2088# 0.018031f
C269 source.n56 a_n1472_n2088# 0.017029f
C270 source.n57 a_n1472_n2088# 0.031691f
C271 source.n58 a_n1472_n2088# 0.031691f
C272 source.n59 a_n1472_n2088# 0.017029f
C273 source.n60 a_n1472_n2088# 0.018031f
C274 source.n61 a_n1472_n2088# 0.040251f
C275 source.n62 a_n1472_n2088# 0.087136f
C276 source.n63 a_n1472_n2088# 0.018031f
C277 source.n64 a_n1472_n2088# 0.017029f
C278 source.n65 a_n1472_n2088# 0.073252f
C279 source.n66 a_n1472_n2088# 0.048756f
C280 source.n67 a_n1472_n2088# 0.15823f
C281 source.t13 a_n1472_n2088# 0.150258f
C282 source.t10 a_n1472_n2088# 0.150258f
C283 source.n68 a_n1472_n2088# 1.17022f
C284 source.n69 a_n1472_n2088# 0.407987f
C285 source.t17 a_n1472_n2088# 0.150258f
C286 source.t19 a_n1472_n2088# 0.150258f
C287 source.n70 a_n1472_n2088# 1.17022f
C288 source.n71 a_n1472_n2088# 1.50106f
C289 source.t4 a_n1472_n2088# 0.150258f
C290 source.t0 a_n1472_n2088# 0.150258f
C291 source.n72 a_n1472_n2088# 1.17021f
C292 source.n73 a_n1472_n2088# 1.50107f
C293 source.t8 a_n1472_n2088# 0.150258f
C294 source.t5 a_n1472_n2088# 0.150258f
C295 source.n74 a_n1472_n2088# 1.17021f
C296 source.n75 a_n1472_n2088# 0.407995f
C297 source.n76 a_n1472_n2088# 0.044544f
C298 source.n77 a_n1472_n2088# 0.031691f
C299 source.n78 a_n1472_n2088# 0.017029f
C300 source.n79 a_n1472_n2088# 0.040251f
C301 source.n80 a_n1472_n2088# 0.018031f
C302 source.n81 a_n1472_n2088# 0.031691f
C303 source.n82 a_n1472_n2088# 0.017029f
C304 source.n83 a_n1472_n2088# 0.040251f
C305 source.n84 a_n1472_n2088# 0.018031f
C306 source.n85 a_n1472_n2088# 0.135614f
C307 source.t7 a_n1472_n2088# 0.065604f
C308 source.n86 a_n1472_n2088# 0.030188f
C309 source.n87 a_n1472_n2088# 0.023776f
C310 source.n88 a_n1472_n2088# 0.017029f
C311 source.n89 a_n1472_n2088# 0.754049f
C312 source.n90 a_n1472_n2088# 0.031691f
C313 source.n91 a_n1472_n2088# 0.017029f
C314 source.n92 a_n1472_n2088# 0.018031f
C315 source.n93 a_n1472_n2088# 0.040251f
C316 source.n94 a_n1472_n2088# 0.040251f
C317 source.n95 a_n1472_n2088# 0.018031f
C318 source.n96 a_n1472_n2088# 0.017029f
C319 source.n97 a_n1472_n2088# 0.031691f
C320 source.n98 a_n1472_n2088# 0.031691f
C321 source.n99 a_n1472_n2088# 0.017029f
C322 source.n100 a_n1472_n2088# 0.018031f
C323 source.n101 a_n1472_n2088# 0.040251f
C324 source.n102 a_n1472_n2088# 0.087136f
C325 source.n103 a_n1472_n2088# 0.018031f
C326 source.n104 a_n1472_n2088# 0.017029f
C327 source.n105 a_n1472_n2088# 0.073252f
C328 source.n106 a_n1472_n2088# 0.048756f
C329 source.n107 a_n1472_n2088# 0.15823f
C330 source.t16 a_n1472_n2088# 0.150258f
C331 source.t11 a_n1472_n2088# 0.150258f
C332 source.n108 a_n1472_n2088# 1.17021f
C333 source.n109 a_n1472_n2088# 0.428242f
C334 source.t15 a_n1472_n2088# 0.150258f
C335 source.t18 a_n1472_n2088# 0.150258f
C336 source.n110 a_n1472_n2088# 1.17021f
C337 source.n111 a_n1472_n2088# 0.407995f
C338 source.n112 a_n1472_n2088# 0.044544f
C339 source.n113 a_n1472_n2088# 0.031691f
C340 source.n114 a_n1472_n2088# 0.017029f
C341 source.n115 a_n1472_n2088# 0.040251f
C342 source.n116 a_n1472_n2088# 0.018031f
C343 source.n117 a_n1472_n2088# 0.031691f
C344 source.n118 a_n1472_n2088# 0.017029f
C345 source.n119 a_n1472_n2088# 0.040251f
C346 source.n120 a_n1472_n2088# 0.018031f
C347 source.n121 a_n1472_n2088# 0.135614f
C348 source.t12 a_n1472_n2088# 0.065604f
C349 source.n122 a_n1472_n2088# 0.030188f
C350 source.n123 a_n1472_n2088# 0.023776f
C351 source.n124 a_n1472_n2088# 0.017029f
C352 source.n125 a_n1472_n2088# 0.754049f
C353 source.n126 a_n1472_n2088# 0.031691f
C354 source.n127 a_n1472_n2088# 0.017029f
C355 source.n128 a_n1472_n2088# 0.018031f
C356 source.n129 a_n1472_n2088# 0.040251f
C357 source.n130 a_n1472_n2088# 0.040251f
C358 source.n131 a_n1472_n2088# 0.018031f
C359 source.n132 a_n1472_n2088# 0.017029f
C360 source.n133 a_n1472_n2088# 0.031691f
C361 source.n134 a_n1472_n2088# 0.031691f
C362 source.n135 a_n1472_n2088# 0.017029f
C363 source.n136 a_n1472_n2088# 0.018031f
C364 source.n137 a_n1472_n2088# 0.040251f
C365 source.n138 a_n1472_n2088# 0.087136f
C366 source.n139 a_n1472_n2088# 0.018031f
C367 source.n140 a_n1472_n2088# 0.017029f
C368 source.n141 a_n1472_n2088# 0.073252f
C369 source.n142 a_n1472_n2088# 0.048756f
C370 source.n143 a_n1472_n2088# 0.309395f
C371 source.n144 a_n1472_n2088# 1.29673f
C372 minus.n0 a_n1472_n2088# 0.053581f
C373 minus.t8 a_n1472_n2088# 0.282583f
C374 minus.t4 a_n1472_n2088# 0.274792f
C375 minus.t1 a_n1472_n2088# 0.274792f
C376 minus.n1 a_n1472_n2088# 0.022069f
C377 minus.t9 a_n1472_n2088# 0.274792f
C378 minus.n2 a_n1472_n2088# 0.126134f
C379 minus.t5 a_n1472_n2088# 0.282583f
C380 minus.n3 a_n1472_n2088# 0.142468f
C381 minus.n4 a_n1472_n2088# 0.117658f
C382 minus.n5 a_n1472_n2088# 0.053581f
C383 minus.n6 a_n1472_n2088# 0.143908f
C384 minus.n7 a_n1472_n2088# 0.022069f
C385 minus.n8 a_n1472_n2088# 0.126134f
C386 minus.n9 a_n1472_n2088# 0.142393f
C387 minus.n10 a_n1472_n2088# 1.40425f
C388 minus.n11 a_n1472_n2088# 0.053581f
C389 minus.t2 a_n1472_n2088# 0.274792f
C390 minus.t6 a_n1472_n2088# 0.274792f
C391 minus.n12 a_n1472_n2088# 0.022069f
C392 minus.t7 a_n1472_n2088# 0.282583f
C393 minus.t3 a_n1472_n2088# 0.274792f
C394 minus.n13 a_n1472_n2088# 0.126134f
C395 minus.n14 a_n1472_n2088# 0.142468f
C396 minus.n15 a_n1472_n2088# 0.117658f
C397 minus.n16 a_n1472_n2088# 0.053581f
C398 minus.n17 a_n1472_n2088# 0.143908f
C399 minus.n18 a_n1472_n2088# 0.022069f
C400 minus.n19 a_n1472_n2088# 0.126134f
C401 minus.t0 a_n1472_n2088# 0.282583f
C402 minus.n20 a_n1472_n2088# 0.142393f
C403 minus.n21 a_n1472_n2088# 0.348688f
C404 minus.n22 a_n1472_n2088# 1.7328f
.ends

