* NGSPICE file created from diffpair381.ext - technology: sky130A

.subckt diffpair381 minus drain_right drain_left source plus
X0 a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X1 a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X2 source minus drain_right a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X3 source plus drain_left a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X4 a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X5 drain_right minus source a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X6 drain_left plus source a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X7 drain_left plus source a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X8 source plus drain_left a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X9 a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X10 drain_right minus source a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X11 source minus drain_right a_n1334_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
.ends

