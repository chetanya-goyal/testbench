* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t25 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 source.t0 plus.t0 drain_left.t13 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X2 source.t21 minus.t1 drain_right.t12 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X3 drain_right.t11 minus.t2 source.t14 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X4 source.t15 minus.t3 drain_right.t10 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 drain_left.t12 plus.t1 source.t12 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X6 drain_left.t11 plus.t2 source.t2 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X7 a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X8 drain_right.t9 minus.t4 source.t20 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X9 drain_right.t8 minus.t5 source.t26 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X10 a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X11 a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X12 drain_left.t10 plus.t3 source.t8 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X13 drain_left.t9 plus.t4 source.t10 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X14 source.t6 plus.t5 drain_left.t8 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 drain_right.t7 minus.t6 source.t27 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X16 source.t13 plus.t6 drain_left.t7 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 source.t17 minus.t7 drain_right.t6 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X18 source.t7 plus.t7 drain_left.t6 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X19 drain_right.t5 minus.t8 source.t23 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X20 source.t9 plus.t8 drain_left.t5 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X21 source.t19 minus.t9 drain_right.t4 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X22 source.t18 minus.t10 drain_right.t3 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X23 drain_left.t4 plus.t9 source.t11 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X24 drain_left.t3 plus.t10 source.t4 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X25 drain_right.t2 minus.t11 source.t24 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X26 drain_right.t1 minus.t12 source.t16 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X27 a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X28 source.t22 minus.t13 drain_right.t0 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X29 drain_left.t2 plus.t11 source.t1 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X30 drain_left.t1 plus.t12 source.t3 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X31 source.t5 plus.t13 drain_left.t0 a_n1724_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n15 minus.t5 322.065
R1 minus.n3 minus.t8 322.065
R2 minus.n32 minus.t4 322.065
R3 minus.n20 minus.t0 322.065
R4 minus.n1 minus.t7 265.101
R5 minus.n14 minus.t1 265.101
R6 minus.n12 minus.t12 265.101
R7 minus.n6 minus.t2 265.101
R8 minus.n4 minus.t13 265.101
R9 minus.n18 minus.t3 265.101
R10 minus.n31 minus.t9 265.101
R11 minus.n29 minus.t11 265.101
R12 minus.n23 minus.t6 265.101
R13 minus.n21 minus.t10 265.101
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n15 minus.n14 35.055
R41 minus.n4 minus.n3 35.055
R42 minus.n21 minus.n20 35.055
R43 minus.n32 minus.n31 35.055
R44 minus.n34 minus.n16 28.1122
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 source.n50 source.n48 289.615
R62 source.n36 source.n34 289.615
R63 source.n2 source.n0 289.615
R64 source.n16 source.n14 289.615
R65 source.n51 source.n50 185
R66 source.n37 source.n36 185
R67 source.n3 source.n2 185
R68 source.n17 source.n16 185
R69 source.t20 source.n49 167.117
R70 source.t1 source.n35 167.117
R71 source.t3 source.n1 167.117
R72 source.t23 source.n15 167.117
R73 source.n9 source.n8 84.1169
R74 source.n11 source.n10 84.1169
R75 source.n13 source.n12 84.1169
R76 source.n23 source.n22 84.1169
R77 source.n25 source.n24 84.1169
R78 source.n27 source.n26 84.1169
R79 source.n47 source.n46 84.1168
R80 source.n45 source.n44 84.1168
R81 source.n43 source.n42 84.1168
R82 source.n33 source.n32 84.1168
R83 source.n31 source.n30 84.1168
R84 source.n29 source.n28 84.1168
R85 source.n50 source.t20 52.3082
R86 source.n36 source.t1 52.3082
R87 source.n2 source.t3 52.3082
R88 source.n16 source.t23 52.3082
R89 source.n55 source.n54 31.4096
R90 source.n41 source.n40 31.4096
R91 source.n7 source.n6 31.4096
R92 source.n21 source.n20 31.4096
R93 source.n29 source.n27 14.7982
R94 source.n46 source.t24 9.9005
R95 source.n46 source.t19 9.9005
R96 source.n44 source.t27 9.9005
R97 source.n44 source.t15 9.9005
R98 source.n42 source.t25 9.9005
R99 source.n42 source.t18 9.9005
R100 source.n32 source.t8 9.9005
R101 source.n32 source.t13 9.9005
R102 source.n30 source.t11 9.9005
R103 source.n30 source.t0 9.9005
R104 source.n28 source.t12 9.9005
R105 source.n28 source.t7 9.9005
R106 source.n8 source.t10 9.9005
R107 source.n8 source.t9 9.9005
R108 source.n10 source.t4 9.9005
R109 source.n10 source.t5 9.9005
R110 source.n12 source.t2 9.9005
R111 source.n12 source.t6 9.9005
R112 source.n22 source.t14 9.9005
R113 source.n22 source.t22 9.9005
R114 source.n24 source.t16 9.9005
R115 source.n24 source.t17 9.9005
R116 source.n26 source.t26 9.9005
R117 source.n26 source.t21 9.9005
R118 source.n51 source.n49 9.71174
R119 source.n37 source.n35 9.71174
R120 source.n3 source.n1 9.71174
R121 source.n17 source.n15 9.71174
R122 source.n54 source.n53 9.45567
R123 source.n40 source.n39 9.45567
R124 source.n6 source.n5 9.45567
R125 source.n20 source.n19 9.45567
R126 source.n53 source.n52 9.3005
R127 source.n39 source.n38 9.3005
R128 source.n5 source.n4 9.3005
R129 source.n19 source.n18 9.3005
R130 source.n56 source.n7 8.72059
R131 source.n54 source.n48 8.14595
R132 source.n40 source.n34 8.14595
R133 source.n6 source.n0 8.14595
R134 source.n20 source.n14 8.14595
R135 source.n52 source.n51 7.3702
R136 source.n38 source.n37 7.3702
R137 source.n4 source.n3 7.3702
R138 source.n18 source.n17 7.3702
R139 source.n52 source.n48 5.81868
R140 source.n38 source.n34 5.81868
R141 source.n4 source.n0 5.81868
R142 source.n18 source.n14 5.81868
R143 source.n56 source.n55 5.53498
R144 source.n53 source.n49 3.44771
R145 source.n39 source.n35 3.44771
R146 source.n5 source.n1 3.44771
R147 source.n19 source.n15 3.44771
R148 source.n21 source.n13 0.741879
R149 source.n43 source.n41 0.741879
R150 source.n27 source.n25 0.543603
R151 source.n25 source.n23 0.543603
R152 source.n23 source.n21 0.543603
R153 source.n13 source.n11 0.543603
R154 source.n11 source.n9 0.543603
R155 source.n9 source.n7 0.543603
R156 source.n31 source.n29 0.543603
R157 source.n33 source.n31 0.543603
R158 source.n41 source.n33 0.543603
R159 source.n45 source.n43 0.543603
R160 source.n47 source.n45 0.543603
R161 source.n55 source.n47 0.543603
R162 source source.n56 0.188
R163 drain_right.n2 drain_right.n0 289.615
R164 drain_right.n20 drain_right.n18 289.615
R165 drain_right.n3 drain_right.n2 185
R166 drain_right.n21 drain_right.n20 185
R167 drain_right.t13 drain_right.n1 167.117
R168 drain_right.t8 drain_right.n19 167.117
R169 drain_right.n15 drain_right.n13 101.338
R170 drain_right.n11 drain_right.n9 101.338
R171 drain_right.n15 drain_right.n14 100.796
R172 drain_right.n17 drain_right.n16 100.796
R173 drain_right.n11 drain_right.n10 100.796
R174 drain_right.n8 drain_right.n7 100.796
R175 drain_right.n2 drain_right.t13 52.3082
R176 drain_right.n20 drain_right.t8 52.3082
R177 drain_right.n8 drain_right.n6 48.6315
R178 drain_right.n25 drain_right.n24 48.0884
R179 drain_right drain_right.n12 22.3609
R180 drain_right.n9 drain_right.t4 9.9005
R181 drain_right.n9 drain_right.t9 9.9005
R182 drain_right.n10 drain_right.t10 9.9005
R183 drain_right.n10 drain_right.t2 9.9005
R184 drain_right.n7 drain_right.t3 9.9005
R185 drain_right.n7 drain_right.t7 9.9005
R186 drain_right.n13 drain_right.t0 9.9005
R187 drain_right.n13 drain_right.t5 9.9005
R188 drain_right.n14 drain_right.t6 9.9005
R189 drain_right.n14 drain_right.t11 9.9005
R190 drain_right.n16 drain_right.t12 9.9005
R191 drain_right.n16 drain_right.t1 9.9005
R192 drain_right.n3 drain_right.n1 9.71174
R193 drain_right.n21 drain_right.n19 9.71174
R194 drain_right.n6 drain_right.n5 9.45567
R195 drain_right.n24 drain_right.n23 9.45567
R196 drain_right.n5 drain_right.n4 9.3005
R197 drain_right.n23 drain_right.n22 9.3005
R198 drain_right.n6 drain_right.n0 8.14595
R199 drain_right.n24 drain_right.n18 8.14595
R200 drain_right.n4 drain_right.n3 7.3702
R201 drain_right.n22 drain_right.n21 7.3702
R202 drain_right drain_right.n25 5.92477
R203 drain_right.n4 drain_right.n0 5.81868
R204 drain_right.n22 drain_right.n18 5.81868
R205 drain_right.n5 drain_right.n1 3.44771
R206 drain_right.n23 drain_right.n19 3.44771
R207 drain_right.n25 drain_right.n17 0.543603
R208 drain_right.n17 drain_right.n15 0.543603
R209 drain_right.n12 drain_right.n8 0.352482
R210 drain_right.n12 drain_right.n11 0.0809298
R211 plus.n3 plus.t2 322.065
R212 plus.n15 plus.t12 322.065
R213 plus.n20 plus.t11 322.065
R214 plus.n32 plus.t1 322.065
R215 plus.n1 plus.t13 265.101
R216 plus.n4 plus.t5 265.101
R217 plus.n6 plus.t10 265.101
R218 plus.n12 plus.t4 265.101
R219 plus.n14 plus.t8 265.101
R220 plus.n18 plus.t0 265.101
R221 plus.n21 plus.t6 265.101
R222 plus.n23 plus.t3 265.101
R223 plus.n29 plus.t9 265.101
R224 plus.n31 plus.t7 265.101
R225 plus.n3 plus.n2 161.489
R226 plus.n20 plus.n19 161.489
R227 plus.n5 plus.n2 161.3
R228 plus.n8 plus.n7 161.3
R229 plus.n9 plus.n1 161.3
R230 plus.n11 plus.n10 161.3
R231 plus.n13 plus.n0 161.3
R232 plus.n16 plus.n15 161.3
R233 plus.n22 plus.n19 161.3
R234 plus.n25 plus.n24 161.3
R235 plus.n26 plus.n18 161.3
R236 plus.n28 plus.n27 161.3
R237 plus.n30 plus.n17 161.3
R238 plus.n33 plus.n32 161.3
R239 plus.n7 plus.n1 73.0308
R240 plus.n11 plus.n1 73.0308
R241 plus.n28 plus.n18 73.0308
R242 plus.n24 plus.n18 73.0308
R243 plus.n6 plus.n5 54.0429
R244 plus.n13 plus.n12 54.0429
R245 plus.n30 plus.n29 54.0429
R246 plus.n23 plus.n22 54.0429
R247 plus.n5 plus.n4 37.9763
R248 plus.n14 plus.n13 37.9763
R249 plus.n31 plus.n30 37.9763
R250 plus.n22 plus.n21 37.9763
R251 plus.n4 plus.n3 35.055
R252 plus.n15 plus.n14 35.055
R253 plus.n32 plus.n31 35.055
R254 plus.n21 plus.n20 35.055
R255 plus plus.n33 25.7812
R256 plus.n7 plus.n6 18.9884
R257 plus.n12 plus.n11 18.9884
R258 plus.n29 plus.n28 18.9884
R259 plus.n24 plus.n23 18.9884
R260 plus plus.n16 8.39255
R261 plus.n8 plus.n2 0.189894
R262 plus.n9 plus.n8 0.189894
R263 plus.n10 plus.n9 0.189894
R264 plus.n10 plus.n0 0.189894
R265 plus.n16 plus.n0 0.189894
R266 plus.n33 plus.n17 0.189894
R267 plus.n27 plus.n17 0.189894
R268 plus.n27 plus.n26 0.189894
R269 plus.n26 plus.n25 0.189894
R270 plus.n25 plus.n19 0.189894
R271 drain_left.n2 drain_left.n0 289.615
R272 drain_left.n15 drain_left.n13 289.615
R273 drain_left.n3 drain_left.n2 185
R274 drain_left.n16 drain_left.n15 185
R275 drain_left.t12 drain_left.n1 167.117
R276 drain_left.t11 drain_left.n14 167.117
R277 drain_left.n11 drain_left.n9 101.338
R278 drain_left.n25 drain_left.n24 100.796
R279 drain_left.n23 drain_left.n22 100.796
R280 drain_left.n21 drain_left.n20 100.796
R281 drain_left.n11 drain_left.n10 100.796
R282 drain_left.n8 drain_left.n7 100.796
R283 drain_left.n2 drain_left.t12 52.3082
R284 drain_left.n15 drain_left.t11 52.3082
R285 drain_left.n8 drain_left.n6 48.6315
R286 drain_left.n21 drain_left.n19 48.6315
R287 drain_left drain_left.n12 22.9142
R288 drain_left.n9 drain_left.t7 9.9005
R289 drain_left.n9 drain_left.t2 9.9005
R290 drain_left.n10 drain_left.t13 9.9005
R291 drain_left.n10 drain_left.t10 9.9005
R292 drain_left.n7 drain_left.t6 9.9005
R293 drain_left.n7 drain_left.t4 9.9005
R294 drain_left.n24 drain_left.t5 9.9005
R295 drain_left.n24 drain_left.t1 9.9005
R296 drain_left.n22 drain_left.t0 9.9005
R297 drain_left.n22 drain_left.t9 9.9005
R298 drain_left.n20 drain_left.t8 9.9005
R299 drain_left.n20 drain_left.t3 9.9005
R300 drain_left.n3 drain_left.n1 9.71174
R301 drain_left.n16 drain_left.n14 9.71174
R302 drain_left.n6 drain_left.n5 9.45567
R303 drain_left.n19 drain_left.n18 9.45567
R304 drain_left.n5 drain_left.n4 9.3005
R305 drain_left.n18 drain_left.n17 9.3005
R306 drain_left.n6 drain_left.n0 8.14595
R307 drain_left.n19 drain_left.n13 8.14595
R308 drain_left.n4 drain_left.n3 7.3702
R309 drain_left.n17 drain_left.n16 7.3702
R310 drain_left drain_left.n25 6.19632
R311 drain_left.n4 drain_left.n0 5.81868
R312 drain_left.n17 drain_left.n13 5.81868
R313 drain_left.n5 drain_left.n1 3.44771
R314 drain_left.n18 drain_left.n14 3.44771
R315 drain_left.n23 drain_left.n21 0.543603
R316 drain_left.n25 drain_left.n23 0.543603
R317 drain_left.n12 drain_left.n8 0.352482
R318 drain_left.n12 drain_left.n11 0.0809298
C0 plus minus 3.45514f
C1 minus source 1.46345f
C2 minus drain_right 1.27377f
C3 minus drain_left 0.178085f
C4 plus source 1.47752f
C5 plus drain_right 0.328674f
C6 plus drain_left 1.43992f
C7 source drain_right 6.87065f
C8 source drain_left 6.87304f
C9 drain_left drain_right 0.879696f
C10 drain_right a_n1724_n1288# 3.93216f
C11 drain_left a_n1724_n1288# 4.17774f
C12 source a_n1724_n1288# 2.545505f
C13 minus a_n1724_n1288# 5.899496f
C14 plus a_n1724_n1288# 6.532769f
C15 drain_left.n0 a_n1724_n1288# 0.035689f
C16 drain_left.n1 a_n1724_n1288# 0.078967f
C17 drain_left.t12 a_n1724_n1288# 0.059261f
C18 drain_left.n2 a_n1724_n1288# 0.061803f
C19 drain_left.n3 a_n1724_n1288# 0.019923f
C20 drain_left.n4 a_n1724_n1288# 0.013139f
C21 drain_left.n5 a_n1724_n1288# 0.174062f
C22 drain_left.n6 a_n1724_n1288# 0.057013f
C23 drain_left.t6 a_n1724_n1288# 0.038645f
C24 drain_left.t4 a_n1724_n1288# 0.038645f
C25 drain_left.n7 a_n1724_n1288# 0.242783f
C26 drain_left.n8 a_n1724_n1288# 0.347403f
C27 drain_left.t7 a_n1724_n1288# 0.038645f
C28 drain_left.t2 a_n1724_n1288# 0.038645f
C29 drain_left.n9 a_n1724_n1288# 0.244297f
C30 drain_left.t13 a_n1724_n1288# 0.038645f
C31 drain_left.t10 a_n1724_n1288# 0.038645f
C32 drain_left.n10 a_n1724_n1288# 0.242783f
C33 drain_left.n11 a_n1724_n1288# 0.5244f
C34 drain_left.n12 a_n1724_n1288# 0.664947f
C35 drain_left.n13 a_n1724_n1288# 0.035689f
C36 drain_left.n14 a_n1724_n1288# 0.078967f
C37 drain_left.t11 a_n1724_n1288# 0.059261f
C38 drain_left.n15 a_n1724_n1288# 0.061803f
C39 drain_left.n16 a_n1724_n1288# 0.019923f
C40 drain_left.n17 a_n1724_n1288# 0.013139f
C41 drain_left.n18 a_n1724_n1288# 0.174062f
C42 drain_left.n19 a_n1724_n1288# 0.057013f
C43 drain_left.t8 a_n1724_n1288# 0.038645f
C44 drain_left.t3 a_n1724_n1288# 0.038645f
C45 drain_left.n20 a_n1724_n1288# 0.242784f
C46 drain_left.n21 a_n1724_n1288# 0.36085f
C47 drain_left.t0 a_n1724_n1288# 0.038645f
C48 drain_left.t9 a_n1724_n1288# 0.038645f
C49 drain_left.n22 a_n1724_n1288# 0.242784f
C50 drain_left.n23 a_n1724_n1288# 0.272735f
C51 drain_left.t5 a_n1724_n1288# 0.038645f
C52 drain_left.t1 a_n1724_n1288# 0.038645f
C53 drain_left.n24 a_n1724_n1288# 0.242784f
C54 drain_left.n25 a_n1724_n1288# 0.476264f
C55 plus.n0 a_n1724_n1288# 0.029655f
C56 plus.t8 a_n1724_n1288# 0.052357f
C57 plus.t4 a_n1724_n1288# 0.052357f
C58 plus.t13 a_n1724_n1288# 0.052357f
C59 plus.n1 a_n1724_n1288# 0.046405f
C60 plus.n2 a_n1724_n1288# 0.069867f
C61 plus.t10 a_n1724_n1288# 0.052357f
C62 plus.t5 a_n1724_n1288# 0.052357f
C63 plus.t2 a_n1724_n1288# 0.05944f
C64 plus.n3 a_n1724_n1288# 0.045221f
C65 plus.n4 a_n1724_n1288# 0.036567f
C66 plus.n5 a_n1724_n1288# 0.012214f
C67 plus.n6 a_n1724_n1288# 0.036567f
C68 plus.n7 a_n1724_n1288# 0.012214f
C69 plus.n8 a_n1724_n1288# 0.029655f
C70 plus.n9 a_n1724_n1288# 0.029655f
C71 plus.n10 a_n1724_n1288# 0.029655f
C72 plus.n11 a_n1724_n1288# 0.012214f
C73 plus.n12 a_n1724_n1288# 0.036567f
C74 plus.n13 a_n1724_n1288# 0.012214f
C75 plus.n14 a_n1724_n1288# 0.036567f
C76 plus.t12 a_n1724_n1288# 0.05944f
C77 plus.n15 a_n1724_n1288# 0.045173f
C78 plus.n16 a_n1724_n1288# 0.214683f
C79 plus.n17 a_n1724_n1288# 0.029655f
C80 plus.t1 a_n1724_n1288# 0.05944f
C81 plus.t7 a_n1724_n1288# 0.052357f
C82 plus.t9 a_n1724_n1288# 0.052357f
C83 plus.t0 a_n1724_n1288# 0.052357f
C84 plus.n18 a_n1724_n1288# 0.046405f
C85 plus.n19 a_n1724_n1288# 0.069867f
C86 plus.t3 a_n1724_n1288# 0.052357f
C87 plus.t6 a_n1724_n1288# 0.052357f
C88 plus.t11 a_n1724_n1288# 0.05944f
C89 plus.n20 a_n1724_n1288# 0.045221f
C90 plus.n21 a_n1724_n1288# 0.036567f
C91 plus.n22 a_n1724_n1288# 0.012214f
C92 plus.n23 a_n1724_n1288# 0.036567f
C93 plus.n24 a_n1724_n1288# 0.012214f
C94 plus.n25 a_n1724_n1288# 0.029655f
C95 plus.n26 a_n1724_n1288# 0.029655f
C96 plus.n27 a_n1724_n1288# 0.029655f
C97 plus.n28 a_n1724_n1288# 0.012214f
C98 plus.n29 a_n1724_n1288# 0.036567f
C99 plus.n30 a_n1724_n1288# 0.012214f
C100 plus.n31 a_n1724_n1288# 0.036567f
C101 plus.n32 a_n1724_n1288# 0.045173f
C102 plus.n33 a_n1724_n1288# 0.659769f
C103 drain_right.n0 a_n1724_n1288# 0.036191f
C104 drain_right.n1 a_n1724_n1288# 0.080077f
C105 drain_right.t13 a_n1724_n1288# 0.060094f
C106 drain_right.n2 a_n1724_n1288# 0.062671f
C107 drain_right.n3 a_n1724_n1288# 0.020203f
C108 drain_right.n4 a_n1724_n1288# 0.013324f
C109 drain_right.n5 a_n1724_n1288# 0.176509f
C110 drain_right.n6 a_n1724_n1288# 0.057815f
C111 drain_right.t3 a_n1724_n1288# 0.039189f
C112 drain_right.t7 a_n1724_n1288# 0.039189f
C113 drain_right.n7 a_n1724_n1288# 0.246195f
C114 drain_right.n8 a_n1724_n1288# 0.352287f
C115 drain_right.t4 a_n1724_n1288# 0.039189f
C116 drain_right.t9 a_n1724_n1288# 0.039189f
C117 drain_right.n9 a_n1724_n1288# 0.247731f
C118 drain_right.t10 a_n1724_n1288# 0.039189f
C119 drain_right.t2 a_n1724_n1288# 0.039189f
C120 drain_right.n10 a_n1724_n1288# 0.246195f
C121 drain_right.n11 a_n1724_n1288# 0.531772f
C122 drain_right.n12 a_n1724_n1288# 0.625661f
C123 drain_right.t0 a_n1724_n1288# 0.039189f
C124 drain_right.t5 a_n1724_n1288# 0.039189f
C125 drain_right.n13 a_n1724_n1288# 0.247732f
C126 drain_right.t6 a_n1724_n1288# 0.039189f
C127 drain_right.t11 a_n1724_n1288# 0.039189f
C128 drain_right.n14 a_n1724_n1288# 0.246197f
C129 drain_right.n15 a_n1724_n1288# 0.561589f
C130 drain_right.t12 a_n1724_n1288# 0.039189f
C131 drain_right.t1 a_n1724_n1288# 0.039189f
C132 drain_right.n16 a_n1724_n1288# 0.246197f
C133 drain_right.n17 a_n1724_n1288# 0.276569f
C134 drain_right.n18 a_n1724_n1288# 0.036191f
C135 drain_right.n19 a_n1724_n1288# 0.080077f
C136 drain_right.t8 a_n1724_n1288# 0.060094f
C137 drain_right.n20 a_n1724_n1288# 0.062671f
C138 drain_right.n21 a_n1724_n1288# 0.020203f
C139 drain_right.n22 a_n1724_n1288# 0.013324f
C140 drain_right.n23 a_n1724_n1288# 0.176509f
C141 drain_right.n24 a_n1724_n1288# 0.056806f
C142 drain_right.n25 a_n1724_n1288# 0.297221f
C143 source.n0 a_n1724_n1288# 0.043826f
C144 source.n1 a_n1724_n1288# 0.09697f
C145 source.t3 a_n1724_n1288# 0.072771f
C146 source.n2 a_n1724_n1288# 0.075892f
C147 source.n3 a_n1724_n1288# 0.024465f
C148 source.n4 a_n1724_n1288# 0.016135f
C149 source.n5 a_n1724_n1288# 0.213745f
C150 source.n6 a_n1724_n1288# 0.048043f
C151 source.n7 a_n1724_n1288# 0.453352f
C152 source.t10 a_n1724_n1288# 0.047456f
C153 source.t9 a_n1724_n1288# 0.047456f
C154 source.n8 a_n1724_n1288# 0.253697f
C155 source.n9 a_n1724_n1288# 0.338535f
C156 source.t4 a_n1724_n1288# 0.047456f
C157 source.t5 a_n1724_n1288# 0.047456f
C158 source.n10 a_n1724_n1288# 0.253697f
C159 source.n11 a_n1724_n1288# 0.338535f
C160 source.t2 a_n1724_n1288# 0.047456f
C161 source.t6 a_n1724_n1288# 0.047456f
C162 source.n12 a_n1724_n1288# 0.253697f
C163 source.n13 a_n1724_n1288# 0.357719f
C164 source.n14 a_n1724_n1288# 0.043826f
C165 source.n15 a_n1724_n1288# 0.09697f
C166 source.t23 a_n1724_n1288# 0.072771f
C167 source.n16 a_n1724_n1288# 0.075892f
C168 source.n17 a_n1724_n1288# 0.024465f
C169 source.n18 a_n1724_n1288# 0.016135f
C170 source.n19 a_n1724_n1288# 0.213745f
C171 source.n20 a_n1724_n1288# 0.048043f
C172 source.n21 a_n1724_n1288# 0.148996f
C173 source.t14 a_n1724_n1288# 0.047456f
C174 source.t22 a_n1724_n1288# 0.047456f
C175 source.n22 a_n1724_n1288# 0.253697f
C176 source.n23 a_n1724_n1288# 0.338535f
C177 source.t16 a_n1724_n1288# 0.047456f
C178 source.t17 a_n1724_n1288# 0.047456f
C179 source.n24 a_n1724_n1288# 0.253697f
C180 source.n25 a_n1724_n1288# 0.338535f
C181 source.t26 a_n1724_n1288# 0.047456f
C182 source.t21 a_n1724_n1288# 0.047456f
C183 source.n26 a_n1724_n1288# 0.253697f
C184 source.n27 a_n1724_n1288# 0.99456f
C185 source.t12 a_n1724_n1288# 0.047456f
C186 source.t7 a_n1724_n1288# 0.047456f
C187 source.n28 a_n1724_n1288# 0.253696f
C188 source.n29 a_n1724_n1288# 0.994562f
C189 source.t11 a_n1724_n1288# 0.047456f
C190 source.t0 a_n1724_n1288# 0.047456f
C191 source.n30 a_n1724_n1288# 0.253696f
C192 source.n31 a_n1724_n1288# 0.338537f
C193 source.t8 a_n1724_n1288# 0.047456f
C194 source.t13 a_n1724_n1288# 0.047456f
C195 source.n32 a_n1724_n1288# 0.253696f
C196 source.n33 a_n1724_n1288# 0.338537f
C197 source.n34 a_n1724_n1288# 0.043826f
C198 source.n35 a_n1724_n1288# 0.09697f
C199 source.t1 a_n1724_n1288# 0.072771f
C200 source.n36 a_n1724_n1288# 0.075892f
C201 source.n37 a_n1724_n1288# 0.024465f
C202 source.n38 a_n1724_n1288# 0.016135f
C203 source.n39 a_n1724_n1288# 0.213745f
C204 source.n40 a_n1724_n1288# 0.048043f
C205 source.n41 a_n1724_n1288# 0.148996f
C206 source.t25 a_n1724_n1288# 0.047456f
C207 source.t18 a_n1724_n1288# 0.047456f
C208 source.n42 a_n1724_n1288# 0.253696f
C209 source.n43 a_n1724_n1288# 0.357721f
C210 source.t27 a_n1724_n1288# 0.047456f
C211 source.t15 a_n1724_n1288# 0.047456f
C212 source.n44 a_n1724_n1288# 0.253696f
C213 source.n45 a_n1724_n1288# 0.338537f
C214 source.t24 a_n1724_n1288# 0.047456f
C215 source.t19 a_n1724_n1288# 0.047456f
C216 source.n46 a_n1724_n1288# 0.253696f
C217 source.n47 a_n1724_n1288# 0.338537f
C218 source.n48 a_n1724_n1288# 0.043826f
C219 source.n49 a_n1724_n1288# 0.09697f
C220 source.t20 a_n1724_n1288# 0.072771f
C221 source.n50 a_n1724_n1288# 0.075892f
C222 source.n51 a_n1724_n1288# 0.024465f
C223 source.n52 a_n1724_n1288# 0.016135f
C224 source.n53 a_n1724_n1288# 0.213745f
C225 source.n54 a_n1724_n1288# 0.048043f
C226 source.n55 a_n1724_n1288# 0.292222f
C227 source.n56 a_n1724_n1288# 0.742364f
C228 minus.n0 a_n1724_n1288# 0.029155f
C229 minus.t5 a_n1724_n1288# 0.058438f
C230 minus.t1 a_n1724_n1288# 0.051476f
C231 minus.t12 a_n1724_n1288# 0.051476f
C232 minus.t7 a_n1724_n1288# 0.051476f
C233 minus.n1 a_n1724_n1288# 0.045623f
C234 minus.n2 a_n1724_n1288# 0.06869f
C235 minus.t2 a_n1724_n1288# 0.051476f
C236 minus.t13 a_n1724_n1288# 0.051476f
C237 minus.t8 a_n1724_n1288# 0.058438f
C238 minus.n3 a_n1724_n1288# 0.044459f
C239 minus.n4 a_n1724_n1288# 0.035951f
C240 minus.n5 a_n1724_n1288# 0.012009f
C241 minus.n6 a_n1724_n1288# 0.035951f
C242 minus.n7 a_n1724_n1288# 0.012009f
C243 minus.n8 a_n1724_n1288# 0.029155f
C244 minus.n9 a_n1724_n1288# 0.029155f
C245 minus.n10 a_n1724_n1288# 0.029155f
C246 minus.n11 a_n1724_n1288# 0.012009f
C247 minus.n12 a_n1724_n1288# 0.035951f
C248 minus.n13 a_n1724_n1288# 0.012009f
C249 minus.n14 a_n1724_n1288# 0.035951f
C250 minus.n15 a_n1724_n1288# 0.044412f
C251 minus.n16 a_n1724_n1288# 0.678561f
C252 minus.n17 a_n1724_n1288# 0.029155f
C253 minus.t9 a_n1724_n1288# 0.051476f
C254 minus.t11 a_n1724_n1288# 0.051476f
C255 minus.t3 a_n1724_n1288# 0.051476f
C256 minus.n18 a_n1724_n1288# 0.045623f
C257 minus.n19 a_n1724_n1288# 0.06869f
C258 minus.t6 a_n1724_n1288# 0.051476f
C259 minus.t10 a_n1724_n1288# 0.051476f
C260 minus.t0 a_n1724_n1288# 0.058438f
C261 minus.n20 a_n1724_n1288# 0.044459f
C262 minus.n21 a_n1724_n1288# 0.035951f
C263 minus.n22 a_n1724_n1288# 0.012009f
C264 minus.n23 a_n1724_n1288# 0.035951f
C265 minus.n24 a_n1724_n1288# 0.012009f
C266 minus.n25 a_n1724_n1288# 0.029155f
C267 minus.n26 a_n1724_n1288# 0.029155f
C268 minus.n27 a_n1724_n1288# 0.029155f
C269 minus.n28 a_n1724_n1288# 0.012009f
C270 minus.n29 a_n1724_n1288# 0.035951f
C271 minus.n30 a_n1724_n1288# 0.012009f
C272 minus.n31 a_n1724_n1288# 0.035951f
C273 minus.t4 a_n1724_n1288# 0.058438f
C274 minus.n32 a_n1724_n1288# 0.044412f
C275 minus.n33 a_n1724_n1288# 0.193113f
C276 minus.n34 a_n1724_n1288# 0.83738f
.ends

