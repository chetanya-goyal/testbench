* NGSPICE file created from diffpair89.ext - technology: sky130A

.subckt diffpair89 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t28 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 source.t22 minus.t0 drain_right.t23 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 source.t19 minus.t1 drain_right.t22 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 drain_right.t21 minus.t2 source.t10 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 source.t35 plus.t1 drain_left.t22 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X5 drain_left.t21 plus.t2 source.t46 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X6 source.t14 minus.t3 drain_right.t20 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X7 drain_left.t20 plus.t3 source.t29 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X8 source.t42 plus.t4 drain_left.t19 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X9 drain_right.t19 minus.t4 source.t0 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X11 a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X12 drain_left.t18 plus.t5 source.t25 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 source.t27 plus.t6 drain_left.t17 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t1 minus.t5 drain_right.t18 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X16 source.t5 minus.t6 drain_right.t17 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_right.t16 minus.t7 source.t9 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X18 drain_right.t15 minus.t8 source.t13 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 drain_right.t14 minus.t9 source.t6 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X20 source.t36 plus.t7 drain_left.t16 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X21 drain_left.t15 plus.t8 source.t33 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X22 source.t16 minus.t10 drain_right.t13 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_right.t12 minus.t11 source.t7 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X24 drain_right.t11 minus.t12 source.t20 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X25 drain_right.t10 minus.t13 source.t23 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X26 source.t47 plus.t9 drain_left.t14 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X27 drain_left.t13 plus.t10 source.t39 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X28 source.t45 plus.t11 drain_left.t12 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X29 drain_right.t9 minus.t14 source.t15 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X30 drain_right.t8 minus.t15 source.t2 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X31 source.t24 plus.t12 drain_left.t11 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X32 source.t4 minus.t16 drain_right.t7 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X33 source.t11 minus.t17 drain_right.t6 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X34 source.t18 minus.t18 drain_right.t5 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X35 drain_left.t10 plus.t13 source.t34 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X36 source.t21 minus.t19 drain_right.t4 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X37 source.t32 plus.t14 drain_left.t9 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X38 drain_right.t3 minus.t20 source.t3 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X39 drain_left.t8 plus.t15 source.t26 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X40 drain_left.t7 plus.t16 source.t41 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X41 source.t43 plus.t17 drain_left.t6 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X42 source.t44 plus.t18 drain_left.t5 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X43 source.t8 minus.t21 drain_right.t2 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X44 a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X45 drain_right.t1 minus.t22 source.t12 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X46 source.t31 plus.t19 drain_left.t4 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X47 drain_left.t3 plus.t20 source.t37 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X48 drain_left.t2 plus.t21 source.t38 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X49 drain_left.t1 plus.t22 source.t40 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X50 source.t30 plus.t23 drain_left.t0 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X51 source.t17 minus.t23 drain_right.t0 a_n2406_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 plus.n6 plus.t11 577.67
R1 plus.n35 plus.t22 577.67
R2 plus.n45 plus.t15 577.67
R3 plus.n72 plus.t6 577.67
R4 plus.n7 plus.t21 530.201
R5 plus.n8 plus.t18 530.201
R6 plus.n14 plus.t13 530.201
R7 plus.n16 plus.t23 530.201
R8 plus.n17 plus.t20 530.201
R9 plus.n23 plus.t17 530.201
R10 plus.n25 plus.t10 530.201
R11 plus.n26 plus.t19 530.201
R12 plus.n32 plus.t16 530.201
R13 plus.n34 plus.t12 530.201
R14 plus.n47 plus.t9 530.201
R15 plus.n46 plus.t3 530.201
R16 plus.n53 plus.t1 530.201
R17 plus.n55 plus.t0 530.201
R18 plus.n43 plus.t7 530.201
R19 plus.n61 plus.t5 530.201
R20 plus.n63 plus.t4 530.201
R21 plus.n40 plus.t2 530.201
R22 plus.n69 plus.t14 530.201
R23 plus.n71 plus.t8 530.201
R24 plus.n10 plus.n6 161.489
R25 plus.n49 plus.n45 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n20 plus.n3 161.3
R32 plus.n22 plus.n21 161.3
R33 plus.n24 plus.n2 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n1 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n49 plus.n48 161.3
R40 plus.n50 plus.n44 161.3
R41 plus.n52 plus.n51 161.3
R42 plus.n54 plus.n42 161.3
R43 plus.n57 plus.n56 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n39 161.3
R47 plus.n65 plus.n64 161.3
R48 plus.n66 plus.n38 161.3
R49 plus.n68 plus.n67 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n13 plus.n5 73.0308
R53 plus.n22 plus.n3 73.0308
R54 plus.n31 plus.n1 73.0308
R55 plus.n68 plus.n38 73.0308
R56 plus.n60 plus.n41 73.0308
R57 plus.n52 plus.n44 73.0308
R58 plus.n9 plus.n8 69.3793
R59 plus.n33 plus.n32 69.3793
R60 plus.n70 plus.n69 69.3793
R61 plus.n48 plus.n46 69.3793
R62 plus.n18 plus.n17 62.0763
R63 plus.n24 plus.n23 62.0763
R64 plus.n62 plus.n61 62.0763
R65 plus.n56 plus.n43 62.0763
R66 plus.n15 plus.n14 54.7732
R67 plus.n27 plus.n26 54.7732
R68 plus.n64 plus.n40 54.7732
R69 plus.n54 plus.n53 54.7732
R70 plus.n7 plus.n6 47.4702
R71 plus.n35 plus.n34 47.4702
R72 plus.n72 plus.n71 47.4702
R73 plus.n47 plus.n45 47.4702
R74 plus.n16 plus.n15 40.1672
R75 plus.n27 plus.n25 40.1672
R76 plus.n64 plus.n63 40.1672
R77 plus.n55 plus.n54 40.1672
R78 plus.n18 plus.n16 32.8641
R79 plus.n25 plus.n24 32.8641
R80 plus.n63 plus.n62 32.8641
R81 plus.n56 plus.n55 32.8641
R82 plus plus.n73 28.3513
R83 plus.n9 plus.n7 25.5611
R84 plus.n34 plus.n33 25.5611
R85 plus.n71 plus.n70 25.5611
R86 plus.n48 plus.n47 25.5611
R87 plus.n14 plus.n13 18.2581
R88 plus.n26 plus.n1 18.2581
R89 plus.n40 plus.n38 18.2581
R90 plus.n53 plus.n52 18.2581
R91 plus.n17 plus.n3 10.955
R92 plus.n23 plus.n22 10.955
R93 plus.n61 plus.n60 10.955
R94 plus.n43 plus.n41 10.955
R95 plus plus.n36 8.37929
R96 plus.n8 plus.n5 3.65202
R97 plus.n32 plus.n31 3.65202
R98 plus.n69 plus.n68 3.65202
R99 plus.n46 plus.n44 3.65202
R100 plus.n11 plus.n10 0.189894
R101 plus.n12 plus.n11 0.189894
R102 plus.n12 plus.n4 0.189894
R103 plus.n19 plus.n4 0.189894
R104 plus.n20 plus.n19 0.189894
R105 plus.n21 plus.n20 0.189894
R106 plus.n21 plus.n2 0.189894
R107 plus.n28 plus.n2 0.189894
R108 plus.n29 plus.n28 0.189894
R109 plus.n30 plus.n29 0.189894
R110 plus.n30 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n67 plus.n37 0.189894
R114 plus.n67 plus.n66 0.189894
R115 plus.n66 plus.n65 0.189894
R116 plus.n65 plus.n39 0.189894
R117 plus.n59 plus.n39 0.189894
R118 plus.n59 plus.n58 0.189894
R119 plus.n58 plus.n57 0.189894
R120 plus.n57 plus.n42 0.189894
R121 plus.n51 plus.n42 0.189894
R122 plus.n51 plus.n50 0.189894
R123 plus.n50 plus.n49 0.189894
R124 source.n0 source.t40 99.1169
R125 source.n11 source.t45 99.1169
R126 source.n12 source.t9 99.1169
R127 source.n23 source.t11 99.1169
R128 source.n47 source.t6 99.1168
R129 source.n36 source.t19 99.1168
R130 source.n35 source.t26 99.1168
R131 source.n24 source.t27 99.1168
R132 source.n2 source.n1 84.1169
R133 source.n4 source.n3 84.1169
R134 source.n6 source.n5 84.1169
R135 source.n8 source.n7 84.1169
R136 source.n10 source.n9 84.1169
R137 source.n14 source.n13 84.1169
R138 source.n16 source.n15 84.1169
R139 source.n18 source.n17 84.1169
R140 source.n20 source.n19 84.1169
R141 source.n22 source.n21 84.1169
R142 source.n46 source.n45 84.1168
R143 source.n44 source.n43 84.1168
R144 source.n42 source.n41 84.1168
R145 source.n40 source.n39 84.1168
R146 source.n38 source.n37 84.1168
R147 source.n34 source.n33 84.1168
R148 source.n32 source.n31 84.1168
R149 source.n30 source.n29 84.1168
R150 source.n28 source.n27 84.1168
R151 source.n26 source.n25 84.1168
R152 source.n45 source.t10 15.0005
R153 source.n45 source.t17 15.0005
R154 source.n43 source.t7 15.0005
R155 source.n43 source.t14 15.0005
R156 source.n41 source.t12 15.0005
R157 source.n41 source.t18 15.0005
R158 source.n39 source.t0 15.0005
R159 source.n39 source.t22 15.0005
R160 source.n37 source.t23 15.0005
R161 source.n37 source.t5 15.0005
R162 source.n33 source.t29 15.0005
R163 source.n33 source.t47 15.0005
R164 source.n31 source.t28 15.0005
R165 source.n31 source.t35 15.0005
R166 source.n29 source.t25 15.0005
R167 source.n29 source.t36 15.0005
R168 source.n27 source.t46 15.0005
R169 source.n27 source.t42 15.0005
R170 source.n25 source.t33 15.0005
R171 source.n25 source.t32 15.0005
R172 source.n1 source.t41 15.0005
R173 source.n1 source.t24 15.0005
R174 source.n3 source.t39 15.0005
R175 source.n3 source.t31 15.0005
R176 source.n5 source.t37 15.0005
R177 source.n5 source.t43 15.0005
R178 source.n7 source.t34 15.0005
R179 source.n7 source.t30 15.0005
R180 source.n9 source.t38 15.0005
R181 source.n9 source.t44 15.0005
R182 source.n13 source.t15 15.0005
R183 source.n13 source.t1 15.0005
R184 source.n15 source.t13 15.0005
R185 source.n15 source.t16 15.0005
R186 source.n17 source.t2 15.0005
R187 source.n17 source.t21 15.0005
R188 source.n19 source.t20 15.0005
R189 source.n19 source.t4 15.0005
R190 source.n21 source.t3 15.0005
R191 source.n21 source.t8 15.0005
R192 source.n24 source.n23 14.2723
R193 source.n48 source.n0 8.72921
R194 source.n48 source.n47 5.5436
R195 source.n23 source.n22 0.560845
R196 source.n22 source.n20 0.560845
R197 source.n20 source.n18 0.560845
R198 source.n18 source.n16 0.560845
R199 source.n16 source.n14 0.560845
R200 source.n14 source.n12 0.560845
R201 source.n11 source.n10 0.560845
R202 source.n10 source.n8 0.560845
R203 source.n8 source.n6 0.560845
R204 source.n6 source.n4 0.560845
R205 source.n4 source.n2 0.560845
R206 source.n2 source.n0 0.560845
R207 source.n26 source.n24 0.560845
R208 source.n28 source.n26 0.560845
R209 source.n30 source.n28 0.560845
R210 source.n32 source.n30 0.560845
R211 source.n34 source.n32 0.560845
R212 source.n35 source.n34 0.560845
R213 source.n38 source.n36 0.560845
R214 source.n40 source.n38 0.560845
R215 source.n42 source.n40 0.560845
R216 source.n44 source.n42 0.560845
R217 source.n46 source.n44 0.560845
R218 source.n47 source.n46 0.560845
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 101.356
R223 drain_left.n7 drain_left.n5 101.356
R224 drain_left.n2 drain_left.n0 101.356
R225 drain_left.n21 drain_left.n20 100.796
R226 drain_left.n19 drain_left.n18 100.796
R227 drain_left.n17 drain_left.n16 100.796
R228 drain_left.n15 drain_left.n14 100.796
R229 drain_left.n13 drain_left.n12 100.796
R230 drain_left.n7 drain_left.n6 100.796
R231 drain_left.n9 drain_left.n8 100.796
R232 drain_left.n4 drain_left.n3 100.796
R233 drain_left.n2 drain_left.n1 100.796
R234 drain_left drain_left.n10 25.1146
R235 drain_left.n5 drain_left.t14 15.0005
R236 drain_left.n5 drain_left.t8 15.0005
R237 drain_left.n6 drain_left.t22 15.0005
R238 drain_left.n6 drain_left.t20 15.0005
R239 drain_left.n8 drain_left.t16 15.0005
R240 drain_left.n8 drain_left.t23 15.0005
R241 drain_left.n3 drain_left.t19 15.0005
R242 drain_left.n3 drain_left.t18 15.0005
R243 drain_left.n1 drain_left.t9 15.0005
R244 drain_left.n1 drain_left.t21 15.0005
R245 drain_left.n0 drain_left.t17 15.0005
R246 drain_left.n0 drain_left.t15 15.0005
R247 drain_left.n20 drain_left.t11 15.0005
R248 drain_left.n20 drain_left.t1 15.0005
R249 drain_left.n18 drain_left.t4 15.0005
R250 drain_left.n18 drain_left.t7 15.0005
R251 drain_left.n16 drain_left.t6 15.0005
R252 drain_left.n16 drain_left.t13 15.0005
R253 drain_left.n14 drain_left.t0 15.0005
R254 drain_left.n14 drain_left.t3 15.0005
R255 drain_left.n12 drain_left.t5 15.0005
R256 drain_left.n12 drain_left.t10 15.0005
R257 drain_left.n11 drain_left.t12 15.0005
R258 drain_left.n11 drain_left.t2 15.0005
R259 drain_left drain_left.n21 6.21356
R260 drain_left.n9 drain_left.n7 0.560845
R261 drain_left.n4 drain_left.n2 0.560845
R262 drain_left.n15 drain_left.n13 0.560845
R263 drain_left.n17 drain_left.n15 0.560845
R264 drain_left.n19 drain_left.n17 0.560845
R265 drain_left.n21 drain_left.n19 0.560845
R266 drain_left.n10 drain_left.n9 0.225326
R267 drain_left.n10 drain_left.n4 0.225326
R268 minus.n35 minus.t17 577.67
R269 minus.n8 minus.t7 577.67
R270 minus.n72 minus.t9 577.67
R271 minus.n43 minus.t1 577.67
R272 minus.n34 minus.t20 530.201
R273 minus.n32 minus.t21 530.201
R274 minus.n3 minus.t12 530.201
R275 minus.n26 minus.t16 530.201
R276 minus.n24 minus.t15 530.201
R277 minus.n6 minus.t19 530.201
R278 minus.n18 minus.t8 530.201
R279 minus.n16 minus.t10 530.201
R280 minus.n9 minus.t14 530.201
R281 minus.n10 minus.t5 530.201
R282 minus.n71 minus.t23 530.201
R283 minus.n69 minus.t2 530.201
R284 minus.n63 minus.t3 530.201
R285 minus.n62 minus.t11 530.201
R286 minus.n60 minus.t18 530.201
R287 minus.n54 minus.t22 530.201
R288 minus.n53 minus.t0 530.201
R289 minus.n51 minus.t4 530.201
R290 minus.n45 minus.t6 530.201
R291 minus.n44 minus.t13 530.201
R292 minus.n12 minus.n8 161.489
R293 minus.n47 minus.n43 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n31 minus.n30 161.3
R297 minus.n29 minus.n1 161.3
R298 minus.n28 minus.n27 161.3
R299 minus.n25 minus.n2 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n20 minus.n19 161.3
R303 minus.n17 minus.n5 161.3
R304 minus.n15 minus.n14 161.3
R305 minus.n13 minus.n7 161.3
R306 minus.n12 minus.n11 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n68 minus.n67 161.3
R310 minus.n66 minus.n38 161.3
R311 minus.n65 minus.n64 161.3
R312 minus.n61 minus.n39 161.3
R313 minus.n59 minus.n58 161.3
R314 minus.n57 minus.n40 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n52 minus.n41 161.3
R317 minus.n50 minus.n49 161.3
R318 minus.n48 minus.n42 161.3
R319 minus.n47 minus.n46 161.3
R320 minus.n31 minus.n1 73.0308
R321 minus.n23 minus.n4 73.0308
R322 minus.n15 minus.n7 73.0308
R323 minus.n50 minus.n42 73.0308
R324 minus.n59 minus.n40 73.0308
R325 minus.n68 minus.n38 73.0308
R326 minus.n33 minus.n32 69.3793
R327 minus.n11 minus.n9 69.3793
R328 minus.n46 minus.n45 69.3793
R329 minus.n70 minus.n69 69.3793
R330 minus.n25 minus.n24 62.0763
R331 minus.n19 minus.n6 62.0763
R332 minus.n55 minus.n54 62.0763
R333 minus.n61 minus.n60 62.0763
R334 minus.n27 minus.n3 54.7732
R335 minus.n17 minus.n16 54.7732
R336 minus.n52 minus.n51 54.7732
R337 minus.n64 minus.n63 54.7732
R338 minus.n35 minus.n34 47.4702
R339 minus.n10 minus.n8 47.4702
R340 minus.n44 minus.n43 47.4702
R341 minus.n72 minus.n71 47.4702
R342 minus.n27 minus.n26 40.1672
R343 minus.n18 minus.n17 40.1672
R344 minus.n53 minus.n52 40.1672
R345 minus.n64 minus.n62 40.1672
R346 minus.n26 minus.n25 32.8641
R347 minus.n19 minus.n18 32.8641
R348 minus.n55 minus.n53 32.8641
R349 minus.n62 minus.n61 32.8641
R350 minus.n74 minus.n36 30.6823
R351 minus.n34 minus.n33 25.5611
R352 minus.n11 minus.n10 25.5611
R353 minus.n46 minus.n44 25.5611
R354 minus.n71 minus.n70 25.5611
R355 minus.n3 minus.n1 18.2581
R356 minus.n16 minus.n15 18.2581
R357 minus.n51 minus.n50 18.2581
R358 minus.n63 minus.n38 18.2581
R359 minus.n24 minus.n23 10.955
R360 minus.n6 minus.n4 10.955
R361 minus.n54 minus.n40 10.955
R362 minus.n60 minus.n59 10.955
R363 minus.n74 minus.n73 6.52323
R364 minus.n32 minus.n31 3.65202
R365 minus.n9 minus.n7 3.65202
R366 minus.n45 minus.n42 3.65202
R367 minus.n69 minus.n68 3.65202
R368 minus.n36 minus.n0 0.189894
R369 minus.n30 minus.n0 0.189894
R370 minus.n30 minus.n29 0.189894
R371 minus.n29 minus.n28 0.189894
R372 minus.n28 minus.n2 0.189894
R373 minus.n22 minus.n2 0.189894
R374 minus.n22 minus.n21 0.189894
R375 minus.n21 minus.n20 0.189894
R376 minus.n20 minus.n5 0.189894
R377 minus.n14 minus.n5 0.189894
R378 minus.n14 minus.n13 0.189894
R379 minus.n13 minus.n12 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n49 minus.n48 0.189894
R382 minus.n49 minus.n41 0.189894
R383 minus.n56 minus.n41 0.189894
R384 minus.n57 minus.n56 0.189894
R385 minus.n58 minus.n57 0.189894
R386 minus.n58 minus.n39 0.189894
R387 minus.n65 minus.n39 0.189894
R388 minus.n66 minus.n65 0.189894
R389 minus.n67 minus.n66 0.189894
R390 minus.n67 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 101.356
R394 drain_right.n7 drain_right.n5 101.356
R395 drain_right.n2 drain_right.n0 101.356
R396 drain_right.n13 drain_right.n12 100.796
R397 drain_right.n15 drain_right.n14 100.796
R398 drain_right.n17 drain_right.n16 100.796
R399 drain_right.n19 drain_right.n18 100.796
R400 drain_right.n21 drain_right.n20 100.796
R401 drain_right.n7 drain_right.n6 100.796
R402 drain_right.n9 drain_right.n8 100.796
R403 drain_right.n4 drain_right.n3 100.796
R404 drain_right.n2 drain_right.n1 100.796
R405 drain_right drain_right.n10 24.5614
R406 drain_right.n5 drain_right.t0 15.0005
R407 drain_right.n5 drain_right.t14 15.0005
R408 drain_right.n6 drain_right.t20 15.0005
R409 drain_right.n6 drain_right.t21 15.0005
R410 drain_right.n8 drain_right.t5 15.0005
R411 drain_right.n8 drain_right.t12 15.0005
R412 drain_right.n3 drain_right.t23 15.0005
R413 drain_right.n3 drain_right.t1 15.0005
R414 drain_right.n1 drain_right.t17 15.0005
R415 drain_right.n1 drain_right.t19 15.0005
R416 drain_right.n0 drain_right.t22 15.0005
R417 drain_right.n0 drain_right.t10 15.0005
R418 drain_right.n11 drain_right.t18 15.0005
R419 drain_right.n11 drain_right.t16 15.0005
R420 drain_right.n12 drain_right.t13 15.0005
R421 drain_right.n12 drain_right.t9 15.0005
R422 drain_right.n14 drain_right.t4 15.0005
R423 drain_right.n14 drain_right.t15 15.0005
R424 drain_right.n16 drain_right.t7 15.0005
R425 drain_right.n16 drain_right.t8 15.0005
R426 drain_right.n18 drain_right.t2 15.0005
R427 drain_right.n18 drain_right.t11 15.0005
R428 drain_right.n20 drain_right.t6 15.0005
R429 drain_right.n20 drain_right.t3 15.0005
R430 drain_right drain_right.n21 6.21356
R431 drain_right.n9 drain_right.n7 0.560845
R432 drain_right.n4 drain_right.n2 0.560845
R433 drain_right.n21 drain_right.n19 0.560845
R434 drain_right.n19 drain_right.n17 0.560845
R435 drain_right.n17 drain_right.n15 0.560845
R436 drain_right.n15 drain_right.n13 0.560845
R437 drain_right.n10 drain_right.n9 0.225326
R438 drain_right.n10 drain_right.n4 0.225326
C0 drain_left minus 0.177738f
C1 drain_right minus 1.37585f
C2 plus source 1.58538f
C3 drain_left source 10.8098f
C4 drain_right source 10.8105f
C5 minus source 1.57142f
C6 drain_left plus 1.61355f
C7 plus drain_right 0.399127f
C8 drain_left drain_right 1.29455f
C9 plus minus 4.29827f
C10 drain_right a_n2406_n1288# 4.68345f
C11 drain_left a_n2406_n1288# 5.00789f
C12 source a_n2406_n1288# 3.490712f
C13 minus a_n2406_n1288# 8.104816f
C14 plus a_n2406_n1288# 8.874544f
C15 drain_right.t22 a_n2406_n1288# 0.059991f
C16 drain_right.t10 a_n2406_n1288# 0.059991f
C17 drain_right.n0 a_n2406_n1288# 0.291152f
C18 drain_right.t17 a_n2406_n1288# 0.059991f
C19 drain_right.t19 a_n2406_n1288# 0.059991f
C20 drain_right.n1 a_n2406_n1288# 0.289536f
C21 drain_right.n2 a_n2406_n1288# 0.572902f
C22 drain_right.t23 a_n2406_n1288# 0.059991f
C23 drain_right.t1 a_n2406_n1288# 0.059991f
C24 drain_right.n3 a_n2406_n1288# 0.289536f
C25 drain_right.n4 a_n2406_n1288# 0.257713f
C26 drain_right.t0 a_n2406_n1288# 0.059991f
C27 drain_right.t14 a_n2406_n1288# 0.059991f
C28 drain_right.n5 a_n2406_n1288# 0.291152f
C29 drain_right.t20 a_n2406_n1288# 0.059991f
C30 drain_right.t21 a_n2406_n1288# 0.059991f
C31 drain_right.n6 a_n2406_n1288# 0.289536f
C32 drain_right.n7 a_n2406_n1288# 0.572902f
C33 drain_right.t5 a_n2406_n1288# 0.059991f
C34 drain_right.t12 a_n2406_n1288# 0.059991f
C35 drain_right.n8 a_n2406_n1288# 0.289536f
C36 drain_right.n9 a_n2406_n1288# 0.257713f
C37 drain_right.n10 a_n2406_n1288# 0.805742f
C38 drain_right.t18 a_n2406_n1288# 0.059991f
C39 drain_right.t16 a_n2406_n1288# 0.059991f
C40 drain_right.n11 a_n2406_n1288# 0.291153f
C41 drain_right.t13 a_n2406_n1288# 0.059991f
C42 drain_right.t9 a_n2406_n1288# 0.059991f
C43 drain_right.n12 a_n2406_n1288# 0.289537f
C44 drain_right.n13 a_n2406_n1288# 0.5729f
C45 drain_right.t4 a_n2406_n1288# 0.059991f
C46 drain_right.t15 a_n2406_n1288# 0.059991f
C47 drain_right.n14 a_n2406_n1288# 0.289537f
C48 drain_right.n15 a_n2406_n1288# 0.282213f
C49 drain_right.t7 a_n2406_n1288# 0.059991f
C50 drain_right.t8 a_n2406_n1288# 0.059991f
C51 drain_right.n16 a_n2406_n1288# 0.289537f
C52 drain_right.n17 a_n2406_n1288# 0.282213f
C53 drain_right.t2 a_n2406_n1288# 0.059991f
C54 drain_right.t11 a_n2406_n1288# 0.059991f
C55 drain_right.n18 a_n2406_n1288# 0.289537f
C56 drain_right.n19 a_n2406_n1288# 0.282213f
C57 drain_right.t6 a_n2406_n1288# 0.059991f
C58 drain_right.t3 a_n2406_n1288# 0.059991f
C59 drain_right.n20 a_n2406_n1288# 0.289537f
C60 drain_right.n21 a_n2406_n1288# 0.491425f
C61 minus.n0 a_n2406_n1288# 0.029673f
C62 minus.t17 a_n2406_n1288# 0.028036f
C63 minus.t20 a_n2406_n1288# 0.026195f
C64 minus.t21 a_n2406_n1288# 0.026195f
C65 minus.n1 a_n2406_n1288# 0.01213f
C66 minus.n2 a_n2406_n1288# 0.029673f
C67 minus.t12 a_n2406_n1288# 0.026195f
C68 minus.n3 a_n2406_n1288# 0.022868f
C69 minus.t16 a_n2406_n1288# 0.026195f
C70 minus.t15 a_n2406_n1288# 0.026195f
C71 minus.n4 a_n2406_n1288# 0.011216f
C72 minus.n5 a_n2406_n1288# 0.029673f
C73 minus.t19 a_n2406_n1288# 0.026195f
C74 minus.n6 a_n2406_n1288# 0.022868f
C75 minus.t8 a_n2406_n1288# 0.026195f
C76 minus.t10 a_n2406_n1288# 0.026195f
C77 minus.n7 a_n2406_n1288# 0.010301f
C78 minus.t7 a_n2406_n1288# 0.028036f
C79 minus.n8 a_n2406_n1288# 0.033198f
C80 minus.t14 a_n2406_n1288# 0.026195f
C81 minus.n9 a_n2406_n1288# 0.022868f
C82 minus.t5 a_n2406_n1288# 0.026195f
C83 minus.n10 a_n2406_n1288# 0.022868f
C84 minus.n11 a_n2406_n1288# 0.012588f
C85 minus.n12 a_n2406_n1288# 0.064793f
C86 minus.n13 a_n2406_n1288# 0.029673f
C87 minus.n14 a_n2406_n1288# 0.029673f
C88 minus.n15 a_n2406_n1288# 0.01213f
C89 minus.n16 a_n2406_n1288# 0.022868f
C90 minus.n17 a_n2406_n1288# 0.012588f
C91 minus.n18 a_n2406_n1288# 0.022868f
C92 minus.n19 a_n2406_n1288# 0.012588f
C93 minus.n20 a_n2406_n1288# 0.029673f
C94 minus.n21 a_n2406_n1288# 0.029673f
C95 minus.n22 a_n2406_n1288# 0.029673f
C96 minus.n23 a_n2406_n1288# 0.011216f
C97 minus.n24 a_n2406_n1288# 0.022868f
C98 minus.n25 a_n2406_n1288# 0.012588f
C99 minus.n26 a_n2406_n1288# 0.022868f
C100 minus.n27 a_n2406_n1288# 0.012588f
C101 minus.n28 a_n2406_n1288# 0.029673f
C102 minus.n29 a_n2406_n1288# 0.029673f
C103 minus.n30 a_n2406_n1288# 0.029673f
C104 minus.n31 a_n2406_n1288# 0.010301f
C105 minus.n32 a_n2406_n1288# 0.022868f
C106 minus.n33 a_n2406_n1288# 0.012588f
C107 minus.n34 a_n2406_n1288# 0.022868f
C108 minus.n35 a_n2406_n1288# 0.033157f
C109 minus.n36 a_n2406_n1288# 0.802591f
C110 minus.n37 a_n2406_n1288# 0.029673f
C111 minus.t23 a_n2406_n1288# 0.026195f
C112 minus.t2 a_n2406_n1288# 0.026195f
C113 minus.n38 a_n2406_n1288# 0.01213f
C114 minus.n39 a_n2406_n1288# 0.029673f
C115 minus.t11 a_n2406_n1288# 0.026195f
C116 minus.t18 a_n2406_n1288# 0.026195f
C117 minus.n40 a_n2406_n1288# 0.011216f
C118 minus.n41 a_n2406_n1288# 0.029673f
C119 minus.t0 a_n2406_n1288# 0.026195f
C120 minus.t4 a_n2406_n1288# 0.026195f
C121 minus.n42 a_n2406_n1288# 0.010301f
C122 minus.t1 a_n2406_n1288# 0.028036f
C123 minus.n43 a_n2406_n1288# 0.033198f
C124 minus.t13 a_n2406_n1288# 0.026195f
C125 minus.n44 a_n2406_n1288# 0.022868f
C126 minus.t6 a_n2406_n1288# 0.026195f
C127 minus.n45 a_n2406_n1288# 0.022868f
C128 minus.n46 a_n2406_n1288# 0.012588f
C129 minus.n47 a_n2406_n1288# 0.064793f
C130 minus.n48 a_n2406_n1288# 0.029673f
C131 minus.n49 a_n2406_n1288# 0.029673f
C132 minus.n50 a_n2406_n1288# 0.01213f
C133 minus.n51 a_n2406_n1288# 0.022868f
C134 minus.n52 a_n2406_n1288# 0.012588f
C135 minus.n53 a_n2406_n1288# 0.022868f
C136 minus.t22 a_n2406_n1288# 0.026195f
C137 minus.n54 a_n2406_n1288# 0.022868f
C138 minus.n55 a_n2406_n1288# 0.012588f
C139 minus.n56 a_n2406_n1288# 0.029673f
C140 minus.n57 a_n2406_n1288# 0.029673f
C141 minus.n58 a_n2406_n1288# 0.029673f
C142 minus.n59 a_n2406_n1288# 0.011216f
C143 minus.n60 a_n2406_n1288# 0.022868f
C144 minus.n61 a_n2406_n1288# 0.012588f
C145 minus.n62 a_n2406_n1288# 0.022868f
C146 minus.t3 a_n2406_n1288# 0.026195f
C147 minus.n63 a_n2406_n1288# 0.022868f
C148 minus.n64 a_n2406_n1288# 0.012588f
C149 minus.n65 a_n2406_n1288# 0.029673f
C150 minus.n66 a_n2406_n1288# 0.029673f
C151 minus.n67 a_n2406_n1288# 0.029673f
C152 minus.n68 a_n2406_n1288# 0.010301f
C153 minus.n69 a_n2406_n1288# 0.022868f
C154 minus.n70 a_n2406_n1288# 0.012588f
C155 minus.n71 a_n2406_n1288# 0.022868f
C156 minus.t9 a_n2406_n1288# 0.028036f
C157 minus.n72 a_n2406_n1288# 0.033157f
C158 minus.n73 a_n2406_n1288# 0.195616f
C159 minus.n74 a_n2406_n1288# 0.988161f
C160 drain_left.t17 a_n2406_n1288# 0.059452f
C161 drain_left.t15 a_n2406_n1288# 0.059452f
C162 drain_left.n0 a_n2406_n1288# 0.288534f
C163 drain_left.t9 a_n2406_n1288# 0.059452f
C164 drain_left.t21 a_n2406_n1288# 0.059452f
C165 drain_left.n1 a_n2406_n1288# 0.286932f
C166 drain_left.n2 a_n2406_n1288# 0.56775f
C167 drain_left.t19 a_n2406_n1288# 0.059452f
C168 drain_left.t18 a_n2406_n1288# 0.059452f
C169 drain_left.n3 a_n2406_n1288# 0.286932f
C170 drain_left.n4 a_n2406_n1288# 0.255395f
C171 drain_left.t14 a_n2406_n1288# 0.059452f
C172 drain_left.t8 a_n2406_n1288# 0.059452f
C173 drain_left.n5 a_n2406_n1288# 0.288534f
C174 drain_left.t22 a_n2406_n1288# 0.059452f
C175 drain_left.t20 a_n2406_n1288# 0.059452f
C176 drain_left.n6 a_n2406_n1288# 0.286932f
C177 drain_left.n7 a_n2406_n1288# 0.56775f
C178 drain_left.t16 a_n2406_n1288# 0.059452f
C179 drain_left.t23 a_n2406_n1288# 0.059452f
C180 drain_left.n8 a_n2406_n1288# 0.286932f
C181 drain_left.n9 a_n2406_n1288# 0.255395f
C182 drain_left.n10 a_n2406_n1288# 0.846863f
C183 drain_left.t12 a_n2406_n1288# 0.059452f
C184 drain_left.t2 a_n2406_n1288# 0.059452f
C185 drain_left.n11 a_n2406_n1288# 0.288535f
C186 drain_left.t5 a_n2406_n1288# 0.059452f
C187 drain_left.t10 a_n2406_n1288# 0.059452f
C188 drain_left.n12 a_n2406_n1288# 0.286933f
C189 drain_left.n13 a_n2406_n1288# 0.567748f
C190 drain_left.t0 a_n2406_n1288# 0.059452f
C191 drain_left.t3 a_n2406_n1288# 0.059452f
C192 drain_left.n14 a_n2406_n1288# 0.286933f
C193 drain_left.n15 a_n2406_n1288# 0.279675f
C194 drain_left.t6 a_n2406_n1288# 0.059452f
C195 drain_left.t13 a_n2406_n1288# 0.059452f
C196 drain_left.n16 a_n2406_n1288# 0.286933f
C197 drain_left.n17 a_n2406_n1288# 0.279675f
C198 drain_left.t4 a_n2406_n1288# 0.059452f
C199 drain_left.t7 a_n2406_n1288# 0.059452f
C200 drain_left.n18 a_n2406_n1288# 0.286933f
C201 drain_left.n19 a_n2406_n1288# 0.279675f
C202 drain_left.t11 a_n2406_n1288# 0.059452f
C203 drain_left.t1 a_n2406_n1288# 0.059452f
C204 drain_left.n20 a_n2406_n1288# 0.286933f
C205 drain_left.n21 a_n2406_n1288# 0.487006f
C206 source.t40 a_n2406_n1288# 0.334096f
C207 source.n0 a_n2406_n1288# 0.636779f
C208 source.t41 a_n2406_n1288# 0.063633f
C209 source.t24 a_n2406_n1288# 0.063633f
C210 source.n1 a_n2406_n1288# 0.267788f
C211 source.n2 a_n2406_n1288# 0.302551f
C212 source.t39 a_n2406_n1288# 0.063633f
C213 source.t31 a_n2406_n1288# 0.063633f
C214 source.n3 a_n2406_n1288# 0.267788f
C215 source.n4 a_n2406_n1288# 0.302551f
C216 source.t37 a_n2406_n1288# 0.063633f
C217 source.t43 a_n2406_n1288# 0.063633f
C218 source.n5 a_n2406_n1288# 0.267788f
C219 source.n6 a_n2406_n1288# 0.302551f
C220 source.t34 a_n2406_n1288# 0.063633f
C221 source.t30 a_n2406_n1288# 0.063633f
C222 source.n7 a_n2406_n1288# 0.267788f
C223 source.n8 a_n2406_n1288# 0.302551f
C224 source.t38 a_n2406_n1288# 0.063633f
C225 source.t44 a_n2406_n1288# 0.063633f
C226 source.n9 a_n2406_n1288# 0.267788f
C227 source.n10 a_n2406_n1288# 0.302551f
C228 source.t45 a_n2406_n1288# 0.334096f
C229 source.n11 a_n2406_n1288# 0.343031f
C230 source.t9 a_n2406_n1288# 0.334096f
C231 source.n12 a_n2406_n1288# 0.343031f
C232 source.t15 a_n2406_n1288# 0.063633f
C233 source.t1 a_n2406_n1288# 0.063633f
C234 source.n13 a_n2406_n1288# 0.267788f
C235 source.n14 a_n2406_n1288# 0.302551f
C236 source.t13 a_n2406_n1288# 0.063633f
C237 source.t16 a_n2406_n1288# 0.063633f
C238 source.n15 a_n2406_n1288# 0.267788f
C239 source.n16 a_n2406_n1288# 0.302551f
C240 source.t2 a_n2406_n1288# 0.063633f
C241 source.t21 a_n2406_n1288# 0.063633f
C242 source.n17 a_n2406_n1288# 0.267788f
C243 source.n18 a_n2406_n1288# 0.302551f
C244 source.t20 a_n2406_n1288# 0.063633f
C245 source.t4 a_n2406_n1288# 0.063633f
C246 source.n19 a_n2406_n1288# 0.267788f
C247 source.n20 a_n2406_n1288# 0.302551f
C248 source.t3 a_n2406_n1288# 0.063633f
C249 source.t8 a_n2406_n1288# 0.063633f
C250 source.n21 a_n2406_n1288# 0.267788f
C251 source.n22 a_n2406_n1288# 0.302551f
C252 source.t11 a_n2406_n1288# 0.334096f
C253 source.n23 a_n2406_n1288# 0.884849f
C254 source.t27 a_n2406_n1288# 0.334095f
C255 source.n24 a_n2406_n1288# 0.884851f
C256 source.t33 a_n2406_n1288# 0.063633f
C257 source.t32 a_n2406_n1288# 0.063633f
C258 source.n25 a_n2406_n1288# 0.267787f
C259 source.n26 a_n2406_n1288# 0.302552f
C260 source.t46 a_n2406_n1288# 0.063633f
C261 source.t42 a_n2406_n1288# 0.063633f
C262 source.n27 a_n2406_n1288# 0.267787f
C263 source.n28 a_n2406_n1288# 0.302552f
C264 source.t25 a_n2406_n1288# 0.063633f
C265 source.t36 a_n2406_n1288# 0.063633f
C266 source.n29 a_n2406_n1288# 0.267787f
C267 source.n30 a_n2406_n1288# 0.302552f
C268 source.t28 a_n2406_n1288# 0.063633f
C269 source.t35 a_n2406_n1288# 0.063633f
C270 source.n31 a_n2406_n1288# 0.267787f
C271 source.n32 a_n2406_n1288# 0.302552f
C272 source.t29 a_n2406_n1288# 0.063633f
C273 source.t47 a_n2406_n1288# 0.063633f
C274 source.n33 a_n2406_n1288# 0.267787f
C275 source.n34 a_n2406_n1288# 0.302552f
C276 source.t26 a_n2406_n1288# 0.334095f
C277 source.n35 a_n2406_n1288# 0.343032f
C278 source.t19 a_n2406_n1288# 0.334095f
C279 source.n36 a_n2406_n1288# 0.343032f
C280 source.t23 a_n2406_n1288# 0.063633f
C281 source.t5 a_n2406_n1288# 0.063633f
C282 source.n37 a_n2406_n1288# 0.267787f
C283 source.n38 a_n2406_n1288# 0.302552f
C284 source.t0 a_n2406_n1288# 0.063633f
C285 source.t22 a_n2406_n1288# 0.063633f
C286 source.n39 a_n2406_n1288# 0.267787f
C287 source.n40 a_n2406_n1288# 0.302552f
C288 source.t12 a_n2406_n1288# 0.063633f
C289 source.t18 a_n2406_n1288# 0.063633f
C290 source.n41 a_n2406_n1288# 0.267787f
C291 source.n42 a_n2406_n1288# 0.302552f
C292 source.t7 a_n2406_n1288# 0.063633f
C293 source.t14 a_n2406_n1288# 0.063633f
C294 source.n43 a_n2406_n1288# 0.267787f
C295 source.n44 a_n2406_n1288# 0.302552f
C296 source.t10 a_n2406_n1288# 0.063633f
C297 source.t17 a_n2406_n1288# 0.063633f
C298 source.n45 a_n2406_n1288# 0.267787f
C299 source.n46 a_n2406_n1288# 0.302552f
C300 source.t6 a_n2406_n1288# 0.334095f
C301 source.n47 a_n2406_n1288# 0.494215f
C302 source.n48 a_n2406_n1288# 0.657606f
C303 plus.n0 a_n2406_n1288# 0.030093f
C304 plus.t12 a_n2406_n1288# 0.026565f
C305 plus.t16 a_n2406_n1288# 0.026565f
C306 plus.n1 a_n2406_n1288# 0.012302f
C307 plus.n2 a_n2406_n1288# 0.030093f
C308 plus.t10 a_n2406_n1288# 0.026565f
C309 plus.t17 a_n2406_n1288# 0.026565f
C310 plus.n3 a_n2406_n1288# 0.011374f
C311 plus.n4 a_n2406_n1288# 0.030093f
C312 plus.t23 a_n2406_n1288# 0.026565f
C313 plus.t13 a_n2406_n1288# 0.026565f
C314 plus.n5 a_n2406_n1288# 0.010447f
C315 plus.t11 a_n2406_n1288# 0.028433f
C316 plus.n6 a_n2406_n1288# 0.033668f
C317 plus.t21 a_n2406_n1288# 0.026565f
C318 plus.n7 a_n2406_n1288# 0.023192f
C319 plus.t18 a_n2406_n1288# 0.026565f
C320 plus.n8 a_n2406_n1288# 0.023192f
C321 plus.n9 a_n2406_n1288# 0.012766f
C322 plus.n10 a_n2406_n1288# 0.06571f
C323 plus.n11 a_n2406_n1288# 0.030093f
C324 plus.n12 a_n2406_n1288# 0.030093f
C325 plus.n13 a_n2406_n1288# 0.012302f
C326 plus.n14 a_n2406_n1288# 0.023192f
C327 plus.n15 a_n2406_n1288# 0.012766f
C328 plus.n16 a_n2406_n1288# 0.023192f
C329 plus.t20 a_n2406_n1288# 0.026565f
C330 plus.n17 a_n2406_n1288# 0.023192f
C331 plus.n18 a_n2406_n1288# 0.012766f
C332 plus.n19 a_n2406_n1288# 0.030093f
C333 plus.n20 a_n2406_n1288# 0.030093f
C334 plus.n21 a_n2406_n1288# 0.030093f
C335 plus.n22 a_n2406_n1288# 0.011374f
C336 plus.n23 a_n2406_n1288# 0.023192f
C337 plus.n24 a_n2406_n1288# 0.012766f
C338 plus.n25 a_n2406_n1288# 0.023192f
C339 plus.t19 a_n2406_n1288# 0.026565f
C340 plus.n26 a_n2406_n1288# 0.023192f
C341 plus.n27 a_n2406_n1288# 0.012766f
C342 plus.n28 a_n2406_n1288# 0.030093f
C343 plus.n29 a_n2406_n1288# 0.030093f
C344 plus.n30 a_n2406_n1288# 0.030093f
C345 plus.n31 a_n2406_n1288# 0.010447f
C346 plus.n32 a_n2406_n1288# 0.023192f
C347 plus.n33 a_n2406_n1288# 0.012766f
C348 plus.n34 a_n2406_n1288# 0.023192f
C349 plus.t22 a_n2406_n1288# 0.028433f
C350 plus.n35 a_n2406_n1288# 0.033626f
C351 plus.n36 a_n2406_n1288# 0.216865f
C352 plus.n37 a_n2406_n1288# 0.030093f
C353 plus.t6 a_n2406_n1288# 0.028433f
C354 plus.t8 a_n2406_n1288# 0.026565f
C355 plus.t14 a_n2406_n1288# 0.026565f
C356 plus.n38 a_n2406_n1288# 0.012302f
C357 plus.n39 a_n2406_n1288# 0.030093f
C358 plus.t2 a_n2406_n1288# 0.026565f
C359 plus.n40 a_n2406_n1288# 0.023192f
C360 plus.t4 a_n2406_n1288# 0.026565f
C361 plus.t5 a_n2406_n1288# 0.026565f
C362 plus.n41 a_n2406_n1288# 0.011374f
C363 plus.n42 a_n2406_n1288# 0.030093f
C364 plus.t7 a_n2406_n1288# 0.026565f
C365 plus.n43 a_n2406_n1288# 0.023192f
C366 plus.t0 a_n2406_n1288# 0.026565f
C367 plus.t1 a_n2406_n1288# 0.026565f
C368 plus.n44 a_n2406_n1288# 0.010447f
C369 plus.t15 a_n2406_n1288# 0.028433f
C370 plus.n45 a_n2406_n1288# 0.033668f
C371 plus.t3 a_n2406_n1288# 0.026565f
C372 plus.n46 a_n2406_n1288# 0.023192f
C373 plus.t9 a_n2406_n1288# 0.026565f
C374 plus.n47 a_n2406_n1288# 0.023192f
C375 plus.n48 a_n2406_n1288# 0.012766f
C376 plus.n49 a_n2406_n1288# 0.06571f
C377 plus.n50 a_n2406_n1288# 0.030093f
C378 plus.n51 a_n2406_n1288# 0.030093f
C379 plus.n52 a_n2406_n1288# 0.012302f
C380 plus.n53 a_n2406_n1288# 0.023192f
C381 plus.n54 a_n2406_n1288# 0.012766f
C382 plus.n55 a_n2406_n1288# 0.023192f
C383 plus.n56 a_n2406_n1288# 0.012766f
C384 plus.n57 a_n2406_n1288# 0.030093f
C385 plus.n58 a_n2406_n1288# 0.030093f
C386 plus.n59 a_n2406_n1288# 0.030093f
C387 plus.n60 a_n2406_n1288# 0.011374f
C388 plus.n61 a_n2406_n1288# 0.023192f
C389 plus.n62 a_n2406_n1288# 0.012766f
C390 plus.n63 a_n2406_n1288# 0.023192f
C391 plus.n64 a_n2406_n1288# 0.012766f
C392 plus.n65 a_n2406_n1288# 0.030093f
C393 plus.n66 a_n2406_n1288# 0.030093f
C394 plus.n67 a_n2406_n1288# 0.030093f
C395 plus.n68 a_n2406_n1288# 0.010447f
C396 plus.n69 a_n2406_n1288# 0.023192f
C397 plus.n70 a_n2406_n1288# 0.012766f
C398 plus.n71 a_n2406_n1288# 0.023192f
C399 plus.n72 a_n2406_n1288# 0.033626f
C400 plus.n73 a_n2406_n1288# 0.774517f
.ends

