* NGSPICE file created from diffpair584.ext - technology: sky130A

.subckt diffpair584 minus drain_right drain_left source plus
X0 source.t19 plus.t0 drain_left.t9 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X1 source.t18 plus.t1 drain_left.t0 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X2 drain_left.t2 plus.t2 source.t17 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X3 source.t0 minus.t0 drain_right.t9 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X4 drain_right.t8 minus.t1 source.t5 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X5 source.t3 minus.t2 drain_right.t7 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X6 source.t16 plus.t3 drain_left.t3 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X7 drain_left.t5 plus.t4 source.t15 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X8 a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X9 source.t9 minus.t3 drain_right.t6 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X10 drain_left.t4 plus.t5 source.t14 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X11 drain_right.t5 minus.t4 source.t2 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X12 drain_left.t8 plus.t6 source.t13 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X13 drain_left.t6 plus.t7 source.t12 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X14 a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X15 drain_left.t7 plus.t8 source.t11 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X16 drain_right.t4 minus.t5 source.t6 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X17 drain_right.t3 minus.t6 source.t8 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X18 source.t7 minus.t7 drain_right.t2 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X19 drain_right.t1 minus.t8 source.t1 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X20 a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X21 source.t10 plus.t9 drain_left.t1 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X22 a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X23 drain_right.t0 minus.t9 source.t4 a_n1412_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
R0 plus.n2 plus.t4 2113.2
R1 plus.n8 plus.t6 2113.2
R2 plus.n12 plus.t2 2113.2
R3 plus.n18 plus.t5 2113.2
R4 plus.n1 plus.t1 2053.32
R5 plus.n5 plus.t7 2053.32
R6 plus.n7 plus.t0 2053.32
R7 plus.n11 plus.t9 2053.32
R8 plus.n15 plus.t8 2053.32
R9 plus.n17 plus.t3 2053.32
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 31.3968
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 15.1899
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n5 drain_left.t5 61.3084
R37 drain_left.n1 drain_left.t4 61.3083
R38 drain_left.n3 drain_left.n2 60.1381
R39 drain_left.n7 drain_left.n6 59.8185
R40 drain_left.n5 drain_left.n4 59.8185
R41 drain_left.n1 drain_left.n0 59.8184
R42 drain_left drain_left.n3 35.5527
R43 drain_left drain_left.n7 6.15322
R44 drain_left.n2 drain_left.t1 0.9905
R45 drain_left.n2 drain_left.t2 0.9905
R46 drain_left.n0 drain_left.t3 0.9905
R47 drain_left.n0 drain_left.t7 0.9905
R48 drain_left.n6 drain_left.t9 0.9905
R49 drain_left.n6 drain_left.t8 0.9905
R50 drain_left.n4 drain_left.t0 0.9905
R51 drain_left.n4 drain_left.t6 0.9905
R52 drain_left.n7 drain_left.n5 0.5005
R53 drain_left.n3 drain_left.n1 0.070154
R54 source.n0 source.t13 44.1297
R55 source.n5 source.t8 44.1296
R56 source.n19 source.t2 44.1295
R57 source.n14 source.t17 44.1295
R58 source.n2 source.n1 43.1397
R59 source.n4 source.n3 43.1397
R60 source.n7 source.n6 43.1397
R61 source.n9 source.n8 43.1397
R62 source.n18 source.n17 43.1396
R63 source.n16 source.n15 43.1396
R64 source.n13 source.n12 43.1396
R65 source.n11 source.n10 43.1396
R66 source.n11 source.n9 28.3483
R67 source.n20 source.n0 22.3354
R68 source.n20 source.n19 5.51343
R69 source.n17 source.t4 0.9905
R70 source.n17 source.t7 0.9905
R71 source.n15 source.t5 0.9905
R72 source.n15 source.t9 0.9905
R73 source.n12 source.t11 0.9905
R74 source.n12 source.t10 0.9905
R75 source.n10 source.t14 0.9905
R76 source.n10 source.t16 0.9905
R77 source.n1 source.t12 0.9905
R78 source.n1 source.t19 0.9905
R79 source.n3 source.t15 0.9905
R80 source.n3 source.t18 0.9905
R81 source.n6 source.t6 0.9905
R82 source.n6 source.t3 0.9905
R83 source.n8 source.t1 0.9905
R84 source.n8 source.t0 0.9905
R85 source.n5 source.n4 0.720328
R86 source.n16 source.n14 0.720328
R87 source.n9 source.n7 0.5005
R88 source.n7 source.n5 0.5005
R89 source.n4 source.n2 0.5005
R90 source.n2 source.n0 0.5005
R91 source.n13 source.n11 0.5005
R92 source.n14 source.n13 0.5005
R93 source.n18 source.n16 0.5005
R94 source.n19 source.n18 0.5005
R95 source source.n20 0.188
R96 minus.n8 minus.t8 2113.2
R97 minus.n2 minus.t6 2113.2
R98 minus.n18 minus.t4 2113.2
R99 minus.n12 minus.t1 2113.2
R100 minus.n7 minus.t0 2053.32
R101 minus.n5 minus.t5 2053.32
R102 minus.n1 minus.t2 2053.32
R103 minus.n17 minus.t7 2053.32
R104 minus.n15 minus.t9 2053.32
R105 minus.n11 minus.t3 2053.32
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 48.2005
R115 minus.n4 minus.n1 48.2005
R116 minus.n14 minus.n11 48.2005
R117 minus.n17 minus.n16 48.2005
R118 minus.n20 minus.n9 40.546
R119 minus.n6 minus.n5 36.5157
R120 minus.n5 minus.n4 36.5157
R121 minus.n15 minus.n14 36.5157
R122 minus.n16 minus.n15 36.5157
R123 minus.n8 minus.n7 24.8308
R124 minus.n2 minus.n1 24.8308
R125 minus.n12 minus.n11 24.8308
R126 minus.n18 minus.n17 24.8308
R127 minus.n20 minus.n19 6.51565
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t8 61.3083
R134 drain_right.n7 drain_right.t1 60.8084
R135 drain_right.n6 drain_right.n4 60.3185
R136 drain_right.n3 drain_right.n2 60.1381
R137 drain_right.n6 drain_right.n5 59.8185
R138 drain_right.n1 drain_right.n0 59.8184
R139 drain_right drain_right.n3 34.9995
R140 drain_right drain_right.n7 5.90322
R141 drain_right.n2 drain_right.t2 0.9905
R142 drain_right.n2 drain_right.t5 0.9905
R143 drain_right.n0 drain_right.t6 0.9905
R144 drain_right.n0 drain_right.t0 0.9905
R145 drain_right.n4 drain_right.t7 0.9905
R146 drain_right.n4 drain_right.t3 0.9905
R147 drain_right.n5 drain_right.t9 0.9905
R148 drain_right.n5 drain_right.t4 0.9905
R149 drain_right.n7 drain_right.n6 0.5005
R150 drain_right.n3 drain_right.n1 0.070154
C0 drain_right minus 5.66008f
C1 drain_left source 36.5348f
C2 drain_right source 36.5164f
C3 drain_left plus 5.789431f
C4 drain_right plus 0.291664f
C5 drain_left drain_right 0.697299f
C6 minus source 4.8797f
C7 plus minus 6.39154f
C8 plus source 4.89486f
C9 drain_left minus 0.171039f
C10 drain_right a_n1412_n4888# 9.4025f
C11 drain_left a_n1412_n4888# 9.637111f
C12 source a_n1412_n4888# 8.800015f
C13 minus a_n1412_n4888# 5.979995f
C14 plus a_n1412_n4888# 8.607651f
C15 drain_right.t8 a_n1412_n4888# 5.82712f
C16 drain_right.t6 a_n1412_n4888# 0.498073f
C17 drain_right.t0 a_n1412_n4888# 0.498073f
C18 drain_right.n0 a_n1412_n4888# 4.55349f
C19 drain_right.n1 a_n1412_n4888# 0.74843f
C20 drain_right.t2 a_n1412_n4888# 0.498073f
C21 drain_right.t5 a_n1412_n4888# 0.498073f
C22 drain_right.n2 a_n1412_n4888# 4.55543f
C23 drain_right.n3 a_n1412_n4888# 2.30758f
C24 drain_right.t7 a_n1412_n4888# 0.498073f
C25 drain_right.t3 a_n1412_n4888# 0.498073f
C26 drain_right.n4 a_n1412_n4888# 4.55664f
C27 drain_right.t9 a_n1412_n4888# 0.498073f
C28 drain_right.t4 a_n1412_n4888# 0.498073f
C29 drain_right.n5 a_n1412_n4888# 4.55349f
C30 drain_right.n6 a_n1412_n4888# 0.744521f
C31 drain_right.t1 a_n1412_n4888# 5.82374f
C32 drain_right.n7 a_n1412_n4888# 0.677071f
C33 minus.n0 a_n1412_n4888# 0.056017f
C34 minus.t8 a_n1412_n4888# 0.797394f
C35 minus.t0 a_n1412_n4888# 0.788852f
C36 minus.t5 a_n1412_n4888# 0.788852f
C37 minus.t2 a_n1412_n4888# 0.788852f
C38 minus.n1 a_n1412_n4888# 0.295918f
C39 minus.t6 a_n1412_n4888# 0.797394f
C40 minus.n2 a_n1412_n4888# 0.314335f
C41 minus.n3 a_n1412_n4888# 0.131631f
C42 minus.n4 a_n1412_n4888# 0.021346f
C43 minus.n5 a_n1412_n4888# 0.295918f
C44 minus.n6 a_n1412_n4888# 0.021346f
C45 minus.n7 a_n1412_n4888# 0.295918f
C46 minus.n8 a_n1412_n4888# 0.314247f
C47 minus.n9 a_n1412_n4888# 2.35514f
C48 minus.n10 a_n1412_n4888# 0.056017f
C49 minus.t7 a_n1412_n4888# 0.788852f
C50 minus.t9 a_n1412_n4888# 0.788852f
C51 minus.t3 a_n1412_n4888# 0.788852f
C52 minus.n11 a_n1412_n4888# 0.295918f
C53 minus.t1 a_n1412_n4888# 0.797394f
C54 minus.n12 a_n1412_n4888# 0.314335f
C55 minus.n13 a_n1412_n4888# 0.131631f
C56 minus.n14 a_n1412_n4888# 0.021346f
C57 minus.n15 a_n1412_n4888# 0.295918f
C58 minus.n16 a_n1412_n4888# 0.021346f
C59 minus.n17 a_n1412_n4888# 0.295918f
C60 minus.t4 a_n1412_n4888# 0.797394f
C61 minus.n18 a_n1412_n4888# 0.314247f
C62 minus.n19 a_n1412_n4888# 0.368288f
C63 minus.n20 a_n1412_n4888# 2.82375f
C64 source.t13 a_n1412_n4888# 5.75384f
C65 source.n0 a_n1412_n4888# 2.44033f
C66 source.t12 a_n1412_n4888# 0.50347f
C67 source.t19 a_n1412_n4888# 0.50347f
C68 source.n1 a_n1412_n4888# 4.50123f
C69 source.n2 a_n1412_n4888# 0.429763f
C70 source.t15 a_n1412_n4888# 0.50347f
C71 source.t18 a_n1412_n4888# 0.50347f
C72 source.n3 a_n1412_n4888# 4.50123f
C73 source.n4 a_n1412_n4888# 0.452327f
C74 source.t8 a_n1412_n4888# 5.75386f
C75 source.n5 a_n1412_n4888# 0.572806f
C76 source.t6 a_n1412_n4888# 0.50347f
C77 source.t3 a_n1412_n4888# 0.50347f
C78 source.n6 a_n1412_n4888# 4.50123f
C79 source.n7 a_n1412_n4888# 0.429763f
C80 source.t1 a_n1412_n4888# 0.50347f
C81 source.t0 a_n1412_n4888# 0.50347f
C82 source.n8 a_n1412_n4888# 4.50123f
C83 source.n9 a_n1412_n4888# 2.93382f
C84 source.t14 a_n1412_n4888# 0.50347f
C85 source.t16 a_n1412_n4888# 0.50347f
C86 source.n10 a_n1412_n4888# 4.50124f
C87 source.n11 a_n1412_n4888# 2.93381f
C88 source.t11 a_n1412_n4888# 0.50347f
C89 source.t10 a_n1412_n4888# 0.50347f
C90 source.n12 a_n1412_n4888# 4.50124f
C91 source.n13 a_n1412_n4888# 0.429754f
C92 source.t17 a_n1412_n4888# 5.75382f
C93 source.n14 a_n1412_n4888# 0.572838f
C94 source.t5 a_n1412_n4888# 0.50347f
C95 source.t9 a_n1412_n4888# 0.50347f
C96 source.n15 a_n1412_n4888# 4.50124f
C97 source.n16 a_n1412_n4888# 0.452319f
C98 source.t4 a_n1412_n4888# 0.50347f
C99 source.t7 a_n1412_n4888# 0.50347f
C100 source.n17 a_n1412_n4888# 4.50124f
C101 source.n18 a_n1412_n4888# 0.429754f
C102 source.t2 a_n1412_n4888# 5.75382f
C103 source.n19 a_n1412_n4888# 0.72346f
C104 source.n20 a_n1412_n4888# 2.86487f
C105 drain_left.t4 a_n1412_n4888# 5.82391f
C106 drain_left.t3 a_n1412_n4888# 0.497799f
C107 drain_left.t7 a_n1412_n4888# 0.497799f
C108 drain_left.n0 a_n1412_n4888# 4.55099f
C109 drain_left.n1 a_n1412_n4888# 0.748019f
C110 drain_left.t1 a_n1412_n4888# 0.497799f
C111 drain_left.t2 a_n1412_n4888# 0.497799f
C112 drain_left.n2 a_n1412_n4888# 4.55292f
C113 drain_left.n3 a_n1412_n4888# 2.37231f
C114 drain_left.t5 a_n1412_n4888# 5.82394f
C115 drain_left.t0 a_n1412_n4888# 0.497799f
C116 drain_left.t6 a_n1412_n4888# 0.497799f
C117 drain_left.n4 a_n1412_n4888# 4.55098f
C118 drain_left.n5 a_n1412_n4888# 0.781195f
C119 drain_left.t9 a_n1412_n4888# 0.497799f
C120 drain_left.t8 a_n1412_n4888# 0.497799f
C121 drain_left.n6 a_n1412_n4888# 4.55098f
C122 drain_left.n7 a_n1412_n4888# 0.627274f
C123 plus.n0 a_n1412_n4888# 0.056724f
C124 plus.t0 a_n1412_n4888# 0.798815f
C125 plus.t7 a_n1412_n4888# 0.798815f
C126 plus.t1 a_n1412_n4888# 0.798815f
C127 plus.n1 a_n1412_n4888# 0.299655f
C128 plus.t4 a_n1412_n4888# 0.807466f
C129 plus.n2 a_n1412_n4888# 0.318306f
C130 plus.n3 a_n1412_n4888# 0.133293f
C131 plus.n4 a_n1412_n4888# 0.021615f
C132 plus.n5 a_n1412_n4888# 0.299655f
C133 plus.n6 a_n1412_n4888# 0.021615f
C134 plus.n7 a_n1412_n4888# 0.299655f
C135 plus.t6 a_n1412_n4888# 0.807466f
C136 plus.n8 a_n1412_n4888# 0.318216f
C137 plus.n9 a_n1412_n4888# 0.863363f
C138 plus.n10 a_n1412_n4888# 0.056724f
C139 plus.t5 a_n1412_n4888# 0.807466f
C140 plus.t3 a_n1412_n4888# 0.798815f
C141 plus.t8 a_n1412_n4888# 0.798815f
C142 plus.t9 a_n1412_n4888# 0.798815f
C143 plus.n11 a_n1412_n4888# 0.299655f
C144 plus.t2 a_n1412_n4888# 0.807466f
C145 plus.n12 a_n1412_n4888# 0.318306f
C146 plus.n13 a_n1412_n4888# 0.133293f
C147 plus.n14 a_n1412_n4888# 0.021615f
C148 plus.n15 a_n1412_n4888# 0.299655f
C149 plus.n16 a_n1412_n4888# 0.021615f
C150 plus.n17 a_n1412_n4888# 0.299655f
C151 plus.n18 a_n1412_n4888# 0.318216f
C152 plus.n19 a_n1412_n4888# 1.87518f
.ends

