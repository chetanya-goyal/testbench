* NGSPICE file created from diffpair348.ext - technology: sky130A

.subckt diffpair348 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t34 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 drain_left.t18 plus.t1 source.t27 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 drain_right.t19 minus.t0 source.t7 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X3 drain_right.t18 minus.t1 source.t1 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 drain_left.t17 plus.t2 source.t24 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 drain_left.t16 plus.t3 source.t20 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X6 source.t3 minus.t2 drain_right.t17 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 source.t8 minus.t3 drain_right.t16 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 drain_left.t15 plus.t4 source.t28 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X9 source.t2 minus.t4 drain_right.t15 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X10 source.t36 plus.t5 drain_left.t14 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X11 a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X12 drain_left.t13 plus.t6 source.t32 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X13 source.t30 plus.t7 drain_left.t12 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X14 source.t6 minus.t5 drain_right.t14 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X15 a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X16 source.t10 minus.t6 drain_right.t13 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 source.t12 minus.t7 drain_right.t12 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X18 source.t16 minus.t8 drain_right.t11 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X19 source.t22 plus.t8 drain_left.t11 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X20 source.t29 plus.t9 drain_left.t10 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X21 source.t23 plus.t10 drain_left.t9 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X22 source.t19 plus.t11 drain_left.t8 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X23 drain_right.t10 minus.t9 source.t17 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X24 drain_left.t7 plus.t12 source.t18 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X25 drain_right.t9 minus.t10 source.t38 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X26 source.t31 plus.t13 drain_left.t6 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X27 drain_left.t5 plus.t14 source.t25 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X28 drain_right.t8 minus.t11 source.t39 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X29 source.t5 minus.t12 drain_right.t7 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X30 source.t0 minus.t13 drain_right.t6 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X31 source.t37 plus.t15 drain_left.t4 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X32 drain_right.t5 minus.t14 source.t4 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X33 a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X34 source.t35 plus.t16 drain_left.t3 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X35 drain_left.t2 plus.t17 source.t33 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X36 drain_right.t4 minus.t15 source.t15 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X37 source.t13 minus.t16 drain_right.t3 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X38 a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X39 source.t26 plus.t18 drain_left.t1 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X40 drain_right.t2 minus.t17 source.t9 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X41 drain_right.t1 minus.t18 source.t11 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X42 drain_right.t0 minus.t19 source.t14 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X43 drain_left.t0 plus.t19 source.t21 a_n1992_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
R0 plus.n6 plus.t7 1045.5
R1 plus.n25 plus.t3 1045.5
R2 plus.n33 plus.t17 1045.5
R3 plus.n52 plus.t8 1045.5
R4 plus.n5 plus.t1 992.92
R5 plus.n9 plus.t11 992.92
R6 plus.n11 plus.t0 992.92
R7 plus.n3 plus.t10 992.92
R8 plus.n17 plus.t19 992.92
R9 plus.n1 plus.t9 992.92
R10 plus.n22 plus.t4 992.92
R11 plus.n24 plus.t15 992.92
R12 plus.n32 plus.t13 992.92
R13 plus.n36 plus.t6 992.92
R14 plus.n38 plus.t18 992.92
R15 plus.n30 plus.t2 992.92
R16 plus.n44 plus.t16 992.92
R17 plus.n28 plus.t12 992.92
R18 plus.n49 plus.t5 992.92
R19 plus.n51 plus.t14 992.92
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus plus.n53 29.4081
R63 plus.n10 plus.n9 29.2126
R64 plus.n22 plus.n21 29.2126
R65 plus.n49 plus.n48 29.2126
R66 plus.n37 plus.n36 29.2126
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 11.0043
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n9 source.t30 51.0588
R93 source.n10 source.t4 51.0588
R94 source.n19 source.t12 51.0588
R95 source.n39 source.t7 51.0586
R96 source.n30 source.t13 51.0586
R97 source.n29 source.t33 51.0586
R98 source.n20 source.t22 51.0586
R99 source.n0 source.t20 51.0586
R100 source.n2 source.n1 48.8588
R101 source.n4 source.n3 48.8588
R102 source.n6 source.n5 48.8588
R103 source.n8 source.n7 48.8588
R104 source.n12 source.n11 48.8588
R105 source.n14 source.n13 48.8588
R106 source.n16 source.n15 48.8588
R107 source.n18 source.n17 48.8588
R108 source.n38 source.n37 48.8586
R109 source.n36 source.n35 48.8586
R110 source.n34 source.n33 48.8586
R111 source.n32 source.n31 48.8586
R112 source.n28 source.n27 48.8586
R113 source.n26 source.n25 48.8586
R114 source.n24 source.n23 48.8586
R115 source.n22 source.n21 48.8586
R116 source.n20 source.n19 19.515
R117 source.n40 source.n0 14.0021
R118 source.n40 source.n39 5.51343
R119 source.n37 source.t38 2.2005
R120 source.n37 source.t16 2.2005
R121 source.n35 source.t15 2.2005
R122 source.n35 source.t5 2.2005
R123 source.n33 source.t17 2.2005
R124 source.n33 source.t8 2.2005
R125 source.n31 source.t1 2.2005
R126 source.n31 source.t0 2.2005
R127 source.n27 source.t32 2.2005
R128 source.n27 source.t31 2.2005
R129 source.n25 source.t24 2.2005
R130 source.n25 source.t26 2.2005
R131 source.n23 source.t18 2.2005
R132 source.n23 source.t35 2.2005
R133 source.n21 source.t25 2.2005
R134 source.n21 source.t36 2.2005
R135 source.n1 source.t28 2.2005
R136 source.n1 source.t37 2.2005
R137 source.n3 source.t21 2.2005
R138 source.n3 source.t29 2.2005
R139 source.n5 source.t34 2.2005
R140 source.n5 source.t23 2.2005
R141 source.n7 source.t27 2.2005
R142 source.n7 source.t19 2.2005
R143 source.n11 source.t39 2.2005
R144 source.n11 source.t2 2.2005
R145 source.n13 source.t9 2.2005
R146 source.n13 source.t3 2.2005
R147 source.n15 source.t11 2.2005
R148 source.n15 source.t10 2.2005
R149 source.n17 source.t14 2.2005
R150 source.n17 source.t6 2.2005
R151 source.n19 source.n18 0.5005
R152 source.n18 source.n16 0.5005
R153 source.n16 source.n14 0.5005
R154 source.n14 source.n12 0.5005
R155 source.n12 source.n10 0.5005
R156 source.n9 source.n8 0.5005
R157 source.n8 source.n6 0.5005
R158 source.n6 source.n4 0.5005
R159 source.n4 source.n2 0.5005
R160 source.n2 source.n0 0.5005
R161 source.n22 source.n20 0.5005
R162 source.n24 source.n22 0.5005
R163 source.n26 source.n24 0.5005
R164 source.n28 source.n26 0.5005
R165 source.n29 source.n28 0.5005
R166 source.n32 source.n30 0.5005
R167 source.n34 source.n32 0.5005
R168 source.n36 source.n34 0.5005
R169 source.n38 source.n36 0.5005
R170 source.n39 source.n38 0.5005
R171 source.n10 source.n9 0.470328
R172 source.n30 source.n29 0.470328
R173 source source.n40 0.188
R174 drain_left.n10 drain_left.n8 66.0376
R175 drain_left.n6 drain_left.n4 66.0373
R176 drain_left.n2 drain_left.n0 66.0373
R177 drain_left.n14 drain_left.n13 65.5376
R178 drain_left.n12 drain_left.n11 65.5376
R179 drain_left.n10 drain_left.n9 65.5376
R180 drain_left.n16 drain_left.n15 65.5374
R181 drain_left.n7 drain_left.n3 65.5373
R182 drain_left.n6 drain_left.n5 65.5373
R183 drain_left.n2 drain_left.n1 65.5373
R184 drain_left drain_left.n7 29.0943
R185 drain_left drain_left.n16 6.15322
R186 drain_left.n3 drain_left.t3 2.2005
R187 drain_left.n3 drain_left.t17 2.2005
R188 drain_left.n4 drain_left.t6 2.2005
R189 drain_left.n4 drain_left.t2 2.2005
R190 drain_left.n5 drain_left.t1 2.2005
R191 drain_left.n5 drain_left.t13 2.2005
R192 drain_left.n1 drain_left.t14 2.2005
R193 drain_left.n1 drain_left.t7 2.2005
R194 drain_left.n0 drain_left.t11 2.2005
R195 drain_left.n0 drain_left.t5 2.2005
R196 drain_left.n15 drain_left.t4 2.2005
R197 drain_left.n15 drain_left.t16 2.2005
R198 drain_left.n13 drain_left.t10 2.2005
R199 drain_left.n13 drain_left.t15 2.2005
R200 drain_left.n11 drain_left.t9 2.2005
R201 drain_left.n11 drain_left.t0 2.2005
R202 drain_left.n9 drain_left.t8 2.2005
R203 drain_left.n9 drain_left.t19 2.2005
R204 drain_left.n8 drain_left.t12 2.2005
R205 drain_left.n8 drain_left.t18 2.2005
R206 drain_left.n12 drain_left.n10 0.5005
R207 drain_left.n14 drain_left.n12 0.5005
R208 drain_left.n16 drain_left.n14 0.5005
R209 drain_left.n7 drain_left.n6 0.445154
R210 drain_left.n7 drain_left.n2 0.445154
R211 minus.n25 minus.t7 1045.5
R212 minus.n6 minus.t14 1045.5
R213 minus.n52 minus.t0 1045.5
R214 minus.n33 minus.t16 1045.5
R215 minus.n24 minus.t19 992.92
R216 minus.n22 minus.t5 992.92
R217 minus.n1 minus.t18 992.92
R218 minus.n17 minus.t6 992.92
R219 minus.n3 minus.t17 992.92
R220 minus.n11 minus.t2 992.92
R221 minus.n9 minus.t11 992.92
R222 minus.n5 minus.t4 992.92
R223 minus.n51 minus.t8 992.92
R224 minus.n49 minus.t10 992.92
R225 minus.n28 minus.t12 992.92
R226 minus.n44 minus.t15 992.92
R227 minus.n30 minus.t3 992.92
R228 minus.n38 minus.t9 992.92
R229 minus.n36 minus.t13 992.92
R230 minus.n32 minus.t1 992.92
R231 minus.n7 minus.n6 161.489
R232 minus.n34 minus.n33 161.489
R233 minus.n26 minus.n25 161.3
R234 minus.n23 minus.n0 161.3
R235 minus.n21 minus.n20 161.3
R236 minus.n19 minus.n18 161.3
R237 minus.n16 minus.n2 161.3
R238 minus.n15 minus.n14 161.3
R239 minus.n13 minus.n12 161.3
R240 minus.n10 minus.n4 161.3
R241 minus.n8 minus.n7 161.3
R242 minus.n53 minus.n52 161.3
R243 minus.n50 minus.n27 161.3
R244 minus.n48 minus.n47 161.3
R245 minus.n46 minus.n45 161.3
R246 minus.n43 minus.n29 161.3
R247 minus.n42 minus.n41 161.3
R248 minus.n40 minus.n39 161.3
R249 minus.n37 minus.n31 161.3
R250 minus.n35 minus.n34 161.3
R251 minus.n16 minus.n15 73.0308
R252 minus.n43 minus.n42 73.0308
R253 minus.n18 minus.n17 67.1884
R254 minus.n12 minus.n3 67.1884
R255 minus.n39 minus.n30 67.1884
R256 minus.n45 minus.n44 67.1884
R257 minus.n21 minus.n1 55.5035
R258 minus.n11 minus.n10 55.5035
R259 minus.n38 minus.n37 55.5035
R260 minus.n48 minus.n28 55.5035
R261 minus.n23 minus.n22 43.8187
R262 minus.n9 minus.n8 43.8187
R263 minus.n36 minus.n35 43.8187
R264 minus.n50 minus.n49 43.8187
R265 minus.n24 minus.n23 40.8975
R266 minus.n8 minus.n5 40.8975
R267 minus.n35 minus.n32 40.8975
R268 minus.n51 minus.n50 40.8975
R269 minus.n54 minus.n26 34.3907
R270 minus.n25 minus.n24 32.1338
R271 minus.n6 minus.n5 32.1338
R272 minus.n33 minus.n32 32.1338
R273 minus.n52 minus.n51 32.1338
R274 minus.n22 minus.n21 29.2126
R275 minus.n10 minus.n9 29.2126
R276 minus.n37 minus.n36 29.2126
R277 minus.n49 minus.n48 29.2126
R278 minus.n18 minus.n1 17.5278
R279 minus.n12 minus.n11 17.5278
R280 minus.n39 minus.n38 17.5278
R281 minus.n45 minus.n28 17.5278
R282 minus.n54 minus.n53 6.49671
R283 minus.n17 minus.n16 5.84292
R284 minus.n15 minus.n3 5.84292
R285 minus.n42 minus.n30 5.84292
R286 minus.n44 minus.n43 5.84292
R287 minus.n26 minus.n0 0.189894
R288 minus.n20 minus.n0 0.189894
R289 minus.n20 minus.n19 0.189894
R290 minus.n19 minus.n2 0.189894
R291 minus.n14 minus.n2 0.189894
R292 minus.n14 minus.n13 0.189894
R293 minus.n13 minus.n4 0.189894
R294 minus.n7 minus.n4 0.189894
R295 minus.n34 minus.n31 0.189894
R296 minus.n40 minus.n31 0.189894
R297 minus.n41 minus.n40 0.189894
R298 minus.n41 minus.n29 0.189894
R299 minus.n46 minus.n29 0.189894
R300 minus.n47 minus.n46 0.189894
R301 minus.n47 minus.n27 0.189894
R302 minus.n53 minus.n27 0.189894
R303 minus minus.n54 0.188
R304 drain_right.n10 drain_right.n8 66.0374
R305 drain_right.n6 drain_right.n4 66.0373
R306 drain_right.n2 drain_right.n0 66.0373
R307 drain_right.n10 drain_right.n9 65.5376
R308 drain_right.n12 drain_right.n11 65.5376
R309 drain_right.n14 drain_right.n13 65.5376
R310 drain_right.n16 drain_right.n15 65.5376
R311 drain_right.n7 drain_right.n3 65.5373
R312 drain_right.n6 drain_right.n5 65.5373
R313 drain_right.n2 drain_right.n1 65.5373
R314 drain_right drain_right.n7 28.5411
R315 drain_right drain_right.n16 6.15322
R316 drain_right.n3 drain_right.t16 2.2005
R317 drain_right.n3 drain_right.t4 2.2005
R318 drain_right.n4 drain_right.t11 2.2005
R319 drain_right.n4 drain_right.t19 2.2005
R320 drain_right.n5 drain_right.t7 2.2005
R321 drain_right.n5 drain_right.t9 2.2005
R322 drain_right.n1 drain_right.t6 2.2005
R323 drain_right.n1 drain_right.t10 2.2005
R324 drain_right.n0 drain_right.t3 2.2005
R325 drain_right.n0 drain_right.t18 2.2005
R326 drain_right.n8 drain_right.t15 2.2005
R327 drain_right.n8 drain_right.t5 2.2005
R328 drain_right.n9 drain_right.t17 2.2005
R329 drain_right.n9 drain_right.t8 2.2005
R330 drain_right.n11 drain_right.t13 2.2005
R331 drain_right.n11 drain_right.t2 2.2005
R332 drain_right.n13 drain_right.t14 2.2005
R333 drain_right.n13 drain_right.t1 2.2005
R334 drain_right.n15 drain_right.t12 2.2005
R335 drain_right.n15 drain_right.t0 2.2005
R336 drain_right.n16 drain_right.n14 0.5005
R337 drain_right.n14 drain_right.n12 0.5005
R338 drain_right.n12 drain_right.n10 0.5005
R339 drain_right.n7 drain_right.n6 0.445154
R340 drain_right.n7 drain_right.n2 0.445154
C0 source minus 4.67468f
C1 drain_right minus 4.84776f
C2 minus plus 5.0825f
C3 drain_left minus 0.171712f
C4 drain_right source 31.477198f
C5 source plus 4.68872f
C6 source drain_left 31.477001f
C7 drain_right plus 0.349242f
C8 drain_right drain_left 1.04652f
C9 drain_left plus 5.04226f
C10 drain_right a_n1992_n2688# 6.31462f
C11 drain_left a_n1992_n2688# 6.62519f
C12 source a_n1992_n2688# 7.11378f
C13 minus a_n1992_n2688# 7.57436f
C14 plus a_n1992_n2688# 9.42146f
C15 drain_right.t3 a_n1992_n2688# 0.255126f
C16 drain_right.t18 a_n1992_n2688# 0.255126f
C17 drain_right.n0 a_n1992_n2688# 2.23466f
C18 drain_right.t6 a_n1992_n2688# 0.255126f
C19 drain_right.t10 a_n1992_n2688# 0.255126f
C20 drain_right.n1 a_n1992_n2688# 2.2315f
C21 drain_right.n2 a_n1992_n2688# 0.812619f
C22 drain_right.t16 a_n1992_n2688# 0.255126f
C23 drain_right.t4 a_n1992_n2688# 0.255126f
C24 drain_right.n3 a_n1992_n2688# 2.2315f
C25 drain_right.t11 a_n1992_n2688# 0.255126f
C26 drain_right.t19 a_n1992_n2688# 0.255126f
C27 drain_right.n4 a_n1992_n2688# 2.23466f
C28 drain_right.t7 a_n1992_n2688# 0.255126f
C29 drain_right.t9 a_n1992_n2688# 0.255126f
C30 drain_right.n5 a_n1992_n2688# 2.2315f
C31 drain_right.n6 a_n1992_n2688# 0.812619f
C32 drain_right.n7 a_n1992_n2688# 1.84032f
C33 drain_right.t15 a_n1992_n2688# 0.255126f
C34 drain_right.t5 a_n1992_n2688# 0.255126f
C35 drain_right.n8 a_n1992_n2688# 2.23466f
C36 drain_right.t17 a_n1992_n2688# 0.255126f
C37 drain_right.t8 a_n1992_n2688# 0.255126f
C38 drain_right.n9 a_n1992_n2688# 2.2315f
C39 drain_right.n10 a_n1992_n2688# 0.817147f
C40 drain_right.t13 a_n1992_n2688# 0.255126f
C41 drain_right.t2 a_n1992_n2688# 0.255126f
C42 drain_right.n11 a_n1992_n2688# 2.2315f
C43 drain_right.n12 a_n1992_n2688# 0.402925f
C44 drain_right.t14 a_n1992_n2688# 0.255126f
C45 drain_right.t1 a_n1992_n2688# 0.255126f
C46 drain_right.n13 a_n1992_n2688# 2.2315f
C47 drain_right.n14 a_n1992_n2688# 0.402925f
C48 drain_right.t12 a_n1992_n2688# 0.255126f
C49 drain_right.t0 a_n1992_n2688# 0.255126f
C50 drain_right.n15 a_n1992_n2688# 2.2315f
C51 drain_right.n16 a_n1992_n2688# 0.699025f
C52 minus.n0 a_n1992_n2688# 0.050739f
C53 minus.t7 a_n1992_n2688# 0.330593f
C54 minus.t19 a_n1992_n2688# 0.323495f
C55 minus.t5 a_n1992_n2688# 0.323495f
C56 minus.t18 a_n1992_n2688# 0.323495f
C57 minus.n1 a_n1992_n2688# 0.137693f
C58 minus.n2 a_n1992_n2688# 0.050739f
C59 minus.t6 a_n1992_n2688# 0.323495f
C60 minus.t17 a_n1992_n2688# 0.323495f
C61 minus.n3 a_n1992_n2688# 0.137693f
C62 minus.n4 a_n1992_n2688# 0.050739f
C63 minus.t2 a_n1992_n2688# 0.323495f
C64 minus.t11 a_n1992_n2688# 0.323495f
C65 minus.t4 a_n1992_n2688# 0.323495f
C66 minus.n5 a_n1992_n2688# 0.137693f
C67 minus.t14 a_n1992_n2688# 0.330593f
C68 minus.n6 a_n1992_n2688# 0.153447f
C69 minus.n7 a_n1992_n2688# 0.116105f
C70 minus.n8 a_n1992_n2688# 0.019335f
C71 minus.n9 a_n1992_n2688# 0.137693f
C72 minus.n10 a_n1992_n2688# 0.019335f
C73 minus.n11 a_n1992_n2688# 0.137693f
C74 minus.n12 a_n1992_n2688# 0.019335f
C75 minus.n13 a_n1992_n2688# 0.050739f
C76 minus.n14 a_n1992_n2688# 0.050739f
C77 minus.n15 a_n1992_n2688# 0.018083f
C78 minus.n16 a_n1992_n2688# 0.018083f
C79 minus.n17 a_n1992_n2688# 0.137693f
C80 minus.n18 a_n1992_n2688# 0.019335f
C81 minus.n19 a_n1992_n2688# 0.050739f
C82 minus.n20 a_n1992_n2688# 0.050739f
C83 minus.n21 a_n1992_n2688# 0.019335f
C84 minus.n22 a_n1992_n2688# 0.137693f
C85 minus.n23 a_n1992_n2688# 0.019335f
C86 minus.n24 a_n1992_n2688# 0.137693f
C87 minus.n25 a_n1992_n2688# 0.153371f
C88 minus.n26 a_n1992_n2688# 1.65386f
C89 minus.n27 a_n1992_n2688# 0.050739f
C90 minus.t8 a_n1992_n2688# 0.323495f
C91 minus.t10 a_n1992_n2688# 0.323495f
C92 minus.t12 a_n1992_n2688# 0.323495f
C93 minus.n28 a_n1992_n2688# 0.137693f
C94 minus.n29 a_n1992_n2688# 0.050739f
C95 minus.t15 a_n1992_n2688# 0.323495f
C96 minus.t3 a_n1992_n2688# 0.323495f
C97 minus.n30 a_n1992_n2688# 0.137693f
C98 minus.n31 a_n1992_n2688# 0.050739f
C99 minus.t9 a_n1992_n2688# 0.323495f
C100 minus.t13 a_n1992_n2688# 0.323495f
C101 minus.t1 a_n1992_n2688# 0.323495f
C102 minus.n32 a_n1992_n2688# 0.137693f
C103 minus.t16 a_n1992_n2688# 0.330593f
C104 minus.n33 a_n1992_n2688# 0.153447f
C105 minus.n34 a_n1992_n2688# 0.116105f
C106 minus.n35 a_n1992_n2688# 0.019335f
C107 minus.n36 a_n1992_n2688# 0.137693f
C108 minus.n37 a_n1992_n2688# 0.019335f
C109 minus.n38 a_n1992_n2688# 0.137693f
C110 minus.n39 a_n1992_n2688# 0.019335f
C111 minus.n40 a_n1992_n2688# 0.050739f
C112 minus.n41 a_n1992_n2688# 0.050739f
C113 minus.n42 a_n1992_n2688# 0.018083f
C114 minus.n43 a_n1992_n2688# 0.018083f
C115 minus.n44 a_n1992_n2688# 0.137693f
C116 minus.n45 a_n1992_n2688# 0.019335f
C117 minus.n46 a_n1992_n2688# 0.050739f
C118 minus.n47 a_n1992_n2688# 0.050739f
C119 minus.n48 a_n1992_n2688# 0.019335f
C120 minus.n49 a_n1992_n2688# 0.137693f
C121 minus.n50 a_n1992_n2688# 0.019335f
C122 minus.n51 a_n1992_n2688# 0.137693f
C123 minus.t0 a_n1992_n2688# 0.330593f
C124 minus.n52 a_n1992_n2688# 0.153371f
C125 minus.n53 a_n1992_n2688# 0.331329f
C126 minus.n54 a_n1992_n2688# 2.01956f
C127 drain_left.t11 a_n1992_n2688# 0.255544f
C128 drain_left.t5 a_n1992_n2688# 0.255544f
C129 drain_left.n0 a_n1992_n2688# 2.23832f
C130 drain_left.t14 a_n1992_n2688# 0.255544f
C131 drain_left.t7 a_n1992_n2688# 0.255544f
C132 drain_left.n1 a_n1992_n2688# 2.23515f
C133 drain_left.n2 a_n1992_n2688# 0.81395f
C134 drain_left.t3 a_n1992_n2688# 0.255544f
C135 drain_left.t17 a_n1992_n2688# 0.255544f
C136 drain_left.n3 a_n1992_n2688# 2.23515f
C137 drain_left.t6 a_n1992_n2688# 0.255544f
C138 drain_left.t2 a_n1992_n2688# 0.255544f
C139 drain_left.n4 a_n1992_n2688# 2.23832f
C140 drain_left.t1 a_n1992_n2688# 0.255544f
C141 drain_left.t13 a_n1992_n2688# 0.255544f
C142 drain_left.n5 a_n1992_n2688# 2.23515f
C143 drain_left.n6 a_n1992_n2688# 0.81395f
C144 drain_left.n7 a_n1992_n2688# 1.91709f
C145 drain_left.t12 a_n1992_n2688# 0.255544f
C146 drain_left.t18 a_n1992_n2688# 0.255544f
C147 drain_left.n8 a_n1992_n2688# 2.23832f
C148 drain_left.t8 a_n1992_n2688# 0.255544f
C149 drain_left.t19 a_n1992_n2688# 0.255544f
C150 drain_left.n9 a_n1992_n2688# 2.23516f
C151 drain_left.n10 a_n1992_n2688# 0.818475f
C152 drain_left.t9 a_n1992_n2688# 0.255544f
C153 drain_left.t0 a_n1992_n2688# 0.255544f
C154 drain_left.n11 a_n1992_n2688# 2.23516f
C155 drain_left.n12 a_n1992_n2688# 0.403584f
C156 drain_left.t10 a_n1992_n2688# 0.255544f
C157 drain_left.t15 a_n1992_n2688# 0.255544f
C158 drain_left.n13 a_n1992_n2688# 2.23516f
C159 drain_left.n14 a_n1992_n2688# 0.403584f
C160 drain_left.t4 a_n1992_n2688# 0.255544f
C161 drain_left.t16 a_n1992_n2688# 0.255544f
C162 drain_left.n15 a_n1992_n2688# 2.23515f
C163 drain_left.n16 a_n1992_n2688# 0.700179f
C164 source.t20 a_n1992_n2688# 2.40445f
C165 source.n0 a_n1992_n2688# 1.37525f
C166 source.t28 a_n1992_n2688# 0.225485f
C167 source.t37 a_n1992_n2688# 0.225485f
C168 source.n1 a_n1992_n2688# 1.88761f
C169 source.n2 a_n1992_n2688# 0.397651f
C170 source.t21 a_n1992_n2688# 0.225485f
C171 source.t29 a_n1992_n2688# 0.225485f
C172 source.n3 a_n1992_n2688# 1.88761f
C173 source.n4 a_n1992_n2688# 0.397651f
C174 source.t34 a_n1992_n2688# 0.225485f
C175 source.t23 a_n1992_n2688# 0.225485f
C176 source.n5 a_n1992_n2688# 1.88761f
C177 source.n6 a_n1992_n2688# 0.397651f
C178 source.t27 a_n1992_n2688# 0.225485f
C179 source.t19 a_n1992_n2688# 0.225485f
C180 source.n7 a_n1992_n2688# 1.88761f
C181 source.n8 a_n1992_n2688# 0.397651f
C182 source.t30 a_n1992_n2688# 2.40446f
C183 source.n9 a_n1992_n2688# 0.492684f
C184 source.t4 a_n1992_n2688# 2.40446f
C185 source.n10 a_n1992_n2688# 0.492684f
C186 source.t39 a_n1992_n2688# 0.225485f
C187 source.t2 a_n1992_n2688# 0.225485f
C188 source.n11 a_n1992_n2688# 1.88761f
C189 source.n12 a_n1992_n2688# 0.397651f
C190 source.t9 a_n1992_n2688# 0.225485f
C191 source.t3 a_n1992_n2688# 0.225485f
C192 source.n13 a_n1992_n2688# 1.88761f
C193 source.n14 a_n1992_n2688# 0.397651f
C194 source.t11 a_n1992_n2688# 0.225485f
C195 source.t10 a_n1992_n2688# 0.225485f
C196 source.n15 a_n1992_n2688# 1.88761f
C197 source.n16 a_n1992_n2688# 0.397651f
C198 source.t14 a_n1992_n2688# 0.225485f
C199 source.t6 a_n1992_n2688# 0.225485f
C200 source.n17 a_n1992_n2688# 1.88761f
C201 source.n18 a_n1992_n2688# 0.397651f
C202 source.t12 a_n1992_n2688# 2.40446f
C203 source.n19 a_n1992_n2688# 1.83448f
C204 source.t22 a_n1992_n2688# 2.40445f
C205 source.n20 a_n1992_n2688# 1.83449f
C206 source.t25 a_n1992_n2688# 0.225485f
C207 source.t36 a_n1992_n2688# 0.225485f
C208 source.n21 a_n1992_n2688# 1.88761f
C209 source.n22 a_n1992_n2688# 0.397657f
C210 source.t18 a_n1992_n2688# 0.225485f
C211 source.t35 a_n1992_n2688# 0.225485f
C212 source.n23 a_n1992_n2688# 1.88761f
C213 source.n24 a_n1992_n2688# 0.397657f
C214 source.t24 a_n1992_n2688# 0.225485f
C215 source.t26 a_n1992_n2688# 0.225485f
C216 source.n25 a_n1992_n2688# 1.88761f
C217 source.n26 a_n1992_n2688# 0.397657f
C218 source.t32 a_n1992_n2688# 0.225485f
C219 source.t31 a_n1992_n2688# 0.225485f
C220 source.n27 a_n1992_n2688# 1.88761f
C221 source.n28 a_n1992_n2688# 0.397657f
C222 source.t33 a_n1992_n2688# 2.40445f
C223 source.n29 a_n1992_n2688# 0.49269f
C224 source.t13 a_n1992_n2688# 2.40445f
C225 source.n30 a_n1992_n2688# 0.49269f
C226 source.t1 a_n1992_n2688# 0.225485f
C227 source.t0 a_n1992_n2688# 0.225485f
C228 source.n31 a_n1992_n2688# 1.88761f
C229 source.n32 a_n1992_n2688# 0.397657f
C230 source.t17 a_n1992_n2688# 0.225485f
C231 source.t8 a_n1992_n2688# 0.225485f
C232 source.n33 a_n1992_n2688# 1.88761f
C233 source.n34 a_n1992_n2688# 0.397657f
C234 source.t15 a_n1992_n2688# 0.225485f
C235 source.t5 a_n1992_n2688# 0.225485f
C236 source.n35 a_n1992_n2688# 1.88761f
C237 source.n36 a_n1992_n2688# 0.397657f
C238 source.t38 a_n1992_n2688# 0.225485f
C239 source.t16 a_n1992_n2688# 0.225485f
C240 source.n37 a_n1992_n2688# 1.88761f
C241 source.n38 a_n1992_n2688# 0.397657f
C242 source.t7 a_n1992_n2688# 2.40445f
C243 source.n39 a_n1992_n2688# 0.668137f
C244 source.n40 a_n1992_n2688# 1.64813f
C245 plus.n0 a_n1992_n2688# 0.051799f
C246 plus.t15 a_n1992_n2688# 0.330248f
C247 plus.t4 a_n1992_n2688# 0.330248f
C248 plus.t9 a_n1992_n2688# 0.330248f
C249 plus.n1 a_n1992_n2688# 0.140567f
C250 plus.n2 a_n1992_n2688# 0.051799f
C251 plus.t19 a_n1992_n2688# 0.330248f
C252 plus.t10 a_n1992_n2688# 0.330248f
C253 plus.n3 a_n1992_n2688# 0.140567f
C254 plus.n4 a_n1992_n2688# 0.051799f
C255 plus.t0 a_n1992_n2688# 0.330248f
C256 plus.t11 a_n1992_n2688# 0.330248f
C257 plus.t1 a_n1992_n2688# 0.330248f
C258 plus.n5 a_n1992_n2688# 0.140567f
C259 plus.t7 a_n1992_n2688# 0.337494f
C260 plus.n6 a_n1992_n2688# 0.15665f
C261 plus.n7 a_n1992_n2688# 0.118529f
C262 plus.n8 a_n1992_n2688# 0.019738f
C263 plus.n9 a_n1992_n2688# 0.140567f
C264 plus.n10 a_n1992_n2688# 0.019738f
C265 plus.n11 a_n1992_n2688# 0.140567f
C266 plus.n12 a_n1992_n2688# 0.019738f
C267 plus.n13 a_n1992_n2688# 0.051799f
C268 plus.n14 a_n1992_n2688# 0.051799f
C269 plus.n15 a_n1992_n2688# 0.018461f
C270 plus.n16 a_n1992_n2688# 0.018461f
C271 plus.n17 a_n1992_n2688# 0.140567f
C272 plus.n18 a_n1992_n2688# 0.019738f
C273 plus.n19 a_n1992_n2688# 0.051799f
C274 plus.n20 a_n1992_n2688# 0.051799f
C275 plus.n21 a_n1992_n2688# 0.019738f
C276 plus.n22 a_n1992_n2688# 0.140567f
C277 plus.n23 a_n1992_n2688# 0.019738f
C278 plus.n24 a_n1992_n2688# 0.140567f
C279 plus.t3 a_n1992_n2688# 0.337494f
C280 plus.n25 a_n1992_n2688# 0.156572f
C281 plus.n26 a_n1992_n2688# 0.508403f
C282 plus.n27 a_n1992_n2688# 0.051799f
C283 plus.t8 a_n1992_n2688# 0.337494f
C284 plus.t14 a_n1992_n2688# 0.330248f
C285 plus.t5 a_n1992_n2688# 0.330248f
C286 plus.t12 a_n1992_n2688# 0.330248f
C287 plus.n28 a_n1992_n2688# 0.140567f
C288 plus.n29 a_n1992_n2688# 0.051799f
C289 plus.t16 a_n1992_n2688# 0.330248f
C290 plus.t2 a_n1992_n2688# 0.330248f
C291 plus.n30 a_n1992_n2688# 0.140567f
C292 plus.n31 a_n1992_n2688# 0.051799f
C293 plus.t18 a_n1992_n2688# 0.330248f
C294 plus.t6 a_n1992_n2688# 0.330248f
C295 plus.t13 a_n1992_n2688# 0.330248f
C296 plus.n32 a_n1992_n2688# 0.140567f
C297 plus.t17 a_n1992_n2688# 0.337494f
C298 plus.n33 a_n1992_n2688# 0.15665f
C299 plus.n34 a_n1992_n2688# 0.118529f
C300 plus.n35 a_n1992_n2688# 0.019738f
C301 plus.n36 a_n1992_n2688# 0.140567f
C302 plus.n37 a_n1992_n2688# 0.019738f
C303 plus.n38 a_n1992_n2688# 0.140567f
C304 plus.n39 a_n1992_n2688# 0.019738f
C305 plus.n40 a_n1992_n2688# 0.051799f
C306 plus.n41 a_n1992_n2688# 0.051799f
C307 plus.n42 a_n1992_n2688# 0.018461f
C308 plus.n43 a_n1992_n2688# 0.018461f
C309 plus.n44 a_n1992_n2688# 0.140567f
C310 plus.n45 a_n1992_n2688# 0.019738f
C311 plus.n46 a_n1992_n2688# 0.051799f
C312 plus.n47 a_n1992_n2688# 0.051799f
C313 plus.n48 a_n1992_n2688# 0.019738f
C314 plus.n49 a_n1992_n2688# 0.140567f
C315 plus.n50 a_n1992_n2688# 0.019738f
C316 plus.n51 a_n1992_n2688# 0.140567f
C317 plus.n52 a_n1992_n2688# 0.156572f
C318 plus.n53 a_n1992_n2688# 1.47347f
.ends

