* NGSPICE file created from diffpair312.ext - technology: sky130A

.subckt diffpair312 minus drain_right drain_left source plus
X0 source.t11 plus.t0 drain_left.t2 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X1 source.t2 minus.t0 drain_right.t5 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X3 drain_left.t3 plus.t1 source.t10 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X4 a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X5 drain_right.t4 minus.t1 source.t3 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X6 drain_right.t3 minus.t2 source.t5 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X7 drain_left.t1 plus.t2 source.t9 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X8 source.t0 minus.t3 drain_right.t2 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X9 drain_right.t1 minus.t4 source.t1 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X10 drain_right.t0 minus.t5 source.t4 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X11 drain_left.t0 plus.t3 source.t8 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X12 a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X13 source.t7 plus.t4 drain_left.t5 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X14 drain_left.t4 plus.t5 source.t6 a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X15 a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# a_n1620_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
R0 plus.n1 plus.t5 253.34
R1 plus.n7 plus.t2 253.34
R2 plus.n4 plus.t3 229.855
R3 plus.n2 plus.t4 229.855
R4 plus.n10 plus.t1 229.855
R5 plus.n8 plus.t0 229.855
R6 plus.n3 plus.n0 161.3
R7 plus.n5 plus.n4 161.3
R8 plus.n9 plus.n6 161.3
R9 plus.n11 plus.n10 161.3
R10 plus.n7 plus.n6 44.8973
R11 plus.n1 plus.n0 44.8973
R12 plus.n4 plus.n3 33.5944
R13 plus.n10 plus.n9 33.5944
R14 plus plus.n11 27.088
R15 plus.n8 plus.n7 18.1882
R16 plus.n2 plus.n1 18.1882
R17 plus.n3 plus.n2 14.6066
R18 plus.n9 plus.n8 14.6066
R19 plus plus.n5 10.0933
R20 plus.n5 plus.n0 0.189894
R21 plus.n11 plus.n6 0.189894
R22 drain_left.n26 drain_left.n0 289.615
R23 drain_left.n59 drain_left.n33 289.615
R24 drain_left.n11 drain_left.n10 185
R25 drain_left.n8 drain_left.n7 185
R26 drain_left.n17 drain_left.n16 185
R27 drain_left.n19 drain_left.n18 185
R28 drain_left.n4 drain_left.n3 185
R29 drain_left.n25 drain_left.n24 185
R30 drain_left.n27 drain_left.n26 185
R31 drain_left.n60 drain_left.n59 185
R32 drain_left.n58 drain_left.n57 185
R33 drain_left.n37 drain_left.n36 185
R34 drain_left.n52 drain_left.n51 185
R35 drain_left.n50 drain_left.n49 185
R36 drain_left.n41 drain_left.n40 185
R37 drain_left.n44 drain_left.n43 185
R38 drain_left.t3 drain_left.n9 147.661
R39 drain_left.t4 drain_left.n42 147.661
R40 drain_left.n10 drain_left.n7 104.615
R41 drain_left.n17 drain_left.n7 104.615
R42 drain_left.n18 drain_left.n17 104.615
R43 drain_left.n18 drain_left.n3 104.615
R44 drain_left.n25 drain_left.n3 104.615
R45 drain_left.n26 drain_left.n25 104.615
R46 drain_left.n59 drain_left.n58 104.615
R47 drain_left.n58 drain_left.n36 104.615
R48 drain_left.n51 drain_left.n36 104.615
R49 drain_left.n51 drain_left.n50 104.615
R50 drain_left.n50 drain_left.n40 104.615
R51 drain_left.n43 drain_left.n40 104.615
R52 drain_left.n32 drain_left.n31 67.3788
R53 drain_left.n65 drain_left.n64 67.1907
R54 drain_left.n10 drain_left.t3 52.3082
R55 drain_left.n43 drain_left.t4 52.3082
R56 drain_left.n65 drain_left.n63 49.8383
R57 drain_left.n32 drain_left.n30 49.5394
R58 drain_left drain_left.n32 25.5005
R59 drain_left.n11 drain_left.n9 15.6674
R60 drain_left.n44 drain_left.n42 15.6674
R61 drain_left.n12 drain_left.n8 12.8005
R62 drain_left.n45 drain_left.n41 12.8005
R63 drain_left.n16 drain_left.n15 12.0247
R64 drain_left.n49 drain_left.n48 12.0247
R65 drain_left.n19 drain_left.n6 11.249
R66 drain_left.n52 drain_left.n39 11.249
R67 drain_left.n20 drain_left.n4 10.4732
R68 drain_left.n53 drain_left.n37 10.4732
R69 drain_left.n24 drain_left.n23 9.69747
R70 drain_left.n57 drain_left.n56 9.69747
R71 drain_left.n30 drain_left.n29 9.45567
R72 drain_left.n63 drain_left.n62 9.45567
R73 drain_left.n29 drain_left.n28 9.3005
R74 drain_left.n2 drain_left.n1 9.3005
R75 drain_left.n23 drain_left.n22 9.3005
R76 drain_left.n21 drain_left.n20 9.3005
R77 drain_left.n6 drain_left.n5 9.3005
R78 drain_left.n15 drain_left.n14 9.3005
R79 drain_left.n13 drain_left.n12 9.3005
R80 drain_left.n62 drain_left.n61 9.3005
R81 drain_left.n35 drain_left.n34 9.3005
R82 drain_left.n56 drain_left.n55 9.3005
R83 drain_left.n54 drain_left.n53 9.3005
R84 drain_left.n39 drain_left.n38 9.3005
R85 drain_left.n48 drain_left.n47 9.3005
R86 drain_left.n46 drain_left.n45 9.3005
R87 drain_left.n27 drain_left.n2 8.92171
R88 drain_left.n60 drain_left.n35 8.92171
R89 drain_left.n28 drain_left.n0 8.14595
R90 drain_left.n61 drain_left.n33 8.14595
R91 drain_left drain_left.n65 6.62735
R92 drain_left.n30 drain_left.n0 5.81868
R93 drain_left.n63 drain_left.n33 5.81868
R94 drain_left.n28 drain_left.n27 5.04292
R95 drain_left.n61 drain_left.n60 5.04292
R96 drain_left.n13 drain_left.n9 4.38594
R97 drain_left.n46 drain_left.n42 4.38594
R98 drain_left.n24 drain_left.n2 4.26717
R99 drain_left.n57 drain_left.n35 4.26717
R100 drain_left.n23 drain_left.n4 3.49141
R101 drain_left.n56 drain_left.n37 3.49141
R102 drain_left.n31 drain_left.t2 3.3005
R103 drain_left.n31 drain_left.t1 3.3005
R104 drain_left.n64 drain_left.t5 3.3005
R105 drain_left.n64 drain_left.t0 3.3005
R106 drain_left.n20 drain_left.n19 2.71565
R107 drain_left.n53 drain_left.n52 2.71565
R108 drain_left.n16 drain_left.n6 1.93989
R109 drain_left.n49 drain_left.n39 1.93989
R110 drain_left.n15 drain_left.n8 1.16414
R111 drain_left.n48 drain_left.n41 1.16414
R112 drain_left.n12 drain_left.n11 0.388379
R113 drain_left.n45 drain_left.n44 0.388379
R114 drain_left.n14 drain_left.n13 0.155672
R115 drain_left.n14 drain_left.n5 0.155672
R116 drain_left.n21 drain_left.n5 0.155672
R117 drain_left.n22 drain_left.n21 0.155672
R118 drain_left.n22 drain_left.n1 0.155672
R119 drain_left.n29 drain_left.n1 0.155672
R120 drain_left.n62 drain_left.n34 0.155672
R121 drain_left.n55 drain_left.n34 0.155672
R122 drain_left.n55 drain_left.n54 0.155672
R123 drain_left.n54 drain_left.n38 0.155672
R124 drain_left.n47 drain_left.n38 0.155672
R125 drain_left.n47 drain_left.n46 0.155672
R126 source.n130 source.n104 289.615
R127 source.n96 source.n70 289.615
R128 source.n26 source.n0 289.615
R129 source.n60 source.n34 289.615
R130 source.n115 source.n114 185
R131 source.n112 source.n111 185
R132 source.n121 source.n120 185
R133 source.n123 source.n122 185
R134 source.n108 source.n107 185
R135 source.n129 source.n128 185
R136 source.n131 source.n130 185
R137 source.n81 source.n80 185
R138 source.n78 source.n77 185
R139 source.n87 source.n86 185
R140 source.n89 source.n88 185
R141 source.n74 source.n73 185
R142 source.n95 source.n94 185
R143 source.n97 source.n96 185
R144 source.n27 source.n26 185
R145 source.n25 source.n24 185
R146 source.n4 source.n3 185
R147 source.n19 source.n18 185
R148 source.n17 source.n16 185
R149 source.n8 source.n7 185
R150 source.n11 source.n10 185
R151 source.n61 source.n60 185
R152 source.n59 source.n58 185
R153 source.n38 source.n37 185
R154 source.n53 source.n52 185
R155 source.n51 source.n50 185
R156 source.n42 source.n41 185
R157 source.n45 source.n44 185
R158 source.t3 source.n113 147.661
R159 source.t9 source.n79 147.661
R160 source.t8 source.n9 147.661
R161 source.t4 source.n43 147.661
R162 source.n114 source.n111 104.615
R163 source.n121 source.n111 104.615
R164 source.n122 source.n121 104.615
R165 source.n122 source.n107 104.615
R166 source.n129 source.n107 104.615
R167 source.n130 source.n129 104.615
R168 source.n80 source.n77 104.615
R169 source.n87 source.n77 104.615
R170 source.n88 source.n87 104.615
R171 source.n88 source.n73 104.615
R172 source.n95 source.n73 104.615
R173 source.n96 source.n95 104.615
R174 source.n26 source.n25 104.615
R175 source.n25 source.n3 104.615
R176 source.n18 source.n3 104.615
R177 source.n18 source.n17 104.615
R178 source.n17 source.n7 104.615
R179 source.n10 source.n7 104.615
R180 source.n60 source.n59 104.615
R181 source.n59 source.n37 104.615
R182 source.n52 source.n37 104.615
R183 source.n52 source.n51 104.615
R184 source.n51 source.n41 104.615
R185 source.n44 source.n41 104.615
R186 source.n114 source.t3 52.3082
R187 source.n80 source.t9 52.3082
R188 source.n10 source.t8 52.3082
R189 source.n44 source.t4 52.3082
R190 source.n33 source.n32 50.512
R191 source.n67 source.n66 50.512
R192 source.n103 source.n102 50.5119
R193 source.n69 source.n68 50.5119
R194 source.n135 source.n134 32.1853
R195 source.n101 source.n100 32.1853
R196 source.n31 source.n30 32.1853
R197 source.n65 source.n64 32.1853
R198 source.n69 source.n67 18.6905
R199 source.n115 source.n113 15.6674
R200 source.n81 source.n79 15.6674
R201 source.n11 source.n9 15.6674
R202 source.n45 source.n43 15.6674
R203 source.n116 source.n112 12.8005
R204 source.n82 source.n78 12.8005
R205 source.n12 source.n8 12.8005
R206 source.n46 source.n42 12.8005
R207 source.n120 source.n119 12.0247
R208 source.n86 source.n85 12.0247
R209 source.n16 source.n15 12.0247
R210 source.n50 source.n49 12.0247
R211 source.n136 source.n31 11.9664
R212 source.n123 source.n110 11.249
R213 source.n89 source.n76 11.249
R214 source.n19 source.n6 11.249
R215 source.n53 source.n40 11.249
R216 source.n124 source.n108 10.4732
R217 source.n90 source.n74 10.4732
R218 source.n20 source.n4 10.4732
R219 source.n54 source.n38 10.4732
R220 source.n128 source.n127 9.69747
R221 source.n94 source.n93 9.69747
R222 source.n24 source.n23 9.69747
R223 source.n58 source.n57 9.69747
R224 source.n134 source.n133 9.45567
R225 source.n100 source.n99 9.45567
R226 source.n30 source.n29 9.45567
R227 source.n64 source.n63 9.45567
R228 source.n133 source.n132 9.3005
R229 source.n106 source.n105 9.3005
R230 source.n127 source.n126 9.3005
R231 source.n125 source.n124 9.3005
R232 source.n110 source.n109 9.3005
R233 source.n119 source.n118 9.3005
R234 source.n117 source.n116 9.3005
R235 source.n99 source.n98 9.3005
R236 source.n72 source.n71 9.3005
R237 source.n93 source.n92 9.3005
R238 source.n91 source.n90 9.3005
R239 source.n76 source.n75 9.3005
R240 source.n85 source.n84 9.3005
R241 source.n83 source.n82 9.3005
R242 source.n29 source.n28 9.3005
R243 source.n2 source.n1 9.3005
R244 source.n23 source.n22 9.3005
R245 source.n21 source.n20 9.3005
R246 source.n6 source.n5 9.3005
R247 source.n15 source.n14 9.3005
R248 source.n13 source.n12 9.3005
R249 source.n63 source.n62 9.3005
R250 source.n36 source.n35 9.3005
R251 source.n57 source.n56 9.3005
R252 source.n55 source.n54 9.3005
R253 source.n40 source.n39 9.3005
R254 source.n49 source.n48 9.3005
R255 source.n47 source.n46 9.3005
R256 source.n131 source.n106 8.92171
R257 source.n97 source.n72 8.92171
R258 source.n27 source.n2 8.92171
R259 source.n61 source.n36 8.92171
R260 source.n132 source.n104 8.14595
R261 source.n98 source.n70 8.14595
R262 source.n28 source.n0 8.14595
R263 source.n62 source.n34 8.14595
R264 source.n134 source.n104 5.81868
R265 source.n100 source.n70 5.81868
R266 source.n30 source.n0 5.81868
R267 source.n64 source.n34 5.81868
R268 source.n136 source.n135 5.7505
R269 source.n132 source.n131 5.04292
R270 source.n98 source.n97 5.04292
R271 source.n28 source.n27 5.04292
R272 source.n62 source.n61 5.04292
R273 source.n117 source.n113 4.38594
R274 source.n83 source.n79 4.38594
R275 source.n13 source.n9 4.38594
R276 source.n47 source.n43 4.38594
R277 source.n128 source.n106 4.26717
R278 source.n94 source.n72 4.26717
R279 source.n24 source.n2 4.26717
R280 source.n58 source.n36 4.26717
R281 source.n127 source.n108 3.49141
R282 source.n93 source.n74 3.49141
R283 source.n23 source.n4 3.49141
R284 source.n57 source.n38 3.49141
R285 source.n102 source.t1 3.3005
R286 source.n102 source.t2 3.3005
R287 source.n68 source.t10 3.3005
R288 source.n68 source.t11 3.3005
R289 source.n32 source.t6 3.3005
R290 source.n32 source.t7 3.3005
R291 source.n66 source.t5 3.3005
R292 source.n66 source.t0 3.3005
R293 source.n124 source.n123 2.71565
R294 source.n90 source.n89 2.71565
R295 source.n20 source.n19 2.71565
R296 source.n54 source.n53 2.71565
R297 source.n120 source.n110 1.93989
R298 source.n86 source.n76 1.93989
R299 source.n16 source.n6 1.93989
R300 source.n50 source.n40 1.93989
R301 source.n119 source.n112 1.16414
R302 source.n85 source.n78 1.16414
R303 source.n15 source.n8 1.16414
R304 source.n49 source.n42 1.16414
R305 source.n67 source.n65 0.974638
R306 source.n33 source.n31 0.974638
R307 source.n101 source.n69 0.974638
R308 source.n135 source.n103 0.974638
R309 source.n65 source.n33 0.957397
R310 source.n103 source.n101 0.957397
R311 source.n116 source.n115 0.388379
R312 source.n82 source.n81 0.388379
R313 source.n12 source.n11 0.388379
R314 source.n46 source.n45 0.388379
R315 source source.n136 0.188
R316 source.n118 source.n117 0.155672
R317 source.n118 source.n109 0.155672
R318 source.n125 source.n109 0.155672
R319 source.n126 source.n125 0.155672
R320 source.n126 source.n105 0.155672
R321 source.n133 source.n105 0.155672
R322 source.n84 source.n83 0.155672
R323 source.n84 source.n75 0.155672
R324 source.n91 source.n75 0.155672
R325 source.n92 source.n91 0.155672
R326 source.n92 source.n71 0.155672
R327 source.n99 source.n71 0.155672
R328 source.n29 source.n1 0.155672
R329 source.n22 source.n1 0.155672
R330 source.n22 source.n21 0.155672
R331 source.n21 source.n5 0.155672
R332 source.n14 source.n5 0.155672
R333 source.n14 source.n13 0.155672
R334 source.n63 source.n35 0.155672
R335 source.n56 source.n35 0.155672
R336 source.n56 source.n55 0.155672
R337 source.n55 source.n39 0.155672
R338 source.n48 source.n39 0.155672
R339 source.n48 source.n47 0.155672
R340 minus.n1 minus.t5 253.34
R341 minus.n7 minus.t4 253.34
R342 minus.n2 minus.t3 229.855
R343 minus.n4 minus.t2 229.855
R344 minus.n8 minus.t0 229.855
R345 minus.n10 minus.t1 229.855
R346 minus.n5 minus.n4 161.3
R347 minus.n3 minus.n0 161.3
R348 minus.n11 minus.n10 161.3
R349 minus.n9 minus.n6 161.3
R350 minus.n1 minus.n0 44.8973
R351 minus.n7 minus.n6 44.8973
R352 minus.n4 minus.n3 33.5944
R353 minus.n10 minus.n9 33.5944
R354 minus.n12 minus.n5 30.9342
R355 minus.n2 minus.n1 18.1882
R356 minus.n8 minus.n7 18.1882
R357 minus.n3 minus.n2 14.6066
R358 minus.n9 minus.n8 14.6066
R359 minus.n12 minus.n11 6.72209
R360 minus.n5 minus.n0 0.189894
R361 minus.n11 minus.n6 0.189894
R362 minus minus.n12 0.188
R363 drain_right.n26 drain_right.n0 289.615
R364 drain_right.n60 drain_right.n34 289.615
R365 drain_right.n11 drain_right.n10 185
R366 drain_right.n8 drain_right.n7 185
R367 drain_right.n17 drain_right.n16 185
R368 drain_right.n19 drain_right.n18 185
R369 drain_right.n4 drain_right.n3 185
R370 drain_right.n25 drain_right.n24 185
R371 drain_right.n27 drain_right.n26 185
R372 drain_right.n61 drain_right.n60 185
R373 drain_right.n59 drain_right.n58 185
R374 drain_right.n38 drain_right.n37 185
R375 drain_right.n53 drain_right.n52 185
R376 drain_right.n51 drain_right.n50 185
R377 drain_right.n42 drain_right.n41 185
R378 drain_right.n45 drain_right.n44 185
R379 drain_right.t1 drain_right.n9 147.661
R380 drain_right.t3 drain_right.n43 147.661
R381 drain_right.n10 drain_right.n7 104.615
R382 drain_right.n17 drain_right.n7 104.615
R383 drain_right.n18 drain_right.n17 104.615
R384 drain_right.n18 drain_right.n3 104.615
R385 drain_right.n25 drain_right.n3 104.615
R386 drain_right.n26 drain_right.n25 104.615
R387 drain_right.n60 drain_right.n59 104.615
R388 drain_right.n59 drain_right.n37 104.615
R389 drain_right.n52 drain_right.n37 104.615
R390 drain_right.n52 drain_right.n51 104.615
R391 drain_right.n51 drain_right.n41 104.615
R392 drain_right.n44 drain_right.n41 104.615
R393 drain_right.n65 drain_right.n33 68.1648
R394 drain_right.n32 drain_right.n31 67.3788
R395 drain_right.n10 drain_right.t1 52.3082
R396 drain_right.n44 drain_right.t3 52.3082
R397 drain_right.n32 drain_right.n30 49.5394
R398 drain_right.n65 drain_right.n64 48.8641
R399 drain_right drain_right.n32 24.9473
R400 drain_right.n11 drain_right.n9 15.6674
R401 drain_right.n45 drain_right.n43 15.6674
R402 drain_right.n12 drain_right.n8 12.8005
R403 drain_right.n46 drain_right.n42 12.8005
R404 drain_right.n16 drain_right.n15 12.0247
R405 drain_right.n50 drain_right.n49 12.0247
R406 drain_right.n19 drain_right.n6 11.249
R407 drain_right.n53 drain_right.n40 11.249
R408 drain_right.n20 drain_right.n4 10.4732
R409 drain_right.n54 drain_right.n38 10.4732
R410 drain_right.n24 drain_right.n23 9.69747
R411 drain_right.n58 drain_right.n57 9.69747
R412 drain_right.n30 drain_right.n29 9.45567
R413 drain_right.n64 drain_right.n63 9.45567
R414 drain_right.n29 drain_right.n28 9.3005
R415 drain_right.n2 drain_right.n1 9.3005
R416 drain_right.n23 drain_right.n22 9.3005
R417 drain_right.n21 drain_right.n20 9.3005
R418 drain_right.n6 drain_right.n5 9.3005
R419 drain_right.n15 drain_right.n14 9.3005
R420 drain_right.n13 drain_right.n12 9.3005
R421 drain_right.n63 drain_right.n62 9.3005
R422 drain_right.n36 drain_right.n35 9.3005
R423 drain_right.n57 drain_right.n56 9.3005
R424 drain_right.n55 drain_right.n54 9.3005
R425 drain_right.n40 drain_right.n39 9.3005
R426 drain_right.n49 drain_right.n48 9.3005
R427 drain_right.n47 drain_right.n46 9.3005
R428 drain_right.n27 drain_right.n2 8.92171
R429 drain_right.n61 drain_right.n36 8.92171
R430 drain_right.n28 drain_right.n0 8.14595
R431 drain_right.n62 drain_right.n34 8.14595
R432 drain_right drain_right.n65 6.14028
R433 drain_right.n30 drain_right.n0 5.81868
R434 drain_right.n64 drain_right.n34 5.81868
R435 drain_right.n28 drain_right.n27 5.04292
R436 drain_right.n62 drain_right.n61 5.04292
R437 drain_right.n13 drain_right.n9 4.38594
R438 drain_right.n47 drain_right.n43 4.38594
R439 drain_right.n24 drain_right.n2 4.26717
R440 drain_right.n58 drain_right.n36 4.26717
R441 drain_right.n23 drain_right.n4 3.49141
R442 drain_right.n57 drain_right.n38 3.49141
R443 drain_right.n31 drain_right.t5 3.3005
R444 drain_right.n31 drain_right.t4 3.3005
R445 drain_right.n33 drain_right.t2 3.3005
R446 drain_right.n33 drain_right.t0 3.3005
R447 drain_right.n20 drain_right.n19 2.71565
R448 drain_right.n54 drain_right.n53 2.71565
R449 drain_right.n16 drain_right.n6 1.93989
R450 drain_right.n50 drain_right.n40 1.93989
R451 drain_right.n15 drain_right.n8 1.16414
R452 drain_right.n49 drain_right.n42 1.16414
R453 drain_right.n12 drain_right.n11 0.388379
R454 drain_right.n46 drain_right.n45 0.388379
R455 drain_right.n14 drain_right.n13 0.155672
R456 drain_right.n14 drain_right.n5 0.155672
R457 drain_right.n21 drain_right.n5 0.155672
R458 drain_right.n22 drain_right.n21 0.155672
R459 drain_right.n22 drain_right.n1 0.155672
R460 drain_right.n29 drain_right.n1 0.155672
R461 drain_right.n63 drain_right.n35 0.155672
R462 drain_right.n56 drain_right.n35 0.155672
R463 drain_right.n56 drain_right.n55 0.155672
R464 drain_right.n55 drain_right.n39 0.155672
R465 drain_right.n48 drain_right.n39 0.155672
R466 drain_right.n48 drain_right.n47 0.155672
C0 source minus 2.50993f
C1 minus drain_right 2.49345f
C2 minus drain_left 0.171398f
C3 plus minus 4.04278f
C4 source drain_right 5.80768f
C5 source drain_left 5.81f
C6 drain_left drain_right 0.74366f
C7 source plus 2.52418f
C8 plus drain_right 0.311011f
C9 plus drain_left 2.64803f
C10 drain_right a_n1620_n2088# 4.71352f
C11 drain_left a_n1620_n2088# 4.958321f
C12 source a_n1620_n2088# 4.11118f
C13 minus a_n1620_n2088# 5.697762f
C14 plus a_n1620_n2088# 7.03694f
C15 drain_right.n0 a_n1620_n2088# 0.032082f
C16 drain_right.n1 a_n1620_n2088# 0.022825f
C17 drain_right.n2 a_n1620_n2088# 0.012265f
C18 drain_right.n3 a_n1620_n2088# 0.02899f
C19 drain_right.n4 a_n1620_n2088# 0.012987f
C20 drain_right.n5 a_n1620_n2088# 0.022825f
C21 drain_right.n6 a_n1620_n2088# 0.012265f
C22 drain_right.n7 a_n1620_n2088# 0.02899f
C23 drain_right.n8 a_n1620_n2088# 0.012987f
C24 drain_right.n9 a_n1620_n2088# 0.097674f
C25 drain_right.t1 a_n1620_n2088# 0.04725f
C26 drain_right.n10 a_n1620_n2088# 0.021743f
C27 drain_right.n11 a_n1620_n2088# 0.017124f
C28 drain_right.n12 a_n1620_n2088# 0.012265f
C29 drain_right.n13 a_n1620_n2088# 0.543095f
C30 drain_right.n14 a_n1620_n2088# 0.022825f
C31 drain_right.n15 a_n1620_n2088# 0.012265f
C32 drain_right.n16 a_n1620_n2088# 0.012987f
C33 drain_right.n17 a_n1620_n2088# 0.02899f
C34 drain_right.n18 a_n1620_n2088# 0.02899f
C35 drain_right.n19 a_n1620_n2088# 0.012987f
C36 drain_right.n20 a_n1620_n2088# 0.012265f
C37 drain_right.n21 a_n1620_n2088# 0.022825f
C38 drain_right.n22 a_n1620_n2088# 0.022825f
C39 drain_right.n23 a_n1620_n2088# 0.012265f
C40 drain_right.n24 a_n1620_n2088# 0.012987f
C41 drain_right.n25 a_n1620_n2088# 0.02899f
C42 drain_right.n26 a_n1620_n2088# 0.062759f
C43 drain_right.n27 a_n1620_n2088# 0.012987f
C44 drain_right.n28 a_n1620_n2088# 0.012265f
C45 drain_right.n29 a_n1620_n2088# 0.052759f
C46 drain_right.n30 a_n1620_n2088# 0.052163f
C47 drain_right.t5 a_n1620_n2088# 0.108221f
C48 drain_right.t4 a_n1620_n2088# 0.108221f
C49 drain_right.n31 a_n1620_n2088# 0.903357f
C50 drain_right.n32 a_n1620_n2088# 1.12156f
C51 drain_right.t2 a_n1620_n2088# 0.108221f
C52 drain_right.t0 a_n1620_n2088# 0.108221f
C53 drain_right.n33 a_n1620_n2088# 0.907393f
C54 drain_right.n34 a_n1620_n2088# 0.032082f
C55 drain_right.n35 a_n1620_n2088# 0.022825f
C56 drain_right.n36 a_n1620_n2088# 0.012265f
C57 drain_right.n37 a_n1620_n2088# 0.02899f
C58 drain_right.n38 a_n1620_n2088# 0.012987f
C59 drain_right.n39 a_n1620_n2088# 0.022825f
C60 drain_right.n40 a_n1620_n2088# 0.012265f
C61 drain_right.n41 a_n1620_n2088# 0.02899f
C62 drain_right.n42 a_n1620_n2088# 0.012987f
C63 drain_right.n43 a_n1620_n2088# 0.097674f
C64 drain_right.t3 a_n1620_n2088# 0.04725f
C65 drain_right.n44 a_n1620_n2088# 0.021743f
C66 drain_right.n45 a_n1620_n2088# 0.017124f
C67 drain_right.n46 a_n1620_n2088# 0.012265f
C68 drain_right.n47 a_n1620_n2088# 0.543095f
C69 drain_right.n48 a_n1620_n2088# 0.022825f
C70 drain_right.n49 a_n1620_n2088# 0.012265f
C71 drain_right.n50 a_n1620_n2088# 0.012987f
C72 drain_right.n51 a_n1620_n2088# 0.02899f
C73 drain_right.n52 a_n1620_n2088# 0.02899f
C74 drain_right.n53 a_n1620_n2088# 0.012987f
C75 drain_right.n54 a_n1620_n2088# 0.012265f
C76 drain_right.n55 a_n1620_n2088# 0.022825f
C77 drain_right.n56 a_n1620_n2088# 0.022825f
C78 drain_right.n57 a_n1620_n2088# 0.012265f
C79 drain_right.n58 a_n1620_n2088# 0.012987f
C80 drain_right.n59 a_n1620_n2088# 0.02899f
C81 drain_right.n60 a_n1620_n2088# 0.062759f
C82 drain_right.n61 a_n1620_n2088# 0.012987f
C83 drain_right.n62 a_n1620_n2088# 0.012265f
C84 drain_right.n63 a_n1620_n2088# 0.052759f
C85 drain_right.n64 a_n1620_n2088# 0.050876f
C86 drain_right.n65 a_n1620_n2088# 0.66306f
C87 minus.n0 a_n1620_n2088# 0.194242f
C88 minus.t5 a_n1620_n2088# 0.652168f
C89 minus.n1 a_n1620_n2088# 0.26506f
C90 minus.t3 a_n1620_n2088# 0.625498f
C91 minus.n2 a_n1620_n2088# 0.290128f
C92 minus.n3 a_n1620_n2088# 0.010195f
C93 minus.t2 a_n1620_n2088# 0.625498f
C94 minus.n4 a_n1620_n2088# 0.28576f
C95 minus.n5 a_n1620_n2088# 1.24007f
C96 minus.n6 a_n1620_n2088# 0.194242f
C97 minus.t4 a_n1620_n2088# 0.652168f
C98 minus.n7 a_n1620_n2088# 0.26506f
C99 minus.t0 a_n1620_n2088# 0.625498f
C100 minus.n8 a_n1620_n2088# 0.290128f
C101 minus.n9 a_n1620_n2088# 0.010195f
C102 minus.t1 a_n1620_n2088# 0.625498f
C103 minus.n10 a_n1620_n2088# 0.28576f
C104 minus.n11 a_n1620_n2088# 0.316985f
C105 minus.n12 a_n1620_n2088# 1.51635f
C106 source.n0 a_n1620_n2088# 0.035913f
C107 source.n1 a_n1620_n2088# 0.02555f
C108 source.n2 a_n1620_n2088# 0.01373f
C109 source.n3 a_n1620_n2088# 0.032452f
C110 source.n4 a_n1620_n2088# 0.014537f
C111 source.n5 a_n1620_n2088# 0.02555f
C112 source.n6 a_n1620_n2088# 0.01373f
C113 source.n7 a_n1620_n2088# 0.032452f
C114 source.n8 a_n1620_n2088# 0.014537f
C115 source.n9 a_n1620_n2088# 0.109338f
C116 source.t8 a_n1620_n2088# 0.052892f
C117 source.n10 a_n1620_n2088# 0.024339f
C118 source.n11 a_n1620_n2088# 0.019169f
C119 source.n12 a_n1620_n2088# 0.01373f
C120 source.n13 a_n1620_n2088# 0.607946f
C121 source.n14 a_n1620_n2088# 0.02555f
C122 source.n15 a_n1620_n2088# 0.01373f
C123 source.n16 a_n1620_n2088# 0.014537f
C124 source.n17 a_n1620_n2088# 0.032452f
C125 source.n18 a_n1620_n2088# 0.032452f
C126 source.n19 a_n1620_n2088# 0.014537f
C127 source.n20 a_n1620_n2088# 0.01373f
C128 source.n21 a_n1620_n2088# 0.02555f
C129 source.n22 a_n1620_n2088# 0.02555f
C130 source.n23 a_n1620_n2088# 0.01373f
C131 source.n24 a_n1620_n2088# 0.014537f
C132 source.n25 a_n1620_n2088# 0.032452f
C133 source.n26 a_n1620_n2088# 0.070253f
C134 source.n27 a_n1620_n2088# 0.014537f
C135 source.n28 a_n1620_n2088# 0.01373f
C136 source.n29 a_n1620_n2088# 0.059058f
C137 source.n30 a_n1620_n2088# 0.039309f
C138 source.n31 a_n1620_n2088# 0.679586f
C139 source.t6 a_n1620_n2088# 0.121144f
C140 source.t7 a_n1620_n2088# 0.121144f
C141 source.n32 a_n1620_n2088# 0.943479f
C142 source.n33 a_n1620_n2088# 0.39849f
C143 source.n34 a_n1620_n2088# 0.035913f
C144 source.n35 a_n1620_n2088# 0.02555f
C145 source.n36 a_n1620_n2088# 0.01373f
C146 source.n37 a_n1620_n2088# 0.032452f
C147 source.n38 a_n1620_n2088# 0.014537f
C148 source.n39 a_n1620_n2088# 0.02555f
C149 source.n40 a_n1620_n2088# 0.01373f
C150 source.n41 a_n1620_n2088# 0.032452f
C151 source.n42 a_n1620_n2088# 0.014537f
C152 source.n43 a_n1620_n2088# 0.109338f
C153 source.t4 a_n1620_n2088# 0.052892f
C154 source.n44 a_n1620_n2088# 0.024339f
C155 source.n45 a_n1620_n2088# 0.019169f
C156 source.n46 a_n1620_n2088# 0.01373f
C157 source.n47 a_n1620_n2088# 0.607946f
C158 source.n48 a_n1620_n2088# 0.02555f
C159 source.n49 a_n1620_n2088# 0.01373f
C160 source.n50 a_n1620_n2088# 0.014537f
C161 source.n51 a_n1620_n2088# 0.032452f
C162 source.n52 a_n1620_n2088# 0.032452f
C163 source.n53 a_n1620_n2088# 0.014537f
C164 source.n54 a_n1620_n2088# 0.01373f
C165 source.n55 a_n1620_n2088# 0.02555f
C166 source.n56 a_n1620_n2088# 0.02555f
C167 source.n57 a_n1620_n2088# 0.01373f
C168 source.n58 a_n1620_n2088# 0.014537f
C169 source.n59 a_n1620_n2088# 0.032452f
C170 source.n60 a_n1620_n2088# 0.070253f
C171 source.n61 a_n1620_n2088# 0.014537f
C172 source.n62 a_n1620_n2088# 0.01373f
C173 source.n63 a_n1620_n2088# 0.059058f
C174 source.n64 a_n1620_n2088# 0.039309f
C175 source.n65 a_n1620_n2088# 0.180802f
C176 source.t5 a_n1620_n2088# 0.121144f
C177 source.t0 a_n1620_n2088# 0.121144f
C178 source.n66 a_n1620_n2088# 0.943479f
C179 source.n67 a_n1620_n2088# 1.31668f
C180 source.t10 a_n1620_n2088# 0.121144f
C181 source.t11 a_n1620_n2088# 0.121144f
C182 source.n68 a_n1620_n2088# 0.943473f
C183 source.n69 a_n1620_n2088# 1.31668f
C184 source.n70 a_n1620_n2088# 0.035913f
C185 source.n71 a_n1620_n2088# 0.02555f
C186 source.n72 a_n1620_n2088# 0.01373f
C187 source.n73 a_n1620_n2088# 0.032452f
C188 source.n74 a_n1620_n2088# 0.014537f
C189 source.n75 a_n1620_n2088# 0.02555f
C190 source.n76 a_n1620_n2088# 0.01373f
C191 source.n77 a_n1620_n2088# 0.032452f
C192 source.n78 a_n1620_n2088# 0.014537f
C193 source.n79 a_n1620_n2088# 0.109338f
C194 source.t9 a_n1620_n2088# 0.052892f
C195 source.n80 a_n1620_n2088# 0.024339f
C196 source.n81 a_n1620_n2088# 0.019169f
C197 source.n82 a_n1620_n2088# 0.01373f
C198 source.n83 a_n1620_n2088# 0.607946f
C199 source.n84 a_n1620_n2088# 0.02555f
C200 source.n85 a_n1620_n2088# 0.01373f
C201 source.n86 a_n1620_n2088# 0.014537f
C202 source.n87 a_n1620_n2088# 0.032452f
C203 source.n88 a_n1620_n2088# 0.032452f
C204 source.n89 a_n1620_n2088# 0.014537f
C205 source.n90 a_n1620_n2088# 0.01373f
C206 source.n91 a_n1620_n2088# 0.02555f
C207 source.n92 a_n1620_n2088# 0.02555f
C208 source.n93 a_n1620_n2088# 0.01373f
C209 source.n94 a_n1620_n2088# 0.014537f
C210 source.n95 a_n1620_n2088# 0.032452f
C211 source.n96 a_n1620_n2088# 0.070253f
C212 source.n97 a_n1620_n2088# 0.014537f
C213 source.n98 a_n1620_n2088# 0.01373f
C214 source.n99 a_n1620_n2088# 0.059058f
C215 source.n100 a_n1620_n2088# 0.039309f
C216 source.n101 a_n1620_n2088# 0.180802f
C217 source.t1 a_n1620_n2088# 0.121144f
C218 source.t2 a_n1620_n2088# 0.121144f
C219 source.n102 a_n1620_n2088# 0.943473f
C220 source.n103 a_n1620_n2088# 0.398497f
C221 source.n104 a_n1620_n2088# 0.035913f
C222 source.n105 a_n1620_n2088# 0.02555f
C223 source.n106 a_n1620_n2088# 0.01373f
C224 source.n107 a_n1620_n2088# 0.032452f
C225 source.n108 a_n1620_n2088# 0.014537f
C226 source.n109 a_n1620_n2088# 0.02555f
C227 source.n110 a_n1620_n2088# 0.01373f
C228 source.n111 a_n1620_n2088# 0.032452f
C229 source.n112 a_n1620_n2088# 0.014537f
C230 source.n113 a_n1620_n2088# 0.109338f
C231 source.t3 a_n1620_n2088# 0.052892f
C232 source.n114 a_n1620_n2088# 0.024339f
C233 source.n115 a_n1620_n2088# 0.019169f
C234 source.n116 a_n1620_n2088# 0.01373f
C235 source.n117 a_n1620_n2088# 0.607946f
C236 source.n118 a_n1620_n2088# 0.02555f
C237 source.n119 a_n1620_n2088# 0.01373f
C238 source.n120 a_n1620_n2088# 0.014537f
C239 source.n121 a_n1620_n2088# 0.032452f
C240 source.n122 a_n1620_n2088# 0.032452f
C241 source.n123 a_n1620_n2088# 0.014537f
C242 source.n124 a_n1620_n2088# 0.01373f
C243 source.n125 a_n1620_n2088# 0.02555f
C244 source.n126 a_n1620_n2088# 0.02555f
C245 source.n127 a_n1620_n2088# 0.01373f
C246 source.n128 a_n1620_n2088# 0.014537f
C247 source.n129 a_n1620_n2088# 0.032452f
C248 source.n130 a_n1620_n2088# 0.070253f
C249 source.n131 a_n1620_n2088# 0.014537f
C250 source.n132 a_n1620_n2088# 0.01373f
C251 source.n133 a_n1620_n2088# 0.059058f
C252 source.n134 a_n1620_n2088# 0.039309f
C253 source.n135 a_n1620_n2088# 0.312899f
C254 source.n136 a_n1620_n2088# 1.06326f
C255 drain_left.n0 a_n1620_n2088# 0.032123f
C256 drain_left.n1 a_n1620_n2088# 0.022854f
C257 drain_left.n2 a_n1620_n2088# 0.012281f
C258 drain_left.n3 a_n1620_n2088# 0.029027f
C259 drain_left.n4 a_n1620_n2088# 0.013003f
C260 drain_left.n5 a_n1620_n2088# 0.022854f
C261 drain_left.n6 a_n1620_n2088# 0.012281f
C262 drain_left.n7 a_n1620_n2088# 0.029027f
C263 drain_left.n8 a_n1620_n2088# 0.013003f
C264 drain_left.n9 a_n1620_n2088# 0.097799f
C265 drain_left.t3 a_n1620_n2088# 0.047311f
C266 drain_left.n10 a_n1620_n2088# 0.02177f
C267 drain_left.n11 a_n1620_n2088# 0.017146f
C268 drain_left.n12 a_n1620_n2088# 0.012281f
C269 drain_left.n13 a_n1620_n2088# 0.543789f
C270 drain_left.n14 a_n1620_n2088# 0.022854f
C271 drain_left.n15 a_n1620_n2088# 0.012281f
C272 drain_left.n16 a_n1620_n2088# 0.013003f
C273 drain_left.n17 a_n1620_n2088# 0.029027f
C274 drain_left.n18 a_n1620_n2088# 0.029027f
C275 drain_left.n19 a_n1620_n2088# 0.013003f
C276 drain_left.n20 a_n1620_n2088# 0.012281f
C277 drain_left.n21 a_n1620_n2088# 0.022854f
C278 drain_left.n22 a_n1620_n2088# 0.022854f
C279 drain_left.n23 a_n1620_n2088# 0.012281f
C280 drain_left.n24 a_n1620_n2088# 0.013003f
C281 drain_left.n25 a_n1620_n2088# 0.029027f
C282 drain_left.n26 a_n1620_n2088# 0.062839f
C283 drain_left.n27 a_n1620_n2088# 0.013003f
C284 drain_left.n28 a_n1620_n2088# 0.012281f
C285 drain_left.n29 a_n1620_n2088# 0.052826f
C286 drain_left.n30 a_n1620_n2088# 0.052229f
C287 drain_left.t2 a_n1620_n2088# 0.10836f
C288 drain_left.t1 a_n1620_n2088# 0.10836f
C289 drain_left.n31 a_n1620_n2088# 0.90451f
C290 drain_left.n32 a_n1620_n2088# 1.16958f
C291 drain_left.n33 a_n1620_n2088# 0.032123f
C292 drain_left.n34 a_n1620_n2088# 0.022854f
C293 drain_left.n35 a_n1620_n2088# 0.012281f
C294 drain_left.n36 a_n1620_n2088# 0.029027f
C295 drain_left.n37 a_n1620_n2088# 0.013003f
C296 drain_left.n38 a_n1620_n2088# 0.022854f
C297 drain_left.n39 a_n1620_n2088# 0.012281f
C298 drain_left.n40 a_n1620_n2088# 0.029027f
C299 drain_left.n41 a_n1620_n2088# 0.013003f
C300 drain_left.n42 a_n1620_n2088# 0.097799f
C301 drain_left.t4 a_n1620_n2088# 0.047311f
C302 drain_left.n43 a_n1620_n2088# 0.02177f
C303 drain_left.n44 a_n1620_n2088# 0.017146f
C304 drain_left.n45 a_n1620_n2088# 0.012281f
C305 drain_left.n46 a_n1620_n2088# 0.543789f
C306 drain_left.n47 a_n1620_n2088# 0.022854f
C307 drain_left.n48 a_n1620_n2088# 0.012281f
C308 drain_left.n49 a_n1620_n2088# 0.013003f
C309 drain_left.n50 a_n1620_n2088# 0.029027f
C310 drain_left.n51 a_n1620_n2088# 0.029027f
C311 drain_left.n52 a_n1620_n2088# 0.013003f
C312 drain_left.n53 a_n1620_n2088# 0.012281f
C313 drain_left.n54 a_n1620_n2088# 0.022854f
C314 drain_left.n55 a_n1620_n2088# 0.022854f
C315 drain_left.n56 a_n1620_n2088# 0.012281f
C316 drain_left.n57 a_n1620_n2088# 0.013003f
C317 drain_left.n58 a_n1620_n2088# 0.029027f
C318 drain_left.n59 a_n1620_n2088# 0.062839f
C319 drain_left.n60 a_n1620_n2088# 0.013003f
C320 drain_left.n61 a_n1620_n2088# 0.012281f
C321 drain_left.n62 a_n1620_n2088# 0.052826f
C322 drain_left.n63 a_n1620_n2088# 0.053203f
C323 drain_left.t5 a_n1620_n2088# 0.10836f
C324 drain_left.t0 a_n1620_n2088# 0.10836f
C325 drain_left.n64 a_n1620_n2088# 0.903719f
C326 drain_left.n65 a_n1620_n2088# 0.647375f
C327 plus.n0 a_n1620_n2088# 0.198403f
C328 plus.t3 a_n1620_n2088# 0.638897f
C329 plus.t4 a_n1620_n2088# 0.638897f
C330 plus.t5 a_n1620_n2088# 0.666139f
C331 plus.n1 a_n1620_n2088# 0.270738f
C332 plus.n2 a_n1620_n2088# 0.296344f
C333 plus.n3 a_n1620_n2088# 0.010413f
C334 plus.n4 a_n1620_n2088# 0.291881f
C335 plus.n5 a_n1620_n2088# 0.418078f
C336 plus.n6 a_n1620_n2088# 0.198403f
C337 plus.t1 a_n1620_n2088# 0.638897f
C338 plus.t2 a_n1620_n2088# 0.666139f
C339 plus.n7 a_n1620_n2088# 0.270738f
C340 plus.t0 a_n1620_n2088# 0.638897f
C341 plus.n8 a_n1620_n2088# 0.296344f
C342 plus.n9 a_n1620_n2088# 0.010413f
C343 plus.n10 a_n1620_n2088# 0.291881f
C344 plus.n11 a_n1620_n2088# 1.14653f
.ends

