* NGSPICE file created from diffpair627.ext - technology: sky130A

.subckt diffpair627 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t21 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 source.t7 minus.t0 drain_right.t15 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X2 source.t26 plus.t1 drain_left.t14 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t18 plus.t2 drain_left.t13 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 drain_right.t14 minus.t1 source.t8 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X5 source.t25 plus.t3 drain_left.t12 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 source.t10 minus.t2 drain_right.t13 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 source.t6 minus.t3 drain_right.t12 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X8 a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X9 source.t27 plus.t4 drain_left.t11 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X10 source.t16 plus.t5 drain_left.t10 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X11 source.t24 plus.t6 drain_left.t9 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X12 drain_left.t8 plus.t7 source.t20 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X13 a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X14 drain_right.t11 minus.t4 source.t15 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X15 source.t2 minus.t5 drain_right.t10 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X16 drain_right.t9 minus.t6 source.t1 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X17 drain_right.t8 minus.t7 source.t3 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X18 drain_left.t7 plus.t8 source.t19 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X19 drain_right.t7 minus.t8 source.t4 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X20 drain_left.t6 plus.t9 source.t17 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X21 a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X22 drain_left.t5 plus.t10 source.t28 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 source.t23 plus.t11 drain_left.t4 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X24 drain_left.t3 plus.t12 source.t31 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X25 drain_right.t6 minus.t9 source.t9 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X26 drain_left.t2 plus.t13 source.t30 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X27 drain_right.t5 minus.t10 source.t11 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X28 drain_left.t1 plus.t14 source.t29 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X29 source.t0 minus.t11 drain_right.t4 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X30 a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X31 drain_right.t3 minus.t12 source.t13 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X32 source.t12 minus.t13 drain_right.t2 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X33 source.t14 minus.t14 drain_right.t1 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X34 source.t5 minus.t15 drain_right.t0 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X35 source.t22 plus.t15 drain_left.t0 a_n2570_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n7 plus.t5 769.066
R1 plus.n33 plus.t0 769.066
R2 plus.n24 plus.t8 744.691
R3 plus.n22 plus.t2 744.691
R4 plus.n2 plus.t10 744.691
R5 plus.n16 plus.t4 744.691
R6 plus.n4 plus.t9 744.691
R7 plus.n10 plus.t3 744.691
R8 plus.n6 plus.t13 744.691
R9 plus.n50 plus.t15 744.691
R10 plus.n48 plus.t7 744.691
R11 plus.n28 plus.t6 744.691
R12 plus.n42 plus.t12 744.691
R13 plus.n30 plus.t11 744.691
R14 plus.n36 plus.t14 744.691
R15 plus.n32 plus.t1 744.691
R16 plus.n9 plus.n8 161.3
R17 plus.n10 plus.n5 161.3
R18 plus.n12 plus.n11 161.3
R19 plus.n13 plus.n4 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n16 plus.n3 161.3
R22 plus.n18 plus.n17 161.3
R23 plus.n19 plus.n2 161.3
R24 plus.n21 plus.n20 161.3
R25 plus.n22 plus.n1 161.3
R26 plus.n23 plus.n0 161.3
R27 plus.n25 plus.n24 161.3
R28 plus.n35 plus.n34 161.3
R29 plus.n36 plus.n31 161.3
R30 plus.n38 plus.n37 161.3
R31 plus.n39 plus.n30 161.3
R32 plus.n41 plus.n40 161.3
R33 plus.n42 plus.n29 161.3
R34 plus.n44 plus.n43 161.3
R35 plus.n45 plus.n28 161.3
R36 plus.n47 plus.n46 161.3
R37 plus.n48 plus.n27 161.3
R38 plus.n49 plus.n26 161.3
R39 plus.n51 plus.n50 161.3
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus plus.n51 35.9233
R45 plus.n22 plus.n21 32.8641
R46 plus.n9 plus.n6 32.8641
R47 plus.n48 plus.n47 32.8641
R48 plus.n35 plus.n32 32.8641
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus plus.n25 15.33
R68 plus.n23 plus.n22 10.955
R69 plus.n49 plus.n48 10.955
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n0 source.t19 44.1297
R93 source.n7 source.t16 44.1296
R94 source.n8 source.t9 44.1296
R95 source.n15 source.t0 44.1296
R96 source.n31 source.t11 44.1295
R97 source.n24 source.t2 44.1295
R98 source.n23 source.t21 44.1295
R99 source.n16 source.t22 44.1295
R100 source.n2 source.n1 43.1397
R101 source.n4 source.n3 43.1397
R102 source.n6 source.n5 43.1397
R103 source.n10 source.n9 43.1397
R104 source.n12 source.n11 43.1397
R105 source.n14 source.n13 43.1397
R106 source.n30 source.n29 43.1396
R107 source.n28 source.n27 43.1396
R108 source.n26 source.n25 43.1396
R109 source.n22 source.n21 43.1396
R110 source.n20 source.n19 43.1396
R111 source.n18 source.n17 43.1396
R112 source.n16 source.n15 28.2363
R113 source.n32 source.n0 22.5294
R114 source.n32 source.n31 5.7074
R115 source.n29 source.t13 0.9905
R116 source.n29 source.t5 0.9905
R117 source.n27 source.t8 0.9905
R118 source.n27 source.t6 0.9905
R119 source.n25 source.t15 0.9905
R120 source.n25 source.t7 0.9905
R121 source.n21 source.t29 0.9905
R122 source.n21 source.t26 0.9905
R123 source.n19 source.t31 0.9905
R124 source.n19 source.t23 0.9905
R125 source.n17 source.t20 0.9905
R126 source.n17 source.t24 0.9905
R127 source.n1 source.t28 0.9905
R128 source.n1 source.t18 0.9905
R129 source.n3 source.t17 0.9905
R130 source.n3 source.t27 0.9905
R131 source.n5 source.t30 0.9905
R132 source.n5 source.t25 0.9905
R133 source.n9 source.t4 0.9905
R134 source.n9 source.t10 0.9905
R135 source.n11 source.t3 0.9905
R136 source.n11 source.t12 0.9905
R137 source.n13 source.t1 0.9905
R138 source.n13 source.t14 0.9905
R139 source.n15 source.n14 0.888431
R140 source.n14 source.n12 0.888431
R141 source.n12 source.n10 0.888431
R142 source.n10 source.n8 0.888431
R143 source.n7 source.n6 0.888431
R144 source.n6 source.n4 0.888431
R145 source.n4 source.n2 0.888431
R146 source.n2 source.n0 0.888431
R147 source.n18 source.n16 0.888431
R148 source.n20 source.n18 0.888431
R149 source.n22 source.n20 0.888431
R150 source.n23 source.n22 0.888431
R151 source.n26 source.n24 0.888431
R152 source.n28 source.n26 0.888431
R153 source.n30 source.n28 0.888431
R154 source.n31 source.n30 0.888431
R155 source.n8 source.n7 0.470328
R156 source.n24 source.n23 0.470328
R157 source source.n32 0.188
R158 drain_left.n9 drain_left.n7 60.7064
R159 drain_left.n5 drain_left.n3 60.7063
R160 drain_left.n2 drain_left.n0 60.7063
R161 drain_left.n13 drain_left.n12 59.8185
R162 drain_left.n11 drain_left.n10 59.8185
R163 drain_left.n9 drain_left.n8 59.8185
R164 drain_left.n5 drain_left.n4 59.8184
R165 drain_left.n2 drain_left.n1 59.8184
R166 drain_left drain_left.n6 39.1992
R167 drain_left drain_left.n13 6.54115
R168 drain_left.n3 drain_left.t14 0.9905
R169 drain_left.n3 drain_left.t15 0.9905
R170 drain_left.n4 drain_left.t4 0.9905
R171 drain_left.n4 drain_left.t1 0.9905
R172 drain_left.n1 drain_left.t9 0.9905
R173 drain_left.n1 drain_left.t3 0.9905
R174 drain_left.n0 drain_left.t0 0.9905
R175 drain_left.n0 drain_left.t8 0.9905
R176 drain_left.n12 drain_left.t13 0.9905
R177 drain_left.n12 drain_left.t7 0.9905
R178 drain_left.n10 drain_left.t11 0.9905
R179 drain_left.n10 drain_left.t5 0.9905
R180 drain_left.n8 drain_left.t12 0.9905
R181 drain_left.n8 drain_left.t6 0.9905
R182 drain_left.n7 drain_left.t10 0.9905
R183 drain_left.n7 drain_left.t2 0.9905
R184 drain_left.n11 drain_left.n9 0.888431
R185 drain_left.n13 drain_left.n11 0.888431
R186 drain_left.n6 drain_left.n5 0.389119
R187 drain_left.n6 drain_left.n2 0.389119
R188 minus.n7 minus.t9 769.066
R189 minus.n33 minus.t5 769.066
R190 minus.n6 minus.t2 744.691
R191 minus.n10 minus.t8 744.691
R192 minus.n12 minus.t13 744.691
R193 minus.n16 minus.t7 744.691
R194 minus.n18 minus.t14 744.691
R195 minus.n22 minus.t6 744.691
R196 minus.n24 minus.t11 744.691
R197 minus.n32 minus.t4 744.691
R198 minus.n36 minus.t0 744.691
R199 minus.n38 minus.t1 744.691
R200 minus.n42 minus.t3 744.691
R201 minus.n44 minus.t12 744.691
R202 minus.n48 minus.t15 744.691
R203 minus.n50 minus.t10 744.691
R204 minus.n25 minus.n24 161.3
R205 minus.n23 minus.n0 161.3
R206 minus.n22 minus.n21 161.3
R207 minus.n20 minus.n1 161.3
R208 minus.n19 minus.n18 161.3
R209 minus.n17 minus.n2 161.3
R210 minus.n16 minus.n15 161.3
R211 minus.n14 minus.n3 161.3
R212 minus.n13 minus.n12 161.3
R213 minus.n11 minus.n4 161.3
R214 minus.n10 minus.n9 161.3
R215 minus.n8 minus.n5 161.3
R216 minus.n51 minus.n50 161.3
R217 minus.n49 minus.n26 161.3
R218 minus.n48 minus.n47 161.3
R219 minus.n46 minus.n27 161.3
R220 minus.n45 minus.n44 161.3
R221 minus.n43 minus.n28 161.3
R222 minus.n42 minus.n41 161.3
R223 minus.n40 minus.n29 161.3
R224 minus.n39 minus.n38 161.3
R225 minus.n37 minus.n30 161.3
R226 minus.n36 minus.n35 161.3
R227 minus.n34 minus.n31 161.3
R228 minus.n52 minus.n25 45.0725
R229 minus.n8 minus.n7 44.9377
R230 minus.n34 minus.n33 44.9377
R231 minus.n24 minus.n23 37.246
R232 minus.n50 minus.n49 37.246
R233 minus.n6 minus.n5 32.8641
R234 minus.n22 minus.n1 32.8641
R235 minus.n32 minus.n31 32.8641
R236 minus.n48 minus.n27 32.8641
R237 minus.n11 minus.n10 28.4823
R238 minus.n18 minus.n17 28.4823
R239 minus.n37 minus.n36 28.4823
R240 minus.n44 minus.n43 28.4823
R241 minus.n16 minus.n3 24.1005
R242 minus.n12 minus.n3 24.1005
R243 minus.n38 minus.n29 24.1005
R244 minus.n42 minus.n29 24.1005
R245 minus.n12 minus.n11 19.7187
R246 minus.n17 minus.n16 19.7187
R247 minus.n38 minus.n37 19.7187
R248 minus.n43 minus.n42 19.7187
R249 minus.n7 minus.n6 17.0522
R250 minus.n33 minus.n32 17.0522
R251 minus.n10 minus.n5 15.3369
R252 minus.n18 minus.n1 15.3369
R253 minus.n36 minus.n31 15.3369
R254 minus.n44 minus.n27 15.3369
R255 minus.n23 minus.n22 10.955
R256 minus.n49 minus.n48 10.955
R257 minus.n52 minus.n51 6.6558
R258 minus.n25 minus.n0 0.189894
R259 minus.n21 minus.n0 0.189894
R260 minus.n21 minus.n20 0.189894
R261 minus.n20 minus.n19 0.189894
R262 minus.n19 minus.n2 0.189894
R263 minus.n15 minus.n2 0.189894
R264 minus.n15 minus.n14 0.189894
R265 minus.n14 minus.n13 0.189894
R266 minus.n13 minus.n4 0.189894
R267 minus.n9 minus.n4 0.189894
R268 minus.n9 minus.n8 0.189894
R269 minus.n35 minus.n34 0.189894
R270 minus.n35 minus.n30 0.189894
R271 minus.n39 minus.n30 0.189894
R272 minus.n40 minus.n39 0.189894
R273 minus.n41 minus.n40 0.189894
R274 minus.n41 minus.n28 0.189894
R275 minus.n45 minus.n28 0.189894
R276 minus.n46 minus.n45 0.189894
R277 minus.n47 minus.n46 0.189894
R278 minus.n47 minus.n26 0.189894
R279 minus.n51 minus.n26 0.189894
R280 minus minus.n52 0.188
R281 drain_right.n9 drain_right.n7 60.7064
R282 drain_right.n5 drain_right.n3 60.7063
R283 drain_right.n2 drain_right.n0 60.7063
R284 drain_right.n9 drain_right.n8 59.8185
R285 drain_right.n11 drain_right.n10 59.8185
R286 drain_right.n13 drain_right.n12 59.8185
R287 drain_right.n5 drain_right.n4 59.8184
R288 drain_right.n2 drain_right.n1 59.8184
R289 drain_right drain_right.n6 38.646
R290 drain_right drain_right.n13 6.54115
R291 drain_right.n3 drain_right.t0 0.9905
R292 drain_right.n3 drain_right.t5 0.9905
R293 drain_right.n4 drain_right.t12 0.9905
R294 drain_right.n4 drain_right.t3 0.9905
R295 drain_right.n1 drain_right.t15 0.9905
R296 drain_right.n1 drain_right.t14 0.9905
R297 drain_right.n0 drain_right.t10 0.9905
R298 drain_right.n0 drain_right.t11 0.9905
R299 drain_right.n7 drain_right.t13 0.9905
R300 drain_right.n7 drain_right.t6 0.9905
R301 drain_right.n8 drain_right.t2 0.9905
R302 drain_right.n8 drain_right.t7 0.9905
R303 drain_right.n10 drain_right.t1 0.9905
R304 drain_right.n10 drain_right.t8 0.9905
R305 drain_right.n12 drain_right.t4 0.9905
R306 drain_right.n12 drain_right.t9 0.9905
R307 drain_right.n13 drain_right.n11 0.888431
R308 drain_right.n11 drain_right.n9 0.888431
R309 drain_right.n6 drain_right.n5 0.389119
R310 drain_right.n6 drain_right.n2 0.389119
C0 source minus 16.3872f
C1 source plus 16.4012f
C2 minus plus 7.83164f
C3 drain_left drain_right 1.34352f
C4 source drain_right 30.6804f
C5 source drain_left 30.678198f
C6 minus drain_right 16.6724f
C7 drain_right plus 0.410755f
C8 minus drain_left 0.172697f
C9 drain_left plus 16.927f
C10 drain_right a_n2570_n4888# 8.24999f
C11 drain_left a_n2570_n4888# 8.608211f
C12 source a_n2570_n4888# 13.749782f
C13 minus a_n2570_n4888# 10.794901f
C14 plus a_n2570_n4888# 12.93996f
C15 drain_right.t10 a_n2570_n4888# 0.430645f
C16 drain_right.t11 a_n2570_n4888# 0.430645f
C17 drain_right.n0 a_n2570_n4888# 3.94286f
C18 drain_right.t15 a_n2570_n4888# 0.430645f
C19 drain_right.t14 a_n2570_n4888# 0.430645f
C20 drain_right.n1 a_n2570_n4888# 3.93705f
C21 drain_right.n2 a_n2570_n4888# 0.734666f
C22 drain_right.t0 a_n2570_n4888# 0.430645f
C23 drain_right.t5 a_n2570_n4888# 0.430645f
C24 drain_right.n3 a_n2570_n4888# 3.94286f
C25 drain_right.t12 a_n2570_n4888# 0.430645f
C26 drain_right.t3 a_n2570_n4888# 0.430645f
C27 drain_right.n4 a_n2570_n4888# 3.93705f
C28 drain_right.n5 a_n2570_n4888# 0.734666f
C29 drain_right.n6 a_n2570_n4888# 2.04397f
C30 drain_right.t13 a_n2570_n4888# 0.430645f
C31 drain_right.t6 a_n2570_n4888# 0.430645f
C32 drain_right.n7 a_n2570_n4888# 3.94285f
C33 drain_right.t2 a_n2570_n4888# 0.430645f
C34 drain_right.t7 a_n2570_n4888# 0.430645f
C35 drain_right.n8 a_n2570_n4888# 3.93705f
C36 drain_right.n9 a_n2570_n4888# 0.776891f
C37 drain_right.t1 a_n2570_n4888# 0.430645f
C38 drain_right.t8 a_n2570_n4888# 0.430645f
C39 drain_right.n10 a_n2570_n4888# 3.93705f
C40 drain_right.n11 a_n2570_n4888# 0.38586f
C41 drain_right.t4 a_n2570_n4888# 0.430645f
C42 drain_right.t9 a_n2570_n4888# 0.430645f
C43 drain_right.n12 a_n2570_n4888# 3.93705f
C44 drain_right.n13 a_n2570_n4888# 0.626871f
C45 minus.n0 a_n2570_n4888# 0.040203f
C46 minus.n1 a_n2570_n4888# 0.009123f
C47 minus.t6 a_n2570_n4888# 1.59391f
C48 minus.n2 a_n2570_n4888# 0.040203f
C49 minus.n3 a_n2570_n4888# 0.009123f
C50 minus.t7 a_n2570_n4888# 1.59391f
C51 minus.n4 a_n2570_n4888# 0.040203f
C52 minus.n5 a_n2570_n4888# 0.009123f
C53 minus.t8 a_n2570_n4888# 1.59391f
C54 minus.t9 a_n2570_n4888# 1.61275f
C55 minus.t2 a_n2570_n4888# 1.59391f
C56 minus.n6 a_n2570_n4888# 0.599872f
C57 minus.n7 a_n2570_n4888# 0.578867f
C58 minus.n8 a_n2570_n4888# 0.17013f
C59 minus.n9 a_n2570_n4888# 0.040203f
C60 minus.n10 a_n2570_n4888# 0.594364f
C61 minus.n11 a_n2570_n4888# 0.009123f
C62 minus.t13 a_n2570_n4888# 1.59391f
C63 minus.n12 a_n2570_n4888# 0.594364f
C64 minus.n13 a_n2570_n4888# 0.040203f
C65 minus.n14 a_n2570_n4888# 0.040203f
C66 minus.n15 a_n2570_n4888# 0.040203f
C67 minus.n16 a_n2570_n4888# 0.594364f
C68 minus.n17 a_n2570_n4888# 0.009123f
C69 minus.t14 a_n2570_n4888# 1.59391f
C70 minus.n18 a_n2570_n4888# 0.594364f
C71 minus.n19 a_n2570_n4888# 0.040203f
C72 minus.n20 a_n2570_n4888# 0.040203f
C73 minus.n21 a_n2570_n4888# 0.040203f
C74 minus.n22 a_n2570_n4888# 0.594364f
C75 minus.n23 a_n2570_n4888# 0.009123f
C76 minus.t11 a_n2570_n4888# 1.59391f
C77 minus.n24 a_n2570_n4888# 0.593249f
C78 minus.n25 a_n2570_n4888# 1.97675f
C79 minus.n26 a_n2570_n4888# 0.040203f
C80 minus.n27 a_n2570_n4888# 0.009123f
C81 minus.n28 a_n2570_n4888# 0.040203f
C82 minus.n29 a_n2570_n4888# 0.009123f
C83 minus.n30 a_n2570_n4888# 0.040203f
C84 minus.n31 a_n2570_n4888# 0.009123f
C85 minus.t5 a_n2570_n4888# 1.61275f
C86 minus.t4 a_n2570_n4888# 1.59391f
C87 minus.n32 a_n2570_n4888# 0.599872f
C88 minus.n33 a_n2570_n4888# 0.578867f
C89 minus.n34 a_n2570_n4888# 0.17013f
C90 minus.n35 a_n2570_n4888# 0.040203f
C91 minus.t0 a_n2570_n4888# 1.59391f
C92 minus.n36 a_n2570_n4888# 0.594364f
C93 minus.n37 a_n2570_n4888# 0.009123f
C94 minus.t1 a_n2570_n4888# 1.59391f
C95 minus.n38 a_n2570_n4888# 0.594364f
C96 minus.n39 a_n2570_n4888# 0.040203f
C97 minus.n40 a_n2570_n4888# 0.040203f
C98 minus.n41 a_n2570_n4888# 0.040203f
C99 minus.t3 a_n2570_n4888# 1.59391f
C100 minus.n42 a_n2570_n4888# 0.594364f
C101 minus.n43 a_n2570_n4888# 0.009123f
C102 minus.t12 a_n2570_n4888# 1.59391f
C103 minus.n44 a_n2570_n4888# 0.594364f
C104 minus.n45 a_n2570_n4888# 0.040203f
C105 minus.n46 a_n2570_n4888# 0.040203f
C106 minus.n47 a_n2570_n4888# 0.040203f
C107 minus.t15 a_n2570_n4888# 1.59391f
C108 minus.n48 a_n2570_n4888# 0.594364f
C109 minus.n49 a_n2570_n4888# 0.009123f
C110 minus.t10 a_n2570_n4888# 1.59391f
C111 minus.n50 a_n2570_n4888# 0.593249f
C112 minus.n51 a_n2570_n4888# 0.277487f
C113 minus.n52 a_n2570_n4888# 2.33769f
C114 drain_left.t0 a_n2570_n4888# 0.431492f
C115 drain_left.t8 a_n2570_n4888# 0.431492f
C116 drain_left.n0 a_n2570_n4888# 3.95061f
C117 drain_left.t9 a_n2570_n4888# 0.431492f
C118 drain_left.t3 a_n2570_n4888# 0.431492f
C119 drain_left.n1 a_n2570_n4888# 3.94479f
C120 drain_left.n2 a_n2570_n4888# 0.73611f
C121 drain_left.t14 a_n2570_n4888# 0.431492f
C122 drain_left.t15 a_n2570_n4888# 0.431492f
C123 drain_left.n3 a_n2570_n4888# 3.95061f
C124 drain_left.t4 a_n2570_n4888# 0.431492f
C125 drain_left.t1 a_n2570_n4888# 0.431492f
C126 drain_left.n4 a_n2570_n4888# 3.94479f
C127 drain_left.n5 a_n2570_n4888# 0.73611f
C128 drain_left.n6 a_n2570_n4888# 2.10424f
C129 drain_left.t10 a_n2570_n4888# 0.431492f
C130 drain_left.t2 a_n2570_n4888# 0.431492f
C131 drain_left.n7 a_n2570_n4888# 3.95061f
C132 drain_left.t12 a_n2570_n4888# 0.431492f
C133 drain_left.t6 a_n2570_n4888# 0.431492f
C134 drain_left.n8 a_n2570_n4888# 3.94479f
C135 drain_left.n9 a_n2570_n4888# 0.778418f
C136 drain_left.t11 a_n2570_n4888# 0.431492f
C137 drain_left.t5 a_n2570_n4888# 0.431492f
C138 drain_left.n10 a_n2570_n4888# 3.94479f
C139 drain_left.n11 a_n2570_n4888# 0.386619f
C140 drain_left.t13 a_n2570_n4888# 0.431492f
C141 drain_left.t7 a_n2570_n4888# 0.431492f
C142 drain_left.n12 a_n2570_n4888# 3.94479f
C143 drain_left.n13 a_n2570_n4888# 0.628104f
C144 source.t19 a_n2570_n4888# 4.07539f
C145 source.n0 a_n2570_n4888# 1.77291f
C146 source.t28 a_n2570_n4888# 0.356603f
C147 source.t18 a_n2570_n4888# 0.356603f
C148 source.n1 a_n2570_n4888# 3.18818f
C149 source.n2 a_n2570_n4888# 0.360805f
C150 source.t17 a_n2570_n4888# 0.356603f
C151 source.t27 a_n2570_n4888# 0.356603f
C152 source.n3 a_n2570_n4888# 3.18818f
C153 source.n4 a_n2570_n4888# 0.360805f
C154 source.t30 a_n2570_n4888# 0.356603f
C155 source.t25 a_n2570_n4888# 0.356603f
C156 source.n5 a_n2570_n4888# 3.18818f
C157 source.n6 a_n2570_n4888# 0.360805f
C158 source.t16 a_n2570_n4888# 4.0754f
C159 source.n7 a_n2570_n4888# 0.415741f
C160 source.t9 a_n2570_n4888# 4.0754f
C161 source.n8 a_n2570_n4888# 0.415741f
C162 source.t4 a_n2570_n4888# 0.356603f
C163 source.t10 a_n2570_n4888# 0.356603f
C164 source.n9 a_n2570_n4888# 3.18818f
C165 source.n10 a_n2570_n4888# 0.360805f
C166 source.t3 a_n2570_n4888# 0.356603f
C167 source.t12 a_n2570_n4888# 0.356603f
C168 source.n11 a_n2570_n4888# 3.18818f
C169 source.n12 a_n2570_n4888# 0.360805f
C170 source.t1 a_n2570_n4888# 0.356603f
C171 source.t14 a_n2570_n4888# 0.356603f
C172 source.n13 a_n2570_n4888# 3.18818f
C173 source.n14 a_n2570_n4888# 0.360805f
C174 source.t0 a_n2570_n4888# 4.0754f
C175 source.n15 a_n2570_n4888# 2.18339f
C176 source.t22 a_n2570_n4888# 4.07538f
C177 source.n16 a_n2570_n4888# 2.18341f
C178 source.t20 a_n2570_n4888# 0.356603f
C179 source.t24 a_n2570_n4888# 0.356603f
C180 source.n17 a_n2570_n4888# 3.18819f
C181 source.n18 a_n2570_n4888# 0.360798f
C182 source.t31 a_n2570_n4888# 0.356603f
C183 source.t23 a_n2570_n4888# 0.356603f
C184 source.n19 a_n2570_n4888# 3.18819f
C185 source.n20 a_n2570_n4888# 0.360798f
C186 source.t29 a_n2570_n4888# 0.356603f
C187 source.t26 a_n2570_n4888# 0.356603f
C188 source.n21 a_n2570_n4888# 3.18819f
C189 source.n22 a_n2570_n4888# 0.360798f
C190 source.t21 a_n2570_n4888# 4.07538f
C191 source.n23 a_n2570_n4888# 0.415763f
C192 source.t2 a_n2570_n4888# 4.07538f
C193 source.n24 a_n2570_n4888# 0.415763f
C194 source.t15 a_n2570_n4888# 0.356603f
C195 source.t7 a_n2570_n4888# 0.356603f
C196 source.n25 a_n2570_n4888# 3.18819f
C197 source.n26 a_n2570_n4888# 0.360798f
C198 source.t8 a_n2570_n4888# 0.356603f
C199 source.t6 a_n2570_n4888# 0.356603f
C200 source.n27 a_n2570_n4888# 3.18819f
C201 source.n28 a_n2570_n4888# 0.360798f
C202 source.t13 a_n2570_n4888# 0.356603f
C203 source.t5 a_n2570_n4888# 0.356603f
C204 source.n29 a_n2570_n4888# 3.18819f
C205 source.n30 a_n2570_n4888# 0.360798f
C206 source.t11 a_n2570_n4888# 4.07538f
C207 source.n31 a_n2570_n4888# 0.562944f
C208 source.n32 a_n2570_n4888# 2.047f
C209 plus.n0 a_n2570_n4888# 0.04048f
C210 plus.t8 a_n2570_n4888# 1.60489f
C211 plus.t2 a_n2570_n4888# 1.60489f
C212 plus.n1 a_n2570_n4888# 0.04048f
C213 plus.t10 a_n2570_n4888# 1.60489f
C214 plus.n2 a_n2570_n4888# 0.59846f
C215 plus.n3 a_n2570_n4888# 0.04048f
C216 plus.t4 a_n2570_n4888# 1.60489f
C217 plus.t9 a_n2570_n4888# 1.60489f
C218 plus.n4 a_n2570_n4888# 0.59846f
C219 plus.n5 a_n2570_n4888# 0.04048f
C220 plus.t3 a_n2570_n4888# 1.60489f
C221 plus.t13 a_n2570_n4888# 1.60489f
C222 plus.n6 a_n2570_n4888# 0.604006f
C223 plus.t5 a_n2570_n4888# 1.62387f
C224 plus.n7 a_n2570_n4888# 0.582856f
C225 plus.n8 a_n2570_n4888# 0.171302f
C226 plus.n9 a_n2570_n4888# 0.009186f
C227 plus.n10 a_n2570_n4888# 0.59846f
C228 plus.n11 a_n2570_n4888# 0.009186f
C229 plus.n12 a_n2570_n4888# 0.04048f
C230 plus.n13 a_n2570_n4888# 0.04048f
C231 plus.n14 a_n2570_n4888# 0.04048f
C232 plus.n15 a_n2570_n4888# 0.009186f
C233 plus.n16 a_n2570_n4888# 0.59846f
C234 plus.n17 a_n2570_n4888# 0.009186f
C235 plus.n18 a_n2570_n4888# 0.04048f
C236 plus.n19 a_n2570_n4888# 0.04048f
C237 plus.n20 a_n2570_n4888# 0.04048f
C238 plus.n21 a_n2570_n4888# 0.009186f
C239 plus.n22 a_n2570_n4888# 0.59846f
C240 plus.n23 a_n2570_n4888# 0.009186f
C241 plus.n24 a_n2570_n4888# 0.597337f
C242 plus.n25 a_n2570_n4888# 0.629127f
C243 plus.n26 a_n2570_n4888# 0.04048f
C244 plus.t15 a_n2570_n4888# 1.60489f
C245 plus.n27 a_n2570_n4888# 0.04048f
C246 plus.t7 a_n2570_n4888# 1.60489f
C247 plus.t6 a_n2570_n4888# 1.60489f
C248 plus.n28 a_n2570_n4888# 0.59846f
C249 plus.n29 a_n2570_n4888# 0.04048f
C250 plus.t12 a_n2570_n4888# 1.60489f
C251 plus.t11 a_n2570_n4888# 1.60489f
C252 plus.n30 a_n2570_n4888# 0.59846f
C253 plus.n31 a_n2570_n4888# 0.04048f
C254 plus.t14 a_n2570_n4888# 1.60489f
C255 plus.t1 a_n2570_n4888# 1.60489f
C256 plus.n32 a_n2570_n4888# 0.604006f
C257 plus.t0 a_n2570_n4888# 1.62387f
C258 plus.n33 a_n2570_n4888# 0.582856f
C259 plus.n34 a_n2570_n4888# 0.171302f
C260 plus.n35 a_n2570_n4888# 0.009186f
C261 plus.n36 a_n2570_n4888# 0.59846f
C262 plus.n37 a_n2570_n4888# 0.009186f
C263 plus.n38 a_n2570_n4888# 0.04048f
C264 plus.n39 a_n2570_n4888# 0.04048f
C265 plus.n40 a_n2570_n4888# 0.04048f
C266 plus.n41 a_n2570_n4888# 0.009186f
C267 plus.n42 a_n2570_n4888# 0.59846f
C268 plus.n43 a_n2570_n4888# 0.009186f
C269 plus.n44 a_n2570_n4888# 0.04048f
C270 plus.n45 a_n2570_n4888# 0.04048f
C271 plus.n46 a_n2570_n4888# 0.04048f
C272 plus.n47 a_n2570_n4888# 0.009186f
C273 plus.n48 a_n2570_n4888# 0.59846f
C274 plus.n49 a_n2570_n4888# 0.009186f
C275 plus.n50 a_n2570_n4888# 0.597337f
C276 plus.n51 a_n2570_n4888# 1.59402f
.ends

