* NGSPICE file created from diffpair293.ext - technology: sky130A

.subckt diffpair293 minus drain_right drain_left source plus
X0 a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.6
X1 source.t15 plus.t0 drain_left.t6 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X2 a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X3 source.t1 minus.t0 drain_right.t7 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X4 drain_left.t0 plus.t1 source.t14 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X5 source.t3 minus.t1 drain_right.t6 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X6 drain_right.t5 minus.t2 source.t0 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X7 drain_left.t3 plus.t2 source.t13 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X8 drain_right.t4 minus.t3 source.t7 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X9 source.t12 plus.t3 drain_left.t1 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X10 drain_left.t4 plus.t4 source.t11 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X11 source.t6 minus.t4 drain_right.t3 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X12 source.t10 plus.t5 drain_left.t2 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X13 drain_right.t2 minus.t5 source.t5 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X14 a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X15 drain_left.t7 plus.t6 source.t9 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X16 source.t8 plus.t7 drain_left.t5 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X17 drain_right.t1 minus.t6 source.t2 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X18 a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X19 source.t4 minus.t7 drain_right.t0 a_n1646_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
R0 plus.n1 plus.t7 333.293
R1 plus.n7 plus.t2 333.293
R2 plus.n4 plus.t4 306.473
R3 plus.n3 plus.t5 306.473
R4 plus.n2 plus.t6 306.473
R5 plus.n10 plus.t3 306.473
R6 plus.n9 plus.t1 306.473
R7 plus.n8 plus.t0 306.473
R8 plus.n5 plus.n4 161.3
R9 plus.n11 plus.n10 161.3
R10 plus.n3 plus.n0 80.6037
R11 plus.n9 plus.n6 80.6037
R12 plus.n4 plus.n3 48.2005
R13 plus.n3 plus.n2 48.2005
R14 plus.n10 plus.n9 48.2005
R15 plus.n9 plus.n8 48.2005
R16 plus.n1 plus.n0 45.2318
R17 plus.n7 plus.n6 45.2318
R18 plus plus.n11 27.0786
R19 plus.n2 plus.n1 13.3799
R20 plus.n8 plus.n7 13.3799
R21 plus plus.n5 9.98535
R22 plus.n5 plus.n0 0.285035
R23 plus.n11 plus.n6 0.285035
R24 drain_left.n5 drain_left.n3 67.9925
R25 drain_left.n2 drain_left.n1 67.5362
R26 drain_left.n2 drain_left.n0 67.5362
R27 drain_left.n5 drain_left.n4 67.1907
R28 drain_left drain_left.n2 25.6277
R29 drain_left drain_left.n5 6.45494
R30 drain_left.n1 drain_left.t6 3.3005
R31 drain_left.n1 drain_left.t3 3.3005
R32 drain_left.n0 drain_left.t1 3.3005
R33 drain_left.n0 drain_left.t0 3.3005
R34 drain_left.n4 drain_left.t2 3.3005
R35 drain_left.n4 drain_left.t4 3.3005
R36 drain_left.n3 drain_left.t5 3.3005
R37 drain_left.n3 drain_left.t7 3.3005
R38 source.n258 source.n232 289.615
R39 source.n224 source.n198 289.615
R40 source.n192 source.n166 289.615
R41 source.n158 source.n132 289.615
R42 source.n26 source.n0 289.615
R43 source.n60 source.n34 289.615
R44 source.n92 source.n66 289.615
R45 source.n126 source.n100 289.615
R46 source.n243 source.n242 185
R47 source.n240 source.n239 185
R48 source.n249 source.n248 185
R49 source.n251 source.n250 185
R50 source.n236 source.n235 185
R51 source.n257 source.n256 185
R52 source.n259 source.n258 185
R53 source.n209 source.n208 185
R54 source.n206 source.n205 185
R55 source.n215 source.n214 185
R56 source.n217 source.n216 185
R57 source.n202 source.n201 185
R58 source.n223 source.n222 185
R59 source.n225 source.n224 185
R60 source.n177 source.n176 185
R61 source.n174 source.n173 185
R62 source.n183 source.n182 185
R63 source.n185 source.n184 185
R64 source.n170 source.n169 185
R65 source.n191 source.n190 185
R66 source.n193 source.n192 185
R67 source.n143 source.n142 185
R68 source.n140 source.n139 185
R69 source.n149 source.n148 185
R70 source.n151 source.n150 185
R71 source.n136 source.n135 185
R72 source.n157 source.n156 185
R73 source.n159 source.n158 185
R74 source.n27 source.n26 185
R75 source.n25 source.n24 185
R76 source.n4 source.n3 185
R77 source.n19 source.n18 185
R78 source.n17 source.n16 185
R79 source.n8 source.n7 185
R80 source.n11 source.n10 185
R81 source.n61 source.n60 185
R82 source.n59 source.n58 185
R83 source.n38 source.n37 185
R84 source.n53 source.n52 185
R85 source.n51 source.n50 185
R86 source.n42 source.n41 185
R87 source.n45 source.n44 185
R88 source.n93 source.n92 185
R89 source.n91 source.n90 185
R90 source.n70 source.n69 185
R91 source.n85 source.n84 185
R92 source.n83 source.n82 185
R93 source.n74 source.n73 185
R94 source.n77 source.n76 185
R95 source.n127 source.n126 185
R96 source.n125 source.n124 185
R97 source.n104 source.n103 185
R98 source.n119 source.n118 185
R99 source.n117 source.n116 185
R100 source.n108 source.n107 185
R101 source.n111 source.n110 185
R102 source.t0 source.n241 147.661
R103 source.t1 source.n207 147.661
R104 source.t13 source.n175 147.661
R105 source.t12 source.n141 147.661
R106 source.t11 source.n9 147.661
R107 source.t8 source.n43 147.661
R108 source.t5 source.n75 147.661
R109 source.t3 source.n109 147.661
R110 source.n242 source.n239 104.615
R111 source.n249 source.n239 104.615
R112 source.n250 source.n249 104.615
R113 source.n250 source.n235 104.615
R114 source.n257 source.n235 104.615
R115 source.n258 source.n257 104.615
R116 source.n208 source.n205 104.615
R117 source.n215 source.n205 104.615
R118 source.n216 source.n215 104.615
R119 source.n216 source.n201 104.615
R120 source.n223 source.n201 104.615
R121 source.n224 source.n223 104.615
R122 source.n176 source.n173 104.615
R123 source.n183 source.n173 104.615
R124 source.n184 source.n183 104.615
R125 source.n184 source.n169 104.615
R126 source.n191 source.n169 104.615
R127 source.n192 source.n191 104.615
R128 source.n142 source.n139 104.615
R129 source.n149 source.n139 104.615
R130 source.n150 source.n149 104.615
R131 source.n150 source.n135 104.615
R132 source.n157 source.n135 104.615
R133 source.n158 source.n157 104.615
R134 source.n26 source.n25 104.615
R135 source.n25 source.n3 104.615
R136 source.n18 source.n3 104.615
R137 source.n18 source.n17 104.615
R138 source.n17 source.n7 104.615
R139 source.n10 source.n7 104.615
R140 source.n60 source.n59 104.615
R141 source.n59 source.n37 104.615
R142 source.n52 source.n37 104.615
R143 source.n52 source.n51 104.615
R144 source.n51 source.n41 104.615
R145 source.n44 source.n41 104.615
R146 source.n92 source.n91 104.615
R147 source.n91 source.n69 104.615
R148 source.n84 source.n69 104.615
R149 source.n84 source.n83 104.615
R150 source.n83 source.n73 104.615
R151 source.n76 source.n73 104.615
R152 source.n126 source.n125 104.615
R153 source.n125 source.n103 104.615
R154 source.n118 source.n103 104.615
R155 source.n118 source.n117 104.615
R156 source.n117 source.n107 104.615
R157 source.n110 source.n107 104.615
R158 source.n242 source.t0 52.3082
R159 source.n208 source.t1 52.3082
R160 source.n176 source.t13 52.3082
R161 source.n142 source.t12 52.3082
R162 source.n10 source.t11 52.3082
R163 source.n44 source.t8 52.3082
R164 source.n76 source.t5 52.3082
R165 source.n110 source.t3 52.3082
R166 source.n33 source.n32 50.512
R167 source.n99 source.n98 50.512
R168 source.n231 source.n230 50.5119
R169 source.n165 source.n164 50.5119
R170 source.n263 source.n262 32.1853
R171 source.n229 source.n228 32.1853
R172 source.n197 source.n196 32.1853
R173 source.n163 source.n162 32.1853
R174 source.n31 source.n30 32.1853
R175 source.n65 source.n64 32.1853
R176 source.n97 source.n96 32.1853
R177 source.n131 source.n130 32.1853
R178 source.n163 source.n131 17.544
R179 source.n243 source.n241 15.6674
R180 source.n209 source.n207 15.6674
R181 source.n177 source.n175 15.6674
R182 source.n143 source.n141 15.6674
R183 source.n11 source.n9 15.6674
R184 source.n45 source.n43 15.6674
R185 source.n77 source.n75 15.6674
R186 source.n111 source.n109 15.6674
R187 source.n244 source.n240 12.8005
R188 source.n210 source.n206 12.8005
R189 source.n178 source.n174 12.8005
R190 source.n144 source.n140 12.8005
R191 source.n12 source.n8 12.8005
R192 source.n46 source.n42 12.8005
R193 source.n78 source.n74 12.8005
R194 source.n112 source.n108 12.8005
R195 source.n248 source.n247 12.0247
R196 source.n214 source.n213 12.0247
R197 source.n182 source.n181 12.0247
R198 source.n148 source.n147 12.0247
R199 source.n16 source.n15 12.0247
R200 source.n50 source.n49 12.0247
R201 source.n82 source.n81 12.0247
R202 source.n116 source.n115 12.0247
R203 source.n264 source.n31 11.8802
R204 source.n251 source.n238 11.249
R205 source.n217 source.n204 11.249
R206 source.n185 source.n172 11.249
R207 source.n151 source.n138 11.249
R208 source.n19 source.n6 11.249
R209 source.n53 source.n40 11.249
R210 source.n85 source.n72 11.249
R211 source.n119 source.n106 11.249
R212 source.n252 source.n236 10.4732
R213 source.n218 source.n202 10.4732
R214 source.n186 source.n170 10.4732
R215 source.n152 source.n136 10.4732
R216 source.n20 source.n4 10.4732
R217 source.n54 source.n38 10.4732
R218 source.n86 source.n70 10.4732
R219 source.n120 source.n104 10.4732
R220 source.n256 source.n255 9.69747
R221 source.n222 source.n221 9.69747
R222 source.n190 source.n189 9.69747
R223 source.n156 source.n155 9.69747
R224 source.n24 source.n23 9.69747
R225 source.n58 source.n57 9.69747
R226 source.n90 source.n89 9.69747
R227 source.n124 source.n123 9.69747
R228 source.n262 source.n261 9.45567
R229 source.n228 source.n227 9.45567
R230 source.n196 source.n195 9.45567
R231 source.n162 source.n161 9.45567
R232 source.n30 source.n29 9.45567
R233 source.n64 source.n63 9.45567
R234 source.n96 source.n95 9.45567
R235 source.n130 source.n129 9.45567
R236 source.n261 source.n260 9.3005
R237 source.n234 source.n233 9.3005
R238 source.n255 source.n254 9.3005
R239 source.n253 source.n252 9.3005
R240 source.n238 source.n237 9.3005
R241 source.n247 source.n246 9.3005
R242 source.n245 source.n244 9.3005
R243 source.n227 source.n226 9.3005
R244 source.n200 source.n199 9.3005
R245 source.n221 source.n220 9.3005
R246 source.n219 source.n218 9.3005
R247 source.n204 source.n203 9.3005
R248 source.n213 source.n212 9.3005
R249 source.n211 source.n210 9.3005
R250 source.n195 source.n194 9.3005
R251 source.n168 source.n167 9.3005
R252 source.n189 source.n188 9.3005
R253 source.n187 source.n186 9.3005
R254 source.n172 source.n171 9.3005
R255 source.n181 source.n180 9.3005
R256 source.n179 source.n178 9.3005
R257 source.n161 source.n160 9.3005
R258 source.n134 source.n133 9.3005
R259 source.n155 source.n154 9.3005
R260 source.n153 source.n152 9.3005
R261 source.n138 source.n137 9.3005
R262 source.n147 source.n146 9.3005
R263 source.n145 source.n144 9.3005
R264 source.n29 source.n28 9.3005
R265 source.n2 source.n1 9.3005
R266 source.n23 source.n22 9.3005
R267 source.n21 source.n20 9.3005
R268 source.n6 source.n5 9.3005
R269 source.n15 source.n14 9.3005
R270 source.n13 source.n12 9.3005
R271 source.n63 source.n62 9.3005
R272 source.n36 source.n35 9.3005
R273 source.n57 source.n56 9.3005
R274 source.n55 source.n54 9.3005
R275 source.n40 source.n39 9.3005
R276 source.n49 source.n48 9.3005
R277 source.n47 source.n46 9.3005
R278 source.n95 source.n94 9.3005
R279 source.n68 source.n67 9.3005
R280 source.n89 source.n88 9.3005
R281 source.n87 source.n86 9.3005
R282 source.n72 source.n71 9.3005
R283 source.n81 source.n80 9.3005
R284 source.n79 source.n78 9.3005
R285 source.n129 source.n128 9.3005
R286 source.n102 source.n101 9.3005
R287 source.n123 source.n122 9.3005
R288 source.n121 source.n120 9.3005
R289 source.n106 source.n105 9.3005
R290 source.n115 source.n114 9.3005
R291 source.n113 source.n112 9.3005
R292 source.n259 source.n234 8.92171
R293 source.n225 source.n200 8.92171
R294 source.n193 source.n168 8.92171
R295 source.n159 source.n134 8.92171
R296 source.n27 source.n2 8.92171
R297 source.n61 source.n36 8.92171
R298 source.n93 source.n68 8.92171
R299 source.n127 source.n102 8.92171
R300 source.n260 source.n232 8.14595
R301 source.n226 source.n198 8.14595
R302 source.n194 source.n166 8.14595
R303 source.n160 source.n132 8.14595
R304 source.n28 source.n0 8.14595
R305 source.n62 source.n34 8.14595
R306 source.n94 source.n66 8.14595
R307 source.n128 source.n100 8.14595
R308 source.n262 source.n232 5.81868
R309 source.n228 source.n198 5.81868
R310 source.n196 source.n166 5.81868
R311 source.n162 source.n132 5.81868
R312 source.n30 source.n0 5.81868
R313 source.n64 source.n34 5.81868
R314 source.n96 source.n66 5.81868
R315 source.n130 source.n100 5.81868
R316 source.n264 source.n263 5.66429
R317 source.n260 source.n259 5.04292
R318 source.n226 source.n225 5.04292
R319 source.n194 source.n193 5.04292
R320 source.n160 source.n159 5.04292
R321 source.n28 source.n27 5.04292
R322 source.n62 source.n61 5.04292
R323 source.n94 source.n93 5.04292
R324 source.n128 source.n127 5.04292
R325 source.n245 source.n241 4.38594
R326 source.n211 source.n207 4.38594
R327 source.n179 source.n175 4.38594
R328 source.n145 source.n141 4.38594
R329 source.n13 source.n9 4.38594
R330 source.n47 source.n43 4.38594
R331 source.n79 source.n75 4.38594
R332 source.n113 source.n109 4.38594
R333 source.n256 source.n234 4.26717
R334 source.n222 source.n200 4.26717
R335 source.n190 source.n168 4.26717
R336 source.n156 source.n134 4.26717
R337 source.n24 source.n2 4.26717
R338 source.n58 source.n36 4.26717
R339 source.n90 source.n68 4.26717
R340 source.n124 source.n102 4.26717
R341 source.n255 source.n236 3.49141
R342 source.n221 source.n202 3.49141
R343 source.n189 source.n170 3.49141
R344 source.n155 source.n136 3.49141
R345 source.n23 source.n4 3.49141
R346 source.n57 source.n38 3.49141
R347 source.n89 source.n70 3.49141
R348 source.n123 source.n104 3.49141
R349 source.n230 source.t2 3.3005
R350 source.n230 source.t4 3.3005
R351 source.n164 source.t14 3.3005
R352 source.n164 source.t15 3.3005
R353 source.n32 source.t9 3.3005
R354 source.n32 source.t10 3.3005
R355 source.n98 source.t7 3.3005
R356 source.n98 source.t6 3.3005
R357 source.n252 source.n251 2.71565
R358 source.n218 source.n217 2.71565
R359 source.n186 source.n185 2.71565
R360 source.n152 source.n151 2.71565
R361 source.n20 source.n19 2.71565
R362 source.n54 source.n53 2.71565
R363 source.n86 source.n85 2.71565
R364 source.n120 source.n119 2.71565
R365 source.n248 source.n238 1.93989
R366 source.n214 source.n204 1.93989
R367 source.n182 source.n172 1.93989
R368 source.n148 source.n138 1.93989
R369 source.n16 source.n6 1.93989
R370 source.n50 source.n40 1.93989
R371 source.n82 source.n72 1.93989
R372 source.n116 source.n106 1.93989
R373 source.n247 source.n240 1.16414
R374 source.n213 source.n206 1.16414
R375 source.n181 source.n174 1.16414
R376 source.n147 source.n140 1.16414
R377 source.n15 source.n8 1.16414
R378 source.n49 source.n42 1.16414
R379 source.n81 source.n74 1.16414
R380 source.n115 source.n108 1.16414
R381 source.n131 source.n99 0.802224
R382 source.n99 source.n97 0.802224
R383 source.n65 source.n33 0.802224
R384 source.n33 source.n31 0.802224
R385 source.n165 source.n163 0.802224
R386 source.n197 source.n165 0.802224
R387 source.n231 source.n229 0.802224
R388 source.n263 source.n231 0.802224
R389 source.n97 source.n65 0.470328
R390 source.n229 source.n197 0.470328
R391 source.n244 source.n243 0.388379
R392 source.n210 source.n209 0.388379
R393 source.n178 source.n177 0.388379
R394 source.n144 source.n143 0.388379
R395 source.n12 source.n11 0.388379
R396 source.n46 source.n45 0.388379
R397 source.n78 source.n77 0.388379
R398 source.n112 source.n111 0.388379
R399 source source.n264 0.188
R400 source.n246 source.n245 0.155672
R401 source.n246 source.n237 0.155672
R402 source.n253 source.n237 0.155672
R403 source.n254 source.n253 0.155672
R404 source.n254 source.n233 0.155672
R405 source.n261 source.n233 0.155672
R406 source.n212 source.n211 0.155672
R407 source.n212 source.n203 0.155672
R408 source.n219 source.n203 0.155672
R409 source.n220 source.n219 0.155672
R410 source.n220 source.n199 0.155672
R411 source.n227 source.n199 0.155672
R412 source.n180 source.n179 0.155672
R413 source.n180 source.n171 0.155672
R414 source.n187 source.n171 0.155672
R415 source.n188 source.n187 0.155672
R416 source.n188 source.n167 0.155672
R417 source.n195 source.n167 0.155672
R418 source.n146 source.n145 0.155672
R419 source.n146 source.n137 0.155672
R420 source.n153 source.n137 0.155672
R421 source.n154 source.n153 0.155672
R422 source.n154 source.n133 0.155672
R423 source.n161 source.n133 0.155672
R424 source.n29 source.n1 0.155672
R425 source.n22 source.n1 0.155672
R426 source.n22 source.n21 0.155672
R427 source.n21 source.n5 0.155672
R428 source.n14 source.n5 0.155672
R429 source.n14 source.n13 0.155672
R430 source.n63 source.n35 0.155672
R431 source.n56 source.n35 0.155672
R432 source.n56 source.n55 0.155672
R433 source.n55 source.n39 0.155672
R434 source.n48 source.n39 0.155672
R435 source.n48 source.n47 0.155672
R436 source.n95 source.n67 0.155672
R437 source.n88 source.n67 0.155672
R438 source.n88 source.n87 0.155672
R439 source.n87 source.n71 0.155672
R440 source.n80 source.n71 0.155672
R441 source.n80 source.n79 0.155672
R442 source.n129 source.n101 0.155672
R443 source.n122 source.n101 0.155672
R444 source.n122 source.n121 0.155672
R445 source.n121 source.n105 0.155672
R446 source.n114 source.n105 0.155672
R447 source.n114 source.n113 0.155672
R448 minus.n1 minus.t5 333.293
R449 minus.n7 minus.t0 333.293
R450 minus.n2 minus.t4 306.473
R451 minus.n3 minus.t3 306.473
R452 minus.n4 minus.t1 306.473
R453 minus.n8 minus.t6 306.473
R454 minus.n9 minus.t7 306.473
R455 minus.n10 minus.t2 306.473
R456 minus.n5 minus.n4 161.3
R457 minus.n11 minus.n10 161.3
R458 minus.n3 minus.n0 80.6037
R459 minus.n9 minus.n6 80.6037
R460 minus.n3 minus.n2 48.2005
R461 minus.n4 minus.n3 48.2005
R462 minus.n9 minus.n8 48.2005
R463 minus.n10 minus.n9 48.2005
R464 minus.n1 minus.n0 45.2318
R465 minus.n7 minus.n6 45.2318
R466 minus.n12 minus.n5 30.9247
R467 minus.n2 minus.n1 13.3799
R468 minus.n8 minus.n7 13.3799
R469 minus.n12 minus.n11 6.61414
R470 minus.n5 minus.n0 0.285035
R471 minus.n11 minus.n6 0.285035
R472 minus minus.n12 0.188
R473 drain_right.n5 drain_right.n3 67.9924
R474 drain_right.n2 drain_right.n1 67.5362
R475 drain_right.n2 drain_right.n0 67.5362
R476 drain_right.n5 drain_right.n4 67.1908
R477 drain_right drain_right.n2 25.0744
R478 drain_right drain_right.n5 6.45494
R479 drain_right.n1 drain_right.t0 3.3005
R480 drain_right.n1 drain_right.t5 3.3005
R481 drain_right.n0 drain_right.t7 3.3005
R482 drain_right.n0 drain_right.t1 3.3005
R483 drain_right.n3 drain_right.t3 3.3005
R484 drain_right.n3 drain_right.t2 3.3005
R485 drain_right.n4 drain_right.t6 3.3005
R486 drain_right.n4 drain_right.t4 3.3005
C0 drain_left drain_right 0.775958f
C1 plus drain_left 2.89013f
C2 drain_left source 7.05487f
C3 minus drain_left 0.171399f
C4 plus drain_right 0.312845f
C5 drain_right source 7.05602f
C6 plus source 2.75955f
C7 minus drain_right 2.73169f
C8 plus minus 4.08444f
C9 minus source 2.74553f
C10 drain_right a_n1646_n2088# 4.43201f
C11 drain_left a_n1646_n2088# 4.68944f
C12 source a_n1646_n2088# 5.353122f
C13 minus a_n1646_n2088# 5.880332f
C14 plus a_n1646_n2088# 7.31546f
C15 drain_right.t7 a_n1646_n2088# 0.129488f
C16 drain_right.t1 a_n1646_n2088# 0.129488f
C17 drain_right.n0 a_n1646_n2088# 1.08165f
C18 drain_right.t0 a_n1646_n2088# 0.129488f
C19 drain_right.t5 a_n1646_n2088# 0.129488f
C20 drain_right.n1 a_n1646_n2088# 1.08165f
C21 drain_right.n2 a_n1646_n2088# 1.55709f
C22 drain_right.t3 a_n1646_n2088# 0.129488f
C23 drain_right.t2 a_n1646_n2088# 0.129488f
C24 drain_right.n3 a_n1646_n2088# 1.08434f
C25 drain_right.t6 a_n1646_n2088# 0.129488f
C26 drain_right.t4 a_n1646_n2088# 0.129488f
C27 drain_right.n4 a_n1646_n2088# 1.07994f
C28 drain_right.n5 a_n1646_n2088# 0.970257f
C29 minus.n0 a_n1646_n2088# 0.228649f
C30 minus.t4 a_n1646_n2088# 0.48964f
C31 minus.t5 a_n1646_n2088# 0.50804f
C32 minus.n1 a_n1646_n2088# 0.211525f
C33 minus.n2 a_n1646_n2088# 0.239162f
C34 minus.t3 a_n1646_n2088# 0.48964f
C35 minus.n3 a_n1646_n2088# 0.239162f
C36 minus.t1 a_n1646_n2088# 0.48964f
C37 minus.n4 a_n1646_n2088# 0.228521f
C38 minus.n5 a_n1646_n2088# 1.30475f
C39 minus.n6 a_n1646_n2088# 0.228649f
C40 minus.t0 a_n1646_n2088# 0.50804f
C41 minus.n7 a_n1646_n2088# 0.211525f
C42 minus.t6 a_n1646_n2088# 0.48964f
C43 minus.n8 a_n1646_n2088# 0.239162f
C44 minus.t7 a_n1646_n2088# 0.48964f
C45 minus.n9 a_n1646_n2088# 0.239162f
C46 minus.t2 a_n1646_n2088# 0.48964f
C47 minus.n10 a_n1646_n2088# 0.228521f
C48 minus.n11 a_n1646_n2088# 0.334785f
C49 minus.n12 a_n1646_n2088# 1.58171f
C50 source.n0 a_n1646_n2088# 0.03118f
C51 source.n1 a_n1646_n2088# 0.022183f
C52 source.n2 a_n1646_n2088# 0.01192f
C53 source.n3 a_n1646_n2088# 0.028175f
C54 source.n4 a_n1646_n2088# 0.012621f
C55 source.n5 a_n1646_n2088# 0.022183f
C56 source.n6 a_n1646_n2088# 0.01192f
C57 source.n7 a_n1646_n2088# 0.028175f
C58 source.n8 a_n1646_n2088# 0.012621f
C59 source.n9 a_n1646_n2088# 0.094928f
C60 source.t11 a_n1646_n2088# 0.045922f
C61 source.n10 a_n1646_n2088# 0.021131f
C62 source.n11 a_n1646_n2088# 0.016643f
C63 source.n12 a_n1646_n2088# 0.01192f
C64 source.n13 a_n1646_n2088# 0.527823f
C65 source.n14 a_n1646_n2088# 0.022183f
C66 source.n15 a_n1646_n2088# 0.01192f
C67 source.n16 a_n1646_n2088# 0.012621f
C68 source.n17 a_n1646_n2088# 0.028175f
C69 source.n18 a_n1646_n2088# 0.028175f
C70 source.n19 a_n1646_n2088# 0.012621f
C71 source.n20 a_n1646_n2088# 0.01192f
C72 source.n21 a_n1646_n2088# 0.022183f
C73 source.n22 a_n1646_n2088# 0.022183f
C74 source.n23 a_n1646_n2088# 0.01192f
C75 source.n24 a_n1646_n2088# 0.012621f
C76 source.n25 a_n1646_n2088# 0.028175f
C77 source.n26 a_n1646_n2088# 0.060994f
C78 source.n27 a_n1646_n2088# 0.012621f
C79 source.n28 a_n1646_n2088# 0.01192f
C80 source.n29 a_n1646_n2088# 0.051275f
C81 source.n30 a_n1646_n2088# 0.034129f
C82 source.n31 a_n1646_n2088# 0.568968f
C83 source.t9 a_n1646_n2088# 0.105178f
C84 source.t10 a_n1646_n2088# 0.105178f
C85 source.n32 a_n1646_n2088# 0.819136f
C86 source.n33 a_n1646_n2088# 0.322557f
C87 source.n34 a_n1646_n2088# 0.03118f
C88 source.n35 a_n1646_n2088# 0.022183f
C89 source.n36 a_n1646_n2088# 0.01192f
C90 source.n37 a_n1646_n2088# 0.028175f
C91 source.n38 a_n1646_n2088# 0.012621f
C92 source.n39 a_n1646_n2088# 0.022183f
C93 source.n40 a_n1646_n2088# 0.01192f
C94 source.n41 a_n1646_n2088# 0.028175f
C95 source.n42 a_n1646_n2088# 0.012621f
C96 source.n43 a_n1646_n2088# 0.094928f
C97 source.t8 a_n1646_n2088# 0.045922f
C98 source.n44 a_n1646_n2088# 0.021131f
C99 source.n45 a_n1646_n2088# 0.016643f
C100 source.n46 a_n1646_n2088# 0.01192f
C101 source.n47 a_n1646_n2088# 0.527823f
C102 source.n48 a_n1646_n2088# 0.022183f
C103 source.n49 a_n1646_n2088# 0.01192f
C104 source.n50 a_n1646_n2088# 0.012621f
C105 source.n51 a_n1646_n2088# 0.028175f
C106 source.n52 a_n1646_n2088# 0.028175f
C107 source.n53 a_n1646_n2088# 0.012621f
C108 source.n54 a_n1646_n2088# 0.01192f
C109 source.n55 a_n1646_n2088# 0.022183f
C110 source.n56 a_n1646_n2088# 0.022183f
C111 source.n57 a_n1646_n2088# 0.01192f
C112 source.n58 a_n1646_n2088# 0.012621f
C113 source.n59 a_n1646_n2088# 0.028175f
C114 source.n60 a_n1646_n2088# 0.060994f
C115 source.n61 a_n1646_n2088# 0.012621f
C116 source.n62 a_n1646_n2088# 0.01192f
C117 source.n63 a_n1646_n2088# 0.051275f
C118 source.n64 a_n1646_n2088# 0.034129f
C119 source.n65 a_n1646_n2088# 0.109835f
C120 source.n66 a_n1646_n2088# 0.03118f
C121 source.n67 a_n1646_n2088# 0.022183f
C122 source.n68 a_n1646_n2088# 0.01192f
C123 source.n69 a_n1646_n2088# 0.028175f
C124 source.n70 a_n1646_n2088# 0.012621f
C125 source.n71 a_n1646_n2088# 0.022183f
C126 source.n72 a_n1646_n2088# 0.01192f
C127 source.n73 a_n1646_n2088# 0.028175f
C128 source.n74 a_n1646_n2088# 0.012621f
C129 source.n75 a_n1646_n2088# 0.094928f
C130 source.t5 a_n1646_n2088# 0.045922f
C131 source.n76 a_n1646_n2088# 0.021131f
C132 source.n77 a_n1646_n2088# 0.016643f
C133 source.n78 a_n1646_n2088# 0.01192f
C134 source.n79 a_n1646_n2088# 0.527823f
C135 source.n80 a_n1646_n2088# 0.022183f
C136 source.n81 a_n1646_n2088# 0.01192f
C137 source.n82 a_n1646_n2088# 0.012621f
C138 source.n83 a_n1646_n2088# 0.028175f
C139 source.n84 a_n1646_n2088# 0.028175f
C140 source.n85 a_n1646_n2088# 0.012621f
C141 source.n86 a_n1646_n2088# 0.01192f
C142 source.n87 a_n1646_n2088# 0.022183f
C143 source.n88 a_n1646_n2088# 0.022183f
C144 source.n89 a_n1646_n2088# 0.01192f
C145 source.n90 a_n1646_n2088# 0.012621f
C146 source.n91 a_n1646_n2088# 0.028175f
C147 source.n92 a_n1646_n2088# 0.060994f
C148 source.n93 a_n1646_n2088# 0.012621f
C149 source.n94 a_n1646_n2088# 0.01192f
C150 source.n95 a_n1646_n2088# 0.051275f
C151 source.n96 a_n1646_n2088# 0.034129f
C152 source.n97 a_n1646_n2088# 0.109835f
C153 source.t7 a_n1646_n2088# 0.105178f
C154 source.t6 a_n1646_n2088# 0.105178f
C155 source.n98 a_n1646_n2088# 0.819136f
C156 source.n99 a_n1646_n2088# 0.322557f
C157 source.n100 a_n1646_n2088# 0.03118f
C158 source.n101 a_n1646_n2088# 0.022183f
C159 source.n102 a_n1646_n2088# 0.01192f
C160 source.n103 a_n1646_n2088# 0.028175f
C161 source.n104 a_n1646_n2088# 0.012621f
C162 source.n105 a_n1646_n2088# 0.022183f
C163 source.n106 a_n1646_n2088# 0.01192f
C164 source.n107 a_n1646_n2088# 0.028175f
C165 source.n108 a_n1646_n2088# 0.012621f
C166 source.n109 a_n1646_n2088# 0.094928f
C167 source.t3 a_n1646_n2088# 0.045922f
C168 source.n110 a_n1646_n2088# 0.021131f
C169 source.n111 a_n1646_n2088# 0.016643f
C170 source.n112 a_n1646_n2088# 0.01192f
C171 source.n113 a_n1646_n2088# 0.527823f
C172 source.n114 a_n1646_n2088# 0.022183f
C173 source.n115 a_n1646_n2088# 0.01192f
C174 source.n116 a_n1646_n2088# 0.012621f
C175 source.n117 a_n1646_n2088# 0.028175f
C176 source.n118 a_n1646_n2088# 0.028175f
C177 source.n119 a_n1646_n2088# 0.012621f
C178 source.n120 a_n1646_n2088# 0.01192f
C179 source.n121 a_n1646_n2088# 0.022183f
C180 source.n122 a_n1646_n2088# 0.022183f
C181 source.n123 a_n1646_n2088# 0.01192f
C182 source.n124 a_n1646_n2088# 0.012621f
C183 source.n125 a_n1646_n2088# 0.028175f
C184 source.n126 a_n1646_n2088# 0.060994f
C185 source.n127 a_n1646_n2088# 0.012621f
C186 source.n128 a_n1646_n2088# 0.01192f
C187 source.n129 a_n1646_n2088# 0.051275f
C188 source.n130 a_n1646_n2088# 0.034129f
C189 source.n131 a_n1646_n2088# 0.859871f
C190 source.n132 a_n1646_n2088# 0.03118f
C191 source.n133 a_n1646_n2088# 0.022183f
C192 source.n134 a_n1646_n2088# 0.01192f
C193 source.n135 a_n1646_n2088# 0.028175f
C194 source.n136 a_n1646_n2088# 0.012621f
C195 source.n137 a_n1646_n2088# 0.022183f
C196 source.n138 a_n1646_n2088# 0.01192f
C197 source.n139 a_n1646_n2088# 0.028175f
C198 source.n140 a_n1646_n2088# 0.012621f
C199 source.n141 a_n1646_n2088# 0.094928f
C200 source.t12 a_n1646_n2088# 0.045922f
C201 source.n142 a_n1646_n2088# 0.021131f
C202 source.n143 a_n1646_n2088# 0.016643f
C203 source.n144 a_n1646_n2088# 0.01192f
C204 source.n145 a_n1646_n2088# 0.527823f
C205 source.n146 a_n1646_n2088# 0.022183f
C206 source.n147 a_n1646_n2088# 0.01192f
C207 source.n148 a_n1646_n2088# 0.012621f
C208 source.n149 a_n1646_n2088# 0.028175f
C209 source.n150 a_n1646_n2088# 0.028175f
C210 source.n151 a_n1646_n2088# 0.012621f
C211 source.n152 a_n1646_n2088# 0.01192f
C212 source.n153 a_n1646_n2088# 0.022183f
C213 source.n154 a_n1646_n2088# 0.022183f
C214 source.n155 a_n1646_n2088# 0.01192f
C215 source.n156 a_n1646_n2088# 0.012621f
C216 source.n157 a_n1646_n2088# 0.028175f
C217 source.n158 a_n1646_n2088# 0.060994f
C218 source.n159 a_n1646_n2088# 0.012621f
C219 source.n160 a_n1646_n2088# 0.01192f
C220 source.n161 a_n1646_n2088# 0.051275f
C221 source.n162 a_n1646_n2088# 0.034129f
C222 source.n163 a_n1646_n2088# 0.859871f
C223 source.t14 a_n1646_n2088# 0.105178f
C224 source.t15 a_n1646_n2088# 0.105178f
C225 source.n164 a_n1646_n2088# 0.81913f
C226 source.n165 a_n1646_n2088# 0.322562f
C227 source.n166 a_n1646_n2088# 0.03118f
C228 source.n167 a_n1646_n2088# 0.022183f
C229 source.n168 a_n1646_n2088# 0.01192f
C230 source.n169 a_n1646_n2088# 0.028175f
C231 source.n170 a_n1646_n2088# 0.012621f
C232 source.n171 a_n1646_n2088# 0.022183f
C233 source.n172 a_n1646_n2088# 0.01192f
C234 source.n173 a_n1646_n2088# 0.028175f
C235 source.n174 a_n1646_n2088# 0.012621f
C236 source.n175 a_n1646_n2088# 0.094928f
C237 source.t13 a_n1646_n2088# 0.045922f
C238 source.n176 a_n1646_n2088# 0.021131f
C239 source.n177 a_n1646_n2088# 0.016643f
C240 source.n178 a_n1646_n2088# 0.01192f
C241 source.n179 a_n1646_n2088# 0.527823f
C242 source.n180 a_n1646_n2088# 0.022183f
C243 source.n181 a_n1646_n2088# 0.01192f
C244 source.n182 a_n1646_n2088# 0.012621f
C245 source.n183 a_n1646_n2088# 0.028175f
C246 source.n184 a_n1646_n2088# 0.028175f
C247 source.n185 a_n1646_n2088# 0.012621f
C248 source.n186 a_n1646_n2088# 0.01192f
C249 source.n187 a_n1646_n2088# 0.022183f
C250 source.n188 a_n1646_n2088# 0.022183f
C251 source.n189 a_n1646_n2088# 0.01192f
C252 source.n190 a_n1646_n2088# 0.012621f
C253 source.n191 a_n1646_n2088# 0.028175f
C254 source.n192 a_n1646_n2088# 0.060994f
C255 source.n193 a_n1646_n2088# 0.012621f
C256 source.n194 a_n1646_n2088# 0.01192f
C257 source.n195 a_n1646_n2088# 0.051275f
C258 source.n196 a_n1646_n2088# 0.034129f
C259 source.n197 a_n1646_n2088# 0.109835f
C260 source.n198 a_n1646_n2088# 0.03118f
C261 source.n199 a_n1646_n2088# 0.022183f
C262 source.n200 a_n1646_n2088# 0.01192f
C263 source.n201 a_n1646_n2088# 0.028175f
C264 source.n202 a_n1646_n2088# 0.012621f
C265 source.n203 a_n1646_n2088# 0.022183f
C266 source.n204 a_n1646_n2088# 0.01192f
C267 source.n205 a_n1646_n2088# 0.028175f
C268 source.n206 a_n1646_n2088# 0.012621f
C269 source.n207 a_n1646_n2088# 0.094928f
C270 source.t1 a_n1646_n2088# 0.045922f
C271 source.n208 a_n1646_n2088# 0.021131f
C272 source.n209 a_n1646_n2088# 0.016643f
C273 source.n210 a_n1646_n2088# 0.01192f
C274 source.n211 a_n1646_n2088# 0.527823f
C275 source.n212 a_n1646_n2088# 0.022183f
C276 source.n213 a_n1646_n2088# 0.01192f
C277 source.n214 a_n1646_n2088# 0.012621f
C278 source.n215 a_n1646_n2088# 0.028175f
C279 source.n216 a_n1646_n2088# 0.028175f
C280 source.n217 a_n1646_n2088# 0.012621f
C281 source.n218 a_n1646_n2088# 0.01192f
C282 source.n219 a_n1646_n2088# 0.022183f
C283 source.n220 a_n1646_n2088# 0.022183f
C284 source.n221 a_n1646_n2088# 0.01192f
C285 source.n222 a_n1646_n2088# 0.012621f
C286 source.n223 a_n1646_n2088# 0.028175f
C287 source.n224 a_n1646_n2088# 0.060994f
C288 source.n225 a_n1646_n2088# 0.012621f
C289 source.n226 a_n1646_n2088# 0.01192f
C290 source.n227 a_n1646_n2088# 0.051275f
C291 source.n228 a_n1646_n2088# 0.034129f
C292 source.n229 a_n1646_n2088# 0.109835f
C293 source.t2 a_n1646_n2088# 0.105178f
C294 source.t4 a_n1646_n2088# 0.105178f
C295 source.n230 a_n1646_n2088# 0.81913f
C296 source.n231 a_n1646_n2088# 0.322562f
C297 source.n232 a_n1646_n2088# 0.03118f
C298 source.n233 a_n1646_n2088# 0.022183f
C299 source.n234 a_n1646_n2088# 0.01192f
C300 source.n235 a_n1646_n2088# 0.028175f
C301 source.n236 a_n1646_n2088# 0.012621f
C302 source.n237 a_n1646_n2088# 0.022183f
C303 source.n238 a_n1646_n2088# 0.01192f
C304 source.n239 a_n1646_n2088# 0.028175f
C305 source.n240 a_n1646_n2088# 0.012621f
C306 source.n241 a_n1646_n2088# 0.094928f
C307 source.t0 a_n1646_n2088# 0.045922f
C308 source.n242 a_n1646_n2088# 0.021131f
C309 source.n243 a_n1646_n2088# 0.016643f
C310 source.n244 a_n1646_n2088# 0.01192f
C311 source.n245 a_n1646_n2088# 0.527823f
C312 source.n246 a_n1646_n2088# 0.022183f
C313 source.n247 a_n1646_n2088# 0.01192f
C314 source.n248 a_n1646_n2088# 0.012621f
C315 source.n249 a_n1646_n2088# 0.028175f
C316 source.n250 a_n1646_n2088# 0.028175f
C317 source.n251 a_n1646_n2088# 0.012621f
C318 source.n252 a_n1646_n2088# 0.01192f
C319 source.n253 a_n1646_n2088# 0.022183f
C320 source.n254 a_n1646_n2088# 0.022183f
C321 source.n255 a_n1646_n2088# 0.01192f
C322 source.n256 a_n1646_n2088# 0.012621f
C323 source.n257 a_n1646_n2088# 0.028175f
C324 source.n258 a_n1646_n2088# 0.060994f
C325 source.n259 a_n1646_n2088# 0.012621f
C326 source.n260 a_n1646_n2088# 0.01192f
C327 source.n261 a_n1646_n2088# 0.051275f
C328 source.n262 a_n1646_n2088# 0.034129f
C329 source.n263 a_n1646_n2088# 0.249707f
C330 source.n264 a_n1646_n2088# 0.916847f
C331 drain_left.t1 a_n1646_n2088# 0.130706f
C332 drain_left.t0 a_n1646_n2088# 0.130706f
C333 drain_left.n0 a_n1646_n2088# 1.09182f
C334 drain_left.t6 a_n1646_n2088# 0.130706f
C335 drain_left.t3 a_n1646_n2088# 0.130706f
C336 drain_left.n1 a_n1646_n2088# 1.09182f
C337 drain_left.n2 a_n1646_n2088# 1.62789f
C338 drain_left.t5 a_n1646_n2088# 0.130706f
C339 drain_left.t7 a_n1646_n2088# 0.130706f
C340 drain_left.n3 a_n1646_n2088# 1.09454f
C341 drain_left.t2 a_n1646_n2088# 0.130706f
C342 drain_left.t4 a_n1646_n2088# 0.130706f
C343 drain_left.n4 a_n1646_n2088# 1.09009f
C344 drain_left.n5 a_n1646_n2088# 0.979382f
C345 plus.n0 a_n1646_n2088# 0.238247f
C346 plus.t4 a_n1646_n2088# 0.510195f
C347 plus.t5 a_n1646_n2088# 0.510195f
C348 plus.t6 a_n1646_n2088# 0.510195f
C349 plus.t7 a_n1646_n2088# 0.529368f
C350 plus.n1 a_n1646_n2088# 0.220405f
C351 plus.n2 a_n1646_n2088# 0.249202f
C352 plus.n3 a_n1646_n2088# 0.249202f
C353 plus.n4 a_n1646_n2088# 0.238115f
C354 plus.n5 a_n1646_n2088# 0.448666f
C355 plus.n6 a_n1646_n2088# 0.238247f
C356 plus.t3 a_n1646_n2088# 0.510195f
C357 plus.t1 a_n1646_n2088# 0.510195f
C358 plus.t2 a_n1646_n2088# 0.529368f
C359 plus.n7 a_n1646_n2088# 0.220405f
C360 plus.t0 a_n1646_n2088# 0.510195f
C361 plus.n8 a_n1646_n2088# 0.249202f
C362 plus.n9 a_n1646_n2088# 0.249202f
C363 plus.n10 a_n1646_n2088# 0.238115f
C364 plus.n11 a_n1646_n2088# 1.23105f
.ends

