* NGSPICE file created from diffpair327.ext - technology: sky130A

.subckt diffpair327 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t25 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 drain_left.t14 plus.t1 source.t29 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 source.t26 plus.t2 drain_left.t13 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X3 source.t24 plus.t3 drain_left.t12 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X4 a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X5 source.t7 minus.t0 drain_right.t15 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X6 drain_left.t11 plus.t4 source.t21 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X7 a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X8 drain_right.t14 minus.t1 source.t9 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 drain_left.t10 plus.t5 source.t31 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X11 drain_right.t13 minus.t2 source.t11 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X12 source.t6 minus.t3 drain_right.t12 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X13 source.t28 plus.t6 drain_left.t9 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X14 a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X15 drain_right.t11 minus.t4 source.t8 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X16 drain_right.t10 minus.t5 source.t2 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X17 source.t1 minus.t6 drain_right.t9 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 source.t3 minus.t7 drain_right.t8 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t5 minus.t8 drain_right.t7 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X20 drain_left.t8 plus.t7 source.t27 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X21 source.t23 plus.t8 drain_left.t7 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X22 drain_right.t6 minus.t9 source.t10 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X23 drain_right.t5 minus.t10 source.t12 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X24 source.t0 minus.t11 drain_right.t4 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X25 drain_left.t6 plus.t9 source.t16 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X26 source.t14 minus.t12 drain_right.t3 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X27 drain_right.t2 minus.t13 source.t4 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X28 source.t22 plus.t10 drain_left.t5 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X29 source.t20 plus.t11 drain_left.t4 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X30 drain_right.t1 minus.t14 source.t13 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X31 drain_left.t3 plus.t12 source.t17 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X32 drain_left.t2 plus.t13 source.t18 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X33 source.t15 minus.t15 drain_right.t0 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X34 source.t30 plus.t14 drain_left.t1 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X35 source.t19 plus.t15 drain_left.t0 a_n1886_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n5 plus.t8 1695.03
R1 plus.n21 plus.t7 1695.03
R2 plus.n28 plus.t4 1695.03
R3 plus.n44 plus.t2 1695.03
R4 plus.n6 plus.t13 1654.87
R5 plus.n3 plus.t11 1654.87
R6 plus.n12 plus.t9 1654.87
R7 plus.n14 plus.t15 1654.87
R8 plus.n1 plus.t12 1654.87
R9 plus.n20 plus.t10 1654.87
R10 plus.n29 plus.t6 1654.87
R11 plus.n26 plus.t0 1654.87
R12 plus.n35 plus.t3 1654.87
R13 plus.n37 plus.t5 1654.87
R14 plus.n24 plus.t14 1654.87
R15 plus.n43 plus.t1 1654.87
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 69.3793
R39 plus.n15 plus.n1 69.3793
R40 plus.n38 plus.n24 69.3793
R41 plus.n34 plus.n26 69.3793
R42 plus.n6 plus.n5 54.7732
R43 plus.n21 plus.n20 54.7732
R44 plus.n44 plus.n43 54.7732
R45 plus.n29 plus.n28 54.7732
R46 plus.n13 plus.n12 47.4702
R47 plus.n14 plus.n13 47.4702
R48 plus.n37 plus.n36 47.4702
R49 plus.n36 plus.n35 47.4702
R50 plus plus.n45 29.0142
R51 plus.n12 plus.n11 25.5611
R52 plus.n15 plus.n14 25.5611
R53 plus.n38 plus.n37 25.5611
R54 plus.n35 plus.n34 25.5611
R55 plus.n7 plus.n6 18.2581
R56 plus.n20 plus.n19 18.2581
R57 plus.n43 plus.n42 18.2581
R58 plus.n30 plus.n29 18.2581
R59 plus plus.n22 11.0119
R60 plus.n8 plus.n3 3.65202
R61 plus.n18 plus.n1 3.65202
R62 plus.n41 plus.n24 3.65202
R63 plus.n31 plus.n26 3.65202
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 source.n7 source.t23 52.1921
R79 source.n8 source.t8 52.1921
R80 source.n15 source.t0 52.1921
R81 source.n31 source.t13 52.1919
R82 source.n24 source.t15 52.1919
R83 source.n23 source.t21 52.1919
R84 source.n16 source.t26 52.1919
R85 source.n0 source.t27 52.1919
R86 source.n2 source.n1 48.8588
R87 source.n4 source.n3 48.8588
R88 source.n6 source.n5 48.8588
R89 source.n10 source.n9 48.8588
R90 source.n12 source.n11 48.8588
R91 source.n14 source.n13 48.8588
R92 source.n30 source.n29 48.8586
R93 source.n28 source.n27 48.8586
R94 source.n26 source.n25 48.8586
R95 source.n22 source.n21 48.8586
R96 source.n20 source.n19 48.8586
R97 source.n18 source.n17 48.8586
R98 source.n16 source.n15 19.5753
R99 source.n32 source.n0 14.0322
R100 source.n32 source.n31 5.5436
R101 source.n29 source.t11 3.33383
R102 source.n29 source.t5 3.33383
R103 source.n27 source.t4 3.33383
R104 source.n27 source.t7 3.33383
R105 source.n25 source.t9 3.33383
R106 source.n25 source.t1 3.33383
R107 source.n21 source.t25 3.33383
R108 source.n21 source.t28 3.33383
R109 source.n19 source.t31 3.33383
R110 source.n19 source.t24 3.33383
R111 source.n17 source.t29 3.33383
R112 source.n17 source.t30 3.33383
R113 source.n1 source.t17 3.33383
R114 source.n1 source.t22 3.33383
R115 source.n3 source.t16 3.33383
R116 source.n3 source.t19 3.33383
R117 source.n5 source.t18 3.33383
R118 source.n5 source.t20 3.33383
R119 source.n9 source.t10 3.33383
R120 source.n9 source.t6 3.33383
R121 source.n11 source.t2 3.33383
R122 source.n11 source.t3 3.33383
R123 source.n13 source.t12 3.33383
R124 source.n13 source.t14 3.33383
R125 source.n15 source.n14 0.560845
R126 source.n14 source.n12 0.560845
R127 source.n12 source.n10 0.560845
R128 source.n10 source.n8 0.560845
R129 source.n7 source.n6 0.560845
R130 source.n6 source.n4 0.560845
R131 source.n4 source.n2 0.560845
R132 source.n2 source.n0 0.560845
R133 source.n18 source.n16 0.560845
R134 source.n20 source.n18 0.560845
R135 source.n22 source.n20 0.560845
R136 source.n23 source.n22 0.560845
R137 source.n26 source.n24 0.560845
R138 source.n28 source.n26 0.560845
R139 source.n30 source.n28 0.560845
R140 source.n31 source.n30 0.560845
R141 source.n8 source.n7 0.470328
R142 source.n24 source.n23 0.470328
R143 source source.n32 0.188
R144 drain_left.n9 drain_left.n7 66.0979
R145 drain_left.n5 drain_left.n3 66.0977
R146 drain_left.n2 drain_left.n0 66.0977
R147 drain_left.n11 drain_left.n10 65.5376
R148 drain_left.n9 drain_left.n8 65.5376
R149 drain_left.n13 drain_left.n12 65.5374
R150 drain_left.n5 drain_left.n4 65.5373
R151 drain_left.n2 drain_left.n1 65.5373
R152 drain_left drain_left.n6 28.7366
R153 drain_left drain_left.n13 6.21356
R154 drain_left.n3 drain_left.t9 3.33383
R155 drain_left.n3 drain_left.t11 3.33383
R156 drain_left.n4 drain_left.t12 3.33383
R157 drain_left.n4 drain_left.t15 3.33383
R158 drain_left.n1 drain_left.t1 3.33383
R159 drain_left.n1 drain_left.t10 3.33383
R160 drain_left.n0 drain_left.t13 3.33383
R161 drain_left.n0 drain_left.t14 3.33383
R162 drain_left.n12 drain_left.t5 3.33383
R163 drain_left.n12 drain_left.t8 3.33383
R164 drain_left.n10 drain_left.t0 3.33383
R165 drain_left.n10 drain_left.t3 3.33383
R166 drain_left.n8 drain_left.t4 3.33383
R167 drain_left.n8 drain_left.t6 3.33383
R168 drain_left.n7 drain_left.t7 3.33383
R169 drain_left.n7 drain_left.t2 3.33383
R170 drain_left.n11 drain_left.n9 0.560845
R171 drain_left.n13 drain_left.n11 0.560845
R172 drain_left.n6 drain_left.n5 0.225326
R173 drain_left.n6 drain_left.n2 0.225326
R174 minus.n21 minus.t11 1695.03
R175 minus.n5 minus.t4 1695.03
R176 minus.n44 minus.t14 1695.03
R177 minus.n28 minus.t15 1695.03
R178 minus.n20 minus.t10 1654.87
R179 minus.n1 minus.t12 1654.87
R180 minus.n14 minus.t5 1654.87
R181 minus.n12 minus.t7 1654.87
R182 minus.n3 minus.t9 1654.87
R183 minus.n6 minus.t3 1654.87
R184 minus.n43 minus.t8 1654.87
R185 minus.n24 minus.t2 1654.87
R186 minus.n37 minus.t0 1654.87
R187 minus.n35 minus.t13 1654.87
R188 minus.n26 minus.t6 1654.87
R189 minus.n29 minus.t1 1654.87
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 69.3793
R213 minus.n11 minus.n3 69.3793
R214 minus.n34 minus.n26 69.3793
R215 minus.n38 minus.n24 69.3793
R216 minus.n21 minus.n20 54.7732
R217 minus.n6 minus.n5 54.7732
R218 minus.n29 minus.n28 54.7732
R219 minus.n44 minus.n43 54.7732
R220 minus.n14 minus.n13 47.4702
R221 minus.n13 minus.n12 47.4702
R222 minus.n36 minus.n35 47.4702
R223 minus.n37 minus.n36 47.4702
R224 minus.n46 minus.n22 33.9967
R225 minus.n15 minus.n14 25.5611
R226 minus.n12 minus.n11 25.5611
R227 minus.n35 minus.n34 25.5611
R228 minus.n38 minus.n37 25.5611
R229 minus.n20 minus.n19 18.2581
R230 minus.n7 minus.n6 18.2581
R231 minus.n30 minus.n29 18.2581
R232 minus.n43 minus.n42 18.2581
R233 minus.n46 minus.n45 6.50429
R234 minus.n18 minus.n1 3.65202
R235 minus.n8 minus.n3 3.65202
R236 minus.n31 minus.n26 3.65202
R237 minus.n41 minus.n24 3.65202
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 66.0978
R254 drain_right.n5 drain_right.n3 66.0977
R255 drain_right.n2 drain_right.n0 66.0977
R256 drain_right.n9 drain_right.n8 65.5376
R257 drain_right.n11 drain_right.n10 65.5376
R258 drain_right.n13 drain_right.n12 65.5376
R259 drain_right.n5 drain_right.n4 65.5373
R260 drain_right.n2 drain_right.n1 65.5373
R261 drain_right drain_right.n6 28.1834
R262 drain_right drain_right.n13 6.21356
R263 drain_right.n3 drain_right.t7 3.33383
R264 drain_right.n3 drain_right.t1 3.33383
R265 drain_right.n4 drain_right.t15 3.33383
R266 drain_right.n4 drain_right.t13 3.33383
R267 drain_right.n1 drain_right.t9 3.33383
R268 drain_right.n1 drain_right.t2 3.33383
R269 drain_right.n0 drain_right.t0 3.33383
R270 drain_right.n0 drain_right.t14 3.33383
R271 drain_right.n7 drain_right.t12 3.33383
R272 drain_right.n7 drain_right.t11 3.33383
R273 drain_right.n8 drain_right.t8 3.33383
R274 drain_right.n8 drain_right.t6 3.33383
R275 drain_right.n10 drain_right.t3 3.33383
R276 drain_right.n10 drain_right.t10 3.33383
R277 drain_right.n12 drain_right.t4 3.33383
R278 drain_right.n12 drain_right.t5 3.33383
R279 drain_right.n13 drain_right.n11 0.560845
R280 drain_right.n11 drain_right.n9 0.560845
R281 drain_right.n6 drain_right.n5 0.225326
R282 drain_right.n6 drain_right.n2 0.225326
C0 plus drain_left 2.97211f
C1 drain_left minus 0.170952f
C2 drain_right source 24.084099f
C3 plus source 2.44816f
C4 minus source 2.43413f
C5 drain_right plus 0.337321f
C6 drain_left source 24.0837f
C7 drain_right minus 2.78852f
C8 drain_right drain_left 0.96779f
C9 plus minus 4.9368f
C10 drain_right a_n1886_n2688# 5.51471f
C11 drain_left a_n1886_n2688# 5.79913f
C12 source a_n1886_n2688# 7.171509f
C13 minus a_n1886_n2688# 6.763806f
C14 plus a_n1886_n2688# 8.67968f
C15 drain_right.t0 a_n1886_n2688# 0.303581f
C16 drain_right.t14 a_n1886_n2688# 0.303581f
C17 drain_right.n0 a_n1886_n2688# 1.96182f
C18 drain_right.t9 a_n1886_n2688# 0.303581f
C19 drain_right.t2 a_n1886_n2688# 0.303581f
C20 drain_right.n1 a_n1886_n2688# 1.95894f
C21 drain_right.n2 a_n1886_n2688# 0.635715f
C22 drain_right.t7 a_n1886_n2688# 0.303581f
C23 drain_right.t1 a_n1886_n2688# 0.303581f
C24 drain_right.n3 a_n1886_n2688# 1.96182f
C25 drain_right.t15 a_n1886_n2688# 0.303581f
C26 drain_right.t13 a_n1886_n2688# 0.303581f
C27 drain_right.n4 a_n1886_n2688# 1.95894f
C28 drain_right.n5 a_n1886_n2688# 0.635715f
C29 drain_right.n6 a_n1886_n2688# 1.14455f
C30 drain_right.t12 a_n1886_n2688# 0.303581f
C31 drain_right.t11 a_n1886_n2688# 0.303581f
C32 drain_right.n7 a_n1886_n2688# 1.96181f
C33 drain_right.t8 a_n1886_n2688# 0.303581f
C34 drain_right.t6 a_n1886_n2688# 0.303581f
C35 drain_right.n8 a_n1886_n2688# 1.95895f
C36 drain_right.n9 a_n1886_n2688# 0.663268f
C37 drain_right.t3 a_n1886_n2688# 0.303581f
C38 drain_right.t10 a_n1886_n2688# 0.303581f
C39 drain_right.n10 a_n1886_n2688# 1.95895f
C40 drain_right.n11 a_n1886_n2688# 0.327393f
C41 drain_right.t4 a_n1886_n2688# 0.303581f
C42 drain_right.t5 a_n1886_n2688# 0.303581f
C43 drain_right.n12 a_n1886_n2688# 1.95895f
C44 drain_right.n13 a_n1886_n2688# 0.562661f
C45 minus.n0 a_n1886_n2688# 0.052911f
C46 minus.t11 a_n1886_n2688# 0.204544f
C47 minus.t10 a_n1886_n2688# 0.202406f
C48 minus.t12 a_n1886_n2688# 0.202406f
C49 minus.n1 a_n1886_n2688# 0.092677f
C50 minus.n2 a_n1886_n2688# 0.052911f
C51 minus.t5 a_n1886_n2688# 0.202406f
C52 minus.t7 a_n1886_n2688# 0.202406f
C53 minus.t9 a_n1886_n2688# 0.202406f
C54 minus.n3 a_n1886_n2688# 0.092677f
C55 minus.n4 a_n1886_n2688# 0.112278f
C56 minus.t3 a_n1886_n2688# 0.202406f
C57 minus.t4 a_n1886_n2688# 0.204544f
C58 minus.n5 a_n1886_n2688# 0.110607f
C59 minus.n6 a_n1886_n2688# 0.092677f
C60 minus.n7 a_n1886_n2688# 0.02163f
C61 minus.n8 a_n1886_n2688# 0.018368f
C62 minus.n9 a_n1886_n2688# 0.052911f
C63 minus.n10 a_n1886_n2688# 0.052911f
C64 minus.n11 a_n1886_n2688# 0.022446f
C65 minus.n12 a_n1886_n2688# 0.092677f
C66 minus.n13 a_n1886_n2688# 0.022446f
C67 minus.n14 a_n1886_n2688# 0.092677f
C68 minus.n15 a_n1886_n2688# 0.022446f
C69 minus.n16 a_n1886_n2688# 0.052911f
C70 minus.n17 a_n1886_n2688# 0.052911f
C71 minus.n18 a_n1886_n2688# 0.018368f
C72 minus.n19 a_n1886_n2688# 0.02163f
C73 minus.n20 a_n1886_n2688# 0.092677f
C74 minus.n21 a_n1886_n2688# 0.110538f
C75 minus.n22 a_n1886_n2688# 1.69342f
C76 minus.n23 a_n1886_n2688# 0.052911f
C77 minus.t8 a_n1886_n2688# 0.202406f
C78 minus.t2 a_n1886_n2688# 0.202406f
C79 minus.n24 a_n1886_n2688# 0.092677f
C80 minus.n25 a_n1886_n2688# 0.052911f
C81 minus.t0 a_n1886_n2688# 0.202406f
C82 minus.t13 a_n1886_n2688# 0.202406f
C83 minus.t6 a_n1886_n2688# 0.202406f
C84 minus.n26 a_n1886_n2688# 0.092677f
C85 minus.n27 a_n1886_n2688# 0.112278f
C86 minus.t1 a_n1886_n2688# 0.202406f
C87 minus.t15 a_n1886_n2688# 0.204544f
C88 minus.n28 a_n1886_n2688# 0.110607f
C89 minus.n29 a_n1886_n2688# 0.092677f
C90 minus.n30 a_n1886_n2688# 0.02163f
C91 minus.n31 a_n1886_n2688# 0.018368f
C92 minus.n32 a_n1886_n2688# 0.052911f
C93 minus.n33 a_n1886_n2688# 0.052911f
C94 minus.n34 a_n1886_n2688# 0.022446f
C95 minus.n35 a_n1886_n2688# 0.092677f
C96 minus.n36 a_n1886_n2688# 0.022446f
C97 minus.n37 a_n1886_n2688# 0.092677f
C98 minus.n38 a_n1886_n2688# 0.022446f
C99 minus.n39 a_n1886_n2688# 0.052911f
C100 minus.n40 a_n1886_n2688# 0.052911f
C101 minus.n41 a_n1886_n2688# 0.018368f
C102 minus.n42 a_n1886_n2688# 0.02163f
C103 minus.n43 a_n1886_n2688# 0.092677f
C104 minus.t14 a_n1886_n2688# 0.204544f
C105 minus.n44 a_n1886_n2688# 0.110538f
C106 minus.n45 a_n1886_n2688# 0.346456f
C107 minus.n46 a_n1886_n2688# 2.06976f
C108 drain_left.t13 a_n1886_n2688# 0.30459f
C109 drain_left.t14 a_n1886_n2688# 0.30459f
C110 drain_left.n0 a_n1886_n2688# 1.96834f
C111 drain_left.t1 a_n1886_n2688# 0.30459f
C112 drain_left.t10 a_n1886_n2688# 0.30459f
C113 drain_left.n1 a_n1886_n2688# 1.96546f
C114 drain_left.n2 a_n1886_n2688# 0.637829f
C115 drain_left.t9 a_n1886_n2688# 0.30459f
C116 drain_left.t11 a_n1886_n2688# 0.30459f
C117 drain_left.n3 a_n1886_n2688# 1.96834f
C118 drain_left.t12 a_n1886_n2688# 0.30459f
C119 drain_left.t15 a_n1886_n2688# 0.30459f
C120 drain_left.n4 a_n1886_n2688# 1.96546f
C121 drain_left.n5 a_n1886_n2688# 0.637829f
C122 drain_left.n6 a_n1886_n2688# 1.20649f
C123 drain_left.t7 a_n1886_n2688# 0.30459f
C124 drain_left.t2 a_n1886_n2688# 0.30459f
C125 drain_left.n7 a_n1886_n2688# 1.96834f
C126 drain_left.t4 a_n1886_n2688# 0.30459f
C127 drain_left.t6 a_n1886_n2688# 0.30459f
C128 drain_left.n8 a_n1886_n2688# 1.96546f
C129 drain_left.n9 a_n1886_n2688# 0.665466f
C130 drain_left.t0 a_n1886_n2688# 0.30459f
C131 drain_left.t3 a_n1886_n2688# 0.30459f
C132 drain_left.n10 a_n1886_n2688# 1.96546f
C133 drain_left.n11 a_n1886_n2688# 0.328481f
C134 drain_left.t5 a_n1886_n2688# 0.30459f
C135 drain_left.t8 a_n1886_n2688# 0.30459f
C136 drain_left.n12 a_n1886_n2688# 1.96545f
C137 drain_left.n13 a_n1886_n2688# 0.564539f
C138 source.t27 a_n1886_n2688# 1.98011f
C139 source.n0 a_n1886_n2688# 1.10454f
C140 source.t17 a_n1886_n2688# 0.262f
C141 source.t22 a_n1886_n2688# 0.262f
C142 source.n1 a_n1886_n2688# 1.62573f
C143 source.n2 a_n1886_n2688# 0.314406f
C144 source.t16 a_n1886_n2688# 0.262f
C145 source.t19 a_n1886_n2688# 0.262f
C146 source.n3 a_n1886_n2688# 1.62573f
C147 source.n4 a_n1886_n2688# 0.314406f
C148 source.t18 a_n1886_n2688# 0.262f
C149 source.t20 a_n1886_n2688# 0.262f
C150 source.n5 a_n1886_n2688# 1.62573f
C151 source.n6 a_n1886_n2688# 0.314406f
C152 source.t23 a_n1886_n2688# 1.98012f
C153 source.n7 a_n1886_n2688# 0.424532f
C154 source.t8 a_n1886_n2688# 1.98012f
C155 source.n8 a_n1886_n2688# 0.424532f
C156 source.t10 a_n1886_n2688# 0.262f
C157 source.t6 a_n1886_n2688# 0.262f
C158 source.n9 a_n1886_n2688# 1.62573f
C159 source.n10 a_n1886_n2688# 0.314406f
C160 source.t2 a_n1886_n2688# 0.262f
C161 source.t3 a_n1886_n2688# 0.262f
C162 source.n11 a_n1886_n2688# 1.62573f
C163 source.n12 a_n1886_n2688# 0.314406f
C164 source.t12 a_n1886_n2688# 0.262f
C165 source.t14 a_n1886_n2688# 0.262f
C166 source.n13 a_n1886_n2688# 1.62573f
C167 source.n14 a_n1886_n2688# 0.314406f
C168 source.t0 a_n1886_n2688# 1.98012f
C169 source.n15 a_n1886_n2688# 1.45826f
C170 source.t26 a_n1886_n2688# 1.98011f
C171 source.n16 a_n1886_n2688# 1.45826f
C172 source.t29 a_n1886_n2688# 0.262f
C173 source.t30 a_n1886_n2688# 0.262f
C174 source.n17 a_n1886_n2688# 1.62573f
C175 source.n18 a_n1886_n2688# 0.31441f
C176 source.t31 a_n1886_n2688# 0.262f
C177 source.t24 a_n1886_n2688# 0.262f
C178 source.n19 a_n1886_n2688# 1.62573f
C179 source.n20 a_n1886_n2688# 0.31441f
C180 source.t25 a_n1886_n2688# 0.262f
C181 source.t28 a_n1886_n2688# 0.262f
C182 source.n21 a_n1886_n2688# 1.62573f
C183 source.n22 a_n1886_n2688# 0.31441f
C184 source.t21 a_n1886_n2688# 1.98011f
C185 source.n23 a_n1886_n2688# 0.424537f
C186 source.t15 a_n1886_n2688# 1.98011f
C187 source.n24 a_n1886_n2688# 0.424537f
C188 source.t9 a_n1886_n2688# 0.262f
C189 source.t1 a_n1886_n2688# 0.262f
C190 source.n25 a_n1886_n2688# 1.62573f
C191 source.n26 a_n1886_n2688# 0.31441f
C192 source.t4 a_n1886_n2688# 0.262f
C193 source.t7 a_n1886_n2688# 0.262f
C194 source.n27 a_n1886_n2688# 1.62573f
C195 source.n28 a_n1886_n2688# 0.31441f
C196 source.t11 a_n1886_n2688# 0.262f
C197 source.t5 a_n1886_n2688# 0.262f
C198 source.n29 a_n1886_n2688# 1.62573f
C199 source.n30 a_n1886_n2688# 0.31441f
C200 source.t13 a_n1886_n2688# 1.98011f
C201 source.n31 a_n1886_n2688# 0.562866f
C202 source.n32 a_n1886_n2688# 1.26641f
C203 plus.n0 a_n1886_n2688# 0.054537f
C204 plus.t10 a_n1886_n2688# 0.208624f
C205 plus.t12 a_n1886_n2688# 0.208624f
C206 plus.n1 a_n1886_n2688# 0.095524f
C207 plus.n2 a_n1886_n2688# 0.054537f
C208 plus.t15 a_n1886_n2688# 0.208624f
C209 plus.t9 a_n1886_n2688# 0.208624f
C210 plus.t11 a_n1886_n2688# 0.208624f
C211 plus.n3 a_n1886_n2688# 0.095524f
C212 plus.n4 a_n1886_n2688# 0.115727f
C213 plus.t13 a_n1886_n2688# 0.208624f
C214 plus.t8 a_n1886_n2688# 0.210828f
C215 plus.n5 a_n1886_n2688# 0.114006f
C216 plus.n6 a_n1886_n2688# 0.095524f
C217 plus.n7 a_n1886_n2688# 0.022295f
C218 plus.n8 a_n1886_n2688# 0.018932f
C219 plus.n9 a_n1886_n2688# 0.054537f
C220 plus.n10 a_n1886_n2688# 0.054537f
C221 plus.n11 a_n1886_n2688# 0.023135f
C222 plus.n12 a_n1886_n2688# 0.095524f
C223 plus.n13 a_n1886_n2688# 0.023135f
C224 plus.n14 a_n1886_n2688# 0.095524f
C225 plus.n15 a_n1886_n2688# 0.023135f
C226 plus.n16 a_n1886_n2688# 0.054537f
C227 plus.n17 a_n1886_n2688# 0.054537f
C228 plus.n18 a_n1886_n2688# 0.018932f
C229 plus.n19 a_n1886_n2688# 0.022295f
C230 plus.n20 a_n1886_n2688# 0.095524f
C231 plus.t7 a_n1886_n2688# 0.210828f
C232 plus.n21 a_n1886_n2688# 0.113934f
C233 plus.n22 a_n1886_n2688# 0.536283f
C234 plus.n23 a_n1886_n2688# 0.054537f
C235 plus.t2 a_n1886_n2688# 0.210828f
C236 plus.t1 a_n1886_n2688# 0.208624f
C237 plus.t14 a_n1886_n2688# 0.208624f
C238 plus.n24 a_n1886_n2688# 0.095524f
C239 plus.n25 a_n1886_n2688# 0.054537f
C240 plus.t5 a_n1886_n2688# 0.208624f
C241 plus.t3 a_n1886_n2688# 0.208624f
C242 plus.t0 a_n1886_n2688# 0.208624f
C243 plus.n26 a_n1886_n2688# 0.095524f
C244 plus.n27 a_n1886_n2688# 0.115727f
C245 plus.t6 a_n1886_n2688# 0.208624f
C246 plus.t4 a_n1886_n2688# 0.210828f
C247 plus.n28 a_n1886_n2688# 0.114006f
C248 plus.n29 a_n1886_n2688# 0.095524f
C249 plus.n30 a_n1886_n2688# 0.022295f
C250 plus.n31 a_n1886_n2688# 0.018932f
C251 plus.n32 a_n1886_n2688# 0.054537f
C252 plus.n33 a_n1886_n2688# 0.054537f
C253 plus.n34 a_n1886_n2688# 0.023135f
C254 plus.n35 a_n1886_n2688# 0.095524f
C255 plus.n36 a_n1886_n2688# 0.023135f
C256 plus.n37 a_n1886_n2688# 0.095524f
C257 plus.n38 a_n1886_n2688# 0.023135f
C258 plus.n39 a_n1886_n2688# 0.054537f
C259 plus.n40 a_n1886_n2688# 0.054537f
C260 plus.n41 a_n1886_n2688# 0.018932f
C261 plus.n42 a_n1886_n2688# 0.022295f
C262 plus.n43 a_n1886_n2688# 0.095524f
C263 plus.n44 a_n1886_n2688# 0.113934f
C264 plus.n45 a_n1886_n2688# 1.52257f
.ends

