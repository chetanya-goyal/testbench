* NGSPICE file created from diffpair217.ext - technology: sky130A

.subckt diffpair217 minus drain_right drain_left source plus
X0 a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X1 drain_right.t15 minus.t0 source.t23 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X2 source.t28 minus.t1 drain_right.t14 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X3 drain_left.t15 plus.t0 source.t9 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X4 source.t6 plus.t1 drain_left.t14 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X5 drain_left.t13 plus.t2 source.t14 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X6 source.t26 minus.t2 drain_right.t13 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X7 source.t21 minus.t3 drain_right.t12 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X8 drain_right.t11 minus.t4 source.t27 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X9 source.t31 plus.t3 drain_left.t12 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X10 drain_right.t10 minus.t5 source.t24 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X11 drain_right.t9 minus.t6 source.t16 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 source.t22 minus.t7 drain_right.t8 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X13 drain_left.t11 plus.t4 source.t3 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X14 drain_left.t10 plus.t5 source.t10 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X15 source.t4 plus.t6 drain_left.t9 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X16 source.t25 minus.t8 drain_right.t7 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X17 source.t18 minus.t9 drain_right.t6 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X18 drain_right.t5 minus.t10 source.t17 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X19 source.t8 plus.t7 drain_left.t8 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X20 a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X21 drain_left.t7 plus.t8 source.t11 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X22 source.t19 minus.t11 drain_right.t4 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X23 drain_right.t3 minus.t12 source.t15 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X24 drain_right.t2 minus.t13 source.t29 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X25 source.t0 plus.t9 drain_left.t6 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X26 a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X27 source.t12 plus.t10 drain_left.t5 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X28 drain_right.t1 minus.t14 source.t30 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X29 source.t20 minus.t15 drain_right.t0 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X30 drain_left.t4 plus.t11 source.t1 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X31 source.t7 plus.t12 drain_left.t3 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X32 a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X33 drain_left.t2 plus.t13 source.t2 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X34 drain_left.t1 plus.t14 source.t13 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X35 source.t5 plus.t15 drain_left.t0 a_n2390_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n6 minus.t14 206.953
R1 minus.n30 minus.t15 206.953
R2 minus.n5 minus.t11 185.972
R3 minus.n9 minus.t10 185.972
R4 minus.n3 minus.t8 185.972
R5 minus.n15 minus.t5 185.972
R6 minus.n1 minus.t7 185.972
R7 minus.n21 minus.t6 185.972
R8 minus.n22 minus.t2 185.972
R9 minus.n29 minus.t4 185.972
R10 minus.n33 minus.t1 185.972
R11 minus.n27 minus.t13 185.972
R12 minus.n39 minus.t9 185.972
R13 minus.n25 minus.t12 185.972
R14 minus.n45 minus.t3 185.972
R15 minus.n46 minus.t0 185.972
R16 minus.n23 minus.n22 161.3
R17 minus.n21 minus.n0 161.3
R18 minus.n20 minus.n19 161.3
R19 minus.n18 minus.n1 161.3
R20 minus.n17 minus.n16 161.3
R21 minus.n15 minus.n2 161.3
R22 minus.n14 minus.n13 161.3
R23 minus.n12 minus.n3 161.3
R24 minus.n11 minus.n10 161.3
R25 minus.n9 minus.n4 161.3
R26 minus.n8 minus.n7 161.3
R27 minus.n47 minus.n46 161.3
R28 minus.n45 minus.n24 161.3
R29 minus.n44 minus.n43 161.3
R30 minus.n42 minus.n25 161.3
R31 minus.n41 minus.n40 161.3
R32 minus.n39 minus.n26 161.3
R33 minus.n38 minus.n37 161.3
R34 minus.n36 minus.n27 161.3
R35 minus.n35 minus.n34 161.3
R36 minus.n33 minus.n28 161.3
R37 minus.n32 minus.n31 161.3
R38 minus.n7 minus.n6 70.4033
R39 minus.n31 minus.n30 70.4033
R40 minus.n22 minus.n21 48.2005
R41 minus.n46 minus.n45 48.2005
R42 minus.n9 minus.n8 44.549
R43 minus.n20 minus.n1 44.549
R44 minus.n33 minus.n32 44.549
R45 minus.n44 minus.n25 44.549
R46 minus.n10 minus.n3 34.3247
R47 minus.n16 minus.n15 34.3247
R48 minus.n34 minus.n27 34.3247
R49 minus.n40 minus.n39 34.3247
R50 minus.n48 minus.n23 31.5119
R51 minus.n15 minus.n14 24.1005
R52 minus.n14 minus.n3 24.1005
R53 minus.n38 minus.n27 24.1005
R54 minus.n39 minus.n38 24.1005
R55 minus.n6 minus.n5 20.9576
R56 minus.n30 minus.n29 20.9576
R57 minus.n10 minus.n9 13.8763
R58 minus.n16 minus.n1 13.8763
R59 minus.n34 minus.n33 13.8763
R60 minus.n40 minus.n25 13.8763
R61 minus.n48 minus.n47 6.6558
R62 minus.n8 minus.n5 3.65202
R63 minus.n21 minus.n20 3.65202
R64 minus.n32 minus.n29 3.65202
R65 minus.n45 minus.n44 3.65202
R66 minus.n23 minus.n0 0.189894
R67 minus.n19 minus.n0 0.189894
R68 minus.n19 minus.n18 0.189894
R69 minus.n18 minus.n17 0.189894
R70 minus.n17 minus.n2 0.189894
R71 minus.n13 minus.n2 0.189894
R72 minus.n13 minus.n12 0.189894
R73 minus.n12 minus.n11 0.189894
R74 minus.n11 minus.n4 0.189894
R75 minus.n7 minus.n4 0.189894
R76 minus.n31 minus.n28 0.189894
R77 minus.n35 minus.n28 0.189894
R78 minus.n36 minus.n35 0.189894
R79 minus.n37 minus.n36 0.189894
R80 minus.n37 minus.n26 0.189894
R81 minus.n41 minus.n26 0.189894
R82 minus.n42 minus.n41 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n24 0.189894
R85 minus.n47 minus.n24 0.189894
R86 minus minus.n48 0.188
R87 source.n0 source.t9 69.6943
R88 source.n7 source.t7 69.6943
R89 source.n8 source.t30 69.6943
R90 source.n15 source.t26 69.6943
R91 source.n31 source.t23 69.6942
R92 source.n24 source.t20 69.6942
R93 source.n23 source.t3 69.6942
R94 source.n16 source.t0 69.6942
R95 source.n2 source.n1 63.0943
R96 source.n4 source.n3 63.0943
R97 source.n6 source.n5 63.0943
R98 source.n10 source.n9 63.0943
R99 source.n12 source.n11 63.0943
R100 source.n14 source.n13 63.0943
R101 source.n30 source.n29 63.0942
R102 source.n28 source.n27 63.0942
R103 source.n26 source.n25 63.0942
R104 source.n22 source.n21 63.0942
R105 source.n20 source.n19 63.0942
R106 source.n18 source.n17 63.0942
R107 source.n16 source.n15 15.2713
R108 source.n32 source.n0 9.60747
R109 source.n29 source.t15 6.6005
R110 source.n29 source.t21 6.6005
R111 source.n27 source.t29 6.6005
R112 source.n27 source.t18 6.6005
R113 source.n25 source.t27 6.6005
R114 source.n25 source.t28 6.6005
R115 source.n21 source.t2 6.6005
R116 source.n21 source.t5 6.6005
R117 source.n19 source.t10 6.6005
R118 source.n19 source.t8 6.6005
R119 source.n17 source.t13 6.6005
R120 source.n17 source.t31 6.6005
R121 source.n1 source.t14 6.6005
R122 source.n1 source.t6 6.6005
R123 source.n3 source.t11 6.6005
R124 source.n3 source.t4 6.6005
R125 source.n5 source.t1 6.6005
R126 source.n5 source.t12 6.6005
R127 source.n9 source.t17 6.6005
R128 source.n9 source.t19 6.6005
R129 source.n11 source.t24 6.6005
R130 source.n11 source.t25 6.6005
R131 source.n13 source.t16 6.6005
R132 source.n13 source.t22 6.6005
R133 source.n32 source.n31 5.66429
R134 source.n15 source.n14 0.802224
R135 source.n14 source.n12 0.802224
R136 source.n12 source.n10 0.802224
R137 source.n10 source.n8 0.802224
R138 source.n7 source.n6 0.802224
R139 source.n6 source.n4 0.802224
R140 source.n4 source.n2 0.802224
R141 source.n2 source.n0 0.802224
R142 source.n18 source.n16 0.802224
R143 source.n20 source.n18 0.802224
R144 source.n22 source.n20 0.802224
R145 source.n23 source.n22 0.802224
R146 source.n26 source.n24 0.802224
R147 source.n28 source.n26 0.802224
R148 source.n30 source.n28 0.802224
R149 source.n31 source.n30 0.802224
R150 source.n8 source.n7 0.470328
R151 source.n24 source.n23 0.470328
R152 source source.n32 0.188
R153 drain_right.n9 drain_right.n7 80.5748
R154 drain_right.n5 drain_right.n3 80.5747
R155 drain_right.n2 drain_right.n0 80.5747
R156 drain_right.n9 drain_right.n8 79.7731
R157 drain_right.n11 drain_right.n10 79.7731
R158 drain_right.n13 drain_right.n12 79.7731
R159 drain_right.n5 drain_right.n4 79.773
R160 drain_right.n2 drain_right.n1 79.773
R161 drain_right drain_right.n6 25.2069
R162 drain_right.n3 drain_right.t12 6.6005
R163 drain_right.n3 drain_right.t15 6.6005
R164 drain_right.n4 drain_right.t6 6.6005
R165 drain_right.n4 drain_right.t3 6.6005
R166 drain_right.n1 drain_right.t14 6.6005
R167 drain_right.n1 drain_right.t2 6.6005
R168 drain_right.n0 drain_right.t0 6.6005
R169 drain_right.n0 drain_right.t11 6.6005
R170 drain_right.n7 drain_right.t4 6.6005
R171 drain_right.n7 drain_right.t1 6.6005
R172 drain_right.n8 drain_right.t7 6.6005
R173 drain_right.n8 drain_right.t5 6.6005
R174 drain_right.n10 drain_right.t8 6.6005
R175 drain_right.n10 drain_right.t10 6.6005
R176 drain_right.n12 drain_right.t13 6.6005
R177 drain_right.n12 drain_right.t9 6.6005
R178 drain_right drain_right.n13 6.45494
R179 drain_right.n13 drain_right.n11 0.802224
R180 drain_right.n11 drain_right.n9 0.802224
R181 drain_right.n6 drain_right.n5 0.346016
R182 drain_right.n6 drain_right.n2 0.346016
R183 plus.n6 plus.t12 206.953
R184 plus.n30 plus.t4 206.953
R185 plus.n22 plus.t0 185.972
R186 plus.n21 plus.t1 185.972
R187 plus.n1 plus.t2 185.972
R188 plus.n15 plus.t6 185.972
R189 plus.n3 plus.t8 185.972
R190 plus.n9 plus.t10 185.972
R191 plus.n5 plus.t11 185.972
R192 plus.n46 plus.t9 185.972
R193 plus.n45 plus.t14 185.972
R194 plus.n25 plus.t3 185.972
R195 plus.n39 plus.t5 185.972
R196 plus.n27 plus.t7 185.972
R197 plus.n33 plus.t13 185.972
R198 plus.n29 plus.t15 185.972
R199 plus.n8 plus.n7 161.3
R200 plus.n9 plus.n4 161.3
R201 plus.n11 plus.n10 161.3
R202 plus.n12 plus.n3 161.3
R203 plus.n14 plus.n13 161.3
R204 plus.n15 plus.n2 161.3
R205 plus.n17 plus.n16 161.3
R206 plus.n18 plus.n1 161.3
R207 plus.n20 plus.n19 161.3
R208 plus.n21 plus.n0 161.3
R209 plus.n23 plus.n22 161.3
R210 plus.n32 plus.n31 161.3
R211 plus.n33 plus.n28 161.3
R212 plus.n35 plus.n34 161.3
R213 plus.n36 plus.n27 161.3
R214 plus.n38 plus.n37 161.3
R215 plus.n39 plus.n26 161.3
R216 plus.n41 plus.n40 161.3
R217 plus.n42 plus.n25 161.3
R218 plus.n44 plus.n43 161.3
R219 plus.n45 plus.n24 161.3
R220 plus.n47 plus.n46 161.3
R221 plus.n7 plus.n6 70.4033
R222 plus.n31 plus.n30 70.4033
R223 plus.n22 plus.n21 48.2005
R224 plus.n46 plus.n45 48.2005
R225 plus.n20 plus.n1 44.549
R226 plus.n9 plus.n8 44.549
R227 plus.n44 plus.n25 44.549
R228 plus.n33 plus.n32 44.549
R229 plus.n16 plus.n15 34.3247
R230 plus.n10 plus.n3 34.3247
R231 plus.n40 plus.n39 34.3247
R232 plus.n34 plus.n27 34.3247
R233 plus plus.n47 28.8021
R234 plus.n14 plus.n3 24.1005
R235 plus.n15 plus.n14 24.1005
R236 plus.n39 plus.n38 24.1005
R237 plus.n38 plus.n27 24.1005
R238 plus.n6 plus.n5 20.9576
R239 plus.n30 plus.n29 20.9576
R240 plus.n16 plus.n1 13.8763
R241 plus.n10 plus.n9 13.8763
R242 plus.n40 plus.n25 13.8763
R243 plus.n34 plus.n33 13.8763
R244 plus plus.n23 8.89065
R245 plus.n21 plus.n20 3.65202
R246 plus.n8 plus.n5 3.65202
R247 plus.n45 plus.n44 3.65202
R248 plus.n32 plus.n29 3.65202
R249 plus.n7 plus.n4 0.189894
R250 plus.n11 plus.n4 0.189894
R251 plus.n12 plus.n11 0.189894
R252 plus.n13 plus.n12 0.189894
R253 plus.n13 plus.n2 0.189894
R254 plus.n17 plus.n2 0.189894
R255 plus.n18 plus.n17 0.189894
R256 plus.n19 plus.n18 0.189894
R257 plus.n19 plus.n0 0.189894
R258 plus.n23 plus.n0 0.189894
R259 plus.n47 plus.n24 0.189894
R260 plus.n43 plus.n24 0.189894
R261 plus.n43 plus.n42 0.189894
R262 plus.n42 plus.n41 0.189894
R263 plus.n41 plus.n26 0.189894
R264 plus.n37 plus.n26 0.189894
R265 plus.n37 plus.n36 0.189894
R266 plus.n36 plus.n35 0.189894
R267 plus.n35 plus.n28 0.189894
R268 plus.n31 plus.n28 0.189894
R269 drain_left.n9 drain_left.n7 80.5748
R270 drain_left.n5 drain_left.n3 80.5747
R271 drain_left.n2 drain_left.n0 80.5747
R272 drain_left.n13 drain_left.n12 79.7731
R273 drain_left.n11 drain_left.n10 79.7731
R274 drain_left.n9 drain_left.n8 79.7731
R275 drain_left.n5 drain_left.n4 79.773
R276 drain_left.n2 drain_left.n1 79.773
R277 drain_left drain_left.n6 25.7601
R278 drain_left.n3 drain_left.t0 6.6005
R279 drain_left.n3 drain_left.t11 6.6005
R280 drain_left.n4 drain_left.t8 6.6005
R281 drain_left.n4 drain_left.t2 6.6005
R282 drain_left.n1 drain_left.t12 6.6005
R283 drain_left.n1 drain_left.t10 6.6005
R284 drain_left.n0 drain_left.t6 6.6005
R285 drain_left.n0 drain_left.t1 6.6005
R286 drain_left.n12 drain_left.t14 6.6005
R287 drain_left.n12 drain_left.t15 6.6005
R288 drain_left.n10 drain_left.t9 6.6005
R289 drain_left.n10 drain_left.t13 6.6005
R290 drain_left.n8 drain_left.t5 6.6005
R291 drain_left.n8 drain_left.t7 6.6005
R292 drain_left.n7 drain_left.t3 6.6005
R293 drain_left.n7 drain_left.t4 6.6005
R294 drain_left drain_left.n13 6.45494
R295 drain_left.n11 drain_left.n9 0.802224
R296 drain_left.n13 drain_left.n11 0.802224
R297 drain_left.n6 drain_left.n5 0.346016
R298 drain_left.n6 drain_left.n2 0.346016
C0 drain_left minus 0.177775f
C1 drain_left plus 3.00399f
C2 source minus 3.19711f
C3 drain_right minus 2.76814f
C4 source plus 3.21111f
C5 drain_right plus 0.397563f
C6 drain_left source 7.81889f
C7 drain_left drain_right 1.24373f
C8 plus minus 4.46428f
C9 source drain_right 7.82061f
C10 drain_right a_n2390_n1488# 4.86645f
C11 drain_left a_n2390_n1488# 5.21621f
C12 source a_n2390_n1488# 3.893904f
C13 minus a_n2390_n1488# 8.742348f
C14 plus a_n2390_n1488# 10.096221f
C15 drain_left.t6 a_n2390_n1488# 0.065628f
C16 drain_left.t1 a_n2390_n1488# 0.065628f
C17 drain_left.n0 a_n2390_n1488# 0.477041f
C18 drain_left.t12 a_n2390_n1488# 0.065628f
C19 drain_left.t10 a_n2390_n1488# 0.065628f
C20 drain_left.n1 a_n2390_n1488# 0.473302f
C21 drain_left.n2 a_n2390_n1488# 0.69783f
C22 drain_left.t0 a_n2390_n1488# 0.065628f
C23 drain_left.t11 a_n2390_n1488# 0.065628f
C24 drain_left.n3 a_n2390_n1488# 0.477041f
C25 drain_left.t8 a_n2390_n1488# 0.065628f
C26 drain_left.t2 a_n2390_n1488# 0.065628f
C27 drain_left.n4 a_n2390_n1488# 0.473302f
C28 drain_left.n5 a_n2390_n1488# 0.69783f
C29 drain_left.n6 a_n2390_n1488# 1.00767f
C30 drain_left.t3 a_n2390_n1488# 0.065628f
C31 drain_left.t4 a_n2390_n1488# 0.065628f
C32 drain_left.n7 a_n2390_n1488# 0.477043f
C33 drain_left.t5 a_n2390_n1488# 0.065628f
C34 drain_left.t7 a_n2390_n1488# 0.065628f
C35 drain_left.n8 a_n2390_n1488# 0.473304f
C36 drain_left.n9 a_n2390_n1488# 0.736662f
C37 drain_left.t9 a_n2390_n1488# 0.065628f
C38 drain_left.t13 a_n2390_n1488# 0.065628f
C39 drain_left.n10 a_n2390_n1488# 0.473304f
C40 drain_left.n11 a_n2390_n1488# 0.364625f
C41 drain_left.t14 a_n2390_n1488# 0.065628f
C42 drain_left.t15 a_n2390_n1488# 0.065628f
C43 drain_left.n12 a_n2390_n1488# 0.473304f
C44 drain_left.n13 a_n2390_n1488# 0.606019f
C45 plus.n0 a_n2390_n1488# 0.045811f
C46 plus.t0 a_n2390_n1488# 0.247267f
C47 plus.t1 a_n2390_n1488# 0.247267f
C48 plus.t2 a_n2390_n1488# 0.247267f
C49 plus.n1 a_n2390_n1488# 0.148203f
C50 plus.n2 a_n2390_n1488# 0.045811f
C51 plus.t6 a_n2390_n1488# 0.247267f
C52 plus.t8 a_n2390_n1488# 0.247267f
C53 plus.n3 a_n2390_n1488# 0.148203f
C54 plus.n4 a_n2390_n1488# 0.045811f
C55 plus.t10 a_n2390_n1488# 0.247267f
C56 plus.t11 a_n2390_n1488# 0.247267f
C57 plus.n5 a_n2390_n1488# 0.146932f
C58 plus.t12 a_n2390_n1488# 0.262099f
C59 plus.n6 a_n2390_n1488# 0.13176f
C60 plus.n7 a_n2390_n1488# 0.154295f
C61 plus.n8 a_n2390_n1488# 0.010396f
C62 plus.n9 a_n2390_n1488# 0.148203f
C63 plus.n10 a_n2390_n1488# 0.010396f
C64 plus.n11 a_n2390_n1488# 0.045811f
C65 plus.n12 a_n2390_n1488# 0.045811f
C66 plus.n13 a_n2390_n1488# 0.045811f
C67 plus.n14 a_n2390_n1488# 0.010396f
C68 plus.n15 a_n2390_n1488# 0.148203f
C69 plus.n16 a_n2390_n1488# 0.010396f
C70 plus.n17 a_n2390_n1488# 0.045811f
C71 plus.n18 a_n2390_n1488# 0.045811f
C72 plus.n19 a_n2390_n1488# 0.045811f
C73 plus.n20 a_n2390_n1488# 0.010396f
C74 plus.n21 a_n2390_n1488# 0.146932f
C75 plus.n22 a_n2390_n1488# 0.146225f
C76 plus.n23 a_n2390_n1488# 0.359792f
C77 plus.n24 a_n2390_n1488# 0.045811f
C78 plus.t9 a_n2390_n1488# 0.247267f
C79 plus.t14 a_n2390_n1488# 0.247267f
C80 plus.t3 a_n2390_n1488# 0.247267f
C81 plus.n25 a_n2390_n1488# 0.148203f
C82 plus.n26 a_n2390_n1488# 0.045811f
C83 plus.t5 a_n2390_n1488# 0.247267f
C84 plus.t7 a_n2390_n1488# 0.247267f
C85 plus.n27 a_n2390_n1488# 0.148203f
C86 plus.n28 a_n2390_n1488# 0.045811f
C87 plus.t13 a_n2390_n1488# 0.247267f
C88 plus.t15 a_n2390_n1488# 0.247267f
C89 plus.n29 a_n2390_n1488# 0.146932f
C90 plus.t4 a_n2390_n1488# 0.262099f
C91 plus.n30 a_n2390_n1488# 0.13176f
C92 plus.n31 a_n2390_n1488# 0.154295f
C93 plus.n32 a_n2390_n1488# 0.010396f
C94 plus.n33 a_n2390_n1488# 0.148203f
C95 plus.n34 a_n2390_n1488# 0.010396f
C96 plus.n35 a_n2390_n1488# 0.045811f
C97 plus.n36 a_n2390_n1488# 0.045811f
C98 plus.n37 a_n2390_n1488# 0.045811f
C99 plus.n38 a_n2390_n1488# 0.010396f
C100 plus.n39 a_n2390_n1488# 0.148203f
C101 plus.n40 a_n2390_n1488# 0.010396f
C102 plus.n41 a_n2390_n1488# 0.045811f
C103 plus.n42 a_n2390_n1488# 0.045811f
C104 plus.n43 a_n2390_n1488# 0.045811f
C105 plus.n44 a_n2390_n1488# 0.010396f
C106 plus.n45 a_n2390_n1488# 0.146932f
C107 plus.n46 a_n2390_n1488# 0.146225f
C108 plus.n47 a_n2390_n1488# 1.22208f
C109 drain_right.t0 a_n2390_n1488# 0.065065f
C110 drain_right.t11 a_n2390_n1488# 0.065065f
C111 drain_right.n0 a_n2390_n1488# 0.472949f
C112 drain_right.t14 a_n2390_n1488# 0.065065f
C113 drain_right.t2 a_n2390_n1488# 0.065065f
C114 drain_right.n1 a_n2390_n1488# 0.469242f
C115 drain_right.n2 a_n2390_n1488# 0.691844f
C116 drain_right.t12 a_n2390_n1488# 0.065065f
C117 drain_right.t15 a_n2390_n1488# 0.065065f
C118 drain_right.n3 a_n2390_n1488# 0.472949f
C119 drain_right.t6 a_n2390_n1488# 0.065065f
C120 drain_right.t3 a_n2390_n1488# 0.065065f
C121 drain_right.n4 a_n2390_n1488# 0.469242f
C122 drain_right.n5 a_n2390_n1488# 0.691844f
C123 drain_right.n6 a_n2390_n1488# 0.944994f
C124 drain_right.t4 a_n2390_n1488# 0.065065f
C125 drain_right.t1 a_n2390_n1488# 0.065065f
C126 drain_right.n7 a_n2390_n1488# 0.472951f
C127 drain_right.t7 a_n2390_n1488# 0.065065f
C128 drain_right.t5 a_n2390_n1488# 0.065065f
C129 drain_right.n8 a_n2390_n1488# 0.469245f
C130 drain_right.n9 a_n2390_n1488# 0.730343f
C131 drain_right.t8 a_n2390_n1488# 0.065065f
C132 drain_right.t10 a_n2390_n1488# 0.065065f
C133 drain_right.n10 a_n2390_n1488# 0.469245f
C134 drain_right.n11 a_n2390_n1488# 0.361498f
C135 drain_right.t13 a_n2390_n1488# 0.065065f
C136 drain_right.t9 a_n2390_n1488# 0.065065f
C137 drain_right.n12 a_n2390_n1488# 0.469245f
C138 drain_right.n13 a_n2390_n1488# 0.600821f
C139 source.t9 a_n2390_n1488# 0.556694f
C140 source.n0 a_n2390_n1488# 0.800938f
C141 source.t14 a_n2390_n1488# 0.067041f
C142 source.t6 a_n2390_n1488# 0.067041f
C143 source.n1 a_n2390_n1488# 0.425076f
C144 source.n2 a_n2390_n1488# 0.392454f
C145 source.t11 a_n2390_n1488# 0.067041f
C146 source.t4 a_n2390_n1488# 0.067041f
C147 source.n3 a_n2390_n1488# 0.425076f
C148 source.n4 a_n2390_n1488# 0.392454f
C149 source.t1 a_n2390_n1488# 0.067041f
C150 source.t12 a_n2390_n1488# 0.067041f
C151 source.n5 a_n2390_n1488# 0.425076f
C152 source.n6 a_n2390_n1488# 0.392454f
C153 source.t7 a_n2390_n1488# 0.556694f
C154 source.n7 a_n2390_n1488# 0.413432f
C155 source.t30 a_n2390_n1488# 0.556694f
C156 source.n8 a_n2390_n1488# 0.413432f
C157 source.t17 a_n2390_n1488# 0.067041f
C158 source.t19 a_n2390_n1488# 0.067041f
C159 source.n9 a_n2390_n1488# 0.425076f
C160 source.n10 a_n2390_n1488# 0.392454f
C161 source.t24 a_n2390_n1488# 0.067041f
C162 source.t25 a_n2390_n1488# 0.067041f
C163 source.n11 a_n2390_n1488# 0.425076f
C164 source.n12 a_n2390_n1488# 0.392454f
C165 source.t16 a_n2390_n1488# 0.067041f
C166 source.t22 a_n2390_n1488# 0.067041f
C167 source.n13 a_n2390_n1488# 0.425076f
C168 source.n14 a_n2390_n1488# 0.392454f
C169 source.t26 a_n2390_n1488# 0.556694f
C170 source.n15 a_n2390_n1488# 1.10142f
C171 source.t0 a_n2390_n1488# 0.556691f
C172 source.n16 a_n2390_n1488# 1.10142f
C173 source.t13 a_n2390_n1488# 0.067041f
C174 source.t31 a_n2390_n1488# 0.067041f
C175 source.n17 a_n2390_n1488# 0.425073f
C176 source.n18 a_n2390_n1488# 0.392457f
C177 source.t10 a_n2390_n1488# 0.067041f
C178 source.t8 a_n2390_n1488# 0.067041f
C179 source.n19 a_n2390_n1488# 0.425073f
C180 source.n20 a_n2390_n1488# 0.392457f
C181 source.t2 a_n2390_n1488# 0.067041f
C182 source.t5 a_n2390_n1488# 0.067041f
C183 source.n21 a_n2390_n1488# 0.425073f
C184 source.n22 a_n2390_n1488# 0.392457f
C185 source.t3 a_n2390_n1488# 0.556691f
C186 source.n23 a_n2390_n1488# 0.413435f
C187 source.t20 a_n2390_n1488# 0.556691f
C188 source.n24 a_n2390_n1488# 0.413435f
C189 source.t27 a_n2390_n1488# 0.067041f
C190 source.t28 a_n2390_n1488# 0.067041f
C191 source.n25 a_n2390_n1488# 0.425073f
C192 source.n26 a_n2390_n1488# 0.392457f
C193 source.t29 a_n2390_n1488# 0.067041f
C194 source.t18 a_n2390_n1488# 0.067041f
C195 source.n27 a_n2390_n1488# 0.425073f
C196 source.n28 a_n2390_n1488# 0.392457f
C197 source.t15 a_n2390_n1488# 0.067041f
C198 source.t21 a_n2390_n1488# 0.067041f
C199 source.n29 a_n2390_n1488# 0.425073f
C200 source.n30 a_n2390_n1488# 0.392457f
C201 source.t23 a_n2390_n1488# 0.556691f
C202 source.n31 a_n2390_n1488# 0.591744f
C203 source.n32 a_n2390_n1488# 0.830271f
C204 minus.n0 a_n2390_n1488# 0.044569f
C205 minus.t7 a_n2390_n1488# 0.240563f
C206 minus.n1 a_n2390_n1488# 0.144184f
C207 minus.n2 a_n2390_n1488# 0.044569f
C208 minus.t8 a_n2390_n1488# 0.240563f
C209 minus.n3 a_n2390_n1488# 0.144184f
C210 minus.n4 a_n2390_n1488# 0.044569f
C211 minus.t11 a_n2390_n1488# 0.240563f
C212 minus.n5 a_n2390_n1488# 0.142948f
C213 minus.t14 a_n2390_n1488# 0.254993f
C214 minus.n6 a_n2390_n1488# 0.128187f
C215 minus.n7 a_n2390_n1488# 0.150112f
C216 minus.n8 a_n2390_n1488# 0.010114f
C217 minus.t10 a_n2390_n1488# 0.240563f
C218 minus.n9 a_n2390_n1488# 0.144184f
C219 minus.n10 a_n2390_n1488# 0.010114f
C220 minus.n11 a_n2390_n1488# 0.044569f
C221 minus.n12 a_n2390_n1488# 0.044569f
C222 minus.n13 a_n2390_n1488# 0.044569f
C223 minus.n14 a_n2390_n1488# 0.010114f
C224 minus.t5 a_n2390_n1488# 0.240563f
C225 minus.n15 a_n2390_n1488# 0.144184f
C226 minus.n16 a_n2390_n1488# 0.010114f
C227 minus.n17 a_n2390_n1488# 0.044569f
C228 minus.n18 a_n2390_n1488# 0.044569f
C229 minus.n19 a_n2390_n1488# 0.044569f
C230 minus.n20 a_n2390_n1488# 0.010114f
C231 minus.t6 a_n2390_n1488# 0.240563f
C232 minus.n21 a_n2390_n1488# 0.142948f
C233 minus.t2 a_n2390_n1488# 0.240563f
C234 minus.n22 a_n2390_n1488# 0.142261f
C235 minus.n23 a_n2390_n1488# 1.26582f
C236 minus.n24 a_n2390_n1488# 0.044569f
C237 minus.t12 a_n2390_n1488# 0.240563f
C238 minus.n25 a_n2390_n1488# 0.144184f
C239 minus.n26 a_n2390_n1488# 0.044569f
C240 minus.t13 a_n2390_n1488# 0.240563f
C241 minus.n27 a_n2390_n1488# 0.144184f
C242 minus.n28 a_n2390_n1488# 0.044569f
C243 minus.t4 a_n2390_n1488# 0.240563f
C244 minus.n29 a_n2390_n1488# 0.142948f
C245 minus.t15 a_n2390_n1488# 0.254993f
C246 minus.n30 a_n2390_n1488# 0.128187f
C247 minus.n31 a_n2390_n1488# 0.150112f
C248 minus.n32 a_n2390_n1488# 0.010114f
C249 minus.t1 a_n2390_n1488# 0.240563f
C250 minus.n33 a_n2390_n1488# 0.144184f
C251 minus.n34 a_n2390_n1488# 0.010114f
C252 minus.n35 a_n2390_n1488# 0.044569f
C253 minus.n36 a_n2390_n1488# 0.044569f
C254 minus.n37 a_n2390_n1488# 0.044569f
C255 minus.n38 a_n2390_n1488# 0.010114f
C256 minus.t9 a_n2390_n1488# 0.240563f
C257 minus.n39 a_n2390_n1488# 0.144184f
C258 minus.n40 a_n2390_n1488# 0.010114f
C259 minus.n41 a_n2390_n1488# 0.044569f
C260 minus.n42 a_n2390_n1488# 0.044569f
C261 minus.n43 a_n2390_n1488# 0.044569f
C262 minus.n44 a_n2390_n1488# 0.010114f
C263 minus.t3 a_n2390_n1488# 0.240563f
C264 minus.n45 a_n2390_n1488# 0.142948f
C265 minus.t0 a_n2390_n1488# 0.240563f
C266 minus.n46 a_n2390_n1488# 0.142261f
C267 minus.n47 a_n2390_n1488# 0.30762f
C268 minus.n48 a_n2390_n1488# 1.54967f
.ends

