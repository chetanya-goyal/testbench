* NGSPICE file created from diffpair365.ext - technology: sky130A

.subckt diffpair365 minus drain_right drain_left source plus
X0 a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X1 source.t19 minus.t0 drain_right.t4 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 drain_left.t11 plus.t0 source.t1 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 source.t18 minus.t1 drain_right.t10 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 source.t5 plus.t1 drain_left.t10 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X5 drain_right.t1 minus.t2 source.t17 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 source.t7 plus.t2 drain_left.t9 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X7 drain_right.t2 minus.t3 source.t16 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X8 drain_right.t6 minus.t4 source.t15 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 source.t14 minus.t5 drain_right.t8 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X11 drain_left.t8 plus.t3 source.t6 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 drain_right.t0 minus.t6 source.t13 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X13 source.t12 minus.t7 drain_right.t5 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X14 a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X15 drain_right.t7 minus.t8 source.t11 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X16 drain_left.t7 plus.t4 source.t0 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 drain_left.t6 plus.t5 source.t2 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X18 source.t23 plus.t6 drain_left.t5 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 source.t10 minus.t9 drain_right.t11 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 source.t4 plus.t7 drain_left.t4 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X21 source.t3 plus.t8 drain_left.t3 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X22 drain_left.t2 plus.t9 source.t20 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 source.t21 plus.t10 drain_left.t1 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X24 drain_right.t9 minus.t10 source.t9 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 source.t8 minus.t11 drain_right.t3 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X26 drain_left.t0 plus.t11 source.t22 a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X27 a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# a_n1878_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 minus.n3 minus.t8 539.035
R1 minus.n17 minus.t11 539.035
R2 minus.n4 minus.t1 512.366
R3 minus.n5 minus.t4 512.366
R4 minus.n1 minus.t9 512.366
R5 minus.n10 minus.t2 512.366
R6 minus.n12 minus.t7 512.366
R7 minus.n18 minus.t10 512.366
R8 minus.n19 minus.t5 512.366
R9 minus.n15 minus.t3 512.366
R10 minus.n24 minus.t0 512.366
R11 minus.n26 minus.t6 512.366
R12 minus.n13 minus.n12 161.3
R13 minus.n11 minus.n0 161.3
R14 minus.n10 minus.n9 161.3
R15 minus.n8 minus.n1 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n2 161.3
R18 minus.n27 minus.n26 161.3
R19 minus.n25 minus.n14 161.3
R20 minus.n24 minus.n23 161.3
R21 minus.n22 minus.n15 161.3
R22 minus.n21 minus.n20 161.3
R23 minus.n19 minus.n16 161.3
R24 minus.n5 minus.n4 48.2005
R25 minus.n10 minus.n1 48.2005
R26 minus.n19 minus.n18 48.2005
R27 minus.n24 minus.n15 48.2005
R28 minus.n12 minus.n11 47.4702
R29 minus.n26 minus.n25 47.4702
R30 minus.n3 minus.n2 45.1192
R31 minus.n17 minus.n16 45.1192
R32 minus.n28 minus.n13 33.9929
R33 minus.n6 minus.n1 24.1005
R34 minus.n6 minus.n5 24.1005
R35 minus.n20 minus.n19 24.1005
R36 minus.n20 minus.n15 24.1005
R37 minus.n4 minus.n3 13.6377
R38 minus.n18 minus.n17 13.6377
R39 minus.n28 minus.n27 6.5308
R40 minus.n11 minus.n10 0.730803
R41 minus.n25 minus.n24 0.730803
R42 minus.n13 minus.n0 0.189894
R43 minus.n9 minus.n0 0.189894
R44 minus.n9 minus.n8 0.189894
R45 minus.n8 minus.n7 0.189894
R46 minus.n7 minus.n2 0.189894
R47 minus.n21 minus.n16 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n14 0.189894
R51 minus.n27 minus.n14 0.189894
R52 minus minus.n28 0.188
R53 drain_right.n6 drain_right.n4 66.2529
R54 drain_right.n3 drain_right.n2 66.1975
R55 drain_right.n3 drain_right.n0 66.1975
R56 drain_right.n6 drain_right.n5 65.5376
R57 drain_right.n8 drain_right.n7 65.5376
R58 drain_right.n3 drain_right.n1 65.5373
R59 drain_right drain_right.n3 28.1187
R60 drain_right drain_right.n8 6.36873
R61 drain_right.n1 drain_right.t8 2.2005
R62 drain_right.n1 drain_right.t2 2.2005
R63 drain_right.n2 drain_right.t4 2.2005
R64 drain_right.n2 drain_right.t0 2.2005
R65 drain_right.n0 drain_right.t3 2.2005
R66 drain_right.n0 drain_right.t9 2.2005
R67 drain_right.n4 drain_right.t10 2.2005
R68 drain_right.n4 drain_right.t7 2.2005
R69 drain_right.n5 drain_right.t11 2.2005
R70 drain_right.n5 drain_right.t6 2.2005
R71 drain_right.n7 drain_right.t5 2.2005
R72 drain_right.n7 drain_right.t1 2.2005
R73 drain_right.n8 drain_right.n6 0.716017
R74 source.n5 source.t5 51.0588
R75 source.n6 source.t11 51.0588
R76 source.n11 source.t12 51.0588
R77 source.n23 source.t13 51.0586
R78 source.n18 source.t8 51.0586
R79 source.n17 source.t2 51.0586
R80 source.n12 source.t7 51.0586
R81 source.n0 source.t22 51.0586
R82 source.n2 source.n1 48.8588
R83 source.n4 source.n3 48.8588
R84 source.n8 source.n7 48.8588
R85 source.n10 source.n9 48.8588
R86 source.n22 source.n21 48.8586
R87 source.n20 source.n19 48.8586
R88 source.n16 source.n15 48.8586
R89 source.n14 source.n13 48.8586
R90 source.n12 source.n11 19.7305
R91 source.n24 source.n0 14.1098
R92 source.n24 source.n23 5.62119
R93 source.n21 source.t16 2.2005
R94 source.n21 source.t19 2.2005
R95 source.n19 source.t9 2.2005
R96 source.n19 source.t14 2.2005
R97 source.n15 source.t1 2.2005
R98 source.n15 source.t23 2.2005
R99 source.n13 source.t20 2.2005
R100 source.n13 source.t3 2.2005
R101 source.n1 source.t6 2.2005
R102 source.n1 source.t4 2.2005
R103 source.n3 source.t0 2.2005
R104 source.n3 source.t21 2.2005
R105 source.n7 source.t15 2.2005
R106 source.n7 source.t18 2.2005
R107 source.n9 source.t17 2.2005
R108 source.n9 source.t10 2.2005
R109 source.n11 source.n10 0.716017
R110 source.n10 source.n8 0.716017
R111 source.n8 source.n6 0.716017
R112 source.n5 source.n4 0.716017
R113 source.n4 source.n2 0.716017
R114 source.n2 source.n0 0.716017
R115 source.n14 source.n12 0.716017
R116 source.n16 source.n14 0.716017
R117 source.n17 source.n16 0.716017
R118 source.n20 source.n18 0.716017
R119 source.n22 source.n20 0.716017
R120 source.n23 source.n22 0.716017
R121 source.n6 source.n5 0.470328
R122 source.n18 source.n17 0.470328
R123 source source.n24 0.188
R124 plus.n5 plus.t1 539.035
R125 plus.n19 plus.t5 539.035
R126 plus.n12 plus.t11 512.366
R127 plus.n10 plus.t7 512.366
R128 plus.n9 plus.t3 512.366
R129 plus.n3 plus.t10 512.366
R130 plus.n4 plus.t4 512.366
R131 plus.n26 plus.t2 512.366
R132 plus.n24 plus.t9 512.366
R133 plus.n23 plus.t8 512.366
R134 plus.n17 plus.t0 512.366
R135 plus.n18 plus.t6 512.366
R136 plus.n6 plus.n3 161.3
R137 plus.n8 plus.n7 161.3
R138 plus.n9 plus.n2 161.3
R139 plus.n10 plus.n1 161.3
R140 plus.n11 plus.n0 161.3
R141 plus.n13 plus.n12 161.3
R142 plus.n20 plus.n17 161.3
R143 plus.n22 plus.n21 161.3
R144 plus.n23 plus.n16 161.3
R145 plus.n24 plus.n15 161.3
R146 plus.n25 plus.n14 161.3
R147 plus.n27 plus.n26 161.3
R148 plus.n10 plus.n9 48.2005
R149 plus.n4 plus.n3 48.2005
R150 plus.n24 plus.n23 48.2005
R151 plus.n18 plus.n17 48.2005
R152 plus.n12 plus.n11 47.4702
R153 plus.n26 plus.n25 47.4702
R154 plus.n6 plus.n5 45.1192
R155 plus.n20 plus.n19 45.1192
R156 plus plus.n27 29.0104
R157 plus.n8 plus.n3 24.1005
R158 plus.n9 plus.n8 24.1005
R159 plus.n23 plus.n22 24.1005
R160 plus.n22 plus.n17 24.1005
R161 plus.n5 plus.n4 13.6377
R162 plus.n19 plus.n18 13.6377
R163 plus plus.n13 11.0384
R164 plus.n11 plus.n10 0.730803
R165 plus.n25 plus.n24 0.730803
R166 plus.n7 plus.n6 0.189894
R167 plus.n7 plus.n2 0.189894
R168 plus.n2 plus.n1 0.189894
R169 plus.n1 plus.n0 0.189894
R170 plus.n13 plus.n0 0.189894
R171 plus.n27 plus.n14 0.189894
R172 plus.n15 plus.n14 0.189894
R173 plus.n16 plus.n15 0.189894
R174 plus.n21 plus.n16 0.189894
R175 plus.n21 plus.n20 0.189894
R176 drain_left.n6 drain_left.n4 66.2531
R177 drain_left.n3 drain_left.n2 66.1975
R178 drain_left.n3 drain_left.n0 66.1975
R179 drain_left.n6 drain_left.n5 65.5376
R180 drain_left.n8 drain_left.n7 65.5374
R181 drain_left.n3 drain_left.n1 65.5373
R182 drain_left drain_left.n3 28.6719
R183 drain_left drain_left.n8 6.36873
R184 drain_left.n1 drain_left.t3 2.2005
R185 drain_left.n1 drain_left.t11 2.2005
R186 drain_left.n2 drain_left.t5 2.2005
R187 drain_left.n2 drain_left.t6 2.2005
R188 drain_left.n0 drain_left.t9 2.2005
R189 drain_left.n0 drain_left.t2 2.2005
R190 drain_left.n7 drain_left.t4 2.2005
R191 drain_left.n7 drain_left.t0 2.2005
R192 drain_left.n5 drain_left.t1 2.2005
R193 drain_left.n5 drain_left.t8 2.2005
R194 drain_left.n4 drain_left.t10 2.2005
R195 drain_left.n4 drain_left.t7 2.2005
R196 drain_left.n8 drain_left.n6 0.716017
C0 source plus 4.87458f
C1 drain_right minus 4.97303f
C2 drain_right drain_left 0.936346f
C3 drain_right source 14.365099f
C4 minus drain_left 0.171641f
C5 minus source 4.86054f
C6 drain_right plus 0.337327f
C7 minus plus 4.93768f
C8 source drain_left 14.3641f
C9 drain_left plus 5.15563f
C10 drain_right a_n1878_n2688# 5.488019f
C11 drain_left a_n1878_n2688# 5.77204f
C12 source a_n1878_n2688# 7.219103f
C13 minus a_n1878_n2688# 7.159318f
C14 plus a_n1878_n2688# 8.81128f
C15 drain_left.t9 a_n1878_n2688# 0.207593f
C16 drain_left.t2 a_n1878_n2688# 0.207593f
C17 drain_left.n0 a_n1878_n2688# 1.8195f
C18 drain_left.t3 a_n1878_n2688# 0.207593f
C19 drain_left.t11 a_n1878_n2688# 0.207593f
C20 drain_left.n1 a_n1878_n2688# 1.81575f
C21 drain_left.t5 a_n1878_n2688# 0.207593f
C22 drain_left.t6 a_n1878_n2688# 0.207593f
C23 drain_left.n2 a_n1878_n2688# 1.8195f
C24 drain_left.n3 a_n1878_n2688# 2.30397f
C25 drain_left.t10 a_n1878_n2688# 0.207593f
C26 drain_left.t7 a_n1878_n2688# 0.207593f
C27 drain_left.n4 a_n1878_n2688# 1.81986f
C28 drain_left.t1 a_n1878_n2688# 0.207593f
C29 drain_left.t8 a_n1878_n2688# 0.207593f
C30 drain_left.n5 a_n1878_n2688# 1.81575f
C31 drain_left.n6 a_n1878_n2688# 0.744442f
C32 drain_left.t4 a_n1878_n2688# 0.207593f
C33 drain_left.t0 a_n1878_n2688# 0.207593f
C34 drain_left.n7 a_n1878_n2688# 1.81574f
C35 drain_left.n8 a_n1878_n2688# 0.619176f
C36 plus.n0 a_n1878_n2688# 0.047589f
C37 plus.t11 a_n1878_n2688# 0.614154f
C38 plus.t7 a_n1878_n2688# 0.614154f
C39 plus.n1 a_n1878_n2688# 0.047589f
C40 plus.t3 a_n1878_n2688# 0.614154f
C41 plus.n2 a_n1878_n2688# 0.047589f
C42 plus.t10 a_n1878_n2688# 0.614154f
C43 plus.n3 a_n1878_n2688# 0.266592f
C44 plus.t4 a_n1878_n2688# 0.614154f
C45 plus.n4 a_n1878_n2688# 0.272328f
C46 plus.t1 a_n1878_n2688# 0.627106f
C47 plus.n5 a_n1878_n2688# 0.249964f
C48 plus.n6 a_n1878_n2688# 0.193813f
C49 plus.n7 a_n1878_n2688# 0.047589f
C50 plus.n8 a_n1878_n2688# 0.010799f
C51 plus.n9 a_n1878_n2688# 0.266592f
C52 plus.n10 a_n1878_n2688# 0.261897f
C53 plus.n11 a_n1878_n2688# 0.010799f
C54 plus.n12 a_n1878_n2688# 0.261604f
C55 plus.n13 a_n1878_n2688# 0.471018f
C56 plus.n14 a_n1878_n2688# 0.047589f
C57 plus.t2 a_n1878_n2688# 0.614154f
C58 plus.n15 a_n1878_n2688# 0.047589f
C59 plus.t9 a_n1878_n2688# 0.614154f
C60 plus.n16 a_n1878_n2688# 0.047589f
C61 plus.t8 a_n1878_n2688# 0.614154f
C62 plus.t0 a_n1878_n2688# 0.614154f
C63 plus.n17 a_n1878_n2688# 0.266592f
C64 plus.t5 a_n1878_n2688# 0.627106f
C65 plus.t6 a_n1878_n2688# 0.614154f
C66 plus.n18 a_n1878_n2688# 0.272328f
C67 plus.n19 a_n1878_n2688# 0.249964f
C68 plus.n20 a_n1878_n2688# 0.193813f
C69 plus.n21 a_n1878_n2688# 0.047589f
C70 plus.n22 a_n1878_n2688# 0.010799f
C71 plus.n23 a_n1878_n2688# 0.266592f
C72 plus.n24 a_n1878_n2688# 0.261897f
C73 plus.n25 a_n1878_n2688# 0.010799f
C74 plus.n26 a_n1878_n2688# 0.261604f
C75 plus.n27 a_n1878_n2688# 1.32957f
C76 source.t22 a_n1878_n2688# 1.81533f
C77 source.n0 a_n1878_n2688# 1.06612f
C78 source.t6 a_n1878_n2688# 0.170239f
C79 source.t4 a_n1878_n2688# 0.170239f
C80 source.n1 a_n1878_n2688# 1.42513f
C81 source.n2 a_n1878_n2688# 0.333467f
C82 source.t0 a_n1878_n2688# 0.170239f
C83 source.t21 a_n1878_n2688# 0.170239f
C84 source.n3 a_n1878_n2688# 1.42513f
C85 source.n4 a_n1878_n2688# 0.333467f
C86 source.t5 a_n1878_n2688# 1.81534f
C87 source.n5 a_n1878_n2688# 0.388593f
C88 source.t11 a_n1878_n2688# 1.81534f
C89 source.n6 a_n1878_n2688# 0.388593f
C90 source.t15 a_n1878_n2688# 0.170239f
C91 source.t18 a_n1878_n2688# 0.170239f
C92 source.n7 a_n1878_n2688# 1.42513f
C93 source.n8 a_n1878_n2688# 0.333467f
C94 source.t17 a_n1878_n2688# 0.170239f
C95 source.t10 a_n1878_n2688# 0.170239f
C96 source.n9 a_n1878_n2688# 1.42513f
C97 source.n10 a_n1878_n2688# 0.333467f
C98 source.t12 a_n1878_n2688# 1.81534f
C99 source.n11 a_n1878_n2688# 1.41826f
C100 source.t7 a_n1878_n2688# 1.81533f
C101 source.n12 a_n1878_n2688# 1.41826f
C102 source.t20 a_n1878_n2688# 0.170239f
C103 source.t3 a_n1878_n2688# 0.170239f
C104 source.n13 a_n1878_n2688# 1.42512f
C105 source.n14 a_n1878_n2688# 0.333472f
C106 source.t1 a_n1878_n2688# 0.170239f
C107 source.t23 a_n1878_n2688# 0.170239f
C108 source.n15 a_n1878_n2688# 1.42512f
C109 source.n16 a_n1878_n2688# 0.333472f
C110 source.t2 a_n1878_n2688# 1.81533f
C111 source.n17 a_n1878_n2688# 0.388598f
C112 source.t8 a_n1878_n2688# 1.81533f
C113 source.n18 a_n1878_n2688# 0.388598f
C114 source.t9 a_n1878_n2688# 0.170239f
C115 source.t14 a_n1878_n2688# 0.170239f
C116 source.n19 a_n1878_n2688# 1.42512f
C117 source.n20 a_n1878_n2688# 0.333472f
C118 source.t16 a_n1878_n2688# 0.170239f
C119 source.t19 a_n1878_n2688# 0.170239f
C120 source.n21 a_n1878_n2688# 1.42512f
C121 source.n22 a_n1878_n2688# 0.333472f
C122 source.t13 a_n1878_n2688# 1.81533f
C123 source.n23 a_n1878_n2688# 0.534287f
C124 source.n24 a_n1878_n2688# 1.25315f
C125 drain_right.t3 a_n1878_n2688# 0.206679f
C126 drain_right.t9 a_n1878_n2688# 0.206679f
C127 drain_right.n0 a_n1878_n2688# 1.81149f
C128 drain_right.t8 a_n1878_n2688# 0.206679f
C129 drain_right.t2 a_n1878_n2688# 0.206679f
C130 drain_right.n1 a_n1878_n2688# 1.80775f
C131 drain_right.t4 a_n1878_n2688# 0.206679f
C132 drain_right.t0 a_n1878_n2688# 0.206679f
C133 drain_right.n2 a_n1878_n2688# 1.81149f
C134 drain_right.n3 a_n1878_n2688# 2.23404f
C135 drain_right.t10 a_n1878_n2688# 0.206679f
C136 drain_right.t7 a_n1878_n2688# 0.206679f
C137 drain_right.n4 a_n1878_n2688# 1.81184f
C138 drain_right.t11 a_n1878_n2688# 0.206679f
C139 drain_right.t6 a_n1878_n2688# 0.206679f
C140 drain_right.n5 a_n1878_n2688# 1.80776f
C141 drain_right.n6 a_n1878_n2688# 0.741171f
C142 drain_right.t5 a_n1878_n2688# 0.206679f
C143 drain_right.t1 a_n1878_n2688# 0.206679f
C144 drain_right.n7 a_n1878_n2688# 1.80776f
C145 drain_right.n8 a_n1878_n2688# 0.616442f
C146 minus.n0 a_n1878_n2688# 0.046655f
C147 minus.t9 a_n1878_n2688# 0.602102f
C148 minus.n1 a_n1878_n2688# 0.26136f
C149 minus.t2 a_n1878_n2688# 0.602102f
C150 minus.n2 a_n1878_n2688# 0.190009f
C151 minus.t8 a_n1878_n2688# 0.614801f
C152 minus.n3 a_n1878_n2688# 0.245059f
C153 minus.t1 a_n1878_n2688# 0.602102f
C154 minus.n4 a_n1878_n2688# 0.266984f
C155 minus.t4 a_n1878_n2688# 0.602102f
C156 minus.n5 a_n1878_n2688# 0.26136f
C157 minus.n6 a_n1878_n2688# 0.010587f
C158 minus.n7 a_n1878_n2688# 0.046655f
C159 minus.n8 a_n1878_n2688# 0.046655f
C160 minus.n9 a_n1878_n2688# 0.046655f
C161 minus.n10 a_n1878_n2688# 0.256758f
C162 minus.n11 a_n1878_n2688# 0.010587f
C163 minus.t7 a_n1878_n2688# 0.602102f
C164 minus.n12 a_n1878_n2688# 0.25647f
C165 minus.n13 a_n1878_n2688# 1.49393f
C166 minus.n14 a_n1878_n2688# 0.046655f
C167 minus.t3 a_n1878_n2688# 0.602102f
C168 minus.n15 a_n1878_n2688# 0.26136f
C169 minus.n16 a_n1878_n2688# 0.190009f
C170 minus.t11 a_n1878_n2688# 0.614801f
C171 minus.n17 a_n1878_n2688# 0.245059f
C172 minus.t10 a_n1878_n2688# 0.602102f
C173 minus.n18 a_n1878_n2688# 0.266984f
C174 minus.t5 a_n1878_n2688# 0.602102f
C175 minus.n19 a_n1878_n2688# 0.26136f
C176 minus.n20 a_n1878_n2688# 0.010587f
C177 minus.n21 a_n1878_n2688# 0.046655f
C178 minus.n22 a_n1878_n2688# 0.046655f
C179 minus.n23 a_n1878_n2688# 0.046655f
C180 minus.t0 a_n1878_n2688# 0.602102f
C181 minus.n24 a_n1878_n2688# 0.256758f
C182 minus.n25 a_n1878_n2688# 0.010587f
C183 minus.t6 a_n1878_n2688# 0.602102f
C184 minus.n26 a_n1878_n2688# 0.25647f
C185 minus.n27 a_n1878_n2688# 0.3084f
C186 minus.n28 a_n1878_n2688# 1.82482f
.ends

