* NGSPICE file created from diffpair528.ext - technology: sky130A

.subckt diffpair528 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t37 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X1 source.t9 plus.t0 drain_left.t19 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X2 drain_left.t18 plus.t1 source.t13 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X3 a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X4 source.t27 minus.t1 drain_right.t18 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X5 source.t7 plus.t2 drain_left.t17 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X6 source.t29 minus.t2 drain_right.t17 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X7 source.t8 plus.t3 drain_left.t16 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X8 source.t19 plus.t4 drain_left.t15 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X9 source.t25 minus.t3 drain_right.t16 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X10 source.t10 plus.t5 drain_left.t14 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X11 drain_left.t13 plus.t6 source.t3 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X12 drain_right.t15 minus.t4 source.t24 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X13 drain_right.t14 minus.t5 source.t31 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X14 source.t20 minus.t6 drain_right.t13 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X15 drain_right.t12 minus.t7 source.t39 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X16 a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X17 drain_left.t12 plus.t7 source.t5 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X18 source.t30 minus.t8 drain_right.t11 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 drain_left.t11 plus.t8 source.t11 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X20 drain_left.t10 plus.t9 source.t14 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X21 source.t0 plus.t10 drain_left.t9 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X22 source.t38 minus.t9 drain_right.t10 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X23 source.t36 minus.t10 drain_right.t9 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X24 drain_right.t8 minus.t11 source.t28 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X25 source.t16 plus.t11 drain_left.t8 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X26 drain_left.t7 plus.t12 source.t2 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X27 source.t1 plus.t13 drain_left.t6 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X28 drain_left.t5 plus.t14 source.t18 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X29 drain_right.t7 minus.t12 source.t26 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X30 drain_right.t6 minus.t13 source.t32 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X31 source.t22 minus.t14 drain_right.t5 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X32 drain_left.t4 plus.t15 source.t4 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X33 drain_right.t4 minus.t15 source.t23 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X34 a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X35 source.t34 minus.t16 drain_right.t3 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X36 source.t33 minus.t17 drain_right.t2 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X37 drain_right.t1 minus.t18 source.t35 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X38 source.t17 plus.t16 drain_left.t3 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X39 drain_left.t2 plus.t17 source.t6 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X40 source.t12 plus.t18 drain_left.t1 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X41 a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X42 drain_right.t0 minus.t19 source.t21 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X43 drain_left.t0 plus.t19 source.t15 a_n2542_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
R0 minus.n6 minus.t12 822.548
R1 minus.n34 minus.t6 822.548
R2 minus.n7 minus.t1 801.567
R3 minus.n5 minus.t7 801.567
R4 minus.n13 minus.t16 801.567
R5 minus.n14 minus.t4 801.567
R6 minus.n18 minus.t9 801.567
R7 minus.n19 minus.t0 801.567
R8 minus.n1 minus.t10 801.567
R9 minus.n25 minus.t15 801.567
R10 minus.n26 minus.t3 801.567
R11 minus.n35 minus.t5 801.567
R12 minus.n33 minus.t14 801.567
R13 minus.n41 minus.t13 801.567
R14 minus.n42 minus.t8 801.567
R15 minus.n46 minus.t18 801.567
R16 minus.n47 minus.t17 801.567
R17 minus.n29 minus.t11 801.567
R18 minus.n53 minus.t2 801.567
R19 minus.n54 minus.t19 801.567
R20 minus.n27 minus.n26 161.3
R21 minus.n25 minus.n0 161.3
R22 minus.n24 minus.n23 161.3
R23 minus.n22 minus.n1 161.3
R24 minus.n21 minus.n20 161.3
R25 minus.n19 minus.n2 161.3
R26 minus.n18 minus.n17 161.3
R27 minus.n16 minus.n3 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n4 161.3
R30 minus.n12 minus.n11 161.3
R31 minus.n10 minus.n5 161.3
R32 minus.n9 minus.n8 161.3
R33 minus.n55 minus.n54 161.3
R34 minus.n53 minus.n28 161.3
R35 minus.n52 minus.n51 161.3
R36 minus.n50 minus.n29 161.3
R37 minus.n49 minus.n48 161.3
R38 minus.n47 minus.n30 161.3
R39 minus.n46 minus.n45 161.3
R40 minus.n44 minus.n31 161.3
R41 minus.n43 minus.n42 161.3
R42 minus.n41 minus.n32 161.3
R43 minus.n40 minus.n39 161.3
R44 minus.n38 minus.n33 161.3
R45 minus.n37 minus.n36 161.3
R46 minus.n9 minus.n6 70.4033
R47 minus.n37 minus.n34 70.4033
R48 minus.n14 minus.n13 48.2005
R49 minus.n19 minus.n18 48.2005
R50 minus.n26 minus.n25 48.2005
R51 minus.n42 minus.n41 48.2005
R52 minus.n47 minus.n46 48.2005
R53 minus.n54 minus.n53 48.2005
R54 minus.n12 minus.n5 47.4702
R55 minus.n20 minus.n1 47.4702
R56 minus.n40 minus.n33 47.4702
R57 minus.n48 minus.n29 47.4702
R58 minus.n56 minus.n27 41.1141
R59 minus.n8 minus.n5 25.5611
R60 minus.n24 minus.n1 25.5611
R61 minus.n36 minus.n33 25.5611
R62 minus.n52 minus.n29 25.5611
R63 minus.n18 minus.n3 24.1005
R64 minus.n14 minus.n3 24.1005
R65 minus.n42 minus.n31 24.1005
R66 minus.n46 minus.n31 24.1005
R67 minus.n8 minus.n7 22.6399
R68 minus.n25 minus.n24 22.6399
R69 minus.n36 minus.n35 22.6399
R70 minus.n53 minus.n52 22.6399
R71 minus.n7 minus.n6 20.9576
R72 minus.n35 minus.n34 20.9576
R73 minus.n56 minus.n55 6.59141
R74 minus.n13 minus.n12 0.730803
R75 minus.n20 minus.n19 0.730803
R76 minus.n41 minus.n40 0.730803
R77 minus.n48 minus.n47 0.730803
R78 minus.n27 minus.n0 0.189894
R79 minus.n23 minus.n0 0.189894
R80 minus.n23 minus.n22 0.189894
R81 minus.n22 minus.n21 0.189894
R82 minus.n21 minus.n2 0.189894
R83 minus.n17 minus.n2 0.189894
R84 minus.n17 minus.n16 0.189894
R85 minus.n16 minus.n15 0.189894
R86 minus.n15 minus.n4 0.189894
R87 minus.n11 minus.n4 0.189894
R88 minus.n11 minus.n10 0.189894
R89 minus.n10 minus.n9 0.189894
R90 minus.n38 minus.n37 0.189894
R91 minus.n39 minus.n38 0.189894
R92 minus.n39 minus.n32 0.189894
R93 minus.n43 minus.n32 0.189894
R94 minus.n44 minus.n43 0.189894
R95 minus.n45 minus.n44 0.189894
R96 minus.n45 minus.n30 0.189894
R97 minus.n49 minus.n30 0.189894
R98 minus.n50 minus.n49 0.189894
R99 minus.n51 minus.n50 0.189894
R100 minus.n51 minus.n28 0.189894
R101 minus.n55 minus.n28 0.189894
R102 minus minus.n56 0.188
R103 source.n9 source.t19 45.521
R104 source.n10 source.t26 45.521
R105 source.n19 source.t25 45.521
R106 source.n39 source.t21 45.5208
R107 source.n30 source.t20 45.5208
R108 source.n29 source.t13 45.5208
R109 source.n20 source.t16 45.5208
R110 source.n0 source.t18 45.5208
R111 source.n2 source.n1 44.201
R112 source.n4 source.n3 44.201
R113 source.n6 source.n5 44.201
R114 source.n8 source.n7 44.201
R115 source.n12 source.n11 44.201
R116 source.n14 source.n13 44.201
R117 source.n16 source.n15 44.201
R118 source.n18 source.n17 44.201
R119 source.n38 source.n37 44.2008
R120 source.n36 source.n35 44.2008
R121 source.n34 source.n33 44.2008
R122 source.n32 source.n31 44.2008
R123 source.n28 source.n27 44.2008
R124 source.n26 source.n25 44.2008
R125 source.n24 source.n23 44.2008
R126 source.n22 source.n21 44.2008
R127 source.n20 source.n19 24.276
R128 source.n40 source.n0 18.6553
R129 source.n40 source.n39 5.62119
R130 source.n37 source.t28 1.3205
R131 source.n37 source.t29 1.3205
R132 source.n35 source.t35 1.3205
R133 source.n35 source.t33 1.3205
R134 source.n33 source.t32 1.3205
R135 source.n33 source.t30 1.3205
R136 source.n31 source.t31 1.3205
R137 source.n31 source.t22 1.3205
R138 source.n27 source.t14 1.3205
R139 source.n27 source.t9 1.3205
R140 source.n25 source.t3 1.3205
R141 source.n25 source.t10 1.3205
R142 source.n23 source.t11 1.3205
R143 source.n23 source.t1 1.3205
R144 source.n21 source.t2 1.3205
R145 source.n21 source.t8 1.3205
R146 source.n1 source.t6 1.3205
R147 source.n1 source.t7 1.3205
R148 source.n3 source.t15 1.3205
R149 source.n3 source.t0 1.3205
R150 source.n5 source.t5 1.3205
R151 source.n5 source.t17 1.3205
R152 source.n7 source.t4 1.3205
R153 source.n7 source.t12 1.3205
R154 source.n11 source.t39 1.3205
R155 source.n11 source.t27 1.3205
R156 source.n13 source.t24 1.3205
R157 source.n13 source.t34 1.3205
R158 source.n15 source.t37 1.3205
R159 source.n15 source.t38 1.3205
R160 source.n17 source.t23 1.3205
R161 source.n17 source.t36 1.3205
R162 source.n19 source.n18 0.716017
R163 source.n18 source.n16 0.716017
R164 source.n16 source.n14 0.716017
R165 source.n14 source.n12 0.716017
R166 source.n12 source.n10 0.716017
R167 source.n9 source.n8 0.716017
R168 source.n8 source.n6 0.716017
R169 source.n6 source.n4 0.716017
R170 source.n4 source.n2 0.716017
R171 source.n2 source.n0 0.716017
R172 source.n22 source.n20 0.716017
R173 source.n24 source.n22 0.716017
R174 source.n26 source.n24 0.716017
R175 source.n28 source.n26 0.716017
R176 source.n29 source.n28 0.716017
R177 source.n32 source.n30 0.716017
R178 source.n34 source.n32 0.716017
R179 source.n36 source.n34 0.716017
R180 source.n38 source.n36 0.716017
R181 source.n39 source.n38 0.716017
R182 source.n10 source.n9 0.470328
R183 source.n30 source.n29 0.470328
R184 source source.n40 0.188
R185 drain_right.n10 drain_right.n8 61.5952
R186 drain_right.n6 drain_right.n4 61.5951
R187 drain_right.n2 drain_right.n0 61.5951
R188 drain_right.n10 drain_right.n9 60.8798
R189 drain_right.n12 drain_right.n11 60.8798
R190 drain_right.n14 drain_right.n13 60.8798
R191 drain_right.n16 drain_right.n15 60.8798
R192 drain_right.n7 drain_right.n3 60.8796
R193 drain_right.n6 drain_right.n5 60.8796
R194 drain_right.n2 drain_right.n1 60.8796
R195 drain_right drain_right.n7 34.8107
R196 drain_right drain_right.n16 6.36873
R197 drain_right.n3 drain_right.t11 1.3205
R198 drain_right.n3 drain_right.t1 1.3205
R199 drain_right.n4 drain_right.t17 1.3205
R200 drain_right.n4 drain_right.t0 1.3205
R201 drain_right.n5 drain_right.t2 1.3205
R202 drain_right.n5 drain_right.t8 1.3205
R203 drain_right.n1 drain_right.t5 1.3205
R204 drain_right.n1 drain_right.t6 1.3205
R205 drain_right.n0 drain_right.t13 1.3205
R206 drain_right.n0 drain_right.t14 1.3205
R207 drain_right.n8 drain_right.t18 1.3205
R208 drain_right.n8 drain_right.t7 1.3205
R209 drain_right.n9 drain_right.t3 1.3205
R210 drain_right.n9 drain_right.t12 1.3205
R211 drain_right.n11 drain_right.t10 1.3205
R212 drain_right.n11 drain_right.t15 1.3205
R213 drain_right.n13 drain_right.t9 1.3205
R214 drain_right.n13 drain_right.t19 1.3205
R215 drain_right.n15 drain_right.t16 1.3205
R216 drain_right.n15 drain_right.t4 1.3205
R217 drain_right.n16 drain_right.n14 0.716017
R218 drain_right.n14 drain_right.n12 0.716017
R219 drain_right.n12 drain_right.n10 0.716017
R220 drain_right.n7 drain_right.n6 0.660671
R221 drain_right.n7 drain_right.n2 0.660671
R222 plus.n8 plus.t4 822.548
R223 plus.n36 plus.t1 822.548
R224 plus.n26 plus.t14 801.567
R225 plus.n25 plus.t2 801.567
R226 plus.n1 plus.t17 801.567
R227 plus.n19 plus.t10 801.567
R228 plus.n18 plus.t19 801.567
R229 plus.n4 plus.t16 801.567
R230 plus.n13 plus.t7 801.567
R231 plus.n11 plus.t18 801.567
R232 plus.n7 plus.t15 801.567
R233 plus.n54 plus.t11 801.567
R234 plus.n53 plus.t12 801.567
R235 plus.n29 plus.t3 801.567
R236 plus.n47 plus.t8 801.567
R237 plus.n46 plus.t13 801.567
R238 plus.n32 plus.t6 801.567
R239 plus.n41 plus.t5 801.567
R240 plus.n39 plus.t9 801.567
R241 plus.n35 plus.t0 801.567
R242 plus.n10 plus.n9 161.3
R243 plus.n11 plus.n6 161.3
R244 plus.n12 plus.n5 161.3
R245 plus.n14 plus.n13 161.3
R246 plus.n15 plus.n4 161.3
R247 plus.n17 plus.n16 161.3
R248 plus.n18 plus.n3 161.3
R249 plus.n19 plus.n2 161.3
R250 plus.n21 plus.n20 161.3
R251 plus.n22 plus.n1 161.3
R252 plus.n24 plus.n23 161.3
R253 plus.n25 plus.n0 161.3
R254 plus.n27 plus.n26 161.3
R255 plus.n38 plus.n37 161.3
R256 plus.n39 plus.n34 161.3
R257 plus.n40 plus.n33 161.3
R258 plus.n42 plus.n41 161.3
R259 plus.n43 plus.n32 161.3
R260 plus.n45 plus.n44 161.3
R261 plus.n46 plus.n31 161.3
R262 plus.n47 plus.n30 161.3
R263 plus.n49 plus.n48 161.3
R264 plus.n50 plus.n29 161.3
R265 plus.n52 plus.n51 161.3
R266 plus.n53 plus.n28 161.3
R267 plus.n55 plus.n54 161.3
R268 plus.n9 plus.n8 70.4033
R269 plus.n37 plus.n36 70.4033
R270 plus.n26 plus.n25 48.2005
R271 plus.n19 plus.n18 48.2005
R272 plus.n13 plus.n4 48.2005
R273 plus.n54 plus.n53 48.2005
R274 plus.n47 plus.n46 48.2005
R275 plus.n41 plus.n32 48.2005
R276 plus.n20 plus.n1 47.4702
R277 plus.n12 plus.n11 47.4702
R278 plus.n48 plus.n29 47.4702
R279 plus.n40 plus.n39 47.4702
R280 plus plus.n55 33.8589
R281 plus.n24 plus.n1 25.5611
R282 plus.n11 plus.n10 25.5611
R283 plus.n52 plus.n29 25.5611
R284 plus.n39 plus.n38 25.5611
R285 plus.n17 plus.n4 24.1005
R286 plus.n18 plus.n17 24.1005
R287 plus.n46 plus.n45 24.1005
R288 plus.n45 plus.n32 24.1005
R289 plus.n25 plus.n24 22.6399
R290 plus.n10 plus.n7 22.6399
R291 plus.n53 plus.n52 22.6399
R292 plus.n38 plus.n35 22.6399
R293 plus.n8 plus.n7 20.9576
R294 plus.n36 plus.n35 20.9576
R295 plus plus.n27 13.3717
R296 plus.n20 plus.n19 0.730803
R297 plus.n13 plus.n12 0.730803
R298 plus.n48 plus.n47 0.730803
R299 plus.n41 plus.n40 0.730803
R300 plus.n9 plus.n6 0.189894
R301 plus.n6 plus.n5 0.189894
R302 plus.n14 plus.n5 0.189894
R303 plus.n15 plus.n14 0.189894
R304 plus.n16 plus.n15 0.189894
R305 plus.n16 plus.n3 0.189894
R306 plus.n3 plus.n2 0.189894
R307 plus.n21 plus.n2 0.189894
R308 plus.n22 plus.n21 0.189894
R309 plus.n23 plus.n22 0.189894
R310 plus.n23 plus.n0 0.189894
R311 plus.n27 plus.n0 0.189894
R312 plus.n55 plus.n28 0.189894
R313 plus.n51 plus.n28 0.189894
R314 plus.n51 plus.n50 0.189894
R315 plus.n50 plus.n49 0.189894
R316 plus.n49 plus.n30 0.189894
R317 plus.n31 plus.n30 0.189894
R318 plus.n44 plus.n31 0.189894
R319 plus.n44 plus.n43 0.189894
R320 plus.n43 plus.n42 0.189894
R321 plus.n42 plus.n33 0.189894
R322 plus.n34 plus.n33 0.189894
R323 plus.n37 plus.n34 0.189894
R324 drain_left.n10 drain_left.n8 61.5953
R325 drain_left.n6 drain_left.n4 61.5951
R326 drain_left.n2 drain_left.n0 61.5951
R327 drain_left.n14 drain_left.n13 60.8798
R328 drain_left.n12 drain_left.n11 60.8798
R329 drain_left.n10 drain_left.n9 60.8798
R330 drain_left.n16 drain_left.n15 60.8796
R331 drain_left.n7 drain_left.n3 60.8796
R332 drain_left.n6 drain_left.n5 60.8796
R333 drain_left.n2 drain_left.n1 60.8796
R334 drain_left drain_left.n7 35.3639
R335 drain_left drain_left.n16 6.36873
R336 drain_left.n3 drain_left.t6 1.3205
R337 drain_left.n3 drain_left.t13 1.3205
R338 drain_left.n4 drain_left.t19 1.3205
R339 drain_left.n4 drain_left.t18 1.3205
R340 drain_left.n5 drain_left.t14 1.3205
R341 drain_left.n5 drain_left.t10 1.3205
R342 drain_left.n1 drain_left.t16 1.3205
R343 drain_left.n1 drain_left.t11 1.3205
R344 drain_left.n0 drain_left.t8 1.3205
R345 drain_left.n0 drain_left.t7 1.3205
R346 drain_left.n15 drain_left.t17 1.3205
R347 drain_left.n15 drain_left.t5 1.3205
R348 drain_left.n13 drain_left.t9 1.3205
R349 drain_left.n13 drain_left.t2 1.3205
R350 drain_left.n11 drain_left.t3 1.3205
R351 drain_left.n11 drain_left.t0 1.3205
R352 drain_left.n9 drain_left.t1 1.3205
R353 drain_left.n9 drain_left.t12 1.3205
R354 drain_left.n8 drain_left.t15 1.3205
R355 drain_left.n8 drain_left.t4 1.3205
R356 drain_left.n12 drain_left.n10 0.716017
R357 drain_left.n14 drain_left.n12 0.716017
R358 drain_left.n16 drain_left.n14 0.716017
R359 drain_left.n7 drain_left.n6 0.660671
R360 drain_left.n7 drain_left.n2 0.660671
C0 drain_right plus 0.40825f
C1 drain_right minus 12.6451f
C2 drain_right drain_left 1.35855f
C3 source drain_right 35.0103f
C4 minus plus 6.87554f
C5 drain_left plus 12.896901f
C6 drain_left minus 0.173163f
C7 source plus 12.518499f
C8 source minus 12.5044f
C9 source drain_left 35.009f
C10 drain_right a_n2542_n3888# 7.60571f
C11 drain_left a_n2542_n3888# 7.97499f
C12 source a_n2542_n3888# 10.775897f
C13 minus a_n2542_n3888# 10.321439f
C14 plus a_n2542_n3888# 12.404641f
C15 drain_left.t8 a_n2542_n3888# 0.349309f
C16 drain_left.t7 a_n2542_n3888# 0.349309f
C17 drain_left.n0 a_n2542_n3888# 3.16186f
C18 drain_left.t16 a_n2542_n3888# 0.349309f
C19 drain_left.t11 a_n2542_n3888# 0.349309f
C20 drain_left.n1 a_n2542_n3888# 3.15734f
C21 drain_left.n2 a_n2542_n3888# 0.757635f
C22 drain_left.t6 a_n2542_n3888# 0.349309f
C23 drain_left.t13 a_n2542_n3888# 0.349309f
C24 drain_left.n3 a_n2542_n3888# 3.15734f
C25 drain_left.t19 a_n2542_n3888# 0.349309f
C26 drain_left.t18 a_n2542_n3888# 0.349309f
C27 drain_left.n4 a_n2542_n3888# 3.16186f
C28 drain_left.t14 a_n2542_n3888# 0.349309f
C29 drain_left.t10 a_n2542_n3888# 0.349309f
C30 drain_left.n5 a_n2542_n3888# 3.15734f
C31 drain_left.n6 a_n2542_n3888# 0.757635f
C32 drain_left.n7 a_n2542_n3888# 2.19264f
C33 drain_left.t15 a_n2542_n3888# 0.349309f
C34 drain_left.t4 a_n2542_n3888# 0.349309f
C35 drain_left.n8 a_n2542_n3888# 3.16187f
C36 drain_left.t1 a_n2542_n3888# 0.349309f
C37 drain_left.t12 a_n2542_n3888# 0.349309f
C38 drain_left.n9 a_n2542_n3888# 3.15735f
C39 drain_left.n10 a_n2542_n3888# 0.761851f
C40 drain_left.t3 a_n2542_n3888# 0.349309f
C41 drain_left.t0 a_n2542_n3888# 0.349309f
C42 drain_left.n11 a_n2542_n3888# 3.15735f
C43 drain_left.n12 a_n2542_n3888# 0.377251f
C44 drain_left.t9 a_n2542_n3888# 0.349309f
C45 drain_left.t2 a_n2542_n3888# 0.349309f
C46 drain_left.n13 a_n2542_n3888# 3.15735f
C47 drain_left.n14 a_n2542_n3888# 0.377251f
C48 drain_left.t17 a_n2542_n3888# 0.349309f
C49 drain_left.t5 a_n2542_n3888# 0.349309f
C50 drain_left.n15 a_n2542_n3888# 3.15733f
C51 drain_left.n16 a_n2542_n3888# 0.630441f
C52 plus.n0 a_n2542_n3888# 0.044605f
C53 plus.t14 a_n2542_n3888# 0.950653f
C54 plus.t2 a_n2542_n3888# 0.950653f
C55 plus.t17 a_n2542_n3888# 0.950653f
C56 plus.n1 a_n2542_n3888# 0.375016f
C57 plus.n2 a_n2542_n3888# 0.044605f
C58 plus.t10 a_n2542_n3888# 0.950653f
C59 plus.t19 a_n2542_n3888# 0.950653f
C60 plus.n3 a_n2542_n3888# 0.044605f
C61 plus.t16 a_n2542_n3888# 0.950653f
C62 plus.n4 a_n2542_n3888# 0.374878f
C63 plus.n5 a_n2542_n3888# 0.044605f
C64 plus.t7 a_n2542_n3888# 0.950653f
C65 plus.t18 a_n2542_n3888# 0.950653f
C66 plus.n6 a_n2542_n3888# 0.044605f
C67 plus.t15 a_n2542_n3888# 0.950653f
C68 plus.n7 a_n2542_n3888# 0.374603f
C69 plus.t4 a_n2542_n3888# 0.960101f
C70 plus.n8 a_n2542_n3888# 0.361234f
C71 plus.n9 a_n2542_n3888# 0.146398f
C72 plus.n10 a_n2542_n3888# 0.010122f
C73 plus.n11 a_n2542_n3888# 0.375016f
C74 plus.n12 a_n2542_n3888# 0.010122f
C75 plus.n13 a_n2542_n3888# 0.370478f
C76 plus.n14 a_n2542_n3888# 0.044605f
C77 plus.n15 a_n2542_n3888# 0.044605f
C78 plus.n16 a_n2542_n3888# 0.044605f
C79 plus.n17 a_n2542_n3888# 0.010122f
C80 plus.n18 a_n2542_n3888# 0.374878f
C81 plus.n19 a_n2542_n3888# 0.370478f
C82 plus.n20 a_n2542_n3888# 0.010122f
C83 plus.n21 a_n2542_n3888# 0.044605f
C84 plus.n22 a_n2542_n3888# 0.044605f
C85 plus.n23 a_n2542_n3888# 0.044605f
C86 plus.n24 a_n2542_n3888# 0.010122f
C87 plus.n25 a_n2542_n3888# 0.374603f
C88 plus.n26 a_n2542_n3888# 0.370341f
C89 plus.n27 a_n2542_n3888# 0.573249f
C90 plus.n28 a_n2542_n3888# 0.044605f
C91 plus.t11 a_n2542_n3888# 0.950653f
C92 plus.t12 a_n2542_n3888# 0.950653f
C93 plus.t3 a_n2542_n3888# 0.950653f
C94 plus.n29 a_n2542_n3888# 0.375016f
C95 plus.n30 a_n2542_n3888# 0.044605f
C96 plus.t8 a_n2542_n3888# 0.950653f
C97 plus.n31 a_n2542_n3888# 0.044605f
C98 plus.t13 a_n2542_n3888# 0.950653f
C99 plus.t6 a_n2542_n3888# 0.950653f
C100 plus.n32 a_n2542_n3888# 0.374878f
C101 plus.n33 a_n2542_n3888# 0.044605f
C102 plus.t5 a_n2542_n3888# 0.950653f
C103 plus.n34 a_n2542_n3888# 0.044605f
C104 plus.t9 a_n2542_n3888# 0.950653f
C105 plus.t0 a_n2542_n3888# 0.950653f
C106 plus.n35 a_n2542_n3888# 0.374603f
C107 plus.t1 a_n2542_n3888# 0.960101f
C108 plus.n36 a_n2542_n3888# 0.361234f
C109 plus.n37 a_n2542_n3888# 0.146398f
C110 plus.n38 a_n2542_n3888# 0.010122f
C111 plus.n39 a_n2542_n3888# 0.375016f
C112 plus.n40 a_n2542_n3888# 0.010122f
C113 plus.n41 a_n2542_n3888# 0.370478f
C114 plus.n42 a_n2542_n3888# 0.044605f
C115 plus.n43 a_n2542_n3888# 0.044605f
C116 plus.n44 a_n2542_n3888# 0.044605f
C117 plus.n45 a_n2542_n3888# 0.010122f
C118 plus.n46 a_n2542_n3888# 0.374878f
C119 plus.n47 a_n2542_n3888# 0.370478f
C120 plus.n48 a_n2542_n3888# 0.010122f
C121 plus.n49 a_n2542_n3888# 0.044605f
C122 plus.n50 a_n2542_n3888# 0.044605f
C123 plus.n51 a_n2542_n3888# 0.044605f
C124 plus.n52 a_n2542_n3888# 0.010122f
C125 plus.n53 a_n2542_n3888# 0.374603f
C126 plus.n54 a_n2542_n3888# 0.370341f
C127 plus.n55 a_n2542_n3888# 1.59148f
C128 drain_right.t13 a_n2542_n3888# 0.347959f
C129 drain_right.t14 a_n2542_n3888# 0.347959f
C130 drain_right.n0 a_n2542_n3888# 3.14964f
C131 drain_right.t5 a_n2542_n3888# 0.347959f
C132 drain_right.t6 a_n2542_n3888# 0.347959f
C133 drain_right.n1 a_n2542_n3888# 3.14514f
C134 drain_right.n2 a_n2542_n3888# 0.754706f
C135 drain_right.t11 a_n2542_n3888# 0.347959f
C136 drain_right.t1 a_n2542_n3888# 0.347959f
C137 drain_right.n3 a_n2542_n3888# 3.14514f
C138 drain_right.t17 a_n2542_n3888# 0.347959f
C139 drain_right.t0 a_n2542_n3888# 0.347959f
C140 drain_right.n4 a_n2542_n3888# 3.14964f
C141 drain_right.t2 a_n2542_n3888# 0.347959f
C142 drain_right.t8 a_n2542_n3888# 0.347959f
C143 drain_right.n5 a_n2542_n3888# 3.14514f
C144 drain_right.n6 a_n2542_n3888# 0.754706f
C145 drain_right.n7 a_n2542_n3888# 2.12374f
C146 drain_right.t18 a_n2542_n3888# 0.347959f
C147 drain_right.t7 a_n2542_n3888# 0.347959f
C148 drain_right.n8 a_n2542_n3888# 3.14963f
C149 drain_right.t3 a_n2542_n3888# 0.347959f
C150 drain_right.t12 a_n2542_n3888# 0.347959f
C151 drain_right.n9 a_n2542_n3888# 3.14514f
C152 drain_right.n10 a_n2542_n3888# 0.758916f
C153 drain_right.t10 a_n2542_n3888# 0.347959f
C154 drain_right.t15 a_n2542_n3888# 0.347959f
C155 drain_right.n11 a_n2542_n3888# 3.14514f
C156 drain_right.n12 a_n2542_n3888# 0.375792f
C157 drain_right.t9 a_n2542_n3888# 0.347959f
C158 drain_right.t19 a_n2542_n3888# 0.347959f
C159 drain_right.n13 a_n2542_n3888# 3.14514f
C160 drain_right.n14 a_n2542_n3888# 0.375792f
C161 drain_right.t16 a_n2542_n3888# 0.347959f
C162 drain_right.t4 a_n2542_n3888# 0.347959f
C163 drain_right.n15 a_n2542_n3888# 3.14514f
C164 drain_right.n16 a_n2542_n3888# 0.627993f
C165 source.t18 a_n2542_n3888# 3.38512f
C166 source.n0 a_n2542_n3888# 1.59075f
C167 source.t6 a_n2542_n3888# 0.302065f
C168 source.t7 a_n2542_n3888# 0.302065f
C169 source.n1 a_n2542_n3888# 2.65339f
C170 source.n2 a_n2542_n3888# 0.36852f
C171 source.t15 a_n2542_n3888# 0.302065f
C172 source.t0 a_n2542_n3888# 0.302065f
C173 source.n3 a_n2542_n3888# 2.65339f
C174 source.n4 a_n2542_n3888# 0.36852f
C175 source.t5 a_n2542_n3888# 0.302065f
C176 source.t17 a_n2542_n3888# 0.302065f
C177 source.n5 a_n2542_n3888# 2.65339f
C178 source.n6 a_n2542_n3888# 0.36852f
C179 source.t4 a_n2542_n3888# 0.302065f
C180 source.t12 a_n2542_n3888# 0.302065f
C181 source.n7 a_n2542_n3888# 2.65339f
C182 source.n8 a_n2542_n3888# 0.36852f
C183 source.t19 a_n2542_n3888# 3.38513f
C184 source.n9 a_n2542_n3888# 0.440418f
C185 source.t26 a_n2542_n3888# 3.38513f
C186 source.n10 a_n2542_n3888# 0.440418f
C187 source.t39 a_n2542_n3888# 0.302065f
C188 source.t27 a_n2542_n3888# 0.302065f
C189 source.n11 a_n2542_n3888# 2.65339f
C190 source.n12 a_n2542_n3888# 0.36852f
C191 source.t24 a_n2542_n3888# 0.302065f
C192 source.t34 a_n2542_n3888# 0.302065f
C193 source.n13 a_n2542_n3888# 2.65339f
C194 source.n14 a_n2542_n3888# 0.36852f
C195 source.t37 a_n2542_n3888# 0.302065f
C196 source.t38 a_n2542_n3888# 0.302065f
C197 source.n15 a_n2542_n3888# 2.65339f
C198 source.n16 a_n2542_n3888# 0.36852f
C199 source.t23 a_n2542_n3888# 0.302065f
C200 source.t36 a_n2542_n3888# 0.302065f
C201 source.n17 a_n2542_n3888# 2.65339f
C202 source.n18 a_n2542_n3888# 0.36852f
C203 source.t25 a_n2542_n3888# 3.38513f
C204 source.n19 a_n2542_n3888# 2.01992f
C205 source.t16 a_n2542_n3888# 3.38513f
C206 source.n20 a_n2542_n3888# 2.01992f
C207 source.t2 a_n2542_n3888# 0.302065f
C208 source.t8 a_n2542_n3888# 0.302065f
C209 source.n21 a_n2542_n3888# 2.65338f
C210 source.n22 a_n2542_n3888# 0.368523f
C211 source.t11 a_n2542_n3888# 0.302065f
C212 source.t1 a_n2542_n3888# 0.302065f
C213 source.n23 a_n2542_n3888# 2.65338f
C214 source.n24 a_n2542_n3888# 0.368523f
C215 source.t3 a_n2542_n3888# 0.302065f
C216 source.t10 a_n2542_n3888# 0.302065f
C217 source.n25 a_n2542_n3888# 2.65338f
C218 source.n26 a_n2542_n3888# 0.368523f
C219 source.t14 a_n2542_n3888# 0.302065f
C220 source.t9 a_n2542_n3888# 0.302065f
C221 source.n27 a_n2542_n3888# 2.65338f
C222 source.n28 a_n2542_n3888# 0.368523f
C223 source.t13 a_n2542_n3888# 3.38513f
C224 source.n29 a_n2542_n3888# 0.440422f
C225 source.t20 a_n2542_n3888# 3.38513f
C226 source.n30 a_n2542_n3888# 0.440422f
C227 source.t31 a_n2542_n3888# 0.302065f
C228 source.t22 a_n2542_n3888# 0.302065f
C229 source.n31 a_n2542_n3888# 2.65338f
C230 source.n32 a_n2542_n3888# 0.368523f
C231 source.t32 a_n2542_n3888# 0.302065f
C232 source.t30 a_n2542_n3888# 0.302065f
C233 source.n33 a_n2542_n3888# 2.65338f
C234 source.n34 a_n2542_n3888# 0.368523f
C235 source.t35 a_n2542_n3888# 0.302065f
C236 source.t33 a_n2542_n3888# 0.302065f
C237 source.n35 a_n2542_n3888# 2.65338f
C238 source.n36 a_n2542_n3888# 0.368523f
C239 source.t28 a_n2542_n3888# 0.302065f
C240 source.t29 a_n2542_n3888# 0.302065f
C241 source.n37 a_n2542_n3888# 2.65338f
C242 source.n38 a_n2542_n3888# 0.368523f
C243 source.t21 a_n2542_n3888# 3.38513f
C244 source.n39 a_n2542_n3888# 0.595526f
C245 source.n40 a_n2542_n3888# 1.87169f
C246 minus.n0 a_n2542_n3888# 0.044068f
C247 minus.t10 a_n2542_n3888# 0.939201f
C248 minus.n1 a_n2542_n3888# 0.370498f
C249 minus.n2 a_n2542_n3888# 0.044068f
C250 minus.n3 a_n2542_n3888# 0.01f
C251 minus.t9 a_n2542_n3888# 0.939201f
C252 minus.n4 a_n2542_n3888# 0.044068f
C253 minus.t7 a_n2542_n3888# 0.939201f
C254 minus.n5 a_n2542_n3888# 0.370498f
C255 minus.t12 a_n2542_n3888# 0.948535f
C256 minus.n6 a_n2542_n3888# 0.356883f
C257 minus.t1 a_n2542_n3888# 0.939201f
C258 minus.n7 a_n2542_n3888# 0.370091f
C259 minus.n8 a_n2542_n3888# 0.01f
C260 minus.n9 a_n2542_n3888# 0.144634f
C261 minus.n10 a_n2542_n3888# 0.044068f
C262 minus.n11 a_n2542_n3888# 0.044068f
C263 minus.n12 a_n2542_n3888# 0.01f
C264 minus.t16 a_n2542_n3888# 0.939201f
C265 minus.n13 a_n2542_n3888# 0.366015f
C266 minus.t4 a_n2542_n3888# 0.939201f
C267 minus.n14 a_n2542_n3888# 0.370362f
C268 minus.n15 a_n2542_n3888# 0.044068f
C269 minus.n16 a_n2542_n3888# 0.044068f
C270 minus.n17 a_n2542_n3888# 0.044068f
C271 minus.n18 a_n2542_n3888# 0.370362f
C272 minus.t0 a_n2542_n3888# 0.939201f
C273 minus.n19 a_n2542_n3888# 0.366015f
C274 minus.n20 a_n2542_n3888# 0.01f
C275 minus.n21 a_n2542_n3888# 0.044068f
C276 minus.n22 a_n2542_n3888# 0.044068f
C277 minus.n23 a_n2542_n3888# 0.044068f
C278 minus.n24 a_n2542_n3888# 0.01f
C279 minus.t15 a_n2542_n3888# 0.939201f
C280 minus.n25 a_n2542_n3888# 0.370091f
C281 minus.t3 a_n2542_n3888# 0.939201f
C282 minus.n26 a_n2542_n3888# 0.365879f
C283 minus.n27 a_n2542_n3888# 1.89378f
C284 minus.n28 a_n2542_n3888# 0.044068f
C285 minus.t11 a_n2542_n3888# 0.939201f
C286 minus.n29 a_n2542_n3888# 0.370498f
C287 minus.n30 a_n2542_n3888# 0.044068f
C288 minus.n31 a_n2542_n3888# 0.01f
C289 minus.n32 a_n2542_n3888# 0.044068f
C290 minus.t14 a_n2542_n3888# 0.939201f
C291 minus.n33 a_n2542_n3888# 0.370498f
C292 minus.t6 a_n2542_n3888# 0.948535f
C293 minus.n34 a_n2542_n3888# 0.356883f
C294 minus.t5 a_n2542_n3888# 0.939201f
C295 minus.n35 a_n2542_n3888# 0.370091f
C296 minus.n36 a_n2542_n3888# 0.01f
C297 minus.n37 a_n2542_n3888# 0.144634f
C298 minus.n38 a_n2542_n3888# 0.044068f
C299 minus.n39 a_n2542_n3888# 0.044068f
C300 minus.n40 a_n2542_n3888# 0.01f
C301 minus.t13 a_n2542_n3888# 0.939201f
C302 minus.n41 a_n2542_n3888# 0.366015f
C303 minus.t8 a_n2542_n3888# 0.939201f
C304 minus.n42 a_n2542_n3888# 0.370362f
C305 minus.n43 a_n2542_n3888# 0.044068f
C306 minus.n44 a_n2542_n3888# 0.044068f
C307 minus.n45 a_n2542_n3888# 0.044068f
C308 minus.t18 a_n2542_n3888# 0.939201f
C309 minus.n46 a_n2542_n3888# 0.370362f
C310 minus.t17 a_n2542_n3888# 0.939201f
C311 minus.n47 a_n2542_n3888# 0.366015f
C312 minus.n48 a_n2542_n3888# 0.01f
C313 minus.n49 a_n2542_n3888# 0.044068f
C314 minus.n50 a_n2542_n3888# 0.044068f
C315 minus.n51 a_n2542_n3888# 0.044068f
C316 minus.n52 a_n2542_n3888# 0.01f
C317 minus.t2 a_n2542_n3888# 0.939201f
C318 minus.n53 a_n2542_n3888# 0.370091f
C319 minus.t19 a_n2542_n3888# 0.939201f
C320 minus.n54 a_n2542_n3888# 0.365879f
C321 minus.n55 a_n2542_n3888# 0.297551f
C322 minus.n56 a_n2542_n3888# 2.26492f
.ends

