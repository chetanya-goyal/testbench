* NGSPICE file created from diffpair553.ext - technology: sky130A

.subckt diffpair553 minus drain_right drain_left source plus
X0 a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X1 drain_left.t7 plus.t0 source.t13 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X2 source.t3 minus.t0 drain_right.t7 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X3 a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X4 a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X5 drain_right.t6 minus.t1 source.t4 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X6 drain_right.t5 minus.t2 source.t1 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X7 source.t7 plus.t1 drain_left.t6 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X8 source.t0 minus.t3 drain_right.t4 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X9 source.t8 plus.t2 drain_left.t5 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 drain_right.t3 minus.t4 source.t6 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X11 drain_right.t2 minus.t5 source.t5 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X12 source.t15 minus.t6 drain_right.t1 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X13 drain_left.t4 plus.t3 source.t14 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X14 a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X15 source.t10 plus.t4 drain_left.t3 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X16 drain_left.t2 plus.t5 source.t9 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X17 drain_left.t1 plus.t6 source.t11 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X18 source.t12 plus.t7 drain_left.t0 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X19 source.t2 minus.t7 drain_right.t0 a_n1846_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n2 plus.t7 521.582
R1 plus.n10 plus.t0 521.582
R2 plus.n6 plus.t3 500.979
R3 plus.n4 plus.t4 500.979
R4 plus.n3 plus.t5 500.979
R5 plus.n14 plus.t1 500.979
R6 plus.n12 plus.t6 500.979
R7 plus.n11 plus.t2 500.979
R8 plus.n5 plus.n0 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n13 plus.n8 161.3
R11 plus.n15 plus.n14 161.3
R12 plus.n4 plus.n1 80.6037
R13 plus.n12 plus.n9 80.6037
R14 plus.n4 plus.n3 48.2005
R15 plus.n12 plus.n11 48.2005
R16 plus.n5 plus.n4 41.6278
R17 plus.n13 plus.n12 41.6278
R18 plus.n2 plus.n1 31.6158
R19 plus.n10 plus.n9 31.6158
R20 plus plus.n15 31.2831
R21 plus.n3 plus.n2 17.6494
R22 plus.n11 plus.n10 17.6494
R23 plus plus.n7 13.4323
R24 plus.n6 plus.n5 6.57323
R25 plus.n14 plus.n13 6.57323
R26 plus.n1 plus.n0 0.285035
R27 plus.n9 plus.n8 0.285035
R28 plus.n7 plus.n0 0.189894
R29 plus.n15 plus.n8 0.189894
R30 source.n3 source.t12 45.521
R31 source.n4 source.t6 45.521
R32 source.n7 source.t15 45.521
R33 source.n15 source.t1 45.5208
R34 source.n12 source.t3 45.5208
R35 source.n11 source.t13 45.5208
R36 source.n8 source.t7 45.5208
R37 source.n0 source.t14 45.5208
R38 source.n2 source.n1 44.201
R39 source.n6 source.n5 44.201
R40 source.n14 source.n13 44.2008
R41 source.n10 source.n9 44.2008
R42 source.n8 source.n7 24.5346
R43 source.n16 source.n0 18.7846
R44 source.n16 source.n15 5.7505
R45 source.n13 source.t5 1.3205
R46 source.n13 source.t2 1.3205
R47 source.n9 source.t11 1.3205
R48 source.n9 source.t8 1.3205
R49 source.n1 source.t9 1.3205
R50 source.n1 source.t10 1.3205
R51 source.n5 source.t4 1.3205
R52 source.n5 source.t0 1.3205
R53 source.n7 source.n6 0.974638
R54 source.n6 source.n4 0.974638
R55 source.n3 source.n2 0.974638
R56 source.n2 source.n0 0.974638
R57 source.n10 source.n8 0.974638
R58 source.n11 source.n10 0.974638
R59 source.n14 source.n12 0.974638
R60 source.n15 source.n14 0.974638
R61 source.n4 source.n3 0.470328
R62 source.n12 source.n11 0.470328
R63 source source.n16 0.188
R64 drain_left.n5 drain_left.n3 61.8539
R65 drain_left.n2 drain_left.n1 61.3113
R66 drain_left.n2 drain_left.n0 61.3113
R67 drain_left.n5 drain_left.n4 60.8796
R68 drain_left drain_left.n2 33.0493
R69 drain_left drain_left.n5 6.62735
R70 drain_left.n1 drain_left.t5 1.3205
R71 drain_left.n1 drain_left.t7 1.3205
R72 drain_left.n0 drain_left.t6 1.3205
R73 drain_left.n0 drain_left.t1 1.3205
R74 drain_left.n4 drain_left.t3 1.3205
R75 drain_left.n4 drain_left.t4 1.3205
R76 drain_left.n3 drain_left.t0 1.3205
R77 drain_left.n3 drain_left.t2 1.3205
R78 minus.n2 minus.t4 521.582
R79 minus.n10 minus.t0 521.582
R80 minus.n1 minus.t3 500.979
R81 minus.n4 minus.t1 500.979
R82 minus.n6 minus.t6 500.979
R83 minus.n9 minus.t5 500.979
R84 minus.n12 minus.t7 500.979
R85 minus.n14 minus.t2 500.979
R86 minus.n7 minus.n6 161.3
R87 minus.n5 minus.n0 161.3
R88 minus.n15 minus.n14 161.3
R89 minus.n13 minus.n8 161.3
R90 minus.n4 minus.n3 80.6037
R91 minus.n12 minus.n11 80.6037
R92 minus.n4 minus.n1 48.2005
R93 minus.n12 minus.n9 48.2005
R94 minus.n5 minus.n4 41.6278
R95 minus.n13 minus.n12 41.6278
R96 minus.n16 minus.n7 38.5384
R97 minus.n3 minus.n2 31.6158
R98 minus.n11 minus.n10 31.6158
R99 minus.n2 minus.n1 17.6494
R100 minus.n10 minus.n9 17.6494
R101 minus.n16 minus.n15 6.65202
R102 minus.n6 minus.n5 6.57323
R103 minus.n14 minus.n13 6.57323
R104 minus.n3 minus.n0 0.285035
R105 minus.n11 minus.n8 0.285035
R106 minus.n7 minus.n0 0.189894
R107 minus.n15 minus.n8 0.189894
R108 minus minus.n16 0.188
R109 drain_right.n5 drain_right.n3 61.8538
R110 drain_right.n2 drain_right.n1 61.3113
R111 drain_right.n2 drain_right.n0 61.3113
R112 drain_right.n5 drain_right.n4 60.8798
R113 drain_right drain_right.n2 32.4961
R114 drain_right drain_right.n5 6.62735
R115 drain_right.n1 drain_right.t0 1.3205
R116 drain_right.n1 drain_right.t5 1.3205
R117 drain_right.n0 drain_right.t7 1.3205
R118 drain_right.n0 drain_right.t2 1.3205
R119 drain_right.n3 drain_right.t4 1.3205
R120 drain_right.n3 drain_right.t3 1.3205
R121 drain_right.n4 drain_right.t1 1.3205
R122 drain_right.n4 drain_right.t6 1.3205
C0 minus drain_left 0.17159f
C1 drain_right drain_left 0.873724f
C2 drain_left plus 7.46229f
C3 source drain_left 12.6908f
C4 minus drain_right 7.28304f
C5 minus plus 5.99881f
C6 source minus 6.95504f
C7 drain_right plus 0.333957f
C8 source drain_right 12.6932f
C9 source plus 6.96908f
C10 drain_right a_n1846_n3888# 6.30103f
C11 drain_left a_n1846_n3888# 6.57209f
C12 source a_n1846_n3888# 10.779258f
C13 minus a_n1846_n3888# 7.359093f
C14 plus a_n1846_n3888# 9.14303f
C15 drain_right.t7 a_n1846_n3888# 0.315163f
C16 drain_right.t2 a_n1846_n3888# 0.315163f
C17 drain_right.n0 a_n1846_n3888# 2.85117f
C18 drain_right.t0 a_n1846_n3888# 0.315163f
C19 drain_right.t5 a_n1846_n3888# 0.315163f
C20 drain_right.n1 a_n1846_n3888# 2.85117f
C21 drain_right.n2 a_n1846_n3888# 2.16262f
C22 drain_right.t4 a_n1846_n3888# 0.315163f
C23 drain_right.t3 a_n1846_n3888# 0.315163f
C24 drain_right.n3 a_n1846_n3888# 2.85492f
C25 drain_right.t1 a_n1846_n3888# 0.315163f
C26 drain_right.t6 a_n1846_n3888# 0.315163f
C27 drain_right.n4 a_n1846_n3888# 2.84871f
C28 drain_right.n5 a_n1846_n3888# 1.01228f
C29 minus.n0 a_n1846_n3888# 0.055643f
C30 minus.t3 a_n1846_n3888# 1.42197f
C31 minus.n1 a_n1846_n3888# 0.557256f
C32 minus.t1 a_n1846_n3888# 1.42197f
C33 minus.t4 a_n1846_n3888# 1.44364f
C34 minus.n2 a_n1846_n3888# 0.530531f
C35 minus.n3 a_n1846_n3888# 0.238661f
C36 minus.n4 a_n1846_n3888# 0.556577f
C37 minus.n5 a_n1846_n3888# 0.009462f
C38 minus.t6 a_n1846_n3888# 1.42197f
C39 minus.n6 a_n1846_n3888# 0.540944f
C40 minus.n7 a_n1846_n3888# 1.62816f
C41 minus.n8 a_n1846_n3888# 0.055643f
C42 minus.t5 a_n1846_n3888# 1.42197f
C43 minus.n9 a_n1846_n3888# 0.557256f
C44 minus.t0 a_n1846_n3888# 1.44364f
C45 minus.n10 a_n1846_n3888# 0.530531f
C46 minus.n11 a_n1846_n3888# 0.238661f
C47 minus.t7 a_n1846_n3888# 1.42197f
C48 minus.n12 a_n1846_n3888# 0.556577f
C49 minus.n13 a_n1846_n3888# 0.009462f
C50 minus.t2 a_n1846_n3888# 1.42197f
C51 minus.n14 a_n1846_n3888# 0.540944f
C52 minus.n15 a_n1846_n3888# 0.287449f
C53 minus.n16 a_n1846_n3888# 1.95975f
C54 drain_left.t6 a_n1846_n3888# 0.316668f
C55 drain_left.t1 a_n1846_n3888# 0.316668f
C56 drain_left.n0 a_n1846_n3888# 2.86478f
C57 drain_left.t5 a_n1846_n3888# 0.316668f
C58 drain_left.t7 a_n1846_n3888# 0.316668f
C59 drain_left.n1 a_n1846_n3888# 2.86478f
C60 drain_left.n2 a_n1846_n3888# 2.22857f
C61 drain_left.t0 a_n1846_n3888# 0.316668f
C62 drain_left.t2 a_n1846_n3888# 0.316668f
C63 drain_left.n3 a_n1846_n3888# 2.86856f
C64 drain_left.t3 a_n1846_n3888# 0.316668f
C65 drain_left.t4 a_n1846_n3888# 0.316668f
C66 drain_left.n4 a_n1846_n3888# 2.8623f
C67 drain_left.n5 a_n1846_n3888# 1.01712f
C68 source.t14 a_n1846_n3888# 2.56922f
C69 source.n0 a_n1846_n3888# 1.23331f
C70 source.t9 a_n1846_n3888# 0.229259f
C71 source.t10 a_n1846_n3888# 0.229259f
C72 source.n1 a_n1846_n3888# 2.01385f
C73 source.n2 a_n1846_n3888# 0.311932f
C74 source.t12 a_n1846_n3888# 2.56922f
C75 source.n3 a_n1846_n3888# 0.350383f
C76 source.t6 a_n1846_n3888# 2.56922f
C77 source.n4 a_n1846_n3888# 0.350383f
C78 source.t4 a_n1846_n3888# 0.229259f
C79 source.t0 a_n1846_n3888# 0.229259f
C80 source.n5 a_n1846_n3888# 2.01385f
C81 source.n6 a_n1846_n3888# 0.311932f
C82 source.t15 a_n1846_n3888# 2.56922f
C83 source.n7 a_n1846_n3888# 1.5653f
C84 source.t7 a_n1846_n3888# 2.56922f
C85 source.n8 a_n1846_n3888# 1.5653f
C86 source.t11 a_n1846_n3888# 0.229259f
C87 source.t8 a_n1846_n3888# 0.229259f
C88 source.n9 a_n1846_n3888# 2.01385f
C89 source.n10 a_n1846_n3888# 0.311934f
C90 source.t13 a_n1846_n3888# 2.56922f
C91 source.n11 a_n1846_n3888# 0.350386f
C92 source.t3 a_n1846_n3888# 2.56922f
C93 source.n12 a_n1846_n3888# 0.350386f
C94 source.t5 a_n1846_n3888# 0.229259f
C95 source.t2 a_n1846_n3888# 0.229259f
C96 source.n13 a_n1846_n3888# 2.01385f
C97 source.n14 a_n1846_n3888# 0.311934f
C98 source.t1 a_n1846_n3888# 2.56922f
C99 source.n15 a_n1846_n3888# 0.480736f
C100 source.n16 a_n1846_n3888# 1.43032f
C101 plus.n0 a_n1846_n3888# 0.056425f
C102 plus.t3 a_n1846_n3888# 1.44197f
C103 plus.t4 a_n1846_n3888# 1.44197f
C104 plus.n1 a_n1846_n3888# 0.242017f
C105 plus.t5 a_n1846_n3888# 1.44197f
C106 plus.t7 a_n1846_n3888# 1.46395f
C107 plus.n2 a_n1846_n3888# 0.537993f
C108 plus.n3 a_n1846_n3888# 0.565094f
C109 plus.n4 a_n1846_n3888# 0.564405f
C110 plus.n5 a_n1846_n3888# 0.009596f
C111 plus.n6 a_n1846_n3888# 0.548553f
C112 plus.n7 a_n1846_n3888# 0.549451f
C113 plus.n8 a_n1846_n3888# 0.056425f
C114 plus.t1 a_n1846_n3888# 1.44197f
C115 plus.n9 a_n1846_n3888# 0.242017f
C116 plus.t6 a_n1846_n3888# 1.44197f
C117 plus.t0 a_n1846_n3888# 1.46395f
C118 plus.n10 a_n1846_n3888# 0.537993f
C119 plus.t2 a_n1846_n3888# 1.44197f
C120 plus.n11 a_n1846_n3888# 0.565094f
C121 plus.n12 a_n1846_n3888# 0.564405f
C122 plus.n13 a_n1846_n3888# 0.009596f
C123 plus.n14 a_n1846_n3888# 0.548553f
C124 plus.n15 a_n1846_n3888# 1.36088f
.ends

