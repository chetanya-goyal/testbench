* NGSPICE file created from diffpair571.ext - technology: sky130A

.subckt diffpair571 minus drain_right drain_left source plus
X0 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X1 drain_right minus source a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X2 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X3 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X4 a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X5 drain_left plus source a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X6 source plus drain_left a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X7 drain_left plus source a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X8 source minus drain_right a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X9 source minus drain_right a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X10 drain_right minus source a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X11 source plus drain_left a_n1034_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
.ends

