* NGSPICE file created from diffpair569.ext - technology: sky130A

.subckt diffpair569 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t5 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X1 source.t46 minus.t1 drain_right.t4 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 drain_right.t1 minus.t2 source.t45 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X3 source.t0 plus.t0 drain_left.t23 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X4 drain_right.t0 minus.t3 source.t44 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X5 source.t43 minus.t4 drain_right.t7 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X6 source.t15 plus.t1 drain_left.t22 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X7 drain_left.t21 plus.t2 source.t19 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X8 drain_left.t20 plus.t3 source.t23 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X9 a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X10 drain_left.t19 plus.t4 source.t16 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source.t1 plus.t5 drain_left.t18 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X13 source.t5 plus.t6 drain_left.t17 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X14 source.t42 minus.t5 drain_right.t6 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 drain_right.t9 minus.t6 source.t41 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X16 source.t6 plus.t7 drain_left.t16 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_right.t8 minus.t7 source.t40 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X18 drain_right.t23 minus.t8 source.t39 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 drain_left.t15 plus.t8 source.t11 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X20 source.t38 minus.t9 drain_right.t22 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 source.t37 minus.t10 drain_right.t21 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X23 drain_right.t20 minus.t11 source.t36 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X24 source.t35 minus.t12 drain_right.t13 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X25 drain_left.t14 plus.t9 source.t8 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X26 drain_left.t13 plus.t10 source.t2 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 source.t10 plus.t11 drain_left.t12 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X28 drain_right.t12 minus.t13 source.t34 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X29 drain_right.t17 minus.t14 source.t33 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X30 source.t13 plus.t12 drain_left.t11 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X31 source.t32 minus.t15 drain_right.t16 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X32 source.t31 minus.t16 drain_right.t15 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X33 drain_right.t14 minus.t17 source.t30 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X34 drain_left.t10 plus.t13 source.t18 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X35 drain_left.t9 plus.t14 source.t20 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X36 source.t29 minus.t18 drain_right.t19 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X37 drain_right.t18 minus.t19 source.t28 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X38 drain_right.t11 minus.t20 source.t27 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X39 drain_left.t8 plus.t15 source.t12 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X40 source.t17 plus.t16 drain_left.t7 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X41 source.t21 plus.t17 drain_left.t6 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X42 drain_right.t10 minus.t21 source.t26 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X43 source.t22 plus.t18 drain_left.t5 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X44 source.t25 minus.t22 drain_right.t3 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X45 source.t4 plus.t19 drain_left.t4 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X46 drain_left.t3 plus.t20 source.t9 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X47 drain_left.t2 plus.t21 source.t3 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X48 source.t24 minus.t23 drain_right.t2 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X49 a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X50 drain_left.t1 plus.t22 source.t7 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X51 source.t14 plus.t23 drain_left.t0 a_n2406_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n35 minus.t16 3469.67
R1 minus.n8 minus.t7 3469.67
R2 minus.n72 minus.t6 3469.67
R3 minus.n43 minus.t4 3469.67
R4 minus.n34 minus.t19 3422.2
R5 minus.n32 minus.t22 3422.2
R6 minus.n3 minus.t11 3422.2
R7 minus.n26 minus.t15 3422.2
R8 minus.n24 minus.t14 3422.2
R9 minus.n6 minus.t18 3422.2
R10 minus.n18 minus.t8 3422.2
R11 minus.n16 minus.t10 3422.2
R12 minus.n9 minus.t13 3422.2
R13 minus.n10 minus.t5 3422.2
R14 minus.n71 minus.t1 3422.2
R15 minus.n69 minus.t21 3422.2
R16 minus.n63 minus.t12 3422.2
R17 minus.n62 minus.t3 3422.2
R18 minus.n60 minus.t0 3422.2
R19 minus.n54 minus.t20 3422.2
R20 minus.n53 minus.t9 3422.2
R21 minus.n51 minus.t2 3422.2
R22 minus.n45 minus.t23 3422.2
R23 minus.n44 minus.t17 3422.2
R24 minus.n12 minus.n8 161.489
R25 minus.n47 minus.n43 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n31 minus.n30 161.3
R29 minus.n29 minus.n1 161.3
R30 minus.n28 minus.n27 161.3
R31 minus.n25 minus.n2 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n20 minus.n19 161.3
R35 minus.n17 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n7 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n68 minus.n67 161.3
R42 minus.n66 minus.n38 161.3
R43 minus.n65 minus.n64 161.3
R44 minus.n61 minus.n39 161.3
R45 minus.n59 minus.n58 161.3
R46 minus.n57 minus.n40 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n52 minus.n41 161.3
R49 minus.n50 minus.n49 161.3
R50 minus.n48 minus.n42 161.3
R51 minus.n47 minus.n46 161.3
R52 minus.n31 minus.n1 73.0308
R53 minus.n23 minus.n4 73.0308
R54 minus.n15 minus.n7 73.0308
R55 minus.n50 minus.n42 73.0308
R56 minus.n59 minus.n40 73.0308
R57 minus.n68 minus.n38 73.0308
R58 minus.n33 minus.n32 69.3793
R59 minus.n11 minus.n9 69.3793
R60 minus.n46 minus.n45 69.3793
R61 minus.n70 minus.n69 69.3793
R62 minus.n25 minus.n24 62.0763
R63 minus.n19 minus.n6 62.0763
R64 minus.n55 minus.n54 62.0763
R65 minus.n61 minus.n60 62.0763
R66 minus.n27 minus.n3 54.7732
R67 minus.n17 minus.n16 54.7732
R68 minus.n52 minus.n51 54.7732
R69 minus.n64 minus.n63 54.7732
R70 minus.n35 minus.n34 47.4702
R71 minus.n10 minus.n8 47.4702
R72 minus.n44 minus.n43 47.4702
R73 minus.n72 minus.n71 47.4702
R74 minus.n74 minus.n36 44.3187
R75 minus.n27 minus.n26 40.1672
R76 minus.n18 minus.n17 40.1672
R77 minus.n53 minus.n52 40.1672
R78 minus.n64 minus.n62 40.1672
R79 minus.n26 minus.n25 32.8641
R80 minus.n19 minus.n18 32.8641
R81 minus.n55 minus.n53 32.8641
R82 minus.n62 minus.n61 32.8641
R83 minus.n34 minus.n33 25.5611
R84 minus.n11 minus.n10 25.5611
R85 minus.n46 minus.n44 25.5611
R86 minus.n71 minus.n70 25.5611
R87 minus.n3 minus.n1 18.2581
R88 minus.n16 minus.n15 18.2581
R89 minus.n51 minus.n50 18.2581
R90 minus.n63 minus.n38 18.2581
R91 minus.n24 minus.n23 10.955
R92 minus.n6 minus.n4 10.955
R93 minus.n54 minus.n40 10.955
R94 minus.n60 minus.n59 10.955
R95 minus.n74 minus.n73 6.52323
R96 minus.n32 minus.n31 3.65202
R97 minus.n9 minus.n7 3.65202
R98 minus.n45 minus.n42 3.65202
R99 minus.n69 minus.n68 3.65202
R100 minus.n36 minus.n0 0.189894
R101 minus.n30 minus.n0 0.189894
R102 minus.n30 minus.n29 0.189894
R103 minus.n29 minus.n28 0.189894
R104 minus.n28 minus.n2 0.189894
R105 minus.n22 minus.n2 0.189894
R106 minus.n22 minus.n21 0.189894
R107 minus.n21 minus.n20 0.189894
R108 minus.n20 minus.n5 0.189894
R109 minus.n14 minus.n5 0.189894
R110 minus.n14 minus.n13 0.189894
R111 minus.n13 minus.n12 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n49 minus.n48 0.189894
R114 minus.n49 minus.n41 0.189894
R115 minus.n56 minus.n41 0.189894
R116 minus.n57 minus.n56 0.189894
R117 minus.n58 minus.n57 0.189894
R118 minus.n58 minus.n39 0.189894
R119 minus.n65 minus.n39 0.189894
R120 minus.n66 minus.n65 0.189894
R121 minus.n67 minus.n66 0.189894
R122 minus.n67 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 drain_right.n13 drain_right.n11 60.3788
R126 drain_right.n7 drain_right.n5 60.3788
R127 drain_right.n2 drain_right.n0 60.3788
R128 drain_right.n13 drain_right.n12 59.8185
R129 drain_right.n15 drain_right.n14 59.8185
R130 drain_right.n17 drain_right.n16 59.8185
R131 drain_right.n19 drain_right.n18 59.8185
R132 drain_right.n21 drain_right.n20 59.8185
R133 drain_right.n7 drain_right.n6 59.8184
R134 drain_right.n9 drain_right.n8 59.8184
R135 drain_right.n4 drain_right.n3 59.8184
R136 drain_right.n2 drain_right.n1 59.8184
R137 drain_right drain_right.n10 38.1977
R138 drain_right drain_right.n21 6.21356
R139 drain_right.n5 drain_right.t4 1.5005
R140 drain_right.n5 drain_right.t9 1.5005
R141 drain_right.n6 drain_right.t13 1.5005
R142 drain_right.n6 drain_right.t10 1.5005
R143 drain_right.n8 drain_right.t5 1.5005
R144 drain_right.n8 drain_right.t0 1.5005
R145 drain_right.n3 drain_right.t22 1.5005
R146 drain_right.n3 drain_right.t11 1.5005
R147 drain_right.n1 drain_right.t2 1.5005
R148 drain_right.n1 drain_right.t1 1.5005
R149 drain_right.n0 drain_right.t7 1.5005
R150 drain_right.n0 drain_right.t14 1.5005
R151 drain_right.n11 drain_right.t6 1.5005
R152 drain_right.n11 drain_right.t8 1.5005
R153 drain_right.n12 drain_right.t21 1.5005
R154 drain_right.n12 drain_right.t12 1.5005
R155 drain_right.n14 drain_right.t19 1.5005
R156 drain_right.n14 drain_right.t23 1.5005
R157 drain_right.n16 drain_right.t16 1.5005
R158 drain_right.n16 drain_right.t17 1.5005
R159 drain_right.n18 drain_right.t3 1.5005
R160 drain_right.n18 drain_right.t20 1.5005
R161 drain_right.n20 drain_right.t15 1.5005
R162 drain_right.n20 drain_right.t18 1.5005
R163 drain_right.n9 drain_right.n7 0.560845
R164 drain_right.n4 drain_right.n2 0.560845
R165 drain_right.n21 drain_right.n19 0.560845
R166 drain_right.n19 drain_right.n17 0.560845
R167 drain_right.n17 drain_right.n15 0.560845
R168 drain_right.n15 drain_right.n13 0.560845
R169 drain_right.n10 drain_right.n9 0.225326
R170 drain_right.n10 drain_right.n4 0.225326
R171 source.n0 source.t7 44.6397
R172 source.n11 source.t10 44.6396
R173 source.n12 source.t40 44.6396
R174 source.n23 source.t31 44.6396
R175 source.n47 source.t41 44.6395
R176 source.n36 source.t43 44.6395
R177 source.n35 source.t8 44.6395
R178 source.n24 source.t5 44.6395
R179 source.n2 source.n1 43.1397
R180 source.n4 source.n3 43.1397
R181 source.n6 source.n5 43.1397
R182 source.n8 source.n7 43.1397
R183 source.n10 source.n9 43.1397
R184 source.n14 source.n13 43.1397
R185 source.n16 source.n15 43.1397
R186 source.n18 source.n17 43.1397
R187 source.n20 source.n19 43.1397
R188 source.n22 source.n21 43.1397
R189 source.n46 source.n45 43.1396
R190 source.n44 source.n43 43.1396
R191 source.n42 source.n41 43.1396
R192 source.n40 source.n39 43.1396
R193 source.n38 source.n37 43.1396
R194 source.n34 source.n33 43.1396
R195 source.n32 source.n31 43.1396
R196 source.n30 source.n29 43.1396
R197 source.n28 source.n27 43.1396
R198 source.n26 source.n25 43.1396
R199 source.n24 source.n23 27.9087
R200 source.n48 source.n0 22.3656
R201 source.n48 source.n47 5.5436
R202 source.n45 source.t26 1.5005
R203 source.n45 source.t46 1.5005
R204 source.n43 source.t44 1.5005
R205 source.n43 source.t35 1.5005
R206 source.n41 source.t27 1.5005
R207 source.n41 source.t47 1.5005
R208 source.n39 source.t45 1.5005
R209 source.n39 source.t38 1.5005
R210 source.n37 source.t30 1.5005
R211 source.n37 source.t24 1.5005
R212 source.n33 source.t23 1.5005
R213 source.n33 source.t22 1.5005
R214 source.n31 source.t18 1.5005
R215 source.n31 source.t6 1.5005
R216 source.n29 source.t16 1.5005
R217 source.n29 source.t15 1.5005
R218 source.n27 source.t11 1.5005
R219 source.n27 source.t1 1.5005
R220 source.n25 source.t19 1.5005
R221 source.n25 source.t0 1.5005
R222 source.n1 source.t12 1.5005
R223 source.n1 source.t13 1.5005
R224 source.n3 source.t2 1.5005
R225 source.n3 source.t4 1.5005
R226 source.n5 source.t9 1.5005
R227 source.n5 source.t17 1.5005
R228 source.n7 source.t20 1.5005
R229 source.n7 source.t14 1.5005
R230 source.n9 source.t3 1.5005
R231 source.n9 source.t21 1.5005
R232 source.n13 source.t34 1.5005
R233 source.n13 source.t42 1.5005
R234 source.n15 source.t39 1.5005
R235 source.n15 source.t37 1.5005
R236 source.n17 source.t33 1.5005
R237 source.n17 source.t29 1.5005
R238 source.n19 source.t36 1.5005
R239 source.n19 source.t32 1.5005
R240 source.n21 source.t28 1.5005
R241 source.n21 source.t25 1.5005
R242 source.n23 source.n22 0.560845
R243 source.n22 source.n20 0.560845
R244 source.n20 source.n18 0.560845
R245 source.n18 source.n16 0.560845
R246 source.n16 source.n14 0.560845
R247 source.n14 source.n12 0.560845
R248 source.n11 source.n10 0.560845
R249 source.n10 source.n8 0.560845
R250 source.n8 source.n6 0.560845
R251 source.n6 source.n4 0.560845
R252 source.n4 source.n2 0.560845
R253 source.n2 source.n0 0.560845
R254 source.n26 source.n24 0.560845
R255 source.n28 source.n26 0.560845
R256 source.n30 source.n28 0.560845
R257 source.n32 source.n30 0.560845
R258 source.n34 source.n32 0.560845
R259 source.n35 source.n34 0.560845
R260 source.n38 source.n36 0.560845
R261 source.n40 source.n38 0.560845
R262 source.n42 source.n40 0.560845
R263 source.n44 source.n42 0.560845
R264 source.n46 source.n44 0.560845
R265 source.n47 source.n46 0.560845
R266 source.n12 source.n11 0.470328
R267 source.n36 source.n35 0.470328
R268 source source.n48 0.188
R269 plus.n6 plus.t11 3469.67
R270 plus.n35 plus.t22 3469.67
R271 plus.n45 plus.t9 3469.67
R272 plus.n72 plus.t6 3469.67
R273 plus.n7 plus.t21 3422.2
R274 plus.n8 plus.t17 3422.2
R275 plus.n14 plus.t14 3422.2
R276 plus.n16 plus.t23 3422.2
R277 plus.n17 plus.t20 3422.2
R278 plus.n23 plus.t16 3422.2
R279 plus.n25 plus.t10 3422.2
R280 plus.n26 plus.t19 3422.2
R281 plus.n32 plus.t15 3422.2
R282 plus.n34 plus.t12 3422.2
R283 plus.n47 plus.t18 3422.2
R284 plus.n46 plus.t3 3422.2
R285 plus.n53 plus.t7 3422.2
R286 plus.n55 plus.t13 3422.2
R287 plus.n43 plus.t1 3422.2
R288 plus.n61 plus.t4 3422.2
R289 plus.n63 plus.t5 3422.2
R290 plus.n40 plus.t8 3422.2
R291 plus.n69 plus.t0 3422.2
R292 plus.n71 plus.t2 3422.2
R293 plus.n10 plus.n6 161.489
R294 plus.n49 plus.n45 161.489
R295 plus.n10 plus.n9 161.3
R296 plus.n11 plus.n5 161.3
R297 plus.n13 plus.n12 161.3
R298 plus.n15 plus.n4 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n3 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n24 plus.n2 161.3
R303 plus.n28 plus.n27 161.3
R304 plus.n29 plus.n1 161.3
R305 plus.n31 plus.n30 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n49 plus.n48 161.3
R309 plus.n50 plus.n44 161.3
R310 plus.n52 plus.n51 161.3
R311 plus.n54 plus.n42 161.3
R312 plus.n57 plus.n56 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n39 161.3
R316 plus.n65 plus.n64 161.3
R317 plus.n66 plus.n38 161.3
R318 plus.n68 plus.n67 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n13 plus.n5 73.0308
R322 plus.n22 plus.n3 73.0308
R323 plus.n31 plus.n1 73.0308
R324 plus.n68 plus.n38 73.0308
R325 plus.n60 plus.n41 73.0308
R326 plus.n52 plus.n44 73.0308
R327 plus.n9 plus.n8 69.3793
R328 plus.n33 plus.n32 69.3793
R329 plus.n70 plus.n69 69.3793
R330 plus.n48 plus.n46 69.3793
R331 plus.n18 plus.n17 62.0763
R332 plus.n24 plus.n23 62.0763
R333 plus.n62 plus.n61 62.0763
R334 plus.n56 plus.n43 62.0763
R335 plus.n15 plus.n14 54.7732
R336 plus.n27 plus.n26 54.7732
R337 plus.n64 plus.n40 54.7732
R338 plus.n54 plus.n53 54.7732
R339 plus.n7 plus.n6 47.4702
R340 plus.n35 plus.n34 47.4702
R341 plus.n72 plus.n71 47.4702
R342 plus.n47 plus.n45 47.4702
R343 plus.n16 plus.n15 40.1672
R344 plus.n27 plus.n25 40.1672
R345 plus.n64 plus.n63 40.1672
R346 plus.n55 plus.n54 40.1672
R347 plus plus.n73 35.1695
R348 plus.n18 plus.n16 32.8641
R349 plus.n25 plus.n24 32.8641
R350 plus.n63 plus.n62 32.8641
R351 plus.n56 plus.n55 32.8641
R352 plus.n9 plus.n7 25.5611
R353 plus.n34 plus.n33 25.5611
R354 plus.n71 plus.n70 25.5611
R355 plus.n48 plus.n47 25.5611
R356 plus.n14 plus.n13 18.2581
R357 plus.n26 plus.n1 18.2581
R358 plus.n40 plus.n38 18.2581
R359 plus.n53 plus.n52 18.2581
R360 plus plus.n36 15.1975
R361 plus.n17 plus.n3 10.955
R362 plus.n23 plus.n22 10.955
R363 plus.n61 plus.n60 10.955
R364 plus.n43 plus.n41 10.955
R365 plus.n8 plus.n5 3.65202
R366 plus.n32 plus.n31 3.65202
R367 plus.n69 plus.n68 3.65202
R368 plus.n46 plus.n44 3.65202
R369 plus.n11 plus.n10 0.189894
R370 plus.n12 plus.n11 0.189894
R371 plus.n12 plus.n4 0.189894
R372 plus.n19 plus.n4 0.189894
R373 plus.n20 plus.n19 0.189894
R374 plus.n21 plus.n20 0.189894
R375 plus.n21 plus.n2 0.189894
R376 plus.n28 plus.n2 0.189894
R377 plus.n29 plus.n28 0.189894
R378 plus.n30 plus.n29 0.189894
R379 plus.n30 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n67 plus.n37 0.189894
R383 plus.n67 plus.n66 0.189894
R384 plus.n66 plus.n65 0.189894
R385 plus.n65 plus.n39 0.189894
R386 plus.n59 plus.n39 0.189894
R387 plus.n59 plus.n58 0.189894
R388 plus.n58 plus.n57 0.189894
R389 plus.n57 plus.n42 0.189894
R390 plus.n51 plus.n42 0.189894
R391 plus.n51 plus.n50 0.189894
R392 plus.n50 plus.n49 0.189894
R393 drain_left.n13 drain_left.n11 60.3788
R394 drain_left.n7 drain_left.n5 60.3788
R395 drain_left.n2 drain_left.n0 60.3788
R396 drain_left.n21 drain_left.n20 59.8185
R397 drain_left.n19 drain_left.n18 59.8185
R398 drain_left.n17 drain_left.n16 59.8185
R399 drain_left.n15 drain_left.n14 59.8185
R400 drain_left.n13 drain_left.n12 59.8185
R401 drain_left.n7 drain_left.n6 59.8184
R402 drain_left.n9 drain_left.n8 59.8184
R403 drain_left.n4 drain_left.n3 59.8184
R404 drain_left.n2 drain_left.n1 59.8184
R405 drain_left drain_left.n10 38.751
R406 drain_left drain_left.n21 6.21356
R407 drain_left.n5 drain_left.t5 1.5005
R408 drain_left.n5 drain_left.t14 1.5005
R409 drain_left.n6 drain_left.t16 1.5005
R410 drain_left.n6 drain_left.t20 1.5005
R411 drain_left.n8 drain_left.t22 1.5005
R412 drain_left.n8 drain_left.t10 1.5005
R413 drain_left.n3 drain_left.t18 1.5005
R414 drain_left.n3 drain_left.t19 1.5005
R415 drain_left.n1 drain_left.t23 1.5005
R416 drain_left.n1 drain_left.t15 1.5005
R417 drain_left.n0 drain_left.t17 1.5005
R418 drain_left.n0 drain_left.t21 1.5005
R419 drain_left.n20 drain_left.t11 1.5005
R420 drain_left.n20 drain_left.t1 1.5005
R421 drain_left.n18 drain_left.t4 1.5005
R422 drain_left.n18 drain_left.t8 1.5005
R423 drain_left.n16 drain_left.t7 1.5005
R424 drain_left.n16 drain_left.t13 1.5005
R425 drain_left.n14 drain_left.t0 1.5005
R426 drain_left.n14 drain_left.t3 1.5005
R427 drain_left.n12 drain_left.t6 1.5005
R428 drain_left.n12 drain_left.t9 1.5005
R429 drain_left.n11 drain_left.t12 1.5005
R430 drain_left.n11 drain_left.t2 1.5005
R431 drain_left.n9 drain_left.n7 0.560845
R432 drain_left.n4 drain_left.n2 0.560845
R433 drain_left.n15 drain_left.n13 0.560845
R434 drain_left.n17 drain_left.n15 0.560845
R435 drain_left.n19 drain_left.n17 0.560845
R436 drain_left.n21 drain_left.n19 0.560845
R437 drain_left.n10 drain_left.n9 0.225326
R438 drain_left.n10 drain_left.n4 0.225326
C0 source drain_right 73.0208f
C1 drain_left drain_right 1.29455f
C2 source drain_left 73.0201f
C3 plus drain_right 0.392113f
C4 source plus 6.91584f
C5 drain_left plus 7.94982f
C6 minus drain_right 7.71204f
C7 source minus 6.9018f
C8 drain_left minus 0.171476f
C9 plus minus 7.62299f
C10 drain_right a_n2406_n4888# 8.30529f
C11 drain_left a_n2406_n4888# 8.65024f
C12 source a_n2406_n4888# 13.311848f
C13 minus a_n2406_n4888# 9.453521f
C14 plus a_n2406_n4888# 12.198931f
C15 drain_left.t17 a_n2406_n4888# 0.675935f
C16 drain_left.t21 a_n2406_n4888# 0.675935f
C17 drain_left.n0 a_n2406_n4888# 4.5414f
C18 drain_left.t23 a_n2406_n4888# 0.675935f
C19 drain_left.t15 a_n2406_n4888# 0.675935f
C20 drain_left.n1 a_n2406_n4888# 4.53814f
C21 drain_left.n2 a_n2406_n4888# 0.68836f
C22 drain_left.t18 a_n2406_n4888# 0.675935f
C23 drain_left.t19 a_n2406_n4888# 0.675935f
C24 drain_left.n3 a_n2406_n4888# 4.53814f
C25 drain_left.n4 a_n2406_n4888# 0.312521f
C26 drain_left.t5 a_n2406_n4888# 0.675935f
C27 drain_left.t14 a_n2406_n4888# 0.675935f
C28 drain_left.n5 a_n2406_n4888# 4.5414f
C29 drain_left.t16 a_n2406_n4888# 0.675935f
C30 drain_left.t20 a_n2406_n4888# 0.675935f
C31 drain_left.n6 a_n2406_n4888# 4.53814f
C32 drain_left.n7 a_n2406_n4888# 0.68836f
C33 drain_left.t22 a_n2406_n4888# 0.675935f
C34 drain_left.t10 a_n2406_n4888# 0.675935f
C35 drain_left.n8 a_n2406_n4888# 4.53814f
C36 drain_left.n9 a_n2406_n4888# 0.312521f
C37 drain_left.n10 a_n2406_n4888# 2.10266f
C38 drain_left.t12 a_n2406_n4888# 0.675935f
C39 drain_left.t2 a_n2406_n4888# 0.675935f
C40 drain_left.n11 a_n2406_n4888# 4.54139f
C41 drain_left.t6 a_n2406_n4888# 0.675935f
C42 drain_left.t9 a_n2406_n4888# 0.675935f
C43 drain_left.n12 a_n2406_n4888# 4.53813f
C44 drain_left.n13 a_n2406_n4888# 0.688372f
C45 drain_left.t0 a_n2406_n4888# 0.675935f
C46 drain_left.t3 a_n2406_n4888# 0.675935f
C47 drain_left.n14 a_n2406_n4888# 4.53813f
C48 drain_left.n15 a_n2406_n4888# 0.340132f
C49 drain_left.t7 a_n2406_n4888# 0.675935f
C50 drain_left.t13 a_n2406_n4888# 0.675935f
C51 drain_left.n16 a_n2406_n4888# 4.53813f
C52 drain_left.n17 a_n2406_n4888# 0.340132f
C53 drain_left.t4 a_n2406_n4888# 0.675935f
C54 drain_left.t8 a_n2406_n4888# 0.675935f
C55 drain_left.n18 a_n2406_n4888# 4.53813f
C56 drain_left.n19 a_n2406_n4888# 0.340132f
C57 drain_left.t11 a_n2406_n4888# 0.675935f
C58 drain_left.t1 a_n2406_n4888# 0.675935f
C59 drain_left.n20 a_n2406_n4888# 4.53813f
C60 drain_left.n21 a_n2406_n4888# 0.575858f
C61 plus.n0 a_n2406_n4888# 0.052164f
C62 plus.t12 a_n2406_n4888# 0.440757f
C63 plus.t15 a_n2406_n4888# 0.440757f
C64 plus.n1 a_n2406_n4888# 0.021325f
C65 plus.n2 a_n2406_n4888# 0.052164f
C66 plus.t10 a_n2406_n4888# 0.440757f
C67 plus.t16 a_n2406_n4888# 0.440757f
C68 plus.n3 a_n2406_n4888# 0.019717f
C69 plus.n4 a_n2406_n4888# 0.052164f
C70 plus.t23 a_n2406_n4888# 0.440757f
C71 plus.t14 a_n2406_n4888# 0.440757f
C72 plus.n5 a_n2406_n4888# 0.018108f
C73 plus.t11 a_n2406_n4888# 0.443096f
C74 plus.n6 a_n2406_n4888# 0.190829f
C75 plus.t21 a_n2406_n4888# 0.440757f
C76 plus.n7 a_n2406_n4888# 0.171771f
C77 plus.t17 a_n2406_n4888# 0.440757f
C78 plus.n8 a_n2406_n4888# 0.171771f
C79 plus.n9 a_n2406_n4888# 0.022129f
C80 plus.n10 a_n2406_n4888# 0.113904f
C81 plus.n11 a_n2406_n4888# 0.052164f
C82 plus.n12 a_n2406_n4888# 0.052164f
C83 plus.n13 a_n2406_n4888# 0.021325f
C84 plus.n14 a_n2406_n4888# 0.171771f
C85 plus.n15 a_n2406_n4888# 0.022129f
C86 plus.n16 a_n2406_n4888# 0.171771f
C87 plus.t20 a_n2406_n4888# 0.440757f
C88 plus.n17 a_n2406_n4888# 0.171771f
C89 plus.n18 a_n2406_n4888# 0.022129f
C90 plus.n19 a_n2406_n4888# 0.052164f
C91 plus.n20 a_n2406_n4888# 0.052164f
C92 plus.n21 a_n2406_n4888# 0.052164f
C93 plus.n22 a_n2406_n4888# 0.019717f
C94 plus.n23 a_n2406_n4888# 0.171771f
C95 plus.n24 a_n2406_n4888# 0.022129f
C96 plus.n25 a_n2406_n4888# 0.171771f
C97 plus.t19 a_n2406_n4888# 0.440757f
C98 plus.n26 a_n2406_n4888# 0.171771f
C99 plus.n27 a_n2406_n4888# 0.022129f
C100 plus.n28 a_n2406_n4888# 0.052164f
C101 plus.n29 a_n2406_n4888# 0.052164f
C102 plus.n30 a_n2406_n4888# 0.052164f
C103 plus.n31 a_n2406_n4888# 0.018108f
C104 plus.n32 a_n2406_n4888# 0.171771f
C105 plus.n33 a_n2406_n4888# 0.022129f
C106 plus.n34 a_n2406_n4888# 0.171771f
C107 plus.t22 a_n2406_n4888# 0.443096f
C108 plus.n35 a_n2406_n4888# 0.190756f
C109 plus.n36 a_n2406_n4888# 0.794861f
C110 plus.n37 a_n2406_n4888# 0.052164f
C111 plus.t6 a_n2406_n4888# 0.443096f
C112 plus.t2 a_n2406_n4888# 0.440757f
C113 plus.t0 a_n2406_n4888# 0.440757f
C114 plus.n38 a_n2406_n4888# 0.021325f
C115 plus.n39 a_n2406_n4888# 0.052164f
C116 plus.t8 a_n2406_n4888# 0.440757f
C117 plus.n40 a_n2406_n4888# 0.171771f
C118 plus.t5 a_n2406_n4888# 0.440757f
C119 plus.t4 a_n2406_n4888# 0.440757f
C120 plus.n41 a_n2406_n4888# 0.019717f
C121 plus.n42 a_n2406_n4888# 0.052164f
C122 plus.t1 a_n2406_n4888# 0.440757f
C123 plus.n43 a_n2406_n4888# 0.171771f
C124 plus.t13 a_n2406_n4888# 0.440757f
C125 plus.t7 a_n2406_n4888# 0.440757f
C126 plus.n44 a_n2406_n4888# 0.018108f
C127 plus.t9 a_n2406_n4888# 0.443096f
C128 plus.n45 a_n2406_n4888# 0.190829f
C129 plus.t3 a_n2406_n4888# 0.440757f
C130 plus.n46 a_n2406_n4888# 0.171771f
C131 plus.t18 a_n2406_n4888# 0.440757f
C132 plus.n47 a_n2406_n4888# 0.171771f
C133 plus.n48 a_n2406_n4888# 0.022129f
C134 plus.n49 a_n2406_n4888# 0.113904f
C135 plus.n50 a_n2406_n4888# 0.052164f
C136 plus.n51 a_n2406_n4888# 0.052164f
C137 plus.n52 a_n2406_n4888# 0.021325f
C138 plus.n53 a_n2406_n4888# 0.171771f
C139 plus.n54 a_n2406_n4888# 0.022129f
C140 plus.n55 a_n2406_n4888# 0.171771f
C141 plus.n56 a_n2406_n4888# 0.022129f
C142 plus.n57 a_n2406_n4888# 0.052164f
C143 plus.n58 a_n2406_n4888# 0.052164f
C144 plus.n59 a_n2406_n4888# 0.052164f
C145 plus.n60 a_n2406_n4888# 0.019717f
C146 plus.n61 a_n2406_n4888# 0.171771f
C147 plus.n62 a_n2406_n4888# 0.022129f
C148 plus.n63 a_n2406_n4888# 0.171771f
C149 plus.n64 a_n2406_n4888# 0.022129f
C150 plus.n65 a_n2406_n4888# 0.052164f
C151 plus.n66 a_n2406_n4888# 0.052164f
C152 plus.n67 a_n2406_n4888# 0.052164f
C153 plus.n68 a_n2406_n4888# 0.018108f
C154 plus.n69 a_n2406_n4888# 0.171771f
C155 plus.n70 a_n2406_n4888# 0.022129f
C156 plus.n71 a_n2406_n4888# 0.171771f
C157 plus.n72 a_n2406_n4888# 0.190756f
C158 plus.n73 a_n2406_n4888# 1.9937f
C159 source.t7 a_n2406_n4888# 4.852859f
C160 source.n0 a_n2406_n4888# 1.97028f
C161 source.t12 a_n2406_n4888# 0.596712f
C162 source.t13 a_n2406_n4888# 0.596712f
C163 source.n1 a_n2406_n4888# 3.92677f
C164 source.n2 a_n2406_n4888# 0.345865f
C165 source.t2 a_n2406_n4888# 0.596712f
C166 source.t4 a_n2406_n4888# 0.596712f
C167 source.n3 a_n2406_n4888# 3.92677f
C168 source.n4 a_n2406_n4888# 0.345865f
C169 source.t9 a_n2406_n4888# 0.596712f
C170 source.t17 a_n2406_n4888# 0.596712f
C171 source.n5 a_n2406_n4888# 3.92677f
C172 source.n6 a_n2406_n4888# 0.345865f
C173 source.t20 a_n2406_n4888# 0.596712f
C174 source.t14 a_n2406_n4888# 0.596712f
C175 source.n7 a_n2406_n4888# 3.92677f
C176 source.n8 a_n2406_n4888# 0.345865f
C177 source.t3 a_n2406_n4888# 0.596712f
C178 source.t21 a_n2406_n4888# 0.596712f
C179 source.n9 a_n2406_n4888# 3.92677f
C180 source.n10 a_n2406_n4888# 0.345865f
C181 source.t10 a_n2406_n4888# 4.85287f
C182 source.n11 a_n2406_n4888# 0.486579f
C183 source.t40 a_n2406_n4888# 4.85287f
C184 source.n12 a_n2406_n4888# 0.486579f
C185 source.t34 a_n2406_n4888# 0.596712f
C186 source.t42 a_n2406_n4888# 0.596712f
C187 source.n13 a_n2406_n4888# 3.92677f
C188 source.n14 a_n2406_n4888# 0.345865f
C189 source.t39 a_n2406_n4888# 0.596712f
C190 source.t37 a_n2406_n4888# 0.596712f
C191 source.n15 a_n2406_n4888# 3.92677f
C192 source.n16 a_n2406_n4888# 0.345865f
C193 source.t33 a_n2406_n4888# 0.596712f
C194 source.t29 a_n2406_n4888# 0.596712f
C195 source.n17 a_n2406_n4888# 3.92677f
C196 source.n18 a_n2406_n4888# 0.345865f
C197 source.t36 a_n2406_n4888# 0.596712f
C198 source.t32 a_n2406_n4888# 0.596712f
C199 source.n19 a_n2406_n4888# 3.92677f
C200 source.n20 a_n2406_n4888# 0.345865f
C201 source.t28 a_n2406_n4888# 0.596712f
C202 source.t25 a_n2406_n4888# 0.596712f
C203 source.n21 a_n2406_n4888# 3.92677f
C204 source.n22 a_n2406_n4888# 0.345865f
C205 source.t31 a_n2406_n4888# 4.85287f
C206 source.n23 a_n2406_n4888# 2.41245f
C207 source.t5 a_n2406_n4888# 4.85285f
C208 source.n24 a_n2406_n4888# 2.41248f
C209 source.t19 a_n2406_n4888# 0.596712f
C210 source.t0 a_n2406_n4888# 0.596712f
C211 source.n25 a_n2406_n4888# 3.92678f
C212 source.n26 a_n2406_n4888# 0.345858f
C213 source.t11 a_n2406_n4888# 0.596712f
C214 source.t1 a_n2406_n4888# 0.596712f
C215 source.n27 a_n2406_n4888# 3.92678f
C216 source.n28 a_n2406_n4888# 0.345858f
C217 source.t16 a_n2406_n4888# 0.596712f
C218 source.t15 a_n2406_n4888# 0.596712f
C219 source.n29 a_n2406_n4888# 3.92678f
C220 source.n30 a_n2406_n4888# 0.345858f
C221 source.t18 a_n2406_n4888# 0.596712f
C222 source.t6 a_n2406_n4888# 0.596712f
C223 source.n31 a_n2406_n4888# 3.92678f
C224 source.n32 a_n2406_n4888# 0.345858f
C225 source.t23 a_n2406_n4888# 0.596712f
C226 source.t22 a_n2406_n4888# 0.596712f
C227 source.n33 a_n2406_n4888# 3.92678f
C228 source.n34 a_n2406_n4888# 0.345858f
C229 source.t8 a_n2406_n4888# 4.85285f
C230 source.n35 a_n2406_n4888# 0.486603f
C231 source.t43 a_n2406_n4888# 4.85285f
C232 source.n36 a_n2406_n4888# 0.486603f
C233 source.t30 a_n2406_n4888# 0.596712f
C234 source.t24 a_n2406_n4888# 0.596712f
C235 source.n37 a_n2406_n4888# 3.92678f
C236 source.n38 a_n2406_n4888# 0.345858f
C237 source.t45 a_n2406_n4888# 0.596712f
C238 source.t38 a_n2406_n4888# 0.596712f
C239 source.n39 a_n2406_n4888# 3.92678f
C240 source.n40 a_n2406_n4888# 0.345858f
C241 source.t27 a_n2406_n4888# 0.596712f
C242 source.t47 a_n2406_n4888# 0.596712f
C243 source.n41 a_n2406_n4888# 3.92678f
C244 source.n42 a_n2406_n4888# 0.345858f
C245 source.t44 a_n2406_n4888# 0.596712f
C246 source.t35 a_n2406_n4888# 0.596712f
C247 source.n43 a_n2406_n4888# 3.92678f
C248 source.n44 a_n2406_n4888# 0.345858f
C249 source.t26 a_n2406_n4888# 0.596712f
C250 source.t46 a_n2406_n4888# 0.596712f
C251 source.n45 a_n2406_n4888# 3.92678f
C252 source.n46 a_n2406_n4888# 0.345858f
C253 source.t41 a_n2406_n4888# 4.85285f
C254 source.n47 a_n2406_n4888# 0.628375f
C255 source.n48 a_n2406_n4888# 2.24401f
C256 drain_right.t7 a_n2406_n4888# 0.675185f
C257 drain_right.t14 a_n2406_n4888# 0.675185f
C258 drain_right.n0 a_n2406_n4888# 4.53636f
C259 drain_right.t2 a_n2406_n4888# 0.675185f
C260 drain_right.t1 a_n2406_n4888# 0.675185f
C261 drain_right.n1 a_n2406_n4888# 4.5331f
C262 drain_right.n2 a_n2406_n4888# 0.687597f
C263 drain_right.t22 a_n2406_n4888# 0.675185f
C264 drain_right.t11 a_n2406_n4888# 0.675185f
C265 drain_right.n3 a_n2406_n4888# 4.5331f
C266 drain_right.n4 a_n2406_n4888# 0.312174f
C267 drain_right.t4 a_n2406_n4888# 0.675185f
C268 drain_right.t9 a_n2406_n4888# 0.675185f
C269 drain_right.n5 a_n2406_n4888# 4.53636f
C270 drain_right.t13 a_n2406_n4888# 0.675185f
C271 drain_right.t10 a_n2406_n4888# 0.675185f
C272 drain_right.n6 a_n2406_n4888# 4.5331f
C273 drain_right.n7 a_n2406_n4888# 0.687597f
C274 drain_right.t5 a_n2406_n4888# 0.675185f
C275 drain_right.t0 a_n2406_n4888# 0.675185f
C276 drain_right.n8 a_n2406_n4888# 4.5331f
C277 drain_right.n9 a_n2406_n4888# 0.312174f
C278 drain_right.n10 a_n2406_n4888# 2.04212f
C279 drain_right.t6 a_n2406_n4888# 0.675185f
C280 drain_right.t8 a_n2406_n4888# 0.675185f
C281 drain_right.n11 a_n2406_n4888# 4.53636f
C282 drain_right.t21 a_n2406_n4888# 0.675185f
C283 drain_right.t12 a_n2406_n4888# 0.675185f
C284 drain_right.n12 a_n2406_n4888# 4.5331f
C285 drain_right.n13 a_n2406_n4888# 0.687609f
C286 drain_right.t19 a_n2406_n4888# 0.675185f
C287 drain_right.t23 a_n2406_n4888# 0.675185f
C288 drain_right.n14 a_n2406_n4888# 4.5331f
C289 drain_right.n15 a_n2406_n4888# 0.339755f
C290 drain_right.t16 a_n2406_n4888# 0.675185f
C291 drain_right.t17 a_n2406_n4888# 0.675185f
C292 drain_right.n16 a_n2406_n4888# 4.5331f
C293 drain_right.n17 a_n2406_n4888# 0.339755f
C294 drain_right.t3 a_n2406_n4888# 0.675185f
C295 drain_right.t20 a_n2406_n4888# 0.675185f
C296 drain_right.n18 a_n2406_n4888# 4.5331f
C297 drain_right.n19 a_n2406_n4888# 0.339755f
C298 drain_right.t15 a_n2406_n4888# 0.675185f
C299 drain_right.t18 a_n2406_n4888# 0.675185f
C300 drain_right.n20 a_n2406_n4888# 4.5331f
C301 drain_right.n21 a_n2406_n4888# 0.575219f
C302 minus.n0 a_n2406_n4888# 0.051456f
C303 minus.t16 a_n2406_n4888# 0.437081f
C304 minus.t19 a_n2406_n4888# 0.434774f
C305 minus.t22 a_n2406_n4888# 0.434774f
C306 minus.n1 a_n2406_n4888# 0.021035f
C307 minus.n2 a_n2406_n4888# 0.051456f
C308 minus.t11 a_n2406_n4888# 0.434774f
C309 minus.n3 a_n2406_n4888# 0.169439f
C310 minus.t15 a_n2406_n4888# 0.434774f
C311 minus.t14 a_n2406_n4888# 0.434774f
C312 minus.n4 a_n2406_n4888# 0.019449f
C313 minus.n5 a_n2406_n4888# 0.051456f
C314 minus.t18 a_n2406_n4888# 0.434774f
C315 minus.n6 a_n2406_n4888# 0.169439f
C316 minus.t8 a_n2406_n4888# 0.434774f
C317 minus.t10 a_n2406_n4888# 0.434774f
C318 minus.n7 a_n2406_n4888# 0.017863f
C319 minus.t7 a_n2406_n4888# 0.437081f
C320 minus.n8 a_n2406_n4888# 0.188239f
C321 minus.t13 a_n2406_n4888# 0.434774f
C322 minus.n9 a_n2406_n4888# 0.169439f
C323 minus.t5 a_n2406_n4888# 0.434774f
C324 minus.n10 a_n2406_n4888# 0.169439f
C325 minus.n11 a_n2406_n4888# 0.021828f
C326 minus.n12 a_n2406_n4888# 0.112358f
C327 minus.n13 a_n2406_n4888# 0.051456f
C328 minus.n14 a_n2406_n4888# 0.051456f
C329 minus.n15 a_n2406_n4888# 0.021035f
C330 minus.n16 a_n2406_n4888# 0.169439f
C331 minus.n17 a_n2406_n4888# 0.021828f
C332 minus.n18 a_n2406_n4888# 0.169439f
C333 minus.n19 a_n2406_n4888# 0.021828f
C334 minus.n20 a_n2406_n4888# 0.051456f
C335 minus.n21 a_n2406_n4888# 0.051456f
C336 minus.n22 a_n2406_n4888# 0.051456f
C337 minus.n23 a_n2406_n4888# 0.019449f
C338 minus.n24 a_n2406_n4888# 0.169439f
C339 minus.n25 a_n2406_n4888# 0.021828f
C340 minus.n26 a_n2406_n4888# 0.169439f
C341 minus.n27 a_n2406_n4888# 0.021828f
C342 minus.n28 a_n2406_n4888# 0.051456f
C343 minus.n29 a_n2406_n4888# 0.051456f
C344 minus.n30 a_n2406_n4888# 0.051456f
C345 minus.n31 a_n2406_n4888# 0.017863f
C346 minus.n32 a_n2406_n4888# 0.169439f
C347 minus.n33 a_n2406_n4888# 0.021828f
C348 minus.n34 a_n2406_n4888# 0.169439f
C349 minus.n35 a_n2406_n4888# 0.188167f
C350 minus.n36 a_n2406_n4888# 2.46527f
C351 minus.n37 a_n2406_n4888# 0.051456f
C352 minus.t1 a_n2406_n4888# 0.434774f
C353 minus.t21 a_n2406_n4888# 0.434774f
C354 minus.n38 a_n2406_n4888# 0.021035f
C355 minus.n39 a_n2406_n4888# 0.051456f
C356 minus.t3 a_n2406_n4888# 0.434774f
C357 minus.t0 a_n2406_n4888# 0.434774f
C358 minus.n40 a_n2406_n4888# 0.019449f
C359 minus.n41 a_n2406_n4888# 0.051456f
C360 minus.t9 a_n2406_n4888# 0.434774f
C361 minus.t2 a_n2406_n4888# 0.434774f
C362 minus.n42 a_n2406_n4888# 0.017863f
C363 minus.t4 a_n2406_n4888# 0.437081f
C364 minus.n43 a_n2406_n4888# 0.188239f
C365 minus.t17 a_n2406_n4888# 0.434774f
C366 minus.n44 a_n2406_n4888# 0.169439f
C367 minus.t23 a_n2406_n4888# 0.434774f
C368 minus.n45 a_n2406_n4888# 0.169439f
C369 minus.n46 a_n2406_n4888# 0.021828f
C370 minus.n47 a_n2406_n4888# 0.112358f
C371 minus.n48 a_n2406_n4888# 0.051456f
C372 minus.n49 a_n2406_n4888# 0.051456f
C373 minus.n50 a_n2406_n4888# 0.021035f
C374 minus.n51 a_n2406_n4888# 0.169439f
C375 minus.n52 a_n2406_n4888# 0.021828f
C376 minus.n53 a_n2406_n4888# 0.169439f
C377 minus.t20 a_n2406_n4888# 0.434774f
C378 minus.n54 a_n2406_n4888# 0.169439f
C379 minus.n55 a_n2406_n4888# 0.021828f
C380 minus.n56 a_n2406_n4888# 0.051456f
C381 minus.n57 a_n2406_n4888# 0.051456f
C382 minus.n58 a_n2406_n4888# 0.051456f
C383 minus.n59 a_n2406_n4888# 0.019449f
C384 minus.n60 a_n2406_n4888# 0.169439f
C385 minus.n61 a_n2406_n4888# 0.021828f
C386 minus.n62 a_n2406_n4888# 0.169439f
C387 minus.t12 a_n2406_n4888# 0.434774f
C388 minus.n63 a_n2406_n4888# 0.169439f
C389 minus.n64 a_n2406_n4888# 0.021828f
C390 minus.n65 a_n2406_n4888# 0.051456f
C391 minus.n66 a_n2406_n4888# 0.051456f
C392 minus.n67 a_n2406_n4888# 0.051456f
C393 minus.n68 a_n2406_n4888# 0.017863f
C394 minus.n69 a_n2406_n4888# 0.169439f
C395 minus.n70 a_n2406_n4888# 0.021828f
C396 minus.n71 a_n2406_n4888# 0.169439f
C397 minus.t6 a_n2406_n4888# 0.437081f
C398 minus.n72 a_n2406_n4888# 0.188167f
C399 minus.n73 a_n2406_n4888# 0.339218f
C400 minus.n74 a_n2406_n4888# 2.92426f
.ends

