* NGSPICE file created from diffpair344.ext - technology: sky130A

.subckt diffpair344 minus drain_right drain_left source plus
X0 source.t19 plus.t0 drain_left.t6 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 source.t18 plus.t1 drain_left.t4 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 source.t6 minus.t0 drain_right.t9 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_left.t3 plus.t2 source.t17 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X4 source.t4 minus.t1 drain_right.t8 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 drain_right.t7 minus.t2 source.t9 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X6 source.t1 minus.t3 drain_right.t6 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 drain_left.t8 plus.t3 source.t16 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 drain_left.t0 plus.t4 source.t15 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X9 drain_left.t1 plus.t5 source.t14 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X10 drain_left.t9 plus.t6 source.t13 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X11 source.t5 minus.t4 drain_right.t5 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X12 a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X13 source.t12 plus.t7 drain_left.t2 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X14 a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X15 drain_right.t4 minus.t5 source.t8 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X16 drain_right.t3 minus.t6 source.t7 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 drain_right.t2 minus.t7 source.t0 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X18 drain_left.t5 plus.t8 source.t11 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X19 drain_right.t1 minus.t8 source.t3 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X20 source.t10 plus.t9 drain_left.t7 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X21 drain_right.t0 minus.t9 source.t2 a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X22 a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X23 a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# a_n1412_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
R0 plus.n2 plus.t4 1052.8
R1 plus.n8 plus.t5 1052.8
R2 plus.n12 plus.t8 1052.8
R3 plus.n18 plus.t2 1052.8
R4 plus.n1 plus.t1 992.92
R5 plus.n5 plus.t6 992.92
R6 plus.n7 plus.t0 992.92
R7 plus.n11 plus.t7 992.92
R8 plus.n15 plus.t3 992.92
R9 plus.n17 plus.t9 992.92
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 27.2301
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 11.0232
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n5 drain_left.t0 68.2376
R37 drain_left.n1 drain_left.t3 68.2373
R38 drain_left.n3 drain_left.n2 65.857
R39 drain_left.n5 drain_left.n4 65.5376
R40 drain_left.n7 drain_left.n6 65.5374
R41 drain_left.n1 drain_left.n0 65.5373
R42 drain_left drain_left.n3 27.2193
R43 drain_left drain_left.n7 6.15322
R44 drain_left.n2 drain_left.t2 2.2005
R45 drain_left.n2 drain_left.t5 2.2005
R46 drain_left.n0 drain_left.t7 2.2005
R47 drain_left.n0 drain_left.t8 2.2005
R48 drain_left.n6 drain_left.t6 2.2005
R49 drain_left.n6 drain_left.t1 2.2005
R50 drain_left.n4 drain_left.t4 2.2005
R51 drain_left.n4 drain_left.t9 2.2005
R52 drain_left.n7 drain_left.n5 0.5005
R53 drain_left.n3 drain_left.n1 0.070154
R54 source.n5 source.t0 51.0588
R55 source.n19 source.t9 51.0586
R56 source.n14 source.t11 51.0586
R57 source.n0 source.t14 51.0586
R58 source.n2 source.n1 48.8588
R59 source.n4 source.n3 48.8588
R60 source.n7 source.n6 48.8588
R61 source.n9 source.n8 48.8588
R62 source.n18 source.n17 48.8586
R63 source.n16 source.n15 48.8586
R64 source.n13 source.n12 48.8586
R65 source.n11 source.n10 48.8586
R66 source.n11 source.n9 20.015
R67 source.n20 source.n0 14.0021
R68 source.n20 source.n19 5.51343
R69 source.n17 source.t7 2.2005
R70 source.n17 source.t5 2.2005
R71 source.n15 source.t3 2.2005
R72 source.n15 source.t6 2.2005
R73 source.n12 source.t16 2.2005
R74 source.n12 source.t12 2.2005
R75 source.n10 source.t17 2.2005
R76 source.n10 source.t10 2.2005
R77 source.n1 source.t13 2.2005
R78 source.n1 source.t19 2.2005
R79 source.n3 source.t15 2.2005
R80 source.n3 source.t18 2.2005
R81 source.n6 source.t8 2.2005
R82 source.n6 source.t1 2.2005
R83 source.n8 source.t2 2.2005
R84 source.n8 source.t4 2.2005
R85 source.n5 source.n4 0.720328
R86 source.n16 source.n14 0.720328
R87 source.n9 source.n7 0.5005
R88 source.n7 source.n5 0.5005
R89 source.n4 source.n2 0.5005
R90 source.n2 source.n0 0.5005
R91 source.n13 source.n11 0.5005
R92 source.n14 source.n13 0.5005
R93 source.n18 source.n16 0.5005
R94 source.n19 source.n18 0.5005
R95 source source.n20 0.188
R96 minus.n8 minus.t9 1052.8
R97 minus.n2 minus.t7 1052.8
R98 minus.n18 minus.t2 1052.8
R99 minus.n12 minus.t8 1052.8
R100 minus.n7 minus.t1 992.92
R101 minus.n5 minus.t5 992.92
R102 minus.n1 minus.t3 992.92
R103 minus.n17 minus.t4 992.92
R104 minus.n15 minus.t6 992.92
R105 minus.n11 minus.t0 992.92
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 48.2005
R115 minus.n4 minus.n1 48.2005
R116 minus.n14 minus.n11 48.2005
R117 minus.n17 minus.n16 48.2005
R118 minus.n6 minus.n5 36.5157
R119 minus.n5 minus.n4 36.5157
R120 minus.n15 minus.n14 36.5157
R121 minus.n16 minus.n15 36.5157
R122 minus.n20 minus.n9 32.2126
R123 minus.n8 minus.n7 24.8308
R124 minus.n2 minus.n1 24.8308
R125 minus.n12 minus.n11 24.8308
R126 minus.n18 minus.n17 24.8308
R127 minus.n20 minus.n19 6.51565
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t1 68.2373
R134 drain_right.n7 drain_right.t0 67.7376
R135 drain_right.n6 drain_right.n4 66.0374
R136 drain_right.n3 drain_right.n2 65.857
R137 drain_right.n6 drain_right.n5 65.5376
R138 drain_right.n1 drain_right.n0 65.5373
R139 drain_right drain_right.n3 26.6661
R140 drain_right drain_right.n7 5.90322
R141 drain_right.n2 drain_right.t5 2.2005
R142 drain_right.n2 drain_right.t7 2.2005
R143 drain_right.n0 drain_right.t9 2.2005
R144 drain_right.n0 drain_right.t3 2.2005
R145 drain_right.n4 drain_right.t6 2.2005
R146 drain_right.n4 drain_right.t2 2.2005
R147 drain_right.n5 drain_right.t8 2.2005
R148 drain_right.n5 drain_right.t4 2.2005
R149 drain_right.n7 drain_right.n6 0.5005
R150 drain_right.n3 drain_right.n1 0.070154
C0 drain_right source 17.5927f
C1 drain_left plus 2.88861f
C2 drain_right plus 0.289643f
C3 drain_left drain_right 0.692689f
C4 minus source 2.45666f
C5 plus minus 4.354509f
C6 plus source 2.4712f
C7 drain_left minus 0.171039f
C8 drain_right minus 2.75662f
C9 drain_left source 17.6019f
C10 drain_right a_n1412_n2688# 6.03485f
C11 drain_left a_n1412_n2688# 6.26864f
C12 source a_n1412_n2688# 4.996522f
C13 minus a_n1412_n2688# 5.238443f
C14 plus a_n1412_n2688# 7.07142f
C15 drain_right.t1 a_n1412_n2688# 2.4641f
C16 drain_right.t9 a_n1412_n2688# 0.221063f
C17 drain_right.t3 a_n1412_n2688# 0.221063f
C18 drain_right.n0 a_n1412_n2688# 1.93357f
C19 drain_right.n1 a_n1412_n2688# 0.700318f
C20 drain_right.t5 a_n1412_n2688# 0.221063f
C21 drain_right.t7 a_n1412_n2688# 0.221063f
C22 drain_right.n2 a_n1412_n2688# 1.93525f
C23 drain_right.n3 a_n1412_n2688# 1.44363f
C24 drain_right.t6 a_n1412_n2688# 0.221063f
C25 drain_right.t2 a_n1412_n2688# 0.221063f
C26 drain_right.n4 a_n1412_n2688# 1.9363f
C27 drain_right.t8 a_n1412_n2688# 0.221063f
C28 drain_right.t4 a_n1412_n2688# 0.221063f
C29 drain_right.n5 a_n1412_n2688# 1.93357f
C30 drain_right.n6 a_n1412_n2688# 0.708047f
C31 drain_right.t0 a_n1412_n2688# 2.46127f
C32 drain_right.n7 a_n1412_n2688# 0.642747f
C33 minus.n0 a_n1412_n2688# 0.055877f
C34 minus.t9 a_n1412_n2688# 0.36519f
C35 minus.t1 a_n1412_n2688# 0.356251f
C36 minus.t5 a_n1412_n2688# 0.356251f
C37 minus.t3 a_n1412_n2688# 0.356251f
C38 minus.n1 a_n1412_n2688# 0.151635f
C39 minus.t7 a_n1412_n2688# 0.36519f
C40 minus.n2 a_n1412_n2688# 0.16959f
C41 minus.n3 a_n1412_n2688# 0.131303f
C42 minus.n4 a_n1412_n2688# 0.021292f
C43 minus.n5 a_n1412_n2688# 0.151635f
C44 minus.n6 a_n1412_n2688# 0.021292f
C45 minus.n7 a_n1412_n2688# 0.151635f
C46 minus.n8 a_n1412_n2688# 0.169501f
C47 minus.n9 a_n1412_n2688# 1.63867f
C48 minus.n10 a_n1412_n2688# 0.055877f
C49 minus.t4 a_n1412_n2688# 0.356251f
C50 minus.t6 a_n1412_n2688# 0.356251f
C51 minus.t0 a_n1412_n2688# 0.356251f
C52 minus.n11 a_n1412_n2688# 0.151635f
C53 minus.t8 a_n1412_n2688# 0.36519f
C54 minus.n12 a_n1412_n2688# 0.16959f
C55 minus.n13 a_n1412_n2688# 0.131303f
C56 minus.n14 a_n1412_n2688# 0.021292f
C57 minus.n15 a_n1412_n2688# 0.151635f
C58 minus.n16 a_n1412_n2688# 0.021292f
C59 minus.n17 a_n1412_n2688# 0.151635f
C60 minus.t2 a_n1412_n2688# 0.36519f
C61 minus.n18 a_n1412_n2688# 0.169501f
C62 minus.n19 a_n1412_n2688# 0.36737f
C63 minus.n20 a_n1412_n2688# 2.01147f
C64 source.t14 a_n1412_n2688# 2.47124f
C65 source.n0 a_n1412_n2688# 1.41345f
C66 source.t13 a_n1412_n2688# 0.231748f
C67 source.t19 a_n1412_n2688# 0.231748f
C68 source.n1 a_n1412_n2688# 1.94005f
C69 source.n2 a_n1412_n2688# 0.408697f
C70 source.t15 a_n1412_n2688# 0.231748f
C71 source.t18 a_n1412_n2688# 0.231748f
C72 source.n3 a_n1412_n2688# 1.94005f
C73 source.n4 a_n1412_n2688# 0.431778f
C74 source.t0 a_n1412_n2688# 2.47125f
C75 source.n5 a_n1412_n2688# 0.532618f
C76 source.t8 a_n1412_n2688# 0.231748f
C77 source.t1 a_n1412_n2688# 0.231748f
C78 source.n6 a_n1412_n2688# 1.94005f
C79 source.n7 a_n1412_n2688# 0.408697f
C80 source.t2 a_n1412_n2688# 0.231748f
C81 source.t4 a_n1412_n2688# 0.231748f
C82 source.n8 a_n1412_n2688# 1.94005f
C83 source.n9 a_n1412_n2688# 1.83709f
C84 source.t17 a_n1412_n2688# 0.231748f
C85 source.t10 a_n1412_n2688# 0.231748f
C86 source.n10 a_n1412_n2688# 1.94004f
C87 source.n11 a_n1412_n2688# 1.8371f
C88 source.t16 a_n1412_n2688# 0.231748f
C89 source.t12 a_n1412_n2688# 0.231748f
C90 source.n12 a_n1412_n2688# 1.94004f
C91 source.n13 a_n1412_n2688# 0.408702f
C92 source.t11 a_n1412_n2688# 2.47124f
C93 source.n14 a_n1412_n2688# 0.532624f
C94 source.t3 a_n1412_n2688# 0.231748f
C95 source.t6 a_n1412_n2688# 0.231748f
C96 source.n15 a_n1412_n2688# 1.94004f
C97 source.n16 a_n1412_n2688# 0.431784f
C98 source.t7 a_n1412_n2688# 0.231748f
C99 source.t5 a_n1412_n2688# 0.231748f
C100 source.n17 a_n1412_n2688# 1.94004f
C101 source.n18 a_n1412_n2688# 0.408702f
C102 source.t9 a_n1412_n2688# 2.47124f
C103 source.n19 a_n1412_n2688# 0.686696f
C104 source.n20 a_n1412_n2688# 1.69391f
C105 drain_left.t3 a_n1412_n2688# 2.46151f
C106 drain_left.t7 a_n1412_n2688# 0.220831f
C107 drain_left.t8 a_n1412_n2688# 0.220831f
C108 drain_left.n0 a_n1412_n2688# 1.93153f
C109 drain_left.n1 a_n1412_n2688# 0.699581f
C110 drain_left.t2 a_n1412_n2688# 0.220831f
C111 drain_left.t5 a_n1412_n2688# 0.220831f
C112 drain_left.n2 a_n1412_n2688# 1.93321f
C113 drain_left.n3 a_n1412_n2688# 1.50654f
C114 drain_left.t0 a_n1412_n2688# 2.46151f
C115 drain_left.t4 a_n1412_n2688# 0.220831f
C116 drain_left.t9 a_n1412_n2688# 0.220831f
C117 drain_left.n4 a_n1412_n2688# 1.93154f
C118 drain_left.n5 a_n1412_n2688# 0.732295f
C119 drain_left.t6 a_n1412_n2688# 0.220831f
C120 drain_left.t1 a_n1412_n2688# 0.220831f
C121 drain_left.n6 a_n1412_n2688# 1.93153f
C122 drain_left.n7 a_n1412_n2688# 0.605068f
C123 plus.n0 a_n1412_n2688# 0.057119f
C124 plus.t0 a_n1412_n2688# 0.364166f
C125 plus.t6 a_n1412_n2688# 0.364166f
C126 plus.t1 a_n1412_n2688# 0.364166f
C127 plus.n1 a_n1412_n2688# 0.155004f
C128 plus.t4 a_n1412_n2688# 0.373304f
C129 plus.n2 a_n1412_n2688# 0.173357f
C130 plus.n3 a_n1412_n2688# 0.13422f
C131 plus.n4 a_n1412_n2688# 0.021765f
C132 plus.n5 a_n1412_n2688# 0.155004f
C133 plus.n6 a_n1412_n2688# 0.021765f
C134 plus.n7 a_n1412_n2688# 0.155004f
C135 plus.t5 a_n1412_n2688# 0.373304f
C136 plus.n8 a_n1412_n2688# 0.173267f
C137 plus.n9 a_n1412_n2688# 0.563243f
C138 plus.n10 a_n1412_n2688# 0.057119f
C139 plus.t2 a_n1412_n2688# 0.373304f
C140 plus.t9 a_n1412_n2688# 0.364166f
C141 plus.t3 a_n1412_n2688# 0.364166f
C142 plus.t7 a_n1412_n2688# 0.364166f
C143 plus.n11 a_n1412_n2688# 0.155004f
C144 plus.t8 a_n1412_n2688# 0.373304f
C145 plus.n12 a_n1412_n2688# 0.173357f
C146 plus.n13 a_n1412_n2688# 0.13422f
C147 plus.n14 a_n1412_n2688# 0.021765f
C148 plus.n15 a_n1412_n2688# 0.155004f
C149 plus.n16 a_n1412_n2688# 0.021765f
C150 plus.n17 a_n1412_n2688# 0.155004f
C151 plus.n18 a_n1412_n2688# 0.173267f
C152 plus.n19 a_n1412_n2688# 1.45908f
.ends

