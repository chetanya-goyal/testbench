* NGSPICE file created from diffpair41.ext - technology: sky130A

.subckt diffpair41 minus drain_right drain_left source plus
X0 source minus drain_right a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X1 source plus drain_left a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 source minus drain_right a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_left plus source a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X5 drain_right minus source a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X6 drain_right minus source a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X7 drain_left plus source a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X8 source plus drain_left a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X9 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X10 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X11 a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# a_n1214_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
.ends

