* NGSPICE file created from diffpair617.ext - technology: sky130A

.subckt diffpair617 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t23 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X1 drain_left.t15 plus.t0 source.t3 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X2 source.t9 plus.t1 drain_left.t14 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X3 source.t14 plus.t2 drain_left.t13 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X4 drain_left.t12 plus.t3 source.t2 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X5 source.t13 plus.t4 drain_left.t11 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X6 drain_left.t10 plus.t5 source.t4 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X7 source.t18 minus.t1 drain_right.t14 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X8 drain_right.t13 minus.t2 source.t17 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X9 drain_right.t12 minus.t3 source.t16 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X10 drain_right.t11 minus.t4 source.t26 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X11 drain_left.t9 plus.t6 source.t15 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X12 source.t21 minus.t5 drain_right.t10 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X13 source.t30 minus.t6 drain_right.t9 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X14 drain_right.t8 minus.t7 source.t29 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X15 source.t1 plus.t7 drain_left.t8 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X16 a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.6
X17 source.t7 plus.t8 drain_left.t7 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X18 a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X19 source.t28 minus.t8 drain_right.t7 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X20 source.t20 minus.t9 drain_right.t6 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X21 drain_right.t5 minus.t10 source.t31 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X22 source.t11 plus.t9 drain_left.t6 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X23 a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X24 drain_left.t5 plus.t10 source.t5 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X25 source.t24 minus.t11 drain_right.t4 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X26 source.t6 plus.t11 drain_left.t4 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X27 drain_right.t3 minus.t12 source.t25 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
X28 source.t19 minus.t13 drain_right.t2 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X29 drain_left.t3 plus.t12 source.t10 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X30 source.t0 plus.t13 drain_left.t2 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X31 a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.6
X32 source.t27 minus.t14 drain_right.t1 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.6
X33 drain_left.t1 plus.t14 source.t8 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X34 drain_left.t0 plus.t15 source.t12 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.6
X35 drain_right.t0 minus.t15 source.t22 a_n2390_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.6
R0 minus.n6 minus.t12 889.788
R1 minus.n30 minus.t14 889.788
R2 minus.n5 minus.t11 868.806
R3 minus.n9 minus.t10 868.806
R4 minus.n3 minus.t8 868.806
R5 minus.n15 minus.t3 868.806
R6 minus.n1 minus.t5 868.806
R7 minus.n21 minus.t4 868.806
R8 minus.n22 minus.t1 868.806
R9 minus.n29 minus.t7 868.806
R10 minus.n33 minus.t9 868.806
R11 minus.n27 minus.t0 868.806
R12 minus.n39 minus.t6 868.806
R13 minus.n25 minus.t2 868.806
R14 minus.n45 minus.t13 868.806
R15 minus.n46 minus.t15 868.806
R16 minus.n23 minus.n22 161.3
R17 minus.n21 minus.n0 161.3
R18 minus.n20 minus.n19 161.3
R19 minus.n18 minus.n1 161.3
R20 minus.n17 minus.n16 161.3
R21 minus.n15 minus.n2 161.3
R22 minus.n14 minus.n13 161.3
R23 minus.n12 minus.n3 161.3
R24 minus.n11 minus.n10 161.3
R25 minus.n9 minus.n4 161.3
R26 minus.n8 minus.n7 161.3
R27 minus.n47 minus.n46 161.3
R28 minus.n45 minus.n24 161.3
R29 minus.n44 minus.n43 161.3
R30 minus.n42 minus.n25 161.3
R31 minus.n41 minus.n40 161.3
R32 minus.n39 minus.n26 161.3
R33 minus.n38 minus.n37 161.3
R34 minus.n36 minus.n27 161.3
R35 minus.n35 minus.n34 161.3
R36 minus.n33 minus.n28 161.3
R37 minus.n32 minus.n31 161.3
R38 minus.n7 minus.n6 70.4033
R39 minus.n31 minus.n30 70.4033
R40 minus.n22 minus.n21 48.2005
R41 minus.n46 minus.n45 48.2005
R42 minus.n9 minus.n8 44.549
R43 minus.n20 minus.n1 44.549
R44 minus.n33 minus.n32 44.549
R45 minus.n44 minus.n25 44.549
R46 minus.n48 minus.n23 44.3906
R47 minus.n10 minus.n3 34.3247
R48 minus.n16 minus.n15 34.3247
R49 minus.n34 minus.n27 34.3247
R50 minus.n40 minus.n39 34.3247
R51 minus.n15 minus.n14 24.1005
R52 minus.n14 minus.n3 24.1005
R53 minus.n38 minus.n27 24.1005
R54 minus.n39 minus.n38 24.1005
R55 minus.n6 minus.n5 20.9576
R56 minus.n30 minus.n29 20.9576
R57 minus.n10 minus.n9 13.8763
R58 minus.n16 minus.n1 13.8763
R59 minus.n34 minus.n33 13.8763
R60 minus.n40 minus.n25 13.8763
R61 minus.n48 minus.n47 6.6558
R62 minus.n8 minus.n5 3.65202
R63 minus.n21 minus.n20 3.65202
R64 minus.n32 minus.n29 3.65202
R65 minus.n45 minus.n44 3.65202
R66 minus.n23 minus.n0 0.189894
R67 minus.n19 minus.n0 0.189894
R68 minus.n19 minus.n18 0.189894
R69 minus.n18 minus.n17 0.189894
R70 minus.n17 minus.n2 0.189894
R71 minus.n13 minus.n2 0.189894
R72 minus.n13 minus.n12 0.189894
R73 minus.n12 minus.n11 0.189894
R74 minus.n11 minus.n4 0.189894
R75 minus.n7 minus.n4 0.189894
R76 minus.n31 minus.n28 0.189894
R77 minus.n35 minus.n28 0.189894
R78 minus.n36 minus.n35 0.189894
R79 minus.n37 minus.n36 0.189894
R80 minus.n37 minus.n26 0.189894
R81 minus.n41 minus.n26 0.189894
R82 minus.n42 minus.n41 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n24 0.189894
R85 minus.n47 minus.n24 0.189894
R86 minus minus.n48 0.188
R87 source.n0 source.t2 44.1297
R88 source.n7 source.t0 44.1296
R89 source.n8 source.t25 44.1296
R90 source.n15 source.t18 44.1296
R91 source.n31 source.t22 44.1295
R92 source.n24 source.t27 44.1295
R93 source.n23 source.t3 44.1295
R94 source.n16 source.t14 44.1295
R95 source.n2 source.n1 43.1397
R96 source.n4 source.n3 43.1397
R97 source.n6 source.n5 43.1397
R98 source.n10 source.n9 43.1397
R99 source.n12 source.n11 43.1397
R100 source.n14 source.n13 43.1397
R101 source.n30 source.n29 43.1396
R102 source.n28 source.n27 43.1396
R103 source.n26 source.n25 43.1396
R104 source.n22 source.n21 43.1396
R105 source.n20 source.n19 43.1396
R106 source.n18 source.n17 43.1396
R107 source.n16 source.n15 28.1501
R108 source.n32 source.n0 22.4863
R109 source.n32 source.n31 5.66429
R110 source.n29 source.t17 0.9905
R111 source.n29 source.t19 0.9905
R112 source.n27 source.t23 0.9905
R113 source.n27 source.t30 0.9905
R114 source.n25 source.t29 0.9905
R115 source.n25 source.t20 0.9905
R116 source.n21 source.t8 0.9905
R117 source.n21 source.t11 0.9905
R118 source.n19 source.t15 0.9905
R119 source.n19 source.t9 0.9905
R120 source.n17 source.t12 0.9905
R121 source.n17 source.t1 0.9905
R122 source.n1 source.t4 0.9905
R123 source.n1 source.t13 0.9905
R124 source.n3 source.t5 0.9905
R125 source.n3 source.t7 0.9905
R126 source.n5 source.t10 0.9905
R127 source.n5 source.t6 0.9905
R128 source.n9 source.t31 0.9905
R129 source.n9 source.t24 0.9905
R130 source.n11 source.t16 0.9905
R131 source.n11 source.t28 0.9905
R132 source.n13 source.t26 0.9905
R133 source.n13 source.t21 0.9905
R134 source.n15 source.n14 0.802224
R135 source.n14 source.n12 0.802224
R136 source.n12 source.n10 0.802224
R137 source.n10 source.n8 0.802224
R138 source.n7 source.n6 0.802224
R139 source.n6 source.n4 0.802224
R140 source.n4 source.n2 0.802224
R141 source.n2 source.n0 0.802224
R142 source.n18 source.n16 0.802224
R143 source.n20 source.n18 0.802224
R144 source.n22 source.n20 0.802224
R145 source.n23 source.n22 0.802224
R146 source.n26 source.n24 0.802224
R147 source.n28 source.n26 0.802224
R148 source.n30 source.n28 0.802224
R149 source.n31 source.n30 0.802224
R150 source.n8 source.n7 0.470328
R151 source.n24 source.n23 0.470328
R152 source source.n32 0.188
R153 drain_right.n9 drain_right.n7 60.6202
R154 drain_right.n5 drain_right.n3 60.6201
R155 drain_right.n2 drain_right.n0 60.6201
R156 drain_right.n9 drain_right.n8 59.8185
R157 drain_right.n11 drain_right.n10 59.8185
R158 drain_right.n13 drain_right.n12 59.8185
R159 drain_right.n5 drain_right.n4 59.8184
R160 drain_right.n2 drain_right.n1 59.8184
R161 drain_right drain_right.n6 38.0857
R162 drain_right drain_right.n13 6.45494
R163 drain_right.n3 drain_right.t2 0.9905
R164 drain_right.n3 drain_right.t0 0.9905
R165 drain_right.n4 drain_right.t9 0.9905
R166 drain_right.n4 drain_right.t13 0.9905
R167 drain_right.n1 drain_right.t6 0.9905
R168 drain_right.n1 drain_right.t15 0.9905
R169 drain_right.n0 drain_right.t1 0.9905
R170 drain_right.n0 drain_right.t8 0.9905
R171 drain_right.n7 drain_right.t4 0.9905
R172 drain_right.n7 drain_right.t3 0.9905
R173 drain_right.n8 drain_right.t7 0.9905
R174 drain_right.n8 drain_right.t5 0.9905
R175 drain_right.n10 drain_right.t10 0.9905
R176 drain_right.n10 drain_right.t12 0.9905
R177 drain_right.n12 drain_right.t14 0.9905
R178 drain_right.n12 drain_right.t11 0.9905
R179 drain_right.n13 drain_right.n11 0.802224
R180 drain_right.n11 drain_right.n9 0.802224
R181 drain_right.n6 drain_right.n5 0.346016
R182 drain_right.n6 drain_right.n2 0.346016
R183 plus.n6 plus.t13 889.788
R184 plus.n30 plus.t0 889.788
R185 plus.n22 plus.t3 868.806
R186 plus.n21 plus.t4 868.806
R187 plus.n1 plus.t5 868.806
R188 plus.n15 plus.t8 868.806
R189 plus.n3 plus.t10 868.806
R190 plus.n9 plus.t11 868.806
R191 plus.n5 plus.t12 868.806
R192 plus.n46 plus.t2 868.806
R193 plus.n45 plus.t15 868.806
R194 plus.n25 plus.t7 868.806
R195 plus.n39 plus.t6 868.806
R196 plus.n27 plus.t1 868.806
R197 plus.n33 plus.t14 868.806
R198 plus.n29 plus.t9 868.806
R199 plus.n8 plus.n7 161.3
R200 plus.n9 plus.n4 161.3
R201 plus.n11 plus.n10 161.3
R202 plus.n12 plus.n3 161.3
R203 plus.n14 plus.n13 161.3
R204 plus.n15 plus.n2 161.3
R205 plus.n17 plus.n16 161.3
R206 plus.n18 plus.n1 161.3
R207 plus.n20 plus.n19 161.3
R208 plus.n21 plus.n0 161.3
R209 plus.n23 plus.n22 161.3
R210 plus.n32 plus.n31 161.3
R211 plus.n33 plus.n28 161.3
R212 plus.n35 plus.n34 161.3
R213 plus.n36 plus.n27 161.3
R214 plus.n38 plus.n37 161.3
R215 plus.n39 plus.n26 161.3
R216 plus.n41 plus.n40 161.3
R217 plus.n42 plus.n25 161.3
R218 plus.n44 plus.n43 161.3
R219 plus.n45 plus.n24 161.3
R220 plus.n47 plus.n46 161.3
R221 plus.n7 plus.n6 70.4033
R222 plus.n31 plus.n30 70.4033
R223 plus.n22 plus.n21 48.2005
R224 plus.n46 plus.n45 48.2005
R225 plus.n20 plus.n1 44.549
R226 plus.n9 plus.n8 44.549
R227 plus.n44 plus.n25 44.549
R228 plus.n33 plus.n32 44.549
R229 plus plus.n47 35.2414
R230 plus.n16 plus.n15 34.3247
R231 plus.n10 plus.n3 34.3247
R232 plus.n40 plus.n39 34.3247
R233 plus.n34 plus.n27 34.3247
R234 plus.n14 plus.n3 24.1005
R235 plus.n15 plus.n14 24.1005
R236 plus.n39 plus.n38 24.1005
R237 plus.n38 plus.n27 24.1005
R238 plus.n6 plus.n5 20.9576
R239 plus.n30 plus.n29 20.9576
R240 plus plus.n23 15.33
R241 plus.n16 plus.n1 13.8763
R242 plus.n10 plus.n9 13.8763
R243 plus.n40 plus.n25 13.8763
R244 plus.n34 plus.n33 13.8763
R245 plus.n21 plus.n20 3.65202
R246 plus.n8 plus.n5 3.65202
R247 plus.n45 plus.n44 3.65202
R248 plus.n32 plus.n29 3.65202
R249 plus.n7 plus.n4 0.189894
R250 plus.n11 plus.n4 0.189894
R251 plus.n12 plus.n11 0.189894
R252 plus.n13 plus.n12 0.189894
R253 plus.n13 plus.n2 0.189894
R254 plus.n17 plus.n2 0.189894
R255 plus.n18 plus.n17 0.189894
R256 plus.n19 plus.n18 0.189894
R257 plus.n19 plus.n0 0.189894
R258 plus.n23 plus.n0 0.189894
R259 plus.n47 plus.n24 0.189894
R260 plus.n43 plus.n24 0.189894
R261 plus.n43 plus.n42 0.189894
R262 plus.n42 plus.n41 0.189894
R263 plus.n41 plus.n26 0.189894
R264 plus.n37 plus.n26 0.189894
R265 plus.n37 plus.n36 0.189894
R266 plus.n36 plus.n35 0.189894
R267 plus.n35 plus.n28 0.189894
R268 plus.n31 plus.n28 0.189894
R269 drain_left.n9 drain_left.n7 60.6202
R270 drain_left.n5 drain_left.n3 60.6201
R271 drain_left.n2 drain_left.n0 60.6201
R272 drain_left.n13 drain_left.n12 59.8185
R273 drain_left.n11 drain_left.n10 59.8185
R274 drain_left.n9 drain_left.n8 59.8185
R275 drain_left.n5 drain_left.n4 59.8184
R276 drain_left.n2 drain_left.n1 59.8184
R277 drain_left drain_left.n6 38.6389
R278 drain_left drain_left.n13 6.45494
R279 drain_left.n3 drain_left.t6 0.9905
R280 drain_left.n3 drain_left.t15 0.9905
R281 drain_left.n4 drain_left.t14 0.9905
R282 drain_left.n4 drain_left.t1 0.9905
R283 drain_left.n1 drain_left.t8 0.9905
R284 drain_left.n1 drain_left.t9 0.9905
R285 drain_left.n0 drain_left.t13 0.9905
R286 drain_left.n0 drain_left.t0 0.9905
R287 drain_left.n12 drain_left.t11 0.9905
R288 drain_left.n12 drain_left.t12 0.9905
R289 drain_left.n10 drain_left.t7 0.9905
R290 drain_left.n10 drain_left.t10 0.9905
R291 drain_left.n8 drain_left.t4 0.9905
R292 drain_left.n8 drain_left.t5 0.9905
R293 drain_left.n7 drain_left.t2 0.9905
R294 drain_left.n7 drain_left.t3 0.9905
R295 drain_left.n11 drain_left.n9 0.802224
R296 drain_left.n13 drain_left.n11 0.802224
R297 drain_left.n6 drain_left.n5 0.346016
R298 drain_left.n6 drain_left.n2 0.346016
C0 source drain_left 33.486202f
C1 plus source 14.886299f
C2 source minus 14.872299f
C3 plus drain_left 15.4592f
C4 drain_left minus 0.172752f
C5 plus minus 7.605721f
C6 source drain_right 33.4879f
C7 drain_left drain_right 1.24373f
C8 plus drain_right 0.391974f
C9 minus drain_right 15.2233f
C10 drain_right a_n2390_n4888# 8.16399f
C11 drain_left a_n2390_n4888# 8.51099f
C12 source a_n2390_n4888# 13.610124f
C13 minus a_n2390_n4888# 10.022881f
C14 plus a_n2390_n4888# 12.25932f
C15 drain_left.t13 a_n2390_n4888# 0.446316f
C16 drain_left.t0 a_n2390_n4888# 0.446316f
C17 drain_left.n0 a_n2390_n4888# 4.08555f
C18 drain_left.t8 a_n2390_n4888# 0.446316f
C19 drain_left.t9 a_n2390_n4888# 0.446316f
C20 drain_left.n1 a_n2390_n4888# 4.08032f
C21 drain_left.n2 a_n2390_n4888# 0.734939f
C22 drain_left.t6 a_n2390_n4888# 0.446316f
C23 drain_left.t15 a_n2390_n4888# 0.446316f
C24 drain_left.n3 a_n2390_n4888# 4.08555f
C25 drain_left.t14 a_n2390_n4888# 0.446316f
C26 drain_left.t1 a_n2390_n4888# 0.446316f
C27 drain_left.n4 a_n2390_n4888# 4.08032f
C28 drain_left.n5 a_n2390_n4888# 0.734939f
C29 drain_left.n6 a_n2390_n4888# 2.11743f
C30 drain_left.t2 a_n2390_n4888# 0.446316f
C31 drain_left.t3 a_n2390_n4888# 0.446316f
C32 drain_left.n7 a_n2390_n4888# 4.08555f
C33 drain_left.t4 a_n2390_n4888# 0.446316f
C34 drain_left.t5 a_n2390_n4888# 0.446316f
C35 drain_left.n8 a_n2390_n4888# 4.08032f
C36 drain_left.n9 a_n2390_n4888# 0.774568f
C37 drain_left.t7 a_n2390_n4888# 0.446316f
C38 drain_left.t10 a_n2390_n4888# 0.446316f
C39 drain_left.n10 a_n2390_n4888# 4.08032f
C40 drain_left.n11 a_n2390_n4888# 0.384213f
C41 drain_left.t11 a_n2390_n4888# 0.446316f
C42 drain_left.t12 a_n2390_n4888# 0.446316f
C43 drain_left.n12 a_n2390_n4888# 4.08032f
C44 drain_left.n13 a_n2390_n4888# 0.63046f
C45 plus.n0 a_n2390_n4888# 0.042923f
C46 plus.t3 a_n2390_n4888# 1.45863f
C47 plus.t4 a_n2390_n4888# 1.45863f
C48 plus.t5 a_n2390_n4888# 1.45863f
C49 plus.n1 a_n2390_n4888# 0.547844f
C50 plus.n2 a_n2390_n4888# 0.042923f
C51 plus.t8 a_n2390_n4888# 1.45863f
C52 plus.t10 a_n2390_n4888# 1.45863f
C53 plus.n3 a_n2390_n4888# 0.547844f
C54 plus.n4 a_n2390_n4888# 0.042923f
C55 plus.t11 a_n2390_n4888# 1.45863f
C56 plus.t12 a_n2390_n4888# 1.45863f
C57 plus.n5 a_n2390_n4888# 0.546653f
C58 plus.t13 a_n2390_n4888# 1.47151f
C59 plus.n6 a_n2390_n4888# 0.533459f
C60 plus.n7 a_n2390_n4888# 0.144568f
C61 plus.n8 a_n2390_n4888# 0.00974f
C62 plus.n9 a_n2390_n4888# 0.547844f
C63 plus.n10 a_n2390_n4888# 0.00974f
C64 plus.n11 a_n2390_n4888# 0.042923f
C65 plus.n12 a_n2390_n4888# 0.042923f
C66 plus.n13 a_n2390_n4888# 0.042923f
C67 plus.n14 a_n2390_n4888# 0.00974f
C68 plus.n15 a_n2390_n4888# 0.547844f
C69 plus.n16 a_n2390_n4888# 0.00974f
C70 plus.n17 a_n2390_n4888# 0.042923f
C71 plus.n18 a_n2390_n4888# 0.042923f
C72 plus.n19 a_n2390_n4888# 0.042923f
C73 plus.n20 a_n2390_n4888# 0.00974f
C74 plus.n21 a_n2390_n4888# 0.546653f
C75 plus.n22 a_n2390_n4888# 0.545992f
C76 plus.n23 a_n2390_n4888# 0.667091f
C77 plus.n24 a_n2390_n4888# 0.042923f
C78 plus.t2 a_n2390_n4888# 1.45863f
C79 plus.t15 a_n2390_n4888# 1.45863f
C80 plus.t7 a_n2390_n4888# 1.45863f
C81 plus.n25 a_n2390_n4888# 0.547844f
C82 plus.n26 a_n2390_n4888# 0.042923f
C83 plus.t6 a_n2390_n4888# 1.45863f
C84 plus.t1 a_n2390_n4888# 1.45863f
C85 plus.n27 a_n2390_n4888# 0.547844f
C86 plus.n28 a_n2390_n4888# 0.042923f
C87 plus.t14 a_n2390_n4888# 1.45863f
C88 plus.t9 a_n2390_n4888# 1.45863f
C89 plus.n29 a_n2390_n4888# 0.546653f
C90 plus.t0 a_n2390_n4888# 1.47151f
C91 plus.n30 a_n2390_n4888# 0.533459f
C92 plus.n31 a_n2390_n4888# 0.144568f
C93 plus.n32 a_n2390_n4888# 0.00974f
C94 plus.n33 a_n2390_n4888# 0.547844f
C95 plus.n34 a_n2390_n4888# 0.00974f
C96 plus.n35 a_n2390_n4888# 0.042923f
C97 plus.n36 a_n2390_n4888# 0.042923f
C98 plus.n37 a_n2390_n4888# 0.042923f
C99 plus.n38 a_n2390_n4888# 0.00974f
C100 plus.n39 a_n2390_n4888# 0.547844f
C101 plus.n40 a_n2390_n4888# 0.00974f
C102 plus.n41 a_n2390_n4888# 0.042923f
C103 plus.n42 a_n2390_n4888# 0.042923f
C104 plus.n43 a_n2390_n4888# 0.042923f
C105 plus.n44 a_n2390_n4888# 0.00974f
C106 plus.n45 a_n2390_n4888# 0.546653f
C107 plus.n46 a_n2390_n4888# 0.545992f
C108 plus.n47 a_n2390_n4888# 1.64932f
C109 drain_right.t1 a_n2390_n4888# 0.444586f
C110 drain_right.t8 a_n2390_n4888# 0.444586f
C111 drain_right.n0 a_n2390_n4888# 4.06971f
C112 drain_right.t6 a_n2390_n4888# 0.444586f
C113 drain_right.t15 a_n2390_n4888# 0.444586f
C114 drain_right.n1 a_n2390_n4888# 4.0645f
C115 drain_right.n2 a_n2390_n4888# 0.73209f
C116 drain_right.t2 a_n2390_n4888# 0.444586f
C117 drain_right.t0 a_n2390_n4888# 0.444586f
C118 drain_right.n3 a_n2390_n4888# 4.06971f
C119 drain_right.t9 a_n2390_n4888# 0.444586f
C120 drain_right.t13 a_n2390_n4888# 0.444586f
C121 drain_right.n4 a_n2390_n4888# 4.0645f
C122 drain_right.n5 a_n2390_n4888# 0.732089f
C123 drain_right.n6 a_n2390_n4888# 2.05112f
C124 drain_right.t4 a_n2390_n4888# 0.444586f
C125 drain_right.t3 a_n2390_n4888# 0.444586f
C126 drain_right.n7 a_n2390_n4888# 4.06971f
C127 drain_right.t7 a_n2390_n4888# 0.444586f
C128 drain_right.t5 a_n2390_n4888# 0.444586f
C129 drain_right.n8 a_n2390_n4888# 4.0645f
C130 drain_right.n9 a_n2390_n4888# 0.771565f
C131 drain_right.t10 a_n2390_n4888# 0.444586f
C132 drain_right.t12 a_n2390_n4888# 0.444586f
C133 drain_right.n10 a_n2390_n4888# 4.0645f
C134 drain_right.n11 a_n2390_n4888# 0.382723f
C135 drain_right.t14 a_n2390_n4888# 0.444586f
C136 drain_right.t11 a_n2390_n4888# 0.444586f
C137 drain_right.n12 a_n2390_n4888# 4.0645f
C138 drain_right.n13 a_n2390_n4888# 0.628016f
C139 source.t2 a_n2390_n4888# 4.19793f
C140 source.n0 a_n2390_n4888# 1.81604f
C141 source.t4 a_n2390_n4888# 0.367325f
C142 source.t13 a_n2390_n4888# 0.367325f
C143 source.n1 a_n2390_n4888# 3.28404f
C144 source.n2 a_n2390_n4888# 0.358741f
C145 source.t5 a_n2390_n4888# 0.367325f
C146 source.t7 a_n2390_n4888# 0.367325f
C147 source.n3 a_n2390_n4888# 3.28404f
C148 source.n4 a_n2390_n4888# 0.358741f
C149 source.t10 a_n2390_n4888# 0.367325f
C150 source.t6 a_n2390_n4888# 0.367325f
C151 source.n5 a_n2390_n4888# 3.28404f
C152 source.n6 a_n2390_n4888# 0.358741f
C153 source.t0 a_n2390_n4888# 4.19794f
C154 source.n7 a_n2390_n4888# 0.421785f
C155 source.t25 a_n2390_n4888# 4.19794f
C156 source.n8 a_n2390_n4888# 0.421785f
C157 source.t31 a_n2390_n4888# 0.367325f
C158 source.t24 a_n2390_n4888# 0.367325f
C159 source.n9 a_n2390_n4888# 3.28404f
C160 source.n10 a_n2390_n4888# 0.358741f
C161 source.t16 a_n2390_n4888# 0.367325f
C162 source.t28 a_n2390_n4888# 0.367325f
C163 source.n11 a_n2390_n4888# 3.28404f
C164 source.n12 a_n2390_n4888# 0.358741f
C165 source.t26 a_n2390_n4888# 0.367325f
C166 source.t21 a_n2390_n4888# 0.367325f
C167 source.n13 a_n2390_n4888# 3.28404f
C168 source.n14 a_n2390_n4888# 0.358741f
C169 source.t18 a_n2390_n4888# 4.19794f
C170 source.n15 a_n2390_n4888# 2.23613f
C171 source.t14 a_n2390_n4888# 4.19792f
C172 source.n16 a_n2390_n4888# 2.23615f
C173 source.t12 a_n2390_n4888# 0.367325f
C174 source.t1 a_n2390_n4888# 0.367325f
C175 source.n17 a_n2390_n4888# 3.28405f
C176 source.n18 a_n2390_n4888# 0.358735f
C177 source.t15 a_n2390_n4888# 0.367325f
C178 source.t9 a_n2390_n4888# 0.367325f
C179 source.n19 a_n2390_n4888# 3.28405f
C180 source.n20 a_n2390_n4888# 0.358735f
C181 source.t8 a_n2390_n4888# 0.367325f
C182 source.t11 a_n2390_n4888# 0.367325f
C183 source.n21 a_n2390_n4888# 3.28405f
C184 source.n22 a_n2390_n4888# 0.358735f
C185 source.t3 a_n2390_n4888# 4.19792f
C186 source.n23 a_n2390_n4888# 0.421808f
C187 source.t27 a_n2390_n4888# 4.19792f
C188 source.n24 a_n2390_n4888# 0.421808f
C189 source.t29 a_n2390_n4888# 0.367325f
C190 source.t20 a_n2390_n4888# 0.367325f
C191 source.n25 a_n2390_n4888# 3.28405f
C192 source.n26 a_n2390_n4888# 0.358735f
C193 source.t23 a_n2390_n4888# 0.367325f
C194 source.t30 a_n2390_n4888# 0.367325f
C195 source.n27 a_n2390_n4888# 3.28405f
C196 source.n28 a_n2390_n4888# 0.358735f
C197 source.t17 a_n2390_n4888# 0.367325f
C198 source.t19 a_n2390_n4888# 0.367325f
C199 source.n29 a_n2390_n4888# 3.28405f
C200 source.n30 a_n2390_n4888# 0.358735f
C201 source.t22 a_n2390_n4888# 4.19792f
C202 source.n31 a_n2390_n4888# 0.568355f
C203 source.n32 a_n2390_n4888# 2.10441f
C204 minus.n0 a_n2390_n4888# 0.042487f
C205 minus.t5 a_n2390_n4888# 1.44382f
C206 minus.n1 a_n2390_n4888# 0.542281f
C207 minus.n2 a_n2390_n4888# 0.042487f
C208 minus.t8 a_n2390_n4888# 1.44382f
C209 minus.n3 a_n2390_n4888# 0.542281f
C210 minus.n4 a_n2390_n4888# 0.042487f
C211 minus.t11 a_n2390_n4888# 1.44382f
C212 minus.n5 a_n2390_n4888# 0.541102f
C213 minus.t12 a_n2390_n4888# 1.45657f
C214 minus.n6 a_n2390_n4888# 0.528041f
C215 minus.n7 a_n2390_n4888# 0.1431f
C216 minus.n8 a_n2390_n4888# 0.009641f
C217 minus.t10 a_n2390_n4888# 1.44382f
C218 minus.n9 a_n2390_n4888# 0.542281f
C219 minus.n10 a_n2390_n4888# 0.009641f
C220 minus.n11 a_n2390_n4888# 0.042487f
C221 minus.n12 a_n2390_n4888# 0.042487f
C222 minus.n13 a_n2390_n4888# 0.042487f
C223 minus.n14 a_n2390_n4888# 0.009641f
C224 minus.t3 a_n2390_n4888# 1.44382f
C225 minus.n15 a_n2390_n4888# 0.542281f
C226 minus.n16 a_n2390_n4888# 0.009641f
C227 minus.n17 a_n2390_n4888# 0.042487f
C228 minus.n18 a_n2390_n4888# 0.042487f
C229 minus.n19 a_n2390_n4888# 0.042487f
C230 minus.n20 a_n2390_n4888# 0.009641f
C231 minus.t4 a_n2390_n4888# 1.44382f
C232 minus.n21 a_n2390_n4888# 0.541102f
C233 minus.t1 a_n2390_n4888# 1.44382f
C234 minus.n22 a_n2390_n4888# 0.540447f
C235 minus.n23 a_n2390_n4888# 2.04387f
C236 minus.n24 a_n2390_n4888# 0.042487f
C237 minus.t2 a_n2390_n4888# 1.44382f
C238 minus.n25 a_n2390_n4888# 0.542281f
C239 minus.n26 a_n2390_n4888# 0.042487f
C240 minus.t0 a_n2390_n4888# 1.44382f
C241 minus.n27 a_n2390_n4888# 0.542281f
C242 minus.n28 a_n2390_n4888# 0.042487f
C243 minus.t7 a_n2390_n4888# 1.44382f
C244 minus.n29 a_n2390_n4888# 0.541102f
C245 minus.t14 a_n2390_n4888# 1.45657f
C246 minus.n30 a_n2390_n4888# 0.528041f
C247 minus.n31 a_n2390_n4888# 0.1431f
C248 minus.n32 a_n2390_n4888# 0.009641f
C249 minus.t9 a_n2390_n4888# 1.44382f
C250 minus.n33 a_n2390_n4888# 0.542281f
C251 minus.n34 a_n2390_n4888# 0.009641f
C252 minus.n35 a_n2390_n4888# 0.042487f
C253 minus.n36 a_n2390_n4888# 0.042487f
C254 minus.n37 a_n2390_n4888# 0.042487f
C255 minus.n38 a_n2390_n4888# 0.009641f
C256 minus.t6 a_n2390_n4888# 1.44382f
C257 minus.n39 a_n2390_n4888# 0.542281f
C258 minus.n40 a_n2390_n4888# 0.009641f
C259 minus.n41 a_n2390_n4888# 0.042487f
C260 minus.n42 a_n2390_n4888# 0.042487f
C261 minus.n43 a_n2390_n4888# 0.042487f
C262 minus.n44 a_n2390_n4888# 0.009641f
C263 minus.t13 a_n2390_n4888# 1.44382f
C264 minus.n45 a_n2390_n4888# 0.541102f
C265 minus.t15 a_n2390_n4888# 1.44382f
C266 minus.n46 a_n2390_n4888# 0.540447f
C267 minus.n47 a_n2390_n4888# 0.29325f
C268 minus.n48 a_n2390_n4888# 2.42136f
.ends

