* NGSPICE file created from diffpair497.ext - technology: sky130A

.subckt diffpair497 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t25 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t14 plus.t1 source.t19 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X2 a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X3 drain_left.t13 plus.t2 source.t29 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X4 drain_right.t15 minus.t0 source.t8 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 drain_right.t14 minus.t1 source.t7 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 source.t22 plus.t3 drain_left.t12 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X7 a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X8 source.t16 plus.t4 drain_left.t11 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 drain_left.t10 plus.t5 source.t17 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X10 source.t30 minus.t2 drain_right.t13 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X11 source.t31 minus.t3 drain_right.t12 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X12 source.t2 minus.t4 drain_right.t11 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X13 source.t6 minus.t5 drain_right.t10 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X14 drain_left.t9 plus.t6 source.t20 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X15 source.t18 plus.t7 drain_left.t8 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X16 drain_right.t9 minus.t6 source.t1 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X17 drain_right.t8 minus.t7 source.t10 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X18 a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X19 drain_right.t7 minus.t8 source.t12 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X20 a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X21 drain_right.t6 minus.t9 source.t5 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X22 drain_right.t5 minus.t10 source.t9 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X23 drain_right.t4 minus.t11 source.t11 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X24 source.t4 minus.t12 drain_right.t3 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X25 source.t13 minus.t13 drain_right.t2 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X26 source.t28 plus.t8 drain_left.t7 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X27 drain_left.t6 plus.t9 source.t26 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X28 source.t3 minus.t14 drain_right.t1 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X29 source.t0 minus.t15 drain_right.t0 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X30 source.t14 plus.t10 drain_left.t5 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X31 source.t23 plus.t11 drain_left.t4 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X32 source.t27 plus.t12 drain_left.t3 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X33 drain_left.t2 plus.t13 source.t24 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X34 source.t21 plus.t14 drain_left.t1 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X35 drain_left.t0 plus.t15 source.t15 a_n1670_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n4 plus.t7 2016
R1 plus.n17 plus.t13 2016
R2 plus.n23 plus.t2 2016
R3 plus.n36 plus.t10 2016
R4 plus.n3 plus.t5 1964.15
R5 plus.n7 plus.t14 1964.15
R6 plus.n9 plus.t9 1964.15
R7 plus.n1 plus.t8 1964.15
R8 plus.n14 plus.t6 1964.15
R9 plus.n16 plus.t4 1964.15
R10 plus.n22 plus.t3 1964.15
R11 plus.n26 plus.t1 1964.15
R12 plus.n28 plus.t11 1964.15
R13 plus.n20 plus.t0 1964.15
R14 plus.n33 plus.t12 1964.15
R15 plus.n35 plus.t15 1964.15
R16 plus.n5 plus.n4 161.489
R17 plus.n24 plus.n23 161.489
R18 plus.n6 plus.n5 161.3
R19 plus.n8 plus.n2 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n0 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n25 plus.n24 161.3
R25 plus.n27 plus.n21 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n19 161.3
R29 plus.n37 plus.n36 161.3
R30 plus.n6 plus.n3 47.4702
R31 plus.n16 plus.n15 47.4702
R32 plus.n35 plus.n34 47.4702
R33 plus.n25 plus.n22 47.4702
R34 plus.n8 plus.n7 43.0884
R35 plus.n14 plus.n13 43.0884
R36 plus.n33 plus.n32 43.0884
R37 plus.n27 plus.n26 43.0884
R38 plus.n10 plus.n9 38.7066
R39 plus.n10 plus.n1 38.7066
R40 plus.n29 plus.n20 38.7066
R41 plus.n29 plus.n28 38.7066
R42 plus.n9 plus.n8 34.3247
R43 plus.n13 plus.n1 34.3247
R44 plus.n32 plus.n20 34.3247
R45 plus.n28 plus.n27 34.3247
R46 plus plus.n37 30.4308
R47 plus.n7 plus.n6 29.9429
R48 plus.n15 plus.n14 29.9429
R49 plus.n34 plus.n33 29.9429
R50 plus.n26 plus.n25 29.9429
R51 plus.n4 plus.n3 25.5611
R52 plus.n17 plus.n16 25.5611
R53 plus.n36 plus.n35 25.5611
R54 plus.n23 plus.n22 25.5611
R55 plus plus.n18 13.2467
R56 plus.n5 plus.n2 0.189894
R57 plus.n11 plus.n2 0.189894
R58 plus.n12 plus.n11 0.189894
R59 plus.n12 plus.n0 0.189894
R60 plus.n18 plus.n0 0.189894
R61 plus.n37 plus.n19 0.189894
R62 plus.n31 plus.n19 0.189894
R63 plus.n31 plus.n30 0.189894
R64 plus.n30 plus.n21 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n7 source.t18 45.521
R67 source.n8 source.t9 45.521
R68 source.n15 source.t0 45.521
R69 source.n31 source.t12 45.5208
R70 source.n24 source.t6 45.5208
R71 source.n23 source.t29 45.5208
R72 source.n16 source.t14 45.5208
R73 source.n0 source.t24 45.5208
R74 source.n2 source.n1 44.201
R75 source.n4 source.n3 44.201
R76 source.n6 source.n5 44.201
R77 source.n10 source.n9 44.201
R78 source.n12 source.n11 44.201
R79 source.n14 source.n13 44.201
R80 source.n30 source.n29 44.2008
R81 source.n28 source.n27 44.2008
R82 source.n26 source.n25 44.2008
R83 source.n22 source.n21 44.2008
R84 source.n20 source.n19 44.2008
R85 source.n18 source.n17 44.2008
R86 source.n16 source.n15 24.0173
R87 source.n32 source.n0 18.526
R88 source.n32 source.n31 5.49188
R89 source.n29 source.t5 1.3205
R90 source.n29 source.t4 1.3205
R91 source.n27 source.t1 1.3205
R92 source.n27 source.t13 1.3205
R93 source.n25 source.t10 1.3205
R94 source.n25 source.t31 1.3205
R95 source.n21 source.t19 1.3205
R96 source.n21 source.t22 1.3205
R97 source.n19 source.t25 1.3205
R98 source.n19 source.t23 1.3205
R99 source.n17 source.t15 1.3205
R100 source.n17 source.t27 1.3205
R101 source.n1 source.t20 1.3205
R102 source.n1 source.t16 1.3205
R103 source.n3 source.t26 1.3205
R104 source.n3 source.t28 1.3205
R105 source.n5 source.t17 1.3205
R106 source.n5 source.t21 1.3205
R107 source.n9 source.t8 1.3205
R108 source.n9 source.t2 1.3205
R109 source.n11 source.t11 1.3205
R110 source.n11 source.t3 1.3205
R111 source.n13 source.t7 1.3205
R112 source.n13 source.t30 1.3205
R113 source.n8 source.n7 0.470328
R114 source.n24 source.n23 0.470328
R115 source.n15 source.n14 0.457397
R116 source.n14 source.n12 0.457397
R117 source.n12 source.n10 0.457397
R118 source.n10 source.n8 0.457397
R119 source.n7 source.n6 0.457397
R120 source.n6 source.n4 0.457397
R121 source.n4 source.n2 0.457397
R122 source.n2 source.n0 0.457397
R123 source.n18 source.n16 0.457397
R124 source.n20 source.n18 0.457397
R125 source.n22 source.n20 0.457397
R126 source.n23 source.n22 0.457397
R127 source.n26 source.n24 0.457397
R128 source.n28 source.n26 0.457397
R129 source.n30 source.n28 0.457397
R130 source.n31 source.n30 0.457397
R131 source source.n32 0.188
R132 drain_left.n9 drain_left.n7 61.3367
R133 drain_left.n5 drain_left.n3 61.3365
R134 drain_left.n2 drain_left.n0 61.3365
R135 drain_left.n11 drain_left.n10 60.8798
R136 drain_left.n9 drain_left.n8 60.8798
R137 drain_left.n13 drain_left.n12 60.8796
R138 drain_left.n5 drain_left.n4 60.8796
R139 drain_left.n2 drain_left.n1 60.8796
R140 drain_left drain_left.n6 32.6096
R141 drain_left drain_left.n13 6.11011
R142 drain_left.n3 drain_left.t12 1.3205
R143 drain_left.n3 drain_left.t13 1.3205
R144 drain_left.n4 drain_left.t4 1.3205
R145 drain_left.n4 drain_left.t14 1.3205
R146 drain_left.n1 drain_left.t3 1.3205
R147 drain_left.n1 drain_left.t15 1.3205
R148 drain_left.n0 drain_left.t5 1.3205
R149 drain_left.n0 drain_left.t0 1.3205
R150 drain_left.n12 drain_left.t11 1.3205
R151 drain_left.n12 drain_left.t2 1.3205
R152 drain_left.n10 drain_left.t7 1.3205
R153 drain_left.n10 drain_left.t9 1.3205
R154 drain_left.n8 drain_left.t1 1.3205
R155 drain_left.n8 drain_left.t6 1.3205
R156 drain_left.n7 drain_left.t8 1.3205
R157 drain_left.n7 drain_left.t10 1.3205
R158 drain_left.n11 drain_left.n9 0.457397
R159 drain_left.n13 drain_left.n11 0.457397
R160 drain_left.n6 drain_left.n5 0.173602
R161 drain_left.n6 drain_left.n2 0.173602
R162 minus.n17 minus.t15 2016
R163 minus.n4 minus.t10 2016
R164 minus.n36 minus.t8 2016
R165 minus.n23 minus.t5 2016
R166 minus.n16 minus.t1 1964.15
R167 minus.n14 minus.t2 1964.15
R168 minus.n1 minus.t11 1964.15
R169 minus.n9 minus.t14 1964.15
R170 minus.n7 minus.t0 1964.15
R171 minus.n3 minus.t4 1964.15
R172 minus.n35 minus.t12 1964.15
R173 minus.n33 minus.t9 1964.15
R174 minus.n20 minus.t13 1964.15
R175 minus.n28 minus.t6 1964.15
R176 minus.n26 minus.t3 1964.15
R177 minus.n22 minus.t7 1964.15
R178 minus.n5 minus.n4 161.489
R179 minus.n24 minus.n23 161.489
R180 minus.n18 minus.n17 161.3
R181 minus.n15 minus.n0 161.3
R182 minus.n13 minus.n12 161.3
R183 minus.n11 minus.n10 161.3
R184 minus.n8 minus.n2 161.3
R185 minus.n6 minus.n5 161.3
R186 minus.n37 minus.n36 161.3
R187 minus.n34 minus.n19 161.3
R188 minus.n32 minus.n31 161.3
R189 minus.n30 minus.n29 161.3
R190 minus.n27 minus.n21 161.3
R191 minus.n25 minus.n24 161.3
R192 minus.n16 minus.n15 47.4702
R193 minus.n6 minus.n3 47.4702
R194 minus.n25 minus.n22 47.4702
R195 minus.n35 minus.n34 47.4702
R196 minus.n14 minus.n13 43.0884
R197 minus.n8 minus.n7 43.0884
R198 minus.n27 minus.n26 43.0884
R199 minus.n33 minus.n32 43.0884
R200 minus.n10 minus.n1 38.7066
R201 minus.n10 minus.n9 38.7066
R202 minus.n29 minus.n28 38.7066
R203 minus.n29 minus.n20 38.7066
R204 minus.n38 minus.n18 37.6861
R205 minus.n13 minus.n1 34.3247
R206 minus.n9 minus.n8 34.3247
R207 minus.n28 minus.n27 34.3247
R208 minus.n32 minus.n20 34.3247
R209 minus.n15 minus.n14 29.9429
R210 minus.n7 minus.n6 29.9429
R211 minus.n26 minus.n25 29.9429
R212 minus.n34 minus.n33 29.9429
R213 minus.n17 minus.n16 25.5611
R214 minus.n4 minus.n3 25.5611
R215 minus.n23 minus.n22 25.5611
R216 minus.n36 minus.n35 25.5611
R217 minus.n38 minus.n37 6.46641
R218 minus.n18 minus.n0 0.189894
R219 minus.n12 minus.n0 0.189894
R220 minus.n12 minus.n11 0.189894
R221 minus.n11 minus.n2 0.189894
R222 minus.n5 minus.n2 0.189894
R223 minus.n24 minus.n21 0.189894
R224 minus.n30 minus.n21 0.189894
R225 minus.n31 minus.n30 0.189894
R226 minus.n31 minus.n19 0.189894
R227 minus.n37 minus.n19 0.189894
R228 minus minus.n38 0.188
R229 drain_right.n9 drain_right.n7 61.3365
R230 drain_right.n5 drain_right.n3 61.3365
R231 drain_right.n2 drain_right.n0 61.3365
R232 drain_right.n9 drain_right.n8 60.8798
R233 drain_right.n11 drain_right.n10 60.8798
R234 drain_right.n13 drain_right.n12 60.8798
R235 drain_right.n5 drain_right.n4 60.8796
R236 drain_right.n2 drain_right.n1 60.8796
R237 drain_right drain_right.n6 32.0564
R238 drain_right drain_right.n13 6.11011
R239 drain_right.n3 drain_right.t3 1.3205
R240 drain_right.n3 drain_right.t7 1.3205
R241 drain_right.n4 drain_right.t2 1.3205
R242 drain_right.n4 drain_right.t6 1.3205
R243 drain_right.n1 drain_right.t12 1.3205
R244 drain_right.n1 drain_right.t9 1.3205
R245 drain_right.n0 drain_right.t10 1.3205
R246 drain_right.n0 drain_right.t8 1.3205
R247 drain_right.n7 drain_right.t11 1.3205
R248 drain_right.n7 drain_right.t5 1.3205
R249 drain_right.n8 drain_right.t1 1.3205
R250 drain_right.n8 drain_right.t15 1.3205
R251 drain_right.n10 drain_right.t13 1.3205
R252 drain_right.n10 drain_right.t4 1.3205
R253 drain_right.n12 drain_right.t0 1.3205
R254 drain_right.n12 drain_right.t14 1.3205
R255 drain_right.n13 drain_right.n11 0.457397
R256 drain_right.n11 drain_right.n9 0.457397
R257 drain_right.n6 drain_right.n5 0.173602
R258 drain_right.n6 drain_right.n2 0.173602
C0 drain_left drain_right 0.846053f
C1 drain_left source 45.185f
C2 plus drain_right 0.314737f
C3 plus source 4.88171f
C4 minus drain_right 5.40757f
C5 source minus 4.86767f
C6 drain_left plus 5.56853f
C7 drain_left minus 0.170856f
C8 plus minus 5.79278f
C9 source drain_right 45.1847f
C10 drain_right a_n1670_n3888# 7.496319f
C11 drain_left a_n1670_n3888# 7.77098f
C12 source a_n1670_n3888# 10.140311f
C13 minus a_n1670_n3888# 6.674868f
C14 plus a_n1670_n3888# 8.969601f
C15 drain_right.t10 a_n1670_n3888# 0.460554f
C16 drain_right.t8 a_n1670_n3888# 0.460554f
C17 drain_right.n0 a_n1670_n3888# 4.16621f
C18 drain_right.t12 a_n1670_n3888# 0.460554f
C19 drain_right.t9 a_n1670_n3888# 0.460554f
C20 drain_right.n1 a_n1670_n3888# 4.16287f
C21 drain_right.n2 a_n1670_n3888# 0.847267f
C22 drain_right.t3 a_n1670_n3888# 0.460554f
C23 drain_right.t7 a_n1670_n3888# 0.460554f
C24 drain_right.n3 a_n1670_n3888# 4.16621f
C25 drain_right.t2 a_n1670_n3888# 0.460554f
C26 drain_right.t6 a_n1670_n3888# 0.460554f
C27 drain_right.n4 a_n1670_n3888# 4.16287f
C28 drain_right.n5 a_n1670_n3888# 0.847267f
C29 drain_right.n6 a_n1670_n3888# 2.01734f
C30 drain_right.t11 a_n1670_n3888# 0.460554f
C31 drain_right.t5 a_n1670_n3888# 0.460554f
C32 drain_right.n7 a_n1670_n3888# 4.1662f
C33 drain_right.t1 a_n1670_n3888# 0.460554f
C34 drain_right.t15 a_n1670_n3888# 0.460554f
C35 drain_right.n8 a_n1670_n3888# 4.16287f
C36 drain_right.n9 a_n1670_n3888# 0.877601f
C37 drain_right.t13 a_n1670_n3888# 0.460554f
C38 drain_right.t4 a_n1670_n3888# 0.460554f
C39 drain_right.n10 a_n1670_n3888# 4.16287f
C40 drain_right.n11 a_n1670_n3888# 0.432638f
C41 drain_right.t0 a_n1670_n3888# 0.460554f
C42 drain_right.t14 a_n1670_n3888# 0.460554f
C43 drain_right.n12 a_n1670_n3888# 4.16287f
C44 drain_right.n13 a_n1670_n3888# 0.750621f
C45 minus.n0 a_n1670_n3888# 0.05424f
C46 minus.t15 a_n1670_n3888# 0.46378f
C47 minus.t1 a_n1670_n3888# 0.459054f
C48 minus.t2 a_n1670_n3888# 0.459054f
C49 minus.t11 a_n1670_n3888# 0.459054f
C50 minus.n1 a_n1670_n3888# 0.181899f
C51 minus.n2 a_n1670_n3888# 0.05424f
C52 minus.t14 a_n1670_n3888# 0.459054f
C53 minus.t0 a_n1670_n3888# 0.459054f
C54 minus.t4 a_n1670_n3888# 0.459054f
C55 minus.n3 a_n1670_n3888# 0.181899f
C56 minus.t10 a_n1670_n3888# 0.46378f
C57 minus.n4 a_n1670_n3888# 0.198089f
C58 minus.n5 a_n1670_n3888# 0.12211f
C59 minus.n6 a_n1670_n3888# 0.018996f
C60 minus.n7 a_n1670_n3888# 0.181899f
C61 minus.n8 a_n1670_n3888# 0.018996f
C62 minus.n9 a_n1670_n3888# 0.181899f
C63 minus.n10 a_n1670_n3888# 0.018996f
C64 minus.n11 a_n1670_n3888# 0.05424f
C65 minus.n12 a_n1670_n3888# 0.05424f
C66 minus.n13 a_n1670_n3888# 0.018996f
C67 minus.n14 a_n1670_n3888# 0.181899f
C68 minus.n15 a_n1670_n3888# 0.018996f
C69 minus.n16 a_n1670_n3888# 0.181899f
C70 minus.n17 a_n1670_n3888# 0.198009f
C71 minus.n18 a_n1670_n3888# 2.03944f
C72 minus.n19 a_n1670_n3888# 0.05424f
C73 minus.t12 a_n1670_n3888# 0.459054f
C74 minus.t9 a_n1670_n3888# 0.459054f
C75 minus.t13 a_n1670_n3888# 0.459054f
C76 minus.n20 a_n1670_n3888# 0.181899f
C77 minus.n21 a_n1670_n3888# 0.05424f
C78 minus.t6 a_n1670_n3888# 0.459054f
C79 minus.t3 a_n1670_n3888# 0.459054f
C80 minus.t7 a_n1670_n3888# 0.459054f
C81 minus.n22 a_n1670_n3888# 0.181899f
C82 minus.t5 a_n1670_n3888# 0.46378f
C83 minus.n23 a_n1670_n3888# 0.198089f
C84 minus.n24 a_n1670_n3888# 0.12211f
C85 minus.n25 a_n1670_n3888# 0.018996f
C86 minus.n26 a_n1670_n3888# 0.181899f
C87 minus.n27 a_n1670_n3888# 0.018996f
C88 minus.n28 a_n1670_n3888# 0.181899f
C89 minus.n29 a_n1670_n3888# 0.018996f
C90 minus.n30 a_n1670_n3888# 0.05424f
C91 minus.n31 a_n1670_n3888# 0.05424f
C92 minus.n32 a_n1670_n3888# 0.018996f
C93 minus.n33 a_n1670_n3888# 0.181899f
C94 minus.n34 a_n1670_n3888# 0.018996f
C95 minus.n35 a_n1670_n3888# 0.181899f
C96 minus.t8 a_n1670_n3888# 0.46378f
C97 minus.n36 a_n1670_n3888# 0.198009f
C98 minus.n37 a_n1670_n3888# 0.350305f
C99 minus.n38 a_n1670_n3888# 2.46778f
C100 drain_left.t5 a_n1670_n3888# 0.46099f
C101 drain_left.t0 a_n1670_n3888# 0.46099f
C102 drain_left.n0 a_n1670_n3888# 4.17015f
C103 drain_left.t3 a_n1670_n3888# 0.46099f
C104 drain_left.t15 a_n1670_n3888# 0.46099f
C105 drain_left.n1 a_n1670_n3888# 4.16681f
C106 drain_left.n2 a_n1670_n3888# 0.848068f
C107 drain_left.t12 a_n1670_n3888# 0.46099f
C108 drain_left.t13 a_n1670_n3888# 0.46099f
C109 drain_left.n3 a_n1670_n3888# 4.17015f
C110 drain_left.t4 a_n1670_n3888# 0.46099f
C111 drain_left.t14 a_n1670_n3888# 0.46099f
C112 drain_left.n4 a_n1670_n3888# 4.16681f
C113 drain_left.n5 a_n1670_n3888# 0.848068f
C114 drain_left.n6 a_n1670_n3888# 2.10042f
C115 drain_left.t8 a_n1670_n3888# 0.46099f
C116 drain_left.t10 a_n1670_n3888# 0.46099f
C117 drain_left.n7 a_n1670_n3888# 4.17015f
C118 drain_left.t1 a_n1670_n3888# 0.46099f
C119 drain_left.t6 a_n1670_n3888# 0.46099f
C120 drain_left.n8 a_n1670_n3888# 4.16681f
C121 drain_left.n9 a_n1670_n3888# 0.878416f
C122 drain_left.t7 a_n1670_n3888# 0.46099f
C123 drain_left.t9 a_n1670_n3888# 0.46099f
C124 drain_left.n10 a_n1670_n3888# 4.16681f
C125 drain_left.n11 a_n1670_n3888# 0.433047f
C126 drain_left.t11 a_n1670_n3888# 0.46099f
C127 drain_left.t2 a_n1670_n3888# 0.46099f
C128 drain_left.n12 a_n1670_n3888# 4.1668f
C129 drain_left.n13 a_n1670_n3888# 0.751346f
C130 source.t24 a_n1670_n3888# 4.25416f
C131 source.n0 a_n1670_n3888# 1.95609f
C132 source.t20 a_n1670_n3888# 0.379611f
C133 source.t16 a_n1670_n3888# 0.379611f
C134 source.n1 a_n1670_n3888# 3.33457f
C135 source.n2 a_n1670_n3888# 0.409751f
C136 source.t26 a_n1670_n3888# 0.379611f
C137 source.t28 a_n1670_n3888# 0.379611f
C138 source.n3 a_n1670_n3888# 3.33457f
C139 source.n4 a_n1670_n3888# 0.409751f
C140 source.t17 a_n1670_n3888# 0.379611f
C141 source.t21 a_n1670_n3888# 0.379611f
C142 source.n5 a_n1670_n3888# 3.33457f
C143 source.n6 a_n1670_n3888# 0.409751f
C144 source.t18 a_n1670_n3888# 4.25416f
C145 source.n7 a_n1670_n3888# 0.526794f
C146 source.t9 a_n1670_n3888# 4.25416f
C147 source.n8 a_n1670_n3888# 0.526794f
C148 source.t8 a_n1670_n3888# 0.379611f
C149 source.t2 a_n1670_n3888# 0.379611f
C150 source.n9 a_n1670_n3888# 3.33457f
C151 source.n10 a_n1670_n3888# 0.409751f
C152 source.t11 a_n1670_n3888# 0.379611f
C153 source.t3 a_n1670_n3888# 0.379611f
C154 source.n11 a_n1670_n3888# 3.33457f
C155 source.n12 a_n1670_n3888# 0.409751f
C156 source.t7 a_n1670_n3888# 0.379611f
C157 source.t30 a_n1670_n3888# 0.379611f
C158 source.n13 a_n1670_n3888# 3.33457f
C159 source.n14 a_n1670_n3888# 0.409751f
C160 source.t0 a_n1670_n3888# 4.25416f
C161 source.n15 a_n1670_n3888# 2.4851f
C162 source.t14 a_n1670_n3888# 4.25416f
C163 source.n16 a_n1670_n3888# 2.4851f
C164 source.t15 a_n1670_n3888# 0.379611f
C165 source.t27 a_n1670_n3888# 0.379611f
C166 source.n17 a_n1670_n3888# 3.33456f
C167 source.n18 a_n1670_n3888# 0.409755f
C168 source.t25 a_n1670_n3888# 0.379611f
C169 source.t23 a_n1670_n3888# 0.379611f
C170 source.n19 a_n1670_n3888# 3.33456f
C171 source.n20 a_n1670_n3888# 0.409755f
C172 source.t19 a_n1670_n3888# 0.379611f
C173 source.t22 a_n1670_n3888# 0.379611f
C174 source.n21 a_n1670_n3888# 3.33456f
C175 source.n22 a_n1670_n3888# 0.409755f
C176 source.t29 a_n1670_n3888# 4.25416f
C177 source.n23 a_n1670_n3888# 0.526799f
C178 source.t6 a_n1670_n3888# 4.25416f
C179 source.n24 a_n1670_n3888# 0.526799f
C180 source.t10 a_n1670_n3888# 0.379611f
C181 source.t31 a_n1670_n3888# 0.379611f
C182 source.n25 a_n1670_n3888# 3.33456f
C183 source.n26 a_n1670_n3888# 0.409755f
C184 source.t1 a_n1670_n3888# 0.379611f
C185 source.t13 a_n1670_n3888# 0.379611f
C186 source.n27 a_n1670_n3888# 3.33456f
C187 source.n28 a_n1670_n3888# 0.409755f
C188 source.t5 a_n1670_n3888# 0.379611f
C189 source.t4 a_n1670_n3888# 0.379611f
C190 source.n29 a_n1670_n3888# 3.33456f
C191 source.n30 a_n1670_n3888# 0.409755f
C192 source.t12 a_n1670_n3888# 4.25416f
C193 source.n31 a_n1670_n3888# 0.700451f
C194 source.n32 a_n1670_n3888# 2.33644f
C195 plus.n0 a_n1670_n3888# 0.05529f
C196 plus.t4 a_n1670_n3888# 0.467945f
C197 plus.t6 a_n1670_n3888# 0.467945f
C198 plus.t8 a_n1670_n3888# 0.467945f
C199 plus.n1 a_n1670_n3888# 0.185422f
C200 plus.n2 a_n1670_n3888# 0.05529f
C201 plus.t9 a_n1670_n3888# 0.467945f
C202 plus.t14 a_n1670_n3888# 0.467945f
C203 plus.t5 a_n1670_n3888# 0.467945f
C204 plus.n3 a_n1670_n3888# 0.185422f
C205 plus.t7 a_n1670_n3888# 0.472762f
C206 plus.n4 a_n1670_n3888# 0.201925f
C207 plus.n5 a_n1670_n3888# 0.124475f
C208 plus.n6 a_n1670_n3888# 0.019364f
C209 plus.n7 a_n1670_n3888# 0.185422f
C210 plus.n8 a_n1670_n3888# 0.019364f
C211 plus.n9 a_n1670_n3888# 0.185422f
C212 plus.n10 a_n1670_n3888# 0.019364f
C213 plus.n11 a_n1670_n3888# 0.05529f
C214 plus.n12 a_n1670_n3888# 0.05529f
C215 plus.n13 a_n1670_n3888# 0.019364f
C216 plus.n14 a_n1670_n3888# 0.185422f
C217 plus.n15 a_n1670_n3888# 0.019364f
C218 plus.n16 a_n1670_n3888# 0.185422f
C219 plus.t13 a_n1670_n3888# 0.472762f
C220 plus.n17 a_n1670_n3888# 0.201844f
C221 plus.n18 a_n1670_n3888# 0.694312f
C222 plus.n19 a_n1670_n3888# 0.05529f
C223 plus.t10 a_n1670_n3888# 0.472762f
C224 plus.t15 a_n1670_n3888# 0.467945f
C225 plus.t12 a_n1670_n3888# 0.467945f
C226 plus.t0 a_n1670_n3888# 0.467945f
C227 plus.n20 a_n1670_n3888# 0.185422f
C228 plus.n21 a_n1670_n3888# 0.05529f
C229 plus.t11 a_n1670_n3888# 0.467945f
C230 plus.t1 a_n1670_n3888# 0.467945f
C231 plus.t3 a_n1670_n3888# 0.467945f
C232 plus.n22 a_n1670_n3888# 0.185422f
C233 plus.t2 a_n1670_n3888# 0.472762f
C234 plus.n23 a_n1670_n3888# 0.201925f
C235 plus.n24 a_n1670_n3888# 0.124475f
C236 plus.n25 a_n1670_n3888# 0.019364f
C237 plus.n26 a_n1670_n3888# 0.185422f
C238 plus.n27 a_n1670_n3888# 0.019364f
C239 plus.n28 a_n1670_n3888# 0.185422f
C240 plus.n29 a_n1670_n3888# 0.019364f
C241 plus.n30 a_n1670_n3888# 0.05529f
C242 plus.n31 a_n1670_n3888# 0.05529f
C243 plus.n32 a_n1670_n3888# 0.019364f
C244 plus.n33 a_n1670_n3888# 0.185422f
C245 plus.n34 a_n1670_n3888# 0.019364f
C246 plus.n35 a_n1670_n3888# 0.185422f
C247 plus.n36 a_n1670_n3888# 0.201844f
C248 plus.n37 a_n1670_n3888# 1.70642f
.ends

