* NGSPICE file created from diffpair470.ext - technology: sky130A

.subckt diffpair470 minus drain_right drain_left source plus
X0 drain_right minus source a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.8
X1 drain_left plus source a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.8
X2 drain_left plus source a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.8
X3 drain_right minus source a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.8
X4 a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X5 a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X6 a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X7 a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# a_n1168_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
.ends

