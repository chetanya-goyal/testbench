* NGSPICE file created from diffpair529.ext - technology: sky130A

.subckt diffpair529 minus drain_right drain_left source plus
X0 a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X1 drain_right.t23 minus.t0 source.t24 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X2 source.t6 plus.t0 drain_left.t23 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X3 drain_left.t22 plus.t1 source.t35 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X4 source.t37 plus.t2 drain_left.t21 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X5 drain_left.t20 plus.t3 source.t42 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X6 source.t14 minus.t1 drain_right.t22 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X7 source.t2 plus.t4 drain_left.t19 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X8 source.t20 minus.t2 drain_right.t21 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X9 source.t3 plus.t5 drain_left.t18 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X10 source.t47 plus.t6 drain_left.t17 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X11 source.t32 minus.t3 drain_right.t20 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X12 drain_right.t19 minus.t4 source.t12 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X13 source.t5 plus.t7 drain_left.t16 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X14 drain_left.t15 plus.t8 source.t1 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 drain_right.t18 minus.t5 source.t13 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X16 drain_right.t17 minus.t6 source.t31 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X17 source.t29 minus.t7 drain_right.t16 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X18 drain_left.t14 plus.t9 source.t4 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 drain_right.t15 minus.t8 source.t11 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X20 drain_left.t13 plus.t10 source.t41 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X21 source.t27 minus.t9 drain_right.t14 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X22 drain_left.t12 plus.t11 source.t38 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X23 drain_left.t11 plus.t12 source.t43 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X24 source.t46 plus.t13 drain_left.t10 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X25 source.t17 minus.t10 drain_right.t13 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X26 source.t28 minus.t11 drain_right.t12 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X27 drain_right.t11 minus.t12 source.t18 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X28 a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X29 source.t39 plus.t14 drain_left.t9 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X30 drain_left.t8 plus.t15 source.t7 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X31 source.t8 plus.t16 drain_left.t7 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X32 drain_left.t6 plus.t17 source.t45 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X33 drain_right.t10 minus.t13 source.t26 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X34 drain_right.t9 minus.t14 source.t23 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X35 a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X36 source.t15 minus.t15 drain_right.t8 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X37 drain_right.t7 minus.t16 source.t19 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X38 source.t34 minus.t17 drain_right.t6 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X39 drain_left.t5 plus.t18 source.t44 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X40 drain_right.t5 minus.t18 source.t22 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X41 source.t16 minus.t19 drain_right.t4 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X42 source.t25 minus.t20 drain_right.t3 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X43 drain_right.t2 minus.t21 source.t30 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X44 source.t10 plus.t19 drain_left.t4 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X45 source.t21 minus.t22 drain_right.t1 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X46 a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X47 drain_left.t3 plus.t20 source.t9 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X48 source.t36 plus.t21 drain_left.t2 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X49 drain_right.t0 minus.t23 source.t33 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X50 source.t40 plus.t22 drain_left.t1 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X51 drain_left.t0 plus.t23 source.t0 a_n2874_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
R0 minus.n9 minus.t13 827.924
R1 minus.n43 minus.t7 827.924
R2 minus.n8 minus.t1 801.567
R3 minus.n7 minus.t8 801.567
R4 minus.n13 minus.t19 801.567
R5 minus.n5 minus.t5 801.567
R6 minus.n18 minus.t10 801.567
R7 minus.n20 minus.t0 801.567
R8 minus.n3 minus.t11 801.567
R9 minus.n25 minus.t18 801.567
R10 minus.n1 minus.t3 801.567
R11 minus.n30 minus.t14 801.567
R12 minus.n32 minus.t22 801.567
R13 minus.n42 minus.t6 801.567
R14 minus.n41 minus.t17 801.567
R15 minus.n47 minus.t16 801.567
R16 minus.n39 minus.t9 801.567
R17 minus.n52 minus.t21 801.567
R18 minus.n54 minus.t20 801.567
R19 minus.n37 minus.t12 801.567
R20 minus.n59 minus.t2 801.567
R21 minus.n35 minus.t23 801.567
R22 minus.n64 minus.t15 801.567
R23 minus.n66 minus.t4 801.567
R24 minus.n33 minus.n32 161.3
R25 minus.n31 minus.n0 161.3
R26 minus.n30 minus.n29 161.3
R27 minus.n28 minus.n1 161.3
R28 minus.n27 minus.n26 161.3
R29 minus.n25 minus.n2 161.3
R30 minus.n24 minus.n23 161.3
R31 minus.n22 minus.n3 161.3
R32 minus.n21 minus.n20 161.3
R33 minus.n19 minus.n4 161.3
R34 minus.n18 minus.n17 161.3
R35 minus.n16 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n6 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n10 minus.n7 161.3
R40 minus.n67 minus.n66 161.3
R41 minus.n65 minus.n34 161.3
R42 minus.n64 minus.n63 161.3
R43 minus.n62 minus.n35 161.3
R44 minus.n61 minus.n60 161.3
R45 minus.n59 minus.n36 161.3
R46 minus.n58 minus.n57 161.3
R47 minus.n56 minus.n37 161.3
R48 minus.n55 minus.n54 161.3
R49 minus.n53 minus.n38 161.3
R50 minus.n52 minus.n51 161.3
R51 minus.n50 minus.n39 161.3
R52 minus.n49 minus.n48 161.3
R53 minus.n47 minus.n40 161.3
R54 minus.n46 minus.n45 161.3
R55 minus.n44 minus.n41 161.3
R56 minus.n8 minus.n7 48.2005
R57 minus.n18 minus.n5 48.2005
R58 minus.n20 minus.n3 48.2005
R59 minus.n30 minus.n1 48.2005
R60 minus.n42 minus.n41 48.2005
R61 minus.n52 minus.n39 48.2005
R62 minus.n54 minus.n37 48.2005
R63 minus.n64 minus.n35 48.2005
R64 minus.n14 minus.n13 47.4702
R65 minus.n25 minus.n24 47.4702
R66 minus.n48 minus.n47 47.4702
R67 minus.n59 minus.n58 47.4702
R68 minus.n32 minus.n31 46.0096
R69 minus.n66 minus.n65 46.0096
R70 minus.n10 minus.n9 45.0871
R71 minus.n44 minus.n43 45.0871
R72 minus.n68 minus.n33 42.3073
R73 minus.n13 minus.n12 25.5611
R74 minus.n26 minus.n25 25.5611
R75 minus.n47 minus.n46 25.5611
R76 minus.n60 minus.n59 25.5611
R77 minus.n20 minus.n19 24.1005
R78 minus.n19 minus.n18 24.1005
R79 minus.n53 minus.n52 24.1005
R80 minus.n54 minus.n53 24.1005
R81 minus.n12 minus.n7 22.6399
R82 minus.n26 minus.n1 22.6399
R83 minus.n46 minus.n41 22.6399
R84 minus.n60 minus.n35 22.6399
R85 minus.n9 minus.n8 14.1472
R86 minus.n43 minus.n42 14.1472
R87 minus.n68 minus.n67 6.52702
R88 minus.n31 minus.n30 2.19141
R89 minus.n65 minus.n64 2.19141
R90 minus.n14 minus.n5 0.730803
R91 minus.n24 minus.n3 0.730803
R92 minus.n48 minus.n39 0.730803
R93 minus.n58 minus.n37 0.730803
R94 minus.n33 minus.n0 0.189894
R95 minus.n29 minus.n0 0.189894
R96 minus.n29 minus.n28 0.189894
R97 minus.n28 minus.n27 0.189894
R98 minus.n27 minus.n2 0.189894
R99 minus.n23 minus.n2 0.189894
R100 minus.n23 minus.n22 0.189894
R101 minus.n22 minus.n21 0.189894
R102 minus.n21 minus.n4 0.189894
R103 minus.n17 minus.n4 0.189894
R104 minus.n17 minus.n16 0.189894
R105 minus.n16 minus.n15 0.189894
R106 minus.n15 minus.n6 0.189894
R107 minus.n11 minus.n6 0.189894
R108 minus.n11 minus.n10 0.189894
R109 minus.n45 minus.n44 0.189894
R110 minus.n45 minus.n40 0.189894
R111 minus.n49 minus.n40 0.189894
R112 minus.n50 minus.n49 0.189894
R113 minus.n51 minus.n50 0.189894
R114 minus.n51 minus.n38 0.189894
R115 minus.n55 minus.n38 0.189894
R116 minus.n56 minus.n55 0.189894
R117 minus.n57 minus.n56 0.189894
R118 minus.n57 minus.n36 0.189894
R119 minus.n61 minus.n36 0.189894
R120 minus.n62 minus.n61 0.189894
R121 minus.n63 minus.n62 0.189894
R122 minus.n63 minus.n34 0.189894
R123 minus.n67 minus.n34 0.189894
R124 minus minus.n68 0.188
R125 source.n11 source.t47 45.521
R126 source.n12 source.t26 45.521
R127 source.n23 source.t21 45.521
R128 source.n47 source.t12 45.5208
R129 source.n36 source.t29 45.5208
R130 source.n35 source.t42 45.5208
R131 source.n24 source.t40 45.5208
R132 source.n0 source.t35 45.5208
R133 source.n2 source.n1 44.201
R134 source.n4 source.n3 44.201
R135 source.n6 source.n5 44.201
R136 source.n8 source.n7 44.201
R137 source.n10 source.n9 44.201
R138 source.n14 source.n13 44.201
R139 source.n16 source.n15 44.201
R140 source.n18 source.n17 44.201
R141 source.n20 source.n19 44.201
R142 source.n22 source.n21 44.201
R143 source.n46 source.n45 44.2008
R144 source.n44 source.n43 44.2008
R145 source.n42 source.n41 44.2008
R146 source.n40 source.n39 44.2008
R147 source.n38 source.n37 44.2008
R148 source.n34 source.n33 44.2008
R149 source.n32 source.n31 44.2008
R150 source.n30 source.n29 44.2008
R151 source.n28 source.n27 44.2008
R152 source.n26 source.n25 44.2008
R153 source.n24 source.n23 24.276
R154 source.n48 source.n0 18.6553
R155 source.n48 source.n47 5.62119
R156 source.n45 source.t33 1.3205
R157 source.n45 source.t15 1.3205
R158 source.n43 source.t18 1.3205
R159 source.n43 source.t20 1.3205
R160 source.n41 source.t30 1.3205
R161 source.n41 source.t25 1.3205
R162 source.n39 source.t19 1.3205
R163 source.n39 source.t27 1.3205
R164 source.n37 source.t31 1.3205
R165 source.n37 source.t34 1.3205
R166 source.n33 source.t43 1.3205
R167 source.n33 source.t6 1.3205
R168 source.n31 source.t1 1.3205
R169 source.n31 source.t5 1.3205
R170 source.n29 source.t38 1.3205
R171 source.n29 source.t8 1.3205
R172 source.n27 source.t7 1.3205
R173 source.n27 source.t3 1.3205
R174 source.n25 source.t4 1.3205
R175 source.n25 source.t39 1.3205
R176 source.n1 source.t45 1.3205
R177 source.n1 source.t37 1.3205
R178 source.n3 source.t9 1.3205
R179 source.n3 source.t2 1.3205
R180 source.n5 source.t0 1.3205
R181 source.n5 source.t46 1.3205
R182 source.n7 source.t41 1.3205
R183 source.n7 source.t10 1.3205
R184 source.n9 source.t44 1.3205
R185 source.n9 source.t36 1.3205
R186 source.n13 source.t11 1.3205
R187 source.n13 source.t14 1.3205
R188 source.n15 source.t13 1.3205
R189 source.n15 source.t16 1.3205
R190 source.n17 source.t24 1.3205
R191 source.n17 source.t17 1.3205
R192 source.n19 source.t22 1.3205
R193 source.n19 source.t28 1.3205
R194 source.n21 source.t23 1.3205
R195 source.n21 source.t32 1.3205
R196 source.n23 source.n22 0.716017
R197 source.n22 source.n20 0.716017
R198 source.n20 source.n18 0.716017
R199 source.n18 source.n16 0.716017
R200 source.n16 source.n14 0.716017
R201 source.n14 source.n12 0.716017
R202 source.n11 source.n10 0.716017
R203 source.n10 source.n8 0.716017
R204 source.n8 source.n6 0.716017
R205 source.n6 source.n4 0.716017
R206 source.n4 source.n2 0.716017
R207 source.n2 source.n0 0.716017
R208 source.n26 source.n24 0.716017
R209 source.n28 source.n26 0.716017
R210 source.n30 source.n28 0.716017
R211 source.n32 source.n30 0.716017
R212 source.n34 source.n32 0.716017
R213 source.n35 source.n34 0.716017
R214 source.n38 source.n36 0.716017
R215 source.n40 source.n38 0.716017
R216 source.n42 source.n40 0.716017
R217 source.n44 source.n42 0.716017
R218 source.n46 source.n44 0.716017
R219 source.n47 source.n46 0.716017
R220 source.n12 source.n11 0.470328
R221 source.n36 source.n35 0.470328
R222 source source.n48 0.188
R223 drain_right.n13 drain_right.n11 61.5952
R224 drain_right.n7 drain_right.n5 61.5951
R225 drain_right.n2 drain_right.n0 61.5951
R226 drain_right.n13 drain_right.n12 60.8798
R227 drain_right.n15 drain_right.n14 60.8798
R228 drain_right.n17 drain_right.n16 60.8798
R229 drain_right.n19 drain_right.n18 60.8798
R230 drain_right.n21 drain_right.n20 60.8798
R231 drain_right.n7 drain_right.n6 60.8796
R232 drain_right.n9 drain_right.n8 60.8796
R233 drain_right.n4 drain_right.n3 60.8796
R234 drain_right.n2 drain_right.n1 60.8796
R235 drain_right drain_right.n10 35.884
R236 drain_right drain_right.n21 6.36873
R237 drain_right.n5 drain_right.t8 1.3205
R238 drain_right.n5 drain_right.t19 1.3205
R239 drain_right.n6 drain_right.t21 1.3205
R240 drain_right.n6 drain_right.t0 1.3205
R241 drain_right.n8 drain_right.t3 1.3205
R242 drain_right.n8 drain_right.t11 1.3205
R243 drain_right.n3 drain_right.t14 1.3205
R244 drain_right.n3 drain_right.t2 1.3205
R245 drain_right.n1 drain_right.t6 1.3205
R246 drain_right.n1 drain_right.t7 1.3205
R247 drain_right.n0 drain_right.t16 1.3205
R248 drain_right.n0 drain_right.t17 1.3205
R249 drain_right.n11 drain_right.t22 1.3205
R250 drain_right.n11 drain_right.t10 1.3205
R251 drain_right.n12 drain_right.t4 1.3205
R252 drain_right.n12 drain_right.t15 1.3205
R253 drain_right.n14 drain_right.t13 1.3205
R254 drain_right.n14 drain_right.t18 1.3205
R255 drain_right.n16 drain_right.t12 1.3205
R256 drain_right.n16 drain_right.t23 1.3205
R257 drain_right.n18 drain_right.t20 1.3205
R258 drain_right.n18 drain_right.t5 1.3205
R259 drain_right.n20 drain_right.t1 1.3205
R260 drain_right.n20 drain_right.t9 1.3205
R261 drain_right.n9 drain_right.n7 0.716017
R262 drain_right.n4 drain_right.n2 0.716017
R263 drain_right.n21 drain_right.n19 0.716017
R264 drain_right.n19 drain_right.n17 0.716017
R265 drain_right.n17 drain_right.n15 0.716017
R266 drain_right.n15 drain_right.n13 0.716017
R267 drain_right.n10 drain_right.n9 0.302913
R268 drain_right.n10 drain_right.n4 0.302913
R269 plus.n11 plus.t6 827.924
R270 plus.n45 plus.t3 827.924
R271 plus.n32 plus.t1 801.567
R272 plus.n30 plus.t2 801.567
R273 plus.n29 plus.t17 801.567
R274 plus.n3 plus.t4 801.567
R275 plus.n23 plus.t20 801.567
R276 plus.n22 plus.t13 801.567
R277 plus.n6 plus.t23 801.567
R278 plus.n17 plus.t19 801.567
R279 plus.n15 plus.t10 801.567
R280 plus.n9 plus.t21 801.567
R281 plus.n10 plus.t18 801.567
R282 plus.n66 plus.t22 801.567
R283 plus.n64 plus.t9 801.567
R284 plus.n63 plus.t14 801.567
R285 plus.n37 plus.t15 801.567
R286 plus.n57 plus.t5 801.567
R287 plus.n56 plus.t11 801.567
R288 plus.n40 plus.t16 801.567
R289 plus.n51 plus.t8 801.567
R290 plus.n49 plus.t7 801.567
R291 plus.n43 plus.t12 801.567
R292 plus.n44 plus.t0 801.567
R293 plus.n12 plus.n9 161.3
R294 plus.n14 plus.n13 161.3
R295 plus.n15 plus.n8 161.3
R296 plus.n16 plus.n7 161.3
R297 plus.n18 plus.n17 161.3
R298 plus.n19 plus.n6 161.3
R299 plus.n21 plus.n20 161.3
R300 plus.n22 plus.n5 161.3
R301 plus.n23 plus.n4 161.3
R302 plus.n25 plus.n24 161.3
R303 plus.n26 plus.n3 161.3
R304 plus.n28 plus.n27 161.3
R305 plus.n29 plus.n2 161.3
R306 plus.n30 plus.n1 161.3
R307 plus.n31 plus.n0 161.3
R308 plus.n33 plus.n32 161.3
R309 plus.n46 plus.n43 161.3
R310 plus.n48 plus.n47 161.3
R311 plus.n49 plus.n42 161.3
R312 plus.n50 plus.n41 161.3
R313 plus.n52 plus.n51 161.3
R314 plus.n53 plus.n40 161.3
R315 plus.n55 plus.n54 161.3
R316 plus.n56 plus.n39 161.3
R317 plus.n57 plus.n38 161.3
R318 plus.n59 plus.n58 161.3
R319 plus.n60 plus.n37 161.3
R320 plus.n62 plus.n61 161.3
R321 plus.n63 plus.n36 161.3
R322 plus.n64 plus.n35 161.3
R323 plus.n65 plus.n34 161.3
R324 plus.n67 plus.n66 161.3
R325 plus.n30 plus.n29 48.2005
R326 plus.n23 plus.n22 48.2005
R327 plus.n17 plus.n6 48.2005
R328 plus.n10 plus.n9 48.2005
R329 plus.n64 plus.n63 48.2005
R330 plus.n57 plus.n56 48.2005
R331 plus.n51 plus.n40 48.2005
R332 plus.n44 plus.n43 48.2005
R333 plus.n24 plus.n3 47.4702
R334 plus.n16 plus.n15 47.4702
R335 plus.n58 plus.n37 47.4702
R336 plus.n50 plus.n49 47.4702
R337 plus.n32 plus.n31 46.0096
R338 plus.n66 plus.n65 46.0096
R339 plus.n12 plus.n11 45.0871
R340 plus.n46 plus.n45 45.0871
R341 plus plus.n67 35.0521
R342 plus.n28 plus.n3 25.5611
R343 plus.n15 plus.n14 25.5611
R344 plus.n62 plus.n37 25.5611
R345 plus.n49 plus.n48 25.5611
R346 plus.n21 plus.n6 24.1005
R347 plus.n22 plus.n21 24.1005
R348 plus.n56 plus.n55 24.1005
R349 plus.n55 plus.n40 24.1005
R350 plus.n29 plus.n28 22.6399
R351 plus.n14 plus.n9 22.6399
R352 plus.n63 plus.n62 22.6399
R353 plus.n48 plus.n43 22.6399
R354 plus.n11 plus.n10 14.1472
R355 plus.n45 plus.n44 14.1472
R356 plus plus.n33 13.3073
R357 plus.n31 plus.n30 2.19141
R358 plus.n65 plus.n64 2.19141
R359 plus.n24 plus.n23 0.730803
R360 plus.n17 plus.n16 0.730803
R361 plus.n58 plus.n57 0.730803
R362 plus.n51 plus.n50 0.730803
R363 plus.n13 plus.n12 0.189894
R364 plus.n13 plus.n8 0.189894
R365 plus.n8 plus.n7 0.189894
R366 plus.n18 plus.n7 0.189894
R367 plus.n19 plus.n18 0.189894
R368 plus.n20 plus.n19 0.189894
R369 plus.n20 plus.n5 0.189894
R370 plus.n5 plus.n4 0.189894
R371 plus.n25 plus.n4 0.189894
R372 plus.n26 plus.n25 0.189894
R373 plus.n27 plus.n26 0.189894
R374 plus.n27 plus.n2 0.189894
R375 plus.n2 plus.n1 0.189894
R376 plus.n1 plus.n0 0.189894
R377 plus.n33 plus.n0 0.189894
R378 plus.n67 plus.n34 0.189894
R379 plus.n35 plus.n34 0.189894
R380 plus.n36 plus.n35 0.189894
R381 plus.n61 plus.n36 0.189894
R382 plus.n61 plus.n60 0.189894
R383 plus.n60 plus.n59 0.189894
R384 plus.n59 plus.n38 0.189894
R385 plus.n39 plus.n38 0.189894
R386 plus.n54 plus.n39 0.189894
R387 plus.n54 plus.n53 0.189894
R388 plus.n53 plus.n52 0.189894
R389 plus.n52 plus.n41 0.189894
R390 plus.n42 plus.n41 0.189894
R391 plus.n47 plus.n42 0.189894
R392 plus.n47 plus.n46 0.189894
R393 drain_left.n13 drain_left.n11 61.5953
R394 drain_left.n7 drain_left.n5 61.5951
R395 drain_left.n2 drain_left.n0 61.5951
R396 drain_left.n19 drain_left.n18 60.8798
R397 drain_left.n17 drain_left.n16 60.8798
R398 drain_left.n15 drain_left.n14 60.8798
R399 drain_left.n13 drain_left.n12 60.8798
R400 drain_left.n21 drain_left.n20 60.8796
R401 drain_left.n7 drain_left.n6 60.8796
R402 drain_left.n9 drain_left.n8 60.8796
R403 drain_left.n4 drain_left.n3 60.8796
R404 drain_left.n2 drain_left.n1 60.8796
R405 drain_left drain_left.n10 36.4372
R406 drain_left drain_left.n21 6.36873
R407 drain_left.n5 drain_left.t23 1.3205
R408 drain_left.n5 drain_left.t20 1.3205
R409 drain_left.n6 drain_left.t16 1.3205
R410 drain_left.n6 drain_left.t11 1.3205
R411 drain_left.n8 drain_left.t7 1.3205
R412 drain_left.n8 drain_left.t15 1.3205
R413 drain_left.n3 drain_left.t18 1.3205
R414 drain_left.n3 drain_left.t12 1.3205
R415 drain_left.n1 drain_left.t9 1.3205
R416 drain_left.n1 drain_left.t8 1.3205
R417 drain_left.n0 drain_left.t1 1.3205
R418 drain_left.n0 drain_left.t14 1.3205
R419 drain_left.n20 drain_left.t21 1.3205
R420 drain_left.n20 drain_left.t22 1.3205
R421 drain_left.n18 drain_left.t19 1.3205
R422 drain_left.n18 drain_left.t6 1.3205
R423 drain_left.n16 drain_left.t10 1.3205
R424 drain_left.n16 drain_left.t3 1.3205
R425 drain_left.n14 drain_left.t4 1.3205
R426 drain_left.n14 drain_left.t0 1.3205
R427 drain_left.n12 drain_left.t2 1.3205
R428 drain_left.n12 drain_left.t13 1.3205
R429 drain_left.n11 drain_left.t17 1.3205
R430 drain_left.n11 drain_left.t5 1.3205
R431 drain_left.n9 drain_left.n7 0.716017
R432 drain_left.n4 drain_left.n2 0.716017
R433 drain_left.n15 drain_left.n13 0.716017
R434 drain_left.n17 drain_left.n15 0.716017
R435 drain_left.n19 drain_left.n17 0.716017
R436 drain_left.n21 drain_left.n19 0.716017
R437 drain_left.n10 drain_left.n9 0.302913
R438 drain_left.n10 drain_left.n4 0.302913
C0 plus source 14.937599f
C1 minus source 14.923501f
C2 drain_left drain_right 1.55979f
C3 plus minus 7.29709f
C4 source drain_left 41.4001f
C5 plus drain_left 15.2702f
C6 source drain_right 41.4016f
C7 plus drain_right 0.443411f
C8 minus drain_left 0.173624f
C9 minus drain_right 14.983901f
C10 drain_right a_n2874_n3888# 8.09821f
C11 drain_left a_n2874_n3888# 8.5075f
C12 source a_n2874_n3888# 10.91761f
C13 minus a_n2874_n3888# 11.722912f
C14 plus a_n2874_n3888# 13.85483f
C15 drain_left.t1 a_n2874_n3888# 0.35011f
C16 drain_left.t14 a_n2874_n3888# 0.35011f
C17 drain_left.n0 a_n2874_n3888# 3.16912f
C18 drain_left.t9 a_n2874_n3888# 0.35011f
C19 drain_left.t8 a_n2874_n3888# 0.35011f
C20 drain_left.n1 a_n2874_n3888# 3.16458f
C21 drain_left.n2 a_n2874_n3888# 0.763603f
C22 drain_left.t18 a_n2874_n3888# 0.35011f
C23 drain_left.t12 a_n2874_n3888# 0.35011f
C24 drain_left.n3 a_n2874_n3888# 3.16458f
C25 drain_left.n4 a_n2874_n3888# 0.341066f
C26 drain_left.t23 a_n2874_n3888# 0.35011f
C27 drain_left.t20 a_n2874_n3888# 0.35011f
C28 drain_left.n5 a_n2874_n3888# 3.16912f
C29 drain_left.t16 a_n2874_n3888# 0.35011f
C30 drain_left.t11 a_n2874_n3888# 0.35011f
C31 drain_left.n6 a_n2874_n3888# 3.16458f
C32 drain_left.n7 a_n2874_n3888# 0.763603f
C33 drain_left.t7 a_n2874_n3888# 0.35011f
C34 drain_left.t15 a_n2874_n3888# 0.35011f
C35 drain_left.n8 a_n2874_n3888# 3.16458f
C36 drain_left.n9 a_n2874_n3888# 0.341066f
C37 drain_left.n10 a_n2874_n3888# 1.98728f
C38 drain_left.t17 a_n2874_n3888# 0.35011f
C39 drain_left.t5 a_n2874_n3888# 0.35011f
C40 drain_left.n11 a_n2874_n3888# 3.16912f
C41 drain_left.t2 a_n2874_n3888# 0.35011f
C42 drain_left.t13 a_n2874_n3888# 0.35011f
C43 drain_left.n12 a_n2874_n3888# 3.16459f
C44 drain_left.n13 a_n2874_n3888# 0.763598f
C45 drain_left.t4 a_n2874_n3888# 0.35011f
C46 drain_left.t0 a_n2874_n3888# 0.35011f
C47 drain_left.n14 a_n2874_n3888# 3.16459f
C48 drain_left.n15 a_n2874_n3888# 0.378116f
C49 drain_left.t10 a_n2874_n3888# 0.35011f
C50 drain_left.t3 a_n2874_n3888# 0.35011f
C51 drain_left.n16 a_n2874_n3888# 3.16459f
C52 drain_left.n17 a_n2874_n3888# 0.378116f
C53 drain_left.t19 a_n2874_n3888# 0.35011f
C54 drain_left.t6 a_n2874_n3888# 0.35011f
C55 drain_left.n18 a_n2874_n3888# 3.16459f
C56 drain_left.n19 a_n2874_n3888# 0.378116f
C57 drain_left.t21 a_n2874_n3888# 0.35011f
C58 drain_left.t22 a_n2874_n3888# 0.35011f
C59 drain_left.n20 a_n2874_n3888# 3.16458f
C60 drain_left.n21 a_n2874_n3888# 0.631887f
C61 plus.n0 a_n2874_n3888# 0.043872f
C62 plus.t1 a_n2874_n3888# 0.935032f
C63 plus.t2 a_n2874_n3888# 0.935032f
C64 plus.n1 a_n2874_n3888# 0.043872f
C65 plus.t17 a_n2874_n3888# 0.935032f
C66 plus.n2 a_n2874_n3888# 0.043872f
C67 plus.t4 a_n2874_n3888# 0.935032f
C68 plus.n3 a_n2874_n3888# 0.368853f
C69 plus.n4 a_n2874_n3888# 0.043872f
C70 plus.t20 a_n2874_n3888# 0.935032f
C71 plus.t13 a_n2874_n3888# 0.935032f
C72 plus.n5 a_n2874_n3888# 0.043872f
C73 plus.t23 a_n2874_n3888# 0.935032f
C74 plus.n6 a_n2874_n3888# 0.368718f
C75 plus.n7 a_n2874_n3888# 0.043872f
C76 plus.t19 a_n2874_n3888# 0.935032f
C77 plus.t10 a_n2874_n3888# 0.935032f
C78 plus.n8 a_n2874_n3888# 0.043872f
C79 plus.t21 a_n2874_n3888# 0.935032f
C80 plus.n9 a_n2874_n3888# 0.368448f
C81 plus.t18 a_n2874_n3888# 0.935032f
C82 plus.n10 a_n2874_n3888# 0.373639f
C83 plus.t6 a_n2874_n3888# 0.946626f
C84 plus.n11 a_n2874_n3888# 0.354098f
C85 plus.n12 a_n2874_n3888# 0.178138f
C86 plus.n13 a_n2874_n3888# 0.043872f
C87 plus.n14 a_n2874_n3888# 0.009955f
C88 plus.n15 a_n2874_n3888# 0.368853f
C89 plus.n16 a_n2874_n3888# 0.009955f
C90 plus.n17 a_n2874_n3888# 0.36439f
C91 plus.n18 a_n2874_n3888# 0.043872f
C92 plus.n19 a_n2874_n3888# 0.043872f
C93 plus.n20 a_n2874_n3888# 0.043872f
C94 plus.n21 a_n2874_n3888# 0.009955f
C95 plus.n22 a_n2874_n3888# 0.368718f
C96 plus.n23 a_n2874_n3888# 0.36439f
C97 plus.n24 a_n2874_n3888# 0.009955f
C98 plus.n25 a_n2874_n3888# 0.043872f
C99 plus.n26 a_n2874_n3888# 0.043872f
C100 plus.n27 a_n2874_n3888# 0.043872f
C101 plus.n28 a_n2874_n3888# 0.009955f
C102 plus.n29 a_n2874_n3888# 0.368448f
C103 plus.n30 a_n2874_n3888# 0.364661f
C104 plus.n31 a_n2874_n3888# 0.009955f
C105 plus.n32 a_n2874_n3888# 0.363849f
C106 plus.n33 a_n2874_n3888# 0.557192f
C107 plus.n34 a_n2874_n3888# 0.043872f
C108 plus.t22 a_n2874_n3888# 0.935032f
C109 plus.n35 a_n2874_n3888# 0.043872f
C110 plus.t9 a_n2874_n3888# 0.935032f
C111 plus.n36 a_n2874_n3888# 0.043872f
C112 plus.t14 a_n2874_n3888# 0.935032f
C113 plus.t15 a_n2874_n3888# 0.935032f
C114 plus.n37 a_n2874_n3888# 0.368853f
C115 plus.n38 a_n2874_n3888# 0.043872f
C116 plus.t5 a_n2874_n3888# 0.935032f
C117 plus.n39 a_n2874_n3888# 0.043872f
C118 plus.t11 a_n2874_n3888# 0.935032f
C119 plus.t16 a_n2874_n3888# 0.935032f
C120 plus.n40 a_n2874_n3888# 0.368718f
C121 plus.n41 a_n2874_n3888# 0.043872f
C122 plus.t8 a_n2874_n3888# 0.935032f
C123 plus.n42 a_n2874_n3888# 0.043872f
C124 plus.t7 a_n2874_n3888# 0.935032f
C125 plus.t12 a_n2874_n3888# 0.935032f
C126 plus.n43 a_n2874_n3888# 0.368448f
C127 plus.t3 a_n2874_n3888# 0.946626f
C128 plus.t0 a_n2874_n3888# 0.935032f
C129 plus.n44 a_n2874_n3888# 0.373639f
C130 plus.n45 a_n2874_n3888# 0.354098f
C131 plus.n46 a_n2874_n3888# 0.178138f
C132 plus.n47 a_n2874_n3888# 0.043872f
C133 plus.n48 a_n2874_n3888# 0.009955f
C134 plus.n49 a_n2874_n3888# 0.368853f
C135 plus.n50 a_n2874_n3888# 0.009955f
C136 plus.n51 a_n2874_n3888# 0.36439f
C137 plus.n52 a_n2874_n3888# 0.043872f
C138 plus.n53 a_n2874_n3888# 0.043872f
C139 plus.n54 a_n2874_n3888# 0.043872f
C140 plus.n55 a_n2874_n3888# 0.009955f
C141 plus.n56 a_n2874_n3888# 0.368718f
C142 plus.n57 a_n2874_n3888# 0.36439f
C143 plus.n58 a_n2874_n3888# 0.009955f
C144 plus.n59 a_n2874_n3888# 0.043872f
C145 plus.n60 a_n2874_n3888# 0.043872f
C146 plus.n61 a_n2874_n3888# 0.043872f
C147 plus.n62 a_n2874_n3888# 0.009955f
C148 plus.n63 a_n2874_n3888# 0.368448f
C149 plus.n64 a_n2874_n3888# 0.364661f
C150 plus.n65 a_n2874_n3888# 0.009955f
C151 plus.n66 a_n2874_n3888# 0.363849f
C152 plus.n67 a_n2874_n3888# 1.63664f
C153 drain_right.t16 a_n2874_n3888# 0.348969f
C154 drain_right.t17 a_n2874_n3888# 0.348969f
C155 drain_right.n0 a_n2874_n3888# 3.15878f
C156 drain_right.t6 a_n2874_n3888# 0.348969f
C157 drain_right.t7 a_n2874_n3888# 0.348969f
C158 drain_right.n1 a_n2874_n3888# 3.15427f
C159 drain_right.n2 a_n2874_n3888# 0.761114f
C160 drain_right.t14 a_n2874_n3888# 0.348969f
C161 drain_right.t2 a_n2874_n3888# 0.348969f
C162 drain_right.n3 a_n2874_n3888# 3.15427f
C163 drain_right.n4 a_n2874_n3888# 0.339954f
C164 drain_right.t8 a_n2874_n3888# 0.348969f
C165 drain_right.t19 a_n2874_n3888# 0.348969f
C166 drain_right.n5 a_n2874_n3888# 3.15878f
C167 drain_right.t21 a_n2874_n3888# 0.348969f
C168 drain_right.t0 a_n2874_n3888# 0.348969f
C169 drain_right.n6 a_n2874_n3888# 3.15427f
C170 drain_right.n7 a_n2874_n3888# 0.761114f
C171 drain_right.t3 a_n2874_n3888# 0.348969f
C172 drain_right.t11 a_n2874_n3888# 0.348969f
C173 drain_right.n8 a_n2874_n3888# 3.15427f
C174 drain_right.n9 a_n2874_n3888# 0.339954f
C175 drain_right.n10 a_n2874_n3888# 1.92051f
C176 drain_right.t22 a_n2874_n3888# 0.348969f
C177 drain_right.t10 a_n2874_n3888# 0.348969f
C178 drain_right.n11 a_n2874_n3888# 3.15878f
C179 drain_right.t4 a_n2874_n3888# 0.348969f
C180 drain_right.t15 a_n2874_n3888# 0.348969f
C181 drain_right.n12 a_n2874_n3888# 3.15427f
C182 drain_right.n13 a_n2874_n3888# 0.76112f
C183 drain_right.t13 a_n2874_n3888# 0.348969f
C184 drain_right.t18 a_n2874_n3888# 0.348969f
C185 drain_right.n14 a_n2874_n3888# 3.15427f
C186 drain_right.n15 a_n2874_n3888# 0.376883f
C187 drain_right.t12 a_n2874_n3888# 0.348969f
C188 drain_right.t23 a_n2874_n3888# 0.348969f
C189 drain_right.n16 a_n2874_n3888# 3.15427f
C190 drain_right.n17 a_n2874_n3888# 0.376883f
C191 drain_right.t20 a_n2874_n3888# 0.348969f
C192 drain_right.t5 a_n2874_n3888# 0.348969f
C193 drain_right.n18 a_n2874_n3888# 3.15427f
C194 drain_right.n19 a_n2874_n3888# 0.376883f
C195 drain_right.t1 a_n2874_n3888# 0.348969f
C196 drain_right.t9 a_n2874_n3888# 0.348969f
C197 drain_right.n20 a_n2874_n3888# 3.15427f
C198 drain_right.n21 a_n2874_n3888# 0.629816f
C199 source.t35 a_n2874_n3888# 3.48083f
C200 source.n0 a_n2874_n3888# 1.63572f
C201 source.t45 a_n2874_n3888# 0.310605f
C202 source.t37 a_n2874_n3888# 0.310605f
C203 source.n1 a_n2874_n3888# 2.7284f
C204 source.n2 a_n2874_n3888# 0.378938f
C205 source.t9 a_n2874_n3888# 0.310605f
C206 source.t2 a_n2874_n3888# 0.310605f
C207 source.n3 a_n2874_n3888# 2.7284f
C208 source.n4 a_n2874_n3888# 0.378938f
C209 source.t0 a_n2874_n3888# 0.310605f
C210 source.t46 a_n2874_n3888# 0.310605f
C211 source.n5 a_n2874_n3888# 2.7284f
C212 source.n6 a_n2874_n3888# 0.378938f
C213 source.t41 a_n2874_n3888# 0.310605f
C214 source.t10 a_n2874_n3888# 0.310605f
C215 source.n7 a_n2874_n3888# 2.7284f
C216 source.n8 a_n2874_n3888# 0.378938f
C217 source.t44 a_n2874_n3888# 0.310605f
C218 source.t36 a_n2874_n3888# 0.310605f
C219 source.n9 a_n2874_n3888# 2.7284f
C220 source.n10 a_n2874_n3888# 0.378938f
C221 source.t47 a_n2874_n3888# 3.48083f
C222 source.n11 a_n2874_n3888# 0.452869f
C223 source.t26 a_n2874_n3888# 3.48083f
C224 source.n12 a_n2874_n3888# 0.452869f
C225 source.t11 a_n2874_n3888# 0.310605f
C226 source.t14 a_n2874_n3888# 0.310605f
C227 source.n13 a_n2874_n3888# 2.7284f
C228 source.n14 a_n2874_n3888# 0.378938f
C229 source.t13 a_n2874_n3888# 0.310605f
C230 source.t16 a_n2874_n3888# 0.310605f
C231 source.n15 a_n2874_n3888# 2.7284f
C232 source.n16 a_n2874_n3888# 0.378938f
C233 source.t24 a_n2874_n3888# 0.310605f
C234 source.t17 a_n2874_n3888# 0.310605f
C235 source.n17 a_n2874_n3888# 2.7284f
C236 source.n18 a_n2874_n3888# 0.378938f
C237 source.t22 a_n2874_n3888# 0.310605f
C238 source.t28 a_n2874_n3888# 0.310605f
C239 source.n19 a_n2874_n3888# 2.7284f
C240 source.n20 a_n2874_n3888# 0.378938f
C241 source.t23 a_n2874_n3888# 0.310605f
C242 source.t32 a_n2874_n3888# 0.310605f
C243 source.n21 a_n2874_n3888# 2.7284f
C244 source.n22 a_n2874_n3888# 0.378938f
C245 source.t21 a_n2874_n3888# 3.48083f
C246 source.n23 a_n2874_n3888# 2.07702f
C247 source.t40 a_n2874_n3888# 3.48083f
C248 source.n24 a_n2874_n3888# 2.07703f
C249 source.t4 a_n2874_n3888# 0.310605f
C250 source.t39 a_n2874_n3888# 0.310605f
C251 source.n25 a_n2874_n3888# 2.7284f
C252 source.n26 a_n2874_n3888# 0.378942f
C253 source.t7 a_n2874_n3888# 0.310605f
C254 source.t3 a_n2874_n3888# 0.310605f
C255 source.n27 a_n2874_n3888# 2.7284f
C256 source.n28 a_n2874_n3888# 0.378942f
C257 source.t38 a_n2874_n3888# 0.310605f
C258 source.t8 a_n2874_n3888# 0.310605f
C259 source.n29 a_n2874_n3888# 2.7284f
C260 source.n30 a_n2874_n3888# 0.378942f
C261 source.t1 a_n2874_n3888# 0.310605f
C262 source.t5 a_n2874_n3888# 0.310605f
C263 source.n31 a_n2874_n3888# 2.7284f
C264 source.n32 a_n2874_n3888# 0.378942f
C265 source.t43 a_n2874_n3888# 0.310605f
C266 source.t6 a_n2874_n3888# 0.310605f
C267 source.n33 a_n2874_n3888# 2.7284f
C268 source.n34 a_n2874_n3888# 0.378942f
C269 source.t42 a_n2874_n3888# 3.48083f
C270 source.n35 a_n2874_n3888# 0.452873f
C271 source.t29 a_n2874_n3888# 3.48083f
C272 source.n36 a_n2874_n3888# 0.452873f
C273 source.t31 a_n2874_n3888# 0.310605f
C274 source.t34 a_n2874_n3888# 0.310605f
C275 source.n37 a_n2874_n3888# 2.7284f
C276 source.n38 a_n2874_n3888# 0.378942f
C277 source.t19 a_n2874_n3888# 0.310605f
C278 source.t27 a_n2874_n3888# 0.310605f
C279 source.n39 a_n2874_n3888# 2.7284f
C280 source.n40 a_n2874_n3888# 0.378942f
C281 source.t30 a_n2874_n3888# 0.310605f
C282 source.t25 a_n2874_n3888# 0.310605f
C283 source.n41 a_n2874_n3888# 2.7284f
C284 source.n42 a_n2874_n3888# 0.378942f
C285 source.t18 a_n2874_n3888# 0.310605f
C286 source.t20 a_n2874_n3888# 0.310605f
C287 source.n43 a_n2874_n3888# 2.7284f
C288 source.n44 a_n2874_n3888# 0.378942f
C289 source.t33 a_n2874_n3888# 0.310605f
C290 source.t15 a_n2874_n3888# 0.310605f
C291 source.n45 a_n2874_n3888# 2.7284f
C292 source.n46 a_n2874_n3888# 0.378942f
C293 source.t12 a_n2874_n3888# 3.48083f
C294 source.n47 a_n2874_n3888# 0.612362f
C295 source.n48 a_n2874_n3888# 1.92461f
C296 minus.n0 a_n2874_n3888# 0.043418f
C297 minus.t3 a_n2874_n3888# 0.925362f
C298 minus.n1 a_n2874_n3888# 0.364637f
C299 minus.t14 a_n2874_n3888# 0.925362f
C300 minus.n2 a_n2874_n3888# 0.043418f
C301 minus.t11 a_n2874_n3888# 0.925362f
C302 minus.n3 a_n2874_n3888# 0.360622f
C303 minus.n4 a_n2874_n3888# 0.043418f
C304 minus.t5 a_n2874_n3888# 0.925362f
C305 minus.n5 a_n2874_n3888# 0.360622f
C306 minus.t10 a_n2874_n3888# 0.925362f
C307 minus.n6 a_n2874_n3888# 0.043418f
C308 minus.t8 a_n2874_n3888# 0.925362f
C309 minus.n7 a_n2874_n3888# 0.364637f
C310 minus.t13 a_n2874_n3888# 0.936837f
C311 minus.t1 a_n2874_n3888# 0.925362f
C312 minus.n8 a_n2874_n3888# 0.369775f
C313 minus.n9 a_n2874_n3888# 0.350436f
C314 minus.n10 a_n2874_n3888# 0.176296f
C315 minus.n11 a_n2874_n3888# 0.043418f
C316 minus.n12 a_n2874_n3888# 0.009852f
C317 minus.t19 a_n2874_n3888# 0.925362f
C318 minus.n13 a_n2874_n3888# 0.365039f
C319 minus.n14 a_n2874_n3888# 0.009852f
C320 minus.n15 a_n2874_n3888# 0.043418f
C321 minus.n16 a_n2874_n3888# 0.043418f
C322 minus.n17 a_n2874_n3888# 0.043418f
C323 minus.n18 a_n2874_n3888# 0.364905f
C324 minus.n19 a_n2874_n3888# 0.009852f
C325 minus.t0 a_n2874_n3888# 0.925362f
C326 minus.n20 a_n2874_n3888# 0.364905f
C327 minus.n21 a_n2874_n3888# 0.043418f
C328 minus.n22 a_n2874_n3888# 0.043418f
C329 minus.n23 a_n2874_n3888# 0.043418f
C330 minus.n24 a_n2874_n3888# 0.009852f
C331 minus.t18 a_n2874_n3888# 0.925362f
C332 minus.n25 a_n2874_n3888# 0.365039f
C333 minus.n26 a_n2874_n3888# 0.009852f
C334 minus.n27 a_n2874_n3888# 0.043418f
C335 minus.n28 a_n2874_n3888# 0.043418f
C336 minus.n29 a_n2874_n3888# 0.043418f
C337 minus.n30 a_n2874_n3888# 0.36089f
C338 minus.n31 a_n2874_n3888# 0.009852f
C339 minus.t22 a_n2874_n3888# 0.925362f
C340 minus.n32 a_n2874_n3888# 0.360087f
C341 minus.n33 a_n2874_n3888# 1.94434f
C342 minus.n34 a_n2874_n3888# 0.043418f
C343 minus.t23 a_n2874_n3888# 0.925362f
C344 minus.n35 a_n2874_n3888# 0.364637f
C345 minus.n36 a_n2874_n3888# 0.043418f
C346 minus.t12 a_n2874_n3888# 0.925362f
C347 minus.n37 a_n2874_n3888# 0.360622f
C348 minus.n38 a_n2874_n3888# 0.043418f
C349 minus.t9 a_n2874_n3888# 0.925362f
C350 minus.n39 a_n2874_n3888# 0.360622f
C351 minus.n40 a_n2874_n3888# 0.043418f
C352 minus.t17 a_n2874_n3888# 0.925362f
C353 minus.n41 a_n2874_n3888# 0.364637f
C354 minus.t7 a_n2874_n3888# 0.936837f
C355 minus.t6 a_n2874_n3888# 0.925362f
C356 minus.n42 a_n2874_n3888# 0.369775f
C357 minus.n43 a_n2874_n3888# 0.350436f
C358 minus.n44 a_n2874_n3888# 0.176296f
C359 minus.n45 a_n2874_n3888# 0.043418f
C360 minus.n46 a_n2874_n3888# 0.009852f
C361 minus.t16 a_n2874_n3888# 0.925362f
C362 minus.n47 a_n2874_n3888# 0.365039f
C363 minus.n48 a_n2874_n3888# 0.009852f
C364 minus.n49 a_n2874_n3888# 0.043418f
C365 minus.n50 a_n2874_n3888# 0.043418f
C366 minus.n51 a_n2874_n3888# 0.043418f
C367 minus.t21 a_n2874_n3888# 0.925362f
C368 minus.n52 a_n2874_n3888# 0.364905f
C369 minus.n53 a_n2874_n3888# 0.009852f
C370 minus.t20 a_n2874_n3888# 0.925362f
C371 minus.n54 a_n2874_n3888# 0.364905f
C372 minus.n55 a_n2874_n3888# 0.043418f
C373 minus.n56 a_n2874_n3888# 0.043418f
C374 minus.n57 a_n2874_n3888# 0.043418f
C375 minus.n58 a_n2874_n3888# 0.009852f
C376 minus.t2 a_n2874_n3888# 0.925362f
C377 minus.n59 a_n2874_n3888# 0.365039f
C378 minus.n60 a_n2874_n3888# 0.009852f
C379 minus.n61 a_n2874_n3888# 0.043418f
C380 minus.n62 a_n2874_n3888# 0.043418f
C381 minus.n63 a_n2874_n3888# 0.043418f
C382 minus.t15 a_n2874_n3888# 0.925362f
C383 minus.n64 a_n2874_n3888# 0.36089f
C384 minus.n65 a_n2874_n3888# 0.009852f
C385 minus.t4 a_n2874_n3888# 0.925362f
C386 minus.n66 a_n2874_n3888# 0.360087f
C387 minus.n67 a_n2874_n3888# 0.286617f
C388 minus.n68 a_n2874_n3888# 2.31917f
.ends

