* NGSPICE file created from diffpair131.ext - technology: sky130A

.subckt diffpair131 minus drain_right drain_left source plus
X0 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X2 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X3 source.t5 minus.t0 drain_right.t0 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X4 source.t0 plus.t0 drain_left.t3 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t4 minus.t1 drain_right.t3 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right.t2 minus.t2 source.t3 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X7 drain_left.t2 plus.t1 source.t1 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X8 source.t6 plus.t2 drain_left.t1 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X9 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X10 drain_right.t1 minus.t3 source.t2 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X11 drain_left.t0 plus.t3 source.t7 a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
R0 minus.n0 minus.t2 166.787
R1 minus.n1 minus.t0 166.787
R2 minus.n0 minus.t1 166.762
R3 minus.n1 minus.t3 166.762
R4 minus.n2 minus.n0 96.7253
R5 minus.n2 minus.n1 76.854
R6 minus minus.n2 0.188
R7 drain_right drain_right.n0 121.636
R8 drain_right drain_right.n1 107.251
R9 drain_right.n0 drain_right.t0 9.9005
R10 drain_right.n0 drain_right.t1 9.9005
R11 drain_right.n1 drain_right.t3 9.9005
R12 drain_right.n1 drain_right.t2 9.9005
R13 source.n58 source.n56 289.615
R14 source.n50 source.n48 289.615
R15 source.n42 source.n40 289.615
R16 source.n34 source.n32 289.615
R17 source.n2 source.n0 289.615
R18 source.n10 source.n8 289.615
R19 source.n18 source.n16 289.615
R20 source.n26 source.n24 289.615
R21 source.n59 source.n58 185
R22 source.n51 source.n50 185
R23 source.n43 source.n42 185
R24 source.n35 source.n34 185
R25 source.n3 source.n2 185
R26 source.n11 source.n10 185
R27 source.n19 source.n18 185
R28 source.n27 source.n26 185
R29 source.t2 source.n57 167.117
R30 source.t5 source.n49 167.117
R31 source.t7 source.n41 167.117
R32 source.t0 source.n33 167.117
R33 source.t1 source.n1 167.117
R34 source.t6 source.n9 167.117
R35 source.t3 source.n17 167.117
R36 source.t4 source.n25 167.117
R37 source.n58 source.t2 52.3082
R38 source.n50 source.t5 52.3082
R39 source.n42 source.t7 52.3082
R40 source.n34 source.t0 52.3082
R41 source.n2 source.t1 52.3082
R42 source.n10 source.t6 52.3082
R43 source.n18 source.t3 52.3082
R44 source.n26 source.t4 52.3082
R45 source.n63 source.n62 31.4096
R46 source.n55 source.n54 31.4096
R47 source.n47 source.n46 31.4096
R48 source.n39 source.n38 31.4096
R49 source.n7 source.n6 31.4096
R50 source.n15 source.n14 31.4096
R51 source.n23 source.n22 31.4096
R52 source.n31 source.n30 31.4096
R53 source.n39 source.n31 14.5137
R54 source.n59 source.n57 9.71174
R55 source.n51 source.n49 9.71174
R56 source.n43 source.n41 9.71174
R57 source.n35 source.n33 9.71174
R58 source.n3 source.n1 9.71174
R59 source.n11 source.n9 9.71174
R60 source.n19 source.n17 9.71174
R61 source.n27 source.n25 9.71174
R62 source.n62 source.n61 9.45567
R63 source.n54 source.n53 9.45567
R64 source.n46 source.n45 9.45567
R65 source.n38 source.n37 9.45567
R66 source.n6 source.n5 9.45567
R67 source.n14 source.n13 9.45567
R68 source.n22 source.n21 9.45567
R69 source.n30 source.n29 9.45567
R70 source.n61 source.n60 9.3005
R71 source.n53 source.n52 9.3005
R72 source.n45 source.n44 9.3005
R73 source.n37 source.n36 9.3005
R74 source.n5 source.n4 9.3005
R75 source.n13 source.n12 9.3005
R76 source.n21 source.n20 9.3005
R77 source.n29 source.n28 9.3005
R78 source.n64 source.n7 8.8499
R79 source.n62 source.n56 8.14595
R80 source.n54 source.n48 8.14595
R81 source.n46 source.n40 8.14595
R82 source.n38 source.n32 8.14595
R83 source.n6 source.n0 8.14595
R84 source.n14 source.n8 8.14595
R85 source.n22 source.n16 8.14595
R86 source.n30 source.n24 8.14595
R87 source.n60 source.n59 7.3702
R88 source.n52 source.n51 7.3702
R89 source.n44 source.n43 7.3702
R90 source.n36 source.n35 7.3702
R91 source.n4 source.n3 7.3702
R92 source.n12 source.n11 7.3702
R93 source.n20 source.n19 7.3702
R94 source.n28 source.n27 7.3702
R95 source.n60 source.n56 5.81868
R96 source.n52 source.n48 5.81868
R97 source.n44 source.n40 5.81868
R98 source.n36 source.n32 5.81868
R99 source.n4 source.n0 5.81868
R100 source.n12 source.n8 5.81868
R101 source.n20 source.n16 5.81868
R102 source.n28 source.n24 5.81868
R103 source.n64 source.n63 5.66429
R104 source.n61 source.n57 3.44771
R105 source.n53 source.n49 3.44771
R106 source.n45 source.n41 3.44771
R107 source.n37 source.n33 3.44771
R108 source.n5 source.n1 3.44771
R109 source.n13 source.n9 3.44771
R110 source.n21 source.n17 3.44771
R111 source.n29 source.n25 3.44771
R112 source.n31 source.n23 0.802224
R113 source.n15 source.n7 0.802224
R114 source.n47 source.n39 0.802224
R115 source.n63 source.n55 0.802224
R116 source.n23 source.n15 0.470328
R117 source.n55 source.n47 0.470328
R118 source source.n64 0.188
R119 plus.n0 plus.t2 166.787
R120 plus.n1 plus.t3 166.787
R121 plus.n0 plus.t1 166.762
R122 plus.n1 plus.t0 166.762
R123 plus plus.n1 94.3942
R124 plus plus.n0 78.7101
R125 drain_left drain_left.n0 122.189
R126 drain_left drain_left.n1 107.251
R127 drain_left.n0 drain_left.t3 9.9005
R128 drain_left.n0 drain_left.t0 9.9005
R129 drain_left.n1 drain_left.t1 9.9005
R130 drain_left.n1 drain_left.t2 9.9005
C0 minus plus 2.88265f
C1 drain_right plus 0.27946f
C2 drain_left source 2.44363f
C3 drain_right minus 0.730102f
C4 drain_left plus 0.849783f
C5 source plus 0.833091f
C6 minus drain_left 0.176251f
C7 drain_right drain_left 0.54499f
C8 minus source 0.819128f
C9 drain_right source 2.44399f
C10 drain_right a_n1274_n1288# 3.54054f
C11 drain_left a_n1274_n1288# 3.67836f
C12 source a_n1274_n1288# 2.88579f
C13 minus a_n1274_n1288# 3.988958f
C14 plus a_n1274_n1288# 5.56009f
C15 drain_left.t3 a_n1274_n1288# 0.030903f
C16 drain_left.t0 a_n1274_n1288# 0.030903f
C17 drain_left.n0 a_n1274_n1288# 0.279462f
C18 drain_left.t1 a_n1274_n1288# 0.030903f
C19 drain_left.t2 a_n1274_n1288# 0.030903f
C20 drain_left.n1 a_n1274_n1288# 0.219963f
C21 plus.t1 a_n1274_n1288# 0.145918f
C22 plus.t2 a_n1274_n1288# 0.145938f
C23 plus.n0 a_n1274_n1288# 0.200292f
C24 plus.t0 a_n1274_n1288# 0.145918f
C25 plus.t3 a_n1274_n1288# 0.145938f
C26 plus.n1 a_n1274_n1288# 0.365341f
C27 source.n0 a_n1274_n1288# 0.024659f
C28 source.n1 a_n1274_n1288# 0.05456f
C29 source.t1 a_n1274_n1288# 0.040945f
C30 source.n2 a_n1274_n1288# 0.042701f
C31 source.n3 a_n1274_n1288# 0.013765f
C32 source.n4 a_n1274_n1288# 0.009078f
C33 source.n5 a_n1274_n1288# 0.120264f
C34 source.n6 a_n1274_n1288# 0.027032f
C35 source.n7 a_n1274_n1288# 0.280044f
C36 source.n8 a_n1274_n1288# 0.024659f
C37 source.n9 a_n1274_n1288# 0.05456f
C38 source.t6 a_n1274_n1288# 0.040945f
C39 source.n10 a_n1274_n1288# 0.042701f
C40 source.n11 a_n1274_n1288# 0.013765f
C41 source.n12 a_n1274_n1288# 0.009078f
C42 source.n13 a_n1274_n1288# 0.120264f
C43 source.n14 a_n1274_n1288# 0.027032f
C44 source.n15 a_n1274_n1288# 0.083129f
C45 source.n16 a_n1274_n1288# 0.024659f
C46 source.n17 a_n1274_n1288# 0.05456f
C47 source.t3 a_n1274_n1288# 0.040945f
C48 source.n18 a_n1274_n1288# 0.042701f
C49 source.n19 a_n1274_n1288# 0.013765f
C50 source.n20 a_n1274_n1288# 0.009078f
C51 source.n21 a_n1274_n1288# 0.120264f
C52 source.n22 a_n1274_n1288# 0.027032f
C53 source.n23 a_n1274_n1288# 0.083129f
C54 source.n24 a_n1274_n1288# 0.024659f
C55 source.n25 a_n1274_n1288# 0.05456f
C56 source.t4 a_n1274_n1288# 0.040945f
C57 source.n26 a_n1274_n1288# 0.042701f
C58 source.n27 a_n1274_n1288# 0.013765f
C59 source.n28 a_n1274_n1288# 0.009078f
C60 source.n29 a_n1274_n1288# 0.120264f
C61 source.n30 a_n1274_n1288# 0.027032f
C62 source.n31 a_n1274_n1288# 0.440747f
C63 source.n32 a_n1274_n1288# 0.024659f
C64 source.n33 a_n1274_n1288# 0.05456f
C65 source.t0 a_n1274_n1288# 0.040945f
C66 source.n34 a_n1274_n1288# 0.042701f
C67 source.n35 a_n1274_n1288# 0.013765f
C68 source.n36 a_n1274_n1288# 0.009078f
C69 source.n37 a_n1274_n1288# 0.120264f
C70 source.n38 a_n1274_n1288# 0.027032f
C71 source.n39 a_n1274_n1288# 0.440747f
C72 source.n40 a_n1274_n1288# 0.024659f
C73 source.n41 a_n1274_n1288# 0.05456f
C74 source.t7 a_n1274_n1288# 0.040945f
C75 source.n42 a_n1274_n1288# 0.042701f
C76 source.n43 a_n1274_n1288# 0.013765f
C77 source.n44 a_n1274_n1288# 0.009078f
C78 source.n45 a_n1274_n1288# 0.120264f
C79 source.n46 a_n1274_n1288# 0.027032f
C80 source.n47 a_n1274_n1288# 0.083129f
C81 source.n48 a_n1274_n1288# 0.024659f
C82 source.n49 a_n1274_n1288# 0.05456f
C83 source.t5 a_n1274_n1288# 0.040945f
C84 source.n50 a_n1274_n1288# 0.042701f
C85 source.n51 a_n1274_n1288# 0.013765f
C86 source.n52 a_n1274_n1288# 0.009078f
C87 source.n53 a_n1274_n1288# 0.120264f
C88 source.n54 a_n1274_n1288# 0.027032f
C89 source.n55 a_n1274_n1288# 0.083129f
C90 source.n56 a_n1274_n1288# 0.024659f
C91 source.n57 a_n1274_n1288# 0.05456f
C92 source.t2 a_n1274_n1288# 0.040945f
C93 source.n58 a_n1274_n1288# 0.042701f
C94 source.n59 a_n1274_n1288# 0.013765f
C95 source.n60 a_n1274_n1288# 0.009078f
C96 source.n61 a_n1274_n1288# 0.120264f
C97 source.n62 a_n1274_n1288# 0.027032f
C98 source.n63 a_n1274_n1288# 0.189656f
C99 source.n64 a_n1274_n1288# 0.423812f
C100 drain_right.t0 a_n1274_n1288# 0.03192f
C101 drain_right.t1 a_n1274_n1288# 0.03192f
C102 drain_right.n0 a_n1274_n1288# 0.279952f
C103 drain_right.t3 a_n1274_n1288# 0.03192f
C104 drain_right.t2 a_n1274_n1288# 0.03192f
C105 drain_right.n1 a_n1274_n1288# 0.227204f
C106 minus.t2 a_n1274_n1288# 0.142358f
C107 minus.t1 a_n1274_n1288# 0.142339f
C108 minus.n0 a_n1274_n1288# 0.377745f
C109 minus.t0 a_n1274_n1288# 0.142358f
C110 minus.t3 a_n1274_n1288# 0.142339f
C111 minus.n1 a_n1274_n1288# 0.186783f
C112 minus.n2 a_n1274_n1288# 1.74298f
.ends

