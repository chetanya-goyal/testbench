* NGSPICE file created from diffpair218.ext - technology: sky130A

.subckt diffpair218 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t36 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X1 drain_right.t19 minus.t0 source.t12 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X2 source.t26 plus.t1 drain_left.t18 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X3 source.t0 minus.t1 drain_right.t18 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X4 source.t20 plus.t2 drain_left.t17 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X5 drain_left.t16 plus.t3 source.t38 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X6 source.t15 minus.t2 drain_right.t17 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X7 source.t37 plus.t4 drain_left.t15 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X8 drain_right.t16 minus.t3 source.t2 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X9 drain_left.t14 plus.t5 source.t39 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X10 source.t9 minus.t4 drain_right.t15 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X11 source.t3 minus.t5 drain_right.t14 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 drain_right.t13 minus.t6 source.t5 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X13 source.t33 plus.t6 drain_left.t13 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X14 drain_right.t12 minus.t7 source.t16 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X15 drain_right.t11 minus.t8 source.t6 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X16 source.t10 minus.t9 drain_right.t10 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X17 a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X18 drain_left.t12 plus.t7 source.t34 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X19 a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X20 drain_left.t11 plus.t8 source.t29 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X21 drain_right.t9 minus.t10 source.t13 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X22 drain_left.t10 plus.t9 source.t35 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X23 source.t21 plus.t10 drain_left.t9 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X24 source.t4 minus.t11 drain_right.t8 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X25 source.t1 minus.t12 drain_right.t7 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X26 drain_right.t6 minus.t13 source.t17 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X27 source.t31 plus.t11 drain_left.t8 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X28 source.t11 minus.t14 drain_right.t5 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X29 drain_left.t7 plus.t12 source.t27 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X30 source.t8 minus.t15 drain_right.t4 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X31 drain_right.t3 minus.t16 source.t18 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X32 drain_right.t2 minus.t17 source.t19 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X33 source.t30 plus.t13 drain_left.t6 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X34 a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X35 source.t32 plus.t14 drain_left.t5 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X36 drain_right.t1 minus.t18 source.t7 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X37 source.t14 minus.t19 drain_right.t0 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X38 drain_left.t4 plus.t15 source.t23 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X39 source.t28 plus.t16 drain_left.t3 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X40 drain_left.t2 plus.t17 source.t24 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X41 a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X42 drain_left.t1 plus.t18 source.t25 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X43 source.t22 plus.t19 drain_left.t0 a_n2762_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 plus.n8 plus.t16 212.793
R1 plus.n36 plus.t7 212.793
R2 plus.n26 plus.t0 185.972
R3 plus.n25 plus.t2 185.972
R4 plus.n24 plus.t3 185.972
R5 plus.n2 plus.t4 185.972
R6 plus.n18 plus.t5 185.972
R7 plus.n4 plus.t10 185.972
R8 plus.n12 plus.t12 185.972
R9 plus.n6 plus.t14 185.972
R10 plus.n7 plus.t15 185.972
R11 plus.n54 plus.t1 185.972
R12 plus.n53 plus.t9 185.972
R13 plus.n52 plus.t13 185.972
R14 plus.n30 plus.t18 185.972
R15 plus.n46 plus.t6 185.972
R16 plus.n32 plus.t8 185.972
R17 plus.n40 plus.t11 185.972
R18 plus.n34 plus.t17 185.972
R19 plus.n35 plus.t19 185.972
R20 plus.n9 plus.n6 161.3
R21 plus.n11 plus.n10 161.3
R22 plus.n12 plus.n5 161.3
R23 plus.n14 plus.n13 161.3
R24 plus.n15 plus.n4 161.3
R25 plus.n17 plus.n16 161.3
R26 plus.n18 plus.n3 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n2 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n24 plus.n1 161.3
R31 plus.n27 plus.n26 161.3
R32 plus.n37 plus.n34 161.3
R33 plus.n39 plus.n38 161.3
R34 plus.n40 plus.n33 161.3
R35 plus.n42 plus.n41 161.3
R36 plus.n43 plus.n32 161.3
R37 plus.n45 plus.n44 161.3
R38 plus.n46 plus.n31 161.3
R39 plus.n48 plus.n47 161.3
R40 plus.n49 plus.n30 161.3
R41 plus.n51 plus.n50 161.3
R42 plus.n52 plus.n29 161.3
R43 plus.n55 plus.n54 161.3
R44 plus.n25 plus.n0 80.6037
R45 plus.n53 plus.n28 80.6037
R46 plus.n26 plus.n25 48.2005
R47 plus.n25 plus.n24 48.2005
R48 plus.n7 plus.n6 48.2005
R49 plus.n54 plus.n53 48.2005
R50 plus.n53 plus.n52 48.2005
R51 plus.n35 plus.n34 48.2005
R52 plus.n9 plus.n8 45.1367
R53 plus.n37 plus.n36 45.1367
R54 plus.n23 plus.n2 44.549
R55 plus.n12 plus.n11 44.549
R56 plus.n51 plus.n30 44.549
R57 plus.n40 plus.n39 44.549
R58 plus.n19 plus.n18 34.3247
R59 plus.n13 plus.n4 34.3247
R60 plus.n47 plus.n46 34.3247
R61 plus.n41 plus.n32 34.3247
R62 plus plus.n55 30.1846
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n19 plus.n2 13.8763
R68 plus.n13 plus.n12 13.8763
R69 plus.n47 plus.n30 13.8763
R70 plus.n41 plus.n40 13.8763
R71 plus.n8 plus.n7 13.3799
R72 plus.n36 plus.n35 13.3799
R73 plus plus.n27 8.86414
R74 plus.n24 plus.n23 3.65202
R75 plus.n11 plus.n6 3.65202
R76 plus.n52 plus.n51 3.65202
R77 plus.n39 plus.n34 3.65202
R78 plus.n1 plus.n0 0.285035
R79 plus.n27 plus.n0 0.285035
R80 plus.n55 plus.n28 0.285035
R81 plus.n29 plus.n28 0.285035
R82 plus.n10 plus.n9 0.189894
R83 plus.n10 plus.n5 0.189894
R84 plus.n14 plus.n5 0.189894
R85 plus.n15 plus.n14 0.189894
R86 plus.n16 plus.n15 0.189894
R87 plus.n16 plus.n3 0.189894
R88 plus.n20 plus.n3 0.189894
R89 plus.n21 plus.n20 0.189894
R90 plus.n22 plus.n21 0.189894
R91 plus.n22 plus.n1 0.189894
R92 plus.n50 plus.n29 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n48 0.189894
R95 plus.n48 plus.n31 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n38 plus.n33 0.189894
R101 plus.n38 plus.n37 0.189894
R102 source.n0 source.t36 69.6943
R103 source.n9 source.t28 69.6943
R104 source.n10 source.t7 69.6943
R105 source.n19 source.t15 69.6943
R106 source.n39 source.t13 69.6942
R107 source.n30 source.t14 69.6942
R108 source.n29 source.t34 69.6942
R109 source.n20 source.t26 69.6942
R110 source.n2 source.n1 63.0943
R111 source.n4 source.n3 63.0943
R112 source.n6 source.n5 63.0943
R113 source.n8 source.n7 63.0943
R114 source.n12 source.n11 63.0943
R115 source.n14 source.n13 63.0943
R116 source.n16 source.n15 63.0943
R117 source.n18 source.n17 63.0943
R118 source.n38 source.n37 63.0942
R119 source.n36 source.n35 63.0942
R120 source.n34 source.n33 63.0942
R121 source.n32 source.n31 63.0942
R122 source.n28 source.n27 63.0942
R123 source.n26 source.n25 63.0942
R124 source.n24 source.n23 63.0942
R125 source.n22 source.n21 63.0942
R126 source.n20 source.n19 15.2713
R127 source.n40 source.n0 9.60747
R128 source.n37 source.t12 6.6005
R129 source.n37 source.t11 6.6005
R130 source.n35 source.t18 6.6005
R131 source.n35 source.t3 6.6005
R132 source.n33 source.t19 6.6005
R133 source.n33 source.t1 6.6005
R134 source.n31 source.t5 6.6005
R135 source.n31 source.t0 6.6005
R136 source.n27 source.t24 6.6005
R137 source.n27 source.t22 6.6005
R138 source.n25 source.t29 6.6005
R139 source.n25 source.t31 6.6005
R140 source.n23 source.t25 6.6005
R141 source.n23 source.t33 6.6005
R142 source.n21 source.t35 6.6005
R143 source.n21 source.t30 6.6005
R144 source.n1 source.t38 6.6005
R145 source.n1 source.t20 6.6005
R146 source.n3 source.t39 6.6005
R147 source.n3 source.t37 6.6005
R148 source.n5 source.t27 6.6005
R149 source.n5 source.t21 6.6005
R150 source.n7 source.t23 6.6005
R151 source.n7 source.t32 6.6005
R152 source.n11 source.t17 6.6005
R153 source.n11 source.t8 6.6005
R154 source.n13 source.t16 6.6005
R155 source.n13 source.t4 6.6005
R156 source.n15 source.t6 6.6005
R157 source.n15 source.t10 6.6005
R158 source.n17 source.t2 6.6005
R159 source.n17 source.t9 6.6005
R160 source.n40 source.n39 5.66429
R161 source.n19 source.n18 0.802224
R162 source.n18 source.n16 0.802224
R163 source.n16 source.n14 0.802224
R164 source.n14 source.n12 0.802224
R165 source.n12 source.n10 0.802224
R166 source.n9 source.n8 0.802224
R167 source.n8 source.n6 0.802224
R168 source.n6 source.n4 0.802224
R169 source.n4 source.n2 0.802224
R170 source.n2 source.n0 0.802224
R171 source.n22 source.n20 0.802224
R172 source.n24 source.n22 0.802224
R173 source.n26 source.n24 0.802224
R174 source.n28 source.n26 0.802224
R175 source.n29 source.n28 0.802224
R176 source.n32 source.n30 0.802224
R177 source.n34 source.n32 0.802224
R178 source.n36 source.n34 0.802224
R179 source.n38 source.n36 0.802224
R180 source.n39 source.n38 0.802224
R181 source.n10 source.n9 0.470328
R182 source.n30 source.n29 0.470328
R183 source source.n40 0.188
R184 drain_left.n10 drain_left.n8 80.5748
R185 drain_left.n6 drain_left.n4 80.5747
R186 drain_left.n2 drain_left.n0 80.5747
R187 drain_left.n16 drain_left.n15 79.7731
R188 drain_left.n14 drain_left.n13 79.7731
R189 drain_left.n12 drain_left.n11 79.7731
R190 drain_left.n10 drain_left.n9 79.7731
R191 drain_left.n7 drain_left.n3 79.773
R192 drain_left.n6 drain_left.n5 79.773
R193 drain_left.n2 drain_left.n1 79.773
R194 drain_left drain_left.n7 26.9627
R195 drain_left.n3 drain_left.t13 6.6005
R196 drain_left.n3 drain_left.t11 6.6005
R197 drain_left.n4 drain_left.t0 6.6005
R198 drain_left.n4 drain_left.t12 6.6005
R199 drain_left.n5 drain_left.t8 6.6005
R200 drain_left.n5 drain_left.t2 6.6005
R201 drain_left.n1 drain_left.t6 6.6005
R202 drain_left.n1 drain_left.t1 6.6005
R203 drain_left.n0 drain_left.t18 6.6005
R204 drain_left.n0 drain_left.t10 6.6005
R205 drain_left.n15 drain_left.t17 6.6005
R206 drain_left.n15 drain_left.t19 6.6005
R207 drain_left.n13 drain_left.t15 6.6005
R208 drain_left.n13 drain_left.t16 6.6005
R209 drain_left.n11 drain_left.t9 6.6005
R210 drain_left.n11 drain_left.t14 6.6005
R211 drain_left.n9 drain_left.t5 6.6005
R212 drain_left.n9 drain_left.t7 6.6005
R213 drain_left.n8 drain_left.t3 6.6005
R214 drain_left.n8 drain_left.t4 6.6005
R215 drain_left drain_left.n16 6.45494
R216 drain_left.n12 drain_left.n10 0.802224
R217 drain_left.n14 drain_left.n12 0.802224
R218 drain_left.n16 drain_left.n14 0.802224
R219 drain_left.n7 drain_left.n6 0.746878
R220 drain_left.n7 drain_left.n2 0.746878
R221 minus.n6 minus.t18 212.793
R222 minus.n34 minus.t19 212.793
R223 minus.n7 minus.t15 185.972
R224 minus.n8 minus.t13 185.972
R225 minus.n12 minus.t11 185.972
R226 minus.n14 minus.t7 185.972
R227 minus.n18 minus.t9 185.972
R228 minus.n20 minus.t8 185.972
R229 minus.n24 minus.t4 185.972
R230 minus.n25 minus.t3 185.972
R231 minus.n26 minus.t2 185.972
R232 minus.n35 minus.t6 185.972
R233 minus.n36 minus.t1 185.972
R234 minus.n40 minus.t17 185.972
R235 minus.n42 minus.t12 185.972
R236 minus.n46 minus.t16 185.972
R237 minus.n48 minus.t5 185.972
R238 minus.n52 minus.t0 185.972
R239 minus.n53 minus.t14 185.972
R240 minus.n54 minus.t10 185.972
R241 minus.n27 minus.n26 161.3
R242 minus.n24 minus.n23 161.3
R243 minus.n22 minus.n1 161.3
R244 minus.n21 minus.n20 161.3
R245 minus.n19 minus.n2 161.3
R246 minus.n18 minus.n17 161.3
R247 minus.n16 minus.n3 161.3
R248 minus.n15 minus.n14 161.3
R249 minus.n13 minus.n4 161.3
R250 minus.n12 minus.n11 161.3
R251 minus.n10 minus.n5 161.3
R252 minus.n9 minus.n8 161.3
R253 minus.n55 minus.n54 161.3
R254 minus.n52 minus.n51 161.3
R255 minus.n50 minus.n29 161.3
R256 minus.n49 minus.n48 161.3
R257 minus.n47 minus.n30 161.3
R258 minus.n46 minus.n45 161.3
R259 minus.n44 minus.n31 161.3
R260 minus.n43 minus.n42 161.3
R261 minus.n41 minus.n32 161.3
R262 minus.n40 minus.n39 161.3
R263 minus.n38 minus.n33 161.3
R264 minus.n37 minus.n36 161.3
R265 minus.n25 minus.n0 80.6037
R266 minus.n53 minus.n28 80.6037
R267 minus.n8 minus.n7 48.2005
R268 minus.n25 minus.n24 48.2005
R269 minus.n26 minus.n25 48.2005
R270 minus.n36 minus.n35 48.2005
R271 minus.n53 minus.n52 48.2005
R272 minus.n54 minus.n53 48.2005
R273 minus.n9 minus.n6 45.1367
R274 minus.n37 minus.n34 45.1367
R275 minus.n12 minus.n5 44.549
R276 minus.n20 minus.n1 44.549
R277 minus.n40 minus.n33 44.549
R278 minus.n48 minus.n29 44.549
R279 minus.n14 minus.n13 34.3247
R280 minus.n19 minus.n18 34.3247
R281 minus.n42 minus.n41 34.3247
R282 minus.n47 minus.n46 34.3247
R283 minus.n56 minus.n27 32.8944
R284 minus.n18 minus.n3 24.1005
R285 minus.n14 minus.n3 24.1005
R286 minus.n42 minus.n31 24.1005
R287 minus.n46 minus.n31 24.1005
R288 minus.n13 minus.n12 13.8763
R289 minus.n20 minus.n19 13.8763
R290 minus.n41 minus.n40 13.8763
R291 minus.n48 minus.n47 13.8763
R292 minus.n7 minus.n6 13.3799
R293 minus.n35 minus.n34 13.3799
R294 minus.n56 minus.n55 6.62929
R295 minus.n8 minus.n5 3.65202
R296 minus.n24 minus.n1 3.65202
R297 minus.n36 minus.n33 3.65202
R298 minus.n52 minus.n29 3.65202
R299 minus.n27 minus.n0 0.285035
R300 minus.n23 minus.n0 0.285035
R301 minus.n51 minus.n28 0.285035
R302 minus.n55 minus.n28 0.285035
R303 minus.n23 minus.n22 0.189894
R304 minus.n22 minus.n21 0.189894
R305 minus.n21 minus.n2 0.189894
R306 minus.n17 minus.n2 0.189894
R307 minus.n17 minus.n16 0.189894
R308 minus.n16 minus.n15 0.189894
R309 minus.n15 minus.n4 0.189894
R310 minus.n11 minus.n4 0.189894
R311 minus.n11 minus.n10 0.189894
R312 minus.n10 minus.n9 0.189894
R313 minus.n38 minus.n37 0.189894
R314 minus.n39 minus.n38 0.189894
R315 minus.n39 minus.n32 0.189894
R316 minus.n43 minus.n32 0.189894
R317 minus.n44 minus.n43 0.189894
R318 minus.n45 minus.n44 0.189894
R319 minus.n45 minus.n30 0.189894
R320 minus.n49 minus.n30 0.189894
R321 minus.n50 minus.n49 0.189894
R322 minus.n51 minus.n50 0.189894
R323 minus minus.n56 0.188
R324 drain_right.n10 drain_right.n8 80.5748
R325 drain_right.n6 drain_right.n4 80.5747
R326 drain_right.n2 drain_right.n0 80.5747
R327 drain_right.n10 drain_right.n9 79.7731
R328 drain_right.n12 drain_right.n11 79.7731
R329 drain_right.n14 drain_right.n13 79.7731
R330 drain_right.n16 drain_right.n15 79.7731
R331 drain_right.n7 drain_right.n3 79.773
R332 drain_right.n6 drain_right.n5 79.773
R333 drain_right.n2 drain_right.n1 79.773
R334 drain_right drain_right.n7 26.4095
R335 drain_right.n3 drain_right.t7 6.6005
R336 drain_right.n3 drain_right.t3 6.6005
R337 drain_right.n4 drain_right.t5 6.6005
R338 drain_right.n4 drain_right.t9 6.6005
R339 drain_right.n5 drain_right.t14 6.6005
R340 drain_right.n5 drain_right.t19 6.6005
R341 drain_right.n1 drain_right.t18 6.6005
R342 drain_right.n1 drain_right.t2 6.6005
R343 drain_right.n0 drain_right.t0 6.6005
R344 drain_right.n0 drain_right.t13 6.6005
R345 drain_right.n8 drain_right.t4 6.6005
R346 drain_right.n8 drain_right.t1 6.6005
R347 drain_right.n9 drain_right.t8 6.6005
R348 drain_right.n9 drain_right.t6 6.6005
R349 drain_right.n11 drain_right.t10 6.6005
R350 drain_right.n11 drain_right.t12 6.6005
R351 drain_right.n13 drain_right.t15 6.6005
R352 drain_right.n13 drain_right.t11 6.6005
R353 drain_right.n15 drain_right.t17 6.6005
R354 drain_right.n15 drain_right.t16 6.6005
R355 drain_right drain_right.n16 6.45494
R356 drain_right.n16 drain_right.n14 0.802224
R357 drain_right.n14 drain_right.n12 0.802224
R358 drain_right.n12 drain_right.n10 0.802224
R359 drain_right.n7 drain_right.n6 0.746878
R360 drain_right.n7 drain_right.n2 0.746878
C0 plus drain_left 3.64665f
C1 plus source 3.94161f
C2 source drain_left 9.438349f
C3 drain_right minus 3.37209f
C4 drain_right plus 0.437356f
C5 drain_right drain_left 1.48678f
C6 drain_right source 9.44019f
C7 plus minus 4.9329f
C8 minus drain_left 0.178626f
C9 minus source 3.92761f
C10 drain_right a_n2762_n1488# 5.37519f
C11 drain_left a_n2762_n1488# 5.76983f
C12 source a_n2762_n1488# 4.038527f
C13 minus a_n2762_n1488# 10.301899f
C14 plus a_n2762_n1488# 11.70051f
C15 drain_right.t0 a_n2762_n1488# 0.0654f
C16 drain_right.t13 a_n2762_n1488# 0.0654f
C17 drain_right.n0 a_n2762_n1488# 0.475384f
C18 drain_right.t18 a_n2762_n1488# 0.0654f
C19 drain_right.t2 a_n2762_n1488# 0.0654f
C20 drain_right.n1 a_n2762_n1488# 0.471658f
C21 drain_right.n2 a_n2762_n1488# 0.730044f
C22 drain_right.t7 a_n2762_n1488# 0.0654f
C23 drain_right.t3 a_n2762_n1488# 0.0654f
C24 drain_right.n3 a_n2762_n1488# 0.471658f
C25 drain_right.t5 a_n2762_n1488# 0.0654f
C26 drain_right.t9 a_n2762_n1488# 0.0654f
C27 drain_right.n4 a_n2762_n1488# 0.475384f
C28 drain_right.t14 a_n2762_n1488# 0.0654f
C29 drain_right.t19 a_n2762_n1488# 0.0654f
C30 drain_right.n5 a_n2762_n1488# 0.471658f
C31 drain_right.n6 a_n2762_n1488# 0.730044f
C32 drain_right.n7 a_n2762_n1488# 1.34703f
C33 drain_right.t4 a_n2762_n1488# 0.0654f
C34 drain_right.t1 a_n2762_n1488# 0.0654f
C35 drain_right.n8 a_n2762_n1488# 0.475386f
C36 drain_right.t8 a_n2762_n1488# 0.0654f
C37 drain_right.t6 a_n2762_n1488# 0.0654f
C38 drain_right.n9 a_n2762_n1488# 0.47166f
C39 drain_right.n10 a_n2762_n1488# 0.734103f
C40 drain_right.t10 a_n2762_n1488# 0.0654f
C41 drain_right.t12 a_n2762_n1488# 0.0654f
C42 drain_right.n11 a_n2762_n1488# 0.47166f
C43 drain_right.n12 a_n2762_n1488# 0.363359f
C44 drain_right.t15 a_n2762_n1488# 0.0654f
C45 drain_right.t11 a_n2762_n1488# 0.0654f
C46 drain_right.n13 a_n2762_n1488# 0.47166f
C47 drain_right.n14 a_n2762_n1488# 0.363359f
C48 drain_right.t17 a_n2762_n1488# 0.0654f
C49 drain_right.t16 a_n2762_n1488# 0.0654f
C50 drain_right.n15 a_n2762_n1488# 0.47166f
C51 drain_right.n16 a_n2762_n1488# 0.603914f
C52 minus.n0 a_n2762_n1488# 0.05737f
C53 minus.n1 a_n2762_n1488# 0.009779f
C54 minus.t4 a_n2762_n1488# 0.232605f
C55 minus.n2 a_n2762_n1488# 0.043095f
C56 minus.n3 a_n2762_n1488# 0.009779f
C57 minus.t9 a_n2762_n1488# 0.232605f
C58 minus.n4 a_n2762_n1488# 0.043095f
C59 minus.n5 a_n2762_n1488# 0.009779f
C60 minus.t11 a_n2762_n1488# 0.232605f
C61 minus.t18 a_n2762_n1488# 0.249959f
C62 minus.n6 a_n2762_n1488# 0.121127f
C63 minus.t15 a_n2762_n1488# 0.232605f
C64 minus.n7 a_n2762_n1488# 0.147334f
C65 minus.t13 a_n2762_n1488# 0.232605f
C66 minus.n8 a_n2762_n1488# 0.138219f
C67 minus.n9 a_n2762_n1488# 0.183941f
C68 minus.n10 a_n2762_n1488# 0.043095f
C69 minus.n11 a_n2762_n1488# 0.043095f
C70 minus.n12 a_n2762_n1488# 0.139415f
C71 minus.n13 a_n2762_n1488# 0.009779f
C72 minus.t7 a_n2762_n1488# 0.232605f
C73 minus.n14 a_n2762_n1488# 0.139415f
C74 minus.n15 a_n2762_n1488# 0.043095f
C75 minus.n16 a_n2762_n1488# 0.043095f
C76 minus.n17 a_n2762_n1488# 0.043095f
C77 minus.n18 a_n2762_n1488# 0.139415f
C78 minus.n19 a_n2762_n1488# 0.009779f
C79 minus.t8 a_n2762_n1488# 0.232605f
C80 minus.n20 a_n2762_n1488# 0.139415f
C81 minus.n21 a_n2762_n1488# 0.043095f
C82 minus.n22 a_n2762_n1488# 0.043095f
C83 minus.n23 a_n2762_n1488# 0.057504f
C84 minus.n24 a_n2762_n1488# 0.138219f
C85 minus.t3 a_n2762_n1488# 0.232605f
C86 minus.n25 a_n2762_n1488# 0.147334f
C87 minus.t2 a_n2762_n1488# 0.232605f
C88 minus.n26 a_n2762_n1488# 0.137555f
C89 minus.n27 a_n2762_n1488# 1.32652f
C90 minus.n28 a_n2762_n1488# 0.05737f
C91 minus.n29 a_n2762_n1488# 0.009779f
C92 minus.n30 a_n2762_n1488# 0.043095f
C93 minus.n31 a_n2762_n1488# 0.009779f
C94 minus.n32 a_n2762_n1488# 0.043095f
C95 minus.n33 a_n2762_n1488# 0.009779f
C96 minus.t19 a_n2762_n1488# 0.249959f
C97 minus.n34 a_n2762_n1488# 0.121127f
C98 minus.t6 a_n2762_n1488# 0.232605f
C99 minus.n35 a_n2762_n1488# 0.147334f
C100 minus.t1 a_n2762_n1488# 0.232605f
C101 minus.n36 a_n2762_n1488# 0.138219f
C102 minus.n37 a_n2762_n1488# 0.183941f
C103 minus.n38 a_n2762_n1488# 0.043095f
C104 minus.n39 a_n2762_n1488# 0.043095f
C105 minus.t17 a_n2762_n1488# 0.232605f
C106 minus.n40 a_n2762_n1488# 0.139415f
C107 minus.n41 a_n2762_n1488# 0.009779f
C108 minus.t12 a_n2762_n1488# 0.232605f
C109 minus.n42 a_n2762_n1488# 0.139415f
C110 minus.n43 a_n2762_n1488# 0.043095f
C111 minus.n44 a_n2762_n1488# 0.043095f
C112 minus.n45 a_n2762_n1488# 0.043095f
C113 minus.t16 a_n2762_n1488# 0.232605f
C114 minus.n46 a_n2762_n1488# 0.139415f
C115 minus.n47 a_n2762_n1488# 0.009779f
C116 minus.t5 a_n2762_n1488# 0.232605f
C117 minus.n48 a_n2762_n1488# 0.139415f
C118 minus.n49 a_n2762_n1488# 0.043095f
C119 minus.n50 a_n2762_n1488# 0.043095f
C120 minus.n51 a_n2762_n1488# 0.057504f
C121 minus.t0 a_n2762_n1488# 0.232605f
C122 minus.n52 a_n2762_n1488# 0.138219f
C123 minus.t14 a_n2762_n1488# 0.232605f
C124 minus.n53 a_n2762_n1488# 0.147334f
C125 minus.t10 a_n2762_n1488# 0.232605f
C126 minus.n54 a_n2762_n1488# 0.137555f
C127 minus.n55 a_n2762_n1488# 0.309198f
C128 minus.n56 a_n2762_n1488# 1.60316f
C129 drain_left.t18 a_n2762_n1488# 0.065867f
C130 drain_left.t10 a_n2762_n1488# 0.065867f
C131 drain_left.n0 a_n2762_n1488# 0.478775f
C132 drain_left.t6 a_n2762_n1488# 0.065867f
C133 drain_left.t1 a_n2762_n1488# 0.065867f
C134 drain_left.n1 a_n2762_n1488# 0.475022f
C135 drain_left.n2 a_n2762_n1488# 0.735252f
C136 drain_left.t13 a_n2762_n1488# 0.065867f
C137 drain_left.t11 a_n2762_n1488# 0.065867f
C138 drain_left.n3 a_n2762_n1488# 0.475022f
C139 drain_left.t0 a_n2762_n1488# 0.065867f
C140 drain_left.t12 a_n2762_n1488# 0.065867f
C141 drain_left.n4 a_n2762_n1488# 0.478775f
C142 drain_left.t8 a_n2762_n1488# 0.065867f
C143 drain_left.t2 a_n2762_n1488# 0.065867f
C144 drain_left.n5 a_n2762_n1488# 0.475022f
C145 drain_left.n6 a_n2762_n1488# 0.735252f
C146 drain_left.n7 a_n2762_n1488# 1.4111f
C147 drain_left.t3 a_n2762_n1488# 0.065867f
C148 drain_left.t4 a_n2762_n1488# 0.065867f
C149 drain_left.n8 a_n2762_n1488# 0.478777f
C150 drain_left.t5 a_n2762_n1488# 0.065867f
C151 drain_left.t7 a_n2762_n1488# 0.065867f
C152 drain_left.n9 a_n2762_n1488# 0.475025f
C153 drain_left.n10 a_n2762_n1488# 0.73934f
C154 drain_left.t9 a_n2762_n1488# 0.065867f
C155 drain_left.t14 a_n2762_n1488# 0.065867f
C156 drain_left.n11 a_n2762_n1488# 0.475025f
C157 drain_left.n12 a_n2762_n1488# 0.365951f
C158 drain_left.t15 a_n2762_n1488# 0.065867f
C159 drain_left.t16 a_n2762_n1488# 0.065867f
C160 drain_left.n13 a_n2762_n1488# 0.475025f
C161 drain_left.n14 a_n2762_n1488# 0.365951f
C162 drain_left.t17 a_n2762_n1488# 0.065867f
C163 drain_left.t19 a_n2762_n1488# 0.065867f
C164 drain_left.n15 a_n2762_n1488# 0.475025f
C165 drain_left.n16 a_n2762_n1488# 0.608222f
C166 source.t36 a_n2762_n1488# 0.573812f
C167 source.n0 a_n2762_n1488# 0.825567f
C168 source.t38 a_n2762_n1488# 0.069102f
C169 source.t20 a_n2762_n1488# 0.069102f
C170 source.n1 a_n2762_n1488# 0.438147f
C171 source.n2 a_n2762_n1488# 0.404522f
C172 source.t39 a_n2762_n1488# 0.069102f
C173 source.t37 a_n2762_n1488# 0.069102f
C174 source.n3 a_n2762_n1488# 0.438147f
C175 source.n4 a_n2762_n1488# 0.404522f
C176 source.t27 a_n2762_n1488# 0.069102f
C177 source.t21 a_n2762_n1488# 0.069102f
C178 source.n5 a_n2762_n1488# 0.438147f
C179 source.n6 a_n2762_n1488# 0.404522f
C180 source.t23 a_n2762_n1488# 0.069102f
C181 source.t32 a_n2762_n1488# 0.069102f
C182 source.n7 a_n2762_n1488# 0.438147f
C183 source.n8 a_n2762_n1488# 0.404522f
C184 source.t28 a_n2762_n1488# 0.573812f
C185 source.n9 a_n2762_n1488# 0.426145f
C186 source.t7 a_n2762_n1488# 0.573812f
C187 source.n10 a_n2762_n1488# 0.426145f
C188 source.t17 a_n2762_n1488# 0.069102f
C189 source.t8 a_n2762_n1488# 0.069102f
C190 source.n11 a_n2762_n1488# 0.438147f
C191 source.n12 a_n2762_n1488# 0.404522f
C192 source.t16 a_n2762_n1488# 0.069102f
C193 source.t4 a_n2762_n1488# 0.069102f
C194 source.n13 a_n2762_n1488# 0.438147f
C195 source.n14 a_n2762_n1488# 0.404522f
C196 source.t6 a_n2762_n1488# 0.069102f
C197 source.t10 a_n2762_n1488# 0.069102f
C198 source.n15 a_n2762_n1488# 0.438147f
C199 source.n16 a_n2762_n1488# 0.404522f
C200 source.t2 a_n2762_n1488# 0.069102f
C201 source.t9 a_n2762_n1488# 0.069102f
C202 source.n17 a_n2762_n1488# 0.438147f
C203 source.n18 a_n2762_n1488# 0.404522f
C204 source.t15 a_n2762_n1488# 0.573812f
C205 source.n19 a_n2762_n1488# 1.13529f
C206 source.t26 a_n2762_n1488# 0.573809f
C207 source.n20 a_n2762_n1488# 1.13529f
C208 source.t35 a_n2762_n1488# 0.069102f
C209 source.t30 a_n2762_n1488# 0.069102f
C210 source.n21 a_n2762_n1488# 0.438144f
C211 source.n22 a_n2762_n1488# 0.404525f
C212 source.t25 a_n2762_n1488# 0.069102f
C213 source.t33 a_n2762_n1488# 0.069102f
C214 source.n23 a_n2762_n1488# 0.438144f
C215 source.n24 a_n2762_n1488# 0.404525f
C216 source.t29 a_n2762_n1488# 0.069102f
C217 source.t31 a_n2762_n1488# 0.069102f
C218 source.n25 a_n2762_n1488# 0.438144f
C219 source.n26 a_n2762_n1488# 0.404525f
C220 source.t24 a_n2762_n1488# 0.069102f
C221 source.t22 a_n2762_n1488# 0.069102f
C222 source.n27 a_n2762_n1488# 0.438144f
C223 source.n28 a_n2762_n1488# 0.404525f
C224 source.t34 a_n2762_n1488# 0.573809f
C225 source.n29 a_n2762_n1488# 0.426148f
C226 source.t14 a_n2762_n1488# 0.573809f
C227 source.n30 a_n2762_n1488# 0.426148f
C228 source.t5 a_n2762_n1488# 0.069102f
C229 source.t0 a_n2762_n1488# 0.069102f
C230 source.n31 a_n2762_n1488# 0.438144f
C231 source.n32 a_n2762_n1488# 0.404525f
C232 source.t19 a_n2762_n1488# 0.069102f
C233 source.t1 a_n2762_n1488# 0.069102f
C234 source.n33 a_n2762_n1488# 0.438144f
C235 source.n34 a_n2762_n1488# 0.404525f
C236 source.t18 a_n2762_n1488# 0.069102f
C237 source.t3 a_n2762_n1488# 0.069102f
C238 source.n35 a_n2762_n1488# 0.438144f
C239 source.n36 a_n2762_n1488# 0.404525f
C240 source.t12 a_n2762_n1488# 0.069102f
C241 source.t11 a_n2762_n1488# 0.069102f
C242 source.n37 a_n2762_n1488# 0.438144f
C243 source.n38 a_n2762_n1488# 0.404525f
C244 source.t13 a_n2762_n1488# 0.573809f
C245 source.n39 a_n2762_n1488# 0.60994f
C246 source.n40 a_n2762_n1488# 0.855802f
C247 plus.n0 a_n2762_n1488# 0.05873f
C248 plus.t0 a_n2762_n1488# 0.238119f
C249 plus.t2 a_n2762_n1488# 0.238119f
C250 plus.t3 a_n2762_n1488# 0.238119f
C251 plus.n1 a_n2762_n1488# 0.058867f
C252 plus.t4 a_n2762_n1488# 0.238119f
C253 plus.n2 a_n2762_n1488# 0.14272f
C254 plus.n3 a_n2762_n1488# 0.044116f
C255 plus.t5 a_n2762_n1488# 0.238119f
C256 plus.t10 a_n2762_n1488# 0.238119f
C257 plus.n4 a_n2762_n1488# 0.14272f
C258 plus.n5 a_n2762_n1488# 0.044116f
C259 plus.t12 a_n2762_n1488# 0.238119f
C260 plus.t14 a_n2762_n1488# 0.238119f
C261 plus.n6 a_n2762_n1488# 0.141496f
C262 plus.t15 a_n2762_n1488# 0.238119f
C263 plus.n7 a_n2762_n1488# 0.150827f
C264 plus.t16 a_n2762_n1488# 0.255884f
C265 plus.n8 a_n2762_n1488# 0.123998f
C266 plus.n9 a_n2762_n1488# 0.188301f
C267 plus.n10 a_n2762_n1488# 0.044116f
C268 plus.n11 a_n2762_n1488# 0.010011f
C269 plus.n12 a_n2762_n1488# 0.14272f
C270 plus.n13 a_n2762_n1488# 0.010011f
C271 plus.n14 a_n2762_n1488# 0.044116f
C272 plus.n15 a_n2762_n1488# 0.044116f
C273 plus.n16 a_n2762_n1488# 0.044116f
C274 plus.n17 a_n2762_n1488# 0.010011f
C275 plus.n18 a_n2762_n1488# 0.14272f
C276 plus.n19 a_n2762_n1488# 0.010011f
C277 plus.n20 a_n2762_n1488# 0.044116f
C278 plus.n21 a_n2762_n1488# 0.044116f
C279 plus.n22 a_n2762_n1488# 0.044116f
C280 plus.n23 a_n2762_n1488# 0.010011f
C281 plus.n24 a_n2762_n1488# 0.141496f
C282 plus.n25 a_n2762_n1488# 0.150827f
C283 plus.n26 a_n2762_n1488# 0.140816f
C284 plus.n27 a_n2762_n1488# 0.358365f
C285 plus.n28 a_n2762_n1488# 0.05873f
C286 plus.t1 a_n2762_n1488# 0.238119f
C287 plus.t9 a_n2762_n1488# 0.238119f
C288 plus.n29 a_n2762_n1488# 0.058867f
C289 plus.t13 a_n2762_n1488# 0.238119f
C290 plus.t18 a_n2762_n1488# 0.238119f
C291 plus.n30 a_n2762_n1488# 0.14272f
C292 plus.n31 a_n2762_n1488# 0.044116f
C293 plus.t6 a_n2762_n1488# 0.238119f
C294 plus.t8 a_n2762_n1488# 0.238119f
C295 plus.n32 a_n2762_n1488# 0.14272f
C296 plus.n33 a_n2762_n1488# 0.044116f
C297 plus.t11 a_n2762_n1488# 0.238119f
C298 plus.t17 a_n2762_n1488# 0.238119f
C299 plus.n34 a_n2762_n1488# 0.141496f
C300 plus.t19 a_n2762_n1488# 0.238119f
C301 plus.n35 a_n2762_n1488# 0.150827f
C302 plus.t7 a_n2762_n1488# 0.255884f
C303 plus.n36 a_n2762_n1488# 0.123998f
C304 plus.n37 a_n2762_n1488# 0.188301f
C305 plus.n38 a_n2762_n1488# 0.044116f
C306 plus.n39 a_n2762_n1488# 0.010011f
C307 plus.n40 a_n2762_n1488# 0.14272f
C308 plus.n41 a_n2762_n1488# 0.010011f
C309 plus.n42 a_n2762_n1488# 0.044116f
C310 plus.n43 a_n2762_n1488# 0.044116f
C311 plus.n44 a_n2762_n1488# 0.044116f
C312 plus.n45 a_n2762_n1488# 0.010011f
C313 plus.n46 a_n2762_n1488# 0.14272f
C314 plus.n47 a_n2762_n1488# 0.010011f
C315 plus.n48 a_n2762_n1488# 0.044116f
C316 plus.n49 a_n2762_n1488# 0.044116f
C317 plus.n50 a_n2762_n1488# 0.044116f
C318 plus.n51 a_n2762_n1488# 0.010011f
C319 plus.n52 a_n2762_n1488# 0.141496f
C320 plus.n53 a_n2762_n1488# 0.150827f
C321 plus.n54 a_n2762_n1488# 0.140816f
C322 plus.n55 a_n2762_n1488# 1.27563f
.ends

