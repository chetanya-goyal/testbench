* NGSPICE file created from diffpair545.ext - technology: sky130A

.subckt diffpair545 minus drain_right drain_left source plus
X0 source.t17 minus.t0 drain_right.t8 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X1 drain_left.t11 plus.t0 source.t19 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X2 source.t20 plus.t1 drain_left.t10 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X3 source.t21 plus.t2 drain_left.t9 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X4 source.t16 minus.t1 drain_right.t2 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 drain_right.t11 minus.t2 source.t15 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X6 source.t22 plus.t3 drain_left.t8 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X7 source.t2 plus.t4 drain_left.t7 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X8 source.t14 minus.t3 drain_right.t0 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X9 a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X10 source.t23 plus.t5 drain_left.t6 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X11 source.t13 minus.t4 drain_right.t3 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X12 drain_right.t10 minus.t5 source.t12 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X13 drain_right.t9 minus.t6 source.t11 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X14 drain_right.t1 minus.t7 source.t10 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X15 drain_left.t5 plus.t6 source.t5 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X16 drain_left.t4 plus.t7 source.t18 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X17 a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X18 drain_right.t6 minus.t8 source.t9 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X19 source.t4 plus.t8 drain_left.t3 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X20 drain_left.t2 plus.t9 source.t1 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X21 drain_left.t1 plus.t10 source.t3 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X22 drain_left.t0 plus.t11 source.t0 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X23 a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X24 source.t8 minus.t9 drain_right.t7 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X25 source.t7 minus.t10 drain_right.t5 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X26 a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X27 drain_right.t4 minus.t11 source.t6 a_n2158_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
R0 minus.n5 minus.t8 595.851
R1 minus.n23 minus.t4 595.851
R2 minus.n4 minus.t1 572.548
R3 minus.n8 minus.t7 572.548
R4 minus.n10 minus.t9 572.548
R5 minus.n14 minus.t6 572.548
R6 minus.n16 minus.t10 572.548
R7 minus.n22 minus.t5 572.548
R8 minus.n26 minus.t0 572.548
R9 minus.n28 minus.t2 572.548
R10 minus.n32 minus.t3 572.548
R11 minus.n34 minus.t11 572.548
R12 minus.n17 minus.n16 161.3
R13 minus.n15 minus.n0 161.3
R14 minus.n14 minus.n13 161.3
R15 minus.n12 minus.n1 161.3
R16 minus.n11 minus.n10 161.3
R17 minus.n9 minus.n2 161.3
R18 minus.n8 minus.n7 161.3
R19 minus.n6 minus.n3 161.3
R20 minus.n35 minus.n34 161.3
R21 minus.n33 minus.n18 161.3
R22 minus.n32 minus.n31 161.3
R23 minus.n30 minus.n19 161.3
R24 minus.n29 minus.n28 161.3
R25 minus.n27 minus.n20 161.3
R26 minus.n26 minus.n25 161.3
R27 minus.n24 minus.n21 161.3
R28 minus.n6 minus.n5 44.8907
R29 minus.n24 minus.n23 44.8907
R30 minus.n36 minus.n17 39.7126
R31 minus.n16 minus.n15 32.8641
R32 minus.n34 minus.n33 32.8641
R33 minus.n4 minus.n3 28.4823
R34 minus.n14 minus.n1 28.4823
R35 minus.n22 minus.n21 28.4823
R36 minus.n32 minus.n19 28.4823
R37 minus.n10 minus.n9 24.1005
R38 minus.n9 minus.n8 24.1005
R39 minus.n27 minus.n26 24.1005
R40 minus.n28 minus.n27 24.1005
R41 minus.n8 minus.n3 19.7187
R42 minus.n10 minus.n1 19.7187
R43 minus.n26 minus.n21 19.7187
R44 minus.n28 minus.n19 19.7187
R45 minus.n5 minus.n4 18.4104
R46 minus.n23 minus.n22 18.4104
R47 minus.n15 minus.n14 15.3369
R48 minus.n33 minus.n32 15.3369
R49 minus.n36 minus.n35 6.64444
R50 minus.n17 minus.n0 0.189894
R51 minus.n13 minus.n0 0.189894
R52 minus.n13 minus.n12 0.189894
R53 minus.n12 minus.n11 0.189894
R54 minus.n11 minus.n2 0.189894
R55 minus.n7 minus.n2 0.189894
R56 minus.n7 minus.n6 0.189894
R57 minus.n25 minus.n24 0.189894
R58 minus.n25 minus.n20 0.189894
R59 minus.n29 minus.n20 0.189894
R60 minus.n30 minus.n29 0.189894
R61 minus.n31 minus.n30 0.189894
R62 minus.n31 minus.n18 0.189894
R63 minus.n35 minus.n18 0.189894
R64 minus minus.n36 0.188
R65 drain_right.n6 drain_right.n4 61.7676
R66 drain_right.n3 drain_right.n2 61.7121
R67 drain_right.n3 drain_right.n0 61.7121
R68 drain_right.n6 drain_right.n5 60.8798
R69 drain_right.n8 drain_right.n7 60.8798
R70 drain_right.n3 drain_right.n1 60.8796
R71 drain_right drain_right.n3 33.5262
R72 drain_right drain_right.n8 6.54115
R73 drain_right.n1 drain_right.t8 1.3205
R74 drain_right.n1 drain_right.t11 1.3205
R75 drain_right.n2 drain_right.t0 1.3205
R76 drain_right.n2 drain_right.t4 1.3205
R77 drain_right.n0 drain_right.t3 1.3205
R78 drain_right.n0 drain_right.t10 1.3205
R79 drain_right.n4 drain_right.t2 1.3205
R80 drain_right.n4 drain_right.t6 1.3205
R81 drain_right.n5 drain_right.t7 1.3205
R82 drain_right.n5 drain_right.t1 1.3205
R83 drain_right.n7 drain_right.t5 1.3205
R84 drain_right.n7 drain_right.t9 1.3205
R85 drain_right.n8 drain_right.n6 0.888431
R86 source.n5 source.t2 45.521
R87 source.n6 source.t9 45.521
R88 source.n11 source.t7 45.521
R89 source.n23 source.t6 45.5208
R90 source.n18 source.t13 45.5208
R91 source.n17 source.t19 45.5208
R92 source.n12 source.t23 45.5208
R93 source.n0 source.t18 45.5208
R94 source.n2 source.n1 44.201
R95 source.n4 source.n3 44.201
R96 source.n8 source.n7 44.201
R97 source.n10 source.n9 44.201
R98 source.n22 source.n21 44.2008
R99 source.n20 source.n19 44.2008
R100 source.n16 source.n15 44.2008
R101 source.n14 source.n13 44.2008
R102 source.n12 source.n11 24.4484
R103 source.n24 source.n0 18.7415
R104 source.n24 source.n23 5.7074
R105 source.n21 source.t15 1.3205
R106 source.n21 source.t14 1.3205
R107 source.n19 source.t12 1.3205
R108 source.n19 source.t17 1.3205
R109 source.n15 source.t0 1.3205
R110 source.n15 source.t20 1.3205
R111 source.n13 source.t1 1.3205
R112 source.n13 source.t4 1.3205
R113 source.n1 source.t5 1.3205
R114 source.n1 source.t22 1.3205
R115 source.n3 source.t3 1.3205
R116 source.n3 source.t21 1.3205
R117 source.n7 source.t10 1.3205
R118 source.n7 source.t16 1.3205
R119 source.n9 source.t11 1.3205
R120 source.n9 source.t8 1.3205
R121 source.n11 source.n10 0.888431
R122 source.n10 source.n8 0.888431
R123 source.n8 source.n6 0.888431
R124 source.n5 source.n4 0.888431
R125 source.n4 source.n2 0.888431
R126 source.n2 source.n0 0.888431
R127 source.n14 source.n12 0.888431
R128 source.n16 source.n14 0.888431
R129 source.n17 source.n16 0.888431
R130 source.n20 source.n18 0.888431
R131 source.n22 source.n20 0.888431
R132 source.n23 source.n22 0.888431
R133 source.n6 source.n5 0.470328
R134 source.n18 source.n17 0.470328
R135 source source.n24 0.188
R136 plus.n5 plus.t4 595.851
R137 plus.n23 plus.t0 595.851
R138 plus.n16 plus.t7 572.548
R139 plus.n14 plus.t3 572.548
R140 plus.n2 plus.t6 572.548
R141 plus.n8 plus.t2 572.548
R142 plus.n4 plus.t10 572.548
R143 plus.n34 plus.t5 572.548
R144 plus.n32 plus.t9 572.548
R145 plus.n20 plus.t8 572.548
R146 plus.n26 plus.t11 572.548
R147 plus.n22 plus.t1 572.548
R148 plus.n7 plus.n6 161.3
R149 plus.n8 plus.n3 161.3
R150 plus.n10 plus.n9 161.3
R151 plus.n11 plus.n2 161.3
R152 plus.n13 plus.n12 161.3
R153 plus.n14 plus.n1 161.3
R154 plus.n15 plus.n0 161.3
R155 plus.n17 plus.n16 161.3
R156 plus.n25 plus.n24 161.3
R157 plus.n26 plus.n21 161.3
R158 plus.n28 plus.n27 161.3
R159 plus.n29 plus.n20 161.3
R160 plus.n31 plus.n30 161.3
R161 plus.n32 plus.n19 161.3
R162 plus.n33 plus.n18 161.3
R163 plus.n35 plus.n34 161.3
R164 plus.n6 plus.n5 44.8907
R165 plus.n24 plus.n23 44.8907
R166 plus.n16 plus.n15 32.8641
R167 plus.n34 plus.n33 32.8641
R168 plus plus.n35 32.4574
R169 plus.n14 plus.n13 28.4823
R170 plus.n7 plus.n4 28.4823
R171 plus.n32 plus.n31 28.4823
R172 plus.n25 plus.n22 28.4823
R173 plus.n9 plus.n8 24.1005
R174 plus.n9 plus.n2 24.1005
R175 plus.n27 plus.n20 24.1005
R176 plus.n27 plus.n26 24.1005
R177 plus.n13 plus.n2 19.7187
R178 plus.n8 plus.n7 19.7187
R179 plus.n31 plus.n20 19.7187
R180 plus.n26 plus.n25 19.7187
R181 plus.n5 plus.n4 18.4104
R182 plus.n23 plus.n22 18.4104
R183 plus.n15 plus.n14 15.3369
R184 plus.n33 plus.n32 15.3369
R185 plus plus.n17 13.4247
R186 plus.n6 plus.n3 0.189894
R187 plus.n10 plus.n3 0.189894
R188 plus.n11 plus.n10 0.189894
R189 plus.n12 plus.n11 0.189894
R190 plus.n12 plus.n1 0.189894
R191 plus.n1 plus.n0 0.189894
R192 plus.n17 plus.n0 0.189894
R193 plus.n35 plus.n18 0.189894
R194 plus.n19 plus.n18 0.189894
R195 plus.n30 plus.n19 0.189894
R196 plus.n30 plus.n29 0.189894
R197 plus.n29 plus.n28 0.189894
R198 plus.n28 plus.n21 0.189894
R199 plus.n24 plus.n21 0.189894
R200 drain_left.n6 drain_left.n4 61.7677
R201 drain_left.n3 drain_left.n2 61.7121
R202 drain_left.n3 drain_left.n0 61.7121
R203 drain_left.n6 drain_left.n5 60.8798
R204 drain_left.n8 drain_left.n7 60.8796
R205 drain_left.n3 drain_left.n1 60.8796
R206 drain_left drain_left.n3 34.0795
R207 drain_left drain_left.n8 6.54115
R208 drain_left.n1 drain_left.t3 1.3205
R209 drain_left.n1 drain_left.t0 1.3205
R210 drain_left.n2 drain_left.t10 1.3205
R211 drain_left.n2 drain_left.t11 1.3205
R212 drain_left.n0 drain_left.t6 1.3205
R213 drain_left.n0 drain_left.t2 1.3205
R214 drain_left.n7 drain_left.t8 1.3205
R215 drain_left.n7 drain_left.t4 1.3205
R216 drain_left.n5 drain_left.t9 1.3205
R217 drain_left.n5 drain_left.t5 1.3205
R218 drain_left.n4 drain_left.t7 1.3205
R219 drain_left.n4 drain_left.t1 1.3205
R220 drain_left.n8 drain_left.n6 0.888431
C0 minus drain_right 9.736401f
C1 source drain_left 18.6782f
C2 source drain_right 18.680199f
C3 minus plus 6.39035f
C4 drain_left drain_right 1.08491f
C5 source plus 9.52671f
C6 drain_left plus 9.948139f
C7 minus source 9.51267f
C8 minus drain_left 0.17184f
C9 drain_right plus 0.366822f
C10 drain_right a_n2158_n3888# 6.768559f
C11 drain_left a_n2158_n3888# 7.07786f
C12 source a_n2158_n3888# 10.790743f
C13 minus a_n2158_n3888# 8.711685f
C14 plus a_n2158_n3888# 10.56617f
C15 drain_left.t6 a_n2158_n3888# 0.322932f
C16 drain_left.t2 a_n2158_n3888# 0.322932f
C17 drain_left.n0 a_n2158_n3888# 2.92413f
C18 drain_left.t3 a_n2158_n3888# 0.322932f
C19 drain_left.t0 a_n2158_n3888# 0.322932f
C20 drain_left.n1 a_n2158_n3888# 2.91893f
C21 drain_left.t10 a_n2158_n3888# 0.322932f
C22 drain_left.t11 a_n2158_n3888# 0.322932f
C23 drain_left.n2 a_n2158_n3888# 2.92413f
C24 drain_left.n3 a_n2158_n3888# 2.70645f
C25 drain_left.t7 a_n2158_n3888# 0.322932f
C26 drain_left.t1 a_n2158_n3888# 0.322932f
C27 drain_left.n4 a_n2158_n3888# 2.92454f
C28 drain_left.t9 a_n2158_n3888# 0.322932f
C29 drain_left.t5 a_n2158_n3888# 0.322932f
C30 drain_left.n5 a_n2158_n3888# 2.91893f
C31 drain_left.n6 a_n2158_n3888# 0.763436f
C32 drain_left.t8 a_n2158_n3888# 0.322932f
C33 drain_left.t4 a_n2158_n3888# 0.322932f
C34 drain_left.n7 a_n2158_n3888# 2.91892f
C35 drain_left.n8 a_n2158_n3888# 0.620017f
C36 plus.n0 a_n2158_n3888# 0.042012f
C37 plus.t7 a_n2158_n3888# 1.25354f
C38 plus.t3 a_n2158_n3888# 1.25354f
C39 plus.n1 a_n2158_n3888# 0.042012f
C40 plus.t6 a_n2158_n3888# 1.25354f
C41 plus.n2 a_n2158_n3888# 0.483746f
C42 plus.n3 a_n2158_n3888# 0.042012f
C43 plus.t2 a_n2158_n3888# 1.25354f
C44 plus.t10 a_n2158_n3888# 1.25354f
C45 plus.n4 a_n2158_n3888# 0.488445f
C46 plus.t4 a_n2158_n3888# 1.27246f
C47 plus.n5 a_n2158_n3888# 0.46859f
C48 plus.n6 a_n2158_n3888# 0.176245f
C49 plus.n7 a_n2158_n3888# 0.009533f
C50 plus.n8 a_n2158_n3888# 0.483746f
C51 plus.n9 a_n2158_n3888# 0.009533f
C52 plus.n10 a_n2158_n3888# 0.042012f
C53 plus.n11 a_n2158_n3888# 0.042012f
C54 plus.n12 a_n2158_n3888# 0.042012f
C55 plus.n13 a_n2158_n3888# 0.009533f
C56 plus.n14 a_n2158_n3888# 0.483746f
C57 plus.n15 a_n2158_n3888# 0.009533f
C58 plus.n16 a_n2158_n3888# 0.481804f
C59 plus.n17 a_n2158_n3888# 0.545145f
C60 plus.n18 a_n2158_n3888# 0.042012f
C61 plus.t5 a_n2158_n3888# 1.25354f
C62 plus.n19 a_n2158_n3888# 0.042012f
C63 plus.t9 a_n2158_n3888# 1.25354f
C64 plus.t8 a_n2158_n3888# 1.25354f
C65 plus.n20 a_n2158_n3888# 0.483746f
C66 plus.n21 a_n2158_n3888# 0.042012f
C67 plus.t11 a_n2158_n3888# 1.25354f
C68 plus.t1 a_n2158_n3888# 1.25354f
C69 plus.n22 a_n2158_n3888# 0.488445f
C70 plus.t0 a_n2158_n3888# 1.27246f
C71 plus.n23 a_n2158_n3888# 0.46859f
C72 plus.n24 a_n2158_n3888# 0.176245f
C73 plus.n25 a_n2158_n3888# 0.009533f
C74 plus.n26 a_n2158_n3888# 0.483746f
C75 plus.n27 a_n2158_n3888# 0.009533f
C76 plus.n28 a_n2158_n3888# 0.042012f
C77 plus.n29 a_n2158_n3888# 0.042012f
C78 plus.n30 a_n2158_n3888# 0.042012f
C79 plus.n31 a_n2158_n3888# 0.009533f
C80 plus.n32 a_n2158_n3888# 0.483746f
C81 plus.n33 a_n2158_n3888# 0.009533f
C82 plus.n34 a_n2158_n3888# 0.481804f
C83 plus.n35 a_n2158_n3888# 1.41918f
C84 source.t18 a_n2158_n3888# 2.87583f
C85 source.n0 a_n2158_n3888# 1.3708f
C86 source.t5 a_n2158_n3888# 0.256619f
C87 source.t22 a_n2158_n3888# 0.256619f
C88 source.n1 a_n2158_n3888# 2.25418f
C89 source.n2 a_n2158_n3888# 0.337131f
C90 source.t3 a_n2158_n3888# 0.256619f
C91 source.t21 a_n2158_n3888# 0.256619f
C92 source.n3 a_n2158_n3888# 2.25418f
C93 source.n4 a_n2158_n3888# 0.337131f
C94 source.t2 a_n2158_n3888# 2.87583f
C95 source.n5 a_n2158_n3888# 0.386184f
C96 source.t9 a_n2158_n3888# 2.87583f
C97 source.n6 a_n2158_n3888# 0.386184f
C98 source.t10 a_n2158_n3888# 0.256619f
C99 source.t16 a_n2158_n3888# 0.256619f
C100 source.n7 a_n2158_n3888# 2.25418f
C101 source.n8 a_n2158_n3888# 0.337131f
C102 source.t11 a_n2158_n3888# 0.256619f
C103 source.t8 a_n2158_n3888# 0.256619f
C104 source.n9 a_n2158_n3888# 2.25418f
C105 source.n10 a_n2158_n3888# 0.337131f
C106 source.t7 a_n2158_n3888# 2.87583f
C107 source.n11 a_n2158_n3888# 1.74008f
C108 source.t23 a_n2158_n3888# 2.87583f
C109 source.n12 a_n2158_n3888# 1.74008f
C110 source.t1 a_n2158_n3888# 0.256619f
C111 source.t4 a_n2158_n3888# 0.256619f
C112 source.n13 a_n2158_n3888# 2.25418f
C113 source.n14 a_n2158_n3888# 0.337134f
C114 source.t0 a_n2158_n3888# 0.256619f
C115 source.t20 a_n2158_n3888# 0.256619f
C116 source.n15 a_n2158_n3888# 2.25418f
C117 source.n16 a_n2158_n3888# 0.337134f
C118 source.t19 a_n2158_n3888# 2.87583f
C119 source.n17 a_n2158_n3888# 0.386188f
C120 source.t13 a_n2158_n3888# 2.87583f
C121 source.n18 a_n2158_n3888# 0.386188f
C122 source.t12 a_n2158_n3888# 0.256619f
C123 source.t17 a_n2158_n3888# 0.256619f
C124 source.n19 a_n2158_n3888# 2.25418f
C125 source.n20 a_n2158_n3888# 0.337134f
C126 source.t15 a_n2158_n3888# 0.256619f
C127 source.t14 a_n2158_n3888# 0.256619f
C128 source.n21 a_n2158_n3888# 2.25418f
C129 source.n22 a_n2158_n3888# 0.337134f
C130 source.t6 a_n2158_n3888# 2.87583f
C131 source.n23 a_n2158_n3888# 0.527407f
C132 source.n24 a_n2158_n3888# 1.59735f
C133 drain_right.t3 a_n2158_n3888# 0.321873f
C134 drain_right.t10 a_n2158_n3888# 0.321873f
C135 drain_right.n0 a_n2158_n3888# 2.91455f
C136 drain_right.t8 a_n2158_n3888# 0.321873f
C137 drain_right.t11 a_n2158_n3888# 0.321873f
C138 drain_right.n1 a_n2158_n3888# 2.90936f
C139 drain_right.t0 a_n2158_n3888# 0.321873f
C140 drain_right.t4 a_n2158_n3888# 0.321873f
C141 drain_right.n2 a_n2158_n3888# 2.91455f
C142 drain_right.n3 a_n2158_n3888# 2.64133f
C143 drain_right.t2 a_n2158_n3888# 0.321873f
C144 drain_right.t6 a_n2158_n3888# 0.321873f
C145 drain_right.n4 a_n2158_n3888# 2.91494f
C146 drain_right.t7 a_n2158_n3888# 0.321873f
C147 drain_right.t1 a_n2158_n3888# 0.321873f
C148 drain_right.n5 a_n2158_n3888# 2.90936f
C149 drain_right.n6 a_n2158_n3888# 0.760943f
C150 drain_right.t5 a_n2158_n3888# 0.321873f
C151 drain_right.t9 a_n2158_n3888# 0.321873f
C152 drain_right.n7 a_n2158_n3888# 2.90936f
C153 drain_right.n8 a_n2158_n3888# 0.617974f
C154 minus.n0 a_n2158_n3888# 0.041549f
C155 minus.n1 a_n2158_n3888# 0.009428f
C156 minus.t6 a_n2158_n3888# 1.23974f
C157 minus.n2 a_n2158_n3888# 0.041549f
C158 minus.n3 a_n2158_n3888# 0.009428f
C159 minus.t7 a_n2158_n3888# 1.23974f
C160 minus.t8 a_n2158_n3888# 1.25845f
C161 minus.t1 a_n2158_n3888# 1.23974f
C162 minus.n4 a_n2158_n3888# 0.483068f
C163 minus.n5 a_n2158_n3888# 0.463431f
C164 minus.n6 a_n2158_n3888# 0.174304f
C165 minus.n7 a_n2158_n3888# 0.041549f
C166 minus.n8 a_n2158_n3888# 0.478421f
C167 minus.n9 a_n2158_n3888# 0.009428f
C168 minus.t9 a_n2158_n3888# 1.23974f
C169 minus.n10 a_n2158_n3888# 0.478421f
C170 minus.n11 a_n2158_n3888# 0.041549f
C171 minus.n12 a_n2158_n3888# 0.041549f
C172 minus.n13 a_n2158_n3888# 0.041549f
C173 minus.n14 a_n2158_n3888# 0.478421f
C174 minus.n15 a_n2158_n3888# 0.009428f
C175 minus.t10 a_n2158_n3888# 1.23974f
C176 minus.n16 a_n2158_n3888# 0.4765f
C177 minus.n17 a_n2158_n3888# 1.69714f
C178 minus.n18 a_n2158_n3888# 0.041549f
C179 minus.n19 a_n2158_n3888# 0.009428f
C180 minus.n20 a_n2158_n3888# 0.041549f
C181 minus.n21 a_n2158_n3888# 0.009428f
C182 minus.t4 a_n2158_n3888# 1.25845f
C183 minus.t5 a_n2158_n3888# 1.23974f
C184 minus.n22 a_n2158_n3888# 0.483068f
C185 minus.n23 a_n2158_n3888# 0.463431f
C186 minus.n24 a_n2158_n3888# 0.174304f
C187 minus.n25 a_n2158_n3888# 0.041549f
C188 minus.t0 a_n2158_n3888# 1.23974f
C189 minus.n26 a_n2158_n3888# 0.478421f
C190 minus.n27 a_n2158_n3888# 0.009428f
C191 minus.t2 a_n2158_n3888# 1.23974f
C192 minus.n28 a_n2158_n3888# 0.478421f
C193 minus.n29 a_n2158_n3888# 0.041549f
C194 minus.n30 a_n2158_n3888# 0.041549f
C195 minus.n31 a_n2158_n3888# 0.041549f
C196 minus.t3 a_n2158_n3888# 1.23974f
C197 minus.n32 a_n2158_n3888# 0.478421f
C198 minus.n33 a_n2158_n3888# 0.009428f
C199 minus.t11 a_n2158_n3888# 1.23974f
C200 minus.n34 a_n2158_n3888# 0.4765f
C201 minus.n35 a_n2158_n3888# 0.285683f
C202 minus.n36 a_n2158_n3888# 2.03639f
.ends

