* NGSPICE file created from diffpair294.ext - technology: sky130A

.subckt diffpair294 minus drain_right drain_left source plus
X0 a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.6
X1 source.t19 plus.t0 drain_left.t7 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X2 a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X3 drain_right.t9 minus.t0 source.t5 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X4 drain_right.t8 minus.t1 source.t1 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X5 drain_left.t4 plus.t1 source.t18 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X6 drain_left.t0 plus.t2 source.t17 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X7 source.t7 minus.t2 drain_right.t7 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X8 source.t3 minus.t3 drain_right.t6 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X9 drain_left.t5 plus.t3 source.t16 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X10 drain_right.t5 minus.t4 source.t8 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X11 source.t15 plus.t4 drain_left.t2 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X12 source.t14 plus.t5 drain_left.t6 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X13 source.t6 minus.t5 drain_right.t4 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X14 drain_left.t8 plus.t6 source.t13 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X15 drain_right.t3 minus.t6 source.t0 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X16 source.t12 plus.t7 drain_left.t3 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X17 drain_left.t1 plus.t8 source.t11 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X18 drain_left.t9 plus.t9 source.t10 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X19 a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X20 drain_right.t2 minus.t7 source.t9 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X21 source.t2 minus.t8 drain_right.t1 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X22 a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X23 drain_right.t0 minus.t9 source.t4 a_n1832_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
R0 plus.n3 plus.t8 332.673
R1 plus.n13 plus.t3 332.673
R2 plus.n8 plus.t2 306.473
R3 plus.n6 plus.t5 306.473
R4 plus.n5 plus.t6 306.473
R5 plus.n4 plus.t7 306.473
R6 plus.n18 plus.t9 306.473
R7 plus.n16 plus.t4 306.473
R8 plus.n15 plus.t1 306.473
R9 plus.n14 plus.t0 306.473
R10 plus.n6 plus.n1 161.3
R11 plus.n7 plus.n0 161.3
R12 plus.n9 plus.n8 161.3
R13 plus.n16 plus.n11 161.3
R14 plus.n17 plus.n10 161.3
R15 plus.n19 plus.n18 161.3
R16 plus.n5 plus.n2 80.6037
R17 plus.n15 plus.n12 80.6037
R18 plus.n6 plus.n5 48.2005
R19 plus.n5 plus.n4 48.2005
R20 plus.n16 plus.n15 48.2005
R21 plus.n15 plus.n14 48.2005
R22 plus.n8 plus.n7 45.2793
R23 plus.n18 plus.n17 45.2793
R24 plus.n3 plus.n2 45.1669
R25 plus.n13 plus.n12 45.1669
R26 plus plus.n19 27.7699
R27 plus.n4 plus.n3 14.3992
R28 plus.n14 plus.n13 14.3992
R29 plus plus.n9 9.97209
R30 plus.n7 plus.n6 2.92171
R31 plus.n17 plus.n16 2.92171
R32 plus.n2 plus.n1 0.285035
R33 plus.n12 plus.n11 0.285035
R34 plus.n1 plus.n0 0.189894
R35 plus.n9 plus.n0 0.189894
R36 plus.n19 plus.n10 0.189894
R37 plus.n11 plus.n10 0.189894
R38 drain_left.n26 drain_left.n0 289.615
R39 drain_left.n61 drain_left.n35 289.615
R40 drain_left.n11 drain_left.n10 185
R41 drain_left.n8 drain_left.n7 185
R42 drain_left.n17 drain_left.n16 185
R43 drain_left.n19 drain_left.n18 185
R44 drain_left.n4 drain_left.n3 185
R45 drain_left.n25 drain_left.n24 185
R46 drain_left.n27 drain_left.n26 185
R47 drain_left.n62 drain_left.n61 185
R48 drain_left.n60 drain_left.n59 185
R49 drain_left.n39 drain_left.n38 185
R50 drain_left.n54 drain_left.n53 185
R51 drain_left.n52 drain_left.n51 185
R52 drain_left.n43 drain_left.n42 185
R53 drain_left.n46 drain_left.n45 185
R54 drain_left.t9 drain_left.n9 147.661
R55 drain_left.t1 drain_left.n44 147.661
R56 drain_left.n10 drain_left.n7 104.615
R57 drain_left.n17 drain_left.n7 104.615
R58 drain_left.n18 drain_left.n17 104.615
R59 drain_left.n18 drain_left.n3 104.615
R60 drain_left.n25 drain_left.n3 104.615
R61 drain_left.n26 drain_left.n25 104.615
R62 drain_left.n61 drain_left.n60 104.615
R63 drain_left.n60 drain_left.n38 104.615
R64 drain_left.n53 drain_left.n38 104.615
R65 drain_left.n53 drain_left.n52 104.615
R66 drain_left.n52 drain_left.n42 104.615
R67 drain_left.n45 drain_left.n42 104.615
R68 drain_left.n34 drain_left.n33 67.7366
R69 drain_left.n67 drain_left.n66 67.1908
R70 drain_left.n69 drain_left.n68 67.1907
R71 drain_left.n32 drain_left.n31 67.1907
R72 drain_left.n10 drain_left.t9 52.3082
R73 drain_left.n45 drain_left.t1 52.3082
R74 drain_left.n32 drain_left.n30 49.6659
R75 drain_left.n67 drain_left.n65 49.6659
R76 drain_left drain_left.n34 26.2289
R77 drain_left.n11 drain_left.n9 15.6674
R78 drain_left.n46 drain_left.n44 15.6674
R79 drain_left.n12 drain_left.n8 12.8005
R80 drain_left.n47 drain_left.n43 12.8005
R81 drain_left.n16 drain_left.n15 12.0247
R82 drain_left.n51 drain_left.n50 12.0247
R83 drain_left.n19 drain_left.n6 11.249
R84 drain_left.n54 drain_left.n41 11.249
R85 drain_left.n20 drain_left.n4 10.4732
R86 drain_left.n55 drain_left.n39 10.4732
R87 drain_left.n24 drain_left.n23 9.69747
R88 drain_left.n59 drain_left.n58 9.69747
R89 drain_left.n30 drain_left.n29 9.45567
R90 drain_left.n65 drain_left.n64 9.45567
R91 drain_left.n29 drain_left.n28 9.3005
R92 drain_left.n2 drain_left.n1 9.3005
R93 drain_left.n23 drain_left.n22 9.3005
R94 drain_left.n21 drain_left.n20 9.3005
R95 drain_left.n6 drain_left.n5 9.3005
R96 drain_left.n15 drain_left.n14 9.3005
R97 drain_left.n13 drain_left.n12 9.3005
R98 drain_left.n64 drain_left.n63 9.3005
R99 drain_left.n37 drain_left.n36 9.3005
R100 drain_left.n58 drain_left.n57 9.3005
R101 drain_left.n56 drain_left.n55 9.3005
R102 drain_left.n41 drain_left.n40 9.3005
R103 drain_left.n50 drain_left.n49 9.3005
R104 drain_left.n48 drain_left.n47 9.3005
R105 drain_left.n27 drain_left.n2 8.92171
R106 drain_left.n62 drain_left.n37 8.92171
R107 drain_left.n28 drain_left.n0 8.14595
R108 drain_left.n63 drain_left.n35 8.14595
R109 drain_left drain_left.n69 6.45494
R110 drain_left.n30 drain_left.n0 5.81868
R111 drain_left.n65 drain_left.n35 5.81868
R112 drain_left.n28 drain_left.n27 5.04292
R113 drain_left.n63 drain_left.n62 5.04292
R114 drain_left.n13 drain_left.n9 4.38594
R115 drain_left.n48 drain_left.n44 4.38594
R116 drain_left.n24 drain_left.n2 4.26717
R117 drain_left.n59 drain_left.n37 4.26717
R118 drain_left.n23 drain_left.n4 3.49141
R119 drain_left.n58 drain_left.n39 3.49141
R120 drain_left.n33 drain_left.t7 3.3005
R121 drain_left.n33 drain_left.t5 3.3005
R122 drain_left.n31 drain_left.t2 3.3005
R123 drain_left.n31 drain_left.t4 3.3005
R124 drain_left.n68 drain_left.t6 3.3005
R125 drain_left.n68 drain_left.t0 3.3005
R126 drain_left.n66 drain_left.t3 3.3005
R127 drain_left.n66 drain_left.t8 3.3005
R128 drain_left.n20 drain_left.n19 2.71565
R129 drain_left.n55 drain_left.n54 2.71565
R130 drain_left.n16 drain_left.n6 1.93989
R131 drain_left.n51 drain_left.n41 1.93989
R132 drain_left.n15 drain_left.n8 1.16414
R133 drain_left.n50 drain_left.n43 1.16414
R134 drain_left.n69 drain_left.n67 0.802224
R135 drain_left.n12 drain_left.n11 0.388379
R136 drain_left.n47 drain_left.n46 0.388379
R137 drain_left.n14 drain_left.n13 0.155672
R138 drain_left.n14 drain_left.n5 0.155672
R139 drain_left.n21 drain_left.n5 0.155672
R140 drain_left.n22 drain_left.n21 0.155672
R141 drain_left.n22 drain_left.n1 0.155672
R142 drain_left.n29 drain_left.n1 0.155672
R143 drain_left.n64 drain_left.n36 0.155672
R144 drain_left.n57 drain_left.n36 0.155672
R145 drain_left.n57 drain_left.n56 0.155672
R146 drain_left.n56 drain_left.n40 0.155672
R147 drain_left.n49 drain_left.n40 0.155672
R148 drain_left.n49 drain_left.n48 0.155672
R149 drain_left.n34 drain_left.n32 0.145585
R150 source.n138 source.n112 289.615
R151 source.n102 source.n76 289.615
R152 source.n26 source.n0 289.615
R153 source.n62 source.n36 289.615
R154 source.n123 source.n122 185
R155 source.n120 source.n119 185
R156 source.n129 source.n128 185
R157 source.n131 source.n130 185
R158 source.n116 source.n115 185
R159 source.n137 source.n136 185
R160 source.n139 source.n138 185
R161 source.n87 source.n86 185
R162 source.n84 source.n83 185
R163 source.n93 source.n92 185
R164 source.n95 source.n94 185
R165 source.n80 source.n79 185
R166 source.n101 source.n100 185
R167 source.n103 source.n102 185
R168 source.n27 source.n26 185
R169 source.n25 source.n24 185
R170 source.n4 source.n3 185
R171 source.n19 source.n18 185
R172 source.n17 source.n16 185
R173 source.n8 source.n7 185
R174 source.n11 source.n10 185
R175 source.n63 source.n62 185
R176 source.n61 source.n60 185
R177 source.n40 source.n39 185
R178 source.n55 source.n54 185
R179 source.n53 source.n52 185
R180 source.n44 source.n43 185
R181 source.n47 source.n46 185
R182 source.t9 source.n121 147.661
R183 source.t16 source.n85 147.661
R184 source.t17 source.n9 147.661
R185 source.t0 source.n45 147.661
R186 source.n122 source.n119 104.615
R187 source.n129 source.n119 104.615
R188 source.n130 source.n129 104.615
R189 source.n130 source.n115 104.615
R190 source.n137 source.n115 104.615
R191 source.n138 source.n137 104.615
R192 source.n86 source.n83 104.615
R193 source.n93 source.n83 104.615
R194 source.n94 source.n93 104.615
R195 source.n94 source.n79 104.615
R196 source.n101 source.n79 104.615
R197 source.n102 source.n101 104.615
R198 source.n26 source.n25 104.615
R199 source.n25 source.n3 104.615
R200 source.n18 source.n3 104.615
R201 source.n18 source.n17 104.615
R202 source.n17 source.n7 104.615
R203 source.n10 source.n7 104.615
R204 source.n62 source.n61 104.615
R205 source.n61 source.n39 104.615
R206 source.n54 source.n39 104.615
R207 source.n54 source.n53 104.615
R208 source.n53 source.n43 104.615
R209 source.n46 source.n43 104.615
R210 source.n122 source.t9 52.3082
R211 source.n86 source.t16 52.3082
R212 source.n10 source.t17 52.3082
R213 source.n46 source.t0 52.3082
R214 source.n33 source.n32 50.512
R215 source.n35 source.n34 50.512
R216 source.n69 source.n68 50.512
R217 source.n71 source.n70 50.512
R218 source.n111 source.n110 50.5119
R219 source.n109 source.n108 50.5119
R220 source.n75 source.n74 50.5119
R221 source.n73 source.n72 50.5119
R222 source.n143 source.n142 32.1853
R223 source.n107 source.n106 32.1853
R224 source.n31 source.n30 32.1853
R225 source.n67 source.n66 32.1853
R226 source.n73 source.n71 18.3457
R227 source.n123 source.n121 15.6674
R228 source.n87 source.n85 15.6674
R229 source.n11 source.n9 15.6674
R230 source.n47 source.n45 15.6674
R231 source.n124 source.n120 12.8005
R232 source.n88 source.n84 12.8005
R233 source.n12 source.n8 12.8005
R234 source.n48 source.n44 12.8005
R235 source.n128 source.n127 12.0247
R236 source.n92 source.n91 12.0247
R237 source.n16 source.n15 12.0247
R238 source.n52 source.n51 12.0247
R239 source.n144 source.n31 11.8802
R240 source.n131 source.n118 11.249
R241 source.n95 source.n82 11.249
R242 source.n19 source.n6 11.249
R243 source.n55 source.n42 11.249
R244 source.n132 source.n116 10.4732
R245 source.n96 source.n80 10.4732
R246 source.n20 source.n4 10.4732
R247 source.n56 source.n40 10.4732
R248 source.n136 source.n135 9.69747
R249 source.n100 source.n99 9.69747
R250 source.n24 source.n23 9.69747
R251 source.n60 source.n59 9.69747
R252 source.n142 source.n141 9.45567
R253 source.n106 source.n105 9.45567
R254 source.n30 source.n29 9.45567
R255 source.n66 source.n65 9.45567
R256 source.n141 source.n140 9.3005
R257 source.n114 source.n113 9.3005
R258 source.n135 source.n134 9.3005
R259 source.n133 source.n132 9.3005
R260 source.n118 source.n117 9.3005
R261 source.n127 source.n126 9.3005
R262 source.n125 source.n124 9.3005
R263 source.n105 source.n104 9.3005
R264 source.n78 source.n77 9.3005
R265 source.n99 source.n98 9.3005
R266 source.n97 source.n96 9.3005
R267 source.n82 source.n81 9.3005
R268 source.n91 source.n90 9.3005
R269 source.n89 source.n88 9.3005
R270 source.n29 source.n28 9.3005
R271 source.n2 source.n1 9.3005
R272 source.n23 source.n22 9.3005
R273 source.n21 source.n20 9.3005
R274 source.n6 source.n5 9.3005
R275 source.n15 source.n14 9.3005
R276 source.n13 source.n12 9.3005
R277 source.n65 source.n64 9.3005
R278 source.n38 source.n37 9.3005
R279 source.n59 source.n58 9.3005
R280 source.n57 source.n56 9.3005
R281 source.n42 source.n41 9.3005
R282 source.n51 source.n50 9.3005
R283 source.n49 source.n48 9.3005
R284 source.n139 source.n114 8.92171
R285 source.n103 source.n78 8.92171
R286 source.n27 source.n2 8.92171
R287 source.n63 source.n38 8.92171
R288 source.n140 source.n112 8.14595
R289 source.n104 source.n76 8.14595
R290 source.n28 source.n0 8.14595
R291 source.n64 source.n36 8.14595
R292 source.n142 source.n112 5.81868
R293 source.n106 source.n76 5.81868
R294 source.n30 source.n0 5.81868
R295 source.n66 source.n36 5.81868
R296 source.n144 source.n143 5.66429
R297 source.n140 source.n139 5.04292
R298 source.n104 source.n103 5.04292
R299 source.n28 source.n27 5.04292
R300 source.n64 source.n63 5.04292
R301 source.n125 source.n121 4.38594
R302 source.n89 source.n85 4.38594
R303 source.n13 source.n9 4.38594
R304 source.n49 source.n45 4.38594
R305 source.n136 source.n114 4.26717
R306 source.n100 source.n78 4.26717
R307 source.n24 source.n2 4.26717
R308 source.n60 source.n38 4.26717
R309 source.n135 source.n116 3.49141
R310 source.n99 source.n80 3.49141
R311 source.n23 source.n4 3.49141
R312 source.n59 source.n40 3.49141
R313 source.n110 source.t4 3.3005
R314 source.n110 source.t3 3.3005
R315 source.n108 source.t1 3.3005
R316 source.n108 source.t2 3.3005
R317 source.n74 source.t18 3.3005
R318 source.n74 source.t19 3.3005
R319 source.n72 source.t10 3.3005
R320 source.n72 source.t15 3.3005
R321 source.n32 source.t13 3.3005
R322 source.n32 source.t14 3.3005
R323 source.n34 source.t11 3.3005
R324 source.n34 source.t12 3.3005
R325 source.n68 source.t8 3.3005
R326 source.n68 source.t6 3.3005
R327 source.n70 source.t5 3.3005
R328 source.n70 source.t7 3.3005
R329 source.n132 source.n131 2.71565
R330 source.n96 source.n95 2.71565
R331 source.n20 source.n19 2.71565
R332 source.n56 source.n55 2.71565
R333 source.n128 source.n118 1.93989
R334 source.n92 source.n82 1.93989
R335 source.n16 source.n6 1.93989
R336 source.n52 source.n42 1.93989
R337 source.n127 source.n120 1.16414
R338 source.n91 source.n84 1.16414
R339 source.n15 source.n8 1.16414
R340 source.n51 source.n44 1.16414
R341 source.n67 source.n35 0.87119
R342 source.n109 source.n107 0.87119
R343 source.n71 source.n69 0.802224
R344 source.n69 source.n67 0.802224
R345 source.n35 source.n33 0.802224
R346 source.n33 source.n31 0.802224
R347 source.n75 source.n73 0.802224
R348 source.n107 source.n75 0.802224
R349 source.n111 source.n109 0.802224
R350 source.n143 source.n111 0.802224
R351 source.n124 source.n123 0.388379
R352 source.n88 source.n87 0.388379
R353 source.n12 source.n11 0.388379
R354 source.n48 source.n47 0.388379
R355 source source.n144 0.188
R356 source.n126 source.n125 0.155672
R357 source.n126 source.n117 0.155672
R358 source.n133 source.n117 0.155672
R359 source.n134 source.n133 0.155672
R360 source.n134 source.n113 0.155672
R361 source.n141 source.n113 0.155672
R362 source.n90 source.n89 0.155672
R363 source.n90 source.n81 0.155672
R364 source.n97 source.n81 0.155672
R365 source.n98 source.n97 0.155672
R366 source.n98 source.n77 0.155672
R367 source.n105 source.n77 0.155672
R368 source.n29 source.n1 0.155672
R369 source.n22 source.n1 0.155672
R370 source.n22 source.n21 0.155672
R371 source.n21 source.n5 0.155672
R372 source.n14 source.n5 0.155672
R373 source.n14 source.n13 0.155672
R374 source.n65 source.n37 0.155672
R375 source.n58 source.n37 0.155672
R376 source.n58 source.n57 0.155672
R377 source.n57 source.n41 0.155672
R378 source.n50 source.n41 0.155672
R379 source.n50 source.n49 0.155672
R380 minus.n3 minus.t6 332.673
R381 minus.n13 minus.t1 332.673
R382 minus.n2 minus.t5 306.473
R383 minus.n1 minus.t4 306.473
R384 minus.n6 minus.t2 306.473
R385 minus.n8 minus.t0 306.473
R386 minus.n12 minus.t8 306.473
R387 minus.n11 minus.t9 306.473
R388 minus.n16 minus.t3 306.473
R389 minus.n18 minus.t7 306.473
R390 minus.n9 minus.n8 161.3
R391 minus.n7 minus.n0 161.3
R392 minus.n6 minus.n5 161.3
R393 minus.n19 minus.n18 161.3
R394 minus.n17 minus.n10 161.3
R395 minus.n16 minus.n15 161.3
R396 minus.n4 minus.n1 80.6037
R397 minus.n14 minus.n11 80.6037
R398 minus.n2 minus.n1 48.2005
R399 minus.n6 minus.n1 48.2005
R400 minus.n12 minus.n11 48.2005
R401 minus.n16 minus.n11 48.2005
R402 minus.n8 minus.n7 45.2793
R403 minus.n18 minus.n17 45.2793
R404 minus.n4 minus.n3 45.1669
R405 minus.n14 minus.n13 45.1669
R406 minus.n20 minus.n9 31.616
R407 minus.n3 minus.n2 14.3992
R408 minus.n13 minus.n12 14.3992
R409 minus.n20 minus.n19 6.60088
R410 minus.n7 minus.n6 2.92171
R411 minus.n17 minus.n16 2.92171
R412 minus.n5 minus.n4 0.285035
R413 minus.n15 minus.n14 0.285035
R414 minus.n9 minus.n0 0.189894
R415 minus.n5 minus.n0 0.189894
R416 minus.n15 minus.n10 0.189894
R417 minus.n19 minus.n10 0.189894
R418 minus minus.n20 0.188
R419 drain_right.n26 drain_right.n0 289.615
R420 drain_right.n64 drain_right.n38 289.615
R421 drain_right.n11 drain_right.n10 185
R422 drain_right.n8 drain_right.n7 185
R423 drain_right.n17 drain_right.n16 185
R424 drain_right.n19 drain_right.n18 185
R425 drain_right.n4 drain_right.n3 185
R426 drain_right.n25 drain_right.n24 185
R427 drain_right.n27 drain_right.n26 185
R428 drain_right.n65 drain_right.n64 185
R429 drain_right.n63 drain_right.n62 185
R430 drain_right.n42 drain_right.n41 185
R431 drain_right.n57 drain_right.n56 185
R432 drain_right.n55 drain_right.n54 185
R433 drain_right.n46 drain_right.n45 185
R434 drain_right.n49 drain_right.n48 185
R435 drain_right.t8 drain_right.n9 147.661
R436 drain_right.t9 drain_right.n47 147.661
R437 drain_right.n10 drain_right.n7 104.615
R438 drain_right.n17 drain_right.n7 104.615
R439 drain_right.n18 drain_right.n17 104.615
R440 drain_right.n18 drain_right.n3 104.615
R441 drain_right.n25 drain_right.n3 104.615
R442 drain_right.n26 drain_right.n25 104.615
R443 drain_right.n64 drain_right.n63 104.615
R444 drain_right.n63 drain_right.n41 104.615
R445 drain_right.n56 drain_right.n41 104.615
R446 drain_right.n56 drain_right.n55 104.615
R447 drain_right.n55 drain_right.n45 104.615
R448 drain_right.n48 drain_right.n45 104.615
R449 drain_right.n37 drain_right.n35 67.9924
R450 drain_right.n34 drain_right.n33 67.7366
R451 drain_right.n37 drain_right.n36 67.1908
R452 drain_right.n32 drain_right.n31 67.1907
R453 drain_right.n10 drain_right.t8 52.3082
R454 drain_right.n48 drain_right.t9 52.3082
R455 drain_right.n32 drain_right.n30 49.6659
R456 drain_right.n69 drain_right.n68 48.8641
R457 drain_right drain_right.n34 25.6757
R458 drain_right.n11 drain_right.n9 15.6674
R459 drain_right.n49 drain_right.n47 15.6674
R460 drain_right.n12 drain_right.n8 12.8005
R461 drain_right.n50 drain_right.n46 12.8005
R462 drain_right.n16 drain_right.n15 12.0247
R463 drain_right.n54 drain_right.n53 12.0247
R464 drain_right.n19 drain_right.n6 11.249
R465 drain_right.n57 drain_right.n44 11.249
R466 drain_right.n20 drain_right.n4 10.4732
R467 drain_right.n58 drain_right.n42 10.4732
R468 drain_right.n24 drain_right.n23 9.69747
R469 drain_right.n62 drain_right.n61 9.69747
R470 drain_right.n30 drain_right.n29 9.45567
R471 drain_right.n68 drain_right.n67 9.45567
R472 drain_right.n29 drain_right.n28 9.3005
R473 drain_right.n2 drain_right.n1 9.3005
R474 drain_right.n23 drain_right.n22 9.3005
R475 drain_right.n21 drain_right.n20 9.3005
R476 drain_right.n6 drain_right.n5 9.3005
R477 drain_right.n15 drain_right.n14 9.3005
R478 drain_right.n13 drain_right.n12 9.3005
R479 drain_right.n67 drain_right.n66 9.3005
R480 drain_right.n40 drain_right.n39 9.3005
R481 drain_right.n61 drain_right.n60 9.3005
R482 drain_right.n59 drain_right.n58 9.3005
R483 drain_right.n44 drain_right.n43 9.3005
R484 drain_right.n53 drain_right.n52 9.3005
R485 drain_right.n51 drain_right.n50 9.3005
R486 drain_right.n27 drain_right.n2 8.92171
R487 drain_right.n65 drain_right.n40 8.92171
R488 drain_right.n28 drain_right.n0 8.14595
R489 drain_right.n66 drain_right.n38 8.14595
R490 drain_right drain_right.n69 6.05408
R491 drain_right.n30 drain_right.n0 5.81868
R492 drain_right.n68 drain_right.n38 5.81868
R493 drain_right.n28 drain_right.n27 5.04292
R494 drain_right.n66 drain_right.n65 5.04292
R495 drain_right.n13 drain_right.n9 4.38594
R496 drain_right.n51 drain_right.n47 4.38594
R497 drain_right.n24 drain_right.n2 4.26717
R498 drain_right.n62 drain_right.n40 4.26717
R499 drain_right.n23 drain_right.n4 3.49141
R500 drain_right.n61 drain_right.n42 3.49141
R501 drain_right.n33 drain_right.t6 3.3005
R502 drain_right.n33 drain_right.t2 3.3005
R503 drain_right.n31 drain_right.t1 3.3005
R504 drain_right.n31 drain_right.t0 3.3005
R505 drain_right.n35 drain_right.t4 3.3005
R506 drain_right.n35 drain_right.t3 3.3005
R507 drain_right.n36 drain_right.t7 3.3005
R508 drain_right.n36 drain_right.t5 3.3005
R509 drain_right.n20 drain_right.n19 2.71565
R510 drain_right.n58 drain_right.n57 2.71565
R511 drain_right.n16 drain_right.n6 1.93989
R512 drain_right.n54 drain_right.n44 1.93989
R513 drain_right.n15 drain_right.n8 1.16414
R514 drain_right.n53 drain_right.n46 1.16414
R515 drain_right.n69 drain_right.n37 0.802224
R516 drain_right.n12 drain_right.n11 0.388379
R517 drain_right.n50 drain_right.n49 0.388379
R518 drain_right.n14 drain_right.n13 0.155672
R519 drain_right.n14 drain_right.n5 0.155672
R520 drain_right.n21 drain_right.n5 0.155672
R521 drain_right.n22 drain_right.n21 0.155672
R522 drain_right.n22 drain_right.n1 0.155672
R523 drain_right.n29 drain_right.n1 0.155672
R524 drain_right.n67 drain_right.n39 0.155672
R525 drain_right.n60 drain_right.n39 0.155672
R526 drain_right.n60 drain_right.n59 0.155672
R527 drain_right.n59 drain_right.n43 0.155672
R528 drain_right.n52 drain_right.n43 0.155672
R529 drain_right.n52 drain_right.n51 0.155672
R530 drain_right.n34 drain_right.n32 0.145585
C0 source plus 3.39032f
C1 drain_left plus 3.46938f
C2 minus plus 4.31868f
C3 source drain_left 8.91432f
C4 source minus 3.37603f
C5 plus drain_right 0.333958f
C6 drain_left minus 0.172117f
C7 source drain_right 8.910769f
C8 drain_left drain_right 0.907907f
C9 minus drain_right 3.29282f
C10 drain_right a_n1832_n2088# 5.18467f
C11 drain_left a_n1832_n2088# 5.47512f
C12 source a_n1832_n2088# 4.120332f
C13 minus a_n1832_n2088# 6.659752f
C14 plus a_n1832_n2088# 8.094151f
C15 drain_right.n0 a_n1832_n2088# 0.035063f
C16 drain_right.n1 a_n1832_n2088# 0.024946f
C17 drain_right.n2 a_n1832_n2088# 0.013405f
C18 drain_right.n3 a_n1832_n2088# 0.031684f
C19 drain_right.n4 a_n1832_n2088# 0.014193f
C20 drain_right.n5 a_n1832_n2088# 0.024946f
C21 drain_right.n6 a_n1832_n2088# 0.013405f
C22 drain_right.n7 a_n1832_n2088# 0.031684f
C23 drain_right.n8 a_n1832_n2088# 0.014193f
C24 drain_right.n9 a_n1832_n2088# 0.10675f
C25 drain_right.t8 a_n1832_n2088# 0.051641f
C26 drain_right.n10 a_n1832_n2088# 0.023763f
C27 drain_right.n11 a_n1832_n2088# 0.018715f
C28 drain_right.n12 a_n1832_n2088# 0.013405f
C29 drain_right.n13 a_n1832_n2088# 0.593559f
C30 drain_right.n14 a_n1832_n2088# 0.024946f
C31 drain_right.n15 a_n1832_n2088# 0.013405f
C32 drain_right.n16 a_n1832_n2088# 0.014193f
C33 drain_right.n17 a_n1832_n2088# 0.031684f
C34 drain_right.n18 a_n1832_n2088# 0.031684f
C35 drain_right.n19 a_n1832_n2088# 0.014193f
C36 drain_right.n20 a_n1832_n2088# 0.013405f
C37 drain_right.n21 a_n1832_n2088# 0.024946f
C38 drain_right.n22 a_n1832_n2088# 0.024946f
C39 drain_right.n23 a_n1832_n2088# 0.013405f
C40 drain_right.n24 a_n1832_n2088# 0.014193f
C41 drain_right.n25 a_n1832_n2088# 0.031684f
C42 drain_right.n26 a_n1832_n2088# 0.06859f
C43 drain_right.n27 a_n1832_n2088# 0.014193f
C44 drain_right.n28 a_n1832_n2088# 0.013405f
C45 drain_right.n29 a_n1832_n2088# 0.057661f
C46 drain_right.n30 a_n1832_n2088# 0.057419f
C47 drain_right.t1 a_n1832_n2088# 0.118277f
C48 drain_right.t0 a_n1832_n2088# 0.118277f
C49 drain_right.n31 a_n1832_n2088# 0.986432f
C50 drain_right.n32 a_n1832_n2088# 0.393222f
C51 drain_right.t6 a_n1832_n2088# 0.118277f
C52 drain_right.t2 a_n1832_n2088# 0.118277f
C53 drain_right.n33 a_n1832_n2088# 0.989026f
C54 drain_right.n34 a_n1832_n2088# 1.1776f
C55 drain_right.t4 a_n1832_n2088# 0.118277f
C56 drain_right.t3 a_n1832_n2088# 0.118277f
C57 drain_right.n35 a_n1832_n2088# 0.990458f
C58 drain_right.t7 a_n1832_n2088# 0.118277f
C59 drain_right.t5 a_n1832_n2088# 0.118277f
C60 drain_right.n36 a_n1832_n2088# 0.986437f
C61 drain_right.n37 a_n1832_n2088# 0.668726f
C62 drain_right.n38 a_n1832_n2088# 0.035063f
C63 drain_right.n39 a_n1832_n2088# 0.024946f
C64 drain_right.n40 a_n1832_n2088# 0.013405f
C65 drain_right.n41 a_n1832_n2088# 0.031684f
C66 drain_right.n42 a_n1832_n2088# 0.014193f
C67 drain_right.n43 a_n1832_n2088# 0.024946f
C68 drain_right.n44 a_n1832_n2088# 0.013405f
C69 drain_right.n45 a_n1832_n2088# 0.031684f
C70 drain_right.n46 a_n1832_n2088# 0.014193f
C71 drain_right.n47 a_n1832_n2088# 0.10675f
C72 drain_right.t9 a_n1832_n2088# 0.051641f
C73 drain_right.n48 a_n1832_n2088# 0.023763f
C74 drain_right.n49 a_n1832_n2088# 0.018715f
C75 drain_right.n50 a_n1832_n2088# 0.013405f
C76 drain_right.n51 a_n1832_n2088# 0.593559f
C77 drain_right.n52 a_n1832_n2088# 0.024946f
C78 drain_right.n53 a_n1832_n2088# 0.013405f
C79 drain_right.n54 a_n1832_n2088# 0.014193f
C80 drain_right.n55 a_n1832_n2088# 0.031684f
C81 drain_right.n56 a_n1832_n2088# 0.031684f
C82 drain_right.n57 a_n1832_n2088# 0.014193f
C83 drain_right.n58 a_n1832_n2088# 0.013405f
C84 drain_right.n59 a_n1832_n2088# 0.024946f
C85 drain_right.n60 a_n1832_n2088# 0.024946f
C86 drain_right.n61 a_n1832_n2088# 0.013405f
C87 drain_right.n62 a_n1832_n2088# 0.014193f
C88 drain_right.n63 a_n1832_n2088# 0.031684f
C89 drain_right.n64 a_n1832_n2088# 0.06859f
C90 drain_right.n65 a_n1832_n2088# 0.014193f
C91 drain_right.n66 a_n1832_n2088# 0.013405f
C92 drain_right.n67 a_n1832_n2088# 0.057661f
C93 drain_right.n68 a_n1832_n2088# 0.055603f
C94 drain_right.n69 a_n1832_n2088# 0.336493f
C95 minus.n0 a_n1832_n2088# 0.045871f
C96 minus.t4 a_n1832_n2088# 0.478988f
C97 minus.n1 a_n1832_n2088# 0.233959f
C98 minus.t2 a_n1832_n2088# 0.478988f
C99 minus.t6 a_n1832_n2088# 0.496586f
C100 minus.t5 a_n1832_n2088# 0.478988f
C101 minus.n2 a_n1832_n2088# 0.233189f
C102 minus.n3 a_n1832_n2088# 0.208074f
C103 minus.n4 a_n1832_n2088# 0.221717f
C104 minus.n5 a_n1832_n2088# 0.061209f
C105 minus.n6 a_n1832_n2088# 0.224116f
C106 minus.n7 a_n1832_n2088# 0.010409f
C107 minus.t0 a_n1832_n2088# 0.478988f
C108 minus.n8 a_n1832_n2088# 0.222984f
C109 minus.n9 a_n1832_n2088# 1.30771f
C110 minus.n10 a_n1832_n2088# 0.045871f
C111 minus.t9 a_n1832_n2088# 0.478988f
C112 minus.n11 a_n1832_n2088# 0.233959f
C113 minus.t1 a_n1832_n2088# 0.496586f
C114 minus.t8 a_n1832_n2088# 0.478988f
C115 minus.n12 a_n1832_n2088# 0.233189f
C116 minus.n13 a_n1832_n2088# 0.208074f
C117 minus.n14 a_n1832_n2088# 0.221717f
C118 minus.n15 a_n1832_n2088# 0.061209f
C119 minus.t3 a_n1832_n2088# 0.478988f
C120 minus.n16 a_n1832_n2088# 0.224116f
C121 minus.n17 a_n1832_n2088# 0.010409f
C122 minus.t7 a_n1832_n2088# 0.478988f
C123 minus.n18 a_n1832_n2088# 0.222984f
C124 minus.n19 a_n1832_n2088# 0.310745f
C125 minus.n20 a_n1832_n2088# 1.60328f
C126 source.n0 a_n1832_n2088# 0.039088f
C127 source.n1 a_n1832_n2088# 0.027809f
C128 source.n2 a_n1832_n2088# 0.014943f
C129 source.n3 a_n1832_n2088# 0.035321f
C130 source.n4 a_n1832_n2088# 0.015822f
C131 source.n5 a_n1832_n2088# 0.027809f
C132 source.n6 a_n1832_n2088# 0.014943f
C133 source.n7 a_n1832_n2088# 0.035321f
C134 source.n8 a_n1832_n2088# 0.015822f
C135 source.n9 a_n1832_n2088# 0.119003f
C136 source.t17 a_n1832_n2088# 0.057568f
C137 source.n10 a_n1832_n2088# 0.02649f
C138 source.n11 a_n1832_n2088# 0.020863f
C139 source.n12 a_n1832_n2088# 0.014943f
C140 source.n13 a_n1832_n2088# 0.661687f
C141 source.n14 a_n1832_n2088# 0.027809f
C142 source.n15 a_n1832_n2088# 0.014943f
C143 source.n16 a_n1832_n2088# 0.015822f
C144 source.n17 a_n1832_n2088# 0.035321f
C145 source.n18 a_n1832_n2088# 0.035321f
C146 source.n19 a_n1832_n2088# 0.015822f
C147 source.n20 a_n1832_n2088# 0.014943f
C148 source.n21 a_n1832_n2088# 0.027809f
C149 source.n22 a_n1832_n2088# 0.027809f
C150 source.n23 a_n1832_n2088# 0.014943f
C151 source.n24 a_n1832_n2088# 0.015822f
C152 source.n25 a_n1832_n2088# 0.035321f
C153 source.n26 a_n1832_n2088# 0.076463f
C154 source.n27 a_n1832_n2088# 0.015822f
C155 source.n28 a_n1832_n2088# 0.014943f
C156 source.n29 a_n1832_n2088# 0.064279f
C157 source.n30 a_n1832_n2088# 0.042784f
C158 source.n31 a_n1832_n2088# 0.713266f
C159 source.t13 a_n1832_n2088# 0.131853f
C160 source.t14 a_n1832_n2088# 0.131853f
C161 source.n32 a_n1832_n2088# 1.02688f
C162 source.n33 a_n1832_n2088# 0.404362f
C163 source.t11 a_n1832_n2088# 0.131853f
C164 source.t12 a_n1832_n2088# 0.131853f
C165 source.n34 a_n1832_n2088# 1.02688f
C166 source.n35 a_n1832_n2088# 0.410541f
C167 source.n36 a_n1832_n2088# 0.039088f
C168 source.n37 a_n1832_n2088# 0.027809f
C169 source.n38 a_n1832_n2088# 0.014943f
C170 source.n39 a_n1832_n2088# 0.035321f
C171 source.n40 a_n1832_n2088# 0.015822f
C172 source.n41 a_n1832_n2088# 0.027809f
C173 source.n42 a_n1832_n2088# 0.014943f
C174 source.n43 a_n1832_n2088# 0.035321f
C175 source.n44 a_n1832_n2088# 0.015822f
C176 source.n45 a_n1832_n2088# 0.119003f
C177 source.t0 a_n1832_n2088# 0.057568f
C178 source.n46 a_n1832_n2088# 0.02649f
C179 source.n47 a_n1832_n2088# 0.020863f
C180 source.n48 a_n1832_n2088# 0.014943f
C181 source.n49 a_n1832_n2088# 0.661687f
C182 source.n50 a_n1832_n2088# 0.027809f
C183 source.n51 a_n1832_n2088# 0.014943f
C184 source.n52 a_n1832_n2088# 0.015822f
C185 source.n53 a_n1832_n2088# 0.035321f
C186 source.n54 a_n1832_n2088# 0.035321f
C187 source.n55 a_n1832_n2088# 0.015822f
C188 source.n56 a_n1832_n2088# 0.014943f
C189 source.n57 a_n1832_n2088# 0.027809f
C190 source.n58 a_n1832_n2088# 0.027809f
C191 source.n59 a_n1832_n2088# 0.014943f
C192 source.n60 a_n1832_n2088# 0.015822f
C193 source.n61 a_n1832_n2088# 0.035321f
C194 source.n62 a_n1832_n2088# 0.076463f
C195 source.n63 a_n1832_n2088# 0.015822f
C196 source.n64 a_n1832_n2088# 0.014943f
C197 source.n65 a_n1832_n2088# 0.064279f
C198 source.n66 a_n1832_n2088# 0.042784f
C199 source.n67 a_n1832_n2088# 0.17361f
C200 source.t8 a_n1832_n2088# 0.131853f
C201 source.t6 a_n1832_n2088# 0.131853f
C202 source.n68 a_n1832_n2088# 1.02688f
C203 source.n69 a_n1832_n2088# 0.404362f
C204 source.t5 a_n1832_n2088# 0.131853f
C205 source.t7 a_n1832_n2088# 0.131853f
C206 source.n70 a_n1832_n2088# 1.02688f
C207 source.n71 a_n1832_n2088# 1.38672f
C208 source.t10 a_n1832_n2088# 0.131853f
C209 source.t15 a_n1832_n2088# 0.131853f
C210 source.n72 a_n1832_n2088# 1.02687f
C211 source.n73 a_n1832_n2088# 1.38673f
C212 source.t18 a_n1832_n2088# 0.131853f
C213 source.t19 a_n1832_n2088# 0.131853f
C214 source.n74 a_n1832_n2088# 1.02687f
C215 source.n75 a_n1832_n2088# 0.404369f
C216 source.n76 a_n1832_n2088# 0.039088f
C217 source.n77 a_n1832_n2088# 0.027809f
C218 source.n78 a_n1832_n2088# 0.014943f
C219 source.n79 a_n1832_n2088# 0.035321f
C220 source.n80 a_n1832_n2088# 0.015822f
C221 source.n81 a_n1832_n2088# 0.027809f
C222 source.n82 a_n1832_n2088# 0.014943f
C223 source.n83 a_n1832_n2088# 0.035321f
C224 source.n84 a_n1832_n2088# 0.015822f
C225 source.n85 a_n1832_n2088# 0.119003f
C226 source.t16 a_n1832_n2088# 0.057568f
C227 source.n86 a_n1832_n2088# 0.02649f
C228 source.n87 a_n1832_n2088# 0.020863f
C229 source.n88 a_n1832_n2088# 0.014943f
C230 source.n89 a_n1832_n2088# 0.661687f
C231 source.n90 a_n1832_n2088# 0.027809f
C232 source.n91 a_n1832_n2088# 0.014943f
C233 source.n92 a_n1832_n2088# 0.015822f
C234 source.n93 a_n1832_n2088# 0.035321f
C235 source.n94 a_n1832_n2088# 0.035321f
C236 source.n95 a_n1832_n2088# 0.015822f
C237 source.n96 a_n1832_n2088# 0.014943f
C238 source.n97 a_n1832_n2088# 0.027809f
C239 source.n98 a_n1832_n2088# 0.027809f
C240 source.n99 a_n1832_n2088# 0.014943f
C241 source.n100 a_n1832_n2088# 0.015822f
C242 source.n101 a_n1832_n2088# 0.035321f
C243 source.n102 a_n1832_n2088# 0.076463f
C244 source.n103 a_n1832_n2088# 0.015822f
C245 source.n104 a_n1832_n2088# 0.014943f
C246 source.n105 a_n1832_n2088# 0.064279f
C247 source.n106 a_n1832_n2088# 0.042784f
C248 source.n107 a_n1832_n2088# 0.17361f
C249 source.t1 a_n1832_n2088# 0.131853f
C250 source.t2 a_n1832_n2088# 0.131853f
C251 source.n108 a_n1832_n2088# 1.02687f
C252 source.n109 a_n1832_n2088# 0.410548f
C253 source.t4 a_n1832_n2088# 0.131853f
C254 source.t3 a_n1832_n2088# 0.131853f
C255 source.n110 a_n1832_n2088# 1.02687f
C256 source.n111 a_n1832_n2088# 0.404369f
C257 source.n112 a_n1832_n2088# 0.039088f
C258 source.n113 a_n1832_n2088# 0.027809f
C259 source.n114 a_n1832_n2088# 0.014943f
C260 source.n115 a_n1832_n2088# 0.035321f
C261 source.n116 a_n1832_n2088# 0.015822f
C262 source.n117 a_n1832_n2088# 0.027809f
C263 source.n118 a_n1832_n2088# 0.014943f
C264 source.n119 a_n1832_n2088# 0.035321f
C265 source.n120 a_n1832_n2088# 0.015822f
C266 source.n121 a_n1832_n2088# 0.119003f
C267 source.t9 a_n1832_n2088# 0.057568f
C268 source.n122 a_n1832_n2088# 0.02649f
C269 source.n123 a_n1832_n2088# 0.020863f
C270 source.n124 a_n1832_n2088# 0.014943f
C271 source.n125 a_n1832_n2088# 0.661687f
C272 source.n126 a_n1832_n2088# 0.027809f
C273 source.n127 a_n1832_n2088# 0.014943f
C274 source.n128 a_n1832_n2088# 0.015822f
C275 source.n129 a_n1832_n2088# 0.035321f
C276 source.n130 a_n1832_n2088# 0.035321f
C277 source.n131 a_n1832_n2088# 0.015822f
C278 source.n132 a_n1832_n2088# 0.014943f
C279 source.n133 a_n1832_n2088# 0.027809f
C280 source.n134 a_n1832_n2088# 0.027809f
C281 source.n135 a_n1832_n2088# 0.014943f
C282 source.n136 a_n1832_n2088# 0.015822f
C283 source.n137 a_n1832_n2088# 0.035321f
C284 source.n138 a_n1832_n2088# 0.076463f
C285 source.n139 a_n1832_n2088# 0.015822f
C286 source.n140 a_n1832_n2088# 0.014943f
C287 source.n141 a_n1832_n2088# 0.064279f
C288 source.n142 a_n1832_n2088# 0.042784f
C289 source.n143 a_n1832_n2088# 0.313036f
C290 source.n144 a_n1832_n2088# 1.14937f
C291 drain_left.n0 a_n1832_n2088# 0.035355f
C292 drain_left.n1 a_n1832_n2088# 0.025154f
C293 drain_left.n2 a_n1832_n2088# 0.013516f
C294 drain_left.n3 a_n1832_n2088# 0.031948f
C295 drain_left.n4 a_n1832_n2088# 0.014311f
C296 drain_left.n5 a_n1832_n2088# 0.025154f
C297 drain_left.n6 a_n1832_n2088# 0.013516f
C298 drain_left.n7 a_n1832_n2088# 0.031948f
C299 drain_left.n8 a_n1832_n2088# 0.014311f
C300 drain_left.n9 a_n1832_n2088# 0.107639f
C301 drain_left.t9 a_n1832_n2088# 0.052071f
C302 drain_left.n10 a_n1832_n2088# 0.023961f
C303 drain_left.n11 a_n1832_n2088# 0.018871f
C304 drain_left.n12 a_n1832_n2088# 0.013516f
C305 drain_left.n13 a_n1832_n2088# 0.598502f
C306 drain_left.n14 a_n1832_n2088# 0.025154f
C307 drain_left.n15 a_n1832_n2088# 0.013516f
C308 drain_left.n16 a_n1832_n2088# 0.014311f
C309 drain_left.n17 a_n1832_n2088# 0.031948f
C310 drain_left.n18 a_n1832_n2088# 0.031948f
C311 drain_left.n19 a_n1832_n2088# 0.014311f
C312 drain_left.n20 a_n1832_n2088# 0.013516f
C313 drain_left.n21 a_n1832_n2088# 0.025154f
C314 drain_left.n22 a_n1832_n2088# 0.025154f
C315 drain_left.n23 a_n1832_n2088# 0.013516f
C316 drain_left.n24 a_n1832_n2088# 0.014311f
C317 drain_left.n25 a_n1832_n2088# 0.031948f
C318 drain_left.n26 a_n1832_n2088# 0.069162f
C319 drain_left.n27 a_n1832_n2088# 0.014311f
C320 drain_left.n28 a_n1832_n2088# 0.013516f
C321 drain_left.n29 a_n1832_n2088# 0.058141f
C322 drain_left.n30 a_n1832_n2088# 0.057897f
C323 drain_left.t2 a_n1832_n2088# 0.119262f
C324 drain_left.t4 a_n1832_n2088# 0.119262f
C325 drain_left.n31 a_n1832_n2088# 0.994647f
C326 drain_left.n32 a_n1832_n2088# 0.396496f
C327 drain_left.t7 a_n1832_n2088# 0.119262f
C328 drain_left.t5 a_n1832_n2088# 0.119262f
C329 drain_left.n33 a_n1832_n2088# 0.997263f
C330 drain_left.n34 a_n1832_n2088# 1.23848f
C331 drain_left.n35 a_n1832_n2088# 0.035355f
C332 drain_left.n36 a_n1832_n2088# 0.025154f
C333 drain_left.n37 a_n1832_n2088# 0.013516f
C334 drain_left.n38 a_n1832_n2088# 0.031948f
C335 drain_left.n39 a_n1832_n2088# 0.014311f
C336 drain_left.n40 a_n1832_n2088# 0.025154f
C337 drain_left.n41 a_n1832_n2088# 0.013516f
C338 drain_left.n42 a_n1832_n2088# 0.031948f
C339 drain_left.n43 a_n1832_n2088# 0.014311f
C340 drain_left.n44 a_n1832_n2088# 0.107639f
C341 drain_left.t1 a_n1832_n2088# 0.052071f
C342 drain_left.n45 a_n1832_n2088# 0.023961f
C343 drain_left.n46 a_n1832_n2088# 0.018871f
C344 drain_left.n47 a_n1832_n2088# 0.013516f
C345 drain_left.n48 a_n1832_n2088# 0.598502f
C346 drain_left.n49 a_n1832_n2088# 0.025154f
C347 drain_left.n50 a_n1832_n2088# 0.013516f
C348 drain_left.n51 a_n1832_n2088# 0.014311f
C349 drain_left.n52 a_n1832_n2088# 0.031948f
C350 drain_left.n53 a_n1832_n2088# 0.031948f
C351 drain_left.n54 a_n1832_n2088# 0.014311f
C352 drain_left.n55 a_n1832_n2088# 0.013516f
C353 drain_left.n56 a_n1832_n2088# 0.025154f
C354 drain_left.n57 a_n1832_n2088# 0.025154f
C355 drain_left.n58 a_n1832_n2088# 0.013516f
C356 drain_left.n59 a_n1832_n2088# 0.014311f
C357 drain_left.n60 a_n1832_n2088# 0.031948f
C358 drain_left.n61 a_n1832_n2088# 0.069162f
C359 drain_left.n62 a_n1832_n2088# 0.014311f
C360 drain_left.n63 a_n1832_n2088# 0.013516f
C361 drain_left.n64 a_n1832_n2088# 0.058141f
C362 drain_left.n65 a_n1832_n2088# 0.057897f
C363 drain_left.t3 a_n1832_n2088# 0.119262f
C364 drain_left.t8 a_n1832_n2088# 0.119262f
C365 drain_left.n66 a_n1832_n2088# 0.994652f
C366 drain_left.n67 a_n1832_n2088# 0.445693f
C367 drain_left.t6 a_n1832_n2088# 0.119262f
C368 drain_left.t0 a_n1832_n2088# 0.119262f
C369 drain_left.n68 a_n1832_n2088# 0.994647f
C370 drain_left.n69 a_n1832_n2088# 0.55345f
C371 plus.n0 a_n1832_n2088# 0.047103f
C372 plus.t2 a_n1832_n2088# 0.491845f
C373 plus.t5 a_n1832_n2088# 0.491845f
C374 plus.n1 a_n1832_n2088# 0.062853f
C375 plus.t6 a_n1832_n2088# 0.491845f
C376 plus.n2 a_n1832_n2088# 0.227668f
C377 plus.t7 a_n1832_n2088# 0.491845f
C378 plus.t8 a_n1832_n2088# 0.509915f
C379 plus.n3 a_n1832_n2088# 0.213659f
C380 plus.n4 a_n1832_n2088# 0.239448f
C381 plus.n5 a_n1832_n2088# 0.240239f
C382 plus.n6 a_n1832_n2088# 0.230131f
C383 plus.n7 a_n1832_n2088# 0.010689f
C384 plus.n8 a_n1832_n2088# 0.228969f
C385 plus.n9 a_n1832_n2088# 0.415256f
C386 plus.n10 a_n1832_n2088# 0.047103f
C387 plus.t9 a_n1832_n2088# 0.491845f
C388 plus.n11 a_n1832_n2088# 0.062853f
C389 plus.t4 a_n1832_n2088# 0.491845f
C390 plus.n12 a_n1832_n2088# 0.227668f
C391 plus.t1 a_n1832_n2088# 0.491845f
C392 plus.t3 a_n1832_n2088# 0.509915f
C393 plus.n13 a_n1832_n2088# 0.213659f
C394 plus.t0 a_n1832_n2088# 0.491845f
C395 plus.n14 a_n1832_n2088# 0.239448f
C396 plus.n15 a_n1832_n2088# 0.240239f
C397 plus.n16 a_n1832_n2088# 0.230131f
C398 plus.n17 a_n1832_n2088# 0.010689f
C399 plus.n18 a_n1832_n2088# 0.228969f
C400 plus.n19 a_n1832_n2088# 1.214f
.ends

