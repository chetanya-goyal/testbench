* NGSPICE file created from diffpair660.ext - technology: sky130A

.subckt diffpair660 minus drain_right drain_left source plus
X0 drain_right minus source a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.25
X1 a_n948_n5892# a_n948_n5892# a_n948_n5892# a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.25
X2 a_n948_n5892# a_n948_n5892# a_n948_n5892# a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
X3 drain_left plus source a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.25
X4 drain_right minus source a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.25
X5 a_n948_n5892# a_n948_n5892# a_n948_n5892# a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
X6 drain_left plus source a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=9.75 ps=50.78 w=25 l=0.25
X7 a_n948_n5892# a_n948_n5892# a_n948_n5892# a_n948_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
.ends

