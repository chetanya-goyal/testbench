* NGSPICE file created from diffpair519.ext - technology: sky130A

.subckt diffpair519 minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t13 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X1 drain_left.t12 plus.t1 source.t46 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X2 source.t12 minus.t0 drain_right.t23 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X3 drain_left.t17 plus.t2 source.t45 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X4 drain_left.t16 plus.t3 source.t44 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X5 drain_right.t22 minus.t1 source.t5 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X6 drain_right.t21 minus.t2 source.t14 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X7 source.t6 minus.t3 drain_right.t20 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X8 source.t43 plus.t4 drain_left.t23 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X9 source.t19 minus.t4 drain_right.t19 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X10 source.t23 minus.t5 drain_right.t18 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X11 drain_left.t22 plus.t5 source.t42 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X12 drain_right.t17 minus.t6 source.t13 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X13 drain_right.t16 minus.t7 source.t0 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X14 source.t41 plus.t6 drain_left.t19 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X15 a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X16 drain_right.t15 minus.t8 source.t4 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 drain_left.t18 plus.t7 source.t40 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X18 source.t9 minus.t9 drain_right.t14 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X19 drain_left.t1 plus.t8 source.t39 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X20 drain_left.t0 plus.t9 source.t38 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X21 source.t37 plus.t10 drain_left.t15 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X22 drain_left.t14 plus.t11 source.t36 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 source.t16 minus.t10 drain_right.t13 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X24 source.t21 minus.t11 drain_right.t12 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X25 source.t1 minus.t12 drain_right.t11 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X26 source.t35 plus.t12 drain_left.t5 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X27 a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X28 drain_right.t10 minus.t13 source.t8 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X29 drain_left.t4 plus.t13 source.t34 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X30 source.t10 minus.t14 drain_right.t9 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X31 drain_left.t7 plus.t14 source.t33 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X32 source.t32 plus.t15 drain_left.t6 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X33 source.t31 plus.t16 drain_left.t9 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X34 source.t30 plus.t17 drain_left.t8 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X35 source.t29 plus.t18 drain_left.t3 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X36 drain_left.t2 plus.t19 source.t28 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X37 drain_right.t8 minus.t15 source.t15 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X38 drain_right.t7 minus.t16 source.t20 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X39 a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X40 drain_right.t6 minus.t17 source.t11 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X41 drain_right.t5 minus.t18 source.t18 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X42 source.t17 minus.t19 drain_right.t4 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X43 source.t22 minus.t20 drain_right.t3 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X44 source.t3 minus.t21 drain_right.t2 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X45 source.t27 plus.t20 drain_left.t11 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X46 a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X47 drain_right.t1 minus.t22 source.t7 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X48 drain_right.t0 minus.t23 source.t2 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X49 source.t26 plus.t21 drain_left.t10 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X50 source.t25 plus.t22 drain_left.t21 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X51 drain_left.t20 plus.t23 source.t24 a_n2354_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 plus.n9 plus.t4 1340.84
R1 plus.n35 plus.t5 1340.84
R2 plus.n46 plus.t2 1340.84
R3 plus.n72 plus.t6 1340.84
R4 plus.n8 plus.t11 1309.43
R5 plus.n13 plus.t16 1309.43
R6 plus.n15 plus.t23 1309.43
R7 plus.n5 plus.t10 1309.43
R8 plus.n20 plus.t13 1309.43
R9 plus.n3 plus.t20 1309.43
R10 plus.n26 plus.t1 1309.43
R11 plus.n28 plus.t12 1309.43
R12 plus.n1 plus.t19 1309.43
R13 plus.n34 plus.t0 1309.43
R14 plus.n45 plus.t15 1309.43
R15 plus.n50 plus.t3 1309.43
R16 plus.n52 plus.t17 1309.43
R17 plus.n42 plus.t8 1309.43
R18 plus.n57 plus.t18 1309.43
R19 plus.n40 plus.t9 1309.43
R20 plus.n63 plus.t21 1309.43
R21 plus.n65 plus.t7 1309.43
R22 plus.n38 plus.t22 1309.43
R23 plus.n71 plus.t14 1309.43
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 33.0255
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus plus.n36 13.2505
R88 plus.n8 plus.n7 12.4157
R89 plus.n34 plus.n33 12.4157
R90 plus.n71 plus.n70 12.4157
R91 plus.n45 plus.n44 12.4157
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 drain_left.n13 drain_left.n11 61.4229
R125 drain_left.n7 drain_left.n5 61.4227
R126 drain_left.n2 drain_left.n0 61.4227
R127 drain_left.n19 drain_left.n18 60.8798
R128 drain_left.n17 drain_left.n16 60.8798
R129 drain_left.n15 drain_left.n14 60.8798
R130 drain_left.n13 drain_left.n12 60.8798
R131 drain_left.n21 drain_left.n20 60.8796
R132 drain_left.n7 drain_left.n6 60.8796
R133 drain_left.n9 drain_left.n8 60.8796
R134 drain_left.n4 drain_left.n3 60.8796
R135 drain_left.n2 drain_left.n1 60.8796
R136 drain_left drain_left.n10 34.7993
R137 drain_left drain_left.n21 6.19632
R138 drain_left.n5 drain_left.t6 1.3205
R139 drain_left.n5 drain_left.t17 1.3205
R140 drain_left.n6 drain_left.t8 1.3205
R141 drain_left.n6 drain_left.t16 1.3205
R142 drain_left.n8 drain_left.t3 1.3205
R143 drain_left.n8 drain_left.t1 1.3205
R144 drain_left.n3 drain_left.t10 1.3205
R145 drain_left.n3 drain_left.t0 1.3205
R146 drain_left.n1 drain_left.t21 1.3205
R147 drain_left.n1 drain_left.t18 1.3205
R148 drain_left.n0 drain_left.t19 1.3205
R149 drain_left.n0 drain_left.t7 1.3205
R150 drain_left.n20 drain_left.t13 1.3205
R151 drain_left.n20 drain_left.t22 1.3205
R152 drain_left.n18 drain_left.t5 1.3205
R153 drain_left.n18 drain_left.t2 1.3205
R154 drain_left.n16 drain_left.t11 1.3205
R155 drain_left.n16 drain_left.t12 1.3205
R156 drain_left.n14 drain_left.t15 1.3205
R157 drain_left.n14 drain_left.t4 1.3205
R158 drain_left.n12 drain_left.t9 1.3205
R159 drain_left.n12 drain_left.t20 1.3205
R160 drain_left.n11 drain_left.t23 1.3205
R161 drain_left.n11 drain_left.t14 1.3205
R162 drain_left.n9 drain_left.n7 0.543603
R163 drain_left.n4 drain_left.n2 0.543603
R164 drain_left.n15 drain_left.n13 0.543603
R165 drain_left.n17 drain_left.n15 0.543603
R166 drain_left.n19 drain_left.n17 0.543603
R167 drain_left.n21 drain_left.n19 0.543603
R168 drain_left.n10 drain_left.n9 0.216706
R169 drain_left.n10 drain_left.n4 0.216706
R170 source.n11 source.t43 45.521
R171 source.n12 source.t8 45.521
R172 source.n23 source.t6 45.521
R173 source.n47 source.t13 45.5208
R174 source.n36 source.t23 45.5208
R175 source.n35 source.t45 45.5208
R176 source.n24 source.t41 45.5208
R177 source.n0 source.t42 45.5208
R178 source.n2 source.n1 44.201
R179 source.n4 source.n3 44.201
R180 source.n6 source.n5 44.201
R181 source.n8 source.n7 44.201
R182 source.n10 source.n9 44.201
R183 source.n14 source.n13 44.201
R184 source.n16 source.n15 44.201
R185 source.n18 source.n17 44.201
R186 source.n20 source.n19 44.201
R187 source.n22 source.n21 44.201
R188 source.n46 source.n45 44.2008
R189 source.n44 source.n43 44.2008
R190 source.n42 source.n41 44.2008
R191 source.n40 source.n39 44.2008
R192 source.n38 source.n37 44.2008
R193 source.n34 source.n33 44.2008
R194 source.n32 source.n31 44.2008
R195 source.n30 source.n29 44.2008
R196 source.n28 source.n27 44.2008
R197 source.n26 source.n25 44.2008
R198 source.n24 source.n23 24.1036
R199 source.n48 source.n0 18.5691
R200 source.n48 source.n47 5.53498
R201 source.n45 source.t0 1.3205
R202 source.n45 source.t10 1.3205
R203 source.n43 source.t7 1.3205
R204 source.n43 source.t3 1.3205
R205 source.n41 source.t2 1.3205
R206 source.n41 source.t21 1.3205
R207 source.n39 source.t11 1.3205
R208 source.n39 source.t1 1.3205
R209 source.n37 source.t18 1.3205
R210 source.n37 source.t19 1.3205
R211 source.n33 source.t44 1.3205
R212 source.n33 source.t32 1.3205
R213 source.n31 source.t39 1.3205
R214 source.n31 source.t30 1.3205
R215 source.n29 source.t38 1.3205
R216 source.n29 source.t29 1.3205
R217 source.n27 source.t40 1.3205
R218 source.n27 source.t26 1.3205
R219 source.n25 source.t33 1.3205
R220 source.n25 source.t25 1.3205
R221 source.n1 source.t28 1.3205
R222 source.n1 source.t47 1.3205
R223 source.n3 source.t46 1.3205
R224 source.n3 source.t35 1.3205
R225 source.n5 source.t34 1.3205
R226 source.n5 source.t27 1.3205
R227 source.n7 source.t24 1.3205
R228 source.n7 source.t37 1.3205
R229 source.n9 source.t36 1.3205
R230 source.n9 source.t31 1.3205
R231 source.n13 source.t5 1.3205
R232 source.n13 source.t17 1.3205
R233 source.n15 source.t15 1.3205
R234 source.n15 source.t16 1.3205
R235 source.n17 source.t4 1.3205
R236 source.n17 source.t12 1.3205
R237 source.n19 source.t14 1.3205
R238 source.n19 source.t22 1.3205
R239 source.n21 source.t20 1.3205
R240 source.n21 source.t9 1.3205
R241 source.n23 source.n22 0.543603
R242 source.n22 source.n20 0.543603
R243 source.n20 source.n18 0.543603
R244 source.n18 source.n16 0.543603
R245 source.n16 source.n14 0.543603
R246 source.n14 source.n12 0.543603
R247 source.n11 source.n10 0.543603
R248 source.n10 source.n8 0.543603
R249 source.n8 source.n6 0.543603
R250 source.n6 source.n4 0.543603
R251 source.n4 source.n2 0.543603
R252 source.n2 source.n0 0.543603
R253 source.n26 source.n24 0.543603
R254 source.n28 source.n26 0.543603
R255 source.n30 source.n28 0.543603
R256 source.n32 source.n30 0.543603
R257 source.n34 source.n32 0.543603
R258 source.n35 source.n34 0.543603
R259 source.n38 source.n36 0.543603
R260 source.n40 source.n38 0.543603
R261 source.n42 source.n40 0.543603
R262 source.n44 source.n42 0.543603
R263 source.n46 source.n44 0.543603
R264 source.n47 source.n46 0.543603
R265 source.n12 source.n11 0.470328
R266 source.n36 source.n35 0.470328
R267 source source.n48 0.188
R268 minus.n35 minus.t3 1340.84
R269 minus.n9 minus.t13 1340.84
R270 minus.n72 minus.t6 1340.84
R271 minus.n46 minus.t5 1340.84
R272 minus.n34 minus.t16 1309.43
R273 minus.n1 minus.t9 1309.43
R274 minus.n28 minus.t2 1309.43
R275 minus.n26 minus.t20 1309.43
R276 minus.n3 minus.t8 1309.43
R277 minus.n20 minus.t0 1309.43
R278 minus.n5 minus.t15 1309.43
R279 minus.n15 minus.t10 1309.43
R280 minus.n13 minus.t1 1309.43
R281 minus.n8 minus.t19 1309.43
R282 minus.n71 minus.t14 1309.43
R283 minus.n38 minus.t7 1309.43
R284 minus.n65 minus.t21 1309.43
R285 minus.n63 minus.t22 1309.43
R286 minus.n40 minus.t11 1309.43
R287 minus.n57 minus.t23 1309.43
R288 minus.n42 minus.t12 1309.43
R289 minus.n52 minus.t17 1309.43
R290 minus.n50 minus.t4 1309.43
R291 minus.n45 minus.t18 1309.43
R292 minus.n10 minus.n9 161.489
R293 minus.n47 minus.n46 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n32 minus.n31 161.3
R297 minus.n30 minus.n29 161.3
R298 minus.n27 minus.n2 161.3
R299 minus.n25 minus.n24 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n19 minus.n18 161.3
R303 minus.n17 minus.n16 161.3
R304 minus.n14 minus.n6 161.3
R305 minus.n12 minus.n11 161.3
R306 minus.n10 minus.n7 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n69 minus.n68 161.3
R310 minus.n67 minus.n66 161.3
R311 minus.n64 minus.n39 161.3
R312 minus.n62 minus.n61 161.3
R313 minus.n60 minus.n59 161.3
R314 minus.n58 minus.n41 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n54 minus.n53 161.3
R317 minus.n51 minus.n43 161.3
R318 minus.n49 minus.n48 161.3
R319 minus.n47 minus.n44 161.3
R320 minus.n33 minus.n32 73.0308
R321 minus.n22 minus.n21 73.0308
R322 minus.n12 minus.n7 73.0308
R323 minus.n49 minus.n44 73.0308
R324 minus.n59 minus.n58 73.0308
R325 minus.n70 minus.n69 73.0308
R326 minus.n29 minus.n1 66.4581
R327 minus.n14 minus.n13 66.4581
R328 minus.n51 minus.n50 66.4581
R329 minus.n66 minus.n38 66.4581
R330 minus.n25 minus.n3 63.5369
R331 minus.n20 minus.n19 63.5369
R332 minus.n57 minus.n56 63.5369
R333 minus.n62 minus.n40 63.5369
R334 minus.n35 minus.n34 60.6157
R335 minus.n9 minus.n8 60.6157
R336 minus.n46 minus.n45 60.6157
R337 minus.n72 minus.n71 60.6157
R338 minus.n28 minus.n27 47.4702
R339 minus.n16 minus.n15 47.4702
R340 minus.n53 minus.n52 47.4702
R341 minus.n65 minus.n64 47.4702
R342 minus.n27 minus.n26 44.549
R343 minus.n16 minus.n5 44.549
R344 minus.n53 minus.n42 44.549
R345 minus.n64 minus.n63 44.549
R346 minus.n74 minus.n36 40.2808
R347 minus.n26 minus.n25 28.4823
R348 minus.n19 minus.n5 28.4823
R349 minus.n56 minus.n42 28.4823
R350 minus.n63 minus.n62 28.4823
R351 minus.n29 minus.n28 25.5611
R352 minus.n15 minus.n14 25.5611
R353 minus.n52 minus.n51 25.5611
R354 minus.n66 minus.n65 25.5611
R355 minus.n34 minus.n33 12.4157
R356 minus.n8 minus.n7 12.4157
R357 minus.n45 minus.n44 12.4157
R358 minus.n71 minus.n70 12.4157
R359 minus.n22 minus.n3 9.49444
R360 minus.n21 minus.n20 9.49444
R361 minus.n58 minus.n57 9.49444
R362 minus.n59 minus.n40 9.49444
R363 minus.n32 minus.n1 6.57323
R364 minus.n13 minus.n12 6.57323
R365 minus.n50 minus.n49 6.57323
R366 minus.n69 minus.n38 6.57323
R367 minus.n74 minus.n73 6.4702
R368 minus.n36 minus.n0 0.189894
R369 minus.n31 minus.n0 0.189894
R370 minus.n31 minus.n30 0.189894
R371 minus.n30 minus.n2 0.189894
R372 minus.n24 minus.n2 0.189894
R373 minus.n24 minus.n23 0.189894
R374 minus.n23 minus.n4 0.189894
R375 minus.n18 minus.n4 0.189894
R376 minus.n18 minus.n17 0.189894
R377 minus.n17 minus.n6 0.189894
R378 minus.n11 minus.n6 0.189894
R379 minus.n11 minus.n10 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n48 minus.n43 0.189894
R382 minus.n54 minus.n43 0.189894
R383 minus.n55 minus.n54 0.189894
R384 minus.n55 minus.n41 0.189894
R385 minus.n60 minus.n41 0.189894
R386 minus.n61 minus.n60 0.189894
R387 minus.n61 minus.n39 0.189894
R388 minus.n67 minus.n39 0.189894
R389 minus.n68 minus.n67 0.189894
R390 minus.n68 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 61.4227
R394 drain_right.n7 drain_right.n5 61.4227
R395 drain_right.n2 drain_right.n0 61.4227
R396 drain_right.n13 drain_right.n12 60.8798
R397 drain_right.n15 drain_right.n14 60.8798
R398 drain_right.n17 drain_right.n16 60.8798
R399 drain_right.n19 drain_right.n18 60.8798
R400 drain_right.n21 drain_right.n20 60.8798
R401 drain_right.n7 drain_right.n6 60.8796
R402 drain_right.n9 drain_right.n8 60.8796
R403 drain_right.n4 drain_right.n3 60.8796
R404 drain_right.n2 drain_right.n1 60.8796
R405 drain_right drain_right.n10 34.2461
R406 drain_right drain_right.n21 6.19632
R407 drain_right.n5 drain_right.t9 1.3205
R408 drain_right.n5 drain_right.t17 1.3205
R409 drain_right.n6 drain_right.t2 1.3205
R410 drain_right.n6 drain_right.t16 1.3205
R411 drain_right.n8 drain_right.t12 1.3205
R412 drain_right.n8 drain_right.t1 1.3205
R413 drain_right.n3 drain_right.t11 1.3205
R414 drain_right.n3 drain_right.t0 1.3205
R415 drain_right.n1 drain_right.t19 1.3205
R416 drain_right.n1 drain_right.t6 1.3205
R417 drain_right.n0 drain_right.t18 1.3205
R418 drain_right.n0 drain_right.t5 1.3205
R419 drain_right.n11 drain_right.t4 1.3205
R420 drain_right.n11 drain_right.t10 1.3205
R421 drain_right.n12 drain_right.t13 1.3205
R422 drain_right.n12 drain_right.t22 1.3205
R423 drain_right.n14 drain_right.t23 1.3205
R424 drain_right.n14 drain_right.t8 1.3205
R425 drain_right.n16 drain_right.t3 1.3205
R426 drain_right.n16 drain_right.t15 1.3205
R427 drain_right.n18 drain_right.t14 1.3205
R428 drain_right.n18 drain_right.t21 1.3205
R429 drain_right.n20 drain_right.t20 1.3205
R430 drain_right.n20 drain_right.t7 1.3205
R431 drain_right.n9 drain_right.n7 0.543603
R432 drain_right.n4 drain_right.n2 0.543603
R433 drain_right.n21 drain_right.n19 0.543603
R434 drain_right.n19 drain_right.n17 0.543603
R435 drain_right.n17 drain_right.n15 0.543603
R436 drain_right.n15 drain_right.n13 0.543603
R437 drain_right.n10 drain_right.n9 0.216706
R438 drain_right.n10 drain_right.n4 0.216706
C0 drain_left drain_right 1.26597f
C1 plus minus 6.64957f
C2 drain_left minus 0.172624f
C3 drain_right minus 10.378f
C4 plus source 10.086599f
C5 drain_left source 54.584f
C6 drain_right source 54.584602f
C7 minus source 10.072599f
C8 drain_left plus 10.6102f
C9 plus drain_right 0.387992f
C10 drain_right a_n2354_n3888# 8.0035f
C11 drain_left a_n2354_n3888# 8.35359f
C12 source a_n2354_n3888# 10.519634f
C13 minus a_n2354_n3888# 9.480506f
C14 plus a_n2354_n3888# 11.721519f
C15 drain_right.t18 a_n2354_n3888# 0.407378f
C16 drain_right.t5 a_n2354_n3888# 0.407378f
C17 drain_right.n0 a_n2354_n3888# 3.6859f
C18 drain_right.t19 a_n2354_n3888# 0.407378f
C19 drain_right.t6 a_n2354_n3888# 0.407378f
C20 drain_right.n1 a_n2354_n3888# 3.68222f
C21 drain_right.n2 a_n2354_n3888# 0.813731f
C22 drain_right.t11 a_n2354_n3888# 0.407378f
C23 drain_right.t0 a_n2354_n3888# 0.407378f
C24 drain_right.n3 a_n2354_n3888# 3.68222f
C25 drain_right.n4 a_n2354_n3888# 0.369266f
C26 drain_right.t9 a_n2354_n3888# 0.407378f
C27 drain_right.t17 a_n2354_n3888# 0.407378f
C28 drain_right.n5 a_n2354_n3888# 3.6859f
C29 drain_right.t2 a_n2354_n3888# 0.407378f
C30 drain_right.t16 a_n2354_n3888# 0.407378f
C31 drain_right.n6 a_n2354_n3888# 3.68222f
C32 drain_right.n7 a_n2354_n3888# 0.813731f
C33 drain_right.t12 a_n2354_n3888# 0.407378f
C34 drain_right.t1 a_n2354_n3888# 0.407378f
C35 drain_right.n8 a_n2354_n3888# 3.68222f
C36 drain_right.n9 a_n2354_n3888# 0.369266f
C37 drain_right.n10 a_n2354_n3888# 2.03894f
C38 drain_right.t4 a_n2354_n3888# 0.407378f
C39 drain_right.t10 a_n2354_n3888# 0.407378f
C40 drain_right.n11 a_n2354_n3888# 3.68589f
C41 drain_right.t13 a_n2354_n3888# 0.407378f
C42 drain_right.t22 a_n2354_n3888# 0.407378f
C43 drain_right.n12 a_n2354_n3888# 3.68223f
C44 drain_right.n13 a_n2354_n3888# 0.813738f
C45 drain_right.t23 a_n2354_n3888# 0.407378f
C46 drain_right.t8 a_n2354_n3888# 0.407378f
C47 drain_right.n14 a_n2354_n3888# 3.68223f
C48 drain_right.n15 a_n2354_n3888# 0.401779f
C49 drain_right.t3 a_n2354_n3888# 0.407378f
C50 drain_right.t15 a_n2354_n3888# 0.407378f
C51 drain_right.n16 a_n2354_n3888# 3.68223f
C52 drain_right.n17 a_n2354_n3888# 0.401779f
C53 drain_right.t14 a_n2354_n3888# 0.407378f
C54 drain_right.t21 a_n2354_n3888# 0.407378f
C55 drain_right.n18 a_n2354_n3888# 3.68223f
C56 drain_right.n19 a_n2354_n3888# 0.401779f
C57 drain_right.t20 a_n2354_n3888# 0.407378f
C58 drain_right.t7 a_n2354_n3888# 0.407378f
C59 drain_right.n20 a_n2354_n3888# 3.68223f
C60 drain_right.n21 a_n2354_n3888# 0.687844f
C61 minus.n0 a_n2354_n3888# 0.048587f
C62 minus.t3 a_n2354_n3888# 0.622383f
C63 minus.t16 a_n2354_n3888# 0.616823f
C64 minus.t9 a_n2354_n3888# 0.616823f
C65 minus.n1 a_n2354_n3888# 0.236925f
C66 minus.n2 a_n2354_n3888# 0.048587f
C67 minus.t2 a_n2354_n3888# 0.616823f
C68 minus.t20 a_n2354_n3888# 0.616823f
C69 minus.t8 a_n2354_n3888# 0.616823f
C70 minus.n3 a_n2354_n3888# 0.236925f
C71 minus.n4 a_n2354_n3888# 0.048587f
C72 minus.t0 a_n2354_n3888# 0.616823f
C73 minus.t15 a_n2354_n3888# 0.616823f
C74 minus.n5 a_n2354_n3888# 0.236925f
C75 minus.n6 a_n2354_n3888# 0.048587f
C76 minus.t10 a_n2354_n3888# 0.616823f
C77 minus.t1 a_n2354_n3888# 0.616823f
C78 minus.n7 a_n2354_n3888# 0.018664f
C79 minus.t19 a_n2354_n3888# 0.616823f
C80 minus.n8 a_n2354_n3888# 0.236925f
C81 minus.t13 a_n2354_n3888# 0.622383f
C82 minus.n9 a_n2354_n3888# 0.251893f
C83 minus.n10 a_n2354_n3888# 0.103999f
C84 minus.n11 a_n2354_n3888# 0.048587f
C85 minus.n12 a_n2354_n3888# 0.017466f
C86 minus.n13 a_n2354_n3888# 0.236925f
C87 minus.n14 a_n2354_n3888# 0.020012f
C88 minus.n15 a_n2354_n3888# 0.236925f
C89 minus.n16 a_n2354_n3888# 0.020012f
C90 minus.n17 a_n2354_n3888# 0.048587f
C91 minus.n18 a_n2354_n3888# 0.048587f
C92 minus.n19 a_n2354_n3888# 0.020012f
C93 minus.n20 a_n2354_n3888# 0.236925f
C94 minus.n21 a_n2354_n3888# 0.018065f
C95 minus.n22 a_n2354_n3888# 0.018065f
C96 minus.n23 a_n2354_n3888# 0.048587f
C97 minus.n24 a_n2354_n3888# 0.048587f
C98 minus.n25 a_n2354_n3888# 0.020012f
C99 minus.n26 a_n2354_n3888# 0.236925f
C100 minus.n27 a_n2354_n3888# 0.020012f
C101 minus.n28 a_n2354_n3888# 0.236925f
C102 minus.n29 a_n2354_n3888# 0.020012f
C103 minus.n30 a_n2354_n3888# 0.048587f
C104 minus.n31 a_n2354_n3888# 0.048587f
C105 minus.n32 a_n2354_n3888# 0.017466f
C106 minus.n33 a_n2354_n3888# 0.018664f
C107 minus.n34 a_n2354_n3888# 0.236925f
C108 minus.n35 a_n2354_n3888# 0.251828f
C109 minus.n36 a_n2354_n3888# 2.02132f
C110 minus.n37 a_n2354_n3888# 0.048587f
C111 minus.t14 a_n2354_n3888# 0.616823f
C112 minus.t7 a_n2354_n3888# 0.616823f
C113 minus.n38 a_n2354_n3888# 0.236925f
C114 minus.n39 a_n2354_n3888# 0.048587f
C115 minus.t21 a_n2354_n3888# 0.616823f
C116 minus.t22 a_n2354_n3888# 0.616823f
C117 minus.t11 a_n2354_n3888# 0.616823f
C118 minus.n40 a_n2354_n3888# 0.236925f
C119 minus.n41 a_n2354_n3888# 0.048587f
C120 minus.t23 a_n2354_n3888# 0.616823f
C121 minus.t12 a_n2354_n3888# 0.616823f
C122 minus.n42 a_n2354_n3888# 0.236925f
C123 minus.n43 a_n2354_n3888# 0.048587f
C124 minus.t17 a_n2354_n3888# 0.616823f
C125 minus.t4 a_n2354_n3888# 0.616823f
C126 minus.n44 a_n2354_n3888# 0.018664f
C127 minus.t5 a_n2354_n3888# 0.622383f
C128 minus.t18 a_n2354_n3888# 0.616823f
C129 minus.n45 a_n2354_n3888# 0.236925f
C130 minus.n46 a_n2354_n3888# 0.251893f
C131 minus.n47 a_n2354_n3888# 0.103999f
C132 minus.n48 a_n2354_n3888# 0.048587f
C133 minus.n49 a_n2354_n3888# 0.017466f
C134 minus.n50 a_n2354_n3888# 0.236925f
C135 minus.n51 a_n2354_n3888# 0.020012f
C136 minus.n52 a_n2354_n3888# 0.236925f
C137 minus.n53 a_n2354_n3888# 0.020012f
C138 minus.n54 a_n2354_n3888# 0.048587f
C139 minus.n55 a_n2354_n3888# 0.048587f
C140 minus.n56 a_n2354_n3888# 0.020012f
C141 minus.n57 a_n2354_n3888# 0.236925f
C142 minus.n58 a_n2354_n3888# 0.018065f
C143 minus.n59 a_n2354_n3888# 0.018065f
C144 minus.n60 a_n2354_n3888# 0.048587f
C145 minus.n61 a_n2354_n3888# 0.048587f
C146 minus.n62 a_n2354_n3888# 0.020012f
C147 minus.n63 a_n2354_n3888# 0.236925f
C148 minus.n64 a_n2354_n3888# 0.020012f
C149 minus.n65 a_n2354_n3888# 0.236925f
C150 minus.n66 a_n2354_n3888# 0.020012f
C151 minus.n67 a_n2354_n3888# 0.048587f
C152 minus.n68 a_n2354_n3888# 0.048587f
C153 minus.n69 a_n2354_n3888# 0.017466f
C154 minus.n70 a_n2354_n3888# 0.018664f
C155 minus.n71 a_n2354_n3888# 0.236925f
C156 minus.t6 a_n2354_n3888# 0.622383f
C157 minus.n72 a_n2354_n3888# 0.251828f
C158 minus.n73 a_n2354_n3888# 0.314234f
C159 minus.n74 a_n2354_n3888# 2.42676f
C160 source.t42 a_n2354_n3888# 4.02724f
C161 source.n0 a_n2354_n3888# 1.86534f
C162 source.t28 a_n2354_n3888# 0.359363f
C163 source.t47 a_n2354_n3888# 0.359363f
C164 source.n1 a_n2354_n3888# 3.1567f
C165 source.n2 a_n2354_n3888# 0.404738f
C166 source.t46 a_n2354_n3888# 0.359363f
C167 source.t35 a_n2354_n3888# 0.359363f
C168 source.n3 a_n2354_n3888# 3.1567f
C169 source.n4 a_n2354_n3888# 0.404738f
C170 source.t34 a_n2354_n3888# 0.359363f
C171 source.t27 a_n2354_n3888# 0.359363f
C172 source.n5 a_n2354_n3888# 3.1567f
C173 source.n6 a_n2354_n3888# 0.404738f
C174 source.t24 a_n2354_n3888# 0.359363f
C175 source.t37 a_n2354_n3888# 0.359363f
C176 source.n7 a_n2354_n3888# 3.1567f
C177 source.n8 a_n2354_n3888# 0.404738f
C178 source.t36 a_n2354_n3888# 0.359363f
C179 source.t31 a_n2354_n3888# 0.359363f
C180 source.n9 a_n2354_n3888# 3.1567f
C181 source.n10 a_n2354_n3888# 0.404738f
C182 source.t43 a_n2354_n3888# 4.02725f
C183 source.n11 a_n2354_n3888# 0.507117f
C184 source.t8 a_n2354_n3888# 4.02725f
C185 source.n12 a_n2354_n3888# 0.507117f
C186 source.t5 a_n2354_n3888# 0.359363f
C187 source.t17 a_n2354_n3888# 0.359363f
C188 source.n13 a_n2354_n3888# 3.1567f
C189 source.n14 a_n2354_n3888# 0.404738f
C190 source.t15 a_n2354_n3888# 0.359363f
C191 source.t16 a_n2354_n3888# 0.359363f
C192 source.n15 a_n2354_n3888# 3.1567f
C193 source.n16 a_n2354_n3888# 0.404738f
C194 source.t4 a_n2354_n3888# 0.359363f
C195 source.t12 a_n2354_n3888# 0.359363f
C196 source.n17 a_n2354_n3888# 3.1567f
C197 source.n18 a_n2354_n3888# 0.404738f
C198 source.t14 a_n2354_n3888# 0.359363f
C199 source.t22 a_n2354_n3888# 0.359363f
C200 source.n19 a_n2354_n3888# 3.1567f
C201 source.n20 a_n2354_n3888# 0.404738f
C202 source.t20 a_n2354_n3888# 0.359363f
C203 source.t9 a_n2354_n3888# 0.359363f
C204 source.n21 a_n2354_n3888# 3.1567f
C205 source.n22 a_n2354_n3888# 0.404738f
C206 source.t6 a_n2354_n3888# 4.02725f
C207 source.n23 a_n2354_n3888# 2.36939f
C208 source.t41 a_n2354_n3888# 4.02724f
C209 source.n24 a_n2354_n3888# 2.36939f
C210 source.t33 a_n2354_n3888# 0.359363f
C211 source.t25 a_n2354_n3888# 0.359363f
C212 source.n25 a_n2354_n3888# 3.1567f
C213 source.n26 a_n2354_n3888# 0.404742f
C214 source.t40 a_n2354_n3888# 0.359363f
C215 source.t26 a_n2354_n3888# 0.359363f
C216 source.n27 a_n2354_n3888# 3.1567f
C217 source.n28 a_n2354_n3888# 0.404742f
C218 source.t38 a_n2354_n3888# 0.359363f
C219 source.t29 a_n2354_n3888# 0.359363f
C220 source.n29 a_n2354_n3888# 3.1567f
C221 source.n30 a_n2354_n3888# 0.404742f
C222 source.t39 a_n2354_n3888# 0.359363f
C223 source.t30 a_n2354_n3888# 0.359363f
C224 source.n31 a_n2354_n3888# 3.1567f
C225 source.n32 a_n2354_n3888# 0.404742f
C226 source.t44 a_n2354_n3888# 0.359363f
C227 source.t32 a_n2354_n3888# 0.359363f
C228 source.n33 a_n2354_n3888# 3.1567f
C229 source.n34 a_n2354_n3888# 0.404742f
C230 source.t45 a_n2354_n3888# 4.02724f
C231 source.n35 a_n2354_n3888# 0.507122f
C232 source.t23 a_n2354_n3888# 4.02724f
C233 source.n36 a_n2354_n3888# 0.507122f
C234 source.t18 a_n2354_n3888# 0.359363f
C235 source.t19 a_n2354_n3888# 0.359363f
C236 source.n37 a_n2354_n3888# 3.1567f
C237 source.n38 a_n2354_n3888# 0.404742f
C238 source.t11 a_n2354_n3888# 0.359363f
C239 source.t1 a_n2354_n3888# 0.359363f
C240 source.n39 a_n2354_n3888# 3.1567f
C241 source.n40 a_n2354_n3888# 0.404742f
C242 source.t2 a_n2354_n3888# 0.359363f
C243 source.t21 a_n2354_n3888# 0.359363f
C244 source.n41 a_n2354_n3888# 3.1567f
C245 source.n42 a_n2354_n3888# 0.404742f
C246 source.t7 a_n2354_n3888# 0.359363f
C247 source.t3 a_n2354_n3888# 0.359363f
C248 source.n43 a_n2354_n3888# 3.1567f
C249 source.n44 a_n2354_n3888# 0.404742f
C250 source.t0 a_n2354_n3888# 0.359363f
C251 source.t10 a_n2354_n3888# 0.359363f
C252 source.n45 a_n2354_n3888# 3.1567f
C253 source.n46 a_n2354_n3888# 0.404742f
C254 source.t13 a_n2354_n3888# 4.02724f
C255 source.n47 a_n2354_n3888# 0.678262f
C256 source.n48 a_n2354_n3888# 2.21675f
C257 drain_left.t19 a_n2354_n3888# 0.407788f
C258 drain_left.t7 a_n2354_n3888# 0.407788f
C259 drain_left.n0 a_n2354_n3888# 3.68961f
C260 drain_left.t21 a_n2354_n3888# 0.407788f
C261 drain_left.t18 a_n2354_n3888# 0.407788f
C262 drain_left.n1 a_n2354_n3888# 3.68593f
C263 drain_left.n2 a_n2354_n3888# 0.81455f
C264 drain_left.t10 a_n2354_n3888# 0.407788f
C265 drain_left.t0 a_n2354_n3888# 0.407788f
C266 drain_left.n3 a_n2354_n3888# 3.68593f
C267 drain_left.n4 a_n2354_n3888# 0.369638f
C268 drain_left.t6 a_n2354_n3888# 0.407788f
C269 drain_left.t17 a_n2354_n3888# 0.407788f
C270 drain_left.n5 a_n2354_n3888# 3.68961f
C271 drain_left.t8 a_n2354_n3888# 0.407788f
C272 drain_left.t16 a_n2354_n3888# 0.407788f
C273 drain_left.n6 a_n2354_n3888# 3.68593f
C274 drain_left.n7 a_n2354_n3888# 0.81455f
C275 drain_left.t3 a_n2354_n3888# 0.407788f
C276 drain_left.t1 a_n2354_n3888# 0.407788f
C277 drain_left.n8 a_n2354_n3888# 3.68593f
C278 drain_left.n9 a_n2354_n3888# 0.369638f
C279 drain_left.n10 a_n2354_n3888# 2.11199f
C280 drain_left.t23 a_n2354_n3888# 0.407788f
C281 drain_left.t14 a_n2354_n3888# 0.407788f
C282 drain_left.n11 a_n2354_n3888# 3.68961f
C283 drain_left.t9 a_n2354_n3888# 0.407788f
C284 drain_left.t20 a_n2354_n3888# 0.407788f
C285 drain_left.n12 a_n2354_n3888# 3.68593f
C286 drain_left.n13 a_n2354_n3888# 0.814544f
C287 drain_left.t15 a_n2354_n3888# 0.407788f
C288 drain_left.t4 a_n2354_n3888# 0.407788f
C289 drain_left.n14 a_n2354_n3888# 3.68593f
C290 drain_left.n15 a_n2354_n3888# 0.402183f
C291 drain_left.t11 a_n2354_n3888# 0.407788f
C292 drain_left.t12 a_n2354_n3888# 0.407788f
C293 drain_left.n16 a_n2354_n3888# 3.68593f
C294 drain_left.n17 a_n2354_n3888# 0.402183f
C295 drain_left.t5 a_n2354_n3888# 0.407788f
C296 drain_left.t2 a_n2354_n3888# 0.407788f
C297 drain_left.n18 a_n2354_n3888# 3.68593f
C298 drain_left.n19 a_n2354_n3888# 0.402183f
C299 drain_left.t13 a_n2354_n3888# 0.407788f
C300 drain_left.t22 a_n2354_n3888# 0.407788f
C301 drain_left.n20 a_n2354_n3888# 3.68592f
C302 drain_left.n21 a_n2354_n3888# 0.688549f
C303 plus.n0 a_n2354_n3888# 0.049124f
C304 plus.t0 a_n2354_n3888# 0.623636f
C305 plus.t19 a_n2354_n3888# 0.623636f
C306 plus.n1 a_n2354_n3888# 0.239542f
C307 plus.n2 a_n2354_n3888# 0.049124f
C308 plus.t12 a_n2354_n3888# 0.623636f
C309 plus.t1 a_n2354_n3888# 0.623636f
C310 plus.t20 a_n2354_n3888# 0.623636f
C311 plus.n3 a_n2354_n3888# 0.239542f
C312 plus.n4 a_n2354_n3888# 0.049124f
C313 plus.t13 a_n2354_n3888# 0.623636f
C314 plus.t10 a_n2354_n3888# 0.623636f
C315 plus.n5 a_n2354_n3888# 0.239542f
C316 plus.n6 a_n2354_n3888# 0.049124f
C317 plus.t23 a_n2354_n3888# 0.623636f
C318 plus.t16 a_n2354_n3888# 0.623636f
C319 plus.n7 a_n2354_n3888# 0.01887f
C320 plus.t4 a_n2354_n3888# 0.629257f
C321 plus.t11 a_n2354_n3888# 0.623636f
C322 plus.n8 a_n2354_n3888# 0.239542f
C323 plus.n9 a_n2354_n3888# 0.254675f
C324 plus.n10 a_n2354_n3888# 0.105148f
C325 plus.n11 a_n2354_n3888# 0.049124f
C326 plus.n12 a_n2354_n3888# 0.017659f
C327 plus.n13 a_n2354_n3888# 0.239542f
C328 plus.n14 a_n2354_n3888# 0.020233f
C329 plus.n15 a_n2354_n3888# 0.239542f
C330 plus.n16 a_n2354_n3888# 0.020233f
C331 plus.n17 a_n2354_n3888# 0.049124f
C332 plus.n18 a_n2354_n3888# 0.049124f
C333 plus.n19 a_n2354_n3888# 0.020233f
C334 plus.n20 a_n2354_n3888# 0.239542f
C335 plus.n21 a_n2354_n3888# 0.018265f
C336 plus.n22 a_n2354_n3888# 0.018265f
C337 plus.n23 a_n2354_n3888# 0.049124f
C338 plus.n24 a_n2354_n3888# 0.049124f
C339 plus.n25 a_n2354_n3888# 0.020233f
C340 plus.n26 a_n2354_n3888# 0.239542f
C341 plus.n27 a_n2354_n3888# 0.020233f
C342 plus.n28 a_n2354_n3888# 0.239542f
C343 plus.n29 a_n2354_n3888# 0.020233f
C344 plus.n30 a_n2354_n3888# 0.049124f
C345 plus.n31 a_n2354_n3888# 0.049124f
C346 plus.n32 a_n2354_n3888# 0.017659f
C347 plus.n33 a_n2354_n3888# 0.01887f
C348 plus.n34 a_n2354_n3888# 0.239542f
C349 plus.t5 a_n2354_n3888# 0.629257f
C350 plus.n35 a_n2354_n3888# 0.254609f
C351 plus.n36 a_n2354_n3888# 0.617319f
C352 plus.n37 a_n2354_n3888# 0.049124f
C353 plus.t6 a_n2354_n3888# 0.629257f
C354 plus.t14 a_n2354_n3888# 0.623636f
C355 plus.t22 a_n2354_n3888# 0.623636f
C356 plus.n38 a_n2354_n3888# 0.239542f
C357 plus.n39 a_n2354_n3888# 0.049124f
C358 plus.t7 a_n2354_n3888# 0.623636f
C359 plus.t21 a_n2354_n3888# 0.623636f
C360 plus.t9 a_n2354_n3888# 0.623636f
C361 plus.n40 a_n2354_n3888# 0.239542f
C362 plus.n41 a_n2354_n3888# 0.049124f
C363 plus.t18 a_n2354_n3888# 0.623636f
C364 plus.t8 a_n2354_n3888# 0.623636f
C365 plus.n42 a_n2354_n3888# 0.239542f
C366 plus.n43 a_n2354_n3888# 0.049124f
C367 plus.t17 a_n2354_n3888# 0.623636f
C368 plus.t3 a_n2354_n3888# 0.623636f
C369 plus.n44 a_n2354_n3888# 0.01887f
C370 plus.t15 a_n2354_n3888# 0.623636f
C371 plus.n45 a_n2354_n3888# 0.239542f
C372 plus.t2 a_n2354_n3888# 0.629257f
C373 plus.n46 a_n2354_n3888# 0.254675f
C374 plus.n47 a_n2354_n3888# 0.105148f
C375 plus.n48 a_n2354_n3888# 0.049124f
C376 plus.n49 a_n2354_n3888# 0.017659f
C377 plus.n50 a_n2354_n3888# 0.239542f
C378 plus.n51 a_n2354_n3888# 0.020233f
C379 plus.n52 a_n2354_n3888# 0.239542f
C380 plus.n53 a_n2354_n3888# 0.020233f
C381 plus.n54 a_n2354_n3888# 0.049124f
C382 plus.n55 a_n2354_n3888# 0.049124f
C383 plus.n56 a_n2354_n3888# 0.020233f
C384 plus.n57 a_n2354_n3888# 0.239542f
C385 plus.n58 a_n2354_n3888# 0.018265f
C386 plus.n59 a_n2354_n3888# 0.018265f
C387 plus.n60 a_n2354_n3888# 0.049124f
C388 plus.n61 a_n2354_n3888# 0.049124f
C389 plus.n62 a_n2354_n3888# 0.020233f
C390 plus.n63 a_n2354_n3888# 0.239542f
C391 plus.n64 a_n2354_n3888# 0.020233f
C392 plus.n65 a_n2354_n3888# 0.239542f
C393 plus.n66 a_n2354_n3888# 0.020233f
C394 plus.n67 a_n2354_n3888# 0.049124f
C395 plus.n68 a_n2354_n3888# 0.049124f
C396 plus.n69 a_n2354_n3888# 0.017659f
C397 plus.n70 a_n2354_n3888# 0.01887f
C398 plus.n71 a_n2354_n3888# 0.239542f
C399 plus.n72 a_n2354_n3888# 0.254609f
C400 plus.n73 a_n2354_n3888# 1.69071f
.ends

