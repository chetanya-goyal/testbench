* NGSPICE file created from diffpair256.ext - technology: sky130A

.subckt diffpair256 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t14 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X1 drain_right.t12 minus.t1 source.t15 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 drain_right.t11 minus.t2 source.t16 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X3 drain_right.t10 minus.t3 source.t17 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 drain_left.t13 plus.t0 source.t8 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X5 source.t0 plus.t1 drain_left.t12 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X6 source.t10 plus.t2 drain_left.t11 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 source.t18 minus.t4 drain_right.t9 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X8 source.t3 plus.t3 drain_left.t10 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X9 source.t19 minus.t5 drain_right.t8 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X10 a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X11 a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X12 drain_left.t9 plus.t4 source.t1 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X13 source.t2 plus.t5 drain_left.t8 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X14 drain_left.t7 plus.t6 source.t4 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X15 drain_left.t6 plus.t7 source.t6 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X16 drain_left.t5 plus.t8 source.t9 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X17 drain_left.t4 plus.t9 source.t7 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X18 drain_right.t7 minus.t6 source.t20 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X19 drain_right.t6 minus.t7 source.t24 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X20 source.t13 plus.t10 drain_left.t3 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X21 a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X22 drain_left.t2 plus.t11 source.t5 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X23 source.t11 plus.t12 drain_left.t1 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X24 drain_right.t5 minus.t8 source.t25 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X25 drain_right.t4 minus.t9 source.t21 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X26 source.t26 minus.t10 drain_right.t3 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X27 a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X28 source.t22 minus.t11 drain_right.t2 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X29 source.t23 minus.t12 drain_right.t1 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X30 drain_left.t0 plus.t13 source.t12 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X31 source.t27 minus.t13 drain_right.t0 a_n1564_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n14 minus.t2 929.312
R1 minus.n3 minus.t6 929.312
R2 minus.n30 minus.t0 929.312
R3 minus.n19 minus.t9 929.312
R4 minus.n13 minus.t4 879.65
R5 minus.n11 minus.t7 879.65
R6 minus.n1 minus.t10 879.65
R7 minus.n6 minus.t1 879.65
R8 minus.n4 minus.t5 879.65
R9 minus.n29 minus.t13 879.65
R10 minus.n27 minus.t3 879.65
R11 minus.n17 minus.t11 879.65
R12 minus.n22 minus.t8 879.65
R13 minus.n20 minus.t12 879.65
R14 minus.n3 minus.n2 161.489
R15 minus.n19 minus.n18 161.489
R16 minus.n15 minus.n14 161.3
R17 minus.n12 minus.n0 161.3
R18 minus.n10 minus.n9 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n5 minus.n2 161.3
R21 minus.n31 minus.n30 161.3
R22 minus.n28 minus.n16 161.3
R23 minus.n26 minus.n25 161.3
R24 minus.n24 minus.n23 161.3
R25 minus.n21 minus.n18 161.3
R26 minus.n13 minus.n12 45.2793
R27 minus.n5 minus.n4 45.2793
R28 minus.n21 minus.n20 45.2793
R29 minus.n29 minus.n28 45.2793
R30 minus.n11 minus.n10 40.8975
R31 minus.n7 minus.n6 40.8975
R32 minus.n23 minus.n22 40.8975
R33 minus.n27 minus.n26 40.8975
R34 minus.n10 minus.n1 36.5157
R35 minus.n7 minus.n1 36.5157
R36 minus.n23 minus.n17 36.5157
R37 minus.n26 minus.n17 36.5157
R38 minus.n12 minus.n11 32.1338
R39 minus.n6 minus.n5 32.1338
R40 minus.n22 minus.n21 32.1338
R41 minus.n28 minus.n27 32.1338
R42 minus.n32 minus.n15 30.4607
R43 minus.n14 minus.n13 27.752
R44 minus.n4 minus.n3 27.752
R45 minus.n20 minus.n19 27.752
R46 minus.n30 minus.n29 27.752
R47 minus.n32 minus.n31 6.46073
R48 minus.n15 minus.n0 0.189894
R49 minus.n9 minus.n0 0.189894
R50 minus.n9 minus.n8 0.189894
R51 minus.n8 minus.n2 0.189894
R52 minus.n24 minus.n18 0.189894
R53 minus.n25 minus.n24 0.189894
R54 minus.n25 minus.n16 0.189894
R55 minus.n31 minus.n16 0.189894
R56 minus minus.n32 0.188
R57 source.n146 source.n120 289.615
R58 source.n108 source.n82 289.615
R59 source.n26 source.n0 289.615
R60 source.n64 source.n38 289.615
R61 source.n131 source.n130 185
R62 source.n128 source.n127 185
R63 source.n137 source.n136 185
R64 source.n139 source.n138 185
R65 source.n124 source.n123 185
R66 source.n145 source.n144 185
R67 source.n147 source.n146 185
R68 source.n93 source.n92 185
R69 source.n90 source.n89 185
R70 source.n99 source.n98 185
R71 source.n101 source.n100 185
R72 source.n86 source.n85 185
R73 source.n107 source.n106 185
R74 source.n109 source.n108 185
R75 source.n27 source.n26 185
R76 source.n25 source.n24 185
R77 source.n4 source.n3 185
R78 source.n19 source.n18 185
R79 source.n17 source.n16 185
R80 source.n8 source.n7 185
R81 source.n11 source.n10 185
R82 source.n65 source.n64 185
R83 source.n63 source.n62 185
R84 source.n42 source.n41 185
R85 source.n57 source.n56 185
R86 source.n55 source.n54 185
R87 source.n46 source.n45 185
R88 source.n49 source.n48 185
R89 source.t14 source.n129 147.661
R90 source.t7 source.n91 147.661
R91 source.t8 source.n9 147.661
R92 source.t20 source.n47 147.661
R93 source.n130 source.n127 104.615
R94 source.n137 source.n127 104.615
R95 source.n138 source.n137 104.615
R96 source.n138 source.n123 104.615
R97 source.n145 source.n123 104.615
R98 source.n146 source.n145 104.615
R99 source.n92 source.n89 104.615
R100 source.n99 source.n89 104.615
R101 source.n100 source.n99 104.615
R102 source.n100 source.n85 104.615
R103 source.n107 source.n85 104.615
R104 source.n108 source.n107 104.615
R105 source.n26 source.n25 104.615
R106 source.n25 source.n3 104.615
R107 source.n18 source.n3 104.615
R108 source.n18 source.n17 104.615
R109 source.n17 source.n7 104.615
R110 source.n10 source.n7 104.615
R111 source.n64 source.n63 104.615
R112 source.n63 source.n41 104.615
R113 source.n56 source.n41 104.615
R114 source.n56 source.n55 104.615
R115 source.n55 source.n45 104.615
R116 source.n48 source.n45 104.615
R117 source.n130 source.t14 52.3082
R118 source.n92 source.t7 52.3082
R119 source.n10 source.t8 52.3082
R120 source.n48 source.t20 52.3082
R121 source.n33 source.n32 50.512
R122 source.n35 source.n34 50.512
R123 source.n37 source.n36 50.512
R124 source.n71 source.n70 50.512
R125 source.n73 source.n72 50.512
R126 source.n75 source.n74 50.512
R127 source.n119 source.n118 50.5119
R128 source.n117 source.n116 50.5119
R129 source.n115 source.n114 50.5119
R130 source.n81 source.n80 50.5119
R131 source.n79 source.n78 50.5119
R132 source.n77 source.n76 50.5119
R133 source.n151 source.n150 32.1853
R134 source.n113 source.n112 32.1853
R135 source.n31 source.n30 32.1853
R136 source.n69 source.n68 32.1853
R137 source.n77 source.n75 17.6561
R138 source.n131 source.n129 15.6674
R139 source.n93 source.n91 15.6674
R140 source.n11 source.n9 15.6674
R141 source.n49 source.n47 15.6674
R142 source.n132 source.n128 12.8005
R143 source.n94 source.n90 12.8005
R144 source.n12 source.n8 12.8005
R145 source.n50 source.n46 12.8005
R146 source.n136 source.n135 12.0247
R147 source.n98 source.n97 12.0247
R148 source.n16 source.n15 12.0247
R149 source.n54 source.n53 12.0247
R150 source.n152 source.n31 11.7078
R151 source.n139 source.n126 11.249
R152 source.n101 source.n88 11.249
R153 source.n19 source.n6 11.249
R154 source.n57 source.n44 11.249
R155 source.n140 source.n124 10.4732
R156 source.n102 source.n86 10.4732
R157 source.n20 source.n4 10.4732
R158 source.n58 source.n42 10.4732
R159 source.n144 source.n143 9.69747
R160 source.n106 source.n105 9.69747
R161 source.n24 source.n23 9.69747
R162 source.n62 source.n61 9.69747
R163 source.n150 source.n149 9.45567
R164 source.n112 source.n111 9.45567
R165 source.n30 source.n29 9.45567
R166 source.n68 source.n67 9.45567
R167 source.n149 source.n148 9.3005
R168 source.n122 source.n121 9.3005
R169 source.n143 source.n142 9.3005
R170 source.n141 source.n140 9.3005
R171 source.n126 source.n125 9.3005
R172 source.n135 source.n134 9.3005
R173 source.n133 source.n132 9.3005
R174 source.n111 source.n110 9.3005
R175 source.n84 source.n83 9.3005
R176 source.n105 source.n104 9.3005
R177 source.n103 source.n102 9.3005
R178 source.n88 source.n87 9.3005
R179 source.n97 source.n96 9.3005
R180 source.n95 source.n94 9.3005
R181 source.n29 source.n28 9.3005
R182 source.n2 source.n1 9.3005
R183 source.n23 source.n22 9.3005
R184 source.n21 source.n20 9.3005
R185 source.n6 source.n5 9.3005
R186 source.n15 source.n14 9.3005
R187 source.n13 source.n12 9.3005
R188 source.n67 source.n66 9.3005
R189 source.n40 source.n39 9.3005
R190 source.n61 source.n60 9.3005
R191 source.n59 source.n58 9.3005
R192 source.n44 source.n43 9.3005
R193 source.n53 source.n52 9.3005
R194 source.n51 source.n50 9.3005
R195 source.n147 source.n122 8.92171
R196 source.n109 source.n84 8.92171
R197 source.n27 source.n2 8.92171
R198 source.n65 source.n40 8.92171
R199 source.n148 source.n120 8.14595
R200 source.n110 source.n82 8.14595
R201 source.n28 source.n0 8.14595
R202 source.n66 source.n38 8.14595
R203 source.n150 source.n120 5.81868
R204 source.n112 source.n82 5.81868
R205 source.n30 source.n0 5.81868
R206 source.n68 source.n38 5.81868
R207 source.n152 source.n151 5.49188
R208 source.n148 source.n147 5.04292
R209 source.n110 source.n109 5.04292
R210 source.n28 source.n27 5.04292
R211 source.n66 source.n65 5.04292
R212 source.n133 source.n129 4.38594
R213 source.n95 source.n91 4.38594
R214 source.n13 source.n9 4.38594
R215 source.n51 source.n47 4.38594
R216 source.n144 source.n122 4.26717
R217 source.n106 source.n84 4.26717
R218 source.n24 source.n2 4.26717
R219 source.n62 source.n40 4.26717
R220 source.n143 source.n124 3.49141
R221 source.n105 source.n86 3.49141
R222 source.n23 source.n4 3.49141
R223 source.n61 source.n42 3.49141
R224 source.n118 source.t17 3.3005
R225 source.n118 source.t27 3.3005
R226 source.n116 source.t25 3.3005
R227 source.n116 source.t22 3.3005
R228 source.n114 source.t21 3.3005
R229 source.n114 source.t23 3.3005
R230 source.n80 source.t6 3.3005
R231 source.n80 source.t13 3.3005
R232 source.n78 source.t9 3.3005
R233 source.n78 source.t3 3.3005
R234 source.n76 source.t1 3.3005
R235 source.n76 source.t10 3.3005
R236 source.n32 source.t5 3.3005
R237 source.n32 source.t2 3.3005
R238 source.n34 source.t12 3.3005
R239 source.n34 source.t11 3.3005
R240 source.n36 source.t4 3.3005
R241 source.n36 source.t0 3.3005
R242 source.n70 source.t15 3.3005
R243 source.n70 source.t19 3.3005
R244 source.n72 source.t24 3.3005
R245 source.n72 source.t26 3.3005
R246 source.n74 source.t16 3.3005
R247 source.n74 source.t18 3.3005
R248 source.n140 source.n139 2.71565
R249 source.n102 source.n101 2.71565
R250 source.n20 source.n19 2.71565
R251 source.n58 source.n57 2.71565
R252 source.n136 source.n126 1.93989
R253 source.n98 source.n88 1.93989
R254 source.n16 source.n6 1.93989
R255 source.n54 source.n44 1.93989
R256 source.n135 source.n128 1.16414
R257 source.n97 source.n90 1.16414
R258 source.n15 source.n8 1.16414
R259 source.n53 source.n46 1.16414
R260 source.n69 source.n37 0.698776
R261 source.n115 source.n113 0.698776
R262 source.n75 source.n73 0.457397
R263 source.n73 source.n71 0.457397
R264 source.n71 source.n69 0.457397
R265 source.n37 source.n35 0.457397
R266 source.n35 source.n33 0.457397
R267 source.n33 source.n31 0.457397
R268 source.n79 source.n77 0.457397
R269 source.n81 source.n79 0.457397
R270 source.n113 source.n81 0.457397
R271 source.n117 source.n115 0.457397
R272 source.n119 source.n117 0.457397
R273 source.n151 source.n119 0.457397
R274 source.n132 source.n131 0.388379
R275 source.n94 source.n93 0.388379
R276 source.n12 source.n11 0.388379
R277 source.n50 source.n49 0.388379
R278 source source.n152 0.188
R279 source.n134 source.n133 0.155672
R280 source.n134 source.n125 0.155672
R281 source.n141 source.n125 0.155672
R282 source.n142 source.n141 0.155672
R283 source.n142 source.n121 0.155672
R284 source.n149 source.n121 0.155672
R285 source.n96 source.n95 0.155672
R286 source.n96 source.n87 0.155672
R287 source.n103 source.n87 0.155672
R288 source.n104 source.n103 0.155672
R289 source.n104 source.n83 0.155672
R290 source.n111 source.n83 0.155672
R291 source.n29 source.n1 0.155672
R292 source.n22 source.n1 0.155672
R293 source.n22 source.n21 0.155672
R294 source.n21 source.n5 0.155672
R295 source.n14 source.n5 0.155672
R296 source.n14 source.n13 0.155672
R297 source.n67 source.n39 0.155672
R298 source.n60 source.n39 0.155672
R299 source.n60 source.n59 0.155672
R300 source.n59 source.n43 0.155672
R301 source.n52 source.n43 0.155672
R302 source.n52 source.n51 0.155672
R303 drain_right.n26 drain_right.n0 289.615
R304 drain_right.n68 drain_right.n42 289.615
R305 drain_right.n11 drain_right.n10 185
R306 drain_right.n8 drain_right.n7 185
R307 drain_right.n17 drain_right.n16 185
R308 drain_right.n19 drain_right.n18 185
R309 drain_right.n4 drain_right.n3 185
R310 drain_right.n25 drain_right.n24 185
R311 drain_right.n27 drain_right.n26 185
R312 drain_right.n69 drain_right.n68 185
R313 drain_right.n67 drain_right.n66 185
R314 drain_right.n46 drain_right.n45 185
R315 drain_right.n61 drain_right.n60 185
R316 drain_right.n59 drain_right.n58 185
R317 drain_right.n50 drain_right.n49 185
R318 drain_right.n53 drain_right.n52 185
R319 drain_right.t4 drain_right.n9 147.661
R320 drain_right.t11 drain_right.n51 147.661
R321 drain_right.n10 drain_right.n7 104.615
R322 drain_right.n17 drain_right.n7 104.615
R323 drain_right.n18 drain_right.n17 104.615
R324 drain_right.n18 drain_right.n3 104.615
R325 drain_right.n25 drain_right.n3 104.615
R326 drain_right.n26 drain_right.n25 104.615
R327 drain_right.n68 drain_right.n67 104.615
R328 drain_right.n67 drain_right.n45 104.615
R329 drain_right.n60 drain_right.n45 104.615
R330 drain_right.n60 drain_right.n59 104.615
R331 drain_right.n59 drain_right.n49 104.615
R332 drain_right.n52 drain_right.n49 104.615
R333 drain_right.n35 drain_right.n33 67.6476
R334 drain_right.n39 drain_right.n37 67.6476
R335 drain_right.n39 drain_right.n38 67.1908
R336 drain_right.n41 drain_right.n40 67.1908
R337 drain_right.n35 drain_right.n34 67.1907
R338 drain_right.n32 drain_right.n31 67.1907
R339 drain_right.n10 drain_right.t4 52.3082
R340 drain_right.n52 drain_right.t11 52.3082
R341 drain_right.n32 drain_right.n30 49.321
R342 drain_right.n73 drain_right.n72 48.8641
R343 drain_right drain_right.n36 24.8955
R344 drain_right.n11 drain_right.n9 15.6674
R345 drain_right.n53 drain_right.n51 15.6674
R346 drain_right.n12 drain_right.n8 12.8005
R347 drain_right.n54 drain_right.n50 12.8005
R348 drain_right.n16 drain_right.n15 12.0247
R349 drain_right.n58 drain_right.n57 12.0247
R350 drain_right.n19 drain_right.n6 11.249
R351 drain_right.n61 drain_right.n48 11.249
R352 drain_right.n20 drain_right.n4 10.4732
R353 drain_right.n62 drain_right.n46 10.4732
R354 drain_right.n24 drain_right.n23 9.69747
R355 drain_right.n66 drain_right.n65 9.69747
R356 drain_right.n30 drain_right.n29 9.45567
R357 drain_right.n72 drain_right.n71 9.45567
R358 drain_right.n29 drain_right.n28 9.3005
R359 drain_right.n2 drain_right.n1 9.3005
R360 drain_right.n23 drain_right.n22 9.3005
R361 drain_right.n21 drain_right.n20 9.3005
R362 drain_right.n6 drain_right.n5 9.3005
R363 drain_right.n15 drain_right.n14 9.3005
R364 drain_right.n13 drain_right.n12 9.3005
R365 drain_right.n71 drain_right.n70 9.3005
R366 drain_right.n44 drain_right.n43 9.3005
R367 drain_right.n65 drain_right.n64 9.3005
R368 drain_right.n63 drain_right.n62 9.3005
R369 drain_right.n48 drain_right.n47 9.3005
R370 drain_right.n57 drain_right.n56 9.3005
R371 drain_right.n55 drain_right.n54 9.3005
R372 drain_right.n27 drain_right.n2 8.92171
R373 drain_right.n69 drain_right.n44 8.92171
R374 drain_right.n28 drain_right.n0 8.14595
R375 drain_right.n70 drain_right.n42 8.14595
R376 drain_right drain_right.n73 5.88166
R377 drain_right.n30 drain_right.n0 5.81868
R378 drain_right.n72 drain_right.n42 5.81868
R379 drain_right.n28 drain_right.n27 5.04292
R380 drain_right.n70 drain_right.n69 5.04292
R381 drain_right.n13 drain_right.n9 4.38594
R382 drain_right.n55 drain_right.n51 4.38594
R383 drain_right.n24 drain_right.n2 4.26717
R384 drain_right.n66 drain_right.n44 4.26717
R385 drain_right.n23 drain_right.n4 3.49141
R386 drain_right.n65 drain_right.n46 3.49141
R387 drain_right.n33 drain_right.t0 3.3005
R388 drain_right.n33 drain_right.t13 3.3005
R389 drain_right.n34 drain_right.t2 3.3005
R390 drain_right.n34 drain_right.t10 3.3005
R391 drain_right.n31 drain_right.t1 3.3005
R392 drain_right.n31 drain_right.t5 3.3005
R393 drain_right.n37 drain_right.t8 3.3005
R394 drain_right.n37 drain_right.t7 3.3005
R395 drain_right.n38 drain_right.t3 3.3005
R396 drain_right.n38 drain_right.t12 3.3005
R397 drain_right.n40 drain_right.t9 3.3005
R398 drain_right.n40 drain_right.t6 3.3005
R399 drain_right.n20 drain_right.n19 2.71565
R400 drain_right.n62 drain_right.n61 2.71565
R401 drain_right.n16 drain_right.n6 1.93989
R402 drain_right.n58 drain_right.n48 1.93989
R403 drain_right.n15 drain_right.n8 1.16414
R404 drain_right.n57 drain_right.n50 1.16414
R405 drain_right.n73 drain_right.n41 0.457397
R406 drain_right.n41 drain_right.n39 0.457397
R407 drain_right.n12 drain_right.n11 0.388379
R408 drain_right.n54 drain_right.n53 0.388379
R409 drain_right.n36 drain_right.n32 0.287826
R410 drain_right.n14 drain_right.n13 0.155672
R411 drain_right.n14 drain_right.n5 0.155672
R412 drain_right.n21 drain_right.n5 0.155672
R413 drain_right.n22 drain_right.n21 0.155672
R414 drain_right.n22 drain_right.n1 0.155672
R415 drain_right.n29 drain_right.n1 0.155672
R416 drain_right.n71 drain_right.n43 0.155672
R417 drain_right.n64 drain_right.n43 0.155672
R418 drain_right.n64 drain_right.n63 0.155672
R419 drain_right.n63 drain_right.n47 0.155672
R420 drain_right.n56 drain_right.n47 0.155672
R421 drain_right.n56 drain_right.n55 0.155672
R422 drain_right.n36 drain_right.n35 0.0593781
R423 plus.n3 plus.t6 929.312
R424 plus.n14 plus.t0 929.312
R425 plus.n19 plus.t9 929.312
R426 plus.n30 plus.t4 929.312
R427 plus.n4 plus.t1 879.65
R428 plus.n6 plus.t13 879.65
R429 plus.n1 plus.t12 879.65
R430 plus.n11 plus.t11 879.65
R431 plus.n13 plus.t5 879.65
R432 plus.n20 plus.t10 879.65
R433 plus.n22 plus.t7 879.65
R434 plus.n17 plus.t3 879.65
R435 plus.n27 plus.t8 879.65
R436 plus.n29 plus.t2 879.65
R437 plus.n3 plus.n2 161.489
R438 plus.n19 plus.n18 161.489
R439 plus.n5 plus.n2 161.3
R440 plus.n8 plus.n7 161.3
R441 plus.n10 plus.n9 161.3
R442 plus.n12 plus.n0 161.3
R443 plus.n15 plus.n14 161.3
R444 plus.n21 plus.n18 161.3
R445 plus.n24 plus.n23 161.3
R446 plus.n26 plus.n25 161.3
R447 plus.n28 plus.n16 161.3
R448 plus.n31 plus.n30 161.3
R449 plus.n5 plus.n4 45.2793
R450 plus.n13 plus.n12 45.2793
R451 plus.n29 plus.n28 45.2793
R452 plus.n21 plus.n20 45.2793
R453 plus.n7 plus.n6 40.8975
R454 plus.n11 plus.n10 40.8975
R455 plus.n27 plus.n26 40.8975
R456 plus.n23 plus.n22 40.8975
R457 plus.n7 plus.n1 36.5157
R458 plus.n10 plus.n1 36.5157
R459 plus.n26 plus.n17 36.5157
R460 plus.n23 plus.n17 36.5157
R461 plus.n6 plus.n5 32.1338
R462 plus.n12 plus.n11 32.1338
R463 plus.n28 plus.n27 32.1338
R464 plus.n22 plus.n21 32.1338
R465 plus.n4 plus.n3 27.752
R466 plus.n14 plus.n13 27.752
R467 plus.n30 plus.n29 27.752
R468 plus.n20 plus.n19 27.752
R469 plus plus.n31 26.6146
R470 plus plus.n15 9.83194
R471 plus.n8 plus.n2 0.189894
R472 plus.n9 plus.n8 0.189894
R473 plus.n9 plus.n0 0.189894
R474 plus.n15 plus.n0 0.189894
R475 plus.n31 plus.n16 0.189894
R476 plus.n25 plus.n16 0.189894
R477 plus.n25 plus.n24 0.189894
R478 plus.n24 plus.n18 0.189894
R479 drain_left.n26 drain_left.n0 289.615
R480 drain_left.n63 drain_left.n37 289.615
R481 drain_left.n11 drain_left.n10 185
R482 drain_left.n8 drain_left.n7 185
R483 drain_left.n17 drain_left.n16 185
R484 drain_left.n19 drain_left.n18 185
R485 drain_left.n4 drain_left.n3 185
R486 drain_left.n25 drain_left.n24 185
R487 drain_left.n27 drain_left.n26 185
R488 drain_left.n64 drain_left.n63 185
R489 drain_left.n62 drain_left.n61 185
R490 drain_left.n41 drain_left.n40 185
R491 drain_left.n56 drain_left.n55 185
R492 drain_left.n54 drain_left.n53 185
R493 drain_left.n45 drain_left.n44 185
R494 drain_left.n48 drain_left.n47 185
R495 drain_left.t9 drain_left.n9 147.661
R496 drain_left.t7 drain_left.n46 147.661
R497 drain_left.n10 drain_left.n7 104.615
R498 drain_left.n17 drain_left.n7 104.615
R499 drain_left.n18 drain_left.n17 104.615
R500 drain_left.n18 drain_left.n3 104.615
R501 drain_left.n25 drain_left.n3 104.615
R502 drain_left.n26 drain_left.n25 104.615
R503 drain_left.n63 drain_left.n62 104.615
R504 drain_left.n62 drain_left.n40 104.615
R505 drain_left.n55 drain_left.n40 104.615
R506 drain_left.n55 drain_left.n54 104.615
R507 drain_left.n54 drain_left.n44 104.615
R508 drain_left.n47 drain_left.n44 104.615
R509 drain_left.n35 drain_left.n33 67.6476
R510 drain_left.n71 drain_left.n70 67.1908
R511 drain_left.n69 drain_left.n68 67.1908
R512 drain_left.n73 drain_left.n72 67.1907
R513 drain_left.n35 drain_left.n34 67.1907
R514 drain_left.n32 drain_left.n31 67.1907
R515 drain_left.n10 drain_left.t9 52.3082
R516 drain_left.n47 drain_left.t7 52.3082
R517 drain_left.n32 drain_left.n30 49.321
R518 drain_left.n69 drain_left.n67 49.321
R519 drain_left drain_left.n36 25.4488
R520 drain_left.n11 drain_left.n9 15.6674
R521 drain_left.n48 drain_left.n46 15.6674
R522 drain_left.n12 drain_left.n8 12.8005
R523 drain_left.n49 drain_left.n45 12.8005
R524 drain_left.n16 drain_left.n15 12.0247
R525 drain_left.n53 drain_left.n52 12.0247
R526 drain_left.n19 drain_left.n6 11.249
R527 drain_left.n56 drain_left.n43 11.249
R528 drain_left.n20 drain_left.n4 10.4732
R529 drain_left.n57 drain_left.n41 10.4732
R530 drain_left.n24 drain_left.n23 9.69747
R531 drain_left.n61 drain_left.n60 9.69747
R532 drain_left.n30 drain_left.n29 9.45567
R533 drain_left.n67 drain_left.n66 9.45567
R534 drain_left.n29 drain_left.n28 9.3005
R535 drain_left.n2 drain_left.n1 9.3005
R536 drain_left.n23 drain_left.n22 9.3005
R537 drain_left.n21 drain_left.n20 9.3005
R538 drain_left.n6 drain_left.n5 9.3005
R539 drain_left.n15 drain_left.n14 9.3005
R540 drain_left.n13 drain_left.n12 9.3005
R541 drain_left.n66 drain_left.n65 9.3005
R542 drain_left.n39 drain_left.n38 9.3005
R543 drain_left.n60 drain_left.n59 9.3005
R544 drain_left.n58 drain_left.n57 9.3005
R545 drain_left.n43 drain_left.n42 9.3005
R546 drain_left.n52 drain_left.n51 9.3005
R547 drain_left.n50 drain_left.n49 9.3005
R548 drain_left.n27 drain_left.n2 8.92171
R549 drain_left.n64 drain_left.n39 8.92171
R550 drain_left.n28 drain_left.n0 8.14595
R551 drain_left.n65 drain_left.n37 8.14595
R552 drain_left drain_left.n73 6.11011
R553 drain_left.n30 drain_left.n0 5.81868
R554 drain_left.n67 drain_left.n37 5.81868
R555 drain_left.n28 drain_left.n27 5.04292
R556 drain_left.n65 drain_left.n64 5.04292
R557 drain_left.n13 drain_left.n9 4.38594
R558 drain_left.n50 drain_left.n46 4.38594
R559 drain_left.n24 drain_left.n2 4.26717
R560 drain_left.n61 drain_left.n39 4.26717
R561 drain_left.n23 drain_left.n4 3.49141
R562 drain_left.n60 drain_left.n41 3.49141
R563 drain_left.n33 drain_left.t3 3.3005
R564 drain_left.n33 drain_left.t4 3.3005
R565 drain_left.n34 drain_left.t10 3.3005
R566 drain_left.n34 drain_left.t6 3.3005
R567 drain_left.n31 drain_left.t11 3.3005
R568 drain_left.n31 drain_left.t5 3.3005
R569 drain_left.n72 drain_left.t8 3.3005
R570 drain_left.n72 drain_left.t13 3.3005
R571 drain_left.n70 drain_left.t1 3.3005
R572 drain_left.n70 drain_left.t2 3.3005
R573 drain_left.n68 drain_left.t12 3.3005
R574 drain_left.n68 drain_left.t0 3.3005
R575 drain_left.n20 drain_left.n19 2.71565
R576 drain_left.n57 drain_left.n56 2.71565
R577 drain_left.n16 drain_left.n6 1.93989
R578 drain_left.n53 drain_left.n43 1.93989
R579 drain_left.n15 drain_left.n8 1.16414
R580 drain_left.n52 drain_left.n45 1.16414
R581 drain_left.n71 drain_left.n69 0.457397
R582 drain_left.n73 drain_left.n71 0.457397
R583 drain_left.n12 drain_left.n11 0.388379
R584 drain_left.n49 drain_left.n48 0.388379
R585 drain_left.n36 drain_left.n32 0.287826
R586 drain_left.n14 drain_left.n13 0.155672
R587 drain_left.n14 drain_left.n5 0.155672
R588 drain_left.n21 drain_left.n5 0.155672
R589 drain_left.n22 drain_left.n21 0.155672
R590 drain_left.n22 drain_left.n1 0.155672
R591 drain_left.n29 drain_left.n1 0.155672
R592 drain_left.n66 drain_left.n38 0.155672
R593 drain_left.n59 drain_left.n38 0.155672
R594 drain_left.n59 drain_left.n58 0.155672
R595 drain_left.n58 drain_left.n42 0.155672
R596 drain_left.n51 drain_left.n42 0.155672
R597 drain_left.n51 drain_left.n50 0.155672
R598 drain_left.n36 drain_left.n35 0.0593781
C0 plus drain_right 0.305003f
C1 drain_right source 17.9885f
C2 drain_right minus 2.21837f
C3 drain_right drain_left 0.792804f
C4 plus source 2.11939f
C5 plus minus 3.99389f
C6 minus source 2.10502f
C7 plus drain_left 2.36689f
C8 drain_left source 17.9951f
C9 drain_left minus 0.171065f
C10 drain_right a_n1564_n2088# 5.54197f
C11 drain_left a_n1564_n2088# 5.81298f
C12 source a_n1564_n2088# 3.897421f
C13 minus a_n1564_n2088# 5.589329f
C14 plus a_n1564_n2088# 7.22225f
C15 drain_left.n0 a_n1564_n2088# 0.048119f
C16 drain_left.n1 a_n1564_n2088# 0.034234f
C17 drain_left.n2 a_n1564_n2088# 0.018396f
C18 drain_left.n3 a_n1564_n2088# 0.043481f
C19 drain_left.n4 a_n1564_n2088# 0.019478f
C20 drain_left.n5 a_n1564_n2088# 0.034234f
C21 drain_left.n6 a_n1564_n2088# 0.018396f
C22 drain_left.n7 a_n1564_n2088# 0.043481f
C23 drain_left.n8 a_n1564_n2088# 0.019478f
C24 drain_left.n9 a_n1564_n2088# 0.146498f
C25 drain_left.t9 a_n1564_n2088# 0.070869f
C26 drain_left.n10 a_n1564_n2088# 0.032611f
C27 drain_left.n11 a_n1564_n2088# 0.025684f
C28 drain_left.n12 a_n1564_n2088# 0.018396f
C29 drain_left.n13 a_n1564_n2088# 0.814567f
C30 drain_left.n14 a_n1564_n2088# 0.034234f
C31 drain_left.n15 a_n1564_n2088# 0.018396f
C32 drain_left.n16 a_n1564_n2088# 0.019478f
C33 drain_left.n17 a_n1564_n2088# 0.043481f
C34 drain_left.n18 a_n1564_n2088# 0.043481f
C35 drain_left.n19 a_n1564_n2088# 0.019478f
C36 drain_left.n20 a_n1564_n2088# 0.018396f
C37 drain_left.n21 a_n1564_n2088# 0.034234f
C38 drain_left.n22 a_n1564_n2088# 0.034234f
C39 drain_left.n23 a_n1564_n2088# 0.018396f
C40 drain_left.n24 a_n1564_n2088# 0.019478f
C41 drain_left.n25 a_n1564_n2088# 0.043481f
C42 drain_left.n26 a_n1564_n2088# 0.09413f
C43 drain_left.n27 a_n1564_n2088# 0.019478f
C44 drain_left.n28 a_n1564_n2088# 0.018396f
C45 drain_left.n29 a_n1564_n2088# 0.079131f
C46 drain_left.n30 a_n1564_n2088# 0.077385f
C47 drain_left.t11 a_n1564_n2088# 0.162317f
C48 drain_left.t5 a_n1564_n2088# 0.162317f
C49 drain_left.n31 a_n1564_n2088# 1.35372f
C50 drain_left.n32 a_n1564_n2088# 0.477956f
C51 drain_left.t3 a_n1564_n2088# 0.162317f
C52 drain_left.t4 a_n1564_n2088# 0.162317f
C53 drain_left.n33 a_n1564_n2088# 1.35637f
C54 drain_left.t10 a_n1564_n2088# 0.162317f
C55 drain_left.t6 a_n1564_n2088# 0.162317f
C56 drain_left.n34 a_n1564_n2088# 1.35372f
C57 drain_left.n35 a_n1564_n2088# 0.738025f
C58 drain_left.n36 a_n1564_n2088# 1.11595f
C59 drain_left.n37 a_n1564_n2088# 0.048119f
C60 drain_left.n38 a_n1564_n2088# 0.034234f
C61 drain_left.n39 a_n1564_n2088# 0.018396f
C62 drain_left.n40 a_n1564_n2088# 0.043481f
C63 drain_left.n41 a_n1564_n2088# 0.019478f
C64 drain_left.n42 a_n1564_n2088# 0.034234f
C65 drain_left.n43 a_n1564_n2088# 0.018396f
C66 drain_left.n44 a_n1564_n2088# 0.043481f
C67 drain_left.n45 a_n1564_n2088# 0.019478f
C68 drain_left.n46 a_n1564_n2088# 0.146498f
C69 drain_left.t7 a_n1564_n2088# 0.070869f
C70 drain_left.n47 a_n1564_n2088# 0.032611f
C71 drain_left.n48 a_n1564_n2088# 0.025684f
C72 drain_left.n49 a_n1564_n2088# 0.018396f
C73 drain_left.n50 a_n1564_n2088# 0.814567f
C74 drain_left.n51 a_n1564_n2088# 0.034234f
C75 drain_left.n52 a_n1564_n2088# 0.018396f
C76 drain_left.n53 a_n1564_n2088# 0.019478f
C77 drain_left.n54 a_n1564_n2088# 0.043481f
C78 drain_left.n55 a_n1564_n2088# 0.043481f
C79 drain_left.n56 a_n1564_n2088# 0.019478f
C80 drain_left.n57 a_n1564_n2088# 0.018396f
C81 drain_left.n58 a_n1564_n2088# 0.034234f
C82 drain_left.n59 a_n1564_n2088# 0.034234f
C83 drain_left.n60 a_n1564_n2088# 0.018396f
C84 drain_left.n61 a_n1564_n2088# 0.019478f
C85 drain_left.n62 a_n1564_n2088# 0.043481f
C86 drain_left.n63 a_n1564_n2088# 0.09413f
C87 drain_left.n64 a_n1564_n2088# 0.019478f
C88 drain_left.n65 a_n1564_n2088# 0.018396f
C89 drain_left.n66 a_n1564_n2088# 0.079131f
C90 drain_left.n67 a_n1564_n2088# 0.077385f
C91 drain_left.t12 a_n1564_n2088# 0.162317f
C92 drain_left.t0 a_n1564_n2088# 0.162317f
C93 drain_left.n68 a_n1564_n2088# 1.35373f
C94 drain_left.n69 a_n1564_n2088# 0.493893f
C95 drain_left.t1 a_n1564_n2088# 0.162317f
C96 drain_left.t2 a_n1564_n2088# 0.162317f
C97 drain_left.n70 a_n1564_n2088# 1.35373f
C98 drain_left.n71 a_n1564_n2088# 0.37865f
C99 drain_left.t8 a_n1564_n2088# 0.162317f
C100 drain_left.t13 a_n1564_n2088# 0.162317f
C101 drain_left.n72 a_n1564_n2088# 1.35372f
C102 drain_left.n73 a_n1564_n2088# 0.65883f
C103 plus.n0 a_n1564_n2088# 0.056404f
C104 plus.t5 a_n1564_n2088# 0.192847f
C105 plus.t11 a_n1564_n2088# 0.192847f
C106 plus.t12 a_n1564_n2088# 0.192847f
C107 plus.n1 a_n1564_n2088# 0.094316f
C108 plus.n2 a_n1564_n2088# 0.125942f
C109 plus.t13 a_n1564_n2088# 0.192847f
C110 plus.t1 a_n1564_n2088# 0.192847f
C111 plus.t6 a_n1564_n2088# 0.197961f
C112 plus.n3 a_n1564_n2088# 0.110429f
C113 plus.n4 a_n1564_n2088# 0.094316f
C114 plus.n5 a_n1564_n2088# 0.019754f
C115 plus.n6 a_n1564_n2088# 0.094316f
C116 plus.n7 a_n1564_n2088# 0.019754f
C117 plus.n8 a_n1564_n2088# 0.056404f
C118 plus.n9 a_n1564_n2088# 0.056404f
C119 plus.n10 a_n1564_n2088# 0.019754f
C120 plus.n11 a_n1564_n2088# 0.094316f
C121 plus.n12 a_n1564_n2088# 0.019754f
C122 plus.n13 a_n1564_n2088# 0.094316f
C123 plus.t0 a_n1564_n2088# 0.197961f
C124 plus.n14 a_n1564_n2088# 0.110347f
C125 plus.n15 a_n1564_n2088# 0.477875f
C126 plus.n16 a_n1564_n2088# 0.056404f
C127 plus.t4 a_n1564_n2088# 0.197961f
C128 plus.t2 a_n1564_n2088# 0.192847f
C129 plus.t8 a_n1564_n2088# 0.192847f
C130 plus.t3 a_n1564_n2088# 0.192847f
C131 plus.n17 a_n1564_n2088# 0.094316f
C132 plus.n18 a_n1564_n2088# 0.125942f
C133 plus.t7 a_n1564_n2088# 0.192847f
C134 plus.t10 a_n1564_n2088# 0.192847f
C135 plus.t9 a_n1564_n2088# 0.197961f
C136 plus.n19 a_n1564_n2088# 0.110429f
C137 plus.n20 a_n1564_n2088# 0.094316f
C138 plus.n21 a_n1564_n2088# 0.019754f
C139 plus.n22 a_n1564_n2088# 0.094316f
C140 plus.n23 a_n1564_n2088# 0.019754f
C141 plus.n24 a_n1564_n2088# 0.056404f
C142 plus.n25 a_n1564_n2088# 0.056404f
C143 plus.n26 a_n1564_n2088# 0.019754f
C144 plus.n27 a_n1564_n2088# 0.094316f
C145 plus.n28 a_n1564_n2088# 0.019754f
C146 plus.n29 a_n1564_n2088# 0.094316f
C147 plus.n30 a_n1564_n2088# 0.110347f
C148 plus.n31 a_n1564_n2088# 1.35847f
C149 drain_right.n0 a_n1564_n2088# 0.047962f
C150 drain_right.n1 a_n1564_n2088# 0.034123f
C151 drain_right.n2 a_n1564_n2088# 0.018336f
C152 drain_right.n3 a_n1564_n2088# 0.043339f
C153 drain_right.n4 a_n1564_n2088# 0.019414f
C154 drain_right.n5 a_n1564_n2088# 0.034123f
C155 drain_right.n6 a_n1564_n2088# 0.018336f
C156 drain_right.n7 a_n1564_n2088# 0.043339f
C157 drain_right.n8 a_n1564_n2088# 0.019414f
C158 drain_right.n9 a_n1564_n2088# 0.14602f
C159 drain_right.t4 a_n1564_n2088# 0.070638f
C160 drain_right.n10 a_n1564_n2088# 0.032505f
C161 drain_right.n11 a_n1564_n2088# 0.0256f
C162 drain_right.n12 a_n1564_n2088# 0.018336f
C163 drain_right.n13 a_n1564_n2088# 0.811911f
C164 drain_right.n14 a_n1564_n2088# 0.034123f
C165 drain_right.n15 a_n1564_n2088# 0.018336f
C166 drain_right.n16 a_n1564_n2088# 0.019414f
C167 drain_right.n17 a_n1564_n2088# 0.043339f
C168 drain_right.n18 a_n1564_n2088# 0.043339f
C169 drain_right.n19 a_n1564_n2088# 0.019414f
C170 drain_right.n20 a_n1564_n2088# 0.018336f
C171 drain_right.n21 a_n1564_n2088# 0.034123f
C172 drain_right.n22 a_n1564_n2088# 0.034123f
C173 drain_right.n23 a_n1564_n2088# 0.018336f
C174 drain_right.n24 a_n1564_n2088# 0.019414f
C175 drain_right.n25 a_n1564_n2088# 0.043339f
C176 drain_right.n26 a_n1564_n2088# 0.093823f
C177 drain_right.n27 a_n1564_n2088# 0.019414f
C178 drain_right.n28 a_n1564_n2088# 0.018336f
C179 drain_right.n29 a_n1564_n2088# 0.078873f
C180 drain_right.n30 a_n1564_n2088# 0.077132f
C181 drain_right.t1 a_n1564_n2088# 0.161788f
C182 drain_right.t5 a_n1564_n2088# 0.161788f
C183 drain_right.n31 a_n1564_n2088# 1.34931f
C184 drain_right.n32 a_n1564_n2088# 0.476398f
C185 drain_right.t0 a_n1564_n2088# 0.161788f
C186 drain_right.t13 a_n1564_n2088# 0.161788f
C187 drain_right.n33 a_n1564_n2088# 1.35195f
C188 drain_right.t2 a_n1564_n2088# 0.161788f
C189 drain_right.t10 a_n1564_n2088# 0.161788f
C190 drain_right.n34 a_n1564_n2088# 1.34931f
C191 drain_right.n35 a_n1564_n2088# 0.735619f
C192 drain_right.n36 a_n1564_n2088# 1.04272f
C193 drain_right.t8 a_n1564_n2088# 0.161788f
C194 drain_right.t7 a_n1564_n2088# 0.161788f
C195 drain_right.n37 a_n1564_n2088# 1.35195f
C196 drain_right.t3 a_n1564_n2088# 0.161788f
C197 drain_right.t12 a_n1564_n2088# 0.161788f
C198 drain_right.n38 a_n1564_n2088# 1.34932f
C199 drain_right.n39 a_n1564_n2088# 0.765939f
C200 drain_right.t9 a_n1564_n2088# 0.161788f
C201 drain_right.t6 a_n1564_n2088# 0.161788f
C202 drain_right.n40 a_n1564_n2088# 1.34932f
C203 drain_right.n41 a_n1564_n2088# 0.377415f
C204 drain_right.n42 a_n1564_n2088# 0.047962f
C205 drain_right.n43 a_n1564_n2088# 0.034123f
C206 drain_right.n44 a_n1564_n2088# 0.018336f
C207 drain_right.n45 a_n1564_n2088# 0.043339f
C208 drain_right.n46 a_n1564_n2088# 0.019414f
C209 drain_right.n47 a_n1564_n2088# 0.034123f
C210 drain_right.n48 a_n1564_n2088# 0.018336f
C211 drain_right.n49 a_n1564_n2088# 0.043339f
C212 drain_right.n50 a_n1564_n2088# 0.019414f
C213 drain_right.n51 a_n1564_n2088# 0.14602f
C214 drain_right.t11 a_n1564_n2088# 0.070638f
C215 drain_right.n52 a_n1564_n2088# 0.032505f
C216 drain_right.n53 a_n1564_n2088# 0.0256f
C217 drain_right.n54 a_n1564_n2088# 0.018336f
C218 drain_right.n55 a_n1564_n2088# 0.811911f
C219 drain_right.n56 a_n1564_n2088# 0.034123f
C220 drain_right.n57 a_n1564_n2088# 0.018336f
C221 drain_right.n58 a_n1564_n2088# 0.019414f
C222 drain_right.n59 a_n1564_n2088# 0.043339f
C223 drain_right.n60 a_n1564_n2088# 0.043339f
C224 drain_right.n61 a_n1564_n2088# 0.019414f
C225 drain_right.n62 a_n1564_n2088# 0.018336f
C226 drain_right.n63 a_n1564_n2088# 0.034123f
C227 drain_right.n64 a_n1564_n2088# 0.034123f
C228 drain_right.n65 a_n1564_n2088# 0.018336f
C229 drain_right.n66 a_n1564_n2088# 0.019414f
C230 drain_right.n67 a_n1564_n2088# 0.043339f
C231 drain_right.n68 a_n1564_n2088# 0.093823f
C232 drain_right.n69 a_n1564_n2088# 0.019414f
C233 drain_right.n70 a_n1564_n2088# 0.018336f
C234 drain_right.n71 a_n1564_n2088# 0.078873f
C235 drain_right.n72 a_n1564_n2088# 0.076058f
C236 drain_right.n73 a_n1564_n2088# 0.393281f
C237 source.n0 a_n1564_n2088# 0.051704f
C238 source.n1 a_n1564_n2088# 0.036784f
C239 source.n2 a_n1564_n2088# 0.019766f
C240 source.n3 a_n1564_n2088# 0.046721f
C241 source.n4 a_n1564_n2088# 0.020929f
C242 source.n5 a_n1564_n2088# 0.036784f
C243 source.n6 a_n1564_n2088# 0.019766f
C244 source.n7 a_n1564_n2088# 0.046721f
C245 source.n8 a_n1564_n2088# 0.020929f
C246 source.n9 a_n1564_n2088# 0.157412f
C247 source.t8 a_n1564_n2088# 0.076149f
C248 source.n10 a_n1564_n2088# 0.03504f
C249 source.n11 a_n1564_n2088# 0.027597f
C250 source.n12 a_n1564_n2088# 0.019766f
C251 source.n13 a_n1564_n2088# 0.875252f
C252 source.n14 a_n1564_n2088# 0.036784f
C253 source.n15 a_n1564_n2088# 0.019766f
C254 source.n16 a_n1564_n2088# 0.020929f
C255 source.n17 a_n1564_n2088# 0.046721f
C256 source.n18 a_n1564_n2088# 0.046721f
C257 source.n19 a_n1564_n2088# 0.020929f
C258 source.n20 a_n1564_n2088# 0.019766f
C259 source.n21 a_n1564_n2088# 0.036784f
C260 source.n22 a_n1564_n2088# 0.036784f
C261 source.n23 a_n1564_n2088# 0.019766f
C262 source.n24 a_n1564_n2088# 0.020929f
C263 source.n25 a_n1564_n2088# 0.046721f
C264 source.n26 a_n1564_n2088# 0.101142f
C265 source.n27 a_n1564_n2088# 0.020929f
C266 source.n28 a_n1564_n2088# 0.019766f
C267 source.n29 a_n1564_n2088# 0.085026f
C268 source.n30 a_n1564_n2088# 0.056593f
C269 source.n31 a_n1564_n2088# 0.873468f
C270 source.t5 a_n1564_n2088# 0.174409f
C271 source.t2 a_n1564_n2088# 0.174409f
C272 source.n32 a_n1564_n2088# 1.35832f
C273 source.n33 a_n1564_n2088# 0.45313f
C274 source.t12 a_n1564_n2088# 0.174409f
C275 source.t11 a_n1564_n2088# 0.174409f
C276 source.n34 a_n1564_n2088# 1.35832f
C277 source.n35 a_n1564_n2088# 0.45313f
C278 source.t4 a_n1564_n2088# 0.174409f
C279 source.t0 a_n1564_n2088# 0.174409f
C280 source.n36 a_n1564_n2088# 1.35832f
C281 source.n37 a_n1564_n2088# 0.48174f
C282 source.n38 a_n1564_n2088# 0.051704f
C283 source.n39 a_n1564_n2088# 0.036784f
C284 source.n40 a_n1564_n2088# 0.019766f
C285 source.n41 a_n1564_n2088# 0.046721f
C286 source.n42 a_n1564_n2088# 0.020929f
C287 source.n43 a_n1564_n2088# 0.036784f
C288 source.n44 a_n1564_n2088# 0.019766f
C289 source.n45 a_n1564_n2088# 0.046721f
C290 source.n46 a_n1564_n2088# 0.020929f
C291 source.n47 a_n1564_n2088# 0.157412f
C292 source.t20 a_n1564_n2088# 0.076149f
C293 source.n48 a_n1564_n2088# 0.03504f
C294 source.n49 a_n1564_n2088# 0.027597f
C295 source.n50 a_n1564_n2088# 0.019766f
C296 source.n51 a_n1564_n2088# 0.875252f
C297 source.n52 a_n1564_n2088# 0.036784f
C298 source.n53 a_n1564_n2088# 0.019766f
C299 source.n54 a_n1564_n2088# 0.020929f
C300 source.n55 a_n1564_n2088# 0.046721f
C301 source.n56 a_n1564_n2088# 0.046721f
C302 source.n57 a_n1564_n2088# 0.020929f
C303 source.n58 a_n1564_n2088# 0.019766f
C304 source.n59 a_n1564_n2088# 0.036784f
C305 source.n60 a_n1564_n2088# 0.036784f
C306 source.n61 a_n1564_n2088# 0.019766f
C307 source.n62 a_n1564_n2088# 0.020929f
C308 source.n63 a_n1564_n2088# 0.046721f
C309 source.n64 a_n1564_n2088# 0.101142f
C310 source.n65 a_n1564_n2088# 0.020929f
C311 source.n66 a_n1564_n2088# 0.019766f
C312 source.n67 a_n1564_n2088# 0.085026f
C313 source.n68 a_n1564_n2088# 0.056593f
C314 source.n69 a_n1564_n2088# 0.168337f
C315 source.t15 a_n1564_n2088# 0.174409f
C316 source.t19 a_n1564_n2088# 0.174409f
C317 source.n70 a_n1564_n2088# 1.35832f
C318 source.n71 a_n1564_n2088# 0.45313f
C319 source.t24 a_n1564_n2088# 0.174409f
C320 source.t26 a_n1564_n2088# 0.174409f
C321 source.n72 a_n1564_n2088# 1.35832f
C322 source.n73 a_n1564_n2088# 0.45313f
C323 source.t16 a_n1564_n2088# 0.174409f
C324 source.t18 a_n1564_n2088# 0.174409f
C325 source.n74 a_n1564_n2088# 1.35832f
C326 source.n75 a_n1564_n2088# 1.71168f
C327 source.t1 a_n1564_n2088# 0.174409f
C328 source.t10 a_n1564_n2088# 0.174409f
C329 source.n76 a_n1564_n2088# 1.35831f
C330 source.n77 a_n1564_n2088# 1.71169f
C331 source.t9 a_n1564_n2088# 0.174409f
C332 source.t3 a_n1564_n2088# 0.174409f
C333 source.n78 a_n1564_n2088# 1.35831f
C334 source.n79 a_n1564_n2088# 0.453139f
C335 source.t6 a_n1564_n2088# 0.174409f
C336 source.t13 a_n1564_n2088# 0.174409f
C337 source.n80 a_n1564_n2088# 1.35831f
C338 source.n81 a_n1564_n2088# 0.453139f
C339 source.n82 a_n1564_n2088# 0.051704f
C340 source.n83 a_n1564_n2088# 0.036784f
C341 source.n84 a_n1564_n2088# 0.019766f
C342 source.n85 a_n1564_n2088# 0.046721f
C343 source.n86 a_n1564_n2088# 0.020929f
C344 source.n87 a_n1564_n2088# 0.036784f
C345 source.n88 a_n1564_n2088# 0.019766f
C346 source.n89 a_n1564_n2088# 0.046721f
C347 source.n90 a_n1564_n2088# 0.020929f
C348 source.n91 a_n1564_n2088# 0.157412f
C349 source.t7 a_n1564_n2088# 0.076149f
C350 source.n92 a_n1564_n2088# 0.03504f
C351 source.n93 a_n1564_n2088# 0.027597f
C352 source.n94 a_n1564_n2088# 0.019766f
C353 source.n95 a_n1564_n2088# 0.875252f
C354 source.n96 a_n1564_n2088# 0.036784f
C355 source.n97 a_n1564_n2088# 0.019766f
C356 source.n98 a_n1564_n2088# 0.020929f
C357 source.n99 a_n1564_n2088# 0.046721f
C358 source.n100 a_n1564_n2088# 0.046721f
C359 source.n101 a_n1564_n2088# 0.020929f
C360 source.n102 a_n1564_n2088# 0.019766f
C361 source.n103 a_n1564_n2088# 0.036784f
C362 source.n104 a_n1564_n2088# 0.036784f
C363 source.n105 a_n1564_n2088# 0.019766f
C364 source.n106 a_n1564_n2088# 0.020929f
C365 source.n107 a_n1564_n2088# 0.046721f
C366 source.n108 a_n1564_n2088# 0.101142f
C367 source.n109 a_n1564_n2088# 0.020929f
C368 source.n110 a_n1564_n2088# 0.019766f
C369 source.n111 a_n1564_n2088# 0.085026f
C370 source.n112 a_n1564_n2088# 0.056593f
C371 source.n113 a_n1564_n2088# 0.168337f
C372 source.t21 a_n1564_n2088# 0.174409f
C373 source.t23 a_n1564_n2088# 0.174409f
C374 source.n114 a_n1564_n2088# 1.35831f
C375 source.n115 a_n1564_n2088# 0.481749f
C376 source.t25 a_n1564_n2088# 0.174409f
C377 source.t22 a_n1564_n2088# 0.174409f
C378 source.n116 a_n1564_n2088# 1.35831f
C379 source.n117 a_n1564_n2088# 0.453139f
C380 source.t17 a_n1564_n2088# 0.174409f
C381 source.t27 a_n1564_n2088# 0.174409f
C382 source.n118 a_n1564_n2088# 1.35831f
C383 source.n119 a_n1564_n2088# 0.453139f
C384 source.n120 a_n1564_n2088# 0.051704f
C385 source.n121 a_n1564_n2088# 0.036784f
C386 source.n122 a_n1564_n2088# 0.019766f
C387 source.n123 a_n1564_n2088# 0.046721f
C388 source.n124 a_n1564_n2088# 0.020929f
C389 source.n125 a_n1564_n2088# 0.036784f
C390 source.n126 a_n1564_n2088# 0.019766f
C391 source.n127 a_n1564_n2088# 0.046721f
C392 source.n128 a_n1564_n2088# 0.020929f
C393 source.n129 a_n1564_n2088# 0.157412f
C394 source.t14 a_n1564_n2088# 0.076149f
C395 source.n130 a_n1564_n2088# 0.03504f
C396 source.n131 a_n1564_n2088# 0.027597f
C397 source.n132 a_n1564_n2088# 0.019766f
C398 source.n133 a_n1564_n2088# 0.875252f
C399 source.n134 a_n1564_n2088# 0.036784f
C400 source.n135 a_n1564_n2088# 0.019766f
C401 source.n136 a_n1564_n2088# 0.020929f
C402 source.n137 a_n1564_n2088# 0.046721f
C403 source.n138 a_n1564_n2088# 0.046721f
C404 source.n139 a_n1564_n2088# 0.020929f
C405 source.n140 a_n1564_n2088# 0.019766f
C406 source.n141 a_n1564_n2088# 0.036784f
C407 source.n142 a_n1564_n2088# 0.036784f
C408 source.n143 a_n1564_n2088# 0.019766f
C409 source.n144 a_n1564_n2088# 0.020929f
C410 source.n145 a_n1564_n2088# 0.046721f
C411 source.n146 a_n1564_n2088# 0.101142f
C412 source.n147 a_n1564_n2088# 0.020929f
C413 source.n148 a_n1564_n2088# 0.019766f
C414 source.n149 a_n1564_n2088# 0.085026f
C415 source.n150 a_n1564_n2088# 0.056593f
C416 source.n151 a_n1564_n2088# 0.340717f
C417 source.n152 a_n1564_n2088# 1.50022f
C418 minus.n0 a_n1564_n2088# 0.054348f
C419 minus.t2 a_n1564_n2088# 0.190744f
C420 minus.t4 a_n1564_n2088# 0.185816f
C421 minus.t7 a_n1564_n2088# 0.185816f
C422 minus.t10 a_n1564_n2088# 0.185816f
C423 minus.n1 a_n1564_n2088# 0.090877f
C424 minus.n2 a_n1564_n2088# 0.12135f
C425 minus.t1 a_n1564_n2088# 0.185816f
C426 minus.t5 a_n1564_n2088# 0.185816f
C427 minus.t6 a_n1564_n2088# 0.190744f
C428 minus.n3 a_n1564_n2088# 0.106402f
C429 minus.n4 a_n1564_n2088# 0.090877f
C430 minus.n5 a_n1564_n2088# 0.019034f
C431 minus.n6 a_n1564_n2088# 0.090877f
C432 minus.n7 a_n1564_n2088# 0.019034f
C433 minus.n8 a_n1564_n2088# 0.054348f
C434 minus.n9 a_n1564_n2088# 0.054348f
C435 minus.n10 a_n1564_n2088# 0.019034f
C436 minus.n11 a_n1564_n2088# 0.090877f
C437 minus.n12 a_n1564_n2088# 0.019034f
C438 minus.n13 a_n1564_n2088# 0.090877f
C439 minus.n14 a_n1564_n2088# 0.106324f
C440 minus.n15 a_n1564_n2088# 1.44899f
C441 minus.n16 a_n1564_n2088# 0.054348f
C442 minus.t13 a_n1564_n2088# 0.185816f
C443 minus.t3 a_n1564_n2088# 0.185816f
C444 minus.t11 a_n1564_n2088# 0.185816f
C445 minus.n17 a_n1564_n2088# 0.090877f
C446 minus.n18 a_n1564_n2088# 0.12135f
C447 minus.t8 a_n1564_n2088# 0.185816f
C448 minus.t12 a_n1564_n2088# 0.185816f
C449 minus.t9 a_n1564_n2088# 0.190744f
C450 minus.n19 a_n1564_n2088# 0.106402f
C451 minus.n20 a_n1564_n2088# 0.090877f
C452 minus.n21 a_n1564_n2088# 0.019034f
C453 minus.n22 a_n1564_n2088# 0.090877f
C454 minus.n23 a_n1564_n2088# 0.019034f
C455 minus.n24 a_n1564_n2088# 0.054348f
C456 minus.n25 a_n1564_n2088# 0.054348f
C457 minus.n26 a_n1564_n2088# 0.019034f
C458 minus.n27 a_n1564_n2088# 0.090877f
C459 minus.n28 a_n1564_n2088# 0.019034f
C460 minus.n29 a_n1564_n2088# 0.090877f
C461 minus.t0 a_n1564_n2088# 0.190744f
C462 minus.n30 a_n1564_n2088# 0.106324f
C463 minus.n31 a_n1564_n2088# 0.350274f
C464 minus.n32 a_n1564_n2088# 1.78863f
.ends

