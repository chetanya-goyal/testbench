* NGSPICE file created from diffpair523.ext - technology: sky130A

.subckt diffpair523 minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t1 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X1 drain_left.t2 plus.t1 source.t14 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X2 source.t6 minus.t0 drain_right.t7 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X3 source.t13 plus.t2 drain_left.t3 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X4 source.t12 plus.t3 drain_left.t4 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X5 drain_right.t6 minus.t1 source.t4 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X6 source.t5 minus.t2 drain_right.t5 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X7 a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.5
X8 a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X9 drain_right.t4 minus.t3 source.t2 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X10 drain_left.t5 plus.t4 source.t11 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X11 drain_left.t6 plus.t5 source.t10 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X12 drain_right.t3 minus.t4 source.t3 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X13 drain_right.t2 minus.t5 source.t7 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.5
X14 source.t1 minus.t6 drain_right.t1 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X15 drain_left.t0 plus.t6 source.t9 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X16 source.t0 minus.t7 drain_right.t0 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.5
X17 a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
X18 source.t8 plus.t7 drain_left.t7 a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.5
X19 a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# a_n1546_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.5
R0 plus.n2 plus.t2 822.548
R1 plus.n10 plus.t1 822.548
R2 plus.n6 plus.t4 801.567
R3 plus.n5 plus.t7 801.567
R4 plus.n1 plus.t6 801.567
R5 plus.n14 plus.t3 801.567
R6 plus.n13 plus.t5 801.567
R7 plus.n9 plus.t0 801.567
R8 plus.n4 plus.n3 161.3
R9 plus.n5 plus.n0 161.3
R10 plus.n7 plus.n6 161.3
R11 plus.n12 plus.n11 161.3
R12 plus.n13 plus.n8 161.3
R13 plus.n15 plus.n14 161.3
R14 plus.n3 plus.n2 70.4033
R15 plus.n11 plus.n10 70.4033
R16 plus.n6 plus.n5 48.2005
R17 plus.n14 plus.n13 48.2005
R18 plus plus.n15 30.0899
R19 plus.n4 plus.n1 24.1005
R20 plus.n5 plus.n4 24.1005
R21 plus.n13 plus.n12 24.1005
R22 plus.n12 plus.n9 24.1005
R23 plus.n2 plus.n1 20.9576
R24 plus.n10 plus.n9 20.9576
R25 plus plus.n7 13.3755
R26 plus.n3 plus.n0 0.189894
R27 plus.n7 plus.n0 0.189894
R28 plus.n15 plus.n8 0.189894
R29 plus.n11 plus.n8 0.189894
R30 drain_left.n5 drain_left.n3 61.5953
R31 drain_left.n2 drain_left.n1 61.182
R32 drain_left.n2 drain_left.n0 61.182
R33 drain_left.n5 drain_left.n4 60.8796
R34 drain_left drain_left.n2 32.1441
R35 drain_left drain_left.n5 6.36873
R36 drain_left.n1 drain_left.t1 1.3205
R37 drain_left.n1 drain_left.t2 1.3205
R38 drain_left.n0 drain_left.t4 1.3205
R39 drain_left.n0 drain_left.t6 1.3205
R40 drain_left.n4 drain_left.t7 1.3205
R41 drain_left.n4 drain_left.t5 1.3205
R42 drain_left.n3 drain_left.t3 1.3205
R43 drain_left.n3 drain_left.t0 1.3205
R44 source.n3 source.t13 45.521
R45 source.n4 source.t3 45.521
R46 source.n7 source.t0 45.521
R47 source.n15 source.t7 45.5208
R48 source.n12 source.t5 45.5208
R49 source.n11 source.t14 45.5208
R50 source.n8 source.t12 45.5208
R51 source.n0 source.t11 45.5208
R52 source.n2 source.n1 44.201
R53 source.n6 source.n5 44.201
R54 source.n14 source.n13 44.2008
R55 source.n10 source.n9 44.2008
R56 source.n8 source.n7 24.276
R57 source.n16 source.n0 18.6553
R58 source.n16 source.n15 5.62119
R59 source.n13 source.t4 1.3205
R60 source.n13 source.t1 1.3205
R61 source.n9 source.t10 1.3205
R62 source.n9 source.t15 1.3205
R63 source.n1 source.t9 1.3205
R64 source.n1 source.t8 1.3205
R65 source.n5 source.t2 1.3205
R66 source.n5 source.t6 1.3205
R67 source.n7 source.n6 0.716017
R68 source.n6 source.n4 0.716017
R69 source.n3 source.n2 0.716017
R70 source.n2 source.n0 0.716017
R71 source.n10 source.n8 0.716017
R72 source.n11 source.n10 0.716017
R73 source.n14 source.n12 0.716017
R74 source.n15 source.n14 0.716017
R75 source.n4 source.n3 0.470328
R76 source.n12 source.n11 0.470328
R77 source source.n16 0.188
R78 minus.n2 minus.t4 822.548
R79 minus.n10 minus.t2 822.548
R80 minus.n1 minus.t0 801.567
R81 minus.n5 minus.t3 801.567
R82 minus.n6 minus.t7 801.567
R83 minus.n9 minus.t1 801.567
R84 minus.n13 minus.t6 801.567
R85 minus.n14 minus.t5 801.567
R86 minus.n7 minus.n6 161.3
R87 minus.n5 minus.n0 161.3
R88 minus.n4 minus.n3 161.3
R89 minus.n15 minus.n14 161.3
R90 minus.n13 minus.n8 161.3
R91 minus.n12 minus.n11 161.3
R92 minus.n3 minus.n2 70.4033
R93 minus.n11 minus.n10 70.4033
R94 minus.n6 minus.n5 48.2005
R95 minus.n14 minus.n13 48.2005
R96 minus.n16 minus.n7 37.3452
R97 minus.n5 minus.n4 24.1005
R98 minus.n4 minus.n1 24.1005
R99 minus.n12 minus.n9 24.1005
R100 minus.n13 minus.n12 24.1005
R101 minus.n2 minus.n1 20.9576
R102 minus.n10 minus.n9 20.9576
R103 minus.n16 minus.n15 6.5952
R104 minus.n7 minus.n0 0.189894
R105 minus.n3 minus.n0 0.189894
R106 minus.n11 minus.n8 0.189894
R107 minus.n15 minus.n8 0.189894
R108 minus minus.n16 0.188
R109 drain_right.n5 drain_right.n3 61.5952
R110 drain_right.n2 drain_right.n1 61.182
R111 drain_right.n2 drain_right.n0 61.182
R112 drain_right.n5 drain_right.n4 60.8798
R113 drain_right drain_right.n2 31.5909
R114 drain_right drain_right.n5 6.36873
R115 drain_right.n1 drain_right.t1 1.3205
R116 drain_right.n1 drain_right.t2 1.3205
R117 drain_right.n0 drain_right.t5 1.3205
R118 drain_right.n0 drain_right.t6 1.3205
R119 drain_right.n3 drain_right.t7 1.3205
R120 drain_right.n3 drain_right.t3 1.3205
R121 drain_right.n4 drain_right.t0 1.3205
R122 drain_right.n4 drain_right.t4 1.3205
C0 source drain_right 15.865f
C1 source plus 5.21019f
C2 minus drain_left 0.171215f
C3 drain_right drain_left 0.727126f
C4 drain_left plus 5.79114f
C5 source drain_left 15.8645f
C6 minus drain_right 5.64311f
C7 minus plus 5.62723f
C8 source minus 5.19615f
C9 drain_right plus 0.302201f
C10 drain_right a_n1546_n3888# 6.220809f
C11 drain_left a_n1546_n3888# 6.46385f
C12 source a_n1546_n3888# 10.433959f
C13 minus a_n1546_n3888# 6.163311f
C14 plus a_n1546_n3888# 8.18359f
C15 drain_right.t5 a_n1546_n3888# 0.344914f
C16 drain_right.t6 a_n1546_n3888# 0.344914f
C17 drain_right.n0 a_n1546_n3888# 3.11934f
C18 drain_right.t1 a_n1546_n3888# 0.344914f
C19 drain_right.t2 a_n1546_n3888# 0.344914f
C20 drain_right.n1 a_n1546_n3888# 3.11934f
C21 drain_right.n2 a_n1546_n3888# 2.18662f
C22 drain_right.t7 a_n1546_n3888# 0.344914f
C23 drain_right.t3 a_n1546_n3888# 0.344914f
C24 drain_right.n3 a_n1546_n3888# 3.12207f
C25 drain_right.t0 a_n1546_n3888# 0.344914f
C26 drain_right.t4 a_n1546_n3888# 0.344914f
C27 drain_right.n4 a_n1546_n3888# 3.11762f
C28 drain_right.n5 a_n1546_n3888# 1.00227f
C29 minus.n0 a_n1546_n3888# 0.048822f
C30 minus.t0 a_n1546_n3888# 1.04054f
C31 minus.n1 a_n1546_n3888# 0.410324f
C32 minus.t4 a_n1546_n3888# 1.05088f
C33 minus.n2 a_n1546_n3888# 0.395392f
C34 minus.n3 a_n1546_n3888# 0.16084f
C35 minus.n4 a_n1546_n3888# 0.011079f
C36 minus.t3 a_n1546_n3888# 1.04054f
C37 minus.n5 a_n1546_n3888# 0.410324f
C38 minus.t7 a_n1546_n3888# 1.04054f
C39 minus.n6 a_n1546_n3888# 0.405357f
C40 minus.n7 a_n1546_n3888# 1.81491f
C41 minus.n8 a_n1546_n3888# 0.048822f
C42 minus.t1 a_n1546_n3888# 1.04054f
C43 minus.n9 a_n1546_n3888# 0.410324f
C44 minus.t2 a_n1546_n3888# 1.05088f
C45 minus.n10 a_n1546_n3888# 0.395392f
C46 minus.n11 a_n1546_n3888# 0.16084f
C47 minus.n12 a_n1546_n3888# 0.011079f
C48 minus.t6 a_n1546_n3888# 1.04054f
C49 minus.n13 a_n1546_n3888# 0.410324f
C50 minus.t5 a_n1546_n3888# 1.04054f
C51 minus.n14 a_n1546_n3888# 0.405357f
C52 minus.n15 a_n1546_n3888# 0.330089f
C53 minus.n16 a_n1546_n3888# 2.19366f
C54 source.t11 a_n1546_n3888# 2.7745f
C55 source.n0 a_n1546_n3888# 1.3038f
C56 source.t9 a_n1546_n3888# 0.247577f
C57 source.t8 a_n1546_n3888# 0.247577f
C58 source.n1 a_n1546_n3888# 2.17476f
C59 source.n2 a_n1546_n3888# 0.302045f
C60 source.t13 a_n1546_n3888# 2.7745f
C61 source.n3 a_n1546_n3888# 0.360973f
C62 source.t3 a_n1546_n3888# 2.7745f
C63 source.n4 a_n1546_n3888# 0.360973f
C64 source.t2 a_n1546_n3888# 0.247577f
C65 source.t6 a_n1546_n3888# 0.247577f
C66 source.n5 a_n1546_n3888# 2.17476f
C67 source.n6 a_n1546_n3888# 0.302045f
C68 source.t0 a_n1546_n3888# 2.7745f
C69 source.n7 a_n1546_n3888# 1.65556f
C70 source.t12 a_n1546_n3888# 2.7745f
C71 source.n8 a_n1546_n3888# 1.65556f
C72 source.t10 a_n1546_n3888# 0.247577f
C73 source.t15 a_n1546_n3888# 0.247577f
C74 source.n9 a_n1546_n3888# 2.17475f
C75 source.n10 a_n1546_n3888# 0.302047f
C76 source.t14 a_n1546_n3888# 2.7745f
C77 source.n11 a_n1546_n3888# 0.360977f
C78 source.t5 a_n1546_n3888# 2.7745f
C79 source.n12 a_n1546_n3888# 0.360977f
C80 source.t4 a_n1546_n3888# 0.247577f
C81 source.t1 a_n1546_n3888# 0.247577f
C82 source.n13 a_n1546_n3888# 2.17475f
C83 source.n14 a_n1546_n3888# 0.302047f
C84 source.t7 a_n1546_n3888# 2.7745f
C85 source.n15 a_n1546_n3888# 0.488102f
C86 source.n16 a_n1546_n3888# 1.53407f
C87 drain_left.t4 a_n1546_n3888# 0.346289f
C88 drain_left.t6 a_n1546_n3888# 0.346289f
C89 drain_left.n0 a_n1546_n3888# 3.13177f
C90 drain_left.t1 a_n1546_n3888# 0.346289f
C91 drain_left.t2 a_n1546_n3888# 0.346289f
C92 drain_left.n1 a_n1546_n3888# 3.13177f
C93 drain_left.n2 a_n1546_n3888# 2.25647f
C94 drain_left.t3 a_n1546_n3888# 0.346289f
C95 drain_left.t0 a_n1546_n3888# 0.346289f
C96 drain_left.n3 a_n1546_n3888# 3.13453f
C97 drain_left.t7 a_n1546_n3888# 0.346289f
C98 drain_left.t5 a_n1546_n3888# 0.346289f
C99 drain_left.n4 a_n1546_n3888# 3.13004f
C100 drain_left.n5 a_n1546_n3888# 1.00627f
C101 plus.n0 a_n1546_n3888# 0.049717f
C102 plus.t4 a_n1546_n3888# 1.05961f
C103 plus.t7 a_n1546_n3888# 1.05961f
C104 plus.t6 a_n1546_n3888# 1.05961f
C105 plus.n1 a_n1546_n3888# 0.417843f
C106 plus.t2 a_n1546_n3888# 1.07014f
C107 plus.n2 a_n1546_n3888# 0.402638f
C108 plus.n3 a_n1546_n3888# 0.163787f
C109 plus.n4 a_n1546_n3888# 0.011282f
C110 plus.n5 a_n1546_n3888# 0.417843f
C111 plus.n6 a_n1546_n3888# 0.412786f
C112 plus.n7 a_n1546_n3888# 0.639392f
C113 plus.n8 a_n1546_n3888# 0.049717f
C114 plus.t3 a_n1546_n3888# 1.05961f
C115 plus.t5 a_n1546_n3888# 1.05961f
C116 plus.t0 a_n1546_n3888# 1.05961f
C117 plus.n9 a_n1546_n3888# 0.417843f
C118 plus.t1 a_n1546_n3888# 1.07014f
C119 plus.n10 a_n1546_n3888# 0.402638f
C120 plus.n11 a_n1546_n3888# 0.163787f
C121 plus.n12 a_n1546_n3888# 0.011282f
C122 plus.n13 a_n1546_n3888# 0.417843f
C123 plus.n14 a_n1546_n3888# 0.412786f
C124 plus.n15 a_n1546_n3888# 1.5176f
.ends

