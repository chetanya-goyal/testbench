* NGSPICE file created from diffpair375.ext - technology: sky130A

.subckt diffpair375 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t16 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X1 source.t3 minus.t0 drain_right.t11 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X2 drain_right.t10 minus.t1 source.t22 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X3 source.t12 plus.t1 drain_left.t10 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 source.t20 minus.t2 drain_right.t9 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X6 source.t7 minus.t3 drain_right.t8 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X7 a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X8 source.t15 plus.t2 drain_left.t9 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X9 drain_left.t8 plus.t3 source.t8 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 source.t0 minus.t4 drain_right.t7 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 drain_right.t6 minus.t5 source.t23 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X12 drain_left.t7 plus.t4 source.t17 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X13 source.t2 minus.t6 drain_right.t5 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X14 source.t18 plus.t5 drain_left.t6 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X15 drain_right.t4 minus.t7 source.t1 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X16 a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X17 drain_left.t5 plus.t6 source.t10 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X18 source.t9 plus.t7 drain_left.t4 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X19 drain_right.t3 minus.t8 source.t21 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X20 drain_left.t3 plus.t8 source.t19 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X21 source.t13 plus.t9 drain_left.t2 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X22 a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X23 drain_right.t2 minus.t9 source.t4 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X24 drain_left.t1 plus.t10 source.t11 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X25 source.t5 minus.t10 drain_right.t1 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X26 drain_right.t0 minus.t11 source.t6 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X27 source.t14 plus.t11 drain_left.t0 a_n2018_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
R0 plus.n4 plus.t7 452.031
R1 plus.n16 plus.t8 452.031
R2 plus.n10 plus.t0 426.973
R3 plus.n8 plus.t2 426.973
R4 plus.n7 plus.t4 426.973
R5 plus.n6 plus.t5 426.973
R6 plus.n5 plus.t6 426.973
R7 plus.n22 plus.t11 426.973
R8 plus.n20 plus.t10 426.973
R9 plus.n19 plus.t9 426.973
R10 plus.n18 plus.t3 426.973
R11 plus.n17 plus.t1 426.973
R12 plus.n8 plus.n1 161.3
R13 plus.n9 plus.n0 161.3
R14 plus.n11 plus.n10 161.3
R15 plus.n20 plus.n13 161.3
R16 plus.n21 plus.n12 161.3
R17 plus.n23 plus.n22 161.3
R18 plus.n6 plus.n3 80.6037
R19 plus.n7 plus.n2 80.6037
R20 plus.n18 plus.n15 80.6037
R21 plus.n19 plus.n14 80.6037
R22 plus.n8 plus.n7 48.2005
R23 plus.n7 plus.n6 48.2005
R24 plus.n6 plus.n5 48.2005
R25 plus.n20 plus.n19 48.2005
R26 plus.n19 plus.n18 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n4 plus.n3 45.0744
R29 plus.n16 plus.n15 45.0744
R30 plus.n10 plus.n9 40.1672
R31 plus.n22 plus.n21 40.1672
R32 plus plus.n23 29.5975
R33 plus.n5 plus.n4 16.1124
R34 plus.n17 plus.n16 16.1124
R35 plus plus.n11 11.0952
R36 plus.n9 plus.n8 8.03383
R37 plus.n21 plus.n20 8.03383
R38 plus.n3 plus.n2 0.380177
R39 plus.n15 plus.n14 0.380177
R40 plus.n2 plus.n1 0.285035
R41 plus.n14 plus.n13 0.285035
R42 plus.n1 plus.n0 0.189894
R43 plus.n11 plus.n0 0.189894
R44 plus.n23 plus.n12 0.189894
R45 plus.n13 plus.n12 0.189894
R46 source.n5 source.t9 51.0588
R47 source.n6 source.t1 51.0588
R48 source.n11 source.t20 51.0588
R49 source.n23 source.t4 51.0586
R50 source.n18 source.t7 51.0586
R51 source.n17 source.t19 51.0586
R52 source.n12 source.t14 51.0586
R53 source.n0 source.t16 51.0586
R54 source.n2 source.n1 48.8588
R55 source.n4 source.n3 48.8588
R56 source.n8 source.n7 48.8588
R57 source.n10 source.n9 48.8588
R58 source.n22 source.n21 48.8586
R59 source.n20 source.n19 48.8586
R60 source.n16 source.n15 48.8586
R61 source.n14 source.n13 48.8586
R62 source.n12 source.n11 19.8167
R63 source.n24 source.n0 14.1529
R64 source.n24 source.n23 5.66429
R65 source.n21 source.t21 2.2005
R66 source.n21 source.t5 2.2005
R67 source.n19 source.t6 2.2005
R68 source.n19 source.t3 2.2005
R69 source.n15 source.t8 2.2005
R70 source.n15 source.t12 2.2005
R71 source.n13 source.t11 2.2005
R72 source.n13 source.t13 2.2005
R73 source.n1 source.t17 2.2005
R74 source.n1 source.t15 2.2005
R75 source.n3 source.t10 2.2005
R76 source.n3 source.t18 2.2005
R77 source.n7 source.t23 2.2005
R78 source.n7 source.t2 2.2005
R79 source.n9 source.t22 2.2005
R80 source.n9 source.t0 2.2005
R81 source.n11 source.n10 0.802224
R82 source.n10 source.n8 0.802224
R83 source.n8 source.n6 0.802224
R84 source.n5 source.n4 0.802224
R85 source.n4 source.n2 0.802224
R86 source.n2 source.n0 0.802224
R87 source.n14 source.n12 0.802224
R88 source.n16 source.n14 0.802224
R89 source.n17 source.n16 0.802224
R90 source.n20 source.n18 0.802224
R91 source.n22 source.n20 0.802224
R92 source.n23 source.n22 0.802224
R93 source.n6 source.n5 0.470328
R94 source.n18 source.n17 0.470328
R95 source source.n24 0.188
R96 drain_left.n6 drain_left.n4 66.3393
R97 drain_left.n3 drain_left.n2 66.2837
R98 drain_left.n3 drain_left.n0 66.2837
R99 drain_left.n6 drain_left.n5 65.5376
R100 drain_left.n8 drain_left.n7 65.5374
R101 drain_left.n3 drain_left.n1 65.5373
R102 drain_left drain_left.n3 29.103
R103 drain_left drain_left.n8 6.45494
R104 drain_left.n1 drain_left.t2 2.2005
R105 drain_left.n1 drain_left.t8 2.2005
R106 drain_left.n2 drain_left.t10 2.2005
R107 drain_left.n2 drain_left.t3 2.2005
R108 drain_left.n0 drain_left.t0 2.2005
R109 drain_left.n0 drain_left.t1 2.2005
R110 drain_left.n7 drain_left.t9 2.2005
R111 drain_left.n7 drain_left.t11 2.2005
R112 drain_left.n5 drain_left.t6 2.2005
R113 drain_left.n5 drain_left.t7 2.2005
R114 drain_left.n4 drain_left.t4 2.2005
R115 drain_left.n4 drain_left.t5 2.2005
R116 drain_left.n8 drain_left.n6 0.802224
R117 minus.n2 minus.t7 452.031
R118 minus.n14 minus.t3 452.031
R119 minus.n3 minus.t6 426.973
R120 minus.n4 minus.t5 426.973
R121 minus.n1 minus.t4 426.973
R122 minus.n8 minus.t1 426.973
R123 minus.n10 minus.t2 426.973
R124 minus.n15 minus.t11 426.973
R125 minus.n16 minus.t0 426.973
R126 minus.n13 minus.t8 426.973
R127 minus.n20 minus.t10 426.973
R128 minus.n22 minus.t9 426.973
R129 minus.n11 minus.n10 161.3
R130 minus.n9 minus.n0 161.3
R131 minus.n8 minus.n7 161.3
R132 minus.n23 minus.n22 161.3
R133 minus.n21 minus.n12 161.3
R134 minus.n20 minus.n19 161.3
R135 minus.n6 minus.n1 80.6037
R136 minus.n5 minus.n4 80.6037
R137 minus.n18 minus.n13 80.6037
R138 minus.n17 minus.n16 80.6037
R139 minus.n4 minus.n3 48.2005
R140 minus.n4 minus.n1 48.2005
R141 minus.n8 minus.n1 48.2005
R142 minus.n16 minus.n15 48.2005
R143 minus.n16 minus.n13 48.2005
R144 minus.n20 minus.n13 48.2005
R145 minus.n5 minus.n2 45.0744
R146 minus.n17 minus.n14 45.0744
R147 minus.n10 minus.n9 40.1672
R148 minus.n22 minus.n21 40.1672
R149 minus.n24 minus.n11 34.58
R150 minus.n3 minus.n2 16.1124
R151 minus.n15 minus.n14 16.1124
R152 minus.n9 minus.n8 8.03383
R153 minus.n21 minus.n20 8.03383
R154 minus.n24 minus.n23 6.58762
R155 minus.n6 minus.n5 0.380177
R156 minus.n18 minus.n17 0.380177
R157 minus.n7 minus.n6 0.285035
R158 minus.n19 minus.n18 0.285035
R159 minus.n11 minus.n0 0.189894
R160 minus.n7 minus.n0 0.189894
R161 minus.n19 minus.n12 0.189894
R162 minus.n23 minus.n12 0.189894
R163 minus minus.n24 0.188
R164 drain_right.n6 drain_right.n4 66.3391
R165 drain_right.n3 drain_right.n2 66.2837
R166 drain_right.n3 drain_right.n0 66.2837
R167 drain_right.n6 drain_right.n5 65.5376
R168 drain_right.n8 drain_right.n7 65.5376
R169 drain_right.n3 drain_right.n1 65.5373
R170 drain_right drain_right.n3 28.5497
R171 drain_right drain_right.n8 6.45494
R172 drain_right.n1 drain_right.t11 2.2005
R173 drain_right.n1 drain_right.t3 2.2005
R174 drain_right.n2 drain_right.t1 2.2005
R175 drain_right.n2 drain_right.t2 2.2005
R176 drain_right.n0 drain_right.t8 2.2005
R177 drain_right.n0 drain_right.t0 2.2005
R178 drain_right.n4 drain_right.t5 2.2005
R179 drain_right.n4 drain_right.t4 2.2005
R180 drain_right.n5 drain_right.t7 2.2005
R181 drain_right.n5 drain_right.t6 2.2005
R182 drain_right.n7 drain_right.t9 2.2005
R183 drain_right.n7 drain_right.t10 2.2005
R184 drain_right.n8 drain_right.n6 0.802224
C0 minus drain_right 5.53455f
C1 source drain_left 13.2047f
C2 plus drain_right 0.352374f
C3 drain_left drain_right 1.01253f
C4 source drain_right 13.2062f
C5 minus plus 5.10847f
C6 minus drain_left 0.17204f
C7 minus source 5.490799f
C8 plus drain_left 5.73172f
C9 source plus 5.50484f
C10 drain_right a_n2018_n2688# 5.54518f
C11 drain_left a_n2018_n2688# 5.84273f
C12 source a_n2018_n2688# 7.330414f
C13 minus a_n2018_n2688# 7.728847f
C14 plus a_n2018_n2688# 9.3238f
C15 drain_right.t8 a_n2018_n2688# 0.197333f
C16 drain_right.t0 a_n2018_n2688# 0.197333f
C17 drain_right.n0 a_n2018_n2688# 1.7302f
C18 drain_right.t11 a_n2018_n2688# 0.197333f
C19 drain_right.t3 a_n2018_n2688# 0.197333f
C20 drain_right.n1 a_n2018_n2688# 1.72601f
C21 drain_right.t1 a_n2018_n2688# 0.197333f
C22 drain_right.t2 a_n2018_n2688# 0.197333f
C23 drain_right.n2 a_n2018_n2688# 1.7302f
C24 drain_right.n3 a_n2018_n2688# 2.21632f
C25 drain_right.t5 a_n2018_n2688# 0.197333f
C26 drain_right.t4 a_n2018_n2688# 0.197333f
C27 drain_right.n4 a_n2018_n2688# 1.73056f
C28 drain_right.t7 a_n2018_n2688# 0.197333f
C29 drain_right.t6 a_n2018_n2688# 0.197333f
C30 drain_right.n5 a_n2018_n2688# 1.72601f
C31 drain_right.n6 a_n2018_n2688# 0.737834f
C32 drain_right.t9 a_n2018_n2688# 0.197333f
C33 drain_right.t10 a_n2018_n2688# 0.197333f
C34 drain_right.n7 a_n2018_n2688# 1.72601f
C35 drain_right.n8 a_n2018_n2688# 0.607547f
C36 minus.n0 a_n2018_n2688# 0.044096f
C37 minus.t4 a_n2018_n2688# 0.682883f
C38 minus.n1 a_n2018_n2688# 0.299048f
C39 minus.t1 a_n2018_n2688# 0.682883f
C40 minus.t7 a_n2018_n2688# 0.69888f
C41 minus.n2 a_n2018_n2688# 0.275933f
C42 minus.t6 a_n2018_n2688# 0.682883f
C43 minus.n3 a_n2018_n2688# 0.297437f
C44 minus.t5 a_n2018_n2688# 0.682883f
C45 minus.n4 a_n2018_n2688# 0.299048f
C46 minus.n5 a_n2018_n2688# 0.225996f
C47 minus.n6 a_n2018_n2688# 0.073447f
C48 minus.n7 a_n2018_n2688# 0.05884f
C49 minus.n8 a_n2018_n2688# 0.290537f
C50 minus.n9 a_n2018_n2688# 0.010006f
C51 minus.t2 a_n2018_n2688# 0.682883f
C52 minus.n10 a_n2018_n2688# 0.287546f
C53 minus.n11 a_n2018_n2688# 1.4532f
C54 minus.n12 a_n2018_n2688# 0.044096f
C55 minus.t8 a_n2018_n2688# 0.682883f
C56 minus.n13 a_n2018_n2688# 0.299048f
C57 minus.t3 a_n2018_n2688# 0.69888f
C58 minus.n14 a_n2018_n2688# 0.275933f
C59 minus.t11 a_n2018_n2688# 0.682883f
C60 minus.n15 a_n2018_n2688# 0.297437f
C61 minus.t0 a_n2018_n2688# 0.682883f
C62 minus.n16 a_n2018_n2688# 0.299048f
C63 minus.n17 a_n2018_n2688# 0.225996f
C64 minus.n18 a_n2018_n2688# 0.073447f
C65 minus.n19 a_n2018_n2688# 0.05884f
C66 minus.t10 a_n2018_n2688# 0.682883f
C67 minus.n20 a_n2018_n2688# 0.290537f
C68 minus.n21 a_n2018_n2688# 0.010006f
C69 minus.t9 a_n2018_n2688# 0.682883f
C70 minus.n22 a_n2018_n2688# 0.287546f
C71 minus.n23 a_n2018_n2688# 0.29735f
C72 minus.n24 a_n2018_n2688# 1.77004f
C73 drain_left.t0 a_n2018_n2688# 0.198293f
C74 drain_left.t1 a_n2018_n2688# 0.198293f
C75 drain_left.n0 a_n2018_n2688# 1.73862f
C76 drain_left.t2 a_n2018_n2688# 0.198293f
C77 drain_left.t8 a_n2018_n2688# 0.198293f
C78 drain_left.n1 a_n2018_n2688# 1.7344f
C79 drain_left.t10 a_n2018_n2688# 0.198293f
C80 drain_left.t3 a_n2018_n2688# 0.198293f
C81 drain_left.n2 a_n2018_n2688# 1.73862f
C82 drain_left.n3 a_n2018_n2688# 2.28433f
C83 drain_left.t4 a_n2018_n2688# 0.198293f
C84 drain_left.t5 a_n2018_n2688# 0.198293f
C85 drain_left.n4 a_n2018_n2688# 1.73898f
C86 drain_left.t6 a_n2018_n2688# 0.198293f
C87 drain_left.t7 a_n2018_n2688# 0.198293f
C88 drain_left.n5 a_n2018_n2688# 1.7344f
C89 drain_left.n6 a_n2018_n2688# 0.741415f
C90 drain_left.t9 a_n2018_n2688# 0.198293f
C91 drain_left.t11 a_n2018_n2688# 0.198293f
C92 drain_left.n7 a_n2018_n2688# 1.73439f
C93 drain_left.n8 a_n2018_n2688# 0.610509f
C94 source.t16 a_n2018_n2688# 1.75046f
C95 source.n0 a_n2018_n2688# 1.03873f
C96 source.t17 a_n2018_n2688# 0.164155f
C97 source.t15 a_n2018_n2688# 0.164155f
C98 source.n1 a_n2018_n2688# 1.37419f
C99 source.n2 a_n2018_n2688# 0.334372f
C100 source.t10 a_n2018_n2688# 0.164155f
C101 source.t18 a_n2018_n2688# 0.164155f
C102 source.n3 a_n2018_n2688# 1.37419f
C103 source.n4 a_n2018_n2688# 0.334372f
C104 source.t9 a_n2018_n2688# 1.75046f
C105 source.n5 a_n2018_n2688# 0.381117f
C106 source.t1 a_n2018_n2688# 1.75046f
C107 source.n6 a_n2018_n2688# 0.381117f
C108 source.t23 a_n2018_n2688# 0.164155f
C109 source.t2 a_n2018_n2688# 0.164155f
C110 source.n7 a_n2018_n2688# 1.37419f
C111 source.n8 a_n2018_n2688# 0.334372f
C112 source.t22 a_n2018_n2688# 0.164155f
C113 source.t0 a_n2018_n2688# 0.164155f
C114 source.n9 a_n2018_n2688# 1.37419f
C115 source.n10 a_n2018_n2688# 0.334372f
C116 source.t20 a_n2018_n2688# 1.75046f
C117 source.n11 a_n2018_n2688# 1.38039f
C118 source.t14 a_n2018_n2688# 1.75046f
C119 source.n12 a_n2018_n2688# 1.3804f
C120 source.t11 a_n2018_n2688# 0.164155f
C121 source.t13 a_n2018_n2688# 0.164155f
C122 source.n13 a_n2018_n2688# 1.37419f
C123 source.n14 a_n2018_n2688# 0.334376f
C124 source.t8 a_n2018_n2688# 0.164155f
C125 source.t12 a_n2018_n2688# 0.164155f
C126 source.n15 a_n2018_n2688# 1.37419f
C127 source.n16 a_n2018_n2688# 0.334376f
C128 source.t19 a_n2018_n2688# 1.75046f
C129 source.n17 a_n2018_n2688# 0.381121f
C130 source.t7 a_n2018_n2688# 1.75046f
C131 source.n18 a_n2018_n2688# 0.381121f
C132 source.t6 a_n2018_n2688# 0.164155f
C133 source.t3 a_n2018_n2688# 0.164155f
C134 source.n19 a_n2018_n2688# 1.37419f
C135 source.n20 a_n2018_n2688# 0.334376f
C136 source.t21 a_n2018_n2688# 0.164155f
C137 source.t5 a_n2018_n2688# 0.164155f
C138 source.n21 a_n2018_n2688# 1.37419f
C139 source.n22 a_n2018_n2688# 0.334376f
C140 source.t4 a_n2018_n2688# 1.75046f
C141 source.n23 a_n2018_n2688# 0.526656f
C142 source.n24 a_n2018_n2688# 1.21182f
C143 plus.n0 a_n2018_n2688# 0.044892f
C144 plus.t0 a_n2018_n2688# 0.695216f
C145 plus.t2 a_n2018_n2688# 0.695216f
C146 plus.n1 a_n2018_n2688# 0.059903f
C147 plus.t4 a_n2018_n2688# 0.695216f
C148 plus.n2 a_n2018_n2688# 0.074773f
C149 plus.t5 a_n2018_n2688# 0.695216f
C150 plus.n3 a_n2018_n2688# 0.230077f
C151 plus.t6 a_n2018_n2688# 0.695216f
C152 plus.t7 a_n2018_n2688# 0.711503f
C153 plus.n4 a_n2018_n2688# 0.280916f
C154 plus.n5 a_n2018_n2688# 0.30281f
C155 plus.n6 a_n2018_n2688# 0.304449f
C156 plus.n7 a_n2018_n2688# 0.304449f
C157 plus.n8 a_n2018_n2688# 0.295784f
C158 plus.n9 a_n2018_n2688# 0.010187f
C159 plus.n10 a_n2018_n2688# 0.29274f
C160 plus.n11 a_n2018_n2688# 0.450489f
C161 plus.n12 a_n2018_n2688# 0.044892f
C162 plus.t11 a_n2018_n2688# 0.695216f
C163 plus.n13 a_n2018_n2688# 0.059903f
C164 plus.t10 a_n2018_n2688# 0.695216f
C165 plus.n14 a_n2018_n2688# 0.074773f
C166 plus.t9 a_n2018_n2688# 0.695216f
C167 plus.n15 a_n2018_n2688# 0.230077f
C168 plus.t3 a_n2018_n2688# 0.695216f
C169 plus.t8 a_n2018_n2688# 0.711503f
C170 plus.n16 a_n2018_n2688# 0.280916f
C171 plus.t1 a_n2018_n2688# 0.695216f
C172 plus.n17 a_n2018_n2688# 0.30281f
C173 plus.n18 a_n2018_n2688# 0.304449f
C174 plus.n19 a_n2018_n2688# 0.304449f
C175 plus.n20 a_n2018_n2688# 0.295784f
C176 plus.n21 a_n2018_n2688# 0.010187f
C177 plus.n22 a_n2018_n2688# 0.29274f
C178 plus.n23 a_n2018_n2688# 1.29245f
.ends

