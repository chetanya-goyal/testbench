* NGSPICE file created from diffpair45.ext - technology: sky130A

.subckt diffpair45 minus drain_right drain_left source plus
X0 a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X1 drain_left.t11 plus.t0 source.t12 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X2 source.t9 minus.t0 drain_right.t11 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X3 source.t17 plus.t1 drain_left.t10 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_right.t10 minus.t1 source.t5 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X5 a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X6 a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X7 drain_right.t9 minus.t2 source.t4 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 source.t22 minus.t3 drain_right.t8 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 drain_left.t9 plus.t2 source.t20 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 drain_left.t8 plus.t3 source.t14 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 source.t23 minus.t4 drain_right.t7 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X12 source.t3 minus.t5 drain_right.t6 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X13 drain_right.t5 minus.t6 source.t0 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 drain_left.t7 plus.t4 source.t11 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X15 a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X16 drain_right.t4 minus.t7 source.t2 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X17 drain_right.t3 minus.t8 source.t7 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 drain_right.t2 minus.t9 source.t6 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X19 drain_left.t6 plus.t5 source.t13 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X20 source.t21 plus.t6 drain_left.t5 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X21 source.t10 plus.t7 drain_left.t4 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X22 source.t8 minus.t10 drain_right.t1 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 source.t18 plus.t8 drain_left.t3 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X24 source.t16 plus.t9 drain_left.t2 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 source.t19 plus.t10 drain_left.t1 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 source.t1 minus.t11 drain_right.t0 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 drain_left.t0 plus.t11 source.t15 a_n1878_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
R0 plus.n6 plus.n3 161.3
R1 plus.n8 plus.n7 161.3
R2 plus.n9 plus.n2 161.3
R3 plus.n10 plus.n1 161.3
R4 plus.n11 plus.n0 161.3
R5 plus.n13 plus.n12 161.3
R6 plus.n20 plus.n17 161.3
R7 plus.n22 plus.n21 161.3
R8 plus.n23 plus.n16 161.3
R9 plus.n24 plus.n15 161.3
R10 plus.n25 plus.n14 161.3
R11 plus.n27 plus.n26 161.3
R12 plus.n5 plus.t1 153.435
R13 plus.n19 plus.t4 153.435
R14 plus.n12 plus.t11 126.766
R15 plus.n10 plus.t9 126.766
R16 plus.n9 plus.t2 126.766
R17 plus.n3 plus.t10 126.766
R18 plus.n4 plus.t5 126.766
R19 plus.n26 plus.t7 126.766
R20 plus.n24 plus.t0 126.766
R21 plus.n23 plus.t8 126.766
R22 plus.n17 plus.t3 126.766
R23 plus.n18 plus.t6 126.766
R24 plus.n10 plus.n9 48.2005
R25 plus.n4 plus.n3 48.2005
R26 plus.n24 plus.n23 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n12 plus.n11 47.4702
R29 plus.n26 plus.n25 47.4702
R30 plus.n6 plus.n5 45.1192
R31 plus.n20 plus.n19 45.1192
R32 plus plus.n27 25.9801
R33 plus.n8 plus.n3 24.1005
R34 plus.n9 plus.n8 24.1005
R35 plus.n23 plus.n22 24.1005
R36 plus.n22 plus.n17 24.1005
R37 plus.n5 plus.n4 13.6377
R38 plus.n19 plus.n18 13.6377
R39 plus plus.n13 8.00808
R40 plus.n11 plus.n10 0.730803
R41 plus.n25 plus.n24 0.730803
R42 plus.n7 plus.n6 0.189894
R43 plus.n7 plus.n2 0.189894
R44 plus.n2 plus.n1 0.189894
R45 plus.n1 plus.n0 0.189894
R46 plus.n13 plus.n0 0.189894
R47 plus.n27 plus.n14 0.189894
R48 plus.n15 plus.n14 0.189894
R49 plus.n16 plus.n15 0.189894
R50 plus.n21 plus.n16 0.189894
R51 plus.n21 plus.n20 0.189894
R52 source.n0 source.t15 243.255
R53 source.n5 source.t17 243.255
R54 source.n6 source.t2 243.255
R55 source.n11 source.t3 243.255
R56 source.n23 source.t6 243.254
R57 source.n18 source.t23 243.254
R58 source.n17 source.t11 243.254
R59 source.n12 source.t10 243.254
R60 source.n2 source.n1 223.454
R61 source.n4 source.n3 223.454
R62 source.n8 source.n7 223.454
R63 source.n10 source.n9 223.454
R64 source.n22 source.n21 223.453
R65 source.n20 source.n19 223.453
R66 source.n16 source.n15 223.453
R67 source.n14 source.n13 223.453
R68 source.n21 source.t0 19.8005
R69 source.n21 source.t1 19.8005
R70 source.n19 source.t7 19.8005
R71 source.n19 source.t22 19.8005
R72 source.n15 source.t14 19.8005
R73 source.n15 source.t21 19.8005
R74 source.n13 source.t12 19.8005
R75 source.n13 source.t18 19.8005
R76 source.n1 source.t20 19.8005
R77 source.n1 source.t16 19.8005
R78 source.n3 source.t13 19.8005
R79 source.n3 source.t19 19.8005
R80 source.n7 source.t4 19.8005
R81 source.n7 source.t9 19.8005
R82 source.n9 source.t5 19.8005
R83 source.n9 source.t8 19.8005
R84 source.n12 source.n11 13.6699
R85 source.n24 source.n0 8.04922
R86 source.n24 source.n23 5.62119
R87 source.n11 source.n10 0.716017
R88 source.n10 source.n8 0.716017
R89 source.n8 source.n6 0.716017
R90 source.n5 source.n4 0.716017
R91 source.n4 source.n2 0.716017
R92 source.n2 source.n0 0.716017
R93 source.n14 source.n12 0.716017
R94 source.n16 source.n14 0.716017
R95 source.n17 source.n16 0.716017
R96 source.n20 source.n18 0.716017
R97 source.n22 source.n20 0.716017
R98 source.n23 source.n22 0.716017
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 240.849
R103 drain_left.n3 drain_left.n2 240.792
R104 drain_left.n3 drain_left.n0 240.792
R105 drain_left.n8 drain_left.n7 240.132
R106 drain_left.n6 drain_left.n5 240.132
R107 drain_left.n3 drain_left.n1 240.131
R108 drain_left drain_left.n3 22.6113
R109 drain_left.n1 drain_left.t3 19.8005
R110 drain_left.n1 drain_left.t8 19.8005
R111 drain_left.n2 drain_left.t5 19.8005
R112 drain_left.n2 drain_left.t7 19.8005
R113 drain_left.n0 drain_left.t4 19.8005
R114 drain_left.n0 drain_left.t11 19.8005
R115 drain_left.n7 drain_left.t2 19.8005
R116 drain_left.n7 drain_left.t0 19.8005
R117 drain_left.n5 drain_left.t1 19.8005
R118 drain_left.n5 drain_left.t9 19.8005
R119 drain_left.n4 drain_left.t10 19.8005
R120 drain_left.n4 drain_left.t6 19.8005
R121 drain_left drain_left.n8 6.36873
R122 drain_left.n8 drain_left.n6 0.716017
R123 minus.n13 minus.n12 161.3
R124 minus.n11 minus.n0 161.3
R125 minus.n10 minus.n9 161.3
R126 minus.n8 minus.n1 161.3
R127 minus.n7 minus.n6 161.3
R128 minus.n5 minus.n2 161.3
R129 minus.n27 minus.n26 161.3
R130 minus.n25 minus.n14 161.3
R131 minus.n24 minus.n23 161.3
R132 minus.n22 minus.n15 161.3
R133 minus.n21 minus.n20 161.3
R134 minus.n19 minus.n16 161.3
R135 minus.n3 minus.t7 153.435
R136 minus.n17 minus.t4 153.435
R137 minus.n4 minus.t0 126.766
R138 minus.n5 minus.t2 126.766
R139 minus.n1 minus.t10 126.766
R140 minus.n10 minus.t1 126.766
R141 minus.n12 minus.t5 126.766
R142 minus.n18 minus.t8 126.766
R143 minus.n19 minus.t3 126.766
R144 minus.n15 minus.t6 126.766
R145 minus.n24 minus.t11 126.766
R146 minus.n26 minus.t9 126.766
R147 minus.n5 minus.n4 48.2005
R148 minus.n10 minus.n1 48.2005
R149 minus.n19 minus.n18 48.2005
R150 minus.n24 minus.n15 48.2005
R151 minus.n12 minus.n11 47.4702
R152 minus.n26 minus.n25 47.4702
R153 minus.n3 minus.n2 45.1192
R154 minus.n17 minus.n16 45.1192
R155 minus.n28 minus.n13 27.9323
R156 minus.n6 minus.n1 24.1005
R157 minus.n6 minus.n5 24.1005
R158 minus.n20 minus.n19 24.1005
R159 minus.n20 minus.n15 24.1005
R160 minus.n4 minus.n3 13.6377
R161 minus.n18 minus.n17 13.6377
R162 minus.n28 minus.n27 6.5308
R163 minus.n11 minus.n10 0.730803
R164 minus.n25 minus.n24 0.730803
R165 minus.n13 minus.n0 0.189894
R166 minus.n9 minus.n0 0.189894
R167 minus.n9 minus.n8 0.189894
R168 minus.n8 minus.n7 0.189894
R169 minus.n7 minus.n2 0.189894
R170 minus.n21 minus.n16 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n14 0.189894
R174 minus.n27 minus.n14 0.189894
R175 minus minus.n28 0.188
R176 drain_right.n6 drain_right.n4 240.849
R177 drain_right.n3 drain_right.n2 240.792
R178 drain_right.n3 drain_right.n0 240.792
R179 drain_right.n6 drain_right.n5 240.132
R180 drain_right.n8 drain_right.n7 240.132
R181 drain_right.n3 drain_right.n1 240.131
R182 drain_right drain_right.n3 22.0581
R183 drain_right.n1 drain_right.t8 19.8005
R184 drain_right.n1 drain_right.t5 19.8005
R185 drain_right.n2 drain_right.t0 19.8005
R186 drain_right.n2 drain_right.t2 19.8005
R187 drain_right.n0 drain_right.t7 19.8005
R188 drain_right.n0 drain_right.t3 19.8005
R189 drain_right.n4 drain_right.t11 19.8005
R190 drain_right.n4 drain_right.t4 19.8005
R191 drain_right.n5 drain_right.t1 19.8005
R192 drain_right.n5 drain_right.t9 19.8005
R193 drain_right.n7 drain_right.t6 19.8005
R194 drain_right.n7 drain_right.t10 19.8005
R195 drain_right drain_right.n8 6.36873
R196 drain_right.n8 drain_right.n6 0.716017
C0 drain_right drain_left 0.93684f
C1 drain_right source 3.85887f
C2 minus drain_left 0.178785f
C3 minus source 1.34036f
C4 drain_right plus 0.345692f
C5 minus plus 3.46559f
C6 source drain_left 3.85792f
C7 drain_left plus 1.15156f
C8 source plus 1.35423f
C9 drain_right minus 0.969074f
C10 drain_right a_n1878_n1088# 3.46085f
C11 drain_left a_n1878_n1088# 3.69971f
C12 source a_n1878_n1088# 2.503217f
C13 minus a_n1878_n1088# 6.457456f
C14 plus a_n1878_n1088# 7.091947f
C15 drain_right.t7 a_n1878_n1088# 0.017101f
C16 drain_right.t3 a_n1878_n1088# 0.017101f
C17 drain_right.n0 a_n1878_n1088# 0.067152f
C18 drain_right.t8 a_n1878_n1088# 0.017101f
C19 drain_right.t5 a_n1878_n1088# 0.017101f
C20 drain_right.n1 a_n1878_n1088# 0.066448f
C21 drain_right.t0 a_n1878_n1088# 0.017101f
C22 drain_right.t2 a_n1878_n1088# 0.017101f
C23 drain_right.n2 a_n1878_n1088# 0.067152f
C24 drain_right.n3 a_n1878_n1088# 1.27265f
C25 drain_right.t11 a_n1878_n1088# 0.017101f
C26 drain_right.t4 a_n1878_n1088# 0.017101f
C27 drain_right.n4 a_n1878_n1088# 0.06722f
C28 drain_right.t1 a_n1878_n1088# 0.017101f
C29 drain_right.t9 a_n1878_n1088# 0.017101f
C30 drain_right.n5 a_n1878_n1088# 0.066448f
C31 drain_right.n6 a_n1878_n1088# 0.510178f
C32 drain_right.t6 a_n1878_n1088# 0.017101f
C33 drain_right.t10 a_n1878_n1088# 0.017101f
C34 drain_right.n7 a_n1878_n1088# 0.066448f
C35 drain_right.n8 a_n1878_n1088# 0.437036f
C36 minus.n0 a_n1878_n1088# 0.029627f
C37 minus.t10 a_n1878_n1088# 0.050233f
C38 minus.n1 a_n1878_n1088# 0.055265f
C39 minus.t1 a_n1878_n1088# 0.050233f
C40 minus.n2 a_n1878_n1088# 0.120662f
C41 minus.t7 a_n1878_n1088# 0.059321f
C42 minus.n3 a_n1878_n1088# 0.043889f
C43 minus.t0 a_n1878_n1088# 0.050233f
C44 minus.n4 a_n1878_n1088# 0.058836f
C45 minus.t2 a_n1878_n1088# 0.050233f
C46 minus.n5 a_n1878_n1088# 0.055265f
C47 minus.n6 a_n1878_n1088# 0.006723f
C48 minus.n7 a_n1878_n1088# 0.029627f
C49 minus.n8 a_n1878_n1088# 0.029627f
C50 minus.n9 a_n1878_n1088# 0.029627f
C51 minus.n10 a_n1878_n1088# 0.052343f
C52 minus.n11 a_n1878_n1088# 0.006723f
C53 minus.t5 a_n1878_n1088# 0.050233f
C54 minus.n12 a_n1878_n1088# 0.05216f
C55 minus.n13 a_n1878_n1088# 0.681606f
C56 minus.n14 a_n1878_n1088# 0.029627f
C57 minus.t6 a_n1878_n1088# 0.050233f
C58 minus.n15 a_n1878_n1088# 0.055265f
C59 minus.n16 a_n1878_n1088# 0.120662f
C60 minus.t4 a_n1878_n1088# 0.059321f
C61 minus.n17 a_n1878_n1088# 0.043889f
C62 minus.t8 a_n1878_n1088# 0.050233f
C63 minus.n18 a_n1878_n1088# 0.058836f
C64 minus.t3 a_n1878_n1088# 0.050233f
C65 minus.n19 a_n1878_n1088# 0.055265f
C66 minus.n20 a_n1878_n1088# 0.006723f
C67 minus.n21 a_n1878_n1088# 0.029627f
C68 minus.n22 a_n1878_n1088# 0.029627f
C69 minus.n23 a_n1878_n1088# 0.029627f
C70 minus.t11 a_n1878_n1088# 0.050233f
C71 minus.n24 a_n1878_n1088# 0.052343f
C72 minus.n25 a_n1878_n1088# 0.006723f
C73 minus.t9 a_n1878_n1088# 0.050233f
C74 minus.n26 a_n1878_n1088# 0.05216f
C75 minus.n27 a_n1878_n1088# 0.195843f
C76 minus.n28 a_n1878_n1088# 0.84137f
C77 drain_left.t4 a_n1878_n1088# 0.016737f
C78 drain_left.t11 a_n1878_n1088# 0.016737f
C79 drain_left.n0 a_n1878_n1088# 0.065726f
C80 drain_left.t3 a_n1878_n1088# 0.016737f
C81 drain_left.t8 a_n1878_n1088# 0.016737f
C82 drain_left.n1 a_n1878_n1088# 0.065037f
C83 drain_left.t5 a_n1878_n1088# 0.016737f
C84 drain_left.t7 a_n1878_n1088# 0.016737f
C85 drain_left.n2 a_n1878_n1088# 0.065726f
C86 drain_left.n3 a_n1878_n1088# 1.28654f
C87 drain_left.t10 a_n1878_n1088# 0.016737f
C88 drain_left.t6 a_n1878_n1088# 0.016737f
C89 drain_left.n4 a_n1878_n1088# 0.065792f
C90 drain_left.t1 a_n1878_n1088# 0.016737f
C91 drain_left.t9 a_n1878_n1088# 0.016737f
C92 drain_left.n5 a_n1878_n1088# 0.065037f
C93 drain_left.n6 a_n1878_n1088# 0.49934f
C94 drain_left.t2 a_n1878_n1088# 0.016737f
C95 drain_left.t0 a_n1878_n1088# 0.016737f
C96 drain_left.n7 a_n1878_n1088# 0.065037f
C97 drain_left.n8 a_n1878_n1088# 0.427752f
C98 source.t15 a_n1878_n1088# 0.110699f
C99 source.n0 a_n1878_n1088# 0.500334f
C100 source.t20 a_n1878_n1088# 0.019889f
C101 source.t16 a_n1878_n1088# 0.019889f
C102 source.n1 a_n1878_n1088# 0.064503f
C103 source.n2 a_n1878_n1088# 0.270631f
C104 source.t13 a_n1878_n1088# 0.019889f
C105 source.t19 a_n1878_n1088# 0.019889f
C106 source.n3 a_n1878_n1088# 0.064503f
C107 source.n4 a_n1878_n1088# 0.270631f
C108 source.t17 a_n1878_n1088# 0.110699f
C109 source.n5 a_n1878_n1088# 0.258752f
C110 source.t2 a_n1878_n1088# 0.110699f
C111 source.n6 a_n1878_n1088# 0.258752f
C112 source.t4 a_n1878_n1088# 0.019889f
C113 source.t9 a_n1878_n1088# 0.019889f
C114 source.n7 a_n1878_n1088# 0.064503f
C115 source.n8 a_n1878_n1088# 0.270631f
C116 source.t5 a_n1878_n1088# 0.019889f
C117 source.t8 a_n1878_n1088# 0.019889f
C118 source.n9 a_n1878_n1088# 0.064503f
C119 source.n10 a_n1878_n1088# 0.270631f
C120 source.t3 a_n1878_n1088# 0.110699f
C121 source.n11 a_n1878_n1088# 0.704962f
C122 source.t10 a_n1878_n1088# 0.110698f
C123 source.n12 a_n1878_n1088# 0.704962f
C124 source.t12 a_n1878_n1088# 0.019889f
C125 source.t18 a_n1878_n1088# 0.019889f
C126 source.n13 a_n1878_n1088# 0.064503f
C127 source.n14 a_n1878_n1088# 0.270631f
C128 source.t14 a_n1878_n1088# 0.019889f
C129 source.t21 a_n1878_n1088# 0.019889f
C130 source.n15 a_n1878_n1088# 0.064503f
C131 source.n16 a_n1878_n1088# 0.270631f
C132 source.t11 a_n1878_n1088# 0.110698f
C133 source.n17 a_n1878_n1088# 0.258752f
C134 source.t23 a_n1878_n1088# 0.110698f
C135 source.n18 a_n1878_n1088# 0.258752f
C136 source.t7 a_n1878_n1088# 0.019889f
C137 source.t22 a_n1878_n1088# 0.019889f
C138 source.n19 a_n1878_n1088# 0.064503f
C139 source.n20 a_n1878_n1088# 0.270631f
C140 source.t0 a_n1878_n1088# 0.019889f
C141 source.t1 a_n1878_n1088# 0.019889f
C142 source.n21 a_n1878_n1088# 0.064503f
C143 source.n22 a_n1878_n1088# 0.270631f
C144 source.t6 a_n1878_n1088# 0.110698f
C145 source.n23 a_n1878_n1088# 0.41194f
C146 source.n24 a_n1878_n1088# 0.515551f
C147 plus.n0 a_n1878_n1088# 0.030143f
C148 plus.t11 a_n1878_n1088# 0.051108f
C149 plus.t9 a_n1878_n1088# 0.051108f
C150 plus.n1 a_n1878_n1088# 0.030143f
C151 plus.t2 a_n1878_n1088# 0.051108f
C152 plus.n2 a_n1878_n1088# 0.030143f
C153 plus.t10 a_n1878_n1088# 0.051108f
C154 plus.n3 a_n1878_n1088# 0.056228f
C155 plus.t5 a_n1878_n1088# 0.051108f
C156 plus.n4 a_n1878_n1088# 0.059861f
C157 plus.t1 a_n1878_n1088# 0.060354f
C158 plus.n5 a_n1878_n1088# 0.044654f
C159 plus.n6 a_n1878_n1088# 0.122763f
C160 plus.n7 a_n1878_n1088# 0.030143f
C161 plus.n8 a_n1878_n1088# 0.00684f
C162 plus.n9 a_n1878_n1088# 0.056228f
C163 plus.n10 a_n1878_n1088# 0.053254f
C164 plus.n11 a_n1878_n1088# 0.00684f
C165 plus.n12 a_n1878_n1088# 0.053068f
C166 plus.n13 a_n1878_n1088# 0.208965f
C167 plus.n14 a_n1878_n1088# 0.030143f
C168 plus.t7 a_n1878_n1088# 0.051108f
C169 plus.n15 a_n1878_n1088# 0.030143f
C170 plus.t0 a_n1878_n1088# 0.051108f
C171 plus.n16 a_n1878_n1088# 0.030143f
C172 plus.t8 a_n1878_n1088# 0.051108f
C173 plus.t3 a_n1878_n1088# 0.051108f
C174 plus.n17 a_n1878_n1088# 0.056228f
C175 plus.t4 a_n1878_n1088# 0.060354f
C176 plus.t6 a_n1878_n1088# 0.051108f
C177 plus.n18 a_n1878_n1088# 0.059861f
C178 plus.n19 a_n1878_n1088# 0.044654f
C179 plus.n20 a_n1878_n1088# 0.122763f
C180 plus.n21 a_n1878_n1088# 0.030143f
C181 plus.n22 a_n1878_n1088# 0.00684f
C182 plus.n23 a_n1878_n1088# 0.056228f
C183 plus.n24 a_n1878_n1088# 0.053254f
C184 plus.n25 a_n1878_n1088# 0.00684f
C185 plus.n26 a_n1878_n1088# 0.053068f
C186 plus.n27 a_n1878_n1088# 0.672341f
.ends

