* NGSPICE file created from diffpair230.ext - technology: sky130A

.subckt diffpair230 minus drain_right drain_left source plus
X0 drain_right minus source a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.8
X1 a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X2 a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X3 drain_left plus source a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.8
X4 a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X5 drain_left plus source a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.8
X6 a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X7 drain_right minus source a_n1168_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.8
.ends

