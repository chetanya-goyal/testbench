* NGSPICE file created from diffpair397.ext - technology: sky130A

.subckt diffpair397 minus drain_right drain_left source plus
X0 a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X1 drain_right.t15 minus.t0 source.t31 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X2 drain_right.t14 minus.t1 source.t30 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X3 source.t1 plus.t0 drain_left.t15 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X5 source.t6 plus.t1 drain_left.t14 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 drain_right.t13 minus.t2 source.t16 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X7 drain_left.t13 plus.t2 source.t8 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X9 drain_right.t12 minus.t3 source.t17 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 drain_left.t12 plus.t3 source.t10 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X12 drain_left.t11 plus.t4 source.t0 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X13 source.t25 minus.t4 drain_right.t11 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X14 source.t22 minus.t5 drain_right.t10 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X15 drain_right.t9 minus.t6 source.t29 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X16 source.t24 minus.t7 drain_right.t8 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X17 drain_right.t7 minus.t8 source.t18 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X18 source.t26 minus.t9 drain_right.t6 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 drain_left.t10 plus.t5 source.t9 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X20 source.t19 minus.t10 drain_right.t5 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X21 drain_left.t9 plus.t6 source.t11 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X22 drain_right.t4 minus.t11 source.t23 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X23 source.t14 plus.t7 drain_left.t8 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X24 source.t20 minus.t12 drain_right.t3 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X25 drain_left.t7 plus.t8 source.t7 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X26 drain_left.t6 plus.t9 source.t12 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X27 source.t27 minus.t13 drain_right.t2 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X28 source.t28 minus.t14 drain_right.t1 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X29 source.t5 plus.t10 drain_left.t5 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X30 source.t13 plus.t11 drain_left.t4 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X31 drain_right.t0 minus.t15 source.t21 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X32 source.t15 plus.t12 drain_left.t3 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X33 drain_left.t2 plus.t13 source.t4 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X34 source.t2 plus.t14 drain_left.t1 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X35 source.t3 plus.t15 drain_left.t0 a_n2750_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n5 minus.t8 341.252
R1 minus.n27 minus.t14 341.252
R2 minus.n6 minus.t4 320.229
R3 minus.n7 minus.t3 320.229
R4 minus.n3 minus.t10 320.229
R5 minus.n13 minus.t11 320.229
R6 minus.n1 minus.t9 320.229
R7 minus.n18 minus.t6 320.229
R8 minus.n20 minus.t13 320.229
R9 minus.n28 minus.t2 320.229
R10 minus.n29 minus.t7 320.229
R11 minus.n25 minus.t1 320.229
R12 minus.n35 minus.t12 320.229
R13 minus.n23 minus.t0 320.229
R14 minus.n40 minus.t5 320.229
R15 minus.n42 minus.t15 320.229
R16 minus.n21 minus.n20 161.3
R17 minus.n19 minus.n0 161.3
R18 minus.n15 minus.n14 161.3
R19 minus.n13 minus.n2 161.3
R20 minus.n12 minus.n11 161.3
R21 minus.n10 minus.n3 161.3
R22 minus.n9 minus.n8 161.3
R23 minus.n43 minus.n42 161.3
R24 minus.n41 minus.n22 161.3
R25 minus.n37 minus.n36 161.3
R26 minus.n35 minus.n24 161.3
R27 minus.n34 minus.n33 161.3
R28 minus.n32 minus.n25 161.3
R29 minus.n31 minus.n30 161.3
R30 minus.n18 minus.n17 80.6037
R31 minus.n16 minus.n1 80.6037
R32 minus.n7 minus.n4 80.6037
R33 minus.n40 minus.n39 80.6037
R34 minus.n38 minus.n23 80.6037
R35 minus.n29 minus.n26 80.6037
R36 minus.n7 minus.n6 48.2005
R37 minus.n18 minus.n1 48.2005
R38 minus.n29 minus.n28 48.2005
R39 minus.n40 minus.n23 48.2005
R40 minus.n8 minus.n7 43.0884
R41 minus.n14 minus.n1 43.0884
R42 minus.n30 minus.n29 43.0884
R43 minus.n36 minus.n23 43.0884
R44 minus.n19 minus.n18 40.1672
R45 minus.n41 minus.n40 40.1672
R46 minus.n44 minus.n21 37.421
R47 minus.n5 minus.n4 31.6481
R48 minus.n27 minus.n26 31.6481
R49 minus.n13 minus.n12 24.1005
R50 minus.n12 minus.n3 24.1005
R51 minus.n34 minus.n25 24.1005
R52 minus.n35 minus.n34 24.1005
R53 minus.n6 minus.n5 17.444
R54 minus.n28 minus.n27 17.444
R55 minus.n20 minus.n19 8.03383
R56 minus.n42 minus.n41 8.03383
R57 minus.n44 minus.n43 6.6558
R58 minus.n8 minus.n3 5.11262
R59 minus.n14 minus.n13 5.11262
R60 minus.n30 minus.n25 5.11262
R61 minus.n36 minus.n35 5.11262
R62 minus.n17 minus.n16 0.380177
R63 minus.n39 minus.n38 0.380177
R64 minus.n17 minus.n0 0.285035
R65 minus.n16 minus.n15 0.285035
R66 minus.n9 minus.n4 0.285035
R67 minus.n31 minus.n26 0.285035
R68 minus.n38 minus.n37 0.285035
R69 minus.n39 minus.n22 0.285035
R70 minus.n21 minus.n0 0.189894
R71 minus.n15 minus.n2 0.189894
R72 minus.n11 minus.n2 0.189894
R73 minus.n11 minus.n10 0.189894
R74 minus.n10 minus.n9 0.189894
R75 minus.n32 minus.n31 0.189894
R76 minus.n33 minus.n32 0.189894
R77 minus.n33 minus.n24 0.189894
R78 minus.n37 minus.n24 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 source.n7 source.t2 51.0588
R82 source.n8 source.t18 51.0588
R83 source.n15 source.t27 51.0588
R84 source.n31 source.t21 51.0586
R85 source.n24 source.t28 51.0586
R86 source.n23 source.t11 51.0586
R87 source.n16 source.t3 51.0586
R88 source.n0 source.t9 51.0586
R89 source.n2 source.n1 48.8588
R90 source.n4 source.n3 48.8588
R91 source.n6 source.n5 48.8588
R92 source.n10 source.n9 48.8588
R93 source.n12 source.n11 48.8588
R94 source.n14 source.n13 48.8588
R95 source.n30 source.n29 48.8586
R96 source.n28 source.n27 48.8586
R97 source.n26 source.n25 48.8586
R98 source.n22 source.n21 48.8586
R99 source.n20 source.n19 48.8586
R100 source.n18 source.n17 48.8586
R101 source.n16 source.n15 19.9891
R102 source.n32 source.n0 14.2391
R103 source.n32 source.n31 5.7505
R104 source.n29 source.t31 2.2005
R105 source.n29 source.t22 2.2005
R106 source.n27 source.t30 2.2005
R107 source.n27 source.t20 2.2005
R108 source.n25 source.t16 2.2005
R109 source.n25 source.t24 2.2005
R110 source.n21 source.t0 2.2005
R111 source.n21 source.t6 2.2005
R112 source.n19 source.t10 2.2005
R113 source.n19 source.t1 2.2005
R114 source.n17 source.t8 2.2005
R115 source.n17 source.t5 2.2005
R116 source.n1 source.t7 2.2005
R117 source.n1 source.t14 2.2005
R118 source.n3 source.t12 2.2005
R119 source.n3 source.t15 2.2005
R120 source.n5 source.t4 2.2005
R121 source.n5 source.t13 2.2005
R122 source.n9 source.t17 2.2005
R123 source.n9 source.t25 2.2005
R124 source.n11 source.t23 2.2005
R125 source.n11 source.t19 2.2005
R126 source.n13 source.t29 2.2005
R127 source.n13 source.t26 2.2005
R128 source.n15 source.n14 0.974638
R129 source.n14 source.n12 0.974638
R130 source.n12 source.n10 0.974638
R131 source.n10 source.n8 0.974638
R132 source.n7 source.n6 0.974638
R133 source.n6 source.n4 0.974638
R134 source.n4 source.n2 0.974638
R135 source.n2 source.n0 0.974638
R136 source.n18 source.n16 0.974638
R137 source.n20 source.n18 0.974638
R138 source.n22 source.n20 0.974638
R139 source.n23 source.n22 0.974638
R140 source.n26 source.n24 0.974638
R141 source.n28 source.n26 0.974638
R142 source.n30 source.n28 0.974638
R143 source.n31 source.n30 0.974638
R144 source.n8 source.n7 0.470328
R145 source.n24 source.n23 0.470328
R146 source source.n32 0.188
R147 drain_right.n9 drain_right.n7 66.5116
R148 drain_right.n5 drain_right.n3 66.5115
R149 drain_right.n2 drain_right.n0 66.5115
R150 drain_right.n9 drain_right.n8 65.5376
R151 drain_right.n11 drain_right.n10 65.5376
R152 drain_right.n13 drain_right.n12 65.5376
R153 drain_right.n5 drain_right.n4 65.5373
R154 drain_right.n2 drain_right.n1 65.5373
R155 drain_right drain_right.n6 30.873
R156 drain_right drain_right.n13 6.62735
R157 drain_right.n3 drain_right.t10 2.2005
R158 drain_right.n3 drain_right.t0 2.2005
R159 drain_right.n4 drain_right.t3 2.2005
R160 drain_right.n4 drain_right.t15 2.2005
R161 drain_right.n1 drain_right.t8 2.2005
R162 drain_right.n1 drain_right.t14 2.2005
R163 drain_right.n0 drain_right.t1 2.2005
R164 drain_right.n0 drain_right.t13 2.2005
R165 drain_right.n7 drain_right.t11 2.2005
R166 drain_right.n7 drain_right.t7 2.2005
R167 drain_right.n8 drain_right.t5 2.2005
R168 drain_right.n8 drain_right.t12 2.2005
R169 drain_right.n10 drain_right.t6 2.2005
R170 drain_right.n10 drain_right.t4 2.2005
R171 drain_right.n12 drain_right.t2 2.2005
R172 drain_right.n12 drain_right.t9 2.2005
R173 drain_right.n13 drain_right.n11 0.974638
R174 drain_right.n11 drain_right.n9 0.974638
R175 drain_right.n6 drain_right.n5 0.432223
R176 drain_right.n6 drain_right.n2 0.432223
R177 plus.n7 plus.t14 341.252
R178 plus.n29 plus.t6 341.252
R179 plus.n20 plus.t5 320.229
R180 plus.n18 plus.t7 320.229
R181 plus.n17 plus.t8 320.229
R182 plus.n3 plus.t12 320.229
R183 plus.n11 plus.t9 320.229
R184 plus.n5 plus.t11 320.229
R185 plus.n6 plus.t13 320.229
R186 plus.n42 plus.t15 320.229
R187 plus.n40 plus.t2 320.229
R188 plus.n39 plus.t10 320.229
R189 plus.n25 plus.t3 320.229
R190 plus.n33 plus.t0 320.229
R191 plus.n27 plus.t4 320.229
R192 plus.n28 plus.t1 320.229
R193 plus.n10 plus.n9 161.3
R194 plus.n11 plus.n4 161.3
R195 plus.n13 plus.n12 161.3
R196 plus.n14 plus.n3 161.3
R197 plus.n16 plus.n15 161.3
R198 plus.n19 plus.n0 161.3
R199 plus.n21 plus.n20 161.3
R200 plus.n32 plus.n31 161.3
R201 plus.n33 plus.n26 161.3
R202 plus.n35 plus.n34 161.3
R203 plus.n36 plus.n25 161.3
R204 plus.n38 plus.n37 161.3
R205 plus.n41 plus.n22 161.3
R206 plus.n43 plus.n42 161.3
R207 plus.n8 plus.n5 80.6037
R208 plus.n17 plus.n2 80.6037
R209 plus.n18 plus.n1 80.6037
R210 plus.n30 plus.n27 80.6037
R211 plus.n39 plus.n24 80.6037
R212 plus.n40 plus.n23 80.6037
R213 plus.n18 plus.n17 48.2005
R214 plus.n6 plus.n5 48.2005
R215 plus.n40 plus.n39 48.2005
R216 plus.n28 plus.n27 48.2005
R217 plus.n17 plus.n16 43.0884
R218 plus.n10 plus.n5 43.0884
R219 plus.n39 plus.n38 43.0884
R220 plus.n32 plus.n27 43.0884
R221 plus.n19 plus.n18 40.1672
R222 plus.n41 plus.n40 40.1672
R223 plus plus.n43 32.4384
R224 plus.n8 plus.n7 31.6481
R225 plus.n30 plus.n29 31.6481
R226 plus.n12 plus.n11 24.1005
R227 plus.n12 plus.n3 24.1005
R228 plus.n34 plus.n25 24.1005
R229 plus.n34 plus.n33 24.1005
R230 plus.n7 plus.n6 17.444
R231 plus.n29 plus.n28 17.444
R232 plus plus.n21 11.1634
R233 plus.n20 plus.n19 8.03383
R234 plus.n42 plus.n41 8.03383
R235 plus.n16 plus.n3 5.11262
R236 plus.n11 plus.n10 5.11262
R237 plus.n38 plus.n25 5.11262
R238 plus.n33 plus.n32 5.11262
R239 plus.n2 plus.n1 0.380177
R240 plus.n24 plus.n23 0.380177
R241 plus.n9 plus.n8 0.285035
R242 plus.n15 plus.n2 0.285035
R243 plus.n1 plus.n0 0.285035
R244 plus.n23 plus.n22 0.285035
R245 plus.n37 plus.n24 0.285035
R246 plus.n31 plus.n30 0.285035
R247 plus.n9 plus.n4 0.189894
R248 plus.n13 plus.n4 0.189894
R249 plus.n14 plus.n13 0.189894
R250 plus.n15 plus.n14 0.189894
R251 plus.n21 plus.n0 0.189894
R252 plus.n43 plus.n22 0.189894
R253 plus.n37 plus.n36 0.189894
R254 plus.n36 plus.n35 0.189894
R255 plus.n35 plus.n26 0.189894
R256 plus.n31 plus.n26 0.189894
R257 drain_left.n9 drain_left.n7 66.5117
R258 drain_left.n5 drain_left.n3 66.5115
R259 drain_left.n2 drain_left.n0 66.5115
R260 drain_left.n11 drain_left.n10 65.5376
R261 drain_left.n9 drain_left.n8 65.5376
R262 drain_left.n13 drain_left.n12 65.5374
R263 drain_left.n5 drain_left.n4 65.5373
R264 drain_left.n2 drain_left.n1 65.5373
R265 drain_left drain_left.n6 31.4262
R266 drain_left drain_left.n13 6.62735
R267 drain_left.n3 drain_left.t14 2.2005
R268 drain_left.n3 drain_left.t9 2.2005
R269 drain_left.n4 drain_left.t15 2.2005
R270 drain_left.n4 drain_left.t11 2.2005
R271 drain_left.n1 drain_left.t5 2.2005
R272 drain_left.n1 drain_left.t12 2.2005
R273 drain_left.n0 drain_left.t0 2.2005
R274 drain_left.n0 drain_left.t13 2.2005
R275 drain_left.n12 drain_left.t8 2.2005
R276 drain_left.n12 drain_left.t10 2.2005
R277 drain_left.n10 drain_left.t3 2.2005
R278 drain_left.n10 drain_left.t7 2.2005
R279 drain_left.n8 drain_left.t4 2.2005
R280 drain_left.n8 drain_left.t6 2.2005
R281 drain_left.n7 drain_left.t1 2.2005
R282 drain_left.n7 drain_left.t2 2.2005
R283 drain_left.n11 drain_left.n9 0.974638
R284 drain_left.n13 drain_left.n11 0.974638
R285 drain_left.n6 drain_left.n5 0.432223
R286 drain_left.n6 drain_left.n2 0.432223
C0 drain_right source 14.8155f
C1 minus drain_left 0.173489f
C2 minus source 8.607241f
C3 source drain_left 14.8128f
C4 drain_right plus 0.430381f
C5 minus plus 6.02047f
C6 drain_right minus 8.38726f
C7 plus drain_left 8.66064f
C8 plus source 8.62128f
C9 drain_right drain_left 1.44945f
C10 drain_right a_n2750_n2688# 6.37444f
C11 drain_left a_n2750_n2688# 6.76622f
C12 source a_n2750_n2688# 7.698781f
C13 minus a_n2750_n2688# 10.813323f
C14 plus a_n2750_n2688# 12.377789f
C15 drain_left.t0 a_n2750_n2688# 0.189599f
C16 drain_left.t13 a_n2750_n2688# 0.189599f
C17 drain_left.n0 a_n2750_n2688# 1.6641f
C18 drain_left.t5 a_n2750_n2688# 0.189599f
C19 drain_left.t12 a_n2750_n2688# 0.189599f
C20 drain_left.n1 a_n2750_n2688# 1.65836f
C21 drain_left.n2 a_n2750_n2688# 0.721635f
C22 drain_left.t14 a_n2750_n2688# 0.189599f
C23 drain_left.t9 a_n2750_n2688# 0.189599f
C24 drain_left.n3 a_n2750_n2688# 1.6641f
C25 drain_left.t15 a_n2750_n2688# 0.189599f
C26 drain_left.t11 a_n2750_n2688# 0.189599f
C27 drain_left.n4 a_n2750_n2688# 1.65836f
C28 drain_left.n5 a_n2750_n2688# 0.721635f
C29 drain_left.n6 a_n2750_n2688# 1.40522f
C30 drain_left.t1 a_n2750_n2688# 0.189599f
C31 drain_left.t2 a_n2750_n2688# 0.189599f
C32 drain_left.n7 a_n2750_n2688# 1.6641f
C33 drain_left.t4 a_n2750_n2688# 0.189599f
C34 drain_left.t6 a_n2750_n2688# 0.189599f
C35 drain_left.n8 a_n2750_n2688# 1.65836f
C36 drain_left.n9 a_n2750_n2688# 0.766791f
C37 drain_left.t3 a_n2750_n2688# 0.189599f
C38 drain_left.t7 a_n2750_n2688# 0.189599f
C39 drain_left.n10 a_n2750_n2688# 1.65836f
C40 drain_left.n11 a_n2750_n2688# 0.380895f
C41 drain_left.t8 a_n2750_n2688# 0.189599f
C42 drain_left.t10 a_n2750_n2688# 0.189599f
C43 drain_left.n12 a_n2750_n2688# 1.65836f
C44 drain_left.n13 a_n2750_n2688# 0.61995f
C45 plus.n0 a_n2750_n2688# 0.052512f
C46 plus.t5 a_n2750_n2688# 0.81259f
C47 plus.t7 a_n2750_n2688# 0.81259f
C48 plus.n1 a_n2750_n2688# 0.065548f
C49 plus.t8 a_n2750_n2688# 0.81259f
C50 plus.n2 a_n2750_n2688# 0.065548f
C51 plus.t12 a_n2750_n2688# 0.81259f
C52 plus.n3 a_n2750_n2688# 0.337811f
C53 plus.n4 a_n2750_n2688# 0.039353f
C54 plus.t9 a_n2750_n2688# 0.81259f
C55 plus.t11 a_n2750_n2688# 0.81259f
C56 plus.n5 a_n2750_n2688# 0.349047f
C57 plus.t13 a_n2750_n2688# 0.81259f
C58 plus.n6 a_n2750_n2688# 0.349355f
C59 plus.t14 a_n2750_n2688# 0.833613f
C60 plus.n7 a_n2750_n2688# 0.323753f
C61 plus.n8 a_n2750_n2688# 0.22571f
C62 plus.n9 a_n2750_n2688# 0.052512f
C63 plus.n10 a_n2750_n2688# 0.00893f
C64 plus.n11 a_n2750_n2688# 0.337811f
C65 plus.n12 a_n2750_n2688# 0.00893f
C66 plus.n13 a_n2750_n2688# 0.039353f
C67 plus.n14 a_n2750_n2688# 0.039353f
C68 plus.n15 a_n2750_n2688# 0.052512f
C69 plus.n16 a_n2750_n2688# 0.00893f
C70 plus.n17 a_n2750_n2688# 0.349047f
C71 plus.n18 a_n2750_n2688# 0.348561f
C72 plus.n19 a_n2750_n2688# 0.00893f
C73 plus.n20 a_n2750_n2688# 0.334293f
C74 plus.n21 a_n2750_n2688# 0.401372f
C75 plus.n22 a_n2750_n2688# 0.052512f
C76 plus.t15 a_n2750_n2688# 0.81259f
C77 plus.n23 a_n2750_n2688# 0.065548f
C78 plus.t2 a_n2750_n2688# 0.81259f
C79 plus.n24 a_n2750_n2688# 0.065548f
C80 plus.t10 a_n2750_n2688# 0.81259f
C81 plus.t3 a_n2750_n2688# 0.81259f
C82 plus.n25 a_n2750_n2688# 0.337811f
C83 plus.n26 a_n2750_n2688# 0.039353f
C84 plus.t0 a_n2750_n2688# 0.81259f
C85 plus.t4 a_n2750_n2688# 0.81259f
C86 plus.n27 a_n2750_n2688# 0.349047f
C87 plus.t1 a_n2750_n2688# 0.81259f
C88 plus.n28 a_n2750_n2688# 0.349355f
C89 plus.t6 a_n2750_n2688# 0.833613f
C90 plus.n29 a_n2750_n2688# 0.323753f
C91 plus.n30 a_n2750_n2688# 0.22571f
C92 plus.n31 a_n2750_n2688# 0.052512f
C93 plus.n32 a_n2750_n2688# 0.00893f
C94 plus.n33 a_n2750_n2688# 0.337811f
C95 plus.n34 a_n2750_n2688# 0.00893f
C96 plus.n35 a_n2750_n2688# 0.039353f
C97 plus.n36 a_n2750_n2688# 0.039353f
C98 plus.n37 a_n2750_n2688# 0.052512f
C99 plus.n38 a_n2750_n2688# 0.00893f
C100 plus.n39 a_n2750_n2688# 0.349047f
C101 plus.n40 a_n2750_n2688# 0.348561f
C102 plus.n41 a_n2750_n2688# 0.00893f
C103 plus.n42 a_n2750_n2688# 0.334293f
C104 plus.n43 a_n2750_n2688# 1.29025f
C105 drain_right.t1 a_n2750_n2688# 0.188013f
C106 drain_right.t13 a_n2750_n2688# 0.188013f
C107 drain_right.n0 a_n2750_n2688# 1.65018f
C108 drain_right.t8 a_n2750_n2688# 0.188013f
C109 drain_right.t14 a_n2750_n2688# 0.188013f
C110 drain_right.n1 a_n2750_n2688# 1.64449f
C111 drain_right.n2 a_n2750_n2688# 0.715599f
C112 drain_right.t10 a_n2750_n2688# 0.188013f
C113 drain_right.t0 a_n2750_n2688# 0.188013f
C114 drain_right.n3 a_n2750_n2688# 1.65018f
C115 drain_right.t3 a_n2750_n2688# 0.188013f
C116 drain_right.t15 a_n2750_n2688# 0.188013f
C117 drain_right.n4 a_n2750_n2688# 1.64449f
C118 drain_right.n5 a_n2750_n2688# 0.715599f
C119 drain_right.n6 a_n2750_n2688# 1.33984f
C120 drain_right.t11 a_n2750_n2688# 0.188013f
C121 drain_right.t7 a_n2750_n2688# 0.188013f
C122 drain_right.n7 a_n2750_n2688# 1.65017f
C123 drain_right.t5 a_n2750_n2688# 0.188013f
C124 drain_right.t12 a_n2750_n2688# 0.188013f
C125 drain_right.n8 a_n2750_n2688# 1.64449f
C126 drain_right.n9 a_n2750_n2688# 0.760384f
C127 drain_right.t6 a_n2750_n2688# 0.188013f
C128 drain_right.t4 a_n2750_n2688# 0.188013f
C129 drain_right.n10 a_n2750_n2688# 1.64449f
C130 drain_right.n11 a_n2750_n2688# 0.377708f
C131 drain_right.t2 a_n2750_n2688# 0.188013f
C132 drain_right.t9 a_n2750_n2688# 0.188013f
C133 drain_right.n12 a_n2750_n2688# 1.64449f
C134 drain_right.n13 a_n2750_n2688# 0.614757f
C135 source.t9 a_n2750_n2688# 1.78055f
C136 source.n0 a_n2750_n2688# 1.07837f
C137 source.t7 a_n2750_n2688# 0.166976f
C138 source.t14 a_n2750_n2688# 0.166976f
C139 source.n1 a_n2750_n2688# 1.39782f
C140 source.n2 a_n2750_n2688# 0.366207f
C141 source.t12 a_n2750_n2688# 0.166976f
C142 source.t15 a_n2750_n2688# 0.166976f
C143 source.n3 a_n2750_n2688# 1.39782f
C144 source.n4 a_n2750_n2688# 0.366207f
C145 source.t4 a_n2750_n2688# 0.166976f
C146 source.t13 a_n2750_n2688# 0.166976f
C147 source.n5 a_n2750_n2688# 1.39782f
C148 source.n6 a_n2750_n2688# 0.366207f
C149 source.t2 a_n2750_n2688# 1.78055f
C150 source.n7 a_n2750_n2688# 0.400711f
C151 source.t18 a_n2750_n2688# 1.78055f
C152 source.n8 a_n2750_n2688# 0.400711f
C153 source.t17 a_n2750_n2688# 0.166976f
C154 source.t25 a_n2750_n2688# 0.166976f
C155 source.n9 a_n2750_n2688# 1.39782f
C156 source.n10 a_n2750_n2688# 0.366207f
C157 source.t23 a_n2750_n2688# 0.166976f
C158 source.t19 a_n2750_n2688# 0.166976f
C159 source.n11 a_n2750_n2688# 1.39782f
C160 source.n12 a_n2750_n2688# 0.366207f
C161 source.t29 a_n2750_n2688# 0.166976f
C162 source.t26 a_n2750_n2688# 0.166976f
C163 source.n13 a_n2750_n2688# 1.39782f
C164 source.n14 a_n2750_n2688# 0.366207f
C165 source.t27 a_n2750_n2688# 1.78055f
C166 source.n15 a_n2750_n2688# 1.43021f
C167 source.t3 a_n2750_n2688# 1.78055f
C168 source.n16 a_n2750_n2688# 1.43021f
C169 source.t8 a_n2750_n2688# 0.166976f
C170 source.t5 a_n2750_n2688# 0.166976f
C171 source.n17 a_n2750_n2688# 1.39781f
C172 source.n18 a_n2750_n2688# 0.366211f
C173 source.t10 a_n2750_n2688# 0.166976f
C174 source.t1 a_n2750_n2688# 0.166976f
C175 source.n19 a_n2750_n2688# 1.39781f
C176 source.n20 a_n2750_n2688# 0.366211f
C177 source.t0 a_n2750_n2688# 0.166976f
C178 source.t6 a_n2750_n2688# 0.166976f
C179 source.n21 a_n2750_n2688# 1.39781f
C180 source.n22 a_n2750_n2688# 0.366211f
C181 source.t11 a_n2750_n2688# 1.78055f
C182 source.n23 a_n2750_n2688# 0.400716f
C183 source.t28 a_n2750_n2688# 1.78055f
C184 source.n24 a_n2750_n2688# 0.400716f
C185 source.t16 a_n2750_n2688# 0.166976f
C186 source.t24 a_n2750_n2688# 0.166976f
C187 source.n25 a_n2750_n2688# 1.39781f
C188 source.n26 a_n2750_n2688# 0.366211f
C189 source.t30 a_n2750_n2688# 0.166976f
C190 source.t20 a_n2750_n2688# 0.166976f
C191 source.n27 a_n2750_n2688# 1.39781f
C192 source.n28 a_n2750_n2688# 0.366211f
C193 source.t31 a_n2750_n2688# 0.166976f
C194 source.t22 a_n2750_n2688# 0.166976f
C195 source.n29 a_n2750_n2688# 1.39781f
C196 source.n30 a_n2750_n2688# 0.366211f
C197 source.t21 a_n2750_n2688# 1.78055f
C198 source.n31 a_n2750_n2688# 0.558945f
C199 source.n32 a_n2750_n2688# 1.23981f
C200 minus.n0 a_n2750_n2688# 0.05166f
C201 minus.t9 a_n2750_n2688# 0.799397f
C202 minus.n1 a_n2750_n2688# 0.343379f
C203 minus.t6 a_n2750_n2688# 0.799397f
C204 minus.n2 a_n2750_n2688# 0.038714f
C205 minus.t10 a_n2750_n2688# 0.799397f
C206 minus.n3 a_n2750_n2688# 0.332327f
C207 minus.n4 a_n2750_n2688# 0.222046f
C208 minus.t8 a_n2750_n2688# 0.820079f
C209 minus.n5 a_n2750_n2688# 0.318496f
C210 minus.t4 a_n2750_n2688# 0.799397f
C211 minus.n6 a_n2750_n2688# 0.343683f
C212 minus.t3 a_n2750_n2688# 0.799397f
C213 minus.n7 a_n2750_n2688# 0.343379f
C214 minus.n8 a_n2750_n2688# 0.008785f
C215 minus.n9 a_n2750_n2688# 0.05166f
C216 minus.n10 a_n2750_n2688# 0.038714f
C217 minus.n11 a_n2750_n2688# 0.038714f
C218 minus.n12 a_n2750_n2688# 0.008785f
C219 minus.t11 a_n2750_n2688# 0.799397f
C220 minus.n13 a_n2750_n2688# 0.332327f
C221 minus.n14 a_n2750_n2688# 0.008785f
C222 minus.n15 a_n2750_n2688# 0.05166f
C223 minus.n16 a_n2750_n2688# 0.064484f
C224 minus.n17 a_n2750_n2688# 0.064484f
C225 minus.n18 a_n2750_n2688# 0.342902f
C226 minus.n19 a_n2750_n2688# 0.008785f
C227 minus.t13 a_n2750_n2688# 0.799397f
C228 minus.n20 a_n2750_n2688# 0.328866f
C229 minus.n21 a_n2750_n2688# 1.4454f
C230 minus.n22 a_n2750_n2688# 0.05166f
C231 minus.t0 a_n2750_n2688# 0.799397f
C232 minus.n23 a_n2750_n2688# 0.343379f
C233 minus.n24 a_n2750_n2688# 0.038714f
C234 minus.t1 a_n2750_n2688# 0.799397f
C235 minus.n25 a_n2750_n2688# 0.332327f
C236 minus.n26 a_n2750_n2688# 0.222046f
C237 minus.t14 a_n2750_n2688# 0.820079f
C238 minus.n27 a_n2750_n2688# 0.318496f
C239 minus.t2 a_n2750_n2688# 0.799397f
C240 minus.n28 a_n2750_n2688# 0.343683f
C241 minus.t7 a_n2750_n2688# 0.799397f
C242 minus.n29 a_n2750_n2688# 0.343379f
C243 minus.n30 a_n2750_n2688# 0.008785f
C244 minus.n31 a_n2750_n2688# 0.05166f
C245 minus.n32 a_n2750_n2688# 0.038714f
C246 minus.n33 a_n2750_n2688# 0.038714f
C247 minus.n34 a_n2750_n2688# 0.008785f
C248 minus.t12 a_n2750_n2688# 0.799397f
C249 minus.n35 a_n2750_n2688# 0.332327f
C250 minus.n36 a_n2750_n2688# 0.008785f
C251 minus.n37 a_n2750_n2688# 0.05166f
C252 minus.n38 a_n2750_n2688# 0.064484f
C253 minus.n39 a_n2750_n2688# 0.064484f
C254 minus.t5 a_n2750_n2688# 0.799397f
C255 minus.n40 a_n2750_n2688# 0.342902f
C256 minus.n41 a_n2750_n2688# 0.008785f
C257 minus.t15 a_n2750_n2688# 0.799397f
C258 minus.n42 a_n2750_n2688# 0.328866f
C259 minus.n43 a_n2750_n2688# 0.267212f
C260 minus.n44 a_n2750_n2688# 1.74498f
.ends

