* NGSPICE file created from diffpair580.ext - technology: sky130A

.subckt diffpair580 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.25
X1 a_n948_n4892# a_n948_n4892# a_n948_n4892# a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X2 a_n948_n4892# a_n948_n4892# a_n948_n4892# a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X3 drain_left.t1 plus.t0 source.t0 a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.25
X4 drain_right.t0 minus.t1 source.t3 a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.25
X5 drain_left.t0 plus.t1 source.t1 a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.25
X6 a_n948_n4892# a_n948_n4892# a_n948_n4892# a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X7 a_n948_n4892# a_n948_n4892# a_n948_n4892# a_n948_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
R0 minus.n0 minus.t0 2277.37
R1 minus.n0 minus.t1 2245.08
R2 minus minus.n0 0.188
R3 source.n0 source.t1 44.1297
R4 source.n1 source.t2 44.1296
R5 source.n3 source.t3 44.1295
R6 source.n2 source.t0 44.1295
R7 source.n2 source.n1 28.3635
R8 source.n4 source.n0 22.3506
R9 source.n4 source.n3 5.51343
R10 source.n1 source.n0 0.720328
R11 source.n3 source.n2 0.720328
R12 source source.n4 0.188
R13 drain_right drain_right.t0 94.392
R14 drain_right drain_right.t1 66.7112
R15 plus plus.t0 2268.22
R16 plus plus.t1 2253.75
R17 drain_left drain_left.t1 94.9452
R18 drain_left drain_left.t0 66.9612
C0 source plus 1.1545f
C1 drain_right source 11.6436f
C2 drain_left plus 2.2171f
C3 drain_right drain_left 0.425393f
C4 minus plus 5.82481f
C5 drain_right minus 2.13608f
C6 drain_right plus 0.243802f
C7 source drain_left 11.66f
C8 source minus 1.13933f
C9 drain_left minus 0.171641f
C10 drain_right a_n948_n4892# 9.32432f
C11 drain_left a_n948_n4892# 9.52006f
C12 source a_n948_n4892# 8.450951f
C13 minus a_n948_n4892# 4.177542f
C14 plus a_n948_n4892# 10.188411f
C15 drain_left.t1 a_n948_n4892# 5.02002f
C16 drain_left.t0 a_n948_n4892# 4.46697f
C17 plus.t1 a_n948_n4892# 0.903819f
C18 plus.t0 a_n948_n4892# 0.923996f
C19 drain_right.t0 a_n948_n4892# 4.95729f
C20 drain_right.t1 a_n948_n4892# 4.4316f
C21 source.t1 a_n948_n4892# 3.79737f
C22 source.n0 a_n948_n4892# 1.62669f
C23 source.t2 a_n948_n4892# 3.79738f
C24 source.n1 a_n948_n4892# 2.03197f
C25 source.t0 a_n948_n4892# 3.79736f
C26 source.n2 a_n948_n4892# 2.03199f
C27 source.t3 a_n948_n4892# 3.79736f
C28 source.n3 a_n948_n4892# 0.492355f
C29 source.n4 a_n948_n4892# 1.89214f
C30 minus.t0 a_n948_n4892# 0.915557f
C31 minus.t1 a_n948_n4892# 0.872816f
C32 minus.n0 a_n948_n4892# 6.07226f
.ends

