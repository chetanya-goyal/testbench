* NGSPICE file created from diffpair39.ext - technology: sky130A

.subckt diffpair39 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t23 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 source.t20 plus.t0 drain_left.t23 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X2 drain_left.t22 plus.t1 source.t19 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 drain_left.t21 plus.t2 source.t18 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 source.t46 minus.t1 drain_right.t2 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X5 drain_right.t20 minus.t2 source.t45 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X6 drain_right.t19 minus.t3 source.t44 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X7 source.t43 minus.t4 drain_right.t9 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X8 drain_right.t21 minus.t5 source.t42 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X9 source.t41 minus.t6 drain_right.t12 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X10 source.t17 plus.t3 drain_left.t20 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X11 source.t16 plus.t4 drain_left.t19 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X12 source.t21 plus.t5 drain_left.t18 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X13 source.t23 plus.t6 drain_left.t17 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X14 source.t40 minus.t7 drain_right.t22 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X15 drain_right.t3 minus.t8 source.t39 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X16 drain_left.t16 plus.t7 source.t22 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X17 drain_right.t7 minus.t9 source.t38 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X18 drain_left.t15 plus.t8 source.t13 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X19 drain_left.t14 plus.t9 source.t12 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X20 a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X21 drain_right.t18 minus.t10 source.t37 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X22 source.t36 minus.t11 drain_right.t0 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 source.t35 minus.t12 drain_right.t16 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X24 source.t6 plus.t10 drain_left.t13 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X25 source.t11 plus.t11 drain_left.t12 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X26 a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X27 drain_left.t11 plus.t12 source.t3 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X28 drain_left.t10 plus.t13 source.t5 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X29 drain_left.t9 plus.t14 source.t8 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X30 source.t34 minus.t13 drain_right.t4 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X31 source.t10 plus.t15 drain_left.t8 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X32 drain_right.t15 minus.t14 source.t33 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X33 drain_right.t17 minus.t15 source.t32 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X34 source.t31 minus.t16 drain_right.t10 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X35 drain_left.t7 plus.t16 source.t1 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X36 a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X37 source.t2 plus.t17 drain_left.t6 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X38 source.t4 plus.t18 drain_left.t5 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X39 drain_right.t1 minus.t17 source.t30 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X40 drain_left.t4 plus.t19 source.t7 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X41 drain_left.t3 plus.t20 source.t9 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X42 drain_right.t5 minus.t18 source.t29 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X43 drain_right.t14 minus.t19 source.t28 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X44 a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X45 drain_right.t11 minus.t20 source.t27 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X46 source.t26 minus.t21 drain_right.t6 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X47 source.t25 minus.t22 drain_right.t8 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X48 source.t24 minus.t23 drain_right.t13 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X49 source.t14 plus.t21 drain_left.t2 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X50 source.t0 plus.t22 drain_left.t1 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X51 drain_left.t0 plus.t23 source.t15 a_n2354_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
R0 minus.n35 minus.t4 216.171
R1 minus.n9 minus.t15 216.171
R2 minus.n72 minus.t14 216.171
R3 minus.n46 minus.t16 216.171
R4 minus.n34 minus.t19 184.768
R5 minus.n1 minus.t11 184.768
R6 minus.n28 minus.t3 184.768
R7 minus.n26 minus.t22 184.768
R8 minus.n3 minus.t10 184.768
R9 minus.n20 minus.t1 184.768
R10 minus.n5 minus.t18 184.768
R11 minus.n15 minus.t13 184.768
R12 minus.n13 minus.t2 184.768
R13 minus.n8 minus.t21 184.768
R14 minus.n71 minus.t0 184.768
R15 minus.n38 minus.t5 184.768
R16 minus.n65 minus.t7 184.768
R17 minus.n63 minus.t20 184.768
R18 minus.n40 minus.t23 184.768
R19 minus.n57 minus.t9 184.768
R20 minus.n42 minus.t12 184.768
R21 minus.n52 minus.t17 184.768
R22 minus.n50 minus.t6 184.768
R23 minus.n45 minus.t8 184.768
R24 minus.n10 minus.n9 161.489
R25 minus.n47 minus.n46 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n32 minus.n31 161.3
R29 minus.n30 minus.n29 161.3
R30 minus.n27 minus.n2 161.3
R31 minus.n25 minus.n24 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n19 minus.n18 161.3
R35 minus.n17 minus.n16 161.3
R36 minus.n14 minus.n6 161.3
R37 minus.n12 minus.n11 161.3
R38 minus.n10 minus.n7 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n69 minus.n68 161.3
R42 minus.n67 minus.n66 161.3
R43 minus.n64 minus.n39 161.3
R44 minus.n62 minus.n61 161.3
R45 minus.n60 minus.n59 161.3
R46 minus.n58 minus.n41 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n54 minus.n53 161.3
R49 minus.n51 minus.n43 161.3
R50 minus.n49 minus.n48 161.3
R51 minus.n47 minus.n44 161.3
R52 minus.n33 minus.n32 73.0308
R53 minus.n22 minus.n21 73.0308
R54 minus.n12 minus.n7 73.0308
R55 minus.n49 minus.n44 73.0308
R56 minus.n59 minus.n58 73.0308
R57 minus.n70 minus.n69 73.0308
R58 minus.n29 minus.n1 66.4581
R59 minus.n14 minus.n13 66.4581
R60 minus.n51 minus.n50 66.4581
R61 minus.n66 minus.n38 66.4581
R62 minus.n25 minus.n3 63.5369
R63 minus.n20 minus.n19 63.5369
R64 minus.n57 minus.n56 63.5369
R65 minus.n62 minus.n40 63.5369
R66 minus.n35 minus.n34 60.6157
R67 minus.n9 minus.n8 60.6157
R68 minus.n46 minus.n45 60.6157
R69 minus.n72 minus.n71 60.6157
R70 minus.n28 minus.n27 47.4702
R71 minus.n16 minus.n15 47.4702
R72 minus.n53 minus.n52 47.4702
R73 minus.n65 minus.n64 47.4702
R74 minus.n27 minus.n26 44.549
R75 minus.n16 minus.n5 44.549
R76 minus.n53 minus.n42 44.549
R77 minus.n64 minus.n63 44.549
R78 minus.n74 minus.n36 29.6747
R79 minus.n26 minus.n25 28.4823
R80 minus.n19 minus.n5 28.4823
R81 minus.n56 minus.n42 28.4823
R82 minus.n63 minus.n62 28.4823
R83 minus.n29 minus.n28 25.5611
R84 minus.n15 minus.n14 25.5611
R85 minus.n52 minus.n51 25.5611
R86 minus.n66 minus.n65 25.5611
R87 minus.n34 minus.n33 12.4157
R88 minus.n8 minus.n7 12.4157
R89 minus.n45 minus.n44 12.4157
R90 minus.n71 minus.n70 12.4157
R91 minus.n22 minus.n3 9.49444
R92 minus.n21 minus.n20 9.49444
R93 minus.n58 minus.n57 9.49444
R94 minus.n59 minus.n40 9.49444
R95 minus.n32 minus.n1 6.57323
R96 minus.n13 minus.n12 6.57323
R97 minus.n50 minus.n49 6.57323
R98 minus.n69 minus.n38 6.57323
R99 minus.n74 minus.n73 6.4702
R100 minus.n36 minus.n0 0.189894
R101 minus.n31 minus.n0 0.189894
R102 minus.n31 minus.n30 0.189894
R103 minus.n30 minus.n2 0.189894
R104 minus.n24 minus.n2 0.189894
R105 minus.n24 minus.n23 0.189894
R106 minus.n23 minus.n4 0.189894
R107 minus.n18 minus.n4 0.189894
R108 minus.n18 minus.n17 0.189894
R109 minus.n17 minus.n6 0.189894
R110 minus.n11 minus.n6 0.189894
R111 minus.n11 minus.n10 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n48 minus.n43 0.189894
R114 minus.n54 minus.n43 0.189894
R115 minus.n55 minus.n54 0.189894
R116 minus.n55 minus.n41 0.189894
R117 minus.n60 minus.n41 0.189894
R118 minus.n61 minus.n60 0.189894
R119 minus.n61 minus.n39 0.189894
R120 minus.n67 minus.n39 0.189894
R121 minus.n68 minus.n67 0.189894
R122 minus.n68 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 drain_right.n13 drain_right.n11 240.675
R126 drain_right.n7 drain_right.n5 240.674
R127 drain_right.n2 drain_right.n0 240.674
R128 drain_right.n13 drain_right.n12 240.132
R129 drain_right.n15 drain_right.n14 240.132
R130 drain_right.n17 drain_right.n16 240.132
R131 drain_right.n19 drain_right.n18 240.132
R132 drain_right.n21 drain_right.n20 240.132
R133 drain_right.n7 drain_right.n6 240.131
R134 drain_right.n9 drain_right.n8 240.131
R135 drain_right.n4 drain_right.n3 240.131
R136 drain_right.n2 drain_right.n1 240.131
R137 drain_right drain_right.n10 23.64
R138 drain_right.n5 drain_right.t23 19.8005
R139 drain_right.n5 drain_right.t15 19.8005
R140 drain_right.n6 drain_right.t22 19.8005
R141 drain_right.n6 drain_right.t21 19.8005
R142 drain_right.n8 drain_right.t13 19.8005
R143 drain_right.n8 drain_right.t11 19.8005
R144 drain_right.n3 drain_right.t16 19.8005
R145 drain_right.n3 drain_right.t7 19.8005
R146 drain_right.n1 drain_right.t12 19.8005
R147 drain_right.n1 drain_right.t1 19.8005
R148 drain_right.n0 drain_right.t10 19.8005
R149 drain_right.n0 drain_right.t3 19.8005
R150 drain_right.n11 drain_right.t6 19.8005
R151 drain_right.n11 drain_right.t17 19.8005
R152 drain_right.n12 drain_right.t4 19.8005
R153 drain_right.n12 drain_right.t20 19.8005
R154 drain_right.n14 drain_right.t2 19.8005
R155 drain_right.n14 drain_right.t5 19.8005
R156 drain_right.n16 drain_right.t8 19.8005
R157 drain_right.n16 drain_right.t18 19.8005
R158 drain_right.n18 drain_right.t0 19.8005
R159 drain_right.n18 drain_right.t19 19.8005
R160 drain_right.n20 drain_right.t9 19.8005
R161 drain_right.n20 drain_right.t14 19.8005
R162 drain_right drain_right.n21 6.19632
R163 drain_right.n9 drain_right.n7 0.543603
R164 drain_right.n4 drain_right.n2 0.543603
R165 drain_right.n21 drain_right.n19 0.543603
R166 drain_right.n19 drain_right.n17 0.543603
R167 drain_right.n17 drain_right.n15 0.543603
R168 drain_right.n15 drain_right.n13 0.543603
R169 drain_right.n10 drain_right.n9 0.216706
R170 drain_right.n10 drain_right.n4 0.216706
R171 source.n0 source.t22 243.255
R172 source.n11 source.t23 243.255
R173 source.n12 source.t32 243.255
R174 source.n23 source.t43 243.255
R175 source.n47 source.t33 243.254
R176 source.n36 source.t31 243.254
R177 source.n35 source.t5 243.254
R178 source.n24 source.t21 243.254
R179 source.n2 source.n1 223.454
R180 source.n4 source.n3 223.454
R181 source.n6 source.n5 223.454
R182 source.n8 source.n7 223.454
R183 source.n10 source.n9 223.454
R184 source.n14 source.n13 223.454
R185 source.n16 source.n15 223.454
R186 source.n18 source.n17 223.454
R187 source.n20 source.n19 223.454
R188 source.n22 source.n21 223.454
R189 source.n46 source.n45 223.453
R190 source.n44 source.n43 223.453
R191 source.n42 source.n41 223.453
R192 source.n40 source.n39 223.453
R193 source.n38 source.n37 223.453
R194 source.n34 source.n33 223.453
R195 source.n32 source.n31 223.453
R196 source.n30 source.n29 223.453
R197 source.n28 source.n27 223.453
R198 source.n26 source.n25 223.453
R199 source.n45 source.t42 19.8005
R200 source.n45 source.t47 19.8005
R201 source.n43 source.t27 19.8005
R202 source.n43 source.t40 19.8005
R203 source.n41 source.t38 19.8005
R204 source.n41 source.t24 19.8005
R205 source.n39 source.t30 19.8005
R206 source.n39 source.t35 19.8005
R207 source.n37 source.t39 19.8005
R208 source.n37 source.t41 19.8005
R209 source.n33 source.t19 19.8005
R210 source.n33 source.t17 19.8005
R211 source.n31 source.t13 19.8005
R212 source.n31 source.t2 19.8005
R213 source.n29 source.t7 19.8005
R214 source.n29 source.t16 19.8005
R215 source.n27 source.t12 19.8005
R216 source.n27 source.t6 19.8005
R217 source.n25 source.t8 19.8005
R218 source.n25 source.t14 19.8005
R219 source.n1 source.t9 19.8005
R220 source.n1 source.t20 19.8005
R221 source.n3 source.t18 19.8005
R222 source.n3 source.t10 19.8005
R223 source.n5 source.t1 19.8005
R224 source.n5 source.t0 19.8005
R225 source.n7 source.t15 19.8005
R226 source.n7 source.t11 19.8005
R227 source.n9 source.t3 19.8005
R228 source.n9 source.t4 19.8005
R229 source.n13 source.t45 19.8005
R230 source.n13 source.t26 19.8005
R231 source.n15 source.t29 19.8005
R232 source.n15 source.t34 19.8005
R233 source.n17 source.t37 19.8005
R234 source.n17 source.t46 19.8005
R235 source.n19 source.t44 19.8005
R236 source.n19 source.t25 19.8005
R237 source.n21 source.t28 19.8005
R238 source.n21 source.t36 19.8005
R239 source.n24 source.n23 13.4975
R240 source.n48 source.n0 7.96301
R241 source.n48 source.n47 5.53498
R242 source.n23 source.n22 0.543603
R243 source.n22 source.n20 0.543603
R244 source.n20 source.n18 0.543603
R245 source.n18 source.n16 0.543603
R246 source.n16 source.n14 0.543603
R247 source.n14 source.n12 0.543603
R248 source.n11 source.n10 0.543603
R249 source.n10 source.n8 0.543603
R250 source.n8 source.n6 0.543603
R251 source.n6 source.n4 0.543603
R252 source.n4 source.n2 0.543603
R253 source.n2 source.n0 0.543603
R254 source.n26 source.n24 0.543603
R255 source.n28 source.n26 0.543603
R256 source.n30 source.n28 0.543603
R257 source.n32 source.n30 0.543603
R258 source.n34 source.n32 0.543603
R259 source.n35 source.n34 0.543603
R260 source.n38 source.n36 0.543603
R261 source.n40 source.n38 0.543603
R262 source.n42 source.n40 0.543603
R263 source.n44 source.n42 0.543603
R264 source.n46 source.n44 0.543603
R265 source.n47 source.n46 0.543603
R266 source.n12 source.n11 0.470328
R267 source.n36 source.n35 0.470328
R268 source source.n48 0.188
R269 plus.n9 plus.t6 216.171
R270 plus.n35 plus.t7 216.171
R271 plus.n46 plus.t13 216.171
R272 plus.n72 plus.t5 216.171
R273 plus.n8 plus.t12 184.768
R274 plus.n13 plus.t18 184.768
R275 plus.n15 plus.t23 184.768
R276 plus.n5 plus.t11 184.768
R277 plus.n20 plus.t16 184.768
R278 plus.n3 plus.t22 184.768
R279 plus.n26 plus.t2 184.768
R280 plus.n28 plus.t15 184.768
R281 plus.n1 plus.t20 184.768
R282 plus.n34 plus.t0 184.768
R283 plus.n45 plus.t3 184.768
R284 plus.n50 plus.t1 184.768
R285 plus.n52 plus.t17 184.768
R286 plus.n42 plus.t8 184.768
R287 plus.n57 plus.t4 184.768
R288 plus.n40 plus.t19 184.768
R289 plus.n63 plus.t10 184.768
R290 plus.n65 plus.t9 184.768
R291 plus.n38 plus.t21 184.768
R292 plus.n71 plus.t14 184.768
R293 plus.n10 plus.n9 161.489
R294 plus.n47 plus.n46 161.489
R295 plus.n10 plus.n7 161.3
R296 plus.n12 plus.n11 161.3
R297 plus.n14 plus.n6 161.3
R298 plus.n17 plus.n16 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n21 plus.n4 161.3
R301 plus.n23 plus.n22 161.3
R302 plus.n25 plus.n24 161.3
R303 plus.n27 plus.n2 161.3
R304 plus.n30 plus.n29 161.3
R305 plus.n32 plus.n31 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n47 plus.n44 161.3
R309 plus.n49 plus.n48 161.3
R310 plus.n51 plus.n43 161.3
R311 plus.n54 plus.n53 161.3
R312 plus.n56 plus.n55 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n61 161.3
R316 plus.n64 plus.n39 161.3
R317 plus.n67 plus.n66 161.3
R318 plus.n69 plus.n68 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n12 plus.n7 73.0308
R322 plus.n22 plus.n21 73.0308
R323 plus.n33 plus.n32 73.0308
R324 plus.n70 plus.n69 73.0308
R325 plus.n59 plus.n58 73.0308
R326 plus.n49 plus.n44 73.0308
R327 plus.n14 plus.n13 66.4581
R328 plus.n29 plus.n1 66.4581
R329 plus.n66 plus.n38 66.4581
R330 plus.n51 plus.n50 66.4581
R331 plus.n20 plus.n19 63.5369
R332 plus.n25 plus.n3 63.5369
R333 plus.n62 plus.n40 63.5369
R334 plus.n57 plus.n56 63.5369
R335 plus.n9 plus.n8 60.6157
R336 plus.n35 plus.n34 60.6157
R337 plus.n72 plus.n71 60.6157
R338 plus.n46 plus.n45 60.6157
R339 plus.n16 plus.n15 47.4702
R340 plus.n28 plus.n27 47.4702
R341 plus.n65 plus.n64 47.4702
R342 plus.n53 plus.n52 47.4702
R343 plus.n16 plus.n5 44.549
R344 plus.n27 plus.n26 44.549
R345 plus.n64 plus.n63 44.549
R346 plus.n53 plus.n42 44.549
R347 plus.n19 plus.n5 28.4823
R348 plus.n26 plus.n25 28.4823
R349 plus.n63 plus.n62 28.4823
R350 plus.n56 plus.n42 28.4823
R351 plus plus.n73 27.7225
R352 plus.n15 plus.n14 25.5611
R353 plus.n29 plus.n28 25.5611
R354 plus.n66 plus.n65 25.5611
R355 plus.n52 plus.n51 25.5611
R356 plus.n8 plus.n7 12.4157
R357 plus.n34 plus.n33 12.4157
R358 plus.n71 plus.n70 12.4157
R359 plus.n45 plus.n44 12.4157
R360 plus.n21 plus.n20 9.49444
R361 plus.n22 plus.n3 9.49444
R362 plus.n59 plus.n40 9.49444
R363 plus.n58 plus.n57 9.49444
R364 plus plus.n36 7.94747
R365 plus.n13 plus.n12 6.57323
R366 plus.n32 plus.n1 6.57323
R367 plus.n69 plus.n38 6.57323
R368 plus.n50 plus.n49 6.57323
R369 plus.n11 plus.n10 0.189894
R370 plus.n11 plus.n6 0.189894
R371 plus.n17 plus.n6 0.189894
R372 plus.n18 plus.n17 0.189894
R373 plus.n18 plus.n4 0.189894
R374 plus.n23 plus.n4 0.189894
R375 plus.n24 plus.n23 0.189894
R376 plus.n24 plus.n2 0.189894
R377 plus.n30 plus.n2 0.189894
R378 plus.n31 plus.n30 0.189894
R379 plus.n31 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n68 plus.n37 0.189894
R383 plus.n68 plus.n67 0.189894
R384 plus.n67 plus.n39 0.189894
R385 plus.n61 plus.n39 0.189894
R386 plus.n61 plus.n60 0.189894
R387 plus.n60 plus.n41 0.189894
R388 plus.n55 plus.n41 0.189894
R389 plus.n55 plus.n54 0.189894
R390 plus.n54 plus.n43 0.189894
R391 plus.n48 plus.n43 0.189894
R392 plus.n48 plus.n47 0.189894
R393 drain_left.n13 drain_left.n11 240.675
R394 drain_left.n7 drain_left.n5 240.674
R395 drain_left.n2 drain_left.n0 240.674
R396 drain_left.n21 drain_left.n20 240.132
R397 drain_left.n19 drain_left.n18 240.132
R398 drain_left.n17 drain_left.n16 240.132
R399 drain_left.n15 drain_left.n14 240.132
R400 drain_left.n13 drain_left.n12 240.132
R401 drain_left.n7 drain_left.n6 240.131
R402 drain_left.n9 drain_left.n8 240.131
R403 drain_left.n4 drain_left.n3 240.131
R404 drain_left.n2 drain_left.n1 240.131
R405 drain_left drain_left.n10 24.1932
R406 drain_left.n5 drain_left.t20 19.8005
R407 drain_left.n5 drain_left.t10 19.8005
R408 drain_left.n6 drain_left.t6 19.8005
R409 drain_left.n6 drain_left.t22 19.8005
R410 drain_left.n8 drain_left.t19 19.8005
R411 drain_left.n8 drain_left.t15 19.8005
R412 drain_left.n3 drain_left.t13 19.8005
R413 drain_left.n3 drain_left.t4 19.8005
R414 drain_left.n1 drain_left.t2 19.8005
R415 drain_left.n1 drain_left.t14 19.8005
R416 drain_left.n0 drain_left.t18 19.8005
R417 drain_left.n0 drain_left.t9 19.8005
R418 drain_left.n20 drain_left.t23 19.8005
R419 drain_left.n20 drain_left.t16 19.8005
R420 drain_left.n18 drain_left.t8 19.8005
R421 drain_left.n18 drain_left.t3 19.8005
R422 drain_left.n16 drain_left.t1 19.8005
R423 drain_left.n16 drain_left.t21 19.8005
R424 drain_left.n14 drain_left.t12 19.8005
R425 drain_left.n14 drain_left.t7 19.8005
R426 drain_left.n12 drain_left.t5 19.8005
R427 drain_left.n12 drain_left.t0 19.8005
R428 drain_left.n11 drain_left.t17 19.8005
R429 drain_left.n11 drain_left.t11 19.8005
R430 drain_left drain_left.n21 6.19632
R431 drain_left.n9 drain_left.n7 0.543603
R432 drain_left.n4 drain_left.n2 0.543603
R433 drain_left.n15 drain_left.n13 0.543603
R434 drain_left.n17 drain_left.n15 0.543603
R435 drain_left.n19 drain_left.n17 0.543603
R436 drain_left.n21 drain_left.n19 0.543603
R437 drain_left.n10 drain_left.n9 0.216706
R438 drain_left.n10 drain_left.n4 0.216706
C0 drain_left plus 1.55441f
C1 plus drain_right 0.396707f
C2 drain_left drain_right 1.26603f
C3 plus minus 4.06701f
C4 drain_left minus 0.180087f
C5 drain_right minus 1.32237f
C6 plus source 1.78093f
C7 drain_left source 7.1944f
C8 drain_right source 7.19503f
C9 minus source 1.76706f
C10 drain_right a_n2354_n1088# 4.46788f
C11 drain_left a_n2354_n1088# 4.78248f
C12 source a_n2354_n1088# 2.765402f
C13 minus a_n2354_n1088# 8.372579f
C14 plus a_n2354_n1088# 9.037783f
C15 drain_left.t18 a_n2354_n1088# 0.020469f
C16 drain_left.t9 a_n2354_n1088# 0.020469f
C17 drain_left.n0 a_n2354_n1088# 0.080172f
C18 drain_left.t2 a_n2354_n1088# 0.020469f
C19 drain_left.t14 a_n2354_n1088# 0.020469f
C20 drain_left.n1 a_n2354_n1088# 0.079535f
C21 drain_left.n2 a_n2354_n1088# 0.553383f
C22 drain_left.t13 a_n2354_n1088# 0.020469f
C23 drain_left.t4 a_n2354_n1088# 0.020469f
C24 drain_left.n3 a_n2354_n1088# 0.079535f
C25 drain_left.n4 a_n2354_n1088# 0.247287f
C26 drain_left.t20 a_n2354_n1088# 0.020469f
C27 drain_left.t10 a_n2354_n1088# 0.020469f
C28 drain_left.n5 a_n2354_n1088# 0.080172f
C29 drain_left.t6 a_n2354_n1088# 0.020469f
C30 drain_left.t22 a_n2354_n1088# 0.020469f
C31 drain_left.n6 a_n2354_n1088# 0.079535f
C32 drain_left.n7 a_n2354_n1088# 0.553383f
C33 drain_left.t19 a_n2354_n1088# 0.020469f
C34 drain_left.t15 a_n2354_n1088# 0.020469f
C35 drain_left.n8 a_n2354_n1088# 0.079535f
C36 drain_left.n9 a_n2354_n1088# 0.247287f
C37 drain_left.n10 a_n2354_n1088# 0.824972f
C38 drain_left.t17 a_n2354_n1088# 0.020469f
C39 drain_left.t11 a_n2354_n1088# 0.020469f
C40 drain_left.n11 a_n2354_n1088# 0.080172f
C41 drain_left.t5 a_n2354_n1088# 0.020469f
C42 drain_left.t0 a_n2354_n1088# 0.020469f
C43 drain_left.n12 a_n2354_n1088# 0.079535f
C44 drain_left.n13 a_n2354_n1088# 0.553383f
C45 drain_left.t12 a_n2354_n1088# 0.020469f
C46 drain_left.t7 a_n2354_n1088# 0.020469f
C47 drain_left.n14 a_n2354_n1088# 0.079535f
C48 drain_left.n15 a_n2354_n1088# 0.271794f
C49 drain_left.t1 a_n2354_n1088# 0.020469f
C50 drain_left.t21 a_n2354_n1088# 0.020469f
C51 drain_left.n16 a_n2354_n1088# 0.079535f
C52 drain_left.n17 a_n2354_n1088# 0.271794f
C53 drain_left.t8 a_n2354_n1088# 0.020469f
C54 drain_left.t3 a_n2354_n1088# 0.020469f
C55 drain_left.n18 a_n2354_n1088# 0.079535f
C56 drain_left.n19 a_n2354_n1088# 0.271794f
C57 drain_left.t23 a_n2354_n1088# 0.020469f
C58 drain_left.t16 a_n2354_n1088# 0.020469f
C59 drain_left.n20 a_n2354_n1088# 0.079535f
C60 drain_left.n21 a_n2354_n1088# 0.487393f
C61 plus.n0 a_n2354_n1088# 0.028362f
C62 plus.t0 a_n2354_n1088# 0.02623f
C63 plus.t20 a_n2354_n1088# 0.02623f
C64 plus.n1 a_n2354_n1088# 0.027024f
C65 plus.n2 a_n2354_n1088# 0.028362f
C66 plus.t15 a_n2354_n1088# 0.02623f
C67 plus.t2 a_n2354_n1088# 0.02623f
C68 plus.t22 a_n2354_n1088# 0.02623f
C69 plus.n3 a_n2354_n1088# 0.027024f
C70 plus.n4 a_n2354_n1088# 0.028362f
C71 plus.t16 a_n2354_n1088# 0.02623f
C72 plus.t11 a_n2354_n1088# 0.02623f
C73 plus.n5 a_n2354_n1088# 0.027024f
C74 plus.n6 a_n2354_n1088# 0.028362f
C75 plus.t23 a_n2354_n1088# 0.02623f
C76 plus.t18 a_n2354_n1088# 0.02623f
C77 plus.n7 a_n2354_n1088# 0.010895f
C78 plus.t6 a_n2354_n1088# 0.030194f
C79 plus.t12 a_n2354_n1088# 0.02623f
C80 plus.n8 a_n2354_n1088# 0.027024f
C81 plus.n9 a_n2354_n1088# 0.035043f
C82 plus.n10 a_n2354_n1088# 0.060708f
C83 plus.n11 a_n2354_n1088# 0.028362f
C84 plus.n12 a_n2354_n1088# 0.010196f
C85 plus.n13 a_n2354_n1088# 0.027024f
C86 plus.n14 a_n2354_n1088# 0.011682f
C87 plus.n15 a_n2354_n1088# 0.027024f
C88 plus.n16 a_n2354_n1088# 0.011682f
C89 plus.n17 a_n2354_n1088# 0.028362f
C90 plus.n18 a_n2354_n1088# 0.028362f
C91 plus.n19 a_n2354_n1088# 0.011682f
C92 plus.n20 a_n2354_n1088# 0.027024f
C93 plus.n21 a_n2354_n1088# 0.010545f
C94 plus.n22 a_n2354_n1088# 0.010545f
C95 plus.n23 a_n2354_n1088# 0.028362f
C96 plus.n24 a_n2354_n1088# 0.028362f
C97 plus.n25 a_n2354_n1088# 0.011682f
C98 plus.n26 a_n2354_n1088# 0.027024f
C99 plus.n27 a_n2354_n1088# 0.011682f
C100 plus.n28 a_n2354_n1088# 0.027024f
C101 plus.n29 a_n2354_n1088# 0.011682f
C102 plus.n30 a_n2354_n1088# 0.028362f
C103 plus.n31 a_n2354_n1088# 0.028362f
C104 plus.n32 a_n2354_n1088# 0.010196f
C105 plus.n33 a_n2354_n1088# 0.010895f
C106 plus.n34 a_n2354_n1088# 0.027024f
C107 plus.t7 a_n2354_n1088# 0.030194f
C108 plus.n35 a_n2354_n1088# 0.035005f
C109 plus.n36 a_n2354_n1088# 0.192348f
C110 plus.n37 a_n2354_n1088# 0.028362f
C111 plus.t5 a_n2354_n1088# 0.030194f
C112 plus.t14 a_n2354_n1088# 0.02623f
C113 plus.t21 a_n2354_n1088# 0.02623f
C114 plus.n38 a_n2354_n1088# 0.027024f
C115 plus.n39 a_n2354_n1088# 0.028362f
C116 plus.t9 a_n2354_n1088# 0.02623f
C117 plus.t10 a_n2354_n1088# 0.02623f
C118 plus.t19 a_n2354_n1088# 0.02623f
C119 plus.n40 a_n2354_n1088# 0.027024f
C120 plus.n41 a_n2354_n1088# 0.028362f
C121 plus.t4 a_n2354_n1088# 0.02623f
C122 plus.t8 a_n2354_n1088# 0.02623f
C123 plus.n42 a_n2354_n1088# 0.027024f
C124 plus.n43 a_n2354_n1088# 0.028362f
C125 plus.t17 a_n2354_n1088# 0.02623f
C126 plus.t1 a_n2354_n1088# 0.02623f
C127 plus.n44 a_n2354_n1088# 0.010895f
C128 plus.t3 a_n2354_n1088# 0.02623f
C129 plus.n45 a_n2354_n1088# 0.027024f
C130 plus.t13 a_n2354_n1088# 0.030194f
C131 plus.n46 a_n2354_n1088# 0.035043f
C132 plus.n47 a_n2354_n1088# 0.060708f
C133 plus.n48 a_n2354_n1088# 0.028362f
C134 plus.n49 a_n2354_n1088# 0.010196f
C135 plus.n50 a_n2354_n1088# 0.027024f
C136 plus.n51 a_n2354_n1088# 0.011682f
C137 plus.n52 a_n2354_n1088# 0.027024f
C138 plus.n53 a_n2354_n1088# 0.011682f
C139 plus.n54 a_n2354_n1088# 0.028362f
C140 plus.n55 a_n2354_n1088# 0.028362f
C141 plus.n56 a_n2354_n1088# 0.011682f
C142 plus.n57 a_n2354_n1088# 0.027024f
C143 plus.n58 a_n2354_n1088# 0.010545f
C144 plus.n59 a_n2354_n1088# 0.010545f
C145 plus.n60 a_n2354_n1088# 0.028362f
C146 plus.n61 a_n2354_n1088# 0.028362f
C147 plus.n62 a_n2354_n1088# 0.011682f
C148 plus.n63 a_n2354_n1088# 0.027024f
C149 plus.n64 a_n2354_n1088# 0.011682f
C150 plus.n65 a_n2354_n1088# 0.027024f
C151 plus.n66 a_n2354_n1088# 0.011682f
C152 plus.n67 a_n2354_n1088# 0.028362f
C153 plus.n68 a_n2354_n1088# 0.028362f
C154 plus.n69 a_n2354_n1088# 0.010196f
C155 plus.n70 a_n2354_n1088# 0.010895f
C156 plus.n71 a_n2354_n1088# 0.027024f
C157 plus.n72 a_n2354_n1088# 0.035005f
C158 plus.n73 a_n2354_n1088# 0.6984f
C159 source.t22 a_n2354_n1088# 0.137753f
C160 source.n0 a_n2354_n1088# 0.59149f
C161 source.t9 a_n2354_n1088# 0.02475f
C162 source.t20 a_n2354_n1088# 0.02475f
C163 source.n1 a_n2354_n1088# 0.080267f
C164 source.n2 a_n2354_n1088# 0.301973f
C165 source.t18 a_n2354_n1088# 0.02475f
C166 source.t10 a_n2354_n1088# 0.02475f
C167 source.n3 a_n2354_n1088# 0.080267f
C168 source.n4 a_n2354_n1088# 0.301973f
C169 source.t1 a_n2354_n1088# 0.02475f
C170 source.t0 a_n2354_n1088# 0.02475f
C171 source.n5 a_n2354_n1088# 0.080267f
C172 source.n6 a_n2354_n1088# 0.301973f
C173 source.t15 a_n2354_n1088# 0.02475f
C174 source.t11 a_n2354_n1088# 0.02475f
C175 source.n7 a_n2354_n1088# 0.080267f
C176 source.n8 a_n2354_n1088# 0.301973f
C177 source.t3 a_n2354_n1088# 0.02475f
C178 source.t4 a_n2354_n1088# 0.02475f
C179 source.n9 a_n2354_n1088# 0.080267f
C180 source.n10 a_n2354_n1088# 0.301973f
C181 source.t23 a_n2354_n1088# 0.137753f
C182 source.n11 a_n2354_n1088# 0.304591f
C183 source.t32 a_n2354_n1088# 0.137753f
C184 source.n12 a_n2354_n1088# 0.304591f
C185 source.t45 a_n2354_n1088# 0.02475f
C186 source.t26 a_n2354_n1088# 0.02475f
C187 source.n13 a_n2354_n1088# 0.080267f
C188 source.n14 a_n2354_n1088# 0.301973f
C189 source.t29 a_n2354_n1088# 0.02475f
C190 source.t34 a_n2354_n1088# 0.02475f
C191 source.n15 a_n2354_n1088# 0.080267f
C192 source.n16 a_n2354_n1088# 0.301973f
C193 source.t37 a_n2354_n1088# 0.02475f
C194 source.t46 a_n2354_n1088# 0.02475f
C195 source.n17 a_n2354_n1088# 0.080267f
C196 source.n18 a_n2354_n1088# 0.301973f
C197 source.t44 a_n2354_n1088# 0.02475f
C198 source.t25 a_n2354_n1088# 0.02475f
C199 source.n19 a_n2354_n1088# 0.080267f
C200 source.n20 a_n2354_n1088# 0.301973f
C201 source.t28 a_n2354_n1088# 0.02475f
C202 source.t36 a_n2354_n1088# 0.02475f
C203 source.n21 a_n2354_n1088# 0.080267f
C204 source.n22 a_n2354_n1088# 0.301973f
C205 source.t43 a_n2354_n1088# 0.137753f
C206 source.n23 a_n2354_n1088# 0.842455f
C207 source.t21 a_n2354_n1088# 0.137753f
C208 source.n24 a_n2354_n1088# 0.842455f
C209 source.t8 a_n2354_n1088# 0.02475f
C210 source.t14 a_n2354_n1088# 0.02475f
C211 source.n25 a_n2354_n1088# 0.080267f
C212 source.n26 a_n2354_n1088# 0.301973f
C213 source.t12 a_n2354_n1088# 0.02475f
C214 source.t6 a_n2354_n1088# 0.02475f
C215 source.n27 a_n2354_n1088# 0.080267f
C216 source.n28 a_n2354_n1088# 0.301973f
C217 source.t7 a_n2354_n1088# 0.02475f
C218 source.t16 a_n2354_n1088# 0.02475f
C219 source.n29 a_n2354_n1088# 0.080267f
C220 source.n30 a_n2354_n1088# 0.301973f
C221 source.t13 a_n2354_n1088# 0.02475f
C222 source.t2 a_n2354_n1088# 0.02475f
C223 source.n31 a_n2354_n1088# 0.080267f
C224 source.n32 a_n2354_n1088# 0.301973f
C225 source.t19 a_n2354_n1088# 0.02475f
C226 source.t17 a_n2354_n1088# 0.02475f
C227 source.n33 a_n2354_n1088# 0.080267f
C228 source.n34 a_n2354_n1088# 0.301973f
C229 source.t5 a_n2354_n1088# 0.137753f
C230 source.n35 a_n2354_n1088# 0.304591f
C231 source.t31 a_n2354_n1088# 0.137753f
C232 source.n36 a_n2354_n1088# 0.304591f
C233 source.t39 a_n2354_n1088# 0.02475f
C234 source.t41 a_n2354_n1088# 0.02475f
C235 source.n37 a_n2354_n1088# 0.080267f
C236 source.n38 a_n2354_n1088# 0.301973f
C237 source.t30 a_n2354_n1088# 0.02475f
C238 source.t35 a_n2354_n1088# 0.02475f
C239 source.n39 a_n2354_n1088# 0.080267f
C240 source.n40 a_n2354_n1088# 0.301973f
C241 source.t38 a_n2354_n1088# 0.02475f
C242 source.t24 a_n2354_n1088# 0.02475f
C243 source.n41 a_n2354_n1088# 0.080267f
C244 source.n42 a_n2354_n1088# 0.301973f
C245 source.t27 a_n2354_n1088# 0.02475f
C246 source.t40 a_n2354_n1088# 0.02475f
C247 source.n43 a_n2354_n1088# 0.080267f
C248 source.n44 a_n2354_n1088# 0.301973f
C249 source.t42 a_n2354_n1088# 0.02475f
C250 source.t47 a_n2354_n1088# 0.02475f
C251 source.n45 a_n2354_n1088# 0.080267f
C252 source.n46 a_n2354_n1088# 0.301973f
C253 source.t33 a_n2354_n1088# 0.137753f
C254 source.n47 a_n2354_n1088# 0.48139f
C255 source.n48 a_n2354_n1088# 0.634306f
C256 drain_right.t10 a_n2354_n1088# 0.020761f
C257 drain_right.t3 a_n2354_n1088# 0.020761f
C258 drain_right.n0 a_n2354_n1088# 0.081316f
C259 drain_right.t12 a_n2354_n1088# 0.020761f
C260 drain_right.t1 a_n2354_n1088# 0.020761f
C261 drain_right.n1 a_n2354_n1088# 0.08067f
C262 drain_right.n2 a_n2354_n1088# 0.561282f
C263 drain_right.t16 a_n2354_n1088# 0.020761f
C264 drain_right.t7 a_n2354_n1088# 0.020761f
C265 drain_right.n3 a_n2354_n1088# 0.08067f
C266 drain_right.n4 a_n2354_n1088# 0.250817f
C267 drain_right.t23 a_n2354_n1088# 0.020761f
C268 drain_right.t15 a_n2354_n1088# 0.020761f
C269 drain_right.n5 a_n2354_n1088# 0.081316f
C270 drain_right.t22 a_n2354_n1088# 0.020761f
C271 drain_right.t21 a_n2354_n1088# 0.020761f
C272 drain_right.n6 a_n2354_n1088# 0.08067f
C273 drain_right.n7 a_n2354_n1088# 0.561282f
C274 drain_right.t13 a_n2354_n1088# 0.020761f
C275 drain_right.t11 a_n2354_n1088# 0.020761f
C276 drain_right.n8 a_n2354_n1088# 0.08067f
C277 drain_right.n9 a_n2354_n1088# 0.250817f
C278 drain_right.n10 a_n2354_n1088# 0.786152f
C279 drain_right.t6 a_n2354_n1088# 0.020761f
C280 drain_right.t17 a_n2354_n1088# 0.020761f
C281 drain_right.n11 a_n2354_n1088# 0.081316f
C282 drain_right.t4 a_n2354_n1088# 0.020761f
C283 drain_right.t20 a_n2354_n1088# 0.020761f
C284 drain_right.n12 a_n2354_n1088# 0.08067f
C285 drain_right.n13 a_n2354_n1088# 0.561282f
C286 drain_right.t2 a_n2354_n1088# 0.020761f
C287 drain_right.t5 a_n2354_n1088# 0.020761f
C288 drain_right.n14 a_n2354_n1088# 0.08067f
C289 drain_right.n15 a_n2354_n1088# 0.275673f
C290 drain_right.t8 a_n2354_n1088# 0.020761f
C291 drain_right.t18 a_n2354_n1088# 0.020761f
C292 drain_right.n16 a_n2354_n1088# 0.08067f
C293 drain_right.n17 a_n2354_n1088# 0.275673f
C294 drain_right.t0 a_n2354_n1088# 0.020761f
C295 drain_right.t19 a_n2354_n1088# 0.020761f
C296 drain_right.n18 a_n2354_n1088# 0.08067f
C297 drain_right.n19 a_n2354_n1088# 0.275673f
C298 drain_right.t9 a_n2354_n1088# 0.020761f
C299 drain_right.t14 a_n2354_n1088# 0.020761f
C300 drain_right.n20 a_n2354_n1088# 0.08067f
C301 drain_right.n21 a_n2354_n1088# 0.49435f
C302 minus.n0 a_n2354_n1088# 0.027971f
C303 minus.t4 a_n2354_n1088# 0.029777f
C304 minus.t19 a_n2354_n1088# 0.025868f
C305 minus.t11 a_n2354_n1088# 0.025868f
C306 minus.n1 a_n2354_n1088# 0.026652f
C307 minus.n2 a_n2354_n1088# 0.027971f
C308 minus.t3 a_n2354_n1088# 0.025868f
C309 minus.t22 a_n2354_n1088# 0.025868f
C310 minus.t10 a_n2354_n1088# 0.025868f
C311 minus.n3 a_n2354_n1088# 0.026652f
C312 minus.n4 a_n2354_n1088# 0.027971f
C313 minus.t1 a_n2354_n1088# 0.025868f
C314 minus.t18 a_n2354_n1088# 0.025868f
C315 minus.n5 a_n2354_n1088# 0.026652f
C316 minus.n6 a_n2354_n1088# 0.027971f
C317 minus.t13 a_n2354_n1088# 0.025868f
C318 minus.t2 a_n2354_n1088# 0.025868f
C319 minus.n7 a_n2354_n1088# 0.010745f
C320 minus.t21 a_n2354_n1088# 0.025868f
C321 minus.n8 a_n2354_n1088# 0.026652f
C322 minus.t15 a_n2354_n1088# 0.029777f
C323 minus.n9 a_n2354_n1088# 0.034559f
C324 minus.n10 a_n2354_n1088# 0.05987f
C325 minus.n11 a_n2354_n1088# 0.027971f
C326 minus.n12 a_n2354_n1088# 0.010055f
C327 minus.n13 a_n2354_n1088# 0.026652f
C328 minus.n14 a_n2354_n1088# 0.011521f
C329 minus.n15 a_n2354_n1088# 0.026652f
C330 minus.n16 a_n2354_n1088# 0.011521f
C331 minus.n17 a_n2354_n1088# 0.027971f
C332 minus.n18 a_n2354_n1088# 0.027971f
C333 minus.n19 a_n2354_n1088# 0.011521f
C334 minus.n20 a_n2354_n1088# 0.026652f
C335 minus.n21 a_n2354_n1088# 0.0104f
C336 minus.n22 a_n2354_n1088# 0.0104f
C337 minus.n23 a_n2354_n1088# 0.027971f
C338 minus.n24 a_n2354_n1088# 0.027971f
C339 minus.n25 a_n2354_n1088# 0.011521f
C340 minus.n26 a_n2354_n1088# 0.026652f
C341 minus.n27 a_n2354_n1088# 0.011521f
C342 minus.n28 a_n2354_n1088# 0.026652f
C343 minus.n29 a_n2354_n1088# 0.011521f
C344 minus.n30 a_n2354_n1088# 0.027971f
C345 minus.n31 a_n2354_n1088# 0.027971f
C346 minus.n32 a_n2354_n1088# 0.010055f
C347 minus.n33 a_n2354_n1088# 0.010745f
C348 minus.n34 a_n2354_n1088# 0.026652f
C349 minus.n35 a_n2354_n1088# 0.034522f
C350 minus.n36 a_n2354_n1088# 0.713394f
C351 minus.n37 a_n2354_n1088# 0.027971f
C352 minus.t0 a_n2354_n1088# 0.025868f
C353 minus.t5 a_n2354_n1088# 0.025868f
C354 minus.n38 a_n2354_n1088# 0.026652f
C355 minus.n39 a_n2354_n1088# 0.027971f
C356 minus.t7 a_n2354_n1088# 0.025868f
C357 minus.t20 a_n2354_n1088# 0.025868f
C358 minus.t23 a_n2354_n1088# 0.025868f
C359 minus.n40 a_n2354_n1088# 0.026652f
C360 minus.n41 a_n2354_n1088# 0.027971f
C361 minus.t9 a_n2354_n1088# 0.025868f
C362 minus.t12 a_n2354_n1088# 0.025868f
C363 minus.n42 a_n2354_n1088# 0.026652f
C364 minus.n43 a_n2354_n1088# 0.027971f
C365 minus.t17 a_n2354_n1088# 0.025868f
C366 minus.t6 a_n2354_n1088# 0.025868f
C367 minus.n44 a_n2354_n1088# 0.010745f
C368 minus.t16 a_n2354_n1088# 0.029777f
C369 minus.t8 a_n2354_n1088# 0.025868f
C370 minus.n45 a_n2354_n1088# 0.026652f
C371 minus.n46 a_n2354_n1088# 0.034559f
C372 minus.n47 a_n2354_n1088# 0.05987f
C373 minus.n48 a_n2354_n1088# 0.027971f
C374 minus.n49 a_n2354_n1088# 0.010055f
C375 minus.n50 a_n2354_n1088# 0.026652f
C376 minus.n51 a_n2354_n1088# 0.011521f
C377 minus.n52 a_n2354_n1088# 0.026652f
C378 minus.n53 a_n2354_n1088# 0.011521f
C379 minus.n54 a_n2354_n1088# 0.027971f
C380 minus.n55 a_n2354_n1088# 0.027971f
C381 minus.n56 a_n2354_n1088# 0.011521f
C382 minus.n57 a_n2354_n1088# 0.026652f
C383 minus.n58 a_n2354_n1088# 0.0104f
C384 minus.n59 a_n2354_n1088# 0.0104f
C385 minus.n60 a_n2354_n1088# 0.027971f
C386 minus.n61 a_n2354_n1088# 0.027971f
C387 minus.n62 a_n2354_n1088# 0.011521f
C388 minus.n63 a_n2354_n1088# 0.026652f
C389 minus.n64 a_n2354_n1088# 0.011521f
C390 minus.n65 a_n2354_n1088# 0.026652f
C391 minus.n66 a_n2354_n1088# 0.011521f
C392 minus.n67 a_n2354_n1088# 0.027971f
C393 minus.n68 a_n2354_n1088# 0.027971f
C394 minus.n69 a_n2354_n1088# 0.010055f
C395 minus.n70 a_n2354_n1088# 0.010745f
C396 minus.n71 a_n2354_n1088# 0.026652f
C397 minus.t14 a_n2354_n1088# 0.029777f
C398 minus.n72 a_n2354_n1088# 0.034522f
C399 minus.n73 a_n2354_n1088# 0.180898f
C400 minus.n74 a_n2354_n1088# 0.881547f
.ends

