* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 drain_left.t13 plus.t0 source.t16 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X2 drain_right.t13 minus.t0 source.t11 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X3 source.t26 plus.t1 drain_left.t12 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X4 source.t14 plus.t2 drain_left.t11 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t4 minus.t1 drain_right.t12 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right.t11 minus.t2 source.t9 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 drain_right.t10 minus.t3 source.t0 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X8 source.t12 minus.t4 drain_right.t9 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_right.t8 minus.t5 source.t1 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X10 source.t5 minus.t6 drain_right.t7 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X11 drain_left.t10 plus.t3 source.t24 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X12 drain_left.t9 plus.t4 source.t22 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X13 drain_left.t8 plus.t5 source.t20 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 source.t17 plus.t6 drain_left.t7 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 source.t8 minus.t7 drain_right.t6 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 drain_right.t5 minus.t8 source.t3 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 source.t15 plus.t7 drain_left.t6 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X18 source.t6 minus.t9 drain_right.t4 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X20 drain_left.t5 plus.t8 source.t18 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X21 drain_right.t3 minus.t10 source.t13 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X22 drain_right.t2 minus.t11 source.t2 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X23 a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X24 source.t25 plus.t9 drain_left.t4 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X25 drain_left.t3 plus.t10 source.t23 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X26 a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X27 drain_right.t1 minus.t12 source.t7 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X28 source.t21 plus.t11 drain_left.t2 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X29 source.t10 minus.t13 drain_right.t0 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X30 drain_left.t1 plus.t12 source.t27 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X31 drain_left.t0 plus.t13 source.t19 a_n2204_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
R0 plus.n5 plus.t10 169.651
R1 plus.n23 plus.t12 169.651
R2 plus.n7 plus.n6 161.3
R3 plus.n8 plus.n3 161.3
R4 plus.n11 plus.n2 161.3
R5 plus.n13 plus.n12 161.3
R6 plus.n14 plus.n1 161.3
R7 plus.n15 plus.n0 161.3
R8 plus.n17 plus.n16 161.3
R9 plus.n25 plus.n24 161.3
R10 plus.n26 plus.n21 161.3
R11 plus.n29 plus.n20 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n19 161.3
R14 plus.n33 plus.n18 161.3
R15 plus.n35 plus.n34 161.3
R16 plus.n16 plus.t0 145.805
R17 plus.n14 plus.t1 145.805
R18 plus.n2 plus.t5 145.805
R19 plus.n9 plus.t7 145.805
R20 plus.n8 plus.t8 145.805
R21 plus.n4 plus.t9 145.805
R22 plus.n34 plus.t4 145.805
R23 plus.n32 plus.t11 145.805
R24 plus.n20 plus.t13 145.805
R25 plus.n27 plus.t2 145.805
R26 plus.n26 plus.t3 145.805
R27 plus.n22 plus.t6 145.805
R28 plus.n10 plus.n9 80.6037
R29 plus.n28 plus.n27 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n14 plus.n13 45.2793
R35 plus.n7 plus.n4 45.2793
R36 plus.n32 plus.n31 45.2793
R37 plus.n25 plus.n22 45.2793
R38 plus.n24 plus.n23 44.9119
R39 plus.n6 plus.n5 44.9119
R40 plus.n16 plus.n15 35.055
R41 plus.n34 plus.n33 35.055
R42 plus plus.n35 27.6373
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n15 plus.n14 13.146
R46 plus.n33 plus.n32 13.146
R47 plus plus.n17 8.43042
R48 plus.n13 plus.n2 2.92171
R49 plus.n8 plus.n7 2.92171
R50 plus.n31 plus.n20 2.92171
R51 plus.n26 plus.n25 2.92171
R52 plus.n10 plus.n3 0.285035
R53 plus.n11 plus.n10 0.285035
R54 plus.n29 plus.n28 0.285035
R55 plus.n28 plus.n21 0.285035
R56 plus.n6 plus.n3 0.189894
R57 plus.n12 plus.n11 0.189894
R58 plus.n12 plus.n1 0.189894
R59 plus.n1 plus.n0 0.189894
R60 plus.n17 plus.n0 0.189894
R61 plus.n35 plus.n18 0.189894
R62 plus.n19 plus.n18 0.189894
R63 plus.n30 plus.n19 0.189894
R64 plus.n30 plus.n29 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n50 source.n48 289.615
R67 source.n36 source.n34 289.615
R68 source.n2 source.n0 289.615
R69 source.n16 source.n14 289.615
R70 source.n51 source.n50 185
R71 source.n37 source.n36 185
R72 source.n3 source.n2 185
R73 source.n17 source.n16 185
R74 source.t7 source.n49 167.117
R75 source.t27 source.n35 167.117
R76 source.t16 source.n1 167.117
R77 source.t13 source.n15 167.117
R78 source.n9 source.n8 84.1169
R79 source.n11 source.n10 84.1169
R80 source.n13 source.n12 84.1169
R81 source.n23 source.n22 84.1169
R82 source.n25 source.n24 84.1169
R83 source.n27 source.n26 84.1169
R84 source.n47 source.n46 84.1168
R85 source.n45 source.n44 84.1168
R86 source.n43 source.n42 84.1168
R87 source.n33 source.n32 84.1168
R88 source.n31 source.n30 84.1168
R89 source.n29 source.n28 84.1168
R90 source.n50 source.t7 52.3082
R91 source.n36 source.t27 52.3082
R92 source.n2 source.t16 52.3082
R93 source.n16 source.t13 52.3082
R94 source.n55 source.n54 31.4096
R95 source.n41 source.n40 31.4096
R96 source.n7 source.n6 31.4096
R97 source.n21 source.n20 31.4096
R98 source.n29 source.n27 15.3154
R99 source.n46 source.t11 9.9005
R100 source.n46 source.t4 9.9005
R101 source.n44 source.t2 9.9005
R102 source.n44 source.t12 9.9005
R103 source.n42 source.t1 9.9005
R104 source.n42 source.t10 9.9005
R105 source.n32 source.t24 9.9005
R106 source.n32 source.t17 9.9005
R107 source.n30 source.t19 9.9005
R108 source.n30 source.t14 9.9005
R109 source.n28 source.t22 9.9005
R110 source.n28 source.t21 9.9005
R111 source.n8 source.t20 9.9005
R112 source.n8 source.t26 9.9005
R113 source.n10 source.t18 9.9005
R114 source.n10 source.t15 9.9005
R115 source.n12 source.t23 9.9005
R116 source.n12 source.t25 9.9005
R117 source.n22 source.t3 9.9005
R118 source.n22 source.t6 9.9005
R119 source.n24 source.t9 9.9005
R120 source.n24 source.t8 9.9005
R121 source.n26 source.t0 9.9005
R122 source.n26 source.t5 9.9005
R123 source.n51 source.n49 9.71174
R124 source.n37 source.n35 9.71174
R125 source.n3 source.n1 9.71174
R126 source.n17 source.n15 9.71174
R127 source.n54 source.n53 9.45567
R128 source.n40 source.n39 9.45567
R129 source.n6 source.n5 9.45567
R130 source.n20 source.n19 9.45567
R131 source.n53 source.n52 9.3005
R132 source.n39 source.n38 9.3005
R133 source.n5 source.n4 9.3005
R134 source.n19 source.n18 9.3005
R135 source.n56 source.n7 8.8499
R136 source.n54 source.n48 8.14595
R137 source.n40 source.n34 8.14595
R138 source.n6 source.n0 8.14595
R139 source.n20 source.n14 8.14595
R140 source.n52 source.n51 7.3702
R141 source.n38 source.n37 7.3702
R142 source.n4 source.n3 7.3702
R143 source.n18 source.n17 7.3702
R144 source.n52 source.n48 5.81868
R145 source.n38 source.n34 5.81868
R146 source.n4 source.n0 5.81868
R147 source.n18 source.n14 5.81868
R148 source.n56 source.n55 5.66429
R149 source.n53 source.n49 3.44771
R150 source.n39 source.n35 3.44771
R151 source.n5 source.n1 3.44771
R152 source.n19 source.n15 3.44771
R153 source.n21 source.n13 0.87119
R154 source.n43 source.n41 0.87119
R155 source.n27 source.n25 0.802224
R156 source.n25 source.n23 0.802224
R157 source.n23 source.n21 0.802224
R158 source.n13 source.n11 0.802224
R159 source.n11 source.n9 0.802224
R160 source.n9 source.n7 0.802224
R161 source.n31 source.n29 0.802224
R162 source.n33 source.n31 0.802224
R163 source.n41 source.n33 0.802224
R164 source.n45 source.n43 0.802224
R165 source.n47 source.n45 0.802224
R166 source.n55 source.n47 0.802224
R167 source source.n56 0.188
R168 drain_left.n2 drain_left.n0 289.615
R169 drain_left.n15 drain_left.n13 289.615
R170 drain_left.n3 drain_left.n2 185
R171 drain_left.n16 drain_left.n15 185
R172 drain_left.t9 drain_left.n1 167.117
R173 drain_left.t3 drain_left.n14 167.117
R174 drain_left.n11 drain_left.n9 101.597
R175 drain_left.n25 drain_left.n24 100.796
R176 drain_left.n23 drain_left.n22 100.796
R177 drain_left.n21 drain_left.n20 100.796
R178 drain_left.n11 drain_left.n10 100.796
R179 drain_left.n8 drain_left.n7 100.796
R180 drain_left.n2 drain_left.t9 52.3082
R181 drain_left.n15 drain_left.t3 52.3082
R182 drain_left.n8 drain_left.n6 48.8901
R183 drain_left.n21 drain_left.n19 48.8901
R184 drain_left drain_left.n12 24.4012
R185 drain_left.n9 drain_left.t7 9.9005
R186 drain_left.n9 drain_left.t1 9.9005
R187 drain_left.n10 drain_left.t11 9.9005
R188 drain_left.n10 drain_left.t10 9.9005
R189 drain_left.n7 drain_left.t2 9.9005
R190 drain_left.n7 drain_left.t0 9.9005
R191 drain_left.n24 drain_left.t12 9.9005
R192 drain_left.n24 drain_left.t13 9.9005
R193 drain_left.n22 drain_left.t6 9.9005
R194 drain_left.n22 drain_left.t8 9.9005
R195 drain_left.n20 drain_left.t4 9.9005
R196 drain_left.n20 drain_left.t5 9.9005
R197 drain_left.n3 drain_left.n1 9.71174
R198 drain_left.n16 drain_left.n14 9.71174
R199 drain_left.n6 drain_left.n5 9.45567
R200 drain_left.n19 drain_left.n18 9.45567
R201 drain_left.n5 drain_left.n4 9.3005
R202 drain_left.n18 drain_left.n17 9.3005
R203 drain_left.n6 drain_left.n0 8.14595
R204 drain_left.n19 drain_left.n13 8.14595
R205 drain_left.n4 drain_left.n3 7.3702
R206 drain_left.n17 drain_left.n16 7.3702
R207 drain_left drain_left.n25 6.45494
R208 drain_left.n4 drain_left.n0 5.81868
R209 drain_left.n17 drain_left.n13 5.81868
R210 drain_left.n5 drain_left.n1 3.44771
R211 drain_left.n18 drain_left.n14 3.44771
R212 drain_left.n23 drain_left.n21 0.802224
R213 drain_left.n25 drain_left.n23 0.802224
R214 drain_left.n12 drain_left.n8 0.546447
R215 drain_left.n12 drain_left.n11 0.145585
R216 minus.n5 minus.t10 169.651
R217 minus.n23 minus.t5 169.651
R218 minus.n17 minus.n16 161.3
R219 minus.n15 minus.n0 161.3
R220 minus.n14 minus.n13 161.3
R221 minus.n12 minus.n1 161.3
R222 minus.n11 minus.n10 161.3
R223 minus.n8 minus.n7 161.3
R224 minus.n6 minus.n3 161.3
R225 minus.n35 minus.n34 161.3
R226 minus.n33 minus.n18 161.3
R227 minus.n32 minus.n31 161.3
R228 minus.n30 minus.n19 161.3
R229 minus.n29 minus.n28 161.3
R230 minus.n26 minus.n25 161.3
R231 minus.n24 minus.n21 161.3
R232 minus.n4 minus.t9 145.805
R233 minus.n8 minus.t8 145.805
R234 minus.n9 minus.t7 145.805
R235 minus.n10 minus.t2 145.805
R236 minus.n14 minus.t6 145.805
R237 minus.n16 minus.t3 145.805
R238 minus.n22 minus.t13 145.805
R239 minus.n26 minus.t11 145.805
R240 minus.n27 minus.t4 145.805
R241 minus.n28 minus.t0 145.805
R242 minus.n32 minus.t1 145.805
R243 minus.n34 minus.t12 145.805
R244 minus.n9 minus.n2 80.6037
R245 minus.n27 minus.n20 80.6037
R246 minus.n9 minus.n8 48.2005
R247 minus.n10 minus.n9 48.2005
R248 minus.n27 minus.n26 48.2005
R249 minus.n28 minus.n27 48.2005
R250 minus.n4 minus.n3 45.2793
R251 minus.n14 minus.n1 45.2793
R252 minus.n22 minus.n21 45.2793
R253 minus.n32 minus.n19 45.2793
R254 minus.n6 minus.n5 44.9119
R255 minus.n24 minus.n23 44.9119
R256 minus.n16 minus.n15 35.055
R257 minus.n34 minus.n33 35.055
R258 minus.n36 minus.n17 29.9683
R259 minus.n5 minus.n4 17.739
R260 minus.n23 minus.n22 17.739
R261 minus.n15 minus.n14 13.146
R262 minus.n33 minus.n32 13.146
R263 minus.n36 minus.n35 6.57436
R264 minus.n8 minus.n3 2.92171
R265 minus.n10 minus.n1 2.92171
R266 minus.n26 minus.n21 2.92171
R267 minus.n28 minus.n19 2.92171
R268 minus.n11 minus.n2 0.285035
R269 minus.n7 minus.n2 0.285035
R270 minus.n25 minus.n20 0.285035
R271 minus.n29 minus.n20 0.285035
R272 minus.n17 minus.n0 0.189894
R273 minus.n13 minus.n0 0.189894
R274 minus.n13 minus.n12 0.189894
R275 minus.n12 minus.n11 0.189894
R276 minus.n7 minus.n6 0.189894
R277 minus.n25 minus.n24 0.189894
R278 minus.n30 minus.n29 0.189894
R279 minus.n31 minus.n30 0.189894
R280 minus.n31 minus.n18 0.189894
R281 minus.n35 minus.n18 0.189894
R282 minus minus.n36 0.188
R283 drain_right.n2 drain_right.n0 289.615
R284 drain_right.n20 drain_right.n18 289.615
R285 drain_right.n3 drain_right.n2 185
R286 drain_right.n21 drain_right.n20 185
R287 drain_right.t8 drain_right.n1 167.117
R288 drain_right.t10 drain_right.n19 167.117
R289 drain_right.n15 drain_right.n13 101.597
R290 drain_right.n11 drain_right.n9 101.597
R291 drain_right.n15 drain_right.n14 100.796
R292 drain_right.n17 drain_right.n16 100.796
R293 drain_right.n11 drain_right.n10 100.796
R294 drain_right.n8 drain_right.n7 100.796
R295 drain_right.n2 drain_right.t8 52.3082
R296 drain_right.n20 drain_right.t10 52.3082
R297 drain_right.n8 drain_right.n6 48.8901
R298 drain_right.n25 drain_right.n24 48.0884
R299 drain_right drain_right.n12 23.848
R300 drain_right.n9 drain_right.t12 9.9005
R301 drain_right.n9 drain_right.t1 9.9005
R302 drain_right.n10 drain_right.t9 9.9005
R303 drain_right.n10 drain_right.t13 9.9005
R304 drain_right.n7 drain_right.t0 9.9005
R305 drain_right.n7 drain_right.t2 9.9005
R306 drain_right.n13 drain_right.t4 9.9005
R307 drain_right.n13 drain_right.t3 9.9005
R308 drain_right.n14 drain_right.t6 9.9005
R309 drain_right.n14 drain_right.t5 9.9005
R310 drain_right.n16 drain_right.t7 9.9005
R311 drain_right.n16 drain_right.t11 9.9005
R312 drain_right.n3 drain_right.n1 9.71174
R313 drain_right.n21 drain_right.n19 9.71174
R314 drain_right.n6 drain_right.n5 9.45567
R315 drain_right.n24 drain_right.n23 9.45567
R316 drain_right.n5 drain_right.n4 9.3005
R317 drain_right.n23 drain_right.n22 9.3005
R318 drain_right.n6 drain_right.n0 8.14595
R319 drain_right.n24 drain_right.n18 8.14595
R320 drain_right.n4 drain_right.n3 7.3702
R321 drain_right.n22 drain_right.n21 7.3702
R322 drain_right drain_right.n25 6.05408
R323 drain_right.n4 drain_right.n0 5.81868
R324 drain_right.n22 drain_right.n18 5.81868
R325 drain_right.n5 drain_right.n1 3.44771
R326 drain_right.n23 drain_right.n19 3.44771
R327 drain_right.n25 drain_right.n17 0.802224
R328 drain_right.n17 drain_right.n15 0.802224
R329 drain_right.n12 drain_right.n8 0.546447
R330 drain_right.n12 drain_right.n11 0.145585
C0 minus drain_right 1.81704f
C1 minus plus 4.05421f
C2 source drain_right 5.89283f
C3 source plus 2.26507f
C4 minus drain_left 0.179263f
C5 source drain_left 5.89342f
C6 drain_right plus 0.380191f
C7 minus source 2.25102f
C8 drain_right drain_left 1.14494f
C9 drain_left plus 2.03303f
C10 drain_right a_n2204_n1288# 4.20701f
C11 drain_left a_n2204_n1288# 4.895741f
C12 source a_n2204_n1288# 2.732844f
C13 minus a_n2204_n1288# 7.902396f
C14 plus a_n2204_n1288# 9.17912f
C15 drain_right.n0 a_n2204_n1288# 0.028671f
C16 drain_right.n1 a_n2204_n1288# 0.063437f
C17 drain_right.t8 a_n2204_n1288# 0.047606f
C18 drain_right.n2 a_n2204_n1288# 0.049648f
C19 drain_right.n3 a_n2204_n1288# 0.016005f
C20 drain_right.n4 a_n2204_n1288# 0.010556f
C21 drain_right.n5 a_n2204_n1288# 0.139831f
C22 drain_right.n6 a_n2204_n1288# 0.046444f
C23 drain_right.t0 a_n2204_n1288# 0.031046f
C24 drain_right.t2 a_n2204_n1288# 0.031046f
C25 drain_right.n7 a_n2204_n1288# 0.195037f
C26 drain_right.n8 a_n2204_n1288# 0.322996f
C27 drain_right.t12 a_n2204_n1288# 0.031046f
C28 drain_right.t1 a_n2204_n1288# 0.031046f
C29 drain_right.n9 a_n2204_n1288# 0.197087f
C30 drain_right.t9 a_n2204_n1288# 0.031046f
C31 drain_right.t13 a_n2204_n1288# 0.031046f
C32 drain_right.n10 a_n2204_n1288# 0.195037f
C33 drain_right.n11 a_n2204_n1288# 0.471116f
C34 drain_right.n12 a_n2204_n1288# 0.604154f
C35 drain_right.t4 a_n2204_n1288# 0.031046f
C36 drain_right.t3 a_n2204_n1288# 0.031046f
C37 drain_right.n13 a_n2204_n1288# 0.197088f
C38 drain_right.t6 a_n2204_n1288# 0.031046f
C39 drain_right.t5 a_n2204_n1288# 0.031046f
C40 drain_right.n14 a_n2204_n1288# 0.195038f
C41 drain_right.n15 a_n2204_n1288# 0.509538f
C42 drain_right.t7 a_n2204_n1288# 0.031046f
C43 drain_right.t11 a_n2204_n1288# 0.031046f
C44 drain_right.n16 a_n2204_n1288# 0.195038f
C45 drain_right.n17 a_n2204_n1288# 0.251838f
C46 drain_right.n18 a_n2204_n1288# 0.028671f
C47 drain_right.n19 a_n2204_n1288# 0.063437f
C48 drain_right.t10 a_n2204_n1288# 0.047606f
C49 drain_right.n20 a_n2204_n1288# 0.049648f
C50 drain_right.n21 a_n2204_n1288# 0.016005f
C51 drain_right.n22 a_n2204_n1288# 0.010556f
C52 drain_right.n23 a_n2204_n1288# 0.139831f
C53 drain_right.n24 a_n2204_n1288# 0.045002f
C54 drain_right.n25 a_n2204_n1288# 0.264354f
C55 minus.n0 a_n2204_n1288# 0.035795f
C56 minus.n1 a_n2204_n1288# 0.008123f
C57 minus.t6 a_n2204_n1288# 0.133016f
C58 minus.n2 a_n2204_n1288# 0.047652f
C59 minus.n3 a_n2204_n1288# 0.008123f
C60 minus.t8 a_n2204_n1288# 0.133016f
C61 minus.t10 a_n2204_n1288# 0.146167f
C62 minus.t9 a_n2204_n1288# 0.133016f
C63 minus.n4 a_n2204_n1288# 0.10017f
C64 minus.n5 a_n2204_n1288# 0.083454f
C65 minus.n6 a_n2204_n1288# 0.14644f
C66 minus.n7 a_n2204_n1288# 0.047764f
C67 minus.n8 a_n2204_n1288# 0.094633f
C68 minus.t7 a_n2204_n1288# 0.133016f
C69 minus.n9 a_n2204_n1288# 0.102314f
C70 minus.t2 a_n2204_n1288# 0.133016f
C71 minus.n10 a_n2204_n1288# 0.094633f
C72 minus.n11 a_n2204_n1288# 0.047764f
C73 minus.n12 a_n2204_n1288# 0.035795f
C74 minus.n13 a_n2204_n1288# 0.035795f
C75 minus.n14 a_n2204_n1288# 0.095737f
C76 minus.n15 a_n2204_n1288# 0.008123f
C77 minus.t3 a_n2204_n1288# 0.133016f
C78 minus.n16 a_n2204_n1288# 0.092206f
C79 minus.n17 a_n2204_n1288# 0.931973f
C80 minus.n18 a_n2204_n1288# 0.035795f
C81 minus.n19 a_n2204_n1288# 0.008123f
C82 minus.n20 a_n2204_n1288# 0.047652f
C83 minus.n21 a_n2204_n1288# 0.008123f
C84 minus.t5 a_n2204_n1288# 0.146167f
C85 minus.t13 a_n2204_n1288# 0.133016f
C86 minus.n22 a_n2204_n1288# 0.10017f
C87 minus.n23 a_n2204_n1288# 0.083454f
C88 minus.n24 a_n2204_n1288# 0.14644f
C89 minus.n25 a_n2204_n1288# 0.047764f
C90 minus.t11 a_n2204_n1288# 0.133016f
C91 minus.n26 a_n2204_n1288# 0.094633f
C92 minus.t4 a_n2204_n1288# 0.133016f
C93 minus.n27 a_n2204_n1288# 0.102314f
C94 minus.t0 a_n2204_n1288# 0.133016f
C95 minus.n28 a_n2204_n1288# 0.094633f
C96 minus.n29 a_n2204_n1288# 0.047764f
C97 minus.n30 a_n2204_n1288# 0.035795f
C98 minus.n31 a_n2204_n1288# 0.035795f
C99 minus.t1 a_n2204_n1288# 0.133016f
C100 minus.n32 a_n2204_n1288# 0.095737f
C101 minus.n33 a_n2204_n1288# 0.008123f
C102 minus.t12 a_n2204_n1288# 0.133016f
C103 minus.n34 a_n2204_n1288# 0.092206f
C104 minus.n35 a_n2204_n1288# 0.240266f
C105 minus.n36 a_n2204_n1288# 1.14669f
C106 drain_left.n0 a_n2204_n1288# 0.037896f
C107 drain_left.n1 a_n2204_n1288# 0.083849f
C108 drain_left.t9 a_n2204_n1288# 0.062925f
C109 drain_left.n2 a_n2204_n1288# 0.065624f
C110 drain_left.n3 a_n2204_n1288# 0.021155f
C111 drain_left.n4 a_n2204_n1288# 0.013952f
C112 drain_left.n5 a_n2204_n1288# 0.184825f
C113 drain_left.n6 a_n2204_n1288# 0.061388f
C114 drain_left.t2 a_n2204_n1288# 0.041035f
C115 drain_left.t0 a_n2204_n1288# 0.041035f
C116 drain_left.n7 a_n2204_n1288# 0.257794f
C117 drain_left.n8 a_n2204_n1288# 0.426926f
C118 drain_left.t7 a_n2204_n1288# 0.041035f
C119 drain_left.t1 a_n2204_n1288# 0.041035f
C120 drain_left.n9 a_n2204_n1288# 0.260503f
C121 drain_left.t11 a_n2204_n1288# 0.041035f
C122 drain_left.t10 a_n2204_n1288# 0.041035f
C123 drain_left.n10 a_n2204_n1288# 0.257794f
C124 drain_left.n11 a_n2204_n1288# 0.622706f
C125 drain_left.n12 a_n2204_n1288# 0.849242f
C126 drain_left.n13 a_n2204_n1288# 0.037896f
C127 drain_left.n14 a_n2204_n1288# 0.083849f
C128 drain_left.t3 a_n2204_n1288# 0.062925f
C129 drain_left.n15 a_n2204_n1288# 0.065624f
C130 drain_left.n16 a_n2204_n1288# 0.021155f
C131 drain_left.n17 a_n2204_n1288# 0.013952f
C132 drain_left.n18 a_n2204_n1288# 0.184825f
C133 drain_left.n19 a_n2204_n1288# 0.061388f
C134 drain_left.t4 a_n2204_n1288# 0.041035f
C135 drain_left.t5 a_n2204_n1288# 0.041035f
C136 drain_left.n20 a_n2204_n1288# 0.257795f
C137 drain_left.n21 a_n2204_n1288# 0.447221f
C138 drain_left.t6 a_n2204_n1288# 0.041035f
C139 drain_left.t8 a_n2204_n1288# 0.041035f
C140 drain_left.n22 a_n2204_n1288# 0.257795f
C141 drain_left.n23 a_n2204_n1288# 0.332871f
C142 drain_left.t12 a_n2204_n1288# 0.041035f
C143 drain_left.t13 a_n2204_n1288# 0.041035f
C144 drain_left.n24 a_n2204_n1288# 0.257795f
C145 drain_left.n25 a_n2204_n1288# 0.559274f
C146 source.n0 a_n2204_n1288# 0.049226f
C147 source.n1 a_n2204_n1288# 0.108919f
C148 source.t16 a_n2204_n1288# 0.081738f
C149 source.n2 a_n2204_n1288# 0.085245f
C150 source.n3 a_n2204_n1288# 0.02748f
C151 source.n4 a_n2204_n1288# 0.018123f
C152 source.n5 a_n2204_n1288# 0.240085f
C153 source.n6 a_n2204_n1288# 0.053964f
C154 source.n7 a_n2204_n1288# 0.559053f
C155 source.t20 a_n2204_n1288# 0.053304f
C156 source.t26 a_n2204_n1288# 0.053304f
C157 source.n8 a_n2204_n1288# 0.284961f
C158 source.n9 a_n2204_n1288# 0.436466f
C159 source.t18 a_n2204_n1288# 0.053304f
C160 source.t15 a_n2204_n1288# 0.053304f
C161 source.n10 a_n2204_n1288# 0.284961f
C162 source.n11 a_n2204_n1288# 0.436466f
C163 source.t23 a_n2204_n1288# 0.053304f
C164 source.t25 a_n2204_n1288# 0.053304f
C165 source.n12 a_n2204_n1288# 0.284961f
C166 source.n13 a_n2204_n1288# 0.44396f
C167 source.n14 a_n2204_n1288# 0.049226f
C168 source.n15 a_n2204_n1288# 0.108919f
C169 source.t13 a_n2204_n1288# 0.081738f
C170 source.n16 a_n2204_n1288# 0.085245f
C171 source.n17 a_n2204_n1288# 0.02748f
C172 source.n18 a_n2204_n1288# 0.018123f
C173 source.n19 a_n2204_n1288# 0.240085f
C174 source.n20 a_n2204_n1288# 0.053964f
C175 source.n21 a_n2204_n1288# 0.209515f
C176 source.t3 a_n2204_n1288# 0.053304f
C177 source.t6 a_n2204_n1288# 0.053304f
C178 source.n22 a_n2204_n1288# 0.284961f
C179 source.n23 a_n2204_n1288# 0.436466f
C180 source.t9 a_n2204_n1288# 0.053304f
C181 source.t8 a_n2204_n1288# 0.053304f
C182 source.n24 a_n2204_n1288# 0.284961f
C183 source.n25 a_n2204_n1288# 0.436466f
C184 source.t0 a_n2204_n1288# 0.053304f
C185 source.t5 a_n2204_n1288# 0.053304f
C186 source.n26 a_n2204_n1288# 0.284961f
C187 source.n27 a_n2204_n1288# 1.20144f
C188 source.t22 a_n2204_n1288# 0.053304f
C189 source.t21 a_n2204_n1288# 0.053304f
C190 source.n28 a_n2204_n1288# 0.284959f
C191 source.n29 a_n2204_n1288# 1.20144f
C192 source.t19 a_n2204_n1288# 0.053304f
C193 source.t14 a_n2204_n1288# 0.053304f
C194 source.n30 a_n2204_n1288# 0.284959f
C195 source.n31 a_n2204_n1288# 0.436467f
C196 source.t24 a_n2204_n1288# 0.053304f
C197 source.t17 a_n2204_n1288# 0.053304f
C198 source.n32 a_n2204_n1288# 0.284959f
C199 source.n33 a_n2204_n1288# 0.436467f
C200 source.n34 a_n2204_n1288# 0.049226f
C201 source.n35 a_n2204_n1288# 0.108919f
C202 source.t27 a_n2204_n1288# 0.081738f
C203 source.n36 a_n2204_n1288# 0.085245f
C204 source.n37 a_n2204_n1288# 0.02748f
C205 source.n38 a_n2204_n1288# 0.018123f
C206 source.n39 a_n2204_n1288# 0.240085f
C207 source.n40 a_n2204_n1288# 0.053964f
C208 source.n41 a_n2204_n1288# 0.209515f
C209 source.t1 a_n2204_n1288# 0.053304f
C210 source.t10 a_n2204_n1288# 0.053304f
C211 source.n42 a_n2204_n1288# 0.284959f
C212 source.n43 a_n2204_n1288# 0.443962f
C213 source.t2 a_n2204_n1288# 0.053304f
C214 source.t12 a_n2204_n1288# 0.053304f
C215 source.n44 a_n2204_n1288# 0.284959f
C216 source.n45 a_n2204_n1288# 0.436467f
C217 source.t11 a_n2204_n1288# 0.053304f
C218 source.t4 a_n2204_n1288# 0.053304f
C219 source.n46 a_n2204_n1288# 0.284959f
C220 source.n47 a_n2204_n1288# 0.436467f
C221 source.n48 a_n2204_n1288# 0.049226f
C222 source.n49 a_n2204_n1288# 0.108919f
C223 source.t7 a_n2204_n1288# 0.081738f
C224 source.n50 a_n2204_n1288# 0.085245f
C225 source.n51 a_n2204_n1288# 0.02748f
C226 source.n52 a_n2204_n1288# 0.018123f
C227 source.n53 a_n2204_n1288# 0.240085f
C228 source.n54 a_n2204_n1288# 0.053964f
C229 source.n55 a_n2204_n1288# 0.378611f
C230 source.n56 a_n2204_n1288# 0.846059f
C231 plus.n0 a_n2204_n1288# 0.047518f
C232 plus.t0 a_n2204_n1288# 0.176581f
C233 plus.t1 a_n2204_n1288# 0.176581f
C234 plus.n1 a_n2204_n1288# 0.047518f
C235 plus.t5 a_n2204_n1288# 0.176581f
C236 plus.n2 a_n2204_n1288# 0.125627f
C237 plus.n3 a_n2204_n1288# 0.063407f
C238 plus.t7 a_n2204_n1288# 0.176581f
C239 plus.t8 a_n2204_n1288# 0.176581f
C240 plus.t9 a_n2204_n1288# 0.176581f
C241 plus.n4 a_n2204_n1288# 0.132978f
C242 plus.t10 a_n2204_n1288# 0.194039f
C243 plus.n5 a_n2204_n1288# 0.110787f
C244 plus.n6 a_n2204_n1288# 0.194402f
C245 plus.n7 a_n2204_n1288# 0.010783f
C246 plus.n8 a_n2204_n1288# 0.125627f
C247 plus.n9 a_n2204_n1288# 0.135824f
C248 plus.n10 a_n2204_n1288# 0.063258f
C249 plus.n11 a_n2204_n1288# 0.063407f
C250 plus.n12 a_n2204_n1288# 0.047518f
C251 plus.n13 a_n2204_n1288# 0.010783f
C252 plus.n14 a_n2204_n1288# 0.127092f
C253 plus.n15 a_n2204_n1288# 0.010783f
C254 plus.n16 a_n2204_n1288# 0.122404f
C255 plus.n17 a_n2204_n1288# 0.348448f
C256 plus.n18 a_n2204_n1288# 0.047518f
C257 plus.t4 a_n2204_n1288# 0.176581f
C258 plus.n19 a_n2204_n1288# 0.047518f
C259 plus.t11 a_n2204_n1288# 0.176581f
C260 plus.t13 a_n2204_n1288# 0.176581f
C261 plus.n20 a_n2204_n1288# 0.125627f
C262 plus.n21 a_n2204_n1288# 0.063407f
C263 plus.t2 a_n2204_n1288# 0.176581f
C264 plus.t3 a_n2204_n1288# 0.176581f
C265 plus.t6 a_n2204_n1288# 0.176581f
C266 plus.n22 a_n2204_n1288# 0.132978f
C267 plus.t12 a_n2204_n1288# 0.194039f
C268 plus.n23 a_n2204_n1288# 0.110787f
C269 plus.n24 a_n2204_n1288# 0.194402f
C270 plus.n25 a_n2204_n1288# 0.010783f
C271 plus.n26 a_n2204_n1288# 0.125627f
C272 plus.n27 a_n2204_n1288# 0.135824f
C273 plus.n28 a_n2204_n1288# 0.063258f
C274 plus.n29 a_n2204_n1288# 0.063407f
C275 plus.n30 a_n2204_n1288# 0.047518f
C276 plus.n31 a_n2204_n1288# 0.010783f
C277 plus.n32 a_n2204_n1288# 0.127092f
C278 plus.n33 a_n2204_n1288# 0.010783f
C279 plus.n34 a_n2204_n1288# 0.122404f
C280 plus.n35 a_n2204_n1288# 1.1786f
.ends

