* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X1 drain_left.t13 plus.t0 source.t26 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X2 source.t11 minus.t0 drain_right.t13 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 drain_right.t12 minus.t1 source.t12 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 drain_right.t11 minus.t2 source.t13 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X5 source.t21 plus.t1 drain_left.t12 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X6 source.t22 plus.t2 drain_left.t11 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X7 drain_left.t10 plus.t3 source.t23 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X8 source.t3 minus.t3 drain_right.t10 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X9 source.t8 minus.t4 drain_right.t9 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X10 drain_left.t9 plus.t4 source.t25 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X11 drain_right.t8 minus.t5 source.t7 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X12 a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X13 drain_right.t7 minus.t6 source.t10 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 drain_left.t8 plus.t5 source.t27 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X15 source.t24 plus.t6 drain_left.t7 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X16 drain_left.t6 plus.t7 source.t14 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X17 source.t1 minus.t7 drain_right.t6 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X18 drain_right.t5 minus.t8 source.t4 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X19 drain_right.t4 minus.t9 source.t0 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X20 source.t15 plus.t8 drain_left.t5 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X21 source.t16 plus.t9 drain_left.t4 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X22 drain_left.t3 plus.t10 source.t19 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 source.t2 minus.t10 drain_right.t3 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X24 drain_left.t2 plus.t11 source.t17 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X25 a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X26 drain_right.t2 minus.t11 source.t5 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X27 a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X28 source.t6 minus.t12 drain_right.t1 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X29 drain_right.t0 minus.t13 source.t9 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X30 drain_left.t1 plus.t12 source.t18 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X31 source.t20 plus.t13 drain_left.t0 a_n1724_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
R0 plus.n3 plus.t3 241.731
R1 plus.n15 plus.t12 241.731
R2 plus.n20 plus.t7 241.731
R3 plus.n32 plus.t11 241.731
R4 plus.n1 plus.t13 184.768
R5 plus.n4 plus.t6 184.768
R6 plus.n6 plus.t10 184.768
R7 plus.n12 plus.t5 184.768
R8 plus.n14 plus.t8 184.768
R9 plus.n18 plus.t9 184.768
R10 plus.n21 plus.t1 184.768
R11 plus.n23 plus.t0 184.768
R12 plus.n29 plus.t4 184.768
R13 plus.n31 plus.t2 184.768
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 54.0429
R33 plus.n13 plus.n12 54.0429
R34 plus.n30 plus.n29 54.0429
R35 plus.n23 plus.n22 54.0429
R36 plus.n5 plus.n4 37.9763
R37 plus.n14 plus.n13 37.9763
R38 plus.n31 plus.n30 37.9763
R39 plus.n22 plus.n21 37.9763
R40 plus.n4 plus.n3 35.055
R41 plus.n15 plus.n14 35.055
R42 plus.n32 plus.n31 35.055
R43 plus.n21 plus.n20 35.055
R44 plus plus.n33 25.4024
R45 plus.n7 plus.n6 18.9884
R46 plus.n12 plus.n11 18.9884
R47 plus.n29 plus.n28 18.9884
R48 plus.n24 plus.n23 18.9884
R49 plus plus.n16 8.01376
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 source.n0 source.t18 243.255
R61 source.n7 source.t4 243.255
R62 source.n27 source.t9 243.254
R63 source.n20 source.t14 243.254
R64 source.n2 source.n1 223.454
R65 source.n4 source.n3 223.454
R66 source.n6 source.n5 223.454
R67 source.n9 source.n8 223.454
R68 source.n11 source.n10 223.454
R69 source.n13 source.n12 223.454
R70 source.n26 source.n25 223.453
R71 source.n24 source.n23 223.453
R72 source.n22 source.n21 223.453
R73 source.n19 source.n18 223.453
R74 source.n17 source.n16 223.453
R75 source.n15 source.n14 223.453
R76 source.n25 source.t10 19.8005
R77 source.n25 source.t8 19.8005
R78 source.n23 source.t13 19.8005
R79 source.n23 source.t2 19.8005
R80 source.n21 source.t0 19.8005
R81 source.n21 source.t3 19.8005
R82 source.n18 source.t26 19.8005
R83 source.n18 source.t21 19.8005
R84 source.n16 source.t25 19.8005
R85 source.n16 source.t16 19.8005
R86 source.n14 source.t17 19.8005
R87 source.n14 source.t22 19.8005
R88 source.n1 source.t27 19.8005
R89 source.n1 source.t15 19.8005
R90 source.n3 source.t19 19.8005
R91 source.n3 source.t20 19.8005
R92 source.n5 source.t23 19.8005
R93 source.n5 source.t24 19.8005
R94 source.n8 source.t12 19.8005
R95 source.n8 source.t6 19.8005
R96 source.n10 source.t5 19.8005
R97 source.n10 source.t1 19.8005
R98 source.n12 source.t7 19.8005
R99 source.n12 source.t11 19.8005
R100 source.n15 source.n13 14.0406
R101 source.n28 source.n0 7.96301
R102 source.n28 source.n27 5.53498
R103 source.n7 source.n6 0.741879
R104 source.n22 source.n20 0.741879
R105 source.n13 source.n11 0.543603
R106 source.n11 source.n9 0.543603
R107 source.n9 source.n7 0.543603
R108 source.n6 source.n4 0.543603
R109 source.n4 source.n2 0.543603
R110 source.n2 source.n0 0.543603
R111 source.n17 source.n15 0.543603
R112 source.n19 source.n17 0.543603
R113 source.n20 source.n19 0.543603
R114 source.n24 source.n22 0.543603
R115 source.n26 source.n24 0.543603
R116 source.n27 source.n26 0.543603
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t10 260.476
R119 drain_left.n1 drain_left.t2 260.474
R120 drain_left.n4 drain_left.n2 240.674
R121 drain_left.n11 drain_left.n10 240.132
R122 drain_left.n9 drain_left.n8 240.132
R123 drain_left.n7 drain_left.n6 240.132
R124 drain_left.n4 drain_left.n3 240.131
R125 drain_left.n1 drain_left.n0 240.131
R126 drain_left drain_left.n5 22.1566
R127 drain_left.n2 drain_left.t12 19.8005
R128 drain_left.n2 drain_left.t6 19.8005
R129 drain_left.n3 drain_left.t4 19.8005
R130 drain_left.n3 drain_left.t13 19.8005
R131 drain_left.n0 drain_left.t11 19.8005
R132 drain_left.n0 drain_left.t9 19.8005
R133 drain_left.n10 drain_left.t5 19.8005
R134 drain_left.n10 drain_left.t1 19.8005
R135 drain_left.n8 drain_left.t0 19.8005
R136 drain_left.n8 drain_left.t8 19.8005
R137 drain_left.n6 drain_left.t7 19.8005
R138 drain_left.n6 drain_left.t3 19.8005
R139 drain_left drain_left.n11 6.19632
R140 drain_left.n9 drain_left.n7 0.543603
R141 drain_left.n11 drain_left.n9 0.543603
R142 drain_left.n5 drain_left.n1 0.352482
R143 drain_left.n5 drain_left.n4 0.0809298
R144 minus.n15 minus.t5 241.731
R145 minus.n3 minus.t8 241.731
R146 minus.n32 minus.t13 241.731
R147 minus.n20 minus.t9 241.731
R148 minus.n1 minus.t7 184.768
R149 minus.n14 minus.t0 184.768
R150 minus.n12 minus.t11 184.768
R151 minus.n6 minus.t1 184.768
R152 minus.n4 minus.t12 184.768
R153 minus.n18 minus.t10 184.768
R154 minus.n31 minus.t4 184.768
R155 minus.n29 minus.t6 184.768
R156 minus.n23 minus.t2 184.768
R157 minus.n21 minus.t3 184.768
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 54.0429
R177 minus.n6 minus.n5 54.0429
R178 minus.n23 minus.n22 54.0429
R179 minus.n30 minus.n29 54.0429
R180 minus.n14 minus.n13 37.9763
R181 minus.n5 minus.n4 37.9763
R182 minus.n22 minus.n21 37.9763
R183 minus.n31 minus.n30 37.9763
R184 minus.n15 minus.n14 35.055
R185 minus.n4 minus.n3 35.055
R186 minus.n21 minus.n20 35.055
R187 minus.n32 minus.n31 35.055
R188 minus.n34 minus.n16 27.3547
R189 minus.n12 minus.n11 18.9884
R190 minus.n7 minus.n6 18.9884
R191 minus.n24 minus.n23 18.9884
R192 minus.n29 minus.n28 18.9884
R193 minus.n34 minus.n33 6.53648
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t4 260.474
R206 drain_right.n11 drain_right.t8 259.933
R207 drain_right.n8 drain_right.n6 240.675
R208 drain_right.n4 drain_right.n2 240.674
R209 drain_right.n8 drain_right.n7 240.132
R210 drain_right.n10 drain_right.n9 240.132
R211 drain_right.n4 drain_right.n3 240.131
R212 drain_right.n1 drain_right.n0 240.131
R213 drain_right drain_right.n5 21.6034
R214 drain_right.n2 drain_right.t9 19.8005
R215 drain_right.n2 drain_right.t0 19.8005
R216 drain_right.n3 drain_right.t3 19.8005
R217 drain_right.n3 drain_right.t7 19.8005
R218 drain_right.n0 drain_right.t10 19.8005
R219 drain_right.n0 drain_right.t11 19.8005
R220 drain_right.n6 drain_right.t1 19.8005
R221 drain_right.n6 drain_right.t5 19.8005
R222 drain_right.n7 drain_right.t6 19.8005
R223 drain_right.n7 drain_right.t12 19.8005
R224 drain_right.n9 drain_right.t13 19.8005
R225 drain_right.n9 drain_right.t2 19.8005
R226 drain_right drain_right.n11 5.92477
R227 drain_right.n11 drain_right.n10 0.543603
R228 drain_right.n10 drain_right.n8 0.543603
R229 drain_right.n5 drain_right.n1 0.352482
R230 drain_right.n5 drain_right.n4 0.0809298
C0 plus source 1.16338f
C1 source drain_left 4.75612f
C2 drain_right minus 0.874137f
C3 drain_right plus 0.330384f
C4 plus minus 3.27164f
C5 drain_right drain_left 0.879354f
C6 drain_right source 4.75452f
C7 minus drain_left 0.179577f
C8 plus drain_left 1.04049f
C9 minus source 1.14946f
C10 drain_right a_n1724_n1088# 3.60545f
C11 drain_left a_n1724_n1088# 3.84596f
C12 source a_n1724_n1088# 2.150157f
C13 minus a_n1724_n1088# 5.80237f
C14 plus a_n1724_n1088# 6.482839f
C15 drain_right.t4 a_n1724_n1088# 0.118971f
C16 drain_right.t10 a_n1724_n1088# 0.019157f
C17 drain_right.t11 a_n1724_n1088# 0.019157f
C18 drain_right.n0 a_n1724_n1088# 0.074437f
C19 drain_right.n1 a_n1724_n1088# 0.470463f
C20 drain_right.t9 a_n1724_n1088# 0.019157f
C21 drain_right.t0 a_n1724_n1088# 0.019157f
C22 drain_right.n2 a_n1724_n1088# 0.075033f
C23 drain_right.t3 a_n1724_n1088# 0.019157f
C24 drain_right.t7 a_n1724_n1088# 0.019157f
C25 drain_right.n3 a_n1724_n1088# 0.074437f
C26 drain_right.n4 a_n1724_n1088# 0.488758f
C27 drain_right.n5 a_n1724_n1088# 0.573195f
C28 drain_right.t1 a_n1724_n1088# 0.019157f
C29 drain_right.t5 a_n1724_n1088# 0.019157f
C30 drain_right.n6 a_n1724_n1088# 0.075033f
C31 drain_right.t6 a_n1724_n1088# 0.019157f
C32 drain_right.t12 a_n1724_n1088# 0.019157f
C33 drain_right.n7 a_n1724_n1088# 0.074437f
C34 drain_right.n8 a_n1724_n1088# 0.517911f
C35 drain_right.t13 a_n1724_n1088# 0.019157f
C36 drain_right.t2 a_n1724_n1088# 0.019157f
C37 drain_right.n9 a_n1724_n1088# 0.074437f
C38 drain_right.n10 a_n1724_n1088# 0.254371f
C39 drain_right.t8 a_n1724_n1088# 0.118491f
C40 drain_right.n11 a_n1724_n1088# 0.432139f
C41 minus.n0 a_n1724_n1088# 0.032389f
C42 minus.t5 a_n1724_n1088# 0.038121f
C43 minus.t0 a_n1724_n1088# 0.029954f
C44 minus.t11 a_n1724_n1088# 0.029954f
C45 minus.t7 a_n1724_n1088# 0.029954f
C46 minus.n1 a_n1724_n1088# 0.041606f
C47 minus.n2 a_n1724_n1088# 0.076309f
C48 minus.t1 a_n1724_n1088# 0.029954f
C49 minus.t12 a_n1724_n1088# 0.029954f
C50 minus.t8 a_n1724_n1088# 0.038121f
C51 minus.n3 a_n1724_n1088# 0.039881f
C52 minus.n4 a_n1724_n1088# 0.030862f
C53 minus.n5 a_n1724_n1088# 0.013341f
C54 minus.n6 a_n1724_n1088# 0.030862f
C55 minus.n7 a_n1724_n1088# 0.013341f
C56 minus.n8 a_n1724_n1088# 0.032389f
C57 minus.n9 a_n1724_n1088# 0.032389f
C58 minus.n10 a_n1724_n1088# 0.032389f
C59 minus.n11 a_n1724_n1088# 0.013341f
C60 minus.n12 a_n1724_n1088# 0.030862f
C61 minus.n13 a_n1724_n1088# 0.013341f
C62 minus.n14 a_n1724_n1088# 0.030862f
C63 minus.n15 a_n1724_n1088# 0.03983f
C64 minus.n16 a_n1724_n1088# 0.718135f
C65 minus.n17 a_n1724_n1088# 0.032389f
C66 minus.t4 a_n1724_n1088# 0.029954f
C67 minus.t6 a_n1724_n1088# 0.029954f
C68 minus.t10 a_n1724_n1088# 0.029954f
C69 minus.n18 a_n1724_n1088# 0.041606f
C70 minus.n19 a_n1724_n1088# 0.076309f
C71 minus.t2 a_n1724_n1088# 0.029954f
C72 minus.t3 a_n1724_n1088# 0.029954f
C73 minus.t9 a_n1724_n1088# 0.038121f
C74 minus.n20 a_n1724_n1088# 0.039881f
C75 minus.n21 a_n1724_n1088# 0.030862f
C76 minus.n22 a_n1724_n1088# 0.013341f
C77 minus.n23 a_n1724_n1088# 0.030862f
C78 minus.n24 a_n1724_n1088# 0.013341f
C79 minus.n25 a_n1724_n1088# 0.032389f
C80 minus.n26 a_n1724_n1088# 0.032389f
C81 minus.n27 a_n1724_n1088# 0.032389f
C82 minus.n28 a_n1724_n1088# 0.013341f
C83 minus.n29 a_n1724_n1088# 0.030862f
C84 minus.n30 a_n1724_n1088# 0.013341f
C85 minus.n31 a_n1724_n1088# 0.030862f
C86 minus.t13 a_n1724_n1088# 0.038121f
C87 minus.n32 a_n1724_n1088# 0.03983f
C88 minus.n33 a_n1724_n1088# 0.214531f
C89 minus.n34 a_n1724_n1088# 0.886062f
C90 drain_left.t2 a_n1724_n1088# 0.116666f
C91 drain_left.t11 a_n1724_n1088# 0.018785f
C92 drain_left.t9 a_n1724_n1088# 0.018785f
C93 drain_left.n0 a_n1724_n1088# 0.072995f
C94 drain_left.n1 a_n1724_n1088# 0.461348f
C95 drain_left.t12 a_n1724_n1088# 0.018785f
C96 drain_left.t6 a_n1724_n1088# 0.018785f
C97 drain_left.n2 a_n1724_n1088# 0.073579f
C98 drain_left.t4 a_n1724_n1088# 0.018785f
C99 drain_left.t13 a_n1724_n1088# 0.018785f
C100 drain_left.n3 a_n1724_n1088# 0.072995f
C101 drain_left.n4 a_n1724_n1088# 0.479289f
C102 drain_left.n5 a_n1724_n1088# 0.608073f
C103 drain_left.t10 a_n1724_n1088# 0.116666f
C104 drain_left.t7 a_n1724_n1088# 0.018785f
C105 drain_left.t3 a_n1724_n1088# 0.018785f
C106 drain_left.n6 a_n1724_n1088# 0.072995f
C107 drain_left.n7 a_n1724_n1088# 0.474422f
C108 drain_left.t0 a_n1724_n1088# 0.018785f
C109 drain_left.t8 a_n1724_n1088# 0.018785f
C110 drain_left.n8 a_n1724_n1088# 0.072995f
C111 drain_left.n9 a_n1724_n1088# 0.249443f
C112 drain_left.t5 a_n1724_n1088# 0.018785f
C113 drain_left.t1 a_n1724_n1088# 0.018785f
C114 drain_left.n10 a_n1724_n1088# 0.072995f
C115 drain_left.n11 a_n1724_n1088# 0.447313f
C116 source.t18 a_n1724_n1088# 0.141189f
C117 source.n0 a_n1724_n1088# 0.606245f
C118 source.t27 a_n1724_n1088# 0.025367f
C119 source.t15 a_n1724_n1088# 0.025367f
C120 source.n1 a_n1724_n1088# 0.082269f
C121 source.n2 a_n1724_n1088# 0.309506f
C122 source.t19 a_n1724_n1088# 0.025367f
C123 source.t20 a_n1724_n1088# 0.025367f
C124 source.n3 a_n1724_n1088# 0.082269f
C125 source.n4 a_n1724_n1088# 0.309506f
C126 source.t23 a_n1724_n1088# 0.025367f
C127 source.t24 a_n1724_n1088# 0.025367f
C128 source.n5 a_n1724_n1088# 0.082269f
C129 source.n6 a_n1724_n1088# 0.330014f
C130 source.t4 a_n1724_n1088# 0.141189f
C131 source.n7 a_n1724_n1088# 0.340277f
C132 source.t12 a_n1724_n1088# 0.025367f
C133 source.t6 a_n1724_n1088# 0.025367f
C134 source.n8 a_n1724_n1088# 0.082269f
C135 source.n9 a_n1724_n1088# 0.309506f
C136 source.t5 a_n1724_n1088# 0.025367f
C137 source.t1 a_n1724_n1088# 0.025367f
C138 source.n10 a_n1724_n1088# 0.082269f
C139 source.n11 a_n1724_n1088# 0.309506f
C140 source.t7 a_n1724_n1088# 0.025367f
C141 source.t11 a_n1724_n1088# 0.025367f
C142 source.n12 a_n1724_n1088# 0.082269f
C143 source.n13 a_n1724_n1088# 0.909383f
C144 source.t17 a_n1724_n1088# 0.025367f
C145 source.t22 a_n1724_n1088# 0.025367f
C146 source.n14 a_n1724_n1088# 0.082269f
C147 source.n15 a_n1724_n1088# 0.909383f
C148 source.t25 a_n1724_n1088# 0.025367f
C149 source.t16 a_n1724_n1088# 0.025367f
C150 source.n16 a_n1724_n1088# 0.082269f
C151 source.n17 a_n1724_n1088# 0.309506f
C152 source.t26 a_n1724_n1088# 0.025367f
C153 source.t21 a_n1724_n1088# 0.025367f
C154 source.n18 a_n1724_n1088# 0.082269f
C155 source.n19 a_n1724_n1088# 0.309506f
C156 source.t14 a_n1724_n1088# 0.141189f
C157 source.n20 a_n1724_n1088# 0.340277f
C158 source.t0 a_n1724_n1088# 0.025367f
C159 source.t3 a_n1724_n1088# 0.025367f
C160 source.n21 a_n1724_n1088# 0.082269f
C161 source.n22 a_n1724_n1088# 0.330014f
C162 source.t13 a_n1724_n1088# 0.025367f
C163 source.t2 a_n1724_n1088# 0.025367f
C164 source.n23 a_n1724_n1088# 0.082269f
C165 source.n24 a_n1724_n1088# 0.309506f
C166 source.t10 a_n1724_n1088# 0.025367f
C167 source.t8 a_n1724_n1088# 0.025367f
C168 source.n25 a_n1724_n1088# 0.082269f
C169 source.n26 a_n1724_n1088# 0.309506f
C170 source.t9 a_n1724_n1088# 0.141189f
C171 source.n27 a_n1724_n1088# 0.493398f
C172 source.n28 a_n1724_n1088# 0.650128f
C173 plus.n0 a_n1724_n1088# 0.033045f
C174 plus.t8 a_n1724_n1088# 0.03056f
C175 plus.t5 a_n1724_n1088# 0.03056f
C176 plus.t13 a_n1724_n1088# 0.03056f
C177 plus.n1 a_n1724_n1088# 0.042449f
C178 plus.n2 a_n1724_n1088# 0.077854f
C179 plus.t10 a_n1724_n1088# 0.03056f
C180 plus.t6 a_n1724_n1088# 0.03056f
C181 plus.t3 a_n1724_n1088# 0.038893f
C182 plus.n3 a_n1724_n1088# 0.040689f
C183 plus.n4 a_n1724_n1088# 0.031487f
C184 plus.n5 a_n1724_n1088# 0.013611f
C185 plus.n6 a_n1724_n1088# 0.031487f
C186 plus.n7 a_n1724_n1088# 0.013611f
C187 plus.n8 a_n1724_n1088# 0.033045f
C188 plus.n9 a_n1724_n1088# 0.033045f
C189 plus.n10 a_n1724_n1088# 0.033045f
C190 plus.n11 a_n1724_n1088# 0.013611f
C191 plus.n12 a_n1724_n1088# 0.031487f
C192 plus.n13 a_n1724_n1088# 0.013611f
C193 plus.n14 a_n1724_n1088# 0.031487f
C194 plus.t12 a_n1724_n1088# 0.038893f
C195 plus.n15 a_n1724_n1088# 0.040636f
C196 plus.n16 a_n1724_n1088# 0.229544f
C197 plus.n17 a_n1724_n1088# 0.033045f
C198 plus.t11 a_n1724_n1088# 0.038893f
C199 plus.t2 a_n1724_n1088# 0.03056f
C200 plus.t4 a_n1724_n1088# 0.03056f
C201 plus.t9 a_n1724_n1088# 0.03056f
C202 plus.n18 a_n1724_n1088# 0.042449f
C203 plus.n19 a_n1724_n1088# 0.077854f
C204 plus.t0 a_n1724_n1088# 0.03056f
C205 plus.t1 a_n1724_n1088# 0.03056f
C206 plus.t7 a_n1724_n1088# 0.038893f
C207 plus.n20 a_n1724_n1088# 0.040689f
C208 plus.n21 a_n1724_n1088# 0.031487f
C209 plus.n22 a_n1724_n1088# 0.013611f
C210 plus.n23 a_n1724_n1088# 0.031487f
C211 plus.n24 a_n1724_n1088# 0.013611f
C212 plus.n25 a_n1724_n1088# 0.033045f
C213 plus.n26 a_n1724_n1088# 0.033045f
C214 plus.n27 a_n1724_n1088# 0.033045f
C215 plus.n28 a_n1724_n1088# 0.013611f
C216 plus.n29 a_n1724_n1088# 0.031487f
C217 plus.n30 a_n1724_n1088# 0.013611f
C218 plus.n31 a_n1724_n1088# 0.031487f
C219 plus.n32 a_n1724_n1088# 0.040636f
C220 plus.n33 a_n1724_n1088# 0.711638f
.ends

