* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X1 drain_left.t13 plus.t0 source.t14 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X2 drain_left.t12 plus.t1 source.t24 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X3 source.t3 minus.t0 drain_right.t13 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X4 source.t27 plus.t2 drain_left.t11 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X5 drain_left.t10 plus.t3 source.t18 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X6 drain_left.t9 plus.t4 source.t21 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X7 drain_left.t8 plus.t5 source.t15 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X8 source.t5 minus.t1 drain_right.t12 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X9 drain_right.t11 minus.t2 source.t7 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X10 a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X11 drain_right.t10 minus.t3 source.t9 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X12 drain_right.t9 minus.t4 source.t1 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X13 source.t2 minus.t5 drain_right.t8 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X14 drain_right.t7 minus.t6 source.t4 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X15 drain_right.t6 minus.t7 source.t6 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X16 source.t26 plus.t6 drain_left.t7 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X17 drain_right.t5 minus.t8 source.t8 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X18 drain_left.t6 plus.t7 source.t25 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X19 source.t16 plus.t8 drain_left.t5 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X20 a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X21 source.t22 plus.t9 drain_left.t4 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X22 drain_right.t4 minus.t9 source.t11 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X23 a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X24 source.t19 plus.t10 drain_left.t3 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X25 drain_right.t3 minus.t10 source.t0 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X26 source.t10 minus.t11 drain_right.t2 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X27 drain_left.t2 plus.t11 source.t17 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X28 source.t13 minus.t12 drain_right.t1 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X29 source.t12 minus.t13 drain_right.t0 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X30 source.t23 plus.t12 drain_left.t1 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X31 drain_left.t0 plus.t13 source.t20 a_n2364_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n8 plus.n7 161.3
R1 plus.n9 plus.n4 161.3
R2 plus.n11 plus.n10 161.3
R3 plus.n12 plus.n3 161.3
R4 plus.n14 plus.n13 161.3
R5 plus.n15 plus.n2 161.3
R6 plus.n17 plus.n16 161.3
R7 plus.n18 plus.n1 161.3
R8 plus.n19 plus.n0 161.3
R9 plus.n21 plus.n20 161.3
R10 plus.n30 plus.n29 161.3
R11 plus.n31 plus.n26 161.3
R12 plus.n33 plus.n32 161.3
R13 plus.n34 plus.n25 161.3
R14 plus.n36 plus.n35 161.3
R15 plus.n37 plus.n24 161.3
R16 plus.n39 plus.n38 161.3
R17 plus.n40 plus.n23 161.3
R18 plus.n41 plus.n22 161.3
R19 plus.n43 plus.n42 161.3
R20 plus.n5 plus.t5 114.394
R21 plus.n27 plus.t7 114.394
R22 plus.n20 plus.t0 90.5476
R23 plus.n18 plus.t9 90.5476
R24 plus.n2 plus.t4 90.5476
R25 plus.n12 plus.t8 90.5476
R26 plus.n4 plus.t1 90.5476
R27 plus.n6 plus.t10 90.5476
R28 plus.n42 plus.t3 90.5476
R29 plus.n40 plus.t2 90.5476
R30 plus.n24 plus.t13 90.5476
R31 plus.n34 plus.t12 90.5476
R32 plus.n26 plus.t11 90.5476
R33 plus.n28 plus.t6 90.5476
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus.n18 plus.n17 30.6732
R39 plus.n7 plus.n6 30.6732
R40 plus.n40 plus.n39 30.6732
R41 plus.n29 plus.n28 30.6732
R42 plus plus.n43 27.9403
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus.n19 plus.n18 13.146
R58 plus.n41 plus.n40 13.146
R59 plus plus.n21 8.12739
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n0 source.t14 243.255
R79 source.n7 source.t11 243.255
R80 source.n27 source.t0 243.254
R81 source.n20 source.t25 243.254
R82 source.n2 source.n1 223.454
R83 source.n4 source.n3 223.454
R84 source.n6 source.n5 223.454
R85 source.n9 source.n8 223.454
R86 source.n11 source.n10 223.454
R87 source.n13 source.n12 223.454
R88 source.n26 source.n25 223.453
R89 source.n24 source.n23 223.453
R90 source.n22 source.n21 223.453
R91 source.n19 source.n18 223.453
R92 source.n17 source.n16 223.453
R93 source.n15 source.n14 223.453
R94 source.n25 source.t6 19.8005
R95 source.n25 source.t10 19.8005
R96 source.n23 source.t4 19.8005
R97 source.n23 source.t2 19.8005
R98 source.n21 source.t7 19.8005
R99 source.n21 source.t5 19.8005
R100 source.n18 source.t17 19.8005
R101 source.n18 source.t26 19.8005
R102 source.n16 source.t20 19.8005
R103 source.n16 source.t23 19.8005
R104 source.n14 source.t18 19.8005
R105 source.n14 source.t27 19.8005
R106 source.n1 source.t21 19.8005
R107 source.n1 source.t22 19.8005
R108 source.n3 source.t24 19.8005
R109 source.n3 source.t16 19.8005
R110 source.n5 source.t15 19.8005
R111 source.n5 source.t19 19.8005
R112 source.n8 source.t8 19.8005
R113 source.n8 source.t3 19.8005
R114 source.n10 source.t1 19.8005
R115 source.n10 source.t13 19.8005
R116 source.n12 source.t9 19.8005
R117 source.n12 source.t12 19.8005
R118 source.n15 source.n13 14.7303
R119 source.n28 source.n0 8.13543
R120 source.n28 source.n27 5.7074
R121 source.n7 source.n6 0.914293
R122 source.n22 source.n20 0.914293
R123 source.n13 source.n11 0.888431
R124 source.n11 source.n9 0.888431
R125 source.n9 source.n7 0.888431
R126 source.n6 source.n4 0.888431
R127 source.n4 source.n2 0.888431
R128 source.n2 source.n0 0.888431
R129 source.n17 source.n15 0.888431
R130 source.n19 source.n17 0.888431
R131 source.n20 source.n19 0.888431
R132 source.n24 source.n22 0.888431
R133 source.n26 source.n24 0.888431
R134 source.n27 source.n26 0.888431
R135 source source.n28 0.188
R136 drain_left.n7 drain_left.t8 260.82
R137 drain_left.n1 drain_left.t10 260.82
R138 drain_left.n4 drain_left.n2 241.019
R139 drain_left.n11 drain_left.n10 240.132
R140 drain_left.n9 drain_left.n8 240.132
R141 drain_left.n7 drain_left.n6 240.132
R142 drain_left.n4 drain_left.n3 240.131
R143 drain_left.n1 drain_left.n0 240.131
R144 drain_left drain_left.n5 24.1393
R145 drain_left.n2 drain_left.t7 19.8005
R146 drain_left.n2 drain_left.t6 19.8005
R147 drain_left.n3 drain_left.t1 19.8005
R148 drain_left.n3 drain_left.t2 19.8005
R149 drain_left.n0 drain_left.t11 19.8005
R150 drain_left.n0 drain_left.t0 19.8005
R151 drain_left.n10 drain_left.t4 19.8005
R152 drain_left.n10 drain_left.t13 19.8005
R153 drain_left.n8 drain_left.t5 19.8005
R154 drain_left.n8 drain_left.t9 19.8005
R155 drain_left.n6 drain_left.t3 19.8005
R156 drain_left.n6 drain_left.t12 19.8005
R157 drain_left drain_left.n11 6.54115
R158 drain_left.n9 drain_left.n7 0.888431
R159 drain_left.n11 drain_left.n9 0.888431
R160 drain_left.n5 drain_left.n1 0.611102
R161 drain_left.n5 drain_left.n4 0.167137
R162 minus.n21 minus.n20 161.3
R163 minus.n19 minus.n0 161.3
R164 minus.n18 minus.n17 161.3
R165 minus.n16 minus.n1 161.3
R166 minus.n15 minus.n14 161.3
R167 minus.n13 minus.n2 161.3
R168 minus.n12 minus.n11 161.3
R169 minus.n10 minus.n3 161.3
R170 minus.n9 minus.n8 161.3
R171 minus.n7 minus.n4 161.3
R172 minus.n43 minus.n42 161.3
R173 minus.n41 minus.n22 161.3
R174 minus.n40 minus.n39 161.3
R175 minus.n38 minus.n23 161.3
R176 minus.n37 minus.n36 161.3
R177 minus.n35 minus.n24 161.3
R178 minus.n34 minus.n33 161.3
R179 minus.n32 minus.n25 161.3
R180 minus.n31 minus.n30 161.3
R181 minus.n29 minus.n26 161.3
R182 minus.n5 minus.t9 114.394
R183 minus.n27 minus.t2 114.394
R184 minus.n6 minus.t0 90.5476
R185 minus.n8 minus.t8 90.5476
R186 minus.n12 minus.t12 90.5476
R187 minus.n14 minus.t4 90.5476
R188 minus.n18 minus.t13 90.5476
R189 minus.n20 minus.t3 90.5476
R190 minus.n28 minus.t1 90.5476
R191 minus.n30 minus.t6 90.5476
R192 minus.n34 minus.t5 90.5476
R193 minus.n36 minus.t7 90.5476
R194 minus.n40 minus.t11 90.5476
R195 minus.n42 minus.t10 90.5476
R196 minus.n5 minus.n4 44.9119
R197 minus.n27 minus.n26 44.9119
R198 minus.n20 minus.n19 35.055
R199 minus.n42 minus.n41 35.055
R200 minus.n7 minus.n6 30.6732
R201 minus.n18 minus.n1 30.6732
R202 minus.n29 minus.n28 30.6732
R203 minus.n40 minus.n23 30.6732
R204 minus.n44 minus.n21 29.8925
R205 minus.n8 minus.n3 26.2914
R206 minus.n14 minus.n13 26.2914
R207 minus.n30 minus.n25 26.2914
R208 minus.n36 minus.n35 26.2914
R209 minus.n12 minus.n3 21.9096
R210 minus.n13 minus.n12 21.9096
R211 minus.n34 minus.n25 21.9096
R212 minus.n35 minus.n34 21.9096
R213 minus.n6 minus.n5 17.739
R214 minus.n28 minus.n27 17.739
R215 minus.n8 minus.n7 17.5278
R216 minus.n14 minus.n1 17.5278
R217 minus.n30 minus.n29 17.5278
R218 minus.n36 minus.n23 17.5278
R219 minus.n19 minus.n18 13.146
R220 minus.n41 minus.n40 13.146
R221 minus.n44 minus.n43 6.65012
R222 minus.n21 minus.n0 0.189894
R223 minus.n17 minus.n0 0.189894
R224 minus.n17 minus.n16 0.189894
R225 minus.n16 minus.n15 0.189894
R226 minus.n15 minus.n2 0.189894
R227 minus.n11 minus.n2 0.189894
R228 minus.n11 minus.n10 0.189894
R229 minus.n10 minus.n9 0.189894
R230 minus.n9 minus.n4 0.189894
R231 minus.n31 minus.n26 0.189894
R232 minus.n32 minus.n31 0.189894
R233 minus.n33 minus.n32 0.189894
R234 minus.n33 minus.n24 0.189894
R235 minus.n37 minus.n24 0.189894
R236 minus.n38 minus.n37 0.189894
R237 minus.n39 minus.n38 0.189894
R238 minus.n39 minus.n22 0.189894
R239 minus.n43 minus.n22 0.189894
R240 minus minus.n44 0.188
R241 drain_right.n1 drain_right.t11 260.82
R242 drain_right.n11 drain_right.t10 259.933
R243 drain_right.n8 drain_right.n6 241.02
R244 drain_right.n4 drain_right.n2 241.019
R245 drain_right.n8 drain_right.n7 240.132
R246 drain_right.n10 drain_right.n9 240.132
R247 drain_right.n4 drain_right.n3 240.131
R248 drain_right.n1 drain_right.n0 240.131
R249 drain_right drain_right.n5 23.5861
R250 drain_right.n2 drain_right.t2 19.8005
R251 drain_right.n2 drain_right.t3 19.8005
R252 drain_right.n3 drain_right.t8 19.8005
R253 drain_right.n3 drain_right.t6 19.8005
R254 drain_right.n0 drain_right.t12 19.8005
R255 drain_right.n0 drain_right.t7 19.8005
R256 drain_right.n6 drain_right.t13 19.8005
R257 drain_right.n6 drain_right.t4 19.8005
R258 drain_right.n7 drain_right.t1 19.8005
R259 drain_right.n7 drain_right.t5 19.8005
R260 drain_right.n9 drain_right.t0 19.8005
R261 drain_right.n9 drain_right.t9 19.8005
R262 drain_right drain_right.n11 6.09718
R263 drain_right.n11 drain_right.n10 0.888431
R264 drain_right.n10 drain_right.n8 0.888431
R265 drain_right.n5 drain_right.n1 0.611102
R266 drain_right.n5 drain_right.n4 0.167137
C0 plus source 1.87953f
C1 minus drain_right 1.25562f
C2 minus source 1.86562f
C3 drain_left drain_right 1.23045f
C4 drain_left source 4.4989f
C5 plus minus 4.06494f
C6 drain_right source 4.49956f
C7 drain_left plus 1.48844f
C8 drain_left minus 0.180645f
C9 plus drain_right 0.39862f
C10 drain_right a_n2364_n1088# 4.10848f
C11 drain_left a_n2364_n1088# 4.41968f
C12 source a_n2364_n1088# 2.339747f
C13 minus a_n2364_n1088# 8.45389f
C14 plus a_n2364_n1088# 9.062241f
C15 drain_right.t11 a_n2364_n1088# 0.097419f
C16 drain_right.t12 a_n2364_n1088# 0.015634f
C17 drain_right.t7 a_n2364_n1088# 0.015634f
C18 drain_right.n0 a_n2364_n1088# 0.060751f
C19 drain_right.n1 a_n2364_n1088# 0.44354f
C20 drain_right.t2 a_n2364_n1088# 0.015634f
C21 drain_right.t3 a_n2364_n1088# 0.015634f
C22 drain_right.n2 a_n2364_n1088# 0.061707f
C23 drain_right.t8 a_n2364_n1088# 0.015634f
C24 drain_right.t6 a_n2364_n1088# 0.015634f
C25 drain_right.n3 a_n2364_n1088# 0.060751f
C26 drain_right.n4 a_n2364_n1088# 0.466917f
C27 drain_right.n5 a_n2364_n1088# 0.611519f
C28 drain_right.t13 a_n2364_n1088# 0.015634f
C29 drain_right.t4 a_n2364_n1088# 0.015634f
C30 drain_right.n6 a_n2364_n1088# 0.061707f
C31 drain_right.t1 a_n2364_n1088# 0.015634f
C32 drain_right.t5 a_n2364_n1088# 0.015634f
C33 drain_right.n7 a_n2364_n1088# 0.060751f
C34 drain_right.n8 a_n2364_n1088# 0.510147f
C35 drain_right.t0 a_n2364_n1088# 0.015634f
C36 drain_right.t9 a_n2364_n1088# 0.015634f
C37 drain_right.n9 a_n2364_n1088# 0.060751f
C38 drain_right.n10 a_n2364_n1088# 0.251567f
C39 drain_right.t10 a_n2364_n1088# 0.096705f
C40 drain_right.n11 a_n2364_n1088# 0.391446f
C41 minus.n0 a_n2364_n1088# 0.025826f
C42 minus.n1 a_n2364_n1088# 0.005861f
C43 minus.t13 a_n2364_n1088# 0.061304f
C44 minus.n2 a_n2364_n1088# 0.025826f
C45 minus.n3 a_n2364_n1088# 0.005861f
C46 minus.t12 a_n2364_n1088# 0.061304f
C47 minus.n4 a_n2364_n1088# 0.108817f
C48 minus.t9 a_n2364_n1088# 0.074014f
C49 minus.n5 a_n2364_n1088# 0.050479f
C50 minus.t0 a_n2364_n1088# 0.061304f
C51 minus.n6 a_n2364_n1088# 0.064144f
C52 minus.n7 a_n2364_n1088# 0.005861f
C53 minus.t8 a_n2364_n1088# 0.061304f
C54 minus.n8 a_n2364_n1088# 0.060944f
C55 minus.n9 a_n2364_n1088# 0.025826f
C56 minus.n10 a_n2364_n1088# 0.025826f
C57 minus.n11 a_n2364_n1088# 0.025826f
C58 minus.n12 a_n2364_n1088# 0.060944f
C59 minus.n13 a_n2364_n1088# 0.005861f
C60 minus.t4 a_n2364_n1088# 0.061304f
C61 minus.n14 a_n2364_n1088# 0.060944f
C62 minus.n15 a_n2364_n1088# 0.025826f
C63 minus.n16 a_n2364_n1088# 0.025826f
C64 minus.n17 a_n2364_n1088# 0.025826f
C65 minus.n18 a_n2364_n1088# 0.060944f
C66 minus.n19 a_n2364_n1088# 0.005861f
C67 minus.t3 a_n2364_n1088# 0.061304f
C68 minus.n20 a_n2364_n1088# 0.059989f
C69 minus.n21 a_n2364_n1088# 0.671363f
C70 minus.n22 a_n2364_n1088# 0.025826f
C71 minus.n23 a_n2364_n1088# 0.005861f
C72 minus.n24 a_n2364_n1088# 0.025826f
C73 minus.n25 a_n2364_n1088# 0.005861f
C74 minus.n26 a_n2364_n1088# 0.108817f
C75 minus.t2 a_n2364_n1088# 0.074014f
C76 minus.n27 a_n2364_n1088# 0.050479f
C77 minus.t1 a_n2364_n1088# 0.061304f
C78 minus.n28 a_n2364_n1088# 0.064144f
C79 minus.n29 a_n2364_n1088# 0.005861f
C80 minus.t6 a_n2364_n1088# 0.061304f
C81 minus.n30 a_n2364_n1088# 0.060944f
C82 minus.n31 a_n2364_n1088# 0.025826f
C83 minus.n32 a_n2364_n1088# 0.025826f
C84 minus.n33 a_n2364_n1088# 0.025826f
C85 minus.t5 a_n2364_n1088# 0.061304f
C86 minus.n34 a_n2364_n1088# 0.060944f
C87 minus.n35 a_n2364_n1088# 0.005861f
C88 minus.t7 a_n2364_n1088# 0.061304f
C89 minus.n36 a_n2364_n1088# 0.060944f
C90 minus.n37 a_n2364_n1088# 0.025826f
C91 minus.n38 a_n2364_n1088# 0.025826f
C92 minus.n39 a_n2364_n1088# 0.025826f
C93 minus.t11 a_n2364_n1088# 0.061304f
C94 minus.n40 a_n2364_n1088# 0.060944f
C95 minus.n41 a_n2364_n1088# 0.005861f
C96 minus.t10 a_n2364_n1088# 0.061304f
C97 minus.n42 a_n2364_n1088# 0.059989f
C98 minus.n43 a_n2364_n1088# 0.177916f
C99 minus.n44 a_n2364_n1088# 0.823853f
C100 drain_left.t10 a_n2364_n1088# 0.095771f
C101 drain_left.t11 a_n2364_n1088# 0.01537f
C102 drain_left.t0 a_n2364_n1088# 0.01537f
C103 drain_left.n0 a_n2364_n1088# 0.059723f
C104 drain_left.n1 a_n2364_n1088# 0.436041f
C105 drain_left.t7 a_n2364_n1088# 0.01537f
C106 drain_left.t6 a_n2364_n1088# 0.01537f
C107 drain_left.n2 a_n2364_n1088# 0.060663f
C108 drain_left.t1 a_n2364_n1088# 0.01537f
C109 drain_left.t2 a_n2364_n1088# 0.01537f
C110 drain_left.n3 a_n2364_n1088# 0.059723f
C111 drain_left.n4 a_n2364_n1088# 0.459023f
C112 drain_left.n5 a_n2364_n1088# 0.638642f
C113 drain_left.t8 a_n2364_n1088# 0.095772f
C114 drain_left.t3 a_n2364_n1088# 0.01537f
C115 drain_left.t12 a_n2364_n1088# 0.01537f
C116 drain_left.n6 a_n2364_n1088# 0.059723f
C117 drain_left.n7 a_n2364_n1088# 0.452683f
C118 drain_left.t5 a_n2364_n1088# 0.01537f
C119 drain_left.t9 a_n2364_n1088# 0.01537f
C120 drain_left.n8 a_n2364_n1088# 0.059723f
C121 drain_left.n9 a_n2364_n1088# 0.247314f
C122 drain_left.t4 a_n2364_n1088# 0.01537f
C123 drain_left.t13 a_n2364_n1088# 0.01537f
C124 drain_left.n10 a_n2364_n1088# 0.059723f
C125 drain_left.n11 a_n2364_n1088# 0.419351f
C126 source.t14 a_n2364_n1088# 0.1183f
C127 source.n0 a_n2364_n1088# 0.561331f
C128 source.t21 a_n2364_n1088# 0.021255f
C129 source.t22 a_n2364_n1088# 0.021255f
C130 source.n1 a_n2364_n1088# 0.068932f
C131 source.n2 a_n2364_n1088# 0.3191f
C132 source.t24 a_n2364_n1088# 0.021255f
C133 source.t16 a_n2364_n1088# 0.021255f
C134 source.n3 a_n2364_n1088# 0.068932f
C135 source.n4 a_n2364_n1088# 0.3191f
C136 source.t15 a_n2364_n1088# 0.021255f
C137 source.t19 a_n2364_n1088# 0.021255f
C138 source.n5 a_n2364_n1088# 0.068932f
C139 source.n6 a_n2364_n1088# 0.321341f
C140 source.t11 a_n2364_n1088# 0.1183f
C141 source.n7 a_n2364_n1088# 0.32994f
C142 source.t8 a_n2364_n1088# 0.021255f
C143 source.t3 a_n2364_n1088# 0.021255f
C144 source.n8 a_n2364_n1088# 0.068932f
C145 source.n9 a_n2364_n1088# 0.3191f
C146 source.t1 a_n2364_n1088# 0.021255f
C147 source.t13 a_n2364_n1088# 0.021255f
C148 source.n10 a_n2364_n1088# 0.068932f
C149 source.n11 a_n2364_n1088# 0.3191f
C150 source.t9 a_n2364_n1088# 0.021255f
C151 source.t12 a_n2364_n1088# 0.021255f
C152 source.n12 a_n2364_n1088# 0.068932f
C153 source.n13 a_n2364_n1088# 0.851612f
C154 source.t18 a_n2364_n1088# 0.021255f
C155 source.t27 a_n2364_n1088# 0.021255f
C156 source.n14 a_n2364_n1088# 0.068932f
C157 source.n15 a_n2364_n1088# 0.851612f
C158 source.t20 a_n2364_n1088# 0.021255f
C159 source.t23 a_n2364_n1088# 0.021255f
C160 source.n16 a_n2364_n1088# 0.068932f
C161 source.n17 a_n2364_n1088# 0.3191f
C162 source.t17 a_n2364_n1088# 0.021255f
C163 source.t26 a_n2364_n1088# 0.021255f
C164 source.n18 a_n2364_n1088# 0.068932f
C165 source.n19 a_n2364_n1088# 0.3191f
C166 source.t25 a_n2364_n1088# 0.1183f
C167 source.n20 a_n2364_n1088# 0.32994f
C168 source.t7 a_n2364_n1088# 0.021255f
C169 source.t5 a_n2364_n1088# 0.021255f
C170 source.n21 a_n2364_n1088# 0.068932f
C171 source.n22 a_n2364_n1088# 0.321341f
C172 source.t4 a_n2364_n1088# 0.021255f
C173 source.t2 a_n2364_n1088# 0.021255f
C174 source.n23 a_n2364_n1088# 0.068932f
C175 source.n24 a_n2364_n1088# 0.3191f
C176 source.t6 a_n2364_n1088# 0.021255f
C177 source.t10 a_n2364_n1088# 0.021255f
C178 source.n25 a_n2364_n1088# 0.068932f
C179 source.n26 a_n2364_n1088# 0.3191f
C180 source.t0 a_n2364_n1088# 0.1183f
C181 source.n27 a_n2364_n1088# 0.466912f
C182 source.n28 a_n2364_n1088# 0.557401f
C183 plus.n0 a_n2364_n1088# 0.02616f
C184 plus.t0 a_n2364_n1088# 0.062095f
C185 plus.t9 a_n2364_n1088# 0.062095f
C186 plus.n1 a_n2364_n1088# 0.02616f
C187 plus.t4 a_n2364_n1088# 0.062095f
C188 plus.n2 a_n2364_n1088# 0.061731f
C189 plus.n3 a_n2364_n1088# 0.02616f
C190 plus.t8 a_n2364_n1088# 0.062095f
C191 plus.t1 a_n2364_n1088# 0.062095f
C192 plus.n4 a_n2364_n1088# 0.061731f
C193 plus.t5 a_n2364_n1088# 0.074969f
C194 plus.n5 a_n2364_n1088# 0.05113f
C195 plus.t10 a_n2364_n1088# 0.062095f
C196 plus.n6 a_n2364_n1088# 0.064971f
C197 plus.n7 a_n2364_n1088# 0.005936f
C198 plus.n8 a_n2364_n1088# 0.110221f
C199 plus.n9 a_n2364_n1088# 0.02616f
C200 plus.n10 a_n2364_n1088# 0.02616f
C201 plus.n11 a_n2364_n1088# 0.005936f
C202 plus.n12 a_n2364_n1088# 0.061731f
C203 plus.n13 a_n2364_n1088# 0.005936f
C204 plus.n14 a_n2364_n1088# 0.02616f
C205 plus.n15 a_n2364_n1088# 0.02616f
C206 plus.n16 a_n2364_n1088# 0.02616f
C207 plus.n17 a_n2364_n1088# 0.005936f
C208 plus.n18 a_n2364_n1088# 0.061731f
C209 plus.n19 a_n2364_n1088# 0.005936f
C210 plus.n20 a_n2364_n1088# 0.060763f
C211 plus.n21 a_n2364_n1088# 0.189037f
C212 plus.n22 a_n2364_n1088# 0.02616f
C213 plus.t3 a_n2364_n1088# 0.062095f
C214 plus.n23 a_n2364_n1088# 0.02616f
C215 plus.t2 a_n2364_n1088# 0.062095f
C216 plus.t13 a_n2364_n1088# 0.062095f
C217 plus.n24 a_n2364_n1088# 0.061731f
C218 plus.n25 a_n2364_n1088# 0.02616f
C219 plus.t12 a_n2364_n1088# 0.062095f
C220 plus.t11 a_n2364_n1088# 0.062095f
C221 plus.n26 a_n2364_n1088# 0.061731f
C222 plus.t7 a_n2364_n1088# 0.074969f
C223 plus.n27 a_n2364_n1088# 0.05113f
C224 plus.t6 a_n2364_n1088# 0.062095f
C225 plus.n28 a_n2364_n1088# 0.064971f
C226 plus.n29 a_n2364_n1088# 0.005936f
C227 plus.n30 a_n2364_n1088# 0.110221f
C228 plus.n31 a_n2364_n1088# 0.02616f
C229 plus.n32 a_n2364_n1088# 0.02616f
C230 plus.n33 a_n2364_n1088# 0.005936f
C231 plus.n34 a_n2364_n1088# 0.061731f
C232 plus.n35 a_n2364_n1088# 0.005936f
C233 plus.n36 a_n2364_n1088# 0.02616f
C234 plus.n37 a_n2364_n1088# 0.02616f
C235 plus.n38 a_n2364_n1088# 0.02616f
C236 plus.n39 a_n2364_n1088# 0.005936f
C237 plus.n40 a_n2364_n1088# 0.061731f
C238 plus.n41 a_n2364_n1088# 0.005936f
C239 plus.n42 a_n2364_n1088# 0.060763f
C240 plus.n43 a_n2364_n1088# 0.656771f
.ends

