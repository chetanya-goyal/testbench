* NGSPICE file created from diffpair604.ext - technology: sky130A

.subckt diffpair604 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t13 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t14 plus.t1 drain_left.t8 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X3 source.t15 minus.t0 drain_right.t9 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X4 source.t7 plus.t2 drain_left.t7 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X5 drain_left.t6 plus.t3 source.t6 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X6 drain_left.t5 plus.t4 source.t12 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X7 source.t16 minus.t1 drain_right.t8 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X8 drain_right.t7 minus.t2 source.t17 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X9 drain_right.t6 minus.t3 source.t18 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X10 drain_right.t5 minus.t4 source.t0 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X11 a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X12 drain_right.t4 minus.t5 source.t19 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X13 source.t11 plus.t5 drain_left.t4 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X14 drain_left.t3 plus.t6 source.t10 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X15 a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X16 source.t2 minus.t6 drain_right.t3 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X17 drain_right.t2 minus.t7 source.t3 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X18 drain_right.t1 minus.t8 source.t4 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X19 source.t5 plus.t7 drain_left.t2 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X20 source.t1 minus.t9 drain_right.t0 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X21 drain_left.t1 plus.t8 source.t9 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X22 drain_left.t0 plus.t9 source.t8 a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X23 a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# a_n1712_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
R0 plus.n2 plus.t4 1063.55
R1 plus.n14 plus.t0 1063.55
R2 plus.n10 plus.t8 1042.57
R3 plus.n9 plus.t5 1042.57
R4 plus.n1 plus.t9 1042.57
R5 plus.n3 plus.t7 1042.57
R6 plus.n22 plus.t3 1042.57
R7 plus.n21 plus.t2 1042.57
R8 plus.n13 plus.t6 1042.57
R9 plus.n15 plus.t1 1042.57
R10 plus.n5 plus.n4 161.3
R11 plus.n6 plus.n1 161.3
R12 plus.n8 plus.n7 161.3
R13 plus.n9 plus.n0 161.3
R14 plus.n11 plus.n10 161.3
R15 plus.n17 plus.n16 161.3
R16 plus.n18 plus.n13 161.3
R17 plus.n20 plus.n19 161.3
R18 plus.n21 plus.n12 161.3
R19 plus.n23 plus.n22 161.3
R20 plus.n5 plus.n2 70.4033
R21 plus.n17 plus.n14 70.4033
R22 plus.n10 plus.n9 48.2005
R23 plus.n22 plus.n21 48.2005
R24 plus.n8 plus.n1 36.5157
R25 plus.n4 plus.n1 36.5157
R26 plus.n20 plus.n13 36.5157
R27 plus.n16 plus.n13 36.5157
R28 plus plus.n23 32.5805
R29 plus.n3 plus.n2 20.9576
R30 plus.n15 plus.n14 20.9576
R31 plus plus.n11 15.2372
R32 plus.n9 plus.n8 11.6853
R33 plus.n4 plus.n3 11.6853
R34 plus.n21 plus.n20 11.6853
R35 plus.n16 plus.n15 11.6853
R36 plus.n6 plus.n5 0.189894
R37 plus.n7 plus.n6 0.189894
R38 plus.n7 plus.n0 0.189894
R39 plus.n11 plus.n0 0.189894
R40 plus.n23 plus.n12 0.189894
R41 plus.n19 plus.n12 0.189894
R42 plus.n19 plus.n18 0.189894
R43 plus.n18 plus.n17 0.189894
R44 source.n0 source.t9 44.1297
R45 source.n5 source.t3 44.1296
R46 source.n19 source.t19 44.1295
R47 source.n14 source.t13 44.1295
R48 source.n2 source.n1 43.1397
R49 source.n4 source.n3 43.1397
R50 source.n7 source.n6 43.1397
R51 source.n9 source.n8 43.1397
R52 source.n18 source.n17 43.1396
R53 source.n16 source.n15 43.1396
R54 source.n13 source.n12 43.1396
R55 source.n11 source.n10 43.1396
R56 source.n11 source.n9 28.7794
R57 source.n20 source.n0 22.4432
R58 source.n20 source.n19 5.62119
R59 source.n17 source.t4 0.9905
R60 source.n17 source.t2 0.9905
R61 source.n15 source.t17 0.9905
R62 source.n15 source.t16 0.9905
R63 source.n12 source.t10 0.9905
R64 source.n12 source.t14 0.9905
R65 source.n10 source.t6 0.9905
R66 source.n10 source.t7 0.9905
R67 source.n1 source.t8 0.9905
R68 source.n1 source.t11 0.9905
R69 source.n3 source.t12 0.9905
R70 source.n3 source.t5 0.9905
R71 source.n6 source.t0 0.9905
R72 source.n6 source.t15 0.9905
R73 source.n8 source.t18 0.9905
R74 source.n8 source.t1 0.9905
R75 source.n5 source.n4 0.828086
R76 source.n16 source.n14 0.828086
R77 source.n9 source.n7 0.716017
R78 source.n7 source.n5 0.716017
R79 source.n4 source.n2 0.716017
R80 source.n2 source.n0 0.716017
R81 source.n13 source.n11 0.716017
R82 source.n14 source.n13 0.716017
R83 source.n18 source.n16 0.716017
R84 source.n19 source.n18 0.716017
R85 source source.n20 0.188
R86 drain_left.n5 drain_left.t5 61.5239
R87 drain_left.n1 drain_left.t6 61.5238
R88 drain_left.n3 drain_left.n2 60.2997
R89 drain_left.n7 drain_left.n6 59.8185
R90 drain_left.n5 drain_left.n4 59.8185
R91 drain_left.n1 drain_left.n0 59.8184
R92 drain_left drain_left.n3 36.4686
R93 drain_left drain_left.n7 6.36873
R94 drain_left.n2 drain_left.t8 0.9905
R95 drain_left.n2 drain_left.t9 0.9905
R96 drain_left.n0 drain_left.t7 0.9905
R97 drain_left.n0 drain_left.t3 0.9905
R98 drain_left.n6 drain_left.t4 0.9905
R99 drain_left.n6 drain_left.t1 0.9905
R100 drain_left.n4 drain_left.t2 0.9905
R101 drain_left.n4 drain_left.t0 0.9905
R102 drain_left.n7 drain_left.n5 0.716017
R103 drain_left.n3 drain_left.n1 0.124033
R104 minus.n2 minus.t7 1063.55
R105 minus.n14 minus.t2 1063.55
R106 minus.n3 minus.t0 1042.57
R107 minus.n1 minus.t4 1042.57
R108 minus.n9 minus.t9 1042.57
R109 minus.n10 minus.t3 1042.57
R110 minus.n15 minus.t1 1042.57
R111 minus.n13 minus.t8 1042.57
R112 minus.n21 minus.t6 1042.57
R113 minus.n22 minus.t5 1042.57
R114 minus.n11 minus.n10 161.3
R115 minus.n9 minus.n0 161.3
R116 minus.n8 minus.n7 161.3
R117 minus.n6 minus.n1 161.3
R118 minus.n5 minus.n4 161.3
R119 minus.n23 minus.n22 161.3
R120 minus.n21 minus.n12 161.3
R121 minus.n20 minus.n19 161.3
R122 minus.n18 minus.n13 161.3
R123 minus.n17 minus.n16 161.3
R124 minus.n5 minus.n2 70.4033
R125 minus.n17 minus.n14 70.4033
R126 minus.n10 minus.n9 48.2005
R127 minus.n22 minus.n21 48.2005
R128 minus.n24 minus.n11 41.7297
R129 minus.n4 minus.n1 36.5157
R130 minus.n8 minus.n1 36.5157
R131 minus.n16 minus.n13 36.5157
R132 minus.n20 minus.n13 36.5157
R133 minus.n3 minus.n2 20.9576
R134 minus.n15 minus.n14 20.9576
R135 minus.n4 minus.n3 11.6853
R136 minus.n9 minus.n8 11.6853
R137 minus.n16 minus.n15 11.6853
R138 minus.n21 minus.n20 11.6853
R139 minus.n24 minus.n23 6.563
R140 minus.n11 minus.n0 0.189894
R141 minus.n7 minus.n0 0.189894
R142 minus.n7 minus.n6 0.189894
R143 minus.n6 minus.n5 0.189894
R144 minus.n18 minus.n17 0.189894
R145 minus.n19 minus.n18 0.189894
R146 minus.n19 minus.n12 0.189894
R147 minus.n23 minus.n12 0.189894
R148 minus minus.n24 0.188
R149 drain_right.n1 drain_right.t7 61.5238
R150 drain_right.n7 drain_right.t6 60.8084
R151 drain_right.n6 drain_right.n4 60.534
R152 drain_right.n3 drain_right.n2 60.2997
R153 drain_right.n6 drain_right.n5 59.8185
R154 drain_right.n1 drain_right.n0 59.8184
R155 drain_right drain_right.n3 35.9154
R156 drain_right drain_right.n7 6.01097
R157 drain_right.n2 drain_right.t3 0.9905
R158 drain_right.n2 drain_right.t4 0.9905
R159 drain_right.n0 drain_right.t8 0.9905
R160 drain_right.n0 drain_right.t1 0.9905
R161 drain_right.n4 drain_right.t9 0.9905
R162 drain_right.n4 drain_right.t2 0.9905
R163 drain_right.n5 drain_right.t0 0.9905
R164 drain_right.n5 drain_right.t5 0.9905
R165 drain_right.n7 drain_right.n6 0.716017
R166 drain_right.n3 drain_right.n1 0.124033
C0 plus source 8.35949f
C1 drain_left source 26.2633f
C2 drain_right minus 8.953719f
C3 plus drain_right 0.323418f
C4 drain_right drain_left 0.850048f
C5 drain_right source 26.2488f
C6 plus minus 6.76396f
C7 minus drain_left 0.171781f
C8 plus drain_left 9.11475f
C9 minus source 8.344509f
C10 drain_right a_n1712_n4888# 9.091459f
C11 drain_left a_n1712_n4888# 9.36224f
C12 source a_n1712_n4888# 9.220331f
C13 minus a_n1712_n4888# 7.200307f
C14 plus a_n1712_n4888# 9.50828f
C15 drain_right.t7 a_n1712_n4888# 4.81328f
C16 drain_right.t8 a_n1712_n4888# 0.411295f
C17 drain_right.t1 a_n1712_n4888# 0.411295f
C18 drain_right.n0 a_n1712_n4888# 3.76015f
C19 drain_right.n1 a_n1712_n4888# 0.653509f
C20 drain_right.t3 a_n1712_n4888# 0.411295f
C21 drain_right.t4 a_n1712_n4888# 0.411295f
C22 drain_right.n2 a_n1712_n4888# 3.76279f
C23 drain_right.n3 a_n1712_n4888# 2.03475f
C24 drain_right.t9 a_n1712_n4888# 0.411295f
C25 drain_right.t2 a_n1712_n4888# 0.411295f
C26 drain_right.n4 a_n1712_n4888# 3.76428f
C27 drain_right.t0 a_n1712_n4888# 0.411295f
C28 drain_right.t5 a_n1712_n4888# 0.411295f
C29 drain_right.n5 a_n1712_n4888# 3.76014f
C30 drain_right.n6 a_n1712_n4888# 0.685557f
C31 drain_right.t6 a_n1712_n4888# 4.80908f
C32 drain_right.n7 a_n1712_n4888# 0.591058f
C33 minus.n0 a_n1712_n4888# 0.047537f
C34 minus.t4 a_n1712_n4888# 1.34621f
C35 minus.n1 a_n1712_n4888# 0.510688f
C36 minus.t7 a_n1712_n4888# 1.35618f
C37 minus.n2 a_n1712_n4888# 0.496075f
C38 minus.t0 a_n1712_n4888# 1.34621f
C39 minus.n3 a_n1712_n4888# 0.50805f
C40 minus.n4 a_n1712_n4888# 0.010787f
C41 minus.n5 a_n1712_n4888# 0.151643f
C42 minus.n6 a_n1712_n4888# 0.047537f
C43 minus.n7 a_n1712_n4888# 0.047537f
C44 minus.n8 a_n1712_n4888# 0.010787f
C45 minus.t9 a_n1712_n4888# 1.34621f
C46 minus.n9 a_n1712_n4888# 0.50805f
C47 minus.t3 a_n1712_n4888# 1.34621f
C48 minus.n10 a_n1712_n4888# 0.505706f
C49 minus.n11 a_n1712_n4888# 2.08731f
C50 minus.n12 a_n1712_n4888# 0.047537f
C51 minus.t8 a_n1712_n4888# 1.34621f
C52 minus.n13 a_n1712_n4888# 0.510688f
C53 minus.t2 a_n1712_n4888# 1.35618f
C54 minus.n14 a_n1712_n4888# 0.496075f
C55 minus.t1 a_n1712_n4888# 1.34621f
C56 minus.n15 a_n1712_n4888# 0.50805f
C57 minus.n16 a_n1712_n4888# 0.010787f
C58 minus.n17 a_n1712_n4888# 0.151643f
C59 minus.n18 a_n1712_n4888# 0.047537f
C60 minus.n19 a_n1712_n4888# 0.047537f
C61 minus.n20 a_n1712_n4888# 0.010787f
C62 minus.t6 a_n1712_n4888# 1.34621f
C63 minus.n21 a_n1712_n4888# 0.50805f
C64 minus.t5 a_n1712_n4888# 1.34621f
C65 minus.n22 a_n1712_n4888# 0.505706f
C66 minus.n23 a_n1712_n4888# 0.317821f
C67 minus.n24 a_n1712_n4888# 2.49284f
C68 drain_left.t6 a_n1712_n4888# 4.82667f
C69 drain_left.t7 a_n1712_n4888# 0.412439f
C70 drain_left.t3 a_n1712_n4888# 0.412439f
C71 drain_left.n0 a_n1712_n4888# 3.77061f
C72 drain_left.n1 a_n1712_n4888# 0.655327f
C73 drain_left.t8 a_n1712_n4888# 0.412439f
C74 drain_left.t9 a_n1712_n4888# 0.412439f
C75 drain_left.n2 a_n1712_n4888# 3.77326f
C76 drain_left.n3 a_n1712_n4888# 2.09485f
C77 drain_left.t5 a_n1712_n4888# 4.82669f
C78 drain_left.t2 a_n1712_n4888# 0.412439f
C79 drain_left.t0 a_n1712_n4888# 0.412439f
C80 drain_left.n4 a_n1712_n4888# 3.7706f
C81 drain_left.n5 a_n1712_n4888# 0.700195f
C82 drain_left.t4 a_n1712_n4888# 0.412439f
C83 drain_left.t1 a_n1712_n4888# 0.412439f
C84 drain_left.n6 a_n1712_n4888# 3.7706f
C85 drain_left.n7 a_n1712_n4888# 0.564753f
C86 source.t9 a_n1712_n4888# 4.77813f
C87 source.n0 a_n1712_n4888# 2.05546f
C88 source.t8 a_n1712_n4888# 0.418093f
C89 source.t11 a_n1712_n4888# 0.418093f
C90 source.n1 a_n1712_n4888# 3.73793f
C91 source.n2 a_n1712_n4888# 0.393627f
C92 source.t12 a_n1712_n4888# 0.418093f
C93 source.t5 a_n1712_n4888# 0.418093f
C94 source.n3 a_n1712_n4888# 3.73793f
C95 source.n4 a_n1712_n4888# 0.40318f
C96 source.t3 a_n1712_n4888# 4.77814f
C97 source.n5 a_n1712_n4888# 0.503228f
C98 source.t0 a_n1712_n4888# 0.418093f
C99 source.t15 a_n1712_n4888# 0.418093f
C100 source.n6 a_n1712_n4888# 3.73793f
C101 source.n7 a_n1712_n4888# 0.393627f
C102 source.t18 a_n1712_n4888# 0.418093f
C103 source.t1 a_n1712_n4888# 0.418093f
C104 source.n8 a_n1712_n4888# 3.73793f
C105 source.n9 a_n1712_n4888# 2.49143f
C106 source.t6 a_n1712_n4888# 0.418093f
C107 source.t7 a_n1712_n4888# 0.418093f
C108 source.n10 a_n1712_n4888# 3.73794f
C109 source.n11 a_n1712_n4888# 2.49142f
C110 source.t10 a_n1712_n4888# 0.418093f
C111 source.t14 a_n1712_n4888# 0.418093f
C112 source.n12 a_n1712_n4888# 3.73794f
C113 source.n13 a_n1712_n4888# 0.393619f
C114 source.t13 a_n1712_n4888# 4.77811f
C115 source.n14 a_n1712_n4888# 0.503254f
C116 source.t17 a_n1712_n4888# 0.418093f
C117 source.t16 a_n1712_n4888# 0.418093f
C118 source.n15 a_n1712_n4888# 3.73794f
C119 source.n16 a_n1712_n4888# 0.403172f
C120 source.t4 a_n1712_n4888# 0.418093f
C121 source.t2 a_n1712_n4888# 0.418093f
C122 source.n17 a_n1712_n4888# 3.73794f
C123 source.n18 a_n1712_n4888# 0.393619f
C124 source.t19 a_n1712_n4888# 4.77811f
C125 source.n19 a_n1712_n4888# 0.63377f
C126 source.n20 a_n1712_n4888# 2.39059f
C127 plus.n0 a_n1712_n4888# 0.048124f
C128 plus.t8 a_n1712_n4888# 1.36281f
C129 plus.t5 a_n1712_n4888# 1.36281f
C130 plus.t9 a_n1712_n4888# 1.36281f
C131 plus.n1 a_n1712_n4888# 0.516989f
C132 plus.t4 a_n1712_n4888# 1.37291f
C133 plus.n2 a_n1712_n4888# 0.502195f
C134 plus.t7 a_n1712_n4888# 1.36281f
C135 plus.n3 a_n1712_n4888# 0.514318f
C136 plus.n4 a_n1712_n4888# 0.01092f
C137 plus.n5 a_n1712_n4888# 0.153514f
C138 plus.n6 a_n1712_n4888# 0.048124f
C139 plus.n7 a_n1712_n4888# 0.048124f
C140 plus.n8 a_n1712_n4888# 0.01092f
C141 plus.n9 a_n1712_n4888# 0.514318f
C142 plus.n10 a_n1712_n4888# 0.511945f
C143 plus.n11 a_n1712_n4888# 0.737692f
C144 plus.n12 a_n1712_n4888# 0.048124f
C145 plus.t3 a_n1712_n4888# 1.36281f
C146 plus.t2 a_n1712_n4888# 1.36281f
C147 plus.t6 a_n1712_n4888# 1.36281f
C148 plus.n13 a_n1712_n4888# 0.516989f
C149 plus.t0 a_n1712_n4888# 1.37291f
C150 plus.n14 a_n1712_n4888# 0.502195f
C151 plus.t1 a_n1712_n4888# 1.36281f
C152 plus.n15 a_n1712_n4888# 0.514318f
C153 plus.n16 a_n1712_n4888# 0.01092f
C154 plus.n17 a_n1712_n4888# 0.153514f
C155 plus.n18 a_n1712_n4888# 0.048124f
C156 plus.n19 a_n1712_n4888# 0.048124f
C157 plus.n20 a_n1712_n4888# 0.01092f
C158 plus.n21 a_n1712_n4888# 0.514318f
C159 plus.n22 a_n1712_n4888# 0.511945f
C160 plus.n23 a_n1712_n4888# 1.66949f
.ends

