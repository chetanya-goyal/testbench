* NGSPICE file created from diffpair165.ext - technology: sky130A

.subckt diffpair165 minus drain_right drain_left source plus
X0 source.t23 plus.t0 drain_left.t9 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X1 drain_right.t11 minus.t0 source.t9 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 source.t22 plus.t1 drain_left.t11 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X3 drain_left.t6 plus.t2 source.t21 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X4 drain_right.t10 minus.t1 source.t4 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X5 a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X6 a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X7 a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X8 drain_left.t10 plus.t3 source.t20 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X9 source.t8 minus.t2 drain_right.t9 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 source.t0 minus.t3 drain_right.t8 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X11 source.t10 minus.t4 drain_right.t7 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X12 source.t19 plus.t4 drain_left.t7 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X13 drain_right.t6 minus.t5 source.t1 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X14 drain_right.t5 minus.t6 source.t5 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X15 a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X16 source.t7 minus.t7 drain_right.t4 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 drain_left.t0 plus.t5 source.t18 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 source.t17 plus.t6 drain_left.t5 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X19 drain_right.t3 minus.t8 source.t3 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X20 drain_left.t1 plus.t7 source.t16 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X21 source.t6 minus.t9 drain_right.t2 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X22 drain_right.t1 minus.t10 source.t11 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 source.t15 plus.t8 drain_left.t8 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X24 drain_left.t2 plus.t9 source.t14 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X25 drain_left.t3 plus.t10 source.t13 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X26 source.t2 minus.t11 drain_right.t0 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X27 source.t12 plus.t11 drain_left.t4 a_n1626_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
R0 plus.n2 plus.t6 745.639
R1 plus.n13 plus.t9 745.639
R2 plus.n17 plus.t2 745.639
R3 plus.n28 plus.t0 745.639
R4 plus.n3 plus.t10 690.867
R5 plus.n4 plus.t8 690.867
R6 plus.n10 plus.t7 690.867
R7 plus.n12 plus.t11 690.867
R8 plus.n19 plus.t1 690.867
R9 plus.n18 plus.t5 690.867
R10 plus.n25 plus.t4 690.867
R11 plus.n27 plus.t3 690.867
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 62.0763
R27 plus.n11 plus.n10 62.0763
R28 plus.n26 plus.n25 62.0763
R29 plus.n20 plus.n18 62.0763
R30 plus.n3 plus.n2 40.1672
R31 plus.n13 plus.n12 40.1672
R32 plus.n28 plus.n27 40.1672
R33 plus.n19 plus.n17 40.1672
R34 plus.n5 plus.n3 32.8641
R35 plus.n12 plus.n11 32.8641
R36 plus.n27 plus.n26 32.8641
R37 plus.n20 plus.n19 32.8641
R38 plus plus.n29 25.7945
R39 plus.n4 plus.n1 10.955
R40 plus.n10 plus.n9 10.955
R41 plus.n25 plus.n24 10.955
R42 plus.n18 plus.n16 10.955
R43 plus plus.n14 8.77702
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 drain_left.n6 drain_left.n4 80.3335
R53 drain_left.n3 drain_left.n2 80.278
R54 drain_left.n3 drain_left.n0 80.278
R55 drain_left.n8 drain_left.n7 79.7731
R56 drain_left.n6 drain_left.n5 79.7731
R57 drain_left.n3 drain_left.n1 79.773
R58 drain_left drain_left.n3 23.3506
R59 drain_left.n1 drain_left.t7 10.0005
R60 drain_left.n1 drain_left.t0 10.0005
R61 drain_left.n2 drain_left.t11 10.0005
R62 drain_left.n2 drain_left.t6 10.0005
R63 drain_left.n0 drain_left.t9 10.0005
R64 drain_left.n0 drain_left.t10 10.0005
R65 drain_left.n7 drain_left.t4 10.0005
R66 drain_left.n7 drain_left.t2 10.0005
R67 drain_left.n5 drain_left.t8 10.0005
R68 drain_left.n5 drain_left.t1 10.0005
R69 drain_left.n4 drain_left.t5 10.0005
R70 drain_left.n4 drain_left.t3 10.0005
R71 drain_left drain_left.n8 6.21356
R72 drain_left.n8 drain_left.n6 0.560845
R73 source.n0 source.t14 73.0943
R74 source.n5 source.t17 73.0943
R75 source.n6 source.t1 73.0943
R76 source.n11 source.t6 73.0943
R77 source.n23 source.t4 73.0942
R78 source.n18 source.t0 73.0942
R79 source.n17 source.t21 73.0942
R80 source.n12 source.t23 73.0942
R81 source.n2 source.n1 63.0943
R82 source.n4 source.n3 63.0943
R83 source.n8 source.n7 63.0943
R84 source.n10 source.n9 63.0943
R85 source.n22 source.n21 63.0942
R86 source.n20 source.n19 63.0942
R87 source.n16 source.n15 63.0942
R88 source.n14 source.n13 63.0942
R89 source.n12 source.n11 15.0299
R90 source.n21 source.t11 10.0005
R91 source.n21 source.t8 10.0005
R92 source.n19 source.t9 10.0005
R93 source.n19 source.t2 10.0005
R94 source.n15 source.t18 10.0005
R95 source.n15 source.t22 10.0005
R96 source.n13 source.t20 10.0005
R97 source.n13 source.t19 10.0005
R98 source.n1 source.t16 10.0005
R99 source.n1 source.t12 10.0005
R100 source.n3 source.t13 10.0005
R101 source.n3 source.t15 10.0005
R102 source.n7 source.t3 10.0005
R103 source.n7 source.t10 10.0005
R104 source.n9 source.t5 10.0005
R105 source.n9 source.t7 10.0005
R106 source.n24 source.n0 9.48679
R107 source.n24 source.n23 5.5436
R108 source.n11 source.n10 0.560845
R109 source.n10 source.n8 0.560845
R110 source.n8 source.n6 0.560845
R111 source.n5 source.n4 0.560845
R112 source.n4 source.n2 0.560845
R113 source.n2 source.n0 0.560845
R114 source.n14 source.n12 0.560845
R115 source.n16 source.n14 0.560845
R116 source.n17 source.n16 0.560845
R117 source.n20 source.n18 0.560845
R118 source.n22 source.n20 0.560845
R119 source.n23 source.n22 0.560845
R120 source.n6 source.n5 0.470328
R121 source.n18 source.n17 0.470328
R122 source source.n24 0.188
R123 minus.n13 minus.t9 745.639
R124 minus.n2 minus.t5 745.639
R125 minus.n28 minus.t1 745.639
R126 minus.n17 minus.t3 745.639
R127 minus.n12 minus.t6 690.867
R128 minus.n10 minus.t7 690.867
R129 minus.n3 minus.t8 690.867
R130 minus.n4 minus.t4 690.867
R131 minus.n27 minus.t2 690.867
R132 minus.n25 minus.t10 690.867
R133 minus.n19 minus.t11 690.867
R134 minus.n18 minus.t0 690.867
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 62.0763
R150 minus.n5 minus.n3 62.0763
R151 minus.n20 minus.n19 62.0763
R152 minus.n26 minus.n25 62.0763
R153 minus.n13 minus.n12 40.1672
R154 minus.n4 minus.n2 40.1672
R155 minus.n18 minus.n17 40.1672
R156 minus.n28 minus.n27 40.1672
R157 minus.n12 minus.n11 32.8641
R158 minus.n5 minus.n4 32.8641
R159 minus.n20 minus.n18 32.8641
R160 minus.n27 minus.n26 32.8641
R161 minus.n30 minus.n14 28.5043
R162 minus.n10 minus.n9 10.955
R163 minus.n3 minus.n1 10.955
R164 minus.n19 minus.n16 10.955
R165 minus.n25 minus.n24 10.955
R166 minus.n30 minus.n29 6.54217
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 80.3335
R177 drain_right.n3 drain_right.n2 80.278
R178 drain_right.n3 drain_right.n0 80.278
R179 drain_right.n6 drain_right.n5 79.7731
R180 drain_right.n8 drain_right.n7 79.7731
R181 drain_right.n3 drain_right.n1 79.773
R182 drain_right drain_right.n3 22.7974
R183 drain_right.n1 drain_right.t0 10.0005
R184 drain_right.n1 drain_right.t1 10.0005
R185 drain_right.n2 drain_right.t9 10.0005
R186 drain_right.n2 drain_right.t10 10.0005
R187 drain_right.n0 drain_right.t8 10.0005
R188 drain_right.n0 drain_right.t11 10.0005
R189 drain_right.n4 drain_right.t7 10.0005
R190 drain_right.n4 drain_right.t6 10.0005
R191 drain_right.n5 drain_right.t4 10.0005
R192 drain_right.n5 drain_right.t3 10.0005
R193 drain_right.n7 drain_right.t2 10.0005
R194 drain_right.n7 drain_right.t5 10.0005
R195 drain_right drain_right.n8 6.21356
R196 drain_right.n8 drain_right.n6 0.560845
C0 plus drain_right 0.315308f
C1 source drain_left 7.77537f
C2 minus plus 3.5038f
C3 source drain_right 7.77525f
C4 source minus 1.02614f
C5 source plus 1.04014f
C6 drain_right drain_left 0.801552f
C7 minus drain_left 0.175622f
C8 plus drain_left 1.19877f
C9 minus drain_right 1.04229f
C10 drain_right a_n1626_n1488# 3.69947f
C11 drain_left a_n1626_n1488# 3.92132f
C12 source a_n1626_n1488# 3.638657f
C13 minus a_n1626_n1488# 5.264042f
C14 plus a_n1626_n1488# 6.075041f
C15 drain_right.t8 a_n1626_n1488# 0.08759f
C16 drain_right.t11 a_n1626_n1488# 0.08759f
C17 drain_right.n0 a_n1626_n1488# 0.478297f
C18 drain_right.t0 a_n1626_n1488# 0.08759f
C19 drain_right.t1 a_n1626_n1488# 0.08759f
C20 drain_right.n1 a_n1626_n1488# 0.476474f
C21 drain_right.t9 a_n1626_n1488# 0.08759f
C22 drain_right.t10 a_n1626_n1488# 0.08759f
C23 drain_right.n2 a_n1626_n1488# 0.478297f
C24 drain_right.n3 a_n1626_n1488# 1.45545f
C25 drain_right.t7 a_n1626_n1488# 0.08759f
C26 drain_right.t6 a_n1626_n1488# 0.08759f
C27 drain_right.n4 a_n1626_n1488# 0.47852f
C28 drain_right.t4 a_n1626_n1488# 0.08759f
C29 drain_right.t3 a_n1626_n1488# 0.08759f
C30 drain_right.n5 a_n1626_n1488# 0.476476f
C31 drain_right.n6 a_n1626_n1488# 0.574282f
C32 drain_right.t2 a_n1626_n1488# 0.08759f
C33 drain_right.t5 a_n1626_n1488# 0.08759f
C34 drain_right.n7 a_n1626_n1488# 0.476476f
C35 drain_right.n8 a_n1626_n1488# 0.486892f
C36 minus.n0 a_n1626_n1488# 0.034114f
C37 minus.t9 a_n1626_n1488# 0.046776f
C38 minus.t6 a_n1626_n1488# 0.044455f
C39 minus.t7 a_n1626_n1488# 0.044455f
C40 minus.n1 a_n1626_n1488# 0.012894f
C41 minus.t5 a_n1626_n1488# 0.046776f
C42 minus.n2 a_n1626_n1488# 0.043797f
C43 minus.t8 a_n1626_n1488# 0.044455f
C44 minus.n3 a_n1626_n1488# 0.031071f
C45 minus.t4 a_n1626_n1488# 0.044455f
C46 minus.n4 a_n1626_n1488# 0.031071f
C47 minus.n5 a_n1626_n1488# 0.014472f
C48 minus.n6 a_n1626_n1488# 0.076591f
C49 minus.n7 a_n1626_n1488# 0.034114f
C50 minus.n8 a_n1626_n1488# 0.034114f
C51 minus.n9 a_n1626_n1488# 0.012894f
C52 minus.n10 a_n1626_n1488# 0.031071f
C53 minus.n11 a_n1626_n1488# 0.014472f
C54 minus.n12 a_n1626_n1488# 0.031071f
C55 minus.n13 a_n1626_n1488# 0.043747f
C56 minus.n14 a_n1626_n1488# 0.813693f
C57 minus.n15 a_n1626_n1488# 0.034114f
C58 minus.t2 a_n1626_n1488# 0.044455f
C59 minus.t10 a_n1626_n1488# 0.044455f
C60 minus.n16 a_n1626_n1488# 0.012894f
C61 minus.t3 a_n1626_n1488# 0.046776f
C62 minus.n17 a_n1626_n1488# 0.043797f
C63 minus.t0 a_n1626_n1488# 0.044455f
C64 minus.n18 a_n1626_n1488# 0.031071f
C65 minus.t11 a_n1626_n1488# 0.044455f
C66 minus.n19 a_n1626_n1488# 0.031071f
C67 minus.n20 a_n1626_n1488# 0.014472f
C68 minus.n21 a_n1626_n1488# 0.076591f
C69 minus.n22 a_n1626_n1488# 0.034114f
C70 minus.n23 a_n1626_n1488# 0.034114f
C71 minus.n24 a_n1626_n1488# 0.012894f
C72 minus.n25 a_n1626_n1488# 0.031071f
C73 minus.n26 a_n1626_n1488# 0.014472f
C74 minus.n27 a_n1626_n1488# 0.031071f
C75 minus.t1 a_n1626_n1488# 0.046776f
C76 minus.n28 a_n1626_n1488# 0.043747f
C77 minus.n29 a_n1626_n1488# 0.226409f
C78 minus.n30 a_n1626_n1488# 1.00377f
C79 source.t14 a_n1626_n1488# 0.485194f
C80 source.n0 a_n1626_n1488# 0.640518f
C81 source.t16 a_n1626_n1488# 0.082379f
C82 source.t12 a_n1626_n1488# 0.082379f
C83 source.n1 a_n1626_n1488# 0.400756f
C84 source.n2 a_n1626_n1488# 0.282606f
C85 source.t13 a_n1626_n1488# 0.082379f
C86 source.t15 a_n1626_n1488# 0.082379f
C87 source.n3 a_n1626_n1488# 0.400756f
C88 source.n4 a_n1626_n1488# 0.282606f
C89 source.t17 a_n1626_n1488# 0.485194f
C90 source.n5 a_n1626_n1488# 0.33976f
C91 source.t1 a_n1626_n1488# 0.485194f
C92 source.n6 a_n1626_n1488# 0.33976f
C93 source.t3 a_n1626_n1488# 0.082379f
C94 source.t10 a_n1626_n1488# 0.082379f
C95 source.n7 a_n1626_n1488# 0.400756f
C96 source.n8 a_n1626_n1488# 0.282606f
C97 source.t5 a_n1626_n1488# 0.082379f
C98 source.t7 a_n1626_n1488# 0.082379f
C99 source.n9 a_n1626_n1488# 0.400756f
C100 source.n10 a_n1626_n1488# 0.282606f
C101 source.t6 a_n1626_n1488# 0.485194f
C102 source.n11 a_n1626_n1488# 0.879881f
C103 source.t23 a_n1626_n1488# 0.485192f
C104 source.n12 a_n1626_n1488# 0.879884f
C105 source.t20 a_n1626_n1488# 0.082379f
C106 source.t19 a_n1626_n1488# 0.082379f
C107 source.n13 a_n1626_n1488# 0.400753f
C108 source.n14 a_n1626_n1488# 0.282608f
C109 source.t18 a_n1626_n1488# 0.082379f
C110 source.t22 a_n1626_n1488# 0.082379f
C111 source.n15 a_n1626_n1488# 0.400753f
C112 source.n16 a_n1626_n1488# 0.282608f
C113 source.t21 a_n1626_n1488# 0.485192f
C114 source.n17 a_n1626_n1488# 0.339763f
C115 source.t0 a_n1626_n1488# 0.485192f
C116 source.n18 a_n1626_n1488# 0.339763f
C117 source.t9 a_n1626_n1488# 0.082379f
C118 source.t2 a_n1626_n1488# 0.082379f
C119 source.n19 a_n1626_n1488# 0.400753f
C120 source.n20 a_n1626_n1488# 0.282608f
C121 source.t11 a_n1626_n1488# 0.082379f
C122 source.t8 a_n1626_n1488# 0.082379f
C123 source.n21 a_n1626_n1488# 0.400753f
C124 source.n22 a_n1626_n1488# 0.282608f
C125 source.t4 a_n1626_n1488# 0.485192f
C126 source.n23 a_n1626_n1488# 0.470245f
C127 source.n24 a_n1626_n1488# 0.665316f
C128 drain_left.t9 a_n1626_n1488# 0.086531f
C129 drain_left.t10 a_n1626_n1488# 0.086531f
C130 drain_left.n0 a_n1626_n1488# 0.472519f
C131 drain_left.t7 a_n1626_n1488# 0.086531f
C132 drain_left.t0 a_n1626_n1488# 0.086531f
C133 drain_left.n1 a_n1626_n1488# 0.470717f
C134 drain_left.t11 a_n1626_n1488# 0.086531f
C135 drain_left.t6 a_n1626_n1488# 0.086531f
C136 drain_left.n2 a_n1626_n1488# 0.472519f
C137 drain_left.n3 a_n1626_n1488# 1.48573f
C138 drain_left.t5 a_n1626_n1488# 0.086531f
C139 drain_left.t3 a_n1626_n1488# 0.086531f
C140 drain_left.n4 a_n1626_n1488# 0.472739f
C141 drain_left.t8 a_n1626_n1488# 0.086531f
C142 drain_left.t1 a_n1626_n1488# 0.086531f
C143 drain_left.n5 a_n1626_n1488# 0.470719f
C144 drain_left.n6 a_n1626_n1488# 0.567343f
C145 drain_left.t4 a_n1626_n1488# 0.086531f
C146 drain_left.t2 a_n1626_n1488# 0.086531f
C147 drain_left.n7 a_n1626_n1488# 0.470719f
C148 drain_left.n8 a_n1626_n1488# 0.481009f
C149 plus.n0 a_n1626_n1488# 0.0348f
C150 plus.t11 a_n1626_n1488# 0.045349f
C151 plus.t7 a_n1626_n1488# 0.045349f
C152 plus.n1 a_n1626_n1488# 0.013153f
C153 plus.t6 a_n1626_n1488# 0.047717f
C154 plus.n2 a_n1626_n1488# 0.044678f
C155 plus.t10 a_n1626_n1488# 0.045349f
C156 plus.n3 a_n1626_n1488# 0.031696f
C157 plus.t8 a_n1626_n1488# 0.045349f
C158 plus.n4 a_n1626_n1488# 0.031696f
C159 plus.n5 a_n1626_n1488# 0.014763f
C160 plus.n6 a_n1626_n1488# 0.078131f
C161 plus.n7 a_n1626_n1488# 0.0348f
C162 plus.n8 a_n1626_n1488# 0.0348f
C163 plus.n9 a_n1626_n1488# 0.013153f
C164 plus.n10 a_n1626_n1488# 0.031696f
C165 plus.n11 a_n1626_n1488# 0.014763f
C166 plus.n12 a_n1626_n1488# 0.031696f
C167 plus.t9 a_n1626_n1488# 0.047717f
C168 plus.n13 a_n1626_n1488# 0.044627f
C169 plus.n14 a_n1626_n1488# 0.263582f
C170 plus.n15 a_n1626_n1488# 0.0348f
C171 plus.t0 a_n1626_n1488# 0.047717f
C172 plus.t3 a_n1626_n1488# 0.045349f
C173 plus.t4 a_n1626_n1488# 0.045349f
C174 plus.n16 a_n1626_n1488# 0.013153f
C175 plus.t2 a_n1626_n1488# 0.047717f
C176 plus.n17 a_n1626_n1488# 0.044678f
C177 plus.t5 a_n1626_n1488# 0.045349f
C178 plus.n18 a_n1626_n1488# 0.031696f
C179 plus.t1 a_n1626_n1488# 0.045349f
C180 plus.n19 a_n1626_n1488# 0.031696f
C181 plus.n20 a_n1626_n1488# 0.014763f
C182 plus.n21 a_n1626_n1488# 0.078131f
C183 plus.n22 a_n1626_n1488# 0.0348f
C184 plus.n23 a_n1626_n1488# 0.0348f
C185 plus.n24 a_n1626_n1488# 0.013153f
C186 plus.n25 a_n1626_n1488# 0.031696f
C187 plus.n26 a_n1626_n1488# 0.014763f
C188 plus.n27 a_n1626_n1488# 0.031696f
C189 plus.n28 a_n1626_n1488# 0.044627f
C190 plus.n29 a_n1626_n1488# 0.782191f
.ends

