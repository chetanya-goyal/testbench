* NGSPICE file created from diffpair241.ext - technology: sky130A

.subckt diffpair241 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t4 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X1 source.t1 plus.t0 drain_left.t3 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X2 source.t7 minus.t1 drain_right.t2 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X3 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X4 drain_left.t2 plus.t1 source.t2 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X5 drain_left.t1 plus.t2 source.t3 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X6 drain_right.t1 minus.t2 source.t5 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X7 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X8 source.t0 plus.t3 drain_left.t0 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X9 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X10 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X11 source.t6 minus.t3 drain_right.t0 a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
R0 minus.n0 minus.t3 1220.34
R1 minus.n0 minus.t0 1220.34
R2 minus.n1 minus.t2 1220.34
R3 minus.n1 minus.t1 1220.34
R4 minus.n2 minus.n0 190.103
R5 minus.n2 minus.n1 167.823
R6 minus minus.n2 0.188
R7 source.n1 source.t1 55.512
R8 source.n2 source.t4 55.512
R9 source.n3 source.t6 55.512
R10 source.n0 source.t2 55.5119
R11 source.n7 source.t5 55.5119
R12 source.n6 source.t7 55.5119
R13 source.n5 source.t3 55.5119
R14 source.n4 source.t0 55.5119
R15 source.n4 source.n3 17.3178
R16 source.n8 source.n0 11.7747
R17 source.n8 source.n7 5.5436
R18 source.n3 source.n2 0.560845
R19 source.n1 source.n0 0.560845
R20 source.n5 source.n4 0.560845
R21 source.n7 source.n6 0.560845
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 90.5944
R26 drain_right drain_right.n1 73.4037
R27 drain_right.n0 drain_right.t2 5.0005
R28 drain_right.n0 drain_right.t1 5.0005
R29 drain_right.n1 drain_right.t0 5.0005
R30 drain_right.n1 drain_right.t3 5.0005
R31 plus.n0 plus.t0 1220.34
R32 plus.n0 plus.t1 1220.34
R33 plus.n1 plus.t2 1220.34
R34 plus.n1 plus.t3 1220.34
R35 plus plus.n1 186.257
R36 plus plus.n0 171.195
R37 drain_left drain_left.n0 91.1476
R38 drain_left drain_left.n1 73.4037
R39 drain_left.n0 drain_left.t0 5.0005
R40 drain_left.n0 drain_left.t1 5.0005
R41 drain_left.n1 drain_left.t3 5.0005
R42 drain_left.n1 drain_left.t2 5.0005
C0 source minus 0.607949f
C1 plus drain_left 0.9905f
C2 plus drain_right 0.256158f
C3 plus source 0.621967f
C4 plus minus 3.39939f
C5 drain_left drain_right 0.481587f
C6 drain_left source 5.55265f
C7 drain_left minus 0.171192f
C8 source drain_right 5.55131f
C9 minus drain_right 0.888201f
C10 drain_right a_n1106_n2092# 4.49788f
C11 drain_left a_n1106_n2092# 4.6417f
C12 source a_n1106_n2092# 5.129342f
C13 minus a_n1106_n2092# 3.574673f
C14 plus a_n1106_n2092# 5.93346f
C15 drain_left.t0 a_n1106_n2092# 0.170029f
C16 drain_left.t1 a_n1106_n2092# 0.170029f
C17 drain_left.n0 a_n1106_n2092# 1.25457f
C18 drain_left.t3 a_n1106_n2092# 0.170029f
C19 drain_left.t2 a_n1106_n2092# 0.170029f
C20 drain_left.n1 a_n1106_n2092# 1.09256f
C21 plus.t0 a_n1106_n2092# 0.116701f
C22 plus.t1 a_n1106_n2092# 0.116701f
C23 plus.n0 a_n1106_n2092# 0.154501f
C24 plus.t3 a_n1106_n2092# 0.116701f
C25 plus.t2 a_n1106_n2092# 0.116701f
C26 plus.n1 a_n1106_n2092# 0.264395f
C27 drain_right.t2 a_n1106_n2092# 0.172888f
C28 drain_right.t1 a_n1106_n2092# 0.172888f
C29 drain_right.n0 a_n1106_n2092# 1.25934f
C30 drain_right.t0 a_n1106_n2092# 0.172888f
C31 drain_right.t3 a_n1106_n2092# 0.172888f
C32 drain_right.n1 a_n1106_n2092# 1.11093f
C33 source.t2 a_n1106_n2092# 0.838145f
C34 source.n0 a_n1106_n2092# 0.617435f
C35 source.t1 a_n1106_n2092# 0.838149f
C36 source.n1 a_n1106_n2092# 0.282f
C37 source.t4 a_n1106_n2092# 0.838149f
C38 source.n2 a_n1106_n2092# 0.282f
C39 source.t6 a_n1106_n2092# 0.838149f
C40 source.n3 a_n1106_n2092# 0.831757f
C41 source.t0 a_n1106_n2092# 0.838145f
C42 source.n4 a_n1106_n2092# 0.831761f
C43 source.t3 a_n1106_n2092# 0.838145f
C44 source.n5 a_n1106_n2092# 0.282004f
C45 source.t7 a_n1106_n2092# 0.838145f
C46 source.n6 a_n1106_n2092# 0.282004f
C47 source.t5 a_n1106_n2092# 0.838145f
C48 source.n7 a_n1106_n2092# 0.376508f
C49 source.n8 a_n1106_n2092# 0.681394f
C50 minus.t3 a_n1106_n2092# 0.113684f
C51 minus.t0 a_n1106_n2092# 0.113684f
C52 minus.n0 a_n1106_n2092# 0.289395f
C53 minus.t1 a_n1106_n2092# 0.113684f
C54 minus.t2 a_n1106_n2092# 0.113684f
C55 minus.n1 a_n1106_n2092# 0.139823f
C56 minus.n2 a_n1106_n2092# 2.4875f
.ends

