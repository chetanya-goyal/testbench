* NGSPICE file created from diffpair339.ext - technology: sky130A

.subckt diffpair339 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t14 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 source.t46 minus.t1 drain_right.t6 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 drain_right.t23 minus.t2 source.t45 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X3 drain_right.t22 minus.t3 source.t44 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 source.t17 plus.t0 drain_left.t23 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 drain_right.t21 minus.t4 source.t43 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X6 drain_right.t13 minus.t5 source.t42 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X7 drain_right.t5 minus.t6 source.t41 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X8 drain_right.t0 minus.t7 source.t40 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X9 drain_right.t3 minus.t8 source.t39 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X10 a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X11 source.t38 minus.t9 drain_right.t2 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X12 drain_right.t12 minus.t10 source.t37 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X13 source.t16 plus.t1 drain_left.t22 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X14 drain_left.t21 plus.t2 source.t22 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X15 source.t36 minus.t11 drain_right.t1 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X16 source.t35 minus.t12 drain_right.t11 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X17 source.t20 plus.t3 drain_left.t20 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X18 source.t34 minus.t13 drain_right.t4 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X19 source.t33 minus.t14 drain_right.t10 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X20 drain_left.t19 plus.t4 source.t19 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X21 source.t32 minus.t15 drain_right.t20 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X22 drain_left.t18 plus.t5 source.t15 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X23 a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X24 source.t31 minus.t16 drain_right.t18 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X25 drain_right.t9 minus.t17 source.t30 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X26 drain_left.t17 plus.t6 source.t1 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X27 source.t2 plus.t7 drain_left.t16 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X28 a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X29 drain_left.t15 plus.t8 source.t6 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X30 source.t10 plus.t9 drain_left.t14 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X31 source.t12 plus.t10 drain_left.t13 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X32 source.t18 plus.t11 drain_left.t12 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X33 drain_right.t8 minus.t18 source.t29 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X34 source.t0 plus.t12 drain_left.t11 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X35 drain_right.t15 minus.t19 source.t28 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X36 drain_right.t16 minus.t20 source.t27 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X37 drain_left.t10 plus.t13 source.t13 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X38 drain_left.t9 plus.t14 source.t21 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X39 source.t23 plus.t15 drain_left.t8 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X40 drain_left.t7 plus.t16 source.t14 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X41 drain_left.t6 plus.t17 source.t3 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X42 source.t5 plus.t18 drain_left.t5 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X43 drain_left.t4 plus.t19 source.t7 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X44 source.t11 plus.t20 drain_left.t3 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X45 source.t26 minus.t21 drain_right.t17 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X46 source.t25 minus.t22 drain_right.t19 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X47 a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X48 drain_left.t2 plus.t21 source.t8 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X49 drain_left.t1 plus.t22 source.t4 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X50 source.t9 plus.t23 drain_left.t0 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X51 source.t24 minus.t23 drain_right.t7 a_n2094_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n29 minus.t9 1301.77
R1 minus.n6 minus.t19 1301.77
R2 minus.n60 minus.t2 1301.77
R3 minus.n37 minus.t1 1301.77
R4 minus.n28 minus.t17 1241.15
R5 minus.n26 minus.t16 1241.15
R6 minus.n1 minus.t18 1241.15
R7 minus.n21 minus.t22 1241.15
R8 minus.n19 minus.t5 1241.15
R9 minus.n3 minus.t14 1241.15
R10 minus.n14 minus.t20 1241.15
R11 minus.n12 minus.t21 1241.15
R12 minus.n5 minus.t4 1241.15
R13 minus.n7 minus.t15 1241.15
R14 minus.n59 minus.t23 1241.15
R15 minus.n57 minus.t3 1241.15
R16 minus.n32 minus.t11 1241.15
R17 minus.n52 minus.t8 1241.15
R18 minus.n50 minus.t12 1241.15
R19 minus.n34 minus.t10 1241.15
R20 minus.n45 minus.t13 1241.15
R21 minus.n43 minus.t6 1241.15
R22 minus.n36 minus.t0 1241.15
R23 minus.n38 minus.t7 1241.15
R24 minus.n9 minus.n6 161.489
R25 minus.n40 minus.n37 161.489
R26 minus.n30 minus.n29 161.3
R27 minus.n27 minus.n0 161.3
R28 minus.n25 minus.n24 161.3
R29 minus.n23 minus.n22 161.3
R30 minus.n20 minus.n2 161.3
R31 minus.n18 minus.n17 161.3
R32 minus.n16 minus.n15 161.3
R33 minus.n13 minus.n4 161.3
R34 minus.n11 minus.n10 161.3
R35 minus.n9 minus.n8 161.3
R36 minus.n61 minus.n60 161.3
R37 minus.n58 minus.n31 161.3
R38 minus.n56 minus.n55 161.3
R39 minus.n54 minus.n53 161.3
R40 minus.n51 minus.n33 161.3
R41 minus.n49 minus.n48 161.3
R42 minus.n47 minus.n46 161.3
R43 minus.n44 minus.n35 161.3
R44 minus.n42 minus.n41 161.3
R45 minus.n40 minus.n39 161.3
R46 minus.n28 minus.n27 56.2338
R47 minus.n8 minus.n7 56.2338
R48 minus.n39 minus.n38 56.2338
R49 minus.n59 minus.n58 56.2338
R50 minus.n26 minus.n25 51.852
R51 minus.n11 minus.n5 51.852
R52 minus.n42 minus.n36 51.852
R53 minus.n57 minus.n56 51.852
R54 minus.n22 minus.n1 47.4702
R55 minus.n13 minus.n12 47.4702
R56 minus.n44 minus.n43 47.4702
R57 minus.n53 minus.n32 47.4702
R58 minus.n21 minus.n20 43.0884
R59 minus.n15 minus.n14 43.0884
R60 minus.n46 minus.n45 43.0884
R61 minus.n52 minus.n51 43.0884
R62 minus.n19 minus.n18 38.7066
R63 minus.n18 minus.n3 38.7066
R64 minus.n49 minus.n34 38.7066
R65 minus.n50 minus.n49 38.7066
R66 minus.n62 minus.n30 34.7694
R67 minus.n20 minus.n19 34.3247
R68 minus.n15 minus.n3 34.3247
R69 minus.n46 minus.n34 34.3247
R70 minus.n51 minus.n50 34.3247
R71 minus.n22 minus.n21 29.9429
R72 minus.n14 minus.n13 29.9429
R73 minus.n45 minus.n44 29.9429
R74 minus.n53 minus.n52 29.9429
R75 minus.n25 minus.n1 25.5611
R76 minus.n12 minus.n11 25.5611
R77 minus.n43 minus.n42 25.5611
R78 minus.n56 minus.n32 25.5611
R79 minus.n27 minus.n26 21.1793
R80 minus.n8 minus.n5 21.1793
R81 minus.n39 minus.n36 21.1793
R82 minus.n58 minus.n57 21.1793
R83 minus.n29 minus.n28 16.7975
R84 minus.n7 minus.n6 16.7975
R85 minus.n38 minus.n37 16.7975
R86 minus.n60 minus.n59 16.7975
R87 minus.n62 minus.n61 6.48914
R88 minus.n30 minus.n0 0.189894
R89 minus.n24 minus.n0 0.189894
R90 minus.n24 minus.n23 0.189894
R91 minus.n23 minus.n2 0.189894
R92 minus.n17 minus.n2 0.189894
R93 minus.n17 minus.n16 0.189894
R94 minus.n16 minus.n4 0.189894
R95 minus.n10 minus.n4 0.189894
R96 minus.n10 minus.n9 0.189894
R97 minus.n41 minus.n40 0.189894
R98 minus.n41 minus.n35 0.189894
R99 minus.n47 minus.n35 0.189894
R100 minus.n48 minus.n47 0.189894
R101 minus.n48 minus.n33 0.189894
R102 minus.n54 minus.n33 0.189894
R103 minus.n55 minus.n54 0.189894
R104 minus.n55 minus.n31 0.189894
R105 minus.n61 minus.n31 0.189894
R106 minus minus.n62 0.188
R107 drain_right.n13 drain_right.n11 65.9943
R108 drain_right.n7 drain_right.n5 65.9942
R109 drain_right.n2 drain_right.n0 65.9942
R110 drain_right.n13 drain_right.n12 65.5376
R111 drain_right.n15 drain_right.n14 65.5376
R112 drain_right.n17 drain_right.n16 65.5376
R113 drain_right.n19 drain_right.n18 65.5376
R114 drain_right.n21 drain_right.n20 65.5376
R115 drain_right.n7 drain_right.n6 65.5373
R116 drain_right.n9 drain_right.n8 65.5373
R117 drain_right.n4 drain_right.n3 65.5373
R118 drain_right.n2 drain_right.n1 65.5373
R119 drain_right drain_right.n10 28.8816
R120 drain_right drain_right.n21 6.11011
R121 drain_right.n5 drain_right.t7 2.2005
R122 drain_right.n5 drain_right.t23 2.2005
R123 drain_right.n6 drain_right.t1 2.2005
R124 drain_right.n6 drain_right.t22 2.2005
R125 drain_right.n8 drain_right.t11 2.2005
R126 drain_right.n8 drain_right.t3 2.2005
R127 drain_right.n3 drain_right.t4 2.2005
R128 drain_right.n3 drain_right.t12 2.2005
R129 drain_right.n1 drain_right.t14 2.2005
R130 drain_right.n1 drain_right.t5 2.2005
R131 drain_right.n0 drain_right.t6 2.2005
R132 drain_right.n0 drain_right.t0 2.2005
R133 drain_right.n11 drain_right.t20 2.2005
R134 drain_right.n11 drain_right.t15 2.2005
R135 drain_right.n12 drain_right.t17 2.2005
R136 drain_right.n12 drain_right.t21 2.2005
R137 drain_right.n14 drain_right.t10 2.2005
R138 drain_right.n14 drain_right.t16 2.2005
R139 drain_right.n16 drain_right.t19 2.2005
R140 drain_right.n16 drain_right.t13 2.2005
R141 drain_right.n18 drain_right.t18 2.2005
R142 drain_right.n18 drain_right.t8 2.2005
R143 drain_right.n20 drain_right.t2 2.2005
R144 drain_right.n20 drain_right.t9 2.2005
R145 drain_right.n9 drain_right.n7 0.457397
R146 drain_right.n4 drain_right.n2 0.457397
R147 drain_right.n21 drain_right.n19 0.457397
R148 drain_right.n19 drain_right.n17 0.457397
R149 drain_right.n17 drain_right.n15 0.457397
R150 drain_right.n15 drain_right.n13 0.457397
R151 drain_right.n10 drain_right.n9 0.173602
R152 drain_right.n10 drain_right.n4 0.173602
R153 source.n11 source.t2 51.0588
R154 source.n12 source.t28 51.0588
R155 source.n23 source.t38 51.0588
R156 source.n47 source.t45 51.0586
R157 source.n36 source.t46 51.0586
R158 source.n35 source.t14 51.0586
R159 source.n24 source.t0 51.0586
R160 source.n0 source.t8 51.0586
R161 source.n2 source.n1 48.8588
R162 source.n4 source.n3 48.8588
R163 source.n6 source.n5 48.8588
R164 source.n8 source.n7 48.8588
R165 source.n10 source.n9 48.8588
R166 source.n14 source.n13 48.8588
R167 source.n16 source.n15 48.8588
R168 source.n18 source.n17 48.8588
R169 source.n20 source.n19 48.8588
R170 source.n22 source.n21 48.8588
R171 source.n46 source.n45 48.8586
R172 source.n44 source.n43 48.8586
R173 source.n42 source.n41 48.8586
R174 source.n40 source.n39 48.8586
R175 source.n38 source.n37 48.8586
R176 source.n34 source.n33 48.8586
R177 source.n32 source.n31 48.8586
R178 source.n30 source.n29 48.8586
R179 source.n28 source.n27 48.8586
R180 source.n26 source.n25 48.8586
R181 source.n24 source.n23 19.4719
R182 source.n48 source.n0 13.9805
R183 source.n48 source.n47 5.49188
R184 source.n45 source.t44 2.2005
R185 source.n45 source.t24 2.2005
R186 source.n43 source.t39 2.2005
R187 source.n43 source.t36 2.2005
R188 source.n41 source.t37 2.2005
R189 source.n41 source.t35 2.2005
R190 source.n39 source.t41 2.2005
R191 source.n39 source.t34 2.2005
R192 source.n37 source.t40 2.2005
R193 source.n37 source.t47 2.2005
R194 source.n33 source.t3 2.2005
R195 source.n33 source.t11 2.2005
R196 source.n31 source.t21 2.2005
R197 source.n31 source.t12 2.2005
R198 source.n29 source.t13 2.2005
R199 source.n29 source.t18 2.2005
R200 source.n27 source.t19 2.2005
R201 source.n27 source.t10 2.2005
R202 source.n25 source.t6 2.2005
R203 source.n25 source.t20 2.2005
R204 source.n1 source.t15 2.2005
R205 source.n1 source.t17 2.2005
R206 source.n3 source.t4 2.2005
R207 source.n3 source.t23 2.2005
R208 source.n5 source.t1 2.2005
R209 source.n5 source.t16 2.2005
R210 source.n7 source.t7 2.2005
R211 source.n7 source.t5 2.2005
R212 source.n9 source.t22 2.2005
R213 source.n9 source.t9 2.2005
R214 source.n13 source.t43 2.2005
R215 source.n13 source.t32 2.2005
R216 source.n15 source.t27 2.2005
R217 source.n15 source.t26 2.2005
R218 source.n17 source.t42 2.2005
R219 source.n17 source.t33 2.2005
R220 source.n19 source.t29 2.2005
R221 source.n19 source.t25 2.2005
R222 source.n21 source.t30 2.2005
R223 source.n21 source.t31 2.2005
R224 source.n12 source.n11 0.470328
R225 source.n36 source.n35 0.470328
R226 source.n23 source.n22 0.457397
R227 source.n22 source.n20 0.457397
R228 source.n20 source.n18 0.457397
R229 source.n18 source.n16 0.457397
R230 source.n16 source.n14 0.457397
R231 source.n14 source.n12 0.457397
R232 source.n11 source.n10 0.457397
R233 source.n10 source.n8 0.457397
R234 source.n8 source.n6 0.457397
R235 source.n6 source.n4 0.457397
R236 source.n4 source.n2 0.457397
R237 source.n2 source.n0 0.457397
R238 source.n26 source.n24 0.457397
R239 source.n28 source.n26 0.457397
R240 source.n30 source.n28 0.457397
R241 source.n32 source.n30 0.457397
R242 source.n34 source.n32 0.457397
R243 source.n35 source.n34 0.457397
R244 source.n38 source.n36 0.457397
R245 source.n40 source.n38 0.457397
R246 source.n42 source.n40 0.457397
R247 source.n44 source.n42 0.457397
R248 source.n46 source.n44 0.457397
R249 source.n47 source.n46 0.457397
R250 source source.n48 0.188
R251 plus.n6 plus.t7 1301.77
R252 plus.n29 plus.t21 1301.77
R253 plus.n37 plus.t16 1301.77
R254 plus.n60 plus.t12 1301.77
R255 plus.n7 plus.t2 1241.15
R256 plus.n5 plus.t23 1241.15
R257 plus.n12 plus.t19 1241.15
R258 plus.n14 plus.t18 1241.15
R259 plus.n3 plus.t6 1241.15
R260 plus.n19 plus.t1 1241.15
R261 plus.n21 plus.t22 1241.15
R262 plus.n1 plus.t15 1241.15
R263 plus.n26 plus.t5 1241.15
R264 plus.n28 plus.t0 1241.15
R265 plus.n38 plus.t20 1241.15
R266 plus.n36 plus.t17 1241.15
R267 plus.n43 plus.t10 1241.15
R268 plus.n45 plus.t14 1241.15
R269 plus.n34 plus.t11 1241.15
R270 plus.n50 plus.t13 1241.15
R271 plus.n52 plus.t9 1241.15
R272 plus.n32 plus.t4 1241.15
R273 plus.n57 plus.t3 1241.15
R274 plus.n59 plus.t8 1241.15
R275 plus.n9 plus.n6 161.489
R276 plus.n40 plus.n37 161.489
R277 plus.n9 plus.n8 161.3
R278 plus.n11 plus.n10 161.3
R279 plus.n13 plus.n4 161.3
R280 plus.n16 plus.n15 161.3
R281 plus.n18 plus.n17 161.3
R282 plus.n20 plus.n2 161.3
R283 plus.n23 plus.n22 161.3
R284 plus.n25 plus.n24 161.3
R285 plus.n27 plus.n0 161.3
R286 plus.n30 plus.n29 161.3
R287 plus.n40 plus.n39 161.3
R288 plus.n42 plus.n41 161.3
R289 plus.n44 plus.n35 161.3
R290 plus.n47 plus.n46 161.3
R291 plus.n49 plus.n48 161.3
R292 plus.n51 plus.n33 161.3
R293 plus.n54 plus.n53 161.3
R294 plus.n56 plus.n55 161.3
R295 plus.n58 plus.n31 161.3
R296 plus.n61 plus.n60 161.3
R297 plus.n8 plus.n7 56.2338
R298 plus.n28 plus.n27 56.2338
R299 plus.n59 plus.n58 56.2338
R300 plus.n39 plus.n38 56.2338
R301 plus.n11 plus.n5 51.852
R302 plus.n26 plus.n25 51.852
R303 plus.n57 plus.n56 51.852
R304 plus.n42 plus.n36 51.852
R305 plus.n13 plus.n12 47.4702
R306 plus.n22 plus.n1 47.4702
R307 plus.n53 plus.n32 47.4702
R308 plus.n44 plus.n43 47.4702
R309 plus.n15 plus.n14 43.0884
R310 plus.n21 plus.n20 43.0884
R311 plus.n52 plus.n51 43.0884
R312 plus.n46 plus.n45 43.0884
R313 plus.n18 plus.n3 38.7066
R314 plus.n19 plus.n18 38.7066
R315 plus.n50 plus.n49 38.7066
R316 plus.n49 plus.n34 38.7066
R317 plus.n15 plus.n3 34.3247
R318 plus.n20 plus.n19 34.3247
R319 plus.n51 plus.n50 34.3247
R320 plus.n46 plus.n34 34.3247
R321 plus.n14 plus.n13 29.9429
R322 plus.n22 plus.n21 29.9429
R323 plus.n53 plus.n52 29.9429
R324 plus.n45 plus.n44 29.9429
R325 plus plus.n61 29.7869
R326 plus.n12 plus.n11 25.5611
R327 plus.n25 plus.n1 25.5611
R328 plus.n56 plus.n32 25.5611
R329 plus.n43 plus.n42 25.5611
R330 plus.n8 plus.n5 21.1793
R331 plus.n27 plus.n26 21.1793
R332 plus.n58 plus.n57 21.1793
R333 plus.n39 plus.n36 21.1793
R334 plus.n7 plus.n6 16.7975
R335 plus.n29 plus.n28 16.7975
R336 plus.n60 plus.n59 16.7975
R337 plus.n38 plus.n37 16.7975
R338 plus plus.n30 10.9967
R339 plus.n10 plus.n9 0.189894
R340 plus.n10 plus.n4 0.189894
R341 plus.n16 plus.n4 0.189894
R342 plus.n17 plus.n16 0.189894
R343 plus.n17 plus.n2 0.189894
R344 plus.n23 plus.n2 0.189894
R345 plus.n24 plus.n23 0.189894
R346 plus.n24 plus.n0 0.189894
R347 plus.n30 plus.n0 0.189894
R348 plus.n61 plus.n31 0.189894
R349 plus.n55 plus.n31 0.189894
R350 plus.n55 plus.n54 0.189894
R351 plus.n54 plus.n33 0.189894
R352 plus.n48 plus.n33 0.189894
R353 plus.n48 plus.n47 0.189894
R354 plus.n47 plus.n35 0.189894
R355 plus.n41 plus.n35 0.189894
R356 plus.n41 plus.n40 0.189894
R357 drain_left.n13 drain_left.n11 65.9945
R358 drain_left.n7 drain_left.n5 65.9942
R359 drain_left.n2 drain_left.n0 65.9942
R360 drain_left.n19 drain_left.n18 65.5376
R361 drain_left.n17 drain_left.n16 65.5376
R362 drain_left.n15 drain_left.n14 65.5376
R363 drain_left.n13 drain_left.n12 65.5376
R364 drain_left.n21 drain_left.n20 65.5374
R365 drain_left.n7 drain_left.n6 65.5373
R366 drain_left.n9 drain_left.n8 65.5373
R367 drain_left.n4 drain_left.n3 65.5373
R368 drain_left.n2 drain_left.n1 65.5373
R369 drain_left drain_left.n10 29.4349
R370 drain_left drain_left.n21 6.11011
R371 drain_left.n5 drain_left.t3 2.2005
R372 drain_left.n5 drain_left.t7 2.2005
R373 drain_left.n6 drain_left.t13 2.2005
R374 drain_left.n6 drain_left.t6 2.2005
R375 drain_left.n8 drain_left.t12 2.2005
R376 drain_left.n8 drain_left.t9 2.2005
R377 drain_left.n3 drain_left.t14 2.2005
R378 drain_left.n3 drain_left.t10 2.2005
R379 drain_left.n1 drain_left.t20 2.2005
R380 drain_left.n1 drain_left.t19 2.2005
R381 drain_left.n0 drain_left.t11 2.2005
R382 drain_left.n0 drain_left.t15 2.2005
R383 drain_left.n20 drain_left.t23 2.2005
R384 drain_left.n20 drain_left.t2 2.2005
R385 drain_left.n18 drain_left.t8 2.2005
R386 drain_left.n18 drain_left.t18 2.2005
R387 drain_left.n16 drain_left.t22 2.2005
R388 drain_left.n16 drain_left.t1 2.2005
R389 drain_left.n14 drain_left.t5 2.2005
R390 drain_left.n14 drain_left.t17 2.2005
R391 drain_left.n12 drain_left.t0 2.2005
R392 drain_left.n12 drain_left.t4 2.2005
R393 drain_left.n11 drain_left.t16 2.2005
R394 drain_left.n11 drain_left.t21 2.2005
R395 drain_left.n9 drain_left.n7 0.457397
R396 drain_left.n4 drain_left.n2 0.457397
R397 drain_left.n15 drain_left.n13 0.457397
R398 drain_left.n17 drain_left.n15 0.457397
R399 drain_left.n19 drain_left.n17 0.457397
R400 drain_left.n21 drain_left.n19 0.457397
R401 drain_left.n10 drain_left.n9 0.173602
R402 drain_left.n10 drain_left.n4 0.173602
C0 source plus 4.64727f
C1 source drain_right 41.2093f
C2 minus drain_left 0.171754f
C3 plus minus 5.21056f
C4 minus drain_right 4.82475f
C5 plus drain_left 5.02989f
C6 drain_right drain_left 1.11966f
C7 plus drain_right 0.359911f
C8 source minus 4.63323f
C9 source drain_left 41.209f
C10 drain_right a_n2094_n2688# 6.75972f
C11 drain_left a_n2094_n2688# 7.08812f
C12 source a_n2094_n2688# 7.123847f
C13 minus a_n2094_n2688# 7.947259f
C14 plus a_n2094_n2688# 9.844861f
C15 drain_left.t11 a_n2094_n2688# 0.276142f
C16 drain_left.t15 a_n2094_n2688# 0.276142f
C17 drain_left.n0 a_n2094_n2688# 2.41838f
C18 drain_left.t20 a_n2094_n2688# 0.276142f
C19 drain_left.t19 a_n2094_n2688# 0.276142f
C20 drain_left.n1 a_n2094_n2688# 2.41532f
C21 drain_left.n2 a_n2094_n2688# 0.863257f
C22 drain_left.t14 a_n2094_n2688# 0.276142f
C23 drain_left.t10 a_n2094_n2688# 0.276142f
C24 drain_left.n3 a_n2094_n2688# 2.41532f
C25 drain_left.n4 a_n2094_n2688# 0.39503f
C26 drain_left.t3 a_n2094_n2688# 0.276142f
C27 drain_left.t7 a_n2094_n2688# 0.276142f
C28 drain_left.n5 a_n2094_n2688# 2.41838f
C29 drain_left.t13 a_n2094_n2688# 0.276142f
C30 drain_left.t6 a_n2094_n2688# 0.276142f
C31 drain_left.n6 a_n2094_n2688# 2.41532f
C32 drain_left.n7 a_n2094_n2688# 0.863257f
C33 drain_left.t12 a_n2094_n2688# 0.276142f
C34 drain_left.t9 a_n2094_n2688# 0.276142f
C35 drain_left.n8 a_n2094_n2688# 2.41532f
C36 drain_left.n9 a_n2094_n2688# 0.39503f
C37 drain_left.n10 a_n2094_n2688# 1.72855f
C38 drain_left.t16 a_n2094_n2688# 0.276142f
C39 drain_left.t21 a_n2094_n2688# 0.276142f
C40 drain_left.n11 a_n2094_n2688# 2.41838f
C41 drain_left.t0 a_n2094_n2688# 0.276142f
C42 drain_left.t4 a_n2094_n2688# 0.276142f
C43 drain_left.n12 a_n2094_n2688# 2.41533f
C44 drain_left.n13 a_n2094_n2688# 0.863247f
C45 drain_left.t5 a_n2094_n2688# 0.276142f
C46 drain_left.t17 a_n2094_n2688# 0.276142f
C47 drain_left.n14 a_n2094_n2688# 2.41533f
C48 drain_left.n15 a_n2094_n2688# 0.425331f
C49 drain_left.t22 a_n2094_n2688# 0.276142f
C50 drain_left.t1 a_n2094_n2688# 0.276142f
C51 drain_left.n16 a_n2094_n2688# 2.41533f
C52 drain_left.n17 a_n2094_n2688# 0.425331f
C53 drain_left.t8 a_n2094_n2688# 0.276142f
C54 drain_left.t18 a_n2094_n2688# 0.276142f
C55 drain_left.n18 a_n2094_n2688# 2.41533f
C56 drain_left.n19 a_n2094_n2688# 0.425331f
C57 drain_left.t23 a_n2094_n2688# 0.276142f
C58 drain_left.t2 a_n2094_n2688# 0.276142f
C59 drain_left.n20 a_n2094_n2688# 2.41532f
C60 drain_left.n21 a_n2094_n2688# 0.743105f
C61 plus.n0 a_n2094_n2688# 0.052222f
C62 plus.t0 a_n2094_n2688# 0.266356f
C63 plus.t5 a_n2094_n2688# 0.266356f
C64 plus.t15 a_n2094_n2688# 0.266356f
C65 plus.n1 a_n2094_n2688# 0.116592f
C66 plus.n2 a_n2094_n2688# 0.052222f
C67 plus.t22 a_n2094_n2688# 0.266356f
C68 plus.t1 a_n2094_n2688# 0.266356f
C69 plus.t6 a_n2094_n2688# 0.266356f
C70 plus.n3 a_n2094_n2688# 0.116592f
C71 plus.n4 a_n2094_n2688# 0.052222f
C72 plus.t18 a_n2094_n2688# 0.266356f
C73 plus.t19 a_n2094_n2688# 0.266356f
C74 plus.t23 a_n2094_n2688# 0.266356f
C75 plus.n5 a_n2094_n2688# 0.116592f
C76 plus.t7 a_n2094_n2688# 0.271957f
C77 plus.n6 a_n2094_n2688# 0.133064f
C78 plus.t2 a_n2094_n2688# 0.266356f
C79 plus.n7 a_n2094_n2688# 0.116592f
C80 plus.n8 a_n2094_n2688# 0.018289f
C81 plus.n9 a_n2094_n2688# 0.121426f
C82 plus.n10 a_n2094_n2688# 0.052222f
C83 plus.n11 a_n2094_n2688# 0.018289f
C84 plus.n12 a_n2094_n2688# 0.116592f
C85 plus.n13 a_n2094_n2688# 0.018289f
C86 plus.n14 a_n2094_n2688# 0.116592f
C87 plus.n15 a_n2094_n2688# 0.018289f
C88 plus.n16 a_n2094_n2688# 0.052222f
C89 plus.n17 a_n2094_n2688# 0.052222f
C90 plus.n18 a_n2094_n2688# 0.018289f
C91 plus.n19 a_n2094_n2688# 0.116592f
C92 plus.n20 a_n2094_n2688# 0.018289f
C93 plus.n21 a_n2094_n2688# 0.116592f
C94 plus.n22 a_n2094_n2688# 0.018289f
C95 plus.n23 a_n2094_n2688# 0.052222f
C96 plus.n24 a_n2094_n2688# 0.052222f
C97 plus.n25 a_n2094_n2688# 0.018289f
C98 plus.n26 a_n2094_n2688# 0.116592f
C99 plus.n27 a_n2094_n2688# 0.018289f
C100 plus.n28 a_n2094_n2688# 0.116592f
C101 plus.t21 a_n2094_n2688# 0.271957f
C102 plus.n29 a_n2094_n2688# 0.132982f
C103 plus.n30 a_n2094_n2688# 0.511595f
C104 plus.n31 a_n2094_n2688# 0.052222f
C105 plus.t12 a_n2094_n2688# 0.271957f
C106 plus.t8 a_n2094_n2688# 0.266356f
C107 plus.t3 a_n2094_n2688# 0.266356f
C108 plus.t4 a_n2094_n2688# 0.266356f
C109 plus.n32 a_n2094_n2688# 0.116592f
C110 plus.n33 a_n2094_n2688# 0.052222f
C111 plus.t9 a_n2094_n2688# 0.266356f
C112 plus.t13 a_n2094_n2688# 0.266356f
C113 plus.t11 a_n2094_n2688# 0.266356f
C114 plus.n34 a_n2094_n2688# 0.116592f
C115 plus.n35 a_n2094_n2688# 0.052222f
C116 plus.t14 a_n2094_n2688# 0.266356f
C117 plus.t10 a_n2094_n2688# 0.266356f
C118 plus.t17 a_n2094_n2688# 0.266356f
C119 plus.n36 a_n2094_n2688# 0.116592f
C120 plus.t16 a_n2094_n2688# 0.271957f
C121 plus.n37 a_n2094_n2688# 0.133064f
C122 plus.t20 a_n2094_n2688# 0.266356f
C123 plus.n38 a_n2094_n2688# 0.116592f
C124 plus.n39 a_n2094_n2688# 0.018289f
C125 plus.n40 a_n2094_n2688# 0.121426f
C126 plus.n41 a_n2094_n2688# 0.052222f
C127 plus.n42 a_n2094_n2688# 0.018289f
C128 plus.n43 a_n2094_n2688# 0.116592f
C129 plus.n44 a_n2094_n2688# 0.018289f
C130 plus.n45 a_n2094_n2688# 0.116592f
C131 plus.n46 a_n2094_n2688# 0.018289f
C132 plus.n47 a_n2094_n2688# 0.052222f
C133 plus.n48 a_n2094_n2688# 0.052222f
C134 plus.n49 a_n2094_n2688# 0.018289f
C135 plus.n50 a_n2094_n2688# 0.116592f
C136 plus.n51 a_n2094_n2688# 0.018289f
C137 plus.n52 a_n2094_n2688# 0.116592f
C138 plus.n53 a_n2094_n2688# 0.018289f
C139 plus.n54 a_n2094_n2688# 0.052222f
C140 plus.n55 a_n2094_n2688# 0.052222f
C141 plus.n56 a_n2094_n2688# 0.018289f
C142 plus.n57 a_n2094_n2688# 0.116592f
C143 plus.n58 a_n2094_n2688# 0.018289f
C144 plus.n59 a_n2094_n2688# 0.116592f
C145 plus.n60 a_n2094_n2688# 0.132982f
C146 plus.n61 a_n2094_n2688# 1.51214f
C147 source.t8 a_n2094_n2688# 2.64989f
C148 source.n0 a_n2094_n2688# 1.5075f
C149 source.t15 a_n2094_n2688# 0.248501f
C150 source.t17 a_n2094_n2688# 0.248501f
C151 source.n1 a_n2094_n2688# 2.08029f
C152 source.n2 a_n2094_n2688# 0.428535f
C153 source.t4 a_n2094_n2688# 0.248501f
C154 source.t23 a_n2094_n2688# 0.248501f
C155 source.n3 a_n2094_n2688# 2.08029f
C156 source.n4 a_n2094_n2688# 0.428535f
C157 source.t1 a_n2094_n2688# 0.248501f
C158 source.t16 a_n2094_n2688# 0.248501f
C159 source.n5 a_n2094_n2688# 2.08029f
C160 source.n6 a_n2094_n2688# 0.428535f
C161 source.t7 a_n2094_n2688# 0.248501f
C162 source.t5 a_n2094_n2688# 0.248501f
C163 source.n7 a_n2094_n2688# 2.08029f
C164 source.n8 a_n2094_n2688# 0.428535f
C165 source.t22 a_n2094_n2688# 0.248501f
C166 source.t9 a_n2094_n2688# 0.248501f
C167 source.n9 a_n2094_n2688# 2.08029f
C168 source.n10 a_n2094_n2688# 0.428535f
C169 source.t2 a_n2094_n2688# 2.64989f
C170 source.n11 a_n2094_n2688# 0.538121f
C171 source.t28 a_n2094_n2688# 2.64989f
C172 source.n12 a_n2094_n2688# 0.538121f
C173 source.t43 a_n2094_n2688# 0.248501f
C174 source.t32 a_n2094_n2688# 0.248501f
C175 source.n13 a_n2094_n2688# 2.08029f
C176 source.n14 a_n2094_n2688# 0.428535f
C177 source.t27 a_n2094_n2688# 0.248501f
C178 source.t26 a_n2094_n2688# 0.248501f
C179 source.n15 a_n2094_n2688# 2.08029f
C180 source.n16 a_n2094_n2688# 0.428535f
C181 source.t42 a_n2094_n2688# 0.248501f
C182 source.t33 a_n2094_n2688# 0.248501f
C183 source.n17 a_n2094_n2688# 2.08029f
C184 source.n18 a_n2094_n2688# 0.428535f
C185 source.t29 a_n2094_n2688# 0.248501f
C186 source.t25 a_n2094_n2688# 0.248501f
C187 source.n19 a_n2094_n2688# 2.08029f
C188 source.n20 a_n2094_n2688# 0.428535f
C189 source.t30 a_n2094_n2688# 0.248501f
C190 source.t31 a_n2094_n2688# 0.248501f
C191 source.n21 a_n2094_n2688# 2.08029f
C192 source.n22 a_n2094_n2688# 0.428535f
C193 source.t38 a_n2094_n2688# 2.64989f
C194 source.n23 a_n2094_n2688# 2.01203f
C195 source.t0 a_n2094_n2688# 2.64989f
C196 source.n24 a_n2094_n2688# 2.01203f
C197 source.t6 a_n2094_n2688# 0.248501f
C198 source.t20 a_n2094_n2688# 0.248501f
C199 source.n25 a_n2094_n2688# 2.08029f
C200 source.n26 a_n2094_n2688# 0.428542f
C201 source.t19 a_n2094_n2688# 0.248501f
C202 source.t10 a_n2094_n2688# 0.248501f
C203 source.n27 a_n2094_n2688# 2.08029f
C204 source.n28 a_n2094_n2688# 0.428542f
C205 source.t13 a_n2094_n2688# 0.248501f
C206 source.t18 a_n2094_n2688# 0.248501f
C207 source.n29 a_n2094_n2688# 2.08029f
C208 source.n30 a_n2094_n2688# 0.428542f
C209 source.t21 a_n2094_n2688# 0.248501f
C210 source.t12 a_n2094_n2688# 0.248501f
C211 source.n31 a_n2094_n2688# 2.08029f
C212 source.n32 a_n2094_n2688# 0.428542f
C213 source.t3 a_n2094_n2688# 0.248501f
C214 source.t11 a_n2094_n2688# 0.248501f
C215 source.n33 a_n2094_n2688# 2.08029f
C216 source.n34 a_n2094_n2688# 0.428542f
C217 source.t14 a_n2094_n2688# 2.64989f
C218 source.n35 a_n2094_n2688# 0.538128f
C219 source.t46 a_n2094_n2688# 2.64989f
C220 source.n36 a_n2094_n2688# 0.538128f
C221 source.t40 a_n2094_n2688# 0.248501f
C222 source.t47 a_n2094_n2688# 0.248501f
C223 source.n37 a_n2094_n2688# 2.08029f
C224 source.n38 a_n2094_n2688# 0.428542f
C225 source.t41 a_n2094_n2688# 0.248501f
C226 source.t34 a_n2094_n2688# 0.248501f
C227 source.n39 a_n2094_n2688# 2.08029f
C228 source.n40 a_n2094_n2688# 0.428542f
C229 source.t37 a_n2094_n2688# 0.248501f
C230 source.t35 a_n2094_n2688# 0.248501f
C231 source.n41 a_n2094_n2688# 2.08029f
C232 source.n42 a_n2094_n2688# 0.428542f
C233 source.t39 a_n2094_n2688# 0.248501f
C234 source.t36 a_n2094_n2688# 0.248501f
C235 source.n43 a_n2094_n2688# 2.08029f
C236 source.n44 a_n2094_n2688# 0.428542f
C237 source.t44 a_n2094_n2688# 0.248501f
C238 source.t24 a_n2094_n2688# 0.248501f
C239 source.n45 a_n2094_n2688# 2.08029f
C240 source.n46 a_n2094_n2688# 0.428542f
C241 source.t45 a_n2094_n2688# 2.64989f
C242 source.n47 a_n2094_n2688# 0.727588f
C243 source.n48 a_n2094_n2688# 1.81383f
C244 drain_right.t6 a_n2094_n2688# 0.275854f
C245 drain_right.t0 a_n2094_n2688# 0.275854f
C246 drain_right.n0 a_n2094_n2688# 2.41585f
C247 drain_right.t14 a_n2094_n2688# 0.275854f
C248 drain_right.t5 a_n2094_n2688# 0.275854f
C249 drain_right.n1 a_n2094_n2688# 2.4128f
C250 drain_right.n2 a_n2094_n2688# 0.862355f
C251 drain_right.t4 a_n2094_n2688# 0.275854f
C252 drain_right.t12 a_n2094_n2688# 0.275854f
C253 drain_right.n3 a_n2094_n2688# 2.4128f
C254 drain_right.n4 a_n2094_n2688# 0.394617f
C255 drain_right.t7 a_n2094_n2688# 0.275854f
C256 drain_right.t23 a_n2094_n2688# 0.275854f
C257 drain_right.n5 a_n2094_n2688# 2.41585f
C258 drain_right.t1 a_n2094_n2688# 0.275854f
C259 drain_right.t22 a_n2094_n2688# 0.275854f
C260 drain_right.n6 a_n2094_n2688# 2.4128f
C261 drain_right.n7 a_n2094_n2688# 0.862355f
C262 drain_right.t11 a_n2094_n2688# 0.275854f
C263 drain_right.t3 a_n2094_n2688# 0.275854f
C264 drain_right.n8 a_n2094_n2688# 2.4128f
C265 drain_right.n9 a_n2094_n2688# 0.394617f
C266 drain_right.n10 a_n2094_n2688# 1.64727f
C267 drain_right.t20 a_n2094_n2688# 0.275854f
C268 drain_right.t15 a_n2094_n2688# 0.275854f
C269 drain_right.n11 a_n2094_n2688# 2.41584f
C270 drain_right.t17 a_n2094_n2688# 0.275854f
C271 drain_right.t21 a_n2094_n2688# 0.275854f
C272 drain_right.n12 a_n2094_n2688# 2.4128f
C273 drain_right.n13 a_n2094_n2688# 0.862355f
C274 drain_right.t10 a_n2094_n2688# 0.275854f
C275 drain_right.t16 a_n2094_n2688# 0.275854f
C276 drain_right.n14 a_n2094_n2688# 2.4128f
C277 drain_right.n15 a_n2094_n2688# 0.424886f
C278 drain_right.t19 a_n2094_n2688# 0.275854f
C279 drain_right.t13 a_n2094_n2688# 0.275854f
C280 drain_right.n16 a_n2094_n2688# 2.4128f
C281 drain_right.n17 a_n2094_n2688# 0.424886f
C282 drain_right.t18 a_n2094_n2688# 0.275854f
C283 drain_right.t8 a_n2094_n2688# 0.275854f
C284 drain_right.n18 a_n2094_n2688# 2.4128f
C285 drain_right.n19 a_n2094_n2688# 0.424886f
C286 drain_right.t2 a_n2094_n2688# 0.275854f
C287 drain_right.t9 a_n2094_n2688# 0.275854f
C288 drain_right.n20 a_n2094_n2688# 2.4128f
C289 drain_right.n21 a_n2094_n2688# 0.742319f
C290 minus.n0 a_n2094_n2688# 0.051151f
C291 minus.t9 a_n2094_n2688# 0.266381f
C292 minus.t17 a_n2094_n2688# 0.260895f
C293 minus.t16 a_n2094_n2688# 0.260895f
C294 minus.t18 a_n2094_n2688# 0.260895f
C295 minus.n1 a_n2094_n2688# 0.114201f
C296 minus.n2 a_n2094_n2688# 0.051151f
C297 minus.t22 a_n2094_n2688# 0.260895f
C298 minus.t5 a_n2094_n2688# 0.260895f
C299 minus.t14 a_n2094_n2688# 0.260895f
C300 minus.n3 a_n2094_n2688# 0.114201f
C301 minus.n4 a_n2094_n2688# 0.051151f
C302 minus.t20 a_n2094_n2688# 0.260895f
C303 minus.t21 a_n2094_n2688# 0.260895f
C304 minus.t4 a_n2094_n2688# 0.260895f
C305 minus.n5 a_n2094_n2688# 0.114201f
C306 minus.t19 a_n2094_n2688# 0.266381f
C307 minus.n6 a_n2094_n2688# 0.130336f
C308 minus.t15 a_n2094_n2688# 0.260895f
C309 minus.n7 a_n2094_n2688# 0.114201f
C310 minus.n8 a_n2094_n2688# 0.017914f
C311 minus.n9 a_n2094_n2688# 0.118937f
C312 minus.n10 a_n2094_n2688# 0.051151f
C313 minus.n11 a_n2094_n2688# 0.017914f
C314 minus.n12 a_n2094_n2688# 0.114201f
C315 minus.n13 a_n2094_n2688# 0.017914f
C316 minus.n14 a_n2094_n2688# 0.114201f
C317 minus.n15 a_n2094_n2688# 0.017914f
C318 minus.n16 a_n2094_n2688# 0.051151f
C319 minus.n17 a_n2094_n2688# 0.051151f
C320 minus.n18 a_n2094_n2688# 0.017914f
C321 minus.n19 a_n2094_n2688# 0.114201f
C322 minus.n20 a_n2094_n2688# 0.017914f
C323 minus.n21 a_n2094_n2688# 0.114201f
C324 minus.n22 a_n2094_n2688# 0.017914f
C325 minus.n23 a_n2094_n2688# 0.051151f
C326 minus.n24 a_n2094_n2688# 0.051151f
C327 minus.n25 a_n2094_n2688# 0.017914f
C328 minus.n26 a_n2094_n2688# 0.114201f
C329 minus.n27 a_n2094_n2688# 0.017914f
C330 minus.n28 a_n2094_n2688# 0.114201f
C331 minus.n29 a_n2094_n2688# 0.130256f
C332 minus.n30 a_n2094_n2688# 1.69635f
C333 minus.n31 a_n2094_n2688# 0.051151f
C334 minus.t23 a_n2094_n2688# 0.260895f
C335 minus.t3 a_n2094_n2688# 0.260895f
C336 minus.t11 a_n2094_n2688# 0.260895f
C337 minus.n32 a_n2094_n2688# 0.114201f
C338 minus.n33 a_n2094_n2688# 0.051151f
C339 minus.t8 a_n2094_n2688# 0.260895f
C340 minus.t12 a_n2094_n2688# 0.260895f
C341 minus.t10 a_n2094_n2688# 0.260895f
C342 minus.n34 a_n2094_n2688# 0.114201f
C343 minus.n35 a_n2094_n2688# 0.051151f
C344 minus.t13 a_n2094_n2688# 0.260895f
C345 minus.t6 a_n2094_n2688# 0.260895f
C346 minus.t0 a_n2094_n2688# 0.260895f
C347 minus.n36 a_n2094_n2688# 0.114201f
C348 minus.t1 a_n2094_n2688# 0.266381f
C349 minus.n37 a_n2094_n2688# 0.130336f
C350 minus.t7 a_n2094_n2688# 0.260895f
C351 minus.n38 a_n2094_n2688# 0.114201f
C352 minus.n39 a_n2094_n2688# 0.017914f
C353 minus.n40 a_n2094_n2688# 0.118937f
C354 minus.n41 a_n2094_n2688# 0.051151f
C355 minus.n42 a_n2094_n2688# 0.017914f
C356 minus.n43 a_n2094_n2688# 0.114201f
C357 minus.n44 a_n2094_n2688# 0.017914f
C358 minus.n45 a_n2094_n2688# 0.114201f
C359 minus.n46 a_n2094_n2688# 0.017914f
C360 minus.n47 a_n2094_n2688# 0.051151f
C361 minus.n48 a_n2094_n2688# 0.051151f
C362 minus.n49 a_n2094_n2688# 0.017914f
C363 minus.n50 a_n2094_n2688# 0.114201f
C364 minus.n51 a_n2094_n2688# 0.017914f
C365 minus.n52 a_n2094_n2688# 0.114201f
C366 minus.n53 a_n2094_n2688# 0.017914f
C367 minus.n54 a_n2094_n2688# 0.051151f
C368 minus.n55 a_n2094_n2688# 0.051151f
C369 minus.n56 a_n2094_n2688# 0.017914f
C370 minus.n57 a_n2094_n2688# 0.114201f
C371 minus.n58 a_n2094_n2688# 0.017914f
C372 minus.n59 a_n2094_n2688# 0.114201f
C373 minus.t2 a_n2094_n2688# 0.266381f
C374 minus.n60 a_n2094_n2688# 0.130256f
C375 minus.n61 a_n2094_n2688# 0.333102f
C376 minus.n62 a_n2094_n2688# 2.06957f
.ends

