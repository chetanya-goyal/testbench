* NGSPICE file created from diffpair514.ext - technology: sky130A

.subckt diffpair514 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t13 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X1 drain_left.t8 plus.t1 source.t16 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X2 drain_right.t9 minus.t0 source.t19 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X3 a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X4 a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X5 drain_left.t7 plus.t2 source.t8 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X6 drain_right.t8 minus.t1 source.t3 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X7 drain_right.t7 minus.t2 source.t2 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X8 drain_left.t6 plus.t3 source.t10 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X9 drain_left.t5 plus.t4 source.t12 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X10 source.t15 plus.t5 drain_left.t4 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X11 source.t5 minus.t3 drain_right.t6 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X12 drain_right.t5 minus.t4 source.t1 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X13 a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X14 drain_right.t4 minus.t5 source.t18 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X15 source.t9 plus.t6 drain_left.t3 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X16 drain_left.t2 plus.t7 source.t11 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X18 source.t7 plus.t8 drain_left.t1 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X19 drain_right.t3 minus.t6 source.t4 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X20 source.t17 minus.t7 drain_right.t2 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X21 source.t6 minus.t8 drain_right.t1 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X22 source.t0 minus.t9 drain_right.t0 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 source.t14 plus.t9 drain_left.t0 a_n1472_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 plus.n3 plus.t2 1347.41
R1 plus.n9 plus.t4 1347.41
R2 plus.n14 plus.t0 1347.41
R3 plus.n20 plus.t3 1347.41
R4 plus.n6 plus.t7 1309.43
R5 plus.n2 plus.t5 1309.43
R6 plus.n8 plus.t9 1309.43
R7 plus.n17 plus.t1 1309.43
R8 plus.n13 plus.t6 1309.43
R9 plus.n19 plus.t8 1309.43
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 54.0429
R25 plus.n9 plus.n8 54.0429
R26 plus.n20 plus.n19 54.0429
R27 plus.n14 plus.n13 54.0429
R28 plus plus.n21 29.7017
R29 plus.n2 plus.n1 18.9884
R30 plus.n8 plus.n7 18.9884
R31 plus.n19 plus.n18 18.9884
R32 plus.n13 plus.n12 18.9884
R33 plus plus.n10 13.2675
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n5 source.t18 45.521
R41 source.n19 source.t1 45.5208
R42 source.n14 source.t13 45.5208
R43 source.n0 source.t12 45.5208
R44 source.n2 source.n1 44.201
R45 source.n4 source.n3 44.201
R46 source.n7 source.n6 44.201
R47 source.n9 source.n8 44.201
R48 source.n18 source.n17 44.2008
R49 source.n16 source.n15 44.2008
R50 source.n13 source.n12 44.2008
R51 source.n11 source.n10 44.2008
R52 source.n11 source.n9 24.6467
R53 source.n20 source.n0 18.5691
R54 source.n20 source.n19 5.53498
R55 source.n17 source.t3 1.3205
R56 source.n17 source.t17 1.3205
R57 source.n15 source.t2 1.3205
R58 source.n15 source.t6 1.3205
R59 source.n12 source.t16 1.3205
R60 source.n12 source.t9 1.3205
R61 source.n10 source.t10 1.3205
R62 source.n10 source.t7 1.3205
R63 source.n1 source.t11 1.3205
R64 source.n1 source.t14 1.3205
R65 source.n3 source.t8 1.3205
R66 source.n3 source.t15 1.3205
R67 source.n6 source.t19 1.3205
R68 source.n6 source.t0 1.3205
R69 source.n8 source.t4 1.3205
R70 source.n8 source.t5 1.3205
R71 source.n5 source.n4 0.741879
R72 source.n16 source.n14 0.741879
R73 source.n9 source.n7 0.543603
R74 source.n7 source.n5 0.543603
R75 source.n4 source.n2 0.543603
R76 source.n2 source.n0 0.543603
R77 source.n13 source.n11 0.543603
R78 source.n14 source.n13 0.543603
R79 source.n18 source.n16 0.543603
R80 source.n19 source.n18 0.543603
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t7 62.7429
R83 drain_left.n1 drain_left.t6 62.7427
R84 drain_left.n3 drain_left.n2 61.2315
R85 drain_left.n5 drain_left.n4 60.8798
R86 drain_left.n7 drain_left.n6 60.8796
R87 drain_left.n1 drain_left.n0 60.8796
R88 drain_left drain_left.n3 31.948
R89 drain_left drain_left.n7 6.19632
R90 drain_left.n2 drain_left.t3 1.3205
R91 drain_left.n2 drain_left.t9 1.3205
R92 drain_left.n0 drain_left.t1 1.3205
R93 drain_left.n0 drain_left.t8 1.3205
R94 drain_left.n6 drain_left.t0 1.3205
R95 drain_left.n6 drain_left.t5 1.3205
R96 drain_left.n4 drain_left.t4 1.3205
R97 drain_left.n4 drain_left.t2 1.3205
R98 drain_left.n7 drain_left.n5 0.543603
R99 drain_left.n3 drain_left.n1 0.0809298
R100 minus.n9 minus.t6 1347.41
R101 minus.n3 minus.t5 1347.41
R102 minus.n20 minus.t4 1347.41
R103 minus.n14 minus.t2 1347.41
R104 minus.n6 minus.t0 1309.43
R105 minus.n8 minus.t3 1309.43
R106 minus.n2 minus.t9 1309.43
R107 minus.n17 minus.t1 1309.43
R108 minus.n19 minus.t7 1309.43
R109 minus.n13 minus.t8 1309.43
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 54.0429
R125 minus.n3 minus.n2 54.0429
R126 minus.n14 minus.n13 54.0429
R127 minus.n20 minus.n19 54.0429
R128 minus.n22 minus.n10 36.9569
R129 minus.n8 minus.n7 18.9884
R130 minus.n2 minus.n1 18.9884
R131 minus.n13 minus.n12 18.9884
R132 minus.n19 minus.n18 18.9884
R133 minus.n22 minus.n21 6.48724
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t7 62.7427
R142 drain_right.n7 drain_right.t3 62.1998
R143 drain_right.n6 drain_right.n4 61.4227
R144 drain_right.n3 drain_right.n2 61.2315
R145 drain_right.n6 drain_right.n5 60.8798
R146 drain_right.n1 drain_right.n0 60.8796
R147 drain_right drain_right.n3 31.3948
R148 drain_right drain_right.n7 5.92477
R149 drain_right.n2 drain_right.t2 1.3205
R150 drain_right.n2 drain_right.t5 1.3205
R151 drain_right.n0 drain_right.t1 1.3205
R152 drain_right.n0 drain_right.t8 1.3205
R153 drain_right.n4 drain_right.t0 1.3205
R154 drain_right.n4 drain_right.t4 1.3205
R155 drain_right.n5 drain_right.t6 1.3205
R156 drain_right.n5 drain_right.t9 1.3205
R157 drain_right.n7 drain_right.n6 0.543603
R158 drain_right.n3 drain_right.n1 0.0809298
C0 plus minus 5.54342f
C1 drain_right plus 0.297192f
C2 source drain_left 25.7745f
C3 minus drain_left 0.171269f
C4 drain_right drain_left 0.725979f
C5 source minus 4.37285f
C6 drain_right source 25.761f
C7 plus drain_left 5.03748f
C8 drain_right minus 4.90061f
C9 source plus 4.3877f
C10 drain_right a_n1472_n3888# 7.801401f
C11 drain_left a_n1472_n3888# 8.04004f
C12 source a_n1472_n3888# 7.148392f
C13 minus a_n1472_n3888# 5.894818f
C14 plus a_n1472_n3888# 8.07864f
C15 drain_right.t7 a_n1472_n3888# 4.07396f
C16 drain_right.t1 a_n1472_n3888# 0.352811f
C17 drain_right.t8 a_n1472_n3888# 0.352811f
C18 drain_right.n0 a_n1472_n3888# 3.189f
C19 drain_right.n1 a_n1472_n3888# 0.697282f
C20 drain_right.t2 a_n1472_n3888# 0.352811f
C21 drain_right.t5 a_n1472_n3888# 0.352811f
C22 drain_right.n2 a_n1472_n3888# 3.19097f
C23 drain_right.n3 a_n1472_n3888# 1.82906f
C24 drain_right.t0 a_n1472_n3888# 0.352811f
C25 drain_right.t4 a_n1472_n3888# 0.352811f
C26 drain_right.n4 a_n1472_n3888# 3.19217f
C27 drain_right.t6 a_n1472_n3888# 0.352811f
C28 drain_right.t9 a_n1472_n3888# 0.352811f
C29 drain_right.n5 a_n1472_n3888# 3.189f
C30 drain_right.n6 a_n1472_n3888# 0.70474f
C31 drain_right.t3 a_n1472_n3888# 4.0706f
C32 drain_right.n7 a_n1472_n3888# 0.636781f
C33 minus.n0 a_n1472_n3888# 0.053599f
C34 minus.t6 a_n1472_n3888# 0.687874f
C35 minus.t3 a_n1472_n3888# 0.680452f
C36 minus.t0 a_n1472_n3888# 0.680452f
C37 minus.n1 a_n1472_n3888# 0.022077f
C38 minus.t9 a_n1472_n3888# 0.680452f
C39 minus.n2 a_n1472_n3888# 0.261366f
C40 minus.t5 a_n1472_n3888# 0.687874f
C41 minus.n3 a_n1472_n3888# 0.278078f
C42 minus.n4 a_n1472_n3888# 0.117698f
C43 minus.n5 a_n1472_n3888# 0.053599f
C44 minus.n6 a_n1472_n3888# 0.279146f
C45 minus.n7 a_n1472_n3888# 0.022077f
C46 minus.n8 a_n1472_n3888# 0.261366f
C47 minus.n9 a_n1472_n3888# 0.278003f
C48 minus.n10 a_n1472_n3888# 1.95627f
C49 minus.n11 a_n1472_n3888# 0.053599f
C50 minus.t7 a_n1472_n3888# 0.680452f
C51 minus.t1 a_n1472_n3888# 0.680452f
C52 minus.n12 a_n1472_n3888# 0.022077f
C53 minus.t2 a_n1472_n3888# 0.687874f
C54 minus.t8 a_n1472_n3888# 0.680452f
C55 minus.n13 a_n1472_n3888# 0.261366f
C56 minus.n14 a_n1472_n3888# 0.278078f
C57 minus.n15 a_n1472_n3888# 0.117698f
C58 minus.n16 a_n1472_n3888# 0.053599f
C59 minus.n17 a_n1472_n3888# 0.279146f
C60 minus.n18 a_n1472_n3888# 0.022077f
C61 minus.n19 a_n1472_n3888# 0.261366f
C62 minus.t4 a_n1472_n3888# 0.687874f
C63 minus.n20 a_n1472_n3888# 0.278003f
C64 minus.n21 a_n1472_n3888# 0.348806f
C65 minus.n22 a_n1472_n3888# 2.3715f
C66 drain_left.t6 a_n1472_n3888# 4.07179f
C67 drain_left.t1 a_n1472_n3888# 0.352623f
C68 drain_left.t8 a_n1472_n3888# 0.352623f
C69 drain_left.n0 a_n1472_n3888# 3.1873f
C70 drain_left.n1 a_n1472_n3888# 0.69691f
C71 drain_left.t3 a_n1472_n3888# 0.352623f
C72 drain_left.t9 a_n1472_n3888# 0.352623f
C73 drain_left.n2 a_n1472_n3888# 3.18927f
C74 drain_left.n3 a_n1472_n3888# 1.89041f
C75 drain_left.t7 a_n1472_n3888# 4.07179f
C76 drain_left.t4 a_n1472_n3888# 0.352623f
C77 drain_left.t2 a_n1472_n3888# 0.352623f
C78 drain_left.n4 a_n1472_n3888# 3.1873f
C79 drain_left.n5 a_n1472_n3888# 0.73268f
C80 drain_left.t0 a_n1472_n3888# 0.352623f
C81 drain_left.t5 a_n1472_n3888# 0.352623f
C82 drain_left.n6 a_n1472_n3888# 3.18729f
C83 drain_left.n7 a_n1472_n3888# 0.595403f
C84 source.t12 a_n1472_n3888# 4.04842f
C85 source.n0 a_n1472_n3888# 1.87515f
C86 source.t11 a_n1472_n3888# 0.361253f
C87 source.t14 a_n1472_n3888# 0.361253f
C88 source.n1 a_n1472_n3888# 3.1733f
C89 source.n2 a_n1472_n3888# 0.406866f
C90 source.t8 a_n1472_n3888# 0.361253f
C91 source.t15 a_n1472_n3888# 0.361253f
C92 source.n3 a_n1472_n3888# 3.1733f
C93 source.n4 a_n1472_n3888# 0.426337f
C94 source.t18 a_n1472_n3888# 4.04842f
C95 source.n5 a_n1472_n3888# 0.53645f
C96 source.t19 a_n1472_n3888# 0.361253f
C97 source.t0 a_n1472_n3888# 0.361253f
C98 source.n6 a_n1472_n3888# 3.1733f
C99 source.n7 a_n1472_n3888# 0.406866f
C100 source.t4 a_n1472_n3888# 0.361253f
C101 source.t5 a_n1472_n3888# 0.361253f
C102 source.n8 a_n1472_n3888# 3.1733f
C103 source.n9 a_n1472_n3888# 2.32507f
C104 source.t10 a_n1472_n3888# 0.361253f
C105 source.t7 a_n1472_n3888# 0.361253f
C106 source.n10 a_n1472_n3888# 3.1733f
C107 source.n11 a_n1472_n3888# 2.32507f
C108 source.t16 a_n1472_n3888# 0.361253f
C109 source.t9 a_n1472_n3888# 0.361253f
C110 source.n12 a_n1472_n3888# 3.1733f
C111 source.n13 a_n1472_n3888# 0.40687f
C112 source.t13 a_n1472_n3888# 4.04842f
C113 source.n14 a_n1472_n3888# 0.536455f
C114 source.t2 a_n1472_n3888# 0.361253f
C115 source.t6 a_n1472_n3888# 0.361253f
C116 source.n15 a_n1472_n3888# 3.1733f
C117 source.n16 a_n1472_n3888# 0.426341f
C118 source.t3 a_n1472_n3888# 0.361253f
C119 source.t17 a_n1472_n3888# 0.361253f
C120 source.n17 a_n1472_n3888# 3.1733f
C121 source.n18 a_n1472_n3888# 0.40687f
C122 source.t1 a_n1472_n3888# 4.04842f
C123 source.n19 a_n1472_n3888# 0.681828f
C124 source.n20 a_n1472_n3888# 2.2284f
C125 plus.n0 a_n1472_n3888# 0.054359f
C126 plus.t9 a_n1472_n3888# 0.690103f
C127 plus.t7 a_n1472_n3888# 0.690103f
C128 plus.n1 a_n1472_n3888# 0.02239f
C129 plus.t2 a_n1472_n3888# 0.697631f
C130 plus.t5 a_n1472_n3888# 0.690103f
C131 plus.n2 a_n1472_n3888# 0.265073f
C132 plus.n3 a_n1472_n3888# 0.282022f
C133 plus.n4 a_n1472_n3888# 0.119367f
C134 plus.n5 a_n1472_n3888# 0.054359f
C135 plus.n6 a_n1472_n3888# 0.283106f
C136 plus.n7 a_n1472_n3888# 0.02239f
C137 plus.n8 a_n1472_n3888# 0.265073f
C138 plus.t4 a_n1472_n3888# 0.697631f
C139 plus.n9 a_n1472_n3888# 0.281946f
C140 plus.n10 a_n1472_n3888# 0.685298f
C141 plus.n11 a_n1472_n3888# 0.054359f
C142 plus.t3 a_n1472_n3888# 0.697631f
C143 plus.t8 a_n1472_n3888# 0.690103f
C144 plus.t1 a_n1472_n3888# 0.690103f
C145 plus.n12 a_n1472_n3888# 0.02239f
C146 plus.t6 a_n1472_n3888# 0.690103f
C147 plus.n13 a_n1472_n3888# 0.265073f
C148 plus.t0 a_n1472_n3888# 0.697631f
C149 plus.n14 a_n1472_n3888# 0.282022f
C150 plus.n15 a_n1472_n3888# 0.119367f
C151 plus.n16 a_n1472_n3888# 0.054359f
C152 plus.n17 a_n1472_n3888# 0.283106f
C153 plus.n18 a_n1472_n3888# 0.02239f
C154 plus.n19 a_n1472_n3888# 0.265073f
C155 plus.n20 a_n1472_n3888# 0.281946f
C156 plus.n21 a_n1472_n3888# 1.62567f
.ends

