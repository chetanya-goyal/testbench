* NGSPICE file created from diffpair595.ext - technology: sky130A

.subckt diffpair595 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t12 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 drain_left.t10 plus.t1 source.t17 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X2 source.t11 minus.t0 drain_right.t11 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X3 drain_right.t10 minus.t1 source.t6 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X4 a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X5 source.t3 minus.t2 drain_right.t9 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X6 source.t4 minus.t3 drain_right.t8 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X7 source.t23 plus.t2 drain_left.t9 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X8 a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X9 drain_left.t8 plus.t3 source.t21 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X10 source.t16 plus.t4 drain_left.t7 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X11 a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X12 a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X13 drain_left.t6 plus.t5 source.t15 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X14 source.t7 minus.t4 drain_right.t7 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X15 source.t8 minus.t5 drain_right.t6 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X16 drain_right.t5 minus.t6 source.t0 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X17 drain_left.t5 plus.t6 source.t18 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X18 source.t19 plus.t7 drain_left.t4 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X19 source.t20 plus.t8 drain_left.t3 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X20 source.t22 plus.t9 drain_left.t2 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X21 source.t14 plus.t10 drain_left.t1 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X22 drain_right.t4 minus.t7 source.t10 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X23 drain_right.t3 minus.t8 source.t2 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X24 drain_right.t2 minus.t9 source.t1 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X25 source.t5 minus.t10 drain_right.t1 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X26 drain_right.t0 minus.t11 source.t9 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X27 drain_left.t0 plus.t11 source.t13 a_n1598_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
R0 plus.n2 plus.t2 1758.57
R1 plus.n13 plus.t6 1758.57
R2 plus.n17 plus.t0 1758.57
R3 plus.n28 plus.t10 1758.57
R4 plus.n3 plus.t5 1711.1
R5 plus.n4 plus.t8 1711.1
R6 plus.n10 plus.t11 1711.1
R7 plus.n12 plus.t4 1711.1
R8 plus.n19 plus.t7 1711.1
R9 plus.n18 plus.t1 1711.1
R10 plus.n25 plus.t9 1711.1
R11 plus.n27 plus.t3 1711.1
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 63.5369
R27 plus.n11 plus.n10 63.5369
R28 plus.n26 plus.n25 63.5369
R29 plus.n20 plus.n18 63.5369
R30 plus.n3 plus.n2 44.549
R31 plus.n13 plus.n12 44.549
R32 plus.n28 plus.n27 44.549
R33 plus.n19 plus.n17 44.549
R34 plus plus.n29 32.0975
R35 plus.n5 plus.n3 28.4823
R36 plus.n12 plus.n11 28.4823
R37 plus.n27 plus.n26 28.4823
R38 plus.n20 plus.n19 28.4823
R39 plus plus.n14 15.1861
R40 plus.n4 plus.n1 9.49444
R41 plus.n10 plus.n9 9.49444
R42 plus.n25 plus.n24 9.49444
R43 plus.n18 plus.n16 9.49444
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n0 source.t18 44.1297
R53 source.n5 source.t23 44.1296
R54 source.n6 source.t0 44.1296
R55 source.n11 source.t11 44.1296
R56 source.n23 source.t9 44.1295
R57 source.n18 source.t4 44.1295
R58 source.n17 source.t12 44.1295
R59 source.n12 source.t14 44.1295
R60 source.n2 source.n1 43.1397
R61 source.n4 source.n3 43.1397
R62 source.n8 source.n7 43.1397
R63 source.n10 source.n9 43.1397
R64 source.n22 source.n21 43.1396
R65 source.n20 source.n19 43.1396
R66 source.n16 source.n15 43.1396
R67 source.n14 source.n13 43.1396
R68 source.n12 source.n11 27.8914
R69 source.n24 source.n0 22.357
R70 source.n24 source.n23 5.53498
R71 source.n21 source.t10 0.9905
R72 source.n21 source.t7 0.9905
R73 source.n19 source.t2 0.9905
R74 source.n19 source.t3 0.9905
R75 source.n15 source.t17 0.9905
R76 source.n15 source.t19 0.9905
R77 source.n13 source.t21 0.9905
R78 source.n13 source.t22 0.9905
R79 source.n1 source.t13 0.9905
R80 source.n1 source.t16 0.9905
R81 source.n3 source.t15 0.9905
R82 source.n3 source.t20 0.9905
R83 source.n7 source.t6 0.9905
R84 source.n7 source.t5 0.9905
R85 source.n9 source.t1 0.9905
R86 source.n9 source.t8 0.9905
R87 source.n11 source.n10 0.543603
R88 source.n10 source.n8 0.543603
R89 source.n8 source.n6 0.543603
R90 source.n5 source.n4 0.543603
R91 source.n4 source.n2 0.543603
R92 source.n2 source.n0 0.543603
R93 source.n14 source.n12 0.543603
R94 source.n16 source.n14 0.543603
R95 source.n17 source.n16 0.543603
R96 source.n20 source.n18 0.543603
R97 source.n22 source.n20 0.543603
R98 source.n23 source.n22 0.543603
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 60.3616
R103 drain_left.n3 drain_left.n2 60.3062
R104 drain_left.n3 drain_left.n0 60.3062
R105 drain_left.n8 drain_left.n7 59.8185
R106 drain_left.n6 drain_left.n5 59.8185
R107 drain_left.n3 drain_left.n1 59.8184
R108 drain_left drain_left.n3 36.1432
R109 drain_left drain_left.n8 6.19632
R110 drain_left.n1 drain_left.t2 0.9905
R111 drain_left.n1 drain_left.t10 0.9905
R112 drain_left.n2 drain_left.t4 0.9905
R113 drain_left.n2 drain_left.t11 0.9905
R114 drain_left.n0 drain_left.t1 0.9905
R115 drain_left.n0 drain_left.t8 0.9905
R116 drain_left.n7 drain_left.t7 0.9905
R117 drain_left.n7 drain_left.t5 0.9905
R118 drain_left.n5 drain_left.t3 0.9905
R119 drain_left.n5 drain_left.t0 0.9905
R120 drain_left.n4 drain_left.t9 0.9905
R121 drain_left.n4 drain_left.t6 0.9905
R122 drain_left.n8 drain_left.n6 0.543603
R123 minus.n13 minus.t0 1758.57
R124 minus.n2 minus.t6 1758.57
R125 minus.n28 minus.t11 1758.57
R126 minus.n17 minus.t3 1758.57
R127 minus.n12 minus.t9 1711.1
R128 minus.n10 minus.t5 1711.1
R129 minus.n3 minus.t1 1711.1
R130 minus.n4 minus.t10 1711.1
R131 minus.n27 minus.t4 1711.1
R132 minus.n25 minus.t7 1711.1
R133 minus.n19 minus.t2 1711.1
R134 minus.n18 minus.t8 1711.1
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 63.5369
R150 minus.n5 minus.n3 63.5369
R151 minus.n20 minus.n19 63.5369
R152 minus.n26 minus.n25 63.5369
R153 minus.n13 minus.n12 44.549
R154 minus.n4 minus.n2 44.549
R155 minus.n18 minus.n17 44.549
R156 minus.n28 minus.n27 44.549
R157 minus.n30 minus.n14 41.2467
R158 minus.n12 minus.n11 28.4823
R159 minus.n5 minus.n4 28.4823
R160 minus.n20 minus.n18 28.4823
R161 minus.n27 minus.n26 28.4823
R162 minus.n10 minus.n9 9.49444
R163 minus.n3 minus.n1 9.49444
R164 minus.n19 minus.n16 9.49444
R165 minus.n25 minus.n24 9.49444
R166 minus.n30 minus.n29 6.51186
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 60.3616
R177 drain_right.n3 drain_right.n2 60.3062
R178 drain_right.n3 drain_right.n0 60.3062
R179 drain_right.n6 drain_right.n5 59.8185
R180 drain_right.n8 drain_right.n7 59.8185
R181 drain_right.n3 drain_right.n1 59.8184
R182 drain_right drain_right.n3 35.59
R183 drain_right drain_right.n8 6.19632
R184 drain_right.n1 drain_right.t9 0.9905
R185 drain_right.n1 drain_right.t4 0.9905
R186 drain_right.n2 drain_right.t7 0.9905
R187 drain_right.n2 drain_right.t0 0.9905
R188 drain_right.n0 drain_right.t8 0.9905
R189 drain_right.n0 drain_right.t3 0.9905
R190 drain_right.n4 drain_right.t1 0.9905
R191 drain_right.n4 drain_right.t5 0.9905
R192 drain_right.n5 drain_right.t6 0.9905
R193 drain_right.n5 drain_right.t10 0.9905
R194 drain_right.n7 drain_right.t11 0.9905
R195 drain_right.n7 drain_right.t2 0.9905
R196 drain_right.n8 drain_right.n6 0.543603
C0 plus drain_right 0.30725f
C1 source drain_left 37.6634f
C2 minus plus 6.62501f
C3 source drain_right 37.663105f
C4 source minus 6.72243f
C5 source plus 6.73647f
C6 drain_right drain_left 0.785787f
C7 minus drain_left 0.170859f
C8 plus drain_left 7.59121f
C9 minus drain_right 7.43776f
C10 drain_right a_n1598_n4888# 7.87242f
C11 drain_left a_n1598_n4888# 8.12939f
C12 source a_n1598_n4888# 12.979519f
C13 minus a_n1598_n4888# 6.738831f
C14 plus a_n1598_n4888# 9.25458f
C15 drain_right.t8 a_n1598_n4888# 0.537988f
C16 drain_right.t3 a_n1598_n4888# 0.537988f
C17 drain_right.n0 a_n1598_n4888# 4.92176f
C18 drain_right.t9 a_n1598_n4888# 0.537988f
C19 drain_right.t4 a_n1598_n4888# 0.537988f
C20 drain_right.n1 a_n1598_n4888# 4.9184f
C21 drain_right.t7 a_n1598_n4888# 0.537988f
C22 drain_right.t0 a_n1598_n4888# 0.537988f
C23 drain_right.n2 a_n1598_n4888# 4.92176f
C24 drain_right.n3 a_n1598_n4888# 3.3527f
C25 drain_right.t1 a_n1598_n4888# 0.537988f
C26 drain_right.t5 a_n1598_n4888# 0.537988f
C27 drain_right.n4 a_n1598_n4888# 4.92218f
C28 drain_right.t6 a_n1598_n4888# 0.537988f
C29 drain_right.t10 a_n1598_n4888# 0.537988f
C30 drain_right.n5 a_n1598_n4888# 4.9184f
C31 drain_right.n6 a_n1598_n4888# 0.822721f
C32 drain_right.t11 a_n1598_n4888# 0.537988f
C33 drain_right.t2 a_n1598_n4888# 0.537988f
C34 drain_right.n7 a_n1598_n4888# 4.9184f
C35 drain_right.n8 a_n1598_n4888# 0.68973f
C36 minus.n0 a_n1598_n4888# 0.05231f
C37 minus.t0 a_n1598_n4888# 0.89296f
C38 minus.t9 a_n1598_n4888# 0.883987f
C39 minus.t5 a_n1598_n4888# 0.883987f
C40 minus.n1 a_n1598_n4888# 0.019449f
C41 minus.t6 a_n1598_n4888# 0.89296f
C42 minus.n2 a_n1598_n4888# 0.345063f
C43 minus.t1 a_n1598_n4888# 0.883987f
C44 minus.n3 a_n1598_n4888# 0.32838f
C45 minus.t10 a_n1598_n4888# 0.883987f
C46 minus.n4 a_n1598_n4888# 0.32838f
C47 minus.n5 a_n1598_n4888# 0.021546f
C48 minus.n6 a_n1598_n4888# 0.119056f
C49 minus.n7 a_n1598_n4888# 0.05231f
C50 minus.n8 a_n1598_n4888# 0.05231f
C51 minus.n9 a_n1598_n4888# 0.019449f
C52 minus.n10 a_n1598_n4888# 0.32838f
C53 minus.n11 a_n1598_n4888# 0.021546f
C54 minus.n12 a_n1598_n4888# 0.32838f
C55 minus.n13 a_n1598_n4888# 0.344984f
C56 minus.n14 a_n1598_n4888# 2.25593f
C57 minus.n15 a_n1598_n4888# 0.05231f
C58 minus.t4 a_n1598_n4888# 0.883987f
C59 minus.t7 a_n1598_n4888# 0.883987f
C60 minus.n16 a_n1598_n4888# 0.019449f
C61 minus.t3 a_n1598_n4888# 0.89296f
C62 minus.n17 a_n1598_n4888# 0.345063f
C63 minus.t8 a_n1598_n4888# 0.883987f
C64 minus.n18 a_n1598_n4888# 0.32838f
C65 minus.t2 a_n1598_n4888# 0.883987f
C66 minus.n19 a_n1598_n4888# 0.32838f
C67 minus.n20 a_n1598_n4888# 0.021546f
C68 minus.n21 a_n1598_n4888# 0.119056f
C69 minus.n22 a_n1598_n4888# 0.05231f
C70 minus.n23 a_n1598_n4888# 0.05231f
C71 minus.n24 a_n1598_n4888# 0.019449f
C72 minus.n25 a_n1598_n4888# 0.32838f
C73 minus.n26 a_n1598_n4888# 0.021546f
C74 minus.n27 a_n1598_n4888# 0.32838f
C75 minus.t11 a_n1598_n4888# 0.89296f
C76 minus.n28 a_n1598_n4888# 0.344984f
C77 minus.n29 a_n1598_n4888# 0.343453f
C78 minus.n30 a_n1598_n4888# 2.69944f
C79 drain_left.t1 a_n1598_n4888# 0.538783f
C80 drain_left.t8 a_n1598_n4888# 0.538783f
C81 drain_left.n0 a_n1598_n4888# 4.92904f
C82 drain_left.t2 a_n1598_n4888# 0.538783f
C83 drain_left.t10 a_n1598_n4888# 0.538783f
C84 drain_left.n1 a_n1598_n4888# 4.92567f
C85 drain_left.t4 a_n1598_n4888# 0.538783f
C86 drain_left.t11 a_n1598_n4888# 0.538783f
C87 drain_left.n2 a_n1598_n4888# 4.92904f
C88 drain_left.n3 a_n1598_n4888# 3.42888f
C89 drain_left.t9 a_n1598_n4888# 0.538783f
C90 drain_left.t6 a_n1598_n4888# 0.538783f
C91 drain_left.n4 a_n1598_n4888# 4.92945f
C92 drain_left.t3 a_n1598_n4888# 0.538783f
C93 drain_left.t0 a_n1598_n4888# 0.538783f
C94 drain_left.n5 a_n1598_n4888# 4.92566f
C95 drain_left.n6 a_n1598_n4888# 0.823936f
C96 drain_left.t7 a_n1598_n4888# 0.538783f
C97 drain_left.t5 a_n1598_n4888# 0.538783f
C98 drain_left.n7 a_n1598_n4888# 4.92566f
C99 drain_left.n8 a_n1598_n4888# 0.690749f
C100 source.t18 a_n1598_n4888# 4.73379f
C101 source.n0 a_n1598_n4888# 2.01344f
C102 source.t13 a_n1598_n4888# 0.414213f
C103 source.t16 a_n1598_n4888# 0.414213f
C104 source.n1 a_n1598_n4888# 3.70324f
C105 source.n2 a_n1598_n4888# 0.360853f
C106 source.t15 a_n1598_n4888# 0.414213f
C107 source.t20 a_n1598_n4888# 0.414213f
C108 source.n3 a_n1598_n4888# 3.70324f
C109 source.n4 a_n1598_n4888# 0.360853f
C110 source.t23 a_n1598_n4888# 4.7338f
C111 source.n5 a_n1598_n4888# 0.453785f
C112 source.t0 a_n1598_n4888# 4.7338f
C113 source.n6 a_n1598_n4888# 0.453785f
C114 source.t6 a_n1598_n4888# 0.414213f
C115 source.t5 a_n1598_n4888# 0.414213f
C116 source.n7 a_n1598_n4888# 3.70324f
C117 source.n8 a_n1598_n4888# 0.360853f
C118 source.t1 a_n1598_n4888# 0.414213f
C119 source.t8 a_n1598_n4888# 0.414213f
C120 source.n9 a_n1598_n4888# 3.70324f
C121 source.n10 a_n1598_n4888# 0.360853f
C122 source.t11 a_n1598_n4888# 4.7338f
C123 source.n11 a_n1598_n4888# 2.47788f
C124 source.t14 a_n1598_n4888# 4.73377f
C125 source.n12 a_n1598_n4888# 2.47791f
C126 source.t21 a_n1598_n4888# 0.414213f
C127 source.t22 a_n1598_n4888# 0.414213f
C128 source.n13 a_n1598_n4888# 3.70325f
C129 source.n14 a_n1598_n4888# 0.360846f
C130 source.t17 a_n1598_n4888# 0.414213f
C131 source.t19 a_n1598_n4888# 0.414213f
C132 source.n15 a_n1598_n4888# 3.70325f
C133 source.n16 a_n1598_n4888# 0.360846f
C134 source.t12 a_n1598_n4888# 4.73377f
C135 source.n17 a_n1598_n4888# 0.453811f
C136 source.t4 a_n1598_n4888# 4.73377f
C137 source.n18 a_n1598_n4888# 0.453811f
C138 source.t2 a_n1598_n4888# 0.414213f
C139 source.t3 a_n1598_n4888# 0.414213f
C140 source.n19 a_n1598_n4888# 3.70325f
C141 source.n20 a_n1598_n4888# 0.360846f
C142 source.t10 a_n1598_n4888# 0.414213f
C143 source.t7 a_n1598_n4888# 0.414213f
C144 source.n21 a_n1598_n4888# 3.70325f
C145 source.n22 a_n1598_n4888# 0.360846f
C146 source.t9 a_n1598_n4888# 4.73377f
C147 source.n23 a_n1598_n4888# 0.601757f
C148 source.n24 a_n1598_n4888# 2.35925f
C149 plus.n0 a_n1598_n4888# 0.053087f
C150 plus.t4 a_n1598_n4888# 0.897113f
C151 plus.t11 a_n1598_n4888# 0.897113f
C152 plus.n1 a_n1598_n4888# 0.019738f
C153 plus.t2 a_n1598_n4888# 0.906219f
C154 plus.n2 a_n1598_n4888# 0.350186f
C155 plus.t5 a_n1598_n4888# 0.897113f
C156 plus.n3 a_n1598_n4888# 0.333256f
C157 plus.t8 a_n1598_n4888# 0.897113f
C158 plus.n4 a_n1598_n4888# 0.333256f
C159 plus.n5 a_n1598_n4888# 0.021866f
C160 plus.n6 a_n1598_n4888# 0.120823f
C161 plus.n7 a_n1598_n4888# 0.053087f
C162 plus.n8 a_n1598_n4888# 0.053087f
C163 plus.n9 a_n1598_n4888# 0.019738f
C164 plus.n10 a_n1598_n4888# 0.333256f
C165 plus.n11 a_n1598_n4888# 0.021866f
C166 plus.n12 a_n1598_n4888# 0.333256f
C167 plus.t6 a_n1598_n4888# 0.906219f
C168 plus.n13 a_n1598_n4888# 0.350107f
C169 plus.n14 a_n1598_n4888# 0.80754f
C170 plus.n15 a_n1598_n4888# 0.053087f
C171 plus.t10 a_n1598_n4888# 0.906219f
C172 plus.t3 a_n1598_n4888# 0.897113f
C173 plus.t9 a_n1598_n4888# 0.897113f
C174 plus.n16 a_n1598_n4888# 0.019738f
C175 plus.t0 a_n1598_n4888# 0.906219f
C176 plus.n17 a_n1598_n4888# 0.350186f
C177 plus.t1 a_n1598_n4888# 0.897113f
C178 plus.n18 a_n1598_n4888# 0.333256f
C179 plus.t7 a_n1598_n4888# 0.897113f
C180 plus.n19 a_n1598_n4888# 0.333256f
C181 plus.n20 a_n1598_n4888# 0.021866f
C182 plus.n21 a_n1598_n4888# 0.120823f
C183 plus.n22 a_n1598_n4888# 0.053087f
C184 plus.n23 a_n1598_n4888# 0.053087f
C185 plus.n24 a_n1598_n4888# 0.019738f
C186 plus.n25 a_n1598_n4888# 0.333256f
C187 plus.n26 a_n1598_n4888# 0.021866f
C188 plus.n27 a_n1598_n4888# 0.333256f
C189 plus.n28 a_n1598_n4888# 0.350107f
C190 plus.n29 a_n1598_n4888# 1.80468f
.ends

