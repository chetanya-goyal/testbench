* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.78 ps=4.78 w=2 l=0.6
X1 drain_left.t1 plus.t0 source.t1 a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.78 ps=4.78 w=2 l=0.6
X2 drain_left.t0 plus.t1 source.t0 a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.78 ps=4.78 w=2 l=0.6
X3 a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X4 a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X5 a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X6 a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X7 drain_right.t0 minus.t1 source.t3 a_n1088_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.78 ps=4.78 w=2 l=0.6
R0 minus.n0 minus.t0 332.846
R1 minus.n0 minus.t1 313.664
R2 minus minus.n0 0.188
R3 source.n26 source.n24 289.615
R4 source.n18 source.n16 289.615
R5 source.n2 source.n0 289.615
R6 source.n10 source.n8 289.615
R7 source.n27 source.n26 185
R8 source.n19 source.n18 185
R9 source.n3 source.n2 185
R10 source.n11 source.n10 185
R11 source.t3 source.n25 167.117
R12 source.t0 source.n17 167.117
R13 source.t1 source.n1 167.117
R14 source.t2 source.n9 167.117
R15 source.n26 source.t3 52.3082
R16 source.n18 source.t0 52.3082
R17 source.n2 source.t1 52.3082
R18 source.n10 source.t2 52.3082
R19 source.n31 source.n30 31.4096
R20 source.n23 source.n22 31.4096
R21 source.n7 source.n6 31.4096
R22 source.n15 source.n14 31.4096
R23 source.n23 source.n15 15.3306
R24 source.n27 source.n25 9.71174
R25 source.n19 source.n17 9.71174
R26 source.n3 source.n1 9.71174
R27 source.n11 source.n9 9.71174
R28 source.n30 source.n29 9.45567
R29 source.n22 source.n21 9.45567
R30 source.n6 source.n5 9.45567
R31 source.n14 source.n13 9.45567
R32 source.n29 source.n28 9.3005
R33 source.n21 source.n20 9.3005
R34 source.n5 source.n4 9.3005
R35 source.n13 source.n12 9.3005
R36 source.n32 source.n7 8.86505
R37 source.n30 source.n24 8.14595
R38 source.n22 source.n16 8.14595
R39 source.n6 source.n0 8.14595
R40 source.n14 source.n8 8.14595
R41 source.n28 source.n27 7.3702
R42 source.n20 source.n19 7.3702
R43 source.n4 source.n3 7.3702
R44 source.n12 source.n11 7.3702
R45 source.n28 source.n24 5.81868
R46 source.n20 source.n16 5.81868
R47 source.n4 source.n0 5.81868
R48 source.n12 source.n8 5.81868
R49 source.n32 source.n31 5.66429
R50 source.n29 source.n25 3.44771
R51 source.n21 source.n17 3.44771
R52 source.n5 source.n1 3.44771
R53 source.n13 source.n9 3.44771
R54 source.n15 source.n7 0.87119
R55 source.n31 source.n23 0.87119
R56 source source.n32 0.188
R57 drain_right.n2 drain_right.n0 289.615
R58 drain_right.n9 drain_right.n7 289.615
R59 drain_right.n3 drain_right.n2 185
R60 drain_right.n10 drain_right.n9 185
R61 drain_right.t0 drain_right.n1 167.117
R62 drain_right.t1 drain_right.n8 167.117
R63 drain_right drain_right.n6 68.4884
R64 drain_right drain_right.n13 54.142
R65 drain_right.n2 drain_right.t0 52.3082
R66 drain_right.n9 drain_right.t1 52.3082
R67 drain_right.n3 drain_right.n1 9.71174
R68 drain_right.n10 drain_right.n8 9.71174
R69 drain_right.n6 drain_right.n5 9.45567
R70 drain_right.n13 drain_right.n12 9.45567
R71 drain_right.n5 drain_right.n4 9.3005
R72 drain_right.n12 drain_right.n11 9.3005
R73 drain_right.n6 drain_right.n0 8.14595
R74 drain_right.n13 drain_right.n7 8.14595
R75 drain_right.n4 drain_right.n3 7.3702
R76 drain_right.n11 drain_right.n10 7.3702
R77 drain_right.n4 drain_right.n0 5.81868
R78 drain_right.n11 drain_right.n7 5.81868
R79 drain_right.n5 drain_right.n1 3.44771
R80 drain_right.n12 drain_right.n8 3.44771
R81 plus plus.t1 330.514
R82 plus plus.t0 315.521
R83 drain_left.n2 drain_left.n0 289.615
R84 drain_left.n9 drain_left.n7 289.615
R85 drain_left.n3 drain_left.n2 185
R86 drain_left.n10 drain_left.n9 185
R87 drain_left.t0 drain_left.n1 167.117
R88 drain_left.t1 drain_left.n8 167.117
R89 drain_left drain_left.n6 69.0416
R90 drain_left drain_left.n13 54.5428
R91 drain_left.n2 drain_left.t0 52.3082
R92 drain_left.n9 drain_left.t1 52.3082
R93 drain_left.n3 drain_left.n1 9.71174
R94 drain_left.n10 drain_left.n8 9.71174
R95 drain_left.n6 drain_left.n5 9.45567
R96 drain_left.n13 drain_left.n12 9.45567
R97 drain_left.n5 drain_left.n4 9.3005
R98 drain_left.n12 drain_left.n11 9.3005
R99 drain_left.n6 drain_left.n0 8.14595
R100 drain_left.n13 drain_left.n7 8.14595
R101 drain_left.n4 drain_left.n3 7.3702
R102 drain_left.n11 drain_left.n10 7.3702
R103 drain_left.n4 drain_left.n0 5.81868
R104 drain_left.n11 drain_left.n7 5.81868
R105 drain_left.n5 drain_left.n1 3.44771
R106 drain_left.n12 drain_left.n8 3.44771
C0 source minus 0.532395f
C1 plus drain_right 0.262111f
C2 plus minus 2.65252f
C3 source drain_left 2.03924f
C4 drain_right minus 0.514645f
C5 plus drain_left 0.614549f
C6 source plus 0.546446f
C7 drain_right drain_left 0.448937f
C8 source drain_right 2.03705f
C9 drain_left minus 0.178042f
C10 drain_right a_n1088_n1292# 3.04744f
C11 drain_left a_n1088_n1292# 3.16298f
C12 source a_n1088_n1292# 2.350568f
C13 minus a_n1088_n1292# 3.241436f
C14 plus a_n1088_n1292# 5.25589f
C15 drain_left.n0 a_n1088_n1292# 0.023639f
C16 drain_left.n1 a_n1088_n1292# 0.052304f
C17 drain_left.t0 a_n1088_n1292# 0.039251f
C18 drain_left.n2 a_n1088_n1292# 0.040935f
C19 drain_left.n3 a_n1088_n1292# 0.013196f
C20 drain_left.n4 a_n1088_n1292# 0.008703f
C21 drain_left.n5 a_n1088_n1292# 0.115291f
C22 drain_left.n6 a_n1088_n1292# 0.143427f
C23 drain_left.n7 a_n1088_n1292# 0.023639f
C24 drain_left.n8 a_n1088_n1292# 0.052304f
C25 drain_left.t1 a_n1088_n1292# 0.039251f
C26 drain_left.n9 a_n1088_n1292# 0.040935f
C27 drain_left.n10 a_n1088_n1292# 0.013196f
C28 drain_left.n11 a_n1088_n1292# 0.008703f
C29 drain_left.n12 a_n1088_n1292# 0.115291f
C30 drain_left.n13 a_n1088_n1292# 0.062398f
C31 plus.t0 a_n1088_n1292# 0.227176f
C32 plus.t1 a_n1088_n1292# 0.280198f
C33 drain_right.n0 a_n1088_n1292# 0.024412f
C34 drain_right.n1 a_n1088_n1292# 0.054015f
C35 drain_right.t0 a_n1088_n1292# 0.040536f
C36 drain_right.n2 a_n1088_n1292# 0.042274f
C37 drain_right.n3 a_n1088_n1292# 0.013628f
C38 drain_right.n4 a_n1088_n1292# 0.008988f
C39 drain_right.n5 a_n1088_n1292# 0.119063f
C40 drain_right.n6 a_n1088_n1292# 0.136294f
C41 drain_right.n7 a_n1088_n1292# 0.024412f
C42 drain_right.n8 a_n1088_n1292# 0.054015f
C43 drain_right.t1 a_n1088_n1292# 0.040536f
C44 drain_right.n9 a_n1088_n1292# 0.042274f
C45 drain_right.n10 a_n1088_n1292# 0.013628f
C46 drain_right.n11 a_n1088_n1292# 0.008988f
C47 drain_right.n12 a_n1088_n1292# 0.119063f
C48 drain_right.n13 a_n1088_n1292# 0.064238f
C49 source.n0 a_n1088_n1292# 0.030424f
C50 source.n1 a_n1088_n1292# 0.067316f
C51 source.t1 a_n1088_n1292# 0.050517f
C52 source.n2 a_n1088_n1292# 0.052684f
C53 source.n3 a_n1088_n1292# 0.016983f
C54 source.n4 a_n1088_n1292# 0.011201f
C55 source.n5 a_n1088_n1292# 0.148381f
C56 source.n6 a_n1088_n1292# 0.033351f
C57 source.n7 a_n1088_n1292# 0.350962f
C58 source.n8 a_n1088_n1292# 0.030424f
C59 source.n9 a_n1088_n1292# 0.067316f
C60 source.t2 a_n1088_n1292# 0.050517f
C61 source.n10 a_n1088_n1292# 0.052684f
C62 source.n11 a_n1088_n1292# 0.016983f
C63 source.n12 a_n1088_n1292# 0.011201f
C64 source.n13 a_n1088_n1292# 0.148381f
C65 source.n14 a_n1088_n1292# 0.033351f
C66 source.n15 a_n1088_n1292# 0.603587f
C67 source.n16 a_n1088_n1292# 0.030424f
C68 source.n17 a_n1088_n1292# 0.067316f
C69 source.t0 a_n1088_n1292# 0.050517f
C70 source.n18 a_n1088_n1292# 0.052684f
C71 source.n19 a_n1088_n1292# 0.016983f
C72 source.n20 a_n1088_n1292# 0.011201f
C73 source.n21 a_n1088_n1292# 0.148381f
C74 source.n22 a_n1088_n1292# 0.033351f
C75 source.n23 a_n1088_n1292# 0.603587f
C76 source.n24 a_n1088_n1292# 0.030424f
C77 source.n25 a_n1088_n1292# 0.067316f
C78 source.t3 a_n1088_n1292# 0.050517f
C79 source.n26 a_n1088_n1292# 0.052684f
C80 source.n27 a_n1088_n1292# 0.016983f
C81 source.n28 a_n1088_n1292# 0.011201f
C82 source.n29 a_n1088_n1292# 0.148381f
C83 source.n30 a_n1088_n1292# 0.033351f
C84 source.n31 a_n1088_n1292# 0.238627f
C85 source.n32 a_n1088_n1292# 0.524716f
C86 minus.t0 a_n1088_n1292# 0.279171f
C87 minus.t1 a_n1088_n1292# 0.217391f
C88 minus.n0 a_n1088_n1292# 2.17575f
.ends

