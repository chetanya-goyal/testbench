* NGSPICE file created from diffpair27.ext - technology: sky130A

.subckt diffpair27 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t16 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 drain_left.t14 plus.t1 source.t29 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X2 source.t14 minus.t0 drain_right.t15 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 source.t9 minus.t1 drain_right.t14 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X4 a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X5 drain_left.t13 plus.t2 source.t26 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X6 source.t12 minus.t2 drain_right.t13 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X7 a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X8 source.t6 minus.t3 drain_right.t12 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X9 source.t13 minus.t4 drain_right.t11 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X10 source.t21 plus.t3 drain_left.t12 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X11 drain_right.t10 minus.t5 source.t15 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X12 source.t11 minus.t6 drain_right.t9 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X13 source.t2 minus.t7 drain_right.t8 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X14 source.t3 minus.t8 drain_right.t7 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X15 drain_right.t6 minus.t9 source.t5 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X16 source.t19 plus.t4 drain_left.t11 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X17 source.t17 plus.t5 drain_left.t10 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X18 source.t18 plus.t6 drain_left.t9 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X19 source.t31 plus.t7 drain_left.t8 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X20 a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X21 drain_left.t7 plus.t8 source.t22 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X22 drain_left.t6 plus.t9 source.t27 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X23 drain_right.t5 minus.t10 source.t8 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X24 a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X25 drain_left.t5 plus.t10 source.t24 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X26 drain_right.t4 minus.t11 source.t10 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X27 drain_left.t4 plus.t11 source.t23 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X28 source.t28 plus.t12 drain_left.t3 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X29 source.t25 plus.t13 drain_left.t2 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X30 source.t30 plus.t14 drain_left.t1 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X31 drain_right.t3 minus.t12 source.t0 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X32 drain_right.t2 minus.t13 source.t1 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X33 drain_right.t1 minus.t14 source.t4 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X34 drain_left.t0 plus.t15 source.t20 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X35 drain_right.t0 minus.t15 source.t7 a_n1760_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
R0 plus.n4 plus.t3 262.618
R1 plus.n19 plus.t2 262.618
R2 plus.n25 plus.t9 262.618
R3 plus.n40 plus.t13 262.618
R4 plus.n5 plus.t1 221.72
R5 plus.n3 plus.t7 221.72
R6 plus.n10 plus.t0 221.72
R7 plus.n1 plus.t6 221.72
R8 plus.n16 plus.t15 221.72
R9 plus.n18 plus.t5 221.72
R10 plus.n26 plus.t4 221.72
R11 plus.n24 plus.t11 221.72
R12 plus.n31 plus.t14 221.72
R13 plus.n22 plus.t8 221.72
R14 plus.n37 plus.t12 221.72
R15 plus.n39 plus.t10 221.72
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus.n6 plus.n5 29.2126
R47 plus.n18 plus.n17 29.2126
R48 plus.n39 plus.n38 29.2126
R49 plus.n27 plus.n26 29.2126
R50 plus plus.n41 25.4687
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 7.94368
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n0 source.t26 243.255
R73 source.n7 source.t21 243.255
R74 source.n8 source.t10 243.255
R75 source.n15 source.t2 243.255
R76 source.n31 source.t15 243.254
R77 source.n24 source.t13 243.254
R78 source.n23 source.t27 243.254
R79 source.n16 source.t25 243.254
R80 source.n2 source.n1 223.454
R81 source.n4 source.n3 223.454
R82 source.n6 source.n5 223.454
R83 source.n10 source.n9 223.454
R84 source.n12 source.n11 223.454
R85 source.n14 source.n13 223.454
R86 source.n30 source.n29 223.453
R87 source.n28 source.n27 223.453
R88 source.n26 source.n25 223.453
R89 source.n22 source.n21 223.453
R90 source.n20 source.n19 223.453
R91 source.n18 source.n17 223.453
R92 source.n29 source.t5 19.8005
R93 source.n29 source.t11 19.8005
R94 source.n27 source.t7 19.8005
R95 source.n27 source.t6 19.8005
R96 source.n25 source.t4 19.8005
R97 source.n25 source.t14 19.8005
R98 source.n21 source.t23 19.8005
R99 source.n21 source.t19 19.8005
R100 source.n19 source.t22 19.8005
R101 source.n19 source.t30 19.8005
R102 source.n17 source.t24 19.8005
R103 source.n17 source.t28 19.8005
R104 source.n1 source.t20 19.8005
R105 source.n1 source.t17 19.8005
R106 source.n3 source.t16 19.8005
R107 source.n3 source.t18 19.8005
R108 source.n5 source.t29 19.8005
R109 source.n5 source.t31 19.8005
R110 source.n9 source.t8 19.8005
R111 source.n9 source.t12 19.8005
R112 source.n11 source.t0 19.8005
R113 source.n11 source.t9 19.8005
R114 source.n13 source.t1 19.8005
R115 source.n13 source.t3 19.8005
R116 source.n16 source.n15 13.4544
R117 source.n32 source.n0 7.94146
R118 source.n32 source.n31 5.51343
R119 source.n15 source.n14 0.5005
R120 source.n14 source.n12 0.5005
R121 source.n12 source.n10 0.5005
R122 source.n10 source.n8 0.5005
R123 source.n7 source.n6 0.5005
R124 source.n6 source.n4 0.5005
R125 source.n4 source.n2 0.5005
R126 source.n2 source.n0 0.5005
R127 source.n18 source.n16 0.5005
R128 source.n20 source.n18 0.5005
R129 source.n22 source.n20 0.5005
R130 source.n23 source.n22 0.5005
R131 source.n26 source.n24 0.5005
R132 source.n28 source.n26 0.5005
R133 source.n30 source.n28 0.5005
R134 source.n31 source.n30 0.5005
R135 source.n8 source.n7 0.470328
R136 source.n24 source.n23 0.470328
R137 source source.n32 0.188
R138 drain_left.n9 drain_left.n7 240.632
R139 drain_left.n5 drain_left.n3 240.631
R140 drain_left.n2 drain_left.n0 240.631
R141 drain_left.n13 drain_left.n12 240.132
R142 drain_left.n11 drain_left.n10 240.132
R143 drain_left.n9 drain_left.n8 240.132
R144 drain_left.n5 drain_left.n4 240.131
R145 drain_left.n2 drain_left.n1 240.131
R146 drain_left drain_left.n6 22.2837
R147 drain_left.n3 drain_left.t11 19.8005
R148 drain_left.n3 drain_left.t6 19.8005
R149 drain_left.n4 drain_left.t1 19.8005
R150 drain_left.n4 drain_left.t4 19.8005
R151 drain_left.n1 drain_left.t3 19.8005
R152 drain_left.n1 drain_left.t7 19.8005
R153 drain_left.n0 drain_left.t2 19.8005
R154 drain_left.n0 drain_left.t5 19.8005
R155 drain_left.n12 drain_left.t10 19.8005
R156 drain_left.n12 drain_left.t13 19.8005
R157 drain_left.n10 drain_left.t9 19.8005
R158 drain_left.n10 drain_left.t0 19.8005
R159 drain_left.n8 drain_left.t8 19.8005
R160 drain_left.n8 drain_left.t15 19.8005
R161 drain_left.n7 drain_left.t12 19.8005
R162 drain_left.n7 drain_left.t14 19.8005
R163 drain_left drain_left.n13 6.15322
R164 drain_left.n11 drain_left.n9 0.5005
R165 drain_left.n13 drain_left.n11 0.5005
R166 drain_left.n6 drain_left.n5 0.195154
R167 drain_left.n6 drain_left.n2 0.195154
R168 minus.n19 minus.t7 262.618
R169 minus.n4 minus.t11 262.618
R170 minus.n40 minus.t5 262.618
R171 minus.n25 minus.t4 262.618
R172 minus.n18 minus.t13 221.72
R173 minus.n16 minus.t8 221.72
R174 minus.n1 minus.t12 221.72
R175 minus.n10 minus.t1 221.72
R176 minus.n3 minus.t10 221.72
R177 minus.n5 minus.t2 221.72
R178 minus.n39 minus.t6 221.72
R179 minus.n37 minus.t9 221.72
R180 minus.n22 minus.t3 221.72
R181 minus.n31 minus.t15 221.72
R182 minus.n24 minus.t0 221.72
R183 minus.n26 minus.t14 221.72
R184 minus.n7 minus.n4 161.489
R185 minus.n28 minus.n25 161.489
R186 minus.n20 minus.n19 161.3
R187 minus.n17 minus.n0 161.3
R188 minus.n15 minus.n14 161.3
R189 minus.n13 minus.n12 161.3
R190 minus.n11 minus.n2 161.3
R191 minus.n9 minus.n8 161.3
R192 minus.n7 minus.n6 161.3
R193 minus.n41 minus.n40 161.3
R194 minus.n38 minus.n21 161.3
R195 minus.n36 minus.n35 161.3
R196 minus.n34 minus.n33 161.3
R197 minus.n32 minus.n23 161.3
R198 minus.n30 minus.n29 161.3
R199 minus.n28 minus.n27 161.3
R200 minus.n12 minus.n11 73.0308
R201 minus.n33 minus.n32 73.0308
R202 minus.n15 minus.n1 67.1884
R203 minus.n10 minus.n9 67.1884
R204 minus.n31 minus.n30 67.1884
R205 minus.n36 minus.n22 67.1884
R206 minus.n17 minus.n16 55.5035
R207 minus.n6 minus.n3 55.5035
R208 minus.n27 minus.n24 55.5035
R209 minus.n38 minus.n37 55.5035
R210 minus.n19 minus.n18 43.8187
R211 minus.n5 minus.n4 43.8187
R212 minus.n26 minus.n25 43.8187
R213 minus.n40 minus.n39 43.8187
R214 minus.n18 minus.n17 29.2126
R215 minus.n6 minus.n5 29.2126
R216 minus.n27 minus.n26 29.2126
R217 minus.n39 minus.n38 29.2126
R218 minus.n42 minus.n20 27.421
R219 minus.n16 minus.n15 17.5278
R220 minus.n9 minus.n3 17.5278
R221 minus.n30 minus.n24 17.5278
R222 minus.n37 minus.n36 17.5278
R223 minus.n42 minus.n41 6.46641
R224 minus.n12 minus.n1 5.84292
R225 minus.n11 minus.n10 5.84292
R226 minus.n32 minus.n31 5.84292
R227 minus.n33 minus.n22 5.84292
R228 minus.n20 minus.n0 0.189894
R229 minus.n14 minus.n0 0.189894
R230 minus.n14 minus.n13 0.189894
R231 minus.n13 minus.n2 0.189894
R232 minus.n8 minus.n2 0.189894
R233 minus.n8 minus.n7 0.189894
R234 minus.n29 minus.n28 0.189894
R235 minus.n29 minus.n23 0.189894
R236 minus.n34 minus.n23 0.189894
R237 minus.n35 minus.n34 0.189894
R238 minus.n35 minus.n21 0.189894
R239 minus.n41 minus.n21 0.189894
R240 minus minus.n42 0.188
R241 drain_right.n9 drain_right.n7 240.632
R242 drain_right.n5 drain_right.n3 240.631
R243 drain_right.n2 drain_right.n0 240.631
R244 drain_right.n9 drain_right.n8 240.132
R245 drain_right.n11 drain_right.n10 240.132
R246 drain_right.n13 drain_right.n12 240.132
R247 drain_right.n5 drain_right.n4 240.131
R248 drain_right.n2 drain_right.n1 240.131
R249 drain_right drain_right.n6 21.7305
R250 drain_right.n3 drain_right.t9 19.8005
R251 drain_right.n3 drain_right.t10 19.8005
R252 drain_right.n4 drain_right.t12 19.8005
R253 drain_right.n4 drain_right.t6 19.8005
R254 drain_right.n1 drain_right.t15 19.8005
R255 drain_right.n1 drain_right.t0 19.8005
R256 drain_right.n0 drain_right.t11 19.8005
R257 drain_right.n0 drain_right.t1 19.8005
R258 drain_right.n7 drain_right.t13 19.8005
R259 drain_right.n7 drain_right.t4 19.8005
R260 drain_right.n8 drain_right.t14 19.8005
R261 drain_right.n8 drain_right.t5 19.8005
R262 drain_right.n10 drain_right.t7 19.8005
R263 drain_right.n10 drain_right.t3 19.8005
R264 drain_right.n12 drain_right.t8 19.8005
R265 drain_right.n12 drain_right.t2 19.8005
R266 drain_right drain_right.n13 6.15322
R267 drain_right.n13 drain_right.n11 0.5005
R268 drain_right.n11 drain_right.n9 0.5005
R269 drain_right.n6 drain_right.n5 0.195154
R270 drain_right.n6 drain_right.n2 0.195154
C0 drain_left minus 0.178502f
C1 drain_right plus 0.332889f
C2 minus plus 3.32274f
C3 drain_left plus 1.06848f
C4 drain_right source 5.29583f
C5 source minus 1.14512f
C6 source drain_left 5.29588f
C7 drain_right minus 0.898215f
C8 source plus 1.15898f
C9 drain_right drain_left 0.897326f
C10 drain_right a_n1760_n1088# 3.63115f
C11 drain_left a_n1760_n1088# 3.86886f
C12 source a_n1760_n1088# 2.499506f
C13 minus a_n1760_n1088# 5.952677f
C14 plus a_n1760_n1088# 6.626657f
C15 drain_right.t11 a_n1760_n1088# 0.021066f
C16 drain_right.t1 a_n1760_n1088# 0.021066f
C17 drain_right.n0 a_n1760_n1088# 0.082444f
C18 drain_right.t15 a_n1760_n1088# 0.021066f
C19 drain_right.t0 a_n1760_n1088# 0.021066f
C20 drain_right.n1 a_n1760_n1088# 0.081856f
C21 drain_right.n2 a_n1760_n1088# 0.531737f
C22 drain_right.t9 a_n1760_n1088# 0.021066f
C23 drain_right.t10 a_n1760_n1088# 0.021066f
C24 drain_right.n3 a_n1760_n1088# 0.082444f
C25 drain_right.t12 a_n1760_n1088# 0.021066f
C26 drain_right.t6 a_n1760_n1088# 0.021066f
C27 drain_right.n4 a_n1760_n1088# 0.081856f
C28 drain_right.n5 a_n1760_n1088# 0.531737f
C29 drain_right.n6 a_n1760_n1088# 0.639871f
C30 drain_right.t13 a_n1760_n1088# 0.021066f
C31 drain_right.t4 a_n1760_n1088# 0.021066f
C32 drain_right.n7 a_n1760_n1088# 0.082444f
C33 drain_right.t14 a_n1760_n1088# 0.021066f
C34 drain_right.t5 a_n1760_n1088# 0.021066f
C35 drain_right.n8 a_n1760_n1088# 0.081856f
C36 drain_right.n9 a_n1760_n1088# 0.55479f
C37 drain_right.t7 a_n1760_n1088# 0.021066f
C38 drain_right.t3 a_n1760_n1088# 0.021066f
C39 drain_right.n10 a_n1760_n1088# 0.081856f
C40 drain_right.n11 a_n1760_n1088# 0.272321f
C41 drain_right.t8 a_n1760_n1088# 0.021066f
C42 drain_right.t2 a_n1760_n1088# 0.021066f
C43 drain_right.n12 a_n1760_n1088# 0.081856f
C44 drain_right.n13 a_n1760_n1088# 0.492365f
C45 minus.n0 a_n1760_n1088# 0.032005f
C46 minus.t7 a_n1760_n1088# 0.028971f
C47 minus.t13 a_n1760_n1088# 0.024666f
C48 minus.t8 a_n1760_n1088# 0.024666f
C49 minus.t12 a_n1760_n1088# 0.024666f
C50 minus.n1 a_n1760_n1088# 0.027057f
C51 minus.n2 a_n1760_n1088# 0.032005f
C52 minus.t1 a_n1760_n1088# 0.024666f
C53 minus.t10 a_n1760_n1088# 0.024666f
C54 minus.n3 a_n1760_n1088# 0.027057f
C55 minus.t11 a_n1760_n1088# 0.028971f
C56 minus.n4 a_n1760_n1088# 0.035584f
C57 minus.t2 a_n1760_n1088# 0.024666f
C58 minus.n5 a_n1760_n1088# 0.027057f
C59 minus.n6 a_n1760_n1088# 0.012196f
C60 minus.n7 a_n1760_n1088# 0.070082f
C61 minus.n8 a_n1760_n1088# 0.032005f
C62 minus.n9 a_n1760_n1088# 0.012196f
C63 minus.n10 a_n1760_n1088# 0.027057f
C64 minus.n11 a_n1760_n1088# 0.011406f
C65 minus.n12 a_n1760_n1088# 0.011406f
C66 minus.n13 a_n1760_n1088# 0.032005f
C67 minus.n14 a_n1760_n1088# 0.032005f
C68 minus.n15 a_n1760_n1088# 0.012196f
C69 minus.n16 a_n1760_n1088# 0.027057f
C70 minus.n17 a_n1760_n1088# 0.012196f
C71 minus.n18 a_n1760_n1088# 0.027057f
C72 minus.n19 a_n1760_n1088# 0.035539f
C73 minus.n20 a_n1760_n1088# 0.710413f
C74 minus.n21 a_n1760_n1088# 0.032005f
C75 minus.t6 a_n1760_n1088# 0.024666f
C76 minus.t9 a_n1760_n1088# 0.024666f
C77 minus.t3 a_n1760_n1088# 0.024666f
C78 minus.n22 a_n1760_n1088# 0.027057f
C79 minus.n23 a_n1760_n1088# 0.032005f
C80 minus.t15 a_n1760_n1088# 0.024666f
C81 minus.t0 a_n1760_n1088# 0.024666f
C82 minus.n24 a_n1760_n1088# 0.027057f
C83 minus.t4 a_n1760_n1088# 0.028971f
C84 minus.n25 a_n1760_n1088# 0.035584f
C85 minus.t14 a_n1760_n1088# 0.024666f
C86 minus.n26 a_n1760_n1088# 0.027057f
C87 minus.n27 a_n1760_n1088# 0.012196f
C88 minus.n28 a_n1760_n1088# 0.070082f
C89 minus.n29 a_n1760_n1088# 0.032005f
C90 minus.n30 a_n1760_n1088# 0.012196f
C91 minus.n31 a_n1760_n1088# 0.027057f
C92 minus.n32 a_n1760_n1088# 0.011406f
C93 minus.n33 a_n1760_n1088# 0.011406f
C94 minus.n34 a_n1760_n1088# 0.032005f
C95 minus.n35 a_n1760_n1088# 0.032005f
C96 minus.n36 a_n1760_n1088# 0.012196f
C97 minus.n37 a_n1760_n1088# 0.027057f
C98 minus.n38 a_n1760_n1088# 0.012196f
C99 minus.n39 a_n1760_n1088# 0.027057f
C100 minus.t5 a_n1760_n1088# 0.028971f
C101 minus.n40 a_n1760_n1088# 0.035539f
C102 minus.n41 a_n1760_n1088# 0.206704f
C103 minus.n42 a_n1760_n1088# 0.879651f
C104 drain_left.t2 a_n1760_n1088# 0.02066f
C105 drain_left.t5 a_n1760_n1088# 0.02066f
C106 drain_left.n0 a_n1760_n1088# 0.080854f
C107 drain_left.t3 a_n1760_n1088# 0.02066f
C108 drain_left.t7 a_n1760_n1088# 0.02066f
C109 drain_left.n1 a_n1760_n1088# 0.080277f
C110 drain_left.n2 a_n1760_n1088# 0.521476f
C111 drain_left.t11 a_n1760_n1088# 0.02066f
C112 drain_left.t6 a_n1760_n1088# 0.02066f
C113 drain_left.n3 a_n1760_n1088# 0.080854f
C114 drain_left.t1 a_n1760_n1088# 0.02066f
C115 drain_left.t4 a_n1760_n1088# 0.02066f
C116 drain_left.n4 a_n1760_n1088# 0.080277f
C117 drain_left.n5 a_n1760_n1088# 0.521476f
C118 drain_left.n6 a_n1760_n1088# 0.678081f
C119 drain_left.t12 a_n1760_n1088# 0.02066f
C120 drain_left.t14 a_n1760_n1088# 0.02066f
C121 drain_left.n7 a_n1760_n1088# 0.080854f
C122 drain_left.t8 a_n1760_n1088# 0.02066f
C123 drain_left.t15 a_n1760_n1088# 0.02066f
C124 drain_left.n8 a_n1760_n1088# 0.080277f
C125 drain_left.n9 a_n1760_n1088# 0.544085f
C126 drain_left.t9 a_n1760_n1088# 0.02066f
C127 drain_left.t0 a_n1760_n1088# 0.02066f
C128 drain_left.n10 a_n1760_n1088# 0.080277f
C129 drain_left.n11 a_n1760_n1088# 0.267066f
C130 drain_left.t10 a_n1760_n1088# 0.02066f
C131 drain_left.t13 a_n1760_n1088# 0.02066f
C132 drain_left.n12 a_n1760_n1088# 0.080277f
C133 drain_left.n13 a_n1760_n1088# 0.482864f
C134 source.t26 a_n1760_n1088# 0.135334f
C135 source.n0 a_n1760_n1088# 0.573441f
C136 source.t20 a_n1760_n1088# 0.024315f
C137 source.t17 a_n1760_n1088# 0.024315f
C138 source.n1 a_n1760_n1088# 0.078858f
C139 source.n2 a_n1760_n1088# 0.288123f
C140 source.t16 a_n1760_n1088# 0.024315f
C141 source.t18 a_n1760_n1088# 0.024315f
C142 source.n3 a_n1760_n1088# 0.078858f
C143 source.n4 a_n1760_n1088# 0.288123f
C144 source.t29 a_n1760_n1088# 0.024315f
C145 source.t31 a_n1760_n1088# 0.024315f
C146 source.n5 a_n1760_n1088# 0.078858f
C147 source.n6 a_n1760_n1088# 0.288123f
C148 source.t21 a_n1760_n1088# 0.135334f
C149 source.n7 a_n1760_n1088# 0.294968f
C150 source.t10 a_n1760_n1088# 0.135334f
C151 source.n8 a_n1760_n1088# 0.294968f
C152 source.t8 a_n1760_n1088# 0.024315f
C153 source.t12 a_n1760_n1088# 0.024315f
C154 source.n9 a_n1760_n1088# 0.078858f
C155 source.n10 a_n1760_n1088# 0.288123f
C156 source.t0 a_n1760_n1088# 0.024315f
C157 source.t9 a_n1760_n1088# 0.024315f
C158 source.n11 a_n1760_n1088# 0.078858f
C159 source.n12 a_n1760_n1088# 0.288123f
C160 source.t1 a_n1760_n1088# 0.024315f
C161 source.t3 a_n1760_n1088# 0.024315f
C162 source.n13 a_n1760_n1088# 0.078858f
C163 source.n14 a_n1760_n1088# 0.288123f
C164 source.t2 a_n1760_n1088# 0.135334f
C165 source.n15 a_n1760_n1088# 0.819112f
C166 source.t25 a_n1760_n1088# 0.135334f
C167 source.n16 a_n1760_n1088# 0.819112f
C168 source.t24 a_n1760_n1088# 0.024315f
C169 source.t28 a_n1760_n1088# 0.024315f
C170 source.n17 a_n1760_n1088# 0.078857f
C171 source.n18 a_n1760_n1088# 0.288123f
C172 source.t22 a_n1760_n1088# 0.024315f
C173 source.t30 a_n1760_n1088# 0.024315f
C174 source.n19 a_n1760_n1088# 0.078857f
C175 source.n20 a_n1760_n1088# 0.288123f
C176 source.t23 a_n1760_n1088# 0.024315f
C177 source.t19 a_n1760_n1088# 0.024315f
C178 source.n21 a_n1760_n1088# 0.078857f
C179 source.n22 a_n1760_n1088# 0.288123f
C180 source.t27 a_n1760_n1088# 0.135334f
C181 source.n23 a_n1760_n1088# 0.294969f
C182 source.t13 a_n1760_n1088# 0.135334f
C183 source.n24 a_n1760_n1088# 0.294969f
C184 source.t4 a_n1760_n1088# 0.024315f
C185 source.t14 a_n1760_n1088# 0.024315f
C186 source.n25 a_n1760_n1088# 0.078857f
C187 source.n26 a_n1760_n1088# 0.288123f
C188 source.t7 a_n1760_n1088# 0.024315f
C189 source.t6 a_n1760_n1088# 0.024315f
C190 source.n27 a_n1760_n1088# 0.078857f
C191 source.n28 a_n1760_n1088# 0.288123f
C192 source.t5 a_n1760_n1088# 0.024315f
C193 source.t11 a_n1760_n1088# 0.024315f
C194 source.n29 a_n1760_n1088# 0.078857f
C195 source.n30 a_n1760_n1088# 0.288123f
C196 source.t15 a_n1760_n1088# 0.135334f
C197 source.n31 a_n1760_n1088# 0.465242f
C198 source.n32 a_n1760_n1088# 0.621428f
C199 plus.n0 a_n1760_n1088# 0.032645f
C200 plus.t5 a_n1760_n1088# 0.025159f
C201 plus.t15 a_n1760_n1088# 0.025159f
C202 plus.t6 a_n1760_n1088# 0.025159f
C203 plus.n1 a_n1760_n1088# 0.027599f
C204 plus.n2 a_n1760_n1088# 0.032645f
C205 plus.t0 a_n1760_n1088# 0.025159f
C206 plus.t7 a_n1760_n1088# 0.025159f
C207 plus.n3 a_n1760_n1088# 0.027599f
C208 plus.t3 a_n1760_n1088# 0.029551f
C209 plus.n4 a_n1760_n1088# 0.036296f
C210 plus.t1 a_n1760_n1088# 0.025159f
C211 plus.n5 a_n1760_n1088# 0.027599f
C212 plus.n6 a_n1760_n1088# 0.01244f
C213 plus.n7 a_n1760_n1088# 0.071484f
C214 plus.n8 a_n1760_n1088# 0.032645f
C215 plus.n9 a_n1760_n1088# 0.01244f
C216 plus.n10 a_n1760_n1088# 0.027599f
C217 plus.n11 a_n1760_n1088# 0.011635f
C218 plus.n12 a_n1760_n1088# 0.011635f
C219 plus.n13 a_n1760_n1088# 0.032645f
C220 plus.n14 a_n1760_n1088# 0.032645f
C221 plus.n15 a_n1760_n1088# 0.01244f
C222 plus.n16 a_n1760_n1088# 0.027599f
C223 plus.n17 a_n1760_n1088# 0.01244f
C224 plus.n18 a_n1760_n1088# 0.027599f
C225 plus.t2 a_n1760_n1088# 0.029551f
C226 plus.n19 a_n1760_n1088# 0.03625f
C227 plus.n20 a_n1760_n1088# 0.22109f
C228 plus.n21 a_n1760_n1088# 0.032645f
C229 plus.t13 a_n1760_n1088# 0.029551f
C230 plus.t10 a_n1760_n1088# 0.025159f
C231 plus.t12 a_n1760_n1088# 0.025159f
C232 plus.t8 a_n1760_n1088# 0.025159f
C233 plus.n22 a_n1760_n1088# 0.027599f
C234 plus.n23 a_n1760_n1088# 0.032645f
C235 plus.t14 a_n1760_n1088# 0.025159f
C236 plus.t11 a_n1760_n1088# 0.025159f
C237 plus.n24 a_n1760_n1088# 0.027599f
C238 plus.t9 a_n1760_n1088# 0.029551f
C239 plus.n25 a_n1760_n1088# 0.036296f
C240 plus.t4 a_n1760_n1088# 0.025159f
C241 plus.n26 a_n1760_n1088# 0.027599f
C242 plus.n27 a_n1760_n1088# 0.01244f
C243 plus.n28 a_n1760_n1088# 0.071484f
C244 plus.n29 a_n1760_n1088# 0.032645f
C245 plus.n30 a_n1760_n1088# 0.01244f
C246 plus.n31 a_n1760_n1088# 0.027599f
C247 plus.n32 a_n1760_n1088# 0.011635f
C248 plus.n33 a_n1760_n1088# 0.011635f
C249 plus.n34 a_n1760_n1088# 0.032645f
C250 plus.n35 a_n1760_n1088# 0.032645f
C251 plus.n36 a_n1760_n1088# 0.01244f
C252 plus.n37 a_n1760_n1088# 0.027599f
C253 plus.n38 a_n1760_n1088# 0.01244f
C254 plus.n39 a_n1760_n1088# 0.027599f
C255 plus.n40 a_n1760_n1088# 0.03625f
C256 plus.n41 a_n1760_n1088# 0.703416f
.ends

