* NGSPICE file created from diffpair85.ext - technology: sky130A

.subckt diffpair85 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t11 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 source.t5 minus.t0 drain_right.t11 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 source.t8 minus.t1 drain_right.t10 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 source.t16 plus.t1 drain_left.t10 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X5 drain_left.t9 plus.t2 source.t13 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X6 a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X7 a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X8 drain_right.t9 minus.t2 source.t3 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X9 source.t7 minus.t3 drain_right.t8 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 source.t9 minus.t4 drain_right.t7 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 drain_right.t6 minus.t5 source.t0 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X12 drain_right.t5 minus.t6 source.t1 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 source.t14 plus.t3 drain_left.t8 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t2 minus.t7 drain_right.t4 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 drain_right.t3 minus.t8 source.t6 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 source.t22 plus.t4 drain_left.t7 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 source.t12 plus.t5 drain_left.t6 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X18 drain_right.t2 minus.t9 source.t10 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 drain_left.t5 plus.t6 source.t21 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X20 source.t23 minus.t10 drain_right.t1 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X21 drain_left.t4 plus.t7 source.t17 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X22 source.t18 plus.t8 drain_left.t3 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_right.t0 minus.t11 source.t4 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X24 a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X25 drain_left.t2 plus.t9 source.t19 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X26 drain_left.t1 plus.t10 source.t20 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X27 source.t15 plus.t11 drain_left.t0 a_n1626_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 plus.n2 plus.t5 584.973
R1 plus.n13 plus.t9 584.973
R2 plus.n17 plus.t7 584.973
R3 plus.n28 plus.t3 584.973
R4 plus.n3 plus.t10 530.201
R5 plus.n4 plus.t8 530.201
R6 plus.n10 plus.t6 530.201
R7 plus.n12 plus.t11 530.201
R8 plus.n19 plus.t4 530.201
R9 plus.n18 plus.t2 530.201
R10 plus.n25 plus.t1 530.201
R11 plus.n27 plus.t0 530.201
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 62.0763
R27 plus.n11 plus.n10 62.0763
R28 plus.n26 plus.n25 62.0763
R29 plus.n20 plus.n18 62.0763
R30 plus.n3 plus.n2 40.1672
R31 plus.n13 plus.n12 40.1672
R32 plus.n28 plus.n27 40.1672
R33 plus.n19 plus.n17 40.1672
R34 plus.n5 plus.n3 32.8641
R35 plus.n12 plus.n11 32.8641
R36 plus.n27 plus.n26 32.8641
R37 plus.n20 plus.n19 32.8641
R38 plus plus.n29 25.4157
R39 plus.n4 plus.n1 10.955
R40 plus.n10 plus.n9 10.955
R41 plus.n25 plus.n24 10.955
R42 plus.n18 plus.n16 10.955
R43 plus plus.n14 8.39823
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n0 source.t19 99.1169
R53 source.n5 source.t12 99.1169
R54 source.n6 source.t0 99.1169
R55 source.n11 source.t23 99.1169
R56 source.n23 source.t4 99.1168
R57 source.n18 source.t8 99.1168
R58 source.n17 source.t17 99.1168
R59 source.n12 source.t14 99.1168
R60 source.n2 source.n1 84.1169
R61 source.n4 source.n3 84.1169
R62 source.n8 source.n7 84.1169
R63 source.n10 source.n9 84.1169
R64 source.n22 source.n21 84.1168
R65 source.n20 source.n19 84.1168
R66 source.n16 source.n15 84.1168
R67 source.n14 source.n13 84.1168
R68 source.n21 source.t3 15.0005
R69 source.n21 source.t5 15.0005
R70 source.n19 source.t6 15.0005
R71 source.n19 source.t9 15.0005
R72 source.n15 source.t13 15.0005
R73 source.n15 source.t22 15.0005
R74 source.n13 source.t11 15.0005
R75 source.n13 source.t16 15.0005
R76 source.n1 source.t21 15.0005
R77 source.n1 source.t15 15.0005
R78 source.n3 source.t20 15.0005
R79 source.n3 source.t18 15.0005
R80 source.n7 source.t10 15.0005
R81 source.n7 source.t7 15.0005
R82 source.n9 source.t1 15.0005
R83 source.n9 source.t2 15.0005
R84 source.n12 source.n11 14.2723
R85 source.n24 source.n0 8.72921
R86 source.n24 source.n23 5.5436
R87 source.n11 source.n10 0.560845
R88 source.n10 source.n8 0.560845
R89 source.n8 source.n6 0.560845
R90 source.n5 source.n4 0.560845
R91 source.n4 source.n2 0.560845
R92 source.n2 source.n0 0.560845
R93 source.n14 source.n12 0.560845
R94 source.n16 source.n14 0.560845
R95 source.n17 source.n16 0.560845
R96 source.n20 source.n18 0.560845
R97 source.n22 source.n20 0.560845
R98 source.n23 source.n22 0.560845
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 101.356
R103 drain_left.n3 drain_left.n2 101.3
R104 drain_left.n3 drain_left.n0 101.3
R105 drain_left.n8 drain_left.n7 100.796
R106 drain_left.n6 drain_left.n5 100.796
R107 drain_left.n3 drain_left.n1 100.796
R108 drain_left drain_left.n3 22.593
R109 drain_left.n1 drain_left.t10 15.0005
R110 drain_left.n1 drain_left.t9 15.0005
R111 drain_left.n2 drain_left.t7 15.0005
R112 drain_left.n2 drain_left.t4 15.0005
R113 drain_left.n0 drain_left.t8 15.0005
R114 drain_left.n0 drain_left.t11 15.0005
R115 drain_left.n7 drain_left.t0 15.0005
R116 drain_left.n7 drain_left.t2 15.0005
R117 drain_left.n5 drain_left.t3 15.0005
R118 drain_left.n5 drain_left.t5 15.0005
R119 drain_left.n4 drain_left.t6 15.0005
R120 drain_left.n4 drain_left.t1 15.0005
R121 drain_left drain_left.n8 6.21356
R122 drain_left.n8 drain_left.n6 0.560845
R123 minus.n13 minus.t10 584.973
R124 minus.n2 minus.t5 584.973
R125 minus.n28 minus.t11 584.973
R126 minus.n17 minus.t1 584.973
R127 minus.n12 minus.t6 530.201
R128 minus.n10 minus.t7 530.201
R129 minus.n3 minus.t9 530.201
R130 minus.n4 minus.t3 530.201
R131 minus.n27 minus.t0 530.201
R132 minus.n25 minus.t2 530.201
R133 minus.n19 minus.t4 530.201
R134 minus.n18 minus.t8 530.201
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 62.0763
R150 minus.n5 minus.n3 62.0763
R151 minus.n20 minus.n19 62.0763
R152 minus.n26 minus.n25 62.0763
R153 minus.n13 minus.n12 40.1672
R154 minus.n4 minus.n2 40.1672
R155 minus.n18 minus.n17 40.1672
R156 minus.n28 minus.n27 40.1672
R157 minus.n12 minus.n11 32.8641
R158 minus.n5 minus.n4 32.8641
R159 minus.n20 minus.n18 32.8641
R160 minus.n27 minus.n26 32.8641
R161 minus.n30 minus.n14 27.7467
R162 minus.n10 minus.n9 10.955
R163 minus.n3 minus.n1 10.955
R164 minus.n19 minus.n16 10.955
R165 minus.n25 minus.n24 10.955
R166 minus.n30 minus.n29 6.54217
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 101.356
R177 drain_right.n3 drain_right.n2 101.3
R178 drain_right.n3 drain_right.n0 101.3
R179 drain_right.n6 drain_right.n5 100.796
R180 drain_right.n8 drain_right.n7 100.796
R181 drain_right.n3 drain_right.n1 100.796
R182 drain_right drain_right.n3 22.0398
R183 drain_right.n1 drain_right.t7 15.0005
R184 drain_right.n1 drain_right.t9 15.0005
R185 drain_right.n2 drain_right.t11 15.0005
R186 drain_right.n2 drain_right.t0 15.0005
R187 drain_right.n0 drain_right.t10 15.0005
R188 drain_right.n0 drain_right.t3 15.0005
R189 drain_right.n4 drain_right.t8 15.0005
R190 drain_right.n4 drain_right.t6 15.0005
R191 drain_right.n5 drain_right.t4 15.0005
R192 drain_right.n5 drain_right.t2 15.0005
R193 drain_right.n7 drain_right.t1 15.0005
R194 drain_right.n7 drain_right.t5 15.0005
R195 drain_right drain_right.n8 6.21356
R196 drain_right.n8 drain_right.n6 0.560845
C0 minus plus 3.31982f
C1 source drain_right 5.96636f
C2 source minus 0.894177f
C3 source plus 0.90814f
C4 drain_right drain_left 0.801778f
C5 minus drain_left 0.176524f
C6 plus drain_left 0.99297f
C7 minus drain_right 0.83651f
C8 plus drain_right 0.31642f
C9 source drain_left 5.96647f
C10 drain_right a_n1626_n1288# 3.49086f
C11 drain_left a_n1626_n1288# 3.71007f
C12 source a_n1626_n1288# 3.073667f
C13 minus a_n1626_n1288# 5.18409f
C14 plus a_n1626_n1288# 5.970277f
C15 drain_right.t10 a_n1626_n1288# 0.05766f
C16 drain_right.t3 a_n1626_n1288# 0.05766f
C17 drain_right.n0 a_n1626_n1288# 0.279672f
C18 drain_right.t7 a_n1626_n1288# 0.05766f
C19 drain_right.t9 a_n1626_n1288# 0.05766f
C20 drain_right.n1 a_n1626_n1288# 0.278288f
C21 drain_right.t11 a_n1626_n1288# 0.05766f
C22 drain_right.t0 a_n1626_n1288# 0.05766f
C23 drain_right.n2 a_n1626_n1288# 0.279672f
C24 drain_right.n3 a_n1626_n1288# 1.37226f
C25 drain_right.t8 a_n1626_n1288# 0.05766f
C26 drain_right.t6 a_n1626_n1288# 0.05766f
C27 drain_right.n4 a_n1626_n1288# 0.279842f
C28 drain_right.t4 a_n1626_n1288# 0.05766f
C29 drain_right.t2 a_n1626_n1288# 0.05766f
C30 drain_right.n5 a_n1626_n1288# 0.278289f
C31 drain_right.n6 a_n1626_n1288# 0.550644f
C32 drain_right.t1 a_n1626_n1288# 0.05766f
C33 drain_right.t5 a_n1626_n1288# 0.05766f
C34 drain_right.n7 a_n1626_n1288# 0.278289f
C35 drain_right.n8 a_n1626_n1288# 0.472334f
C36 minus.n0 a_n1626_n1288# 0.03533f
C37 minus.t10 a_n1626_n1288# 0.033789f
C38 minus.t6 a_n1626_n1288# 0.031188f
C39 minus.t7 a_n1626_n1288# 0.031188f
C40 minus.n1 a_n1626_n1288# 0.013354f
C41 minus.t5 a_n1626_n1288# 0.033789f
C42 minus.n2 a_n1626_n1288# 0.040211f
C43 minus.t9 a_n1626_n1288# 0.031188f
C44 minus.n3 a_n1626_n1288# 0.027228f
C45 minus.t3 a_n1626_n1288# 0.031188f
C46 minus.n4 a_n1626_n1288# 0.027228f
C47 minus.n5 a_n1626_n1288# 0.014987f
C48 minus.n6 a_n1626_n1288# 0.079321f
C49 minus.n7 a_n1626_n1288# 0.03533f
C50 minus.n8 a_n1626_n1288# 0.03533f
C51 minus.n9 a_n1626_n1288# 0.013354f
C52 minus.n10 a_n1626_n1288# 0.027228f
C53 minus.n11 a_n1626_n1288# 0.014987f
C54 minus.n12 a_n1626_n1288# 0.027228f
C55 minus.n13 a_n1626_n1288# 0.040159f
C56 minus.n14 a_n1626_n1288# 0.803648f
C57 minus.n15 a_n1626_n1288# 0.03533f
C58 minus.t0 a_n1626_n1288# 0.031188f
C59 minus.t2 a_n1626_n1288# 0.031188f
C60 minus.n16 a_n1626_n1288# 0.013354f
C61 minus.t1 a_n1626_n1288# 0.033789f
C62 minus.n17 a_n1626_n1288# 0.040211f
C63 minus.t8 a_n1626_n1288# 0.031188f
C64 minus.n18 a_n1626_n1288# 0.027228f
C65 minus.t4 a_n1626_n1288# 0.031188f
C66 minus.n19 a_n1626_n1288# 0.027228f
C67 minus.n20 a_n1626_n1288# 0.014987f
C68 minus.n21 a_n1626_n1288# 0.079321f
C69 minus.n22 a_n1626_n1288# 0.03533f
C70 minus.n23 a_n1626_n1288# 0.03533f
C71 minus.n24 a_n1626_n1288# 0.013354f
C72 minus.n25 a_n1626_n1288# 0.027228f
C73 minus.n26 a_n1626_n1288# 0.014987f
C74 minus.n27 a_n1626_n1288# 0.027228f
C75 minus.t11 a_n1626_n1288# 0.033789f
C76 minus.n28 a_n1626_n1288# 0.040159f
C77 minus.n29 a_n1626_n1288# 0.234479f
C78 minus.n30 a_n1626_n1288# 0.991465f
C79 drain_left.t8 a_n1626_n1288# 0.056769f
C80 drain_left.t11 a_n1626_n1288# 0.056769f
C81 drain_left.n0 a_n1626_n1288# 0.27535f
C82 drain_left.t10 a_n1626_n1288# 0.056769f
C83 drain_left.t9 a_n1626_n1288# 0.056769f
C84 drain_left.n1 a_n1626_n1288# 0.273986f
C85 drain_left.t7 a_n1626_n1288# 0.056769f
C86 drain_left.t4 a_n1626_n1288# 0.056769f
C87 drain_left.n2 a_n1626_n1288# 0.27535f
C88 drain_left.n3 a_n1626_n1288# 1.3976f
C89 drain_left.t6 a_n1626_n1288# 0.056769f
C90 drain_left.t1 a_n1626_n1288# 0.056769f
C91 drain_left.n4 a_n1626_n1288# 0.275517f
C92 drain_left.t3 a_n1626_n1288# 0.056769f
C93 drain_left.t5 a_n1626_n1288# 0.056769f
C94 drain_left.n5 a_n1626_n1288# 0.273987f
C95 drain_left.n6 a_n1626_n1288# 0.542133f
C96 drain_left.t0 a_n1626_n1288# 0.056769f
C97 drain_left.t2 a_n1626_n1288# 0.056769f
C98 drain_left.n7 a_n1626_n1288# 0.273987f
C99 drain_left.n8 a_n1626_n1288# 0.465033f
C100 source.t19 a_n1626_n1288# 0.303064f
C101 source.n0 a_n1626_n1288# 0.577632f
C102 source.t21 a_n1626_n1288# 0.057722f
C103 source.t15 a_n1626_n1288# 0.057722f
C104 source.n1 a_n1626_n1288# 0.242914f
C105 source.n2 a_n1626_n1288# 0.274448f
C106 source.t20 a_n1626_n1288# 0.057722f
C107 source.t18 a_n1626_n1288# 0.057722f
C108 source.n3 a_n1626_n1288# 0.242914f
C109 source.n4 a_n1626_n1288# 0.274448f
C110 source.t12 a_n1626_n1288# 0.303064f
C111 source.n5 a_n1626_n1288# 0.311168f
C112 source.t0 a_n1626_n1288# 0.303064f
C113 source.n6 a_n1626_n1288# 0.311168f
C114 source.t10 a_n1626_n1288# 0.057722f
C115 source.t7 a_n1626_n1288# 0.057722f
C116 source.n7 a_n1626_n1288# 0.242914f
C117 source.n8 a_n1626_n1288# 0.274448f
C118 source.t1 a_n1626_n1288# 0.057722f
C119 source.t2 a_n1626_n1288# 0.057722f
C120 source.n9 a_n1626_n1288# 0.242914f
C121 source.n10 a_n1626_n1288# 0.274448f
C122 source.t23 a_n1626_n1288# 0.303064f
C123 source.n11 a_n1626_n1288# 0.80266f
C124 source.t14 a_n1626_n1288# 0.303063f
C125 source.n12 a_n1626_n1288# 0.802661f
C126 source.t11 a_n1626_n1288# 0.057722f
C127 source.t16 a_n1626_n1288# 0.057722f
C128 source.n13 a_n1626_n1288# 0.242913f
C129 source.n14 a_n1626_n1288# 0.27445f
C130 source.t13 a_n1626_n1288# 0.057722f
C131 source.t22 a_n1626_n1288# 0.057722f
C132 source.n15 a_n1626_n1288# 0.242913f
C133 source.n16 a_n1626_n1288# 0.27445f
C134 source.t17 a_n1626_n1288# 0.303063f
C135 source.n17 a_n1626_n1288# 0.311169f
C136 source.t8 a_n1626_n1288# 0.303063f
C137 source.n18 a_n1626_n1288# 0.311169f
C138 source.t6 a_n1626_n1288# 0.057722f
C139 source.t9 a_n1626_n1288# 0.057722f
C140 source.n19 a_n1626_n1288# 0.242913f
C141 source.n20 a_n1626_n1288# 0.27445f
C142 source.t3 a_n1626_n1288# 0.057722f
C143 source.t5 a_n1626_n1288# 0.057722f
C144 source.n21 a_n1626_n1288# 0.242913f
C145 source.n22 a_n1626_n1288# 0.27445f
C146 source.t4 a_n1626_n1288# 0.303063f
C147 source.n23 a_n1626_n1288# 0.44831f
C148 source.n24 a_n1626_n1288# 0.596525f
C149 plus.n0 a_n1626_n1288# 0.036112f
C150 plus.t11 a_n1626_n1288# 0.031878f
C151 plus.t6 a_n1626_n1288# 0.031878f
C152 plus.n1 a_n1626_n1288# 0.013649f
C153 plus.t5 a_n1626_n1288# 0.034536f
C154 plus.n2 a_n1626_n1288# 0.041101f
C155 plus.t10 a_n1626_n1288# 0.031878f
C156 plus.n3 a_n1626_n1288# 0.02783f
C157 plus.t8 a_n1626_n1288# 0.031878f
C158 plus.n4 a_n1626_n1288# 0.02783f
C159 plus.n5 a_n1626_n1288# 0.015319f
C160 plus.n6 a_n1626_n1288# 0.081076f
C161 plus.n7 a_n1626_n1288# 0.036112f
C162 plus.n8 a_n1626_n1288# 0.036112f
C163 plus.n9 a_n1626_n1288# 0.013649f
C164 plus.n10 a_n1626_n1288# 0.02783f
C165 plus.n11 a_n1626_n1288# 0.015319f
C166 plus.n12 a_n1626_n1288# 0.02783f
C167 plus.t9 a_n1626_n1288# 0.034536f
C168 plus.n13 a_n1626_n1288# 0.041048f
C169 plus.n14 a_n1626_n1288# 0.261931f
C170 plus.n15 a_n1626_n1288# 0.036112f
C171 plus.t3 a_n1626_n1288# 0.034536f
C172 plus.t0 a_n1626_n1288# 0.031878f
C173 plus.t1 a_n1626_n1288# 0.031878f
C174 plus.n16 a_n1626_n1288# 0.013649f
C175 plus.t7 a_n1626_n1288# 0.034536f
C176 plus.n17 a_n1626_n1288# 0.041101f
C177 plus.t2 a_n1626_n1288# 0.031878f
C178 plus.n18 a_n1626_n1288# 0.02783f
C179 plus.t4 a_n1626_n1288# 0.031878f
C180 plus.n19 a_n1626_n1288# 0.02783f
C181 plus.n20 a_n1626_n1288# 0.015319f
C182 plus.n21 a_n1626_n1288# 0.081076f
C183 plus.n22 a_n1626_n1288# 0.036112f
C184 plus.n23 a_n1626_n1288# 0.036112f
C185 plus.n24 a_n1626_n1288# 0.013649f
C186 plus.n25 a_n1626_n1288# 0.02783f
C187 plus.n26 a_n1626_n1288# 0.015319f
C188 plus.n27 a_n1626_n1288# 0.02783f
C189 plus.n28 a_n1626_n1288# 0.041048f
C190 plus.n29 a_n1626_n1288# 0.786055f
.ends

