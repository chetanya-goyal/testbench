* NGSPICE file created from diffpair426.ext - technology: sky130A

.subckt diffpair426 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t4 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 source.t26 plus.t1 drain_left.t2 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X3 source.t9 minus.t0 drain_right.t13 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X4 source.t0 minus.t1 drain_right.t12 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X5 source.t11 minus.t2 drain_right.t11 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 drain_left.t12 plus.t2 source.t25 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X7 drain_left.t8 plus.t3 source.t24 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X8 drain_right.t10 minus.t3 source.t2 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X9 source.t7 minus.t4 drain_right.t9 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 drain_left.t7 plus.t4 source.t23 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X11 drain_left.t6 plus.t5 source.t22 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X12 drain_left.t13 plus.t6 source.t21 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X13 drain_left.t1 plus.t7 source.t20 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X14 drain_right.t8 minus.t5 source.t3 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X15 a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X16 drain_right.t7 minus.t6 source.t5 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X17 source.t12 minus.t7 drain_right.t6 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X18 a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X19 drain_left.t3 plus.t8 source.t19 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X20 source.t18 plus.t9 drain_left.t9 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X21 drain_right.t5 minus.t8 source.t6 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X22 drain_right.t4 minus.t9 source.t8 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X23 source.t17 plus.t10 drain_left.t11 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X24 drain_right.t3 minus.t10 source.t10 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X25 drain_right.t2 minus.t11 source.t4 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X26 drain_left.t5 plus.t11 source.t16 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X27 source.t1 minus.t12 drain_right.t1 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X28 source.t15 plus.t12 drain_left.t10 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X29 a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X30 drain_right.t0 minus.t13 source.t13 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X31 source.t14 plus.t13 drain_left.t0 a_n1644_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n3 plus.t3 1317.17
R1 plus.n15 plus.t5 1317.17
R2 plus.n20 plus.t11 1317.17
R3 plus.n32 plus.t8 1317.17
R4 plus.n1 plus.t0 1282.12
R5 plus.n4 plus.t1 1282.12
R6 plus.n6 plus.t7 1282.12
R7 plus.n12 plus.t6 1282.12
R8 plus.n14 plus.t12 1282.12
R9 plus.n18 plus.t13 1282.12
R10 plus.n21 plus.t9 1282.12
R11 plus.n23 plus.t4 1282.12
R12 plus.n29 plus.t2 1282.12
R13 plus.n31 plus.t10 1282.12
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 29.1808
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus plus.n16 12.0952
R46 plus.n7 plus.n6 11.6853
R47 plus.n12 plus.n11 11.6853
R48 plus.n29 plus.n28 11.6853
R49 plus.n24 plus.n23 11.6853
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n60 drain_left.n0 289.615
R61 drain_left.n131 drain_left.n71 289.615
R62 drain_left.n20 drain_left.n19 185
R63 drain_left.n25 drain_left.n24 185
R64 drain_left.n27 drain_left.n26 185
R65 drain_left.n16 drain_left.n15 185
R66 drain_left.n33 drain_left.n32 185
R67 drain_left.n35 drain_left.n34 185
R68 drain_left.n12 drain_left.n11 185
R69 drain_left.n42 drain_left.n41 185
R70 drain_left.n43 drain_left.n10 185
R71 drain_left.n45 drain_left.n44 185
R72 drain_left.n8 drain_left.n7 185
R73 drain_left.n51 drain_left.n50 185
R74 drain_left.n53 drain_left.n52 185
R75 drain_left.n4 drain_left.n3 185
R76 drain_left.n59 drain_left.n58 185
R77 drain_left.n61 drain_left.n60 185
R78 drain_left.n132 drain_left.n131 185
R79 drain_left.n130 drain_left.n129 185
R80 drain_left.n75 drain_left.n74 185
R81 drain_left.n124 drain_left.n123 185
R82 drain_left.n122 drain_left.n121 185
R83 drain_left.n79 drain_left.n78 185
R84 drain_left.n116 drain_left.n115 185
R85 drain_left.n114 drain_left.n81 185
R86 drain_left.n113 drain_left.n112 185
R87 drain_left.n84 drain_left.n82 185
R88 drain_left.n107 drain_left.n106 185
R89 drain_left.n105 drain_left.n104 185
R90 drain_left.n88 drain_left.n87 185
R91 drain_left.n99 drain_left.n98 185
R92 drain_left.n97 drain_left.n96 185
R93 drain_left.n92 drain_left.n91 185
R94 drain_left.n21 drain_left.t3 149.524
R95 drain_left.n93 drain_left.t8 149.524
R96 drain_left.n25 drain_left.n19 104.615
R97 drain_left.n26 drain_left.n25 104.615
R98 drain_left.n26 drain_left.n15 104.615
R99 drain_left.n33 drain_left.n15 104.615
R100 drain_left.n34 drain_left.n33 104.615
R101 drain_left.n34 drain_left.n11 104.615
R102 drain_left.n42 drain_left.n11 104.615
R103 drain_left.n43 drain_left.n42 104.615
R104 drain_left.n44 drain_left.n43 104.615
R105 drain_left.n44 drain_left.n7 104.615
R106 drain_left.n51 drain_left.n7 104.615
R107 drain_left.n52 drain_left.n51 104.615
R108 drain_left.n52 drain_left.n3 104.615
R109 drain_left.n59 drain_left.n3 104.615
R110 drain_left.n60 drain_left.n59 104.615
R111 drain_left.n131 drain_left.n130 104.615
R112 drain_left.n130 drain_left.n74 104.615
R113 drain_left.n123 drain_left.n74 104.615
R114 drain_left.n123 drain_left.n122 104.615
R115 drain_left.n122 drain_left.n78 104.615
R116 drain_left.n115 drain_left.n78 104.615
R117 drain_left.n115 drain_left.n114 104.615
R118 drain_left.n114 drain_left.n113 104.615
R119 drain_left.n113 drain_left.n82 104.615
R120 drain_left.n106 drain_left.n82 104.615
R121 drain_left.n106 drain_left.n105 104.615
R122 drain_left.n105 drain_left.n87 104.615
R123 drain_left.n98 drain_left.n87 104.615
R124 drain_left.n98 drain_left.n97 104.615
R125 drain_left.n97 drain_left.n91 104.615
R126 drain_left.n69 drain_left.n67 60.0525
R127 drain_left.n139 drain_left.n138 59.5527
R128 drain_left.n137 drain_left.n136 59.5527
R129 drain_left.n69 drain_left.n68 59.5525
R130 drain_left.n66 drain_left.n65 59.5525
R131 drain_left.n141 drain_left.n140 59.5525
R132 drain_left.t3 drain_left.n19 52.3082
R133 drain_left.t8 drain_left.n91 52.3082
R134 drain_left.n66 drain_left.n64 47.0369
R135 drain_left.n137 drain_left.n135 47.0369
R136 drain_left drain_left.n70 30.2421
R137 drain_left.n45 drain_left.n10 13.1884
R138 drain_left.n116 drain_left.n81 13.1884
R139 drain_left.n41 drain_left.n40 12.8005
R140 drain_left.n46 drain_left.n8 12.8005
R141 drain_left.n117 drain_left.n79 12.8005
R142 drain_left.n112 drain_left.n83 12.8005
R143 drain_left.n39 drain_left.n12 12.0247
R144 drain_left.n50 drain_left.n49 12.0247
R145 drain_left.n121 drain_left.n120 12.0247
R146 drain_left.n111 drain_left.n84 12.0247
R147 drain_left.n36 drain_left.n35 11.249
R148 drain_left.n53 drain_left.n6 11.249
R149 drain_left.n124 drain_left.n77 11.249
R150 drain_left.n108 drain_left.n107 11.249
R151 drain_left.n32 drain_left.n14 10.4732
R152 drain_left.n54 drain_left.n4 10.4732
R153 drain_left.n125 drain_left.n75 10.4732
R154 drain_left.n104 drain_left.n86 10.4732
R155 drain_left.n21 drain_left.n20 10.2747
R156 drain_left.n93 drain_left.n92 10.2747
R157 drain_left.n31 drain_left.n16 9.69747
R158 drain_left.n58 drain_left.n57 9.69747
R159 drain_left.n129 drain_left.n128 9.69747
R160 drain_left.n103 drain_left.n88 9.69747
R161 drain_left.n64 drain_left.n63 9.45567
R162 drain_left.n135 drain_left.n134 9.45567
R163 drain_left.n63 drain_left.n62 9.3005
R164 drain_left.n2 drain_left.n1 9.3005
R165 drain_left.n57 drain_left.n56 9.3005
R166 drain_left.n55 drain_left.n54 9.3005
R167 drain_left.n6 drain_left.n5 9.3005
R168 drain_left.n49 drain_left.n48 9.3005
R169 drain_left.n47 drain_left.n46 9.3005
R170 drain_left.n23 drain_left.n22 9.3005
R171 drain_left.n18 drain_left.n17 9.3005
R172 drain_left.n29 drain_left.n28 9.3005
R173 drain_left.n31 drain_left.n30 9.3005
R174 drain_left.n14 drain_left.n13 9.3005
R175 drain_left.n37 drain_left.n36 9.3005
R176 drain_left.n39 drain_left.n38 9.3005
R177 drain_left.n40 drain_left.n9 9.3005
R178 drain_left.n95 drain_left.n94 9.3005
R179 drain_left.n90 drain_left.n89 9.3005
R180 drain_left.n101 drain_left.n100 9.3005
R181 drain_left.n103 drain_left.n102 9.3005
R182 drain_left.n86 drain_left.n85 9.3005
R183 drain_left.n109 drain_left.n108 9.3005
R184 drain_left.n111 drain_left.n110 9.3005
R185 drain_left.n83 drain_left.n80 9.3005
R186 drain_left.n134 drain_left.n133 9.3005
R187 drain_left.n73 drain_left.n72 9.3005
R188 drain_left.n128 drain_left.n127 9.3005
R189 drain_left.n126 drain_left.n125 9.3005
R190 drain_left.n77 drain_left.n76 9.3005
R191 drain_left.n120 drain_left.n119 9.3005
R192 drain_left.n118 drain_left.n117 9.3005
R193 drain_left.n28 drain_left.n27 8.92171
R194 drain_left.n61 drain_left.n2 8.92171
R195 drain_left.n132 drain_left.n73 8.92171
R196 drain_left.n100 drain_left.n99 8.92171
R197 drain_left.n24 drain_left.n18 8.14595
R198 drain_left.n62 drain_left.n0 8.14595
R199 drain_left.n133 drain_left.n71 8.14595
R200 drain_left.n96 drain_left.n90 8.14595
R201 drain_left.n23 drain_left.n20 7.3702
R202 drain_left.n95 drain_left.n92 7.3702
R203 drain_left drain_left.n141 6.15322
R204 drain_left.n24 drain_left.n23 5.81868
R205 drain_left.n64 drain_left.n0 5.81868
R206 drain_left.n135 drain_left.n71 5.81868
R207 drain_left.n96 drain_left.n95 5.81868
R208 drain_left.n27 drain_left.n18 5.04292
R209 drain_left.n62 drain_left.n61 5.04292
R210 drain_left.n133 drain_left.n132 5.04292
R211 drain_left.n99 drain_left.n90 5.04292
R212 drain_left.n28 drain_left.n16 4.26717
R213 drain_left.n58 drain_left.n2 4.26717
R214 drain_left.n129 drain_left.n73 4.26717
R215 drain_left.n100 drain_left.n88 4.26717
R216 drain_left.n32 drain_left.n31 3.49141
R217 drain_left.n57 drain_left.n4 3.49141
R218 drain_left.n128 drain_left.n75 3.49141
R219 drain_left.n104 drain_left.n103 3.49141
R220 drain_left.n22 drain_left.n21 2.84303
R221 drain_left.n94 drain_left.n93 2.84303
R222 drain_left.n35 drain_left.n14 2.71565
R223 drain_left.n54 drain_left.n53 2.71565
R224 drain_left.n125 drain_left.n124 2.71565
R225 drain_left.n107 drain_left.n86 2.71565
R226 drain_left.n36 drain_left.n12 1.93989
R227 drain_left.n50 drain_left.n6 1.93989
R228 drain_left.n121 drain_left.n77 1.93989
R229 drain_left.n108 drain_left.n84 1.93989
R230 drain_left.n67 drain_left.t9 1.6505
R231 drain_left.n67 drain_left.t5 1.6505
R232 drain_left.n68 drain_left.t0 1.6505
R233 drain_left.n68 drain_left.t7 1.6505
R234 drain_left.n65 drain_left.t11 1.6505
R235 drain_left.n65 drain_left.t12 1.6505
R236 drain_left.n140 drain_left.t10 1.6505
R237 drain_left.n140 drain_left.t6 1.6505
R238 drain_left.n138 drain_left.t4 1.6505
R239 drain_left.n138 drain_left.t13 1.6505
R240 drain_left.n136 drain_left.t2 1.6505
R241 drain_left.n136 drain_left.t1 1.6505
R242 drain_left.n41 drain_left.n39 1.16414
R243 drain_left.n49 drain_left.n8 1.16414
R244 drain_left.n120 drain_left.n79 1.16414
R245 drain_left.n112 drain_left.n111 1.16414
R246 drain_left.n139 drain_left.n137 0.5005
R247 drain_left.n141 drain_left.n139 0.5005
R248 drain_left.n40 drain_left.n10 0.388379
R249 drain_left.n46 drain_left.n45 0.388379
R250 drain_left.n117 drain_left.n116 0.388379
R251 drain_left.n83 drain_left.n81 0.388379
R252 drain_left.n70 drain_left.n66 0.320154
R253 drain_left.n22 drain_left.n17 0.155672
R254 drain_left.n29 drain_left.n17 0.155672
R255 drain_left.n30 drain_left.n29 0.155672
R256 drain_left.n30 drain_left.n13 0.155672
R257 drain_left.n37 drain_left.n13 0.155672
R258 drain_left.n38 drain_left.n37 0.155672
R259 drain_left.n38 drain_left.n9 0.155672
R260 drain_left.n47 drain_left.n9 0.155672
R261 drain_left.n48 drain_left.n47 0.155672
R262 drain_left.n48 drain_left.n5 0.155672
R263 drain_left.n55 drain_left.n5 0.155672
R264 drain_left.n56 drain_left.n55 0.155672
R265 drain_left.n56 drain_left.n1 0.155672
R266 drain_left.n63 drain_left.n1 0.155672
R267 drain_left.n134 drain_left.n72 0.155672
R268 drain_left.n127 drain_left.n72 0.155672
R269 drain_left.n127 drain_left.n126 0.155672
R270 drain_left.n126 drain_left.n76 0.155672
R271 drain_left.n119 drain_left.n76 0.155672
R272 drain_left.n119 drain_left.n118 0.155672
R273 drain_left.n118 drain_left.n80 0.155672
R274 drain_left.n110 drain_left.n80 0.155672
R275 drain_left.n110 drain_left.n109 0.155672
R276 drain_left.n109 drain_left.n85 0.155672
R277 drain_left.n102 drain_left.n85 0.155672
R278 drain_left.n102 drain_left.n101 0.155672
R279 drain_left.n101 drain_left.n89 0.155672
R280 drain_left.n94 drain_left.n89 0.155672
R281 drain_left.n70 drain_left.n69 0.070154
R282 source.n282 source.n222 289.615
R283 source.n210 source.n150 289.615
R284 source.n60 source.n0 289.615
R285 source.n132 source.n72 289.615
R286 source.n242 source.n241 185
R287 source.n247 source.n246 185
R288 source.n249 source.n248 185
R289 source.n238 source.n237 185
R290 source.n255 source.n254 185
R291 source.n257 source.n256 185
R292 source.n234 source.n233 185
R293 source.n264 source.n263 185
R294 source.n265 source.n232 185
R295 source.n267 source.n266 185
R296 source.n230 source.n229 185
R297 source.n273 source.n272 185
R298 source.n275 source.n274 185
R299 source.n226 source.n225 185
R300 source.n281 source.n280 185
R301 source.n283 source.n282 185
R302 source.n170 source.n169 185
R303 source.n175 source.n174 185
R304 source.n177 source.n176 185
R305 source.n166 source.n165 185
R306 source.n183 source.n182 185
R307 source.n185 source.n184 185
R308 source.n162 source.n161 185
R309 source.n192 source.n191 185
R310 source.n193 source.n160 185
R311 source.n195 source.n194 185
R312 source.n158 source.n157 185
R313 source.n201 source.n200 185
R314 source.n203 source.n202 185
R315 source.n154 source.n153 185
R316 source.n209 source.n208 185
R317 source.n211 source.n210 185
R318 source.n61 source.n60 185
R319 source.n59 source.n58 185
R320 source.n4 source.n3 185
R321 source.n53 source.n52 185
R322 source.n51 source.n50 185
R323 source.n8 source.n7 185
R324 source.n45 source.n44 185
R325 source.n43 source.n10 185
R326 source.n42 source.n41 185
R327 source.n13 source.n11 185
R328 source.n36 source.n35 185
R329 source.n34 source.n33 185
R330 source.n17 source.n16 185
R331 source.n28 source.n27 185
R332 source.n26 source.n25 185
R333 source.n21 source.n20 185
R334 source.n133 source.n132 185
R335 source.n131 source.n130 185
R336 source.n76 source.n75 185
R337 source.n125 source.n124 185
R338 source.n123 source.n122 185
R339 source.n80 source.n79 185
R340 source.n117 source.n116 185
R341 source.n115 source.n82 185
R342 source.n114 source.n113 185
R343 source.n85 source.n83 185
R344 source.n108 source.n107 185
R345 source.n106 source.n105 185
R346 source.n89 source.n88 185
R347 source.n100 source.n99 185
R348 source.n98 source.n97 185
R349 source.n93 source.n92 185
R350 source.n243 source.t6 149.524
R351 source.n171 source.t16 149.524
R352 source.n22 source.t22 149.524
R353 source.n94 source.t5 149.524
R354 source.n247 source.n241 104.615
R355 source.n248 source.n247 104.615
R356 source.n248 source.n237 104.615
R357 source.n255 source.n237 104.615
R358 source.n256 source.n255 104.615
R359 source.n256 source.n233 104.615
R360 source.n264 source.n233 104.615
R361 source.n265 source.n264 104.615
R362 source.n266 source.n265 104.615
R363 source.n266 source.n229 104.615
R364 source.n273 source.n229 104.615
R365 source.n274 source.n273 104.615
R366 source.n274 source.n225 104.615
R367 source.n281 source.n225 104.615
R368 source.n282 source.n281 104.615
R369 source.n175 source.n169 104.615
R370 source.n176 source.n175 104.615
R371 source.n176 source.n165 104.615
R372 source.n183 source.n165 104.615
R373 source.n184 source.n183 104.615
R374 source.n184 source.n161 104.615
R375 source.n192 source.n161 104.615
R376 source.n193 source.n192 104.615
R377 source.n194 source.n193 104.615
R378 source.n194 source.n157 104.615
R379 source.n201 source.n157 104.615
R380 source.n202 source.n201 104.615
R381 source.n202 source.n153 104.615
R382 source.n209 source.n153 104.615
R383 source.n210 source.n209 104.615
R384 source.n60 source.n59 104.615
R385 source.n59 source.n3 104.615
R386 source.n52 source.n3 104.615
R387 source.n52 source.n51 104.615
R388 source.n51 source.n7 104.615
R389 source.n44 source.n7 104.615
R390 source.n44 source.n43 104.615
R391 source.n43 source.n42 104.615
R392 source.n42 source.n11 104.615
R393 source.n35 source.n11 104.615
R394 source.n35 source.n34 104.615
R395 source.n34 source.n16 104.615
R396 source.n27 source.n16 104.615
R397 source.n27 source.n26 104.615
R398 source.n26 source.n20 104.615
R399 source.n132 source.n131 104.615
R400 source.n131 source.n75 104.615
R401 source.n124 source.n75 104.615
R402 source.n124 source.n123 104.615
R403 source.n123 source.n79 104.615
R404 source.n116 source.n79 104.615
R405 source.n116 source.n115 104.615
R406 source.n115 source.n114 104.615
R407 source.n114 source.n83 104.615
R408 source.n107 source.n83 104.615
R409 source.n107 source.n106 104.615
R410 source.n106 source.n88 104.615
R411 source.n99 source.n88 104.615
R412 source.n99 source.n98 104.615
R413 source.n98 source.n92 104.615
R414 source.t6 source.n241 52.3082
R415 source.t16 source.n169 52.3082
R416 source.t22 source.n20 52.3082
R417 source.t5 source.n92 52.3082
R418 source.n67 source.n66 42.8739
R419 source.n69 source.n68 42.8739
R420 source.n71 source.n70 42.8739
R421 source.n139 source.n138 42.8739
R422 source.n141 source.n140 42.8739
R423 source.n143 source.n142 42.8739
R424 source.n221 source.n220 42.8737
R425 source.n219 source.n218 42.8737
R426 source.n217 source.n216 42.8737
R427 source.n149 source.n148 42.8737
R428 source.n147 source.n146 42.8737
R429 source.n145 source.n144 42.8737
R430 source.n287 source.n286 29.8581
R431 source.n215 source.n214 29.8581
R432 source.n65 source.n64 29.8581
R433 source.n137 source.n136 29.8581
R434 source.n145 source.n143 22.2877
R435 source.n288 source.n65 16.2748
R436 source.n267 source.n232 13.1884
R437 source.n195 source.n160 13.1884
R438 source.n45 source.n10 13.1884
R439 source.n117 source.n82 13.1884
R440 source.n263 source.n262 12.8005
R441 source.n268 source.n230 12.8005
R442 source.n191 source.n190 12.8005
R443 source.n196 source.n158 12.8005
R444 source.n46 source.n8 12.8005
R445 source.n41 source.n12 12.8005
R446 source.n118 source.n80 12.8005
R447 source.n113 source.n84 12.8005
R448 source.n261 source.n234 12.0247
R449 source.n272 source.n271 12.0247
R450 source.n189 source.n162 12.0247
R451 source.n200 source.n199 12.0247
R452 source.n50 source.n49 12.0247
R453 source.n40 source.n13 12.0247
R454 source.n122 source.n121 12.0247
R455 source.n112 source.n85 12.0247
R456 source.n258 source.n257 11.249
R457 source.n275 source.n228 11.249
R458 source.n186 source.n185 11.249
R459 source.n203 source.n156 11.249
R460 source.n53 source.n6 11.249
R461 source.n37 source.n36 11.249
R462 source.n125 source.n78 11.249
R463 source.n109 source.n108 11.249
R464 source.n254 source.n236 10.4732
R465 source.n276 source.n226 10.4732
R466 source.n182 source.n164 10.4732
R467 source.n204 source.n154 10.4732
R468 source.n54 source.n4 10.4732
R469 source.n33 source.n15 10.4732
R470 source.n126 source.n76 10.4732
R471 source.n105 source.n87 10.4732
R472 source.n243 source.n242 10.2747
R473 source.n171 source.n170 10.2747
R474 source.n22 source.n21 10.2747
R475 source.n94 source.n93 10.2747
R476 source.n253 source.n238 9.69747
R477 source.n280 source.n279 9.69747
R478 source.n181 source.n166 9.69747
R479 source.n208 source.n207 9.69747
R480 source.n58 source.n57 9.69747
R481 source.n32 source.n17 9.69747
R482 source.n130 source.n129 9.69747
R483 source.n104 source.n89 9.69747
R484 source.n286 source.n285 9.45567
R485 source.n214 source.n213 9.45567
R486 source.n64 source.n63 9.45567
R487 source.n136 source.n135 9.45567
R488 source.n285 source.n284 9.3005
R489 source.n224 source.n223 9.3005
R490 source.n279 source.n278 9.3005
R491 source.n277 source.n276 9.3005
R492 source.n228 source.n227 9.3005
R493 source.n271 source.n270 9.3005
R494 source.n269 source.n268 9.3005
R495 source.n245 source.n244 9.3005
R496 source.n240 source.n239 9.3005
R497 source.n251 source.n250 9.3005
R498 source.n253 source.n252 9.3005
R499 source.n236 source.n235 9.3005
R500 source.n259 source.n258 9.3005
R501 source.n261 source.n260 9.3005
R502 source.n262 source.n231 9.3005
R503 source.n213 source.n212 9.3005
R504 source.n152 source.n151 9.3005
R505 source.n207 source.n206 9.3005
R506 source.n205 source.n204 9.3005
R507 source.n156 source.n155 9.3005
R508 source.n199 source.n198 9.3005
R509 source.n197 source.n196 9.3005
R510 source.n173 source.n172 9.3005
R511 source.n168 source.n167 9.3005
R512 source.n179 source.n178 9.3005
R513 source.n181 source.n180 9.3005
R514 source.n164 source.n163 9.3005
R515 source.n187 source.n186 9.3005
R516 source.n189 source.n188 9.3005
R517 source.n190 source.n159 9.3005
R518 source.n24 source.n23 9.3005
R519 source.n19 source.n18 9.3005
R520 source.n30 source.n29 9.3005
R521 source.n32 source.n31 9.3005
R522 source.n15 source.n14 9.3005
R523 source.n38 source.n37 9.3005
R524 source.n40 source.n39 9.3005
R525 source.n12 source.n9 9.3005
R526 source.n63 source.n62 9.3005
R527 source.n2 source.n1 9.3005
R528 source.n57 source.n56 9.3005
R529 source.n55 source.n54 9.3005
R530 source.n6 source.n5 9.3005
R531 source.n49 source.n48 9.3005
R532 source.n47 source.n46 9.3005
R533 source.n96 source.n95 9.3005
R534 source.n91 source.n90 9.3005
R535 source.n102 source.n101 9.3005
R536 source.n104 source.n103 9.3005
R537 source.n87 source.n86 9.3005
R538 source.n110 source.n109 9.3005
R539 source.n112 source.n111 9.3005
R540 source.n84 source.n81 9.3005
R541 source.n135 source.n134 9.3005
R542 source.n74 source.n73 9.3005
R543 source.n129 source.n128 9.3005
R544 source.n127 source.n126 9.3005
R545 source.n78 source.n77 9.3005
R546 source.n121 source.n120 9.3005
R547 source.n119 source.n118 9.3005
R548 source.n250 source.n249 8.92171
R549 source.n283 source.n224 8.92171
R550 source.n178 source.n177 8.92171
R551 source.n211 source.n152 8.92171
R552 source.n61 source.n2 8.92171
R553 source.n29 source.n28 8.92171
R554 source.n133 source.n74 8.92171
R555 source.n101 source.n100 8.92171
R556 source.n246 source.n240 8.14595
R557 source.n284 source.n222 8.14595
R558 source.n174 source.n168 8.14595
R559 source.n212 source.n150 8.14595
R560 source.n62 source.n0 8.14595
R561 source.n25 source.n19 8.14595
R562 source.n134 source.n72 8.14595
R563 source.n97 source.n91 8.14595
R564 source.n245 source.n242 7.3702
R565 source.n173 source.n170 7.3702
R566 source.n24 source.n21 7.3702
R567 source.n96 source.n93 7.3702
R568 source.n246 source.n245 5.81868
R569 source.n286 source.n222 5.81868
R570 source.n174 source.n173 5.81868
R571 source.n214 source.n150 5.81868
R572 source.n64 source.n0 5.81868
R573 source.n25 source.n24 5.81868
R574 source.n136 source.n72 5.81868
R575 source.n97 source.n96 5.81868
R576 source.n288 source.n287 5.51343
R577 source.n249 source.n240 5.04292
R578 source.n284 source.n283 5.04292
R579 source.n177 source.n168 5.04292
R580 source.n212 source.n211 5.04292
R581 source.n62 source.n61 5.04292
R582 source.n28 source.n19 5.04292
R583 source.n134 source.n133 5.04292
R584 source.n100 source.n91 5.04292
R585 source.n250 source.n238 4.26717
R586 source.n280 source.n224 4.26717
R587 source.n178 source.n166 4.26717
R588 source.n208 source.n152 4.26717
R589 source.n58 source.n2 4.26717
R590 source.n29 source.n17 4.26717
R591 source.n130 source.n74 4.26717
R592 source.n101 source.n89 4.26717
R593 source.n254 source.n253 3.49141
R594 source.n279 source.n226 3.49141
R595 source.n182 source.n181 3.49141
R596 source.n207 source.n154 3.49141
R597 source.n57 source.n4 3.49141
R598 source.n33 source.n32 3.49141
R599 source.n129 source.n76 3.49141
R600 source.n105 source.n104 3.49141
R601 source.n244 source.n243 2.84303
R602 source.n172 source.n171 2.84303
R603 source.n23 source.n22 2.84303
R604 source.n95 source.n94 2.84303
R605 source.n257 source.n236 2.71565
R606 source.n276 source.n275 2.71565
R607 source.n185 source.n164 2.71565
R608 source.n204 source.n203 2.71565
R609 source.n54 source.n53 2.71565
R610 source.n36 source.n15 2.71565
R611 source.n126 source.n125 2.71565
R612 source.n108 source.n87 2.71565
R613 source.n258 source.n234 1.93989
R614 source.n272 source.n228 1.93989
R615 source.n186 source.n162 1.93989
R616 source.n200 source.n156 1.93989
R617 source.n50 source.n6 1.93989
R618 source.n37 source.n13 1.93989
R619 source.n122 source.n78 1.93989
R620 source.n109 source.n85 1.93989
R621 source.n220 source.t2 1.6505
R622 source.n220 source.t1 1.6505
R623 source.n218 source.t8 1.6505
R624 source.n218 source.t12 1.6505
R625 source.n216 source.t13 1.6505
R626 source.n216 source.t11 1.6505
R627 source.n148 source.t23 1.6505
R628 source.n148 source.t18 1.6505
R629 source.n146 source.t25 1.6505
R630 source.n146 source.t14 1.6505
R631 source.n144 source.t19 1.6505
R632 source.n144 source.t17 1.6505
R633 source.n66 source.t21 1.6505
R634 source.n66 source.t15 1.6505
R635 source.n68 source.t20 1.6505
R636 source.n68 source.t27 1.6505
R637 source.n70 source.t24 1.6505
R638 source.n70 source.t26 1.6505
R639 source.n138 source.t3 1.6505
R640 source.n138 source.t0 1.6505
R641 source.n140 source.t10 1.6505
R642 source.n140 source.t9 1.6505
R643 source.n142 source.t4 1.6505
R644 source.n142 source.t7 1.6505
R645 source.n263 source.n261 1.16414
R646 source.n271 source.n230 1.16414
R647 source.n191 source.n189 1.16414
R648 source.n199 source.n158 1.16414
R649 source.n49 source.n8 1.16414
R650 source.n41 source.n40 1.16414
R651 source.n121 source.n80 1.16414
R652 source.n113 source.n112 1.16414
R653 source.n137 source.n71 0.720328
R654 source.n217 source.n215 0.720328
R655 source.n143 source.n141 0.5005
R656 source.n141 source.n139 0.5005
R657 source.n139 source.n137 0.5005
R658 source.n71 source.n69 0.5005
R659 source.n69 source.n67 0.5005
R660 source.n67 source.n65 0.5005
R661 source.n147 source.n145 0.5005
R662 source.n149 source.n147 0.5005
R663 source.n215 source.n149 0.5005
R664 source.n219 source.n217 0.5005
R665 source.n221 source.n219 0.5005
R666 source.n287 source.n221 0.5005
R667 source.n262 source.n232 0.388379
R668 source.n268 source.n267 0.388379
R669 source.n190 source.n160 0.388379
R670 source.n196 source.n195 0.388379
R671 source.n46 source.n45 0.388379
R672 source.n12 source.n10 0.388379
R673 source.n118 source.n117 0.388379
R674 source.n84 source.n82 0.388379
R675 source source.n288 0.188
R676 source.n244 source.n239 0.155672
R677 source.n251 source.n239 0.155672
R678 source.n252 source.n251 0.155672
R679 source.n252 source.n235 0.155672
R680 source.n259 source.n235 0.155672
R681 source.n260 source.n259 0.155672
R682 source.n260 source.n231 0.155672
R683 source.n269 source.n231 0.155672
R684 source.n270 source.n269 0.155672
R685 source.n270 source.n227 0.155672
R686 source.n277 source.n227 0.155672
R687 source.n278 source.n277 0.155672
R688 source.n278 source.n223 0.155672
R689 source.n285 source.n223 0.155672
R690 source.n172 source.n167 0.155672
R691 source.n179 source.n167 0.155672
R692 source.n180 source.n179 0.155672
R693 source.n180 source.n163 0.155672
R694 source.n187 source.n163 0.155672
R695 source.n188 source.n187 0.155672
R696 source.n188 source.n159 0.155672
R697 source.n197 source.n159 0.155672
R698 source.n198 source.n197 0.155672
R699 source.n198 source.n155 0.155672
R700 source.n205 source.n155 0.155672
R701 source.n206 source.n205 0.155672
R702 source.n206 source.n151 0.155672
R703 source.n213 source.n151 0.155672
R704 source.n63 source.n1 0.155672
R705 source.n56 source.n1 0.155672
R706 source.n56 source.n55 0.155672
R707 source.n55 source.n5 0.155672
R708 source.n48 source.n5 0.155672
R709 source.n48 source.n47 0.155672
R710 source.n47 source.n9 0.155672
R711 source.n39 source.n9 0.155672
R712 source.n39 source.n38 0.155672
R713 source.n38 source.n14 0.155672
R714 source.n31 source.n14 0.155672
R715 source.n31 source.n30 0.155672
R716 source.n30 source.n18 0.155672
R717 source.n23 source.n18 0.155672
R718 source.n135 source.n73 0.155672
R719 source.n128 source.n73 0.155672
R720 source.n128 source.n127 0.155672
R721 source.n127 source.n77 0.155672
R722 source.n120 source.n77 0.155672
R723 source.n120 source.n119 0.155672
R724 source.n119 source.n81 0.155672
R725 source.n111 source.n81 0.155672
R726 source.n111 source.n110 0.155672
R727 source.n110 source.n86 0.155672
R728 source.n103 source.n86 0.155672
R729 source.n103 source.n102 0.155672
R730 source.n102 source.n90 0.155672
R731 source.n95 source.n90 0.155672
R732 minus.n15 minus.t11 1317.17
R733 minus.n3 minus.t6 1317.17
R734 minus.n32 minus.t8 1317.17
R735 minus.n20 minus.t13 1317.17
R736 minus.n1 minus.t0 1282.12
R737 minus.n14 minus.t4 1282.12
R738 minus.n12 minus.t10 1282.12
R739 minus.n6 minus.t5 1282.12
R740 minus.n4 minus.t1 1282.12
R741 minus.n18 minus.t7 1282.12
R742 minus.n31 minus.t12 1282.12
R743 minus.n29 minus.t3 1282.12
R744 minus.n23 minus.t9 1282.12
R745 minus.n21 minus.t2 1282.12
R746 minus.n3 minus.n2 161.489
R747 minus.n20 minus.n19 161.489
R748 minus.n16 minus.n15 161.3
R749 minus.n13 minus.n0 161.3
R750 minus.n11 minus.n10 161.3
R751 minus.n9 minus.n1 161.3
R752 minus.n8 minus.n7 161.3
R753 minus.n5 minus.n2 161.3
R754 minus.n33 minus.n32 161.3
R755 minus.n30 minus.n17 161.3
R756 minus.n28 minus.n27 161.3
R757 minus.n26 minus.n18 161.3
R758 minus.n25 minus.n24 161.3
R759 minus.n22 minus.n19 161.3
R760 minus.n11 minus.n1 73.0308
R761 minus.n7 minus.n1 73.0308
R762 minus.n24 minus.n18 73.0308
R763 minus.n28 minus.n18 73.0308
R764 minus.n13 minus.n12 61.346
R765 minus.n6 minus.n5 61.346
R766 minus.n23 minus.n22 61.346
R767 minus.n30 minus.n29 61.346
R768 minus.n15 minus.n14 49.6611
R769 minus.n4 minus.n3 49.6611
R770 minus.n21 minus.n20 49.6611
R771 minus.n32 minus.n31 49.6611
R772 minus.n34 minus.n16 35.2997
R773 minus.n14 minus.n13 23.3702
R774 minus.n5 minus.n4 23.3702
R775 minus.n22 minus.n21 23.3702
R776 minus.n31 minus.n30 23.3702
R777 minus.n12 minus.n11 11.6853
R778 minus.n7 minus.n6 11.6853
R779 minus.n24 minus.n23 11.6853
R780 minus.n29 minus.n28 11.6853
R781 minus.n34 minus.n33 6.45126
R782 minus.n16 minus.n0 0.189894
R783 minus.n10 minus.n0 0.189894
R784 minus.n10 minus.n9 0.189894
R785 minus.n9 minus.n8 0.189894
R786 minus.n8 minus.n2 0.189894
R787 minus.n25 minus.n19 0.189894
R788 minus.n26 minus.n25 0.189894
R789 minus.n27 minus.n26 0.189894
R790 minus.n27 minus.n17 0.189894
R791 minus.n33 minus.n17 0.189894
R792 minus minus.n34 0.188
R793 drain_right.n60 drain_right.n0 289.615
R794 drain_right.n136 drain_right.n76 289.615
R795 drain_right.n20 drain_right.n19 185
R796 drain_right.n25 drain_right.n24 185
R797 drain_right.n27 drain_right.n26 185
R798 drain_right.n16 drain_right.n15 185
R799 drain_right.n33 drain_right.n32 185
R800 drain_right.n35 drain_right.n34 185
R801 drain_right.n12 drain_right.n11 185
R802 drain_right.n42 drain_right.n41 185
R803 drain_right.n43 drain_right.n10 185
R804 drain_right.n45 drain_right.n44 185
R805 drain_right.n8 drain_right.n7 185
R806 drain_right.n51 drain_right.n50 185
R807 drain_right.n53 drain_right.n52 185
R808 drain_right.n4 drain_right.n3 185
R809 drain_right.n59 drain_right.n58 185
R810 drain_right.n61 drain_right.n60 185
R811 drain_right.n137 drain_right.n136 185
R812 drain_right.n135 drain_right.n134 185
R813 drain_right.n80 drain_right.n79 185
R814 drain_right.n129 drain_right.n128 185
R815 drain_right.n127 drain_right.n126 185
R816 drain_right.n84 drain_right.n83 185
R817 drain_right.n121 drain_right.n120 185
R818 drain_right.n119 drain_right.n86 185
R819 drain_right.n118 drain_right.n117 185
R820 drain_right.n89 drain_right.n87 185
R821 drain_right.n112 drain_right.n111 185
R822 drain_right.n110 drain_right.n109 185
R823 drain_right.n93 drain_right.n92 185
R824 drain_right.n104 drain_right.n103 185
R825 drain_right.n102 drain_right.n101 185
R826 drain_right.n97 drain_right.n96 185
R827 drain_right.n21 drain_right.t0 149.524
R828 drain_right.n98 drain_right.t2 149.524
R829 drain_right.n25 drain_right.n19 104.615
R830 drain_right.n26 drain_right.n25 104.615
R831 drain_right.n26 drain_right.n15 104.615
R832 drain_right.n33 drain_right.n15 104.615
R833 drain_right.n34 drain_right.n33 104.615
R834 drain_right.n34 drain_right.n11 104.615
R835 drain_right.n42 drain_right.n11 104.615
R836 drain_right.n43 drain_right.n42 104.615
R837 drain_right.n44 drain_right.n43 104.615
R838 drain_right.n44 drain_right.n7 104.615
R839 drain_right.n51 drain_right.n7 104.615
R840 drain_right.n52 drain_right.n51 104.615
R841 drain_right.n52 drain_right.n3 104.615
R842 drain_right.n59 drain_right.n3 104.615
R843 drain_right.n60 drain_right.n59 104.615
R844 drain_right.n136 drain_right.n135 104.615
R845 drain_right.n135 drain_right.n79 104.615
R846 drain_right.n128 drain_right.n79 104.615
R847 drain_right.n128 drain_right.n127 104.615
R848 drain_right.n127 drain_right.n83 104.615
R849 drain_right.n120 drain_right.n83 104.615
R850 drain_right.n120 drain_right.n119 104.615
R851 drain_right.n119 drain_right.n118 104.615
R852 drain_right.n118 drain_right.n87 104.615
R853 drain_right.n111 drain_right.n87 104.615
R854 drain_right.n111 drain_right.n110 104.615
R855 drain_right.n110 drain_right.n92 104.615
R856 drain_right.n103 drain_right.n92 104.615
R857 drain_right.n103 drain_right.n102 104.615
R858 drain_right.n102 drain_right.n96 104.615
R859 drain_right.n69 drain_right.n67 60.0525
R860 drain_right.n73 drain_right.n71 60.0525
R861 drain_right.n73 drain_right.n72 59.5527
R862 drain_right.n75 drain_right.n74 59.5527
R863 drain_right.n69 drain_right.n68 59.5525
R864 drain_right.n66 drain_right.n65 59.5525
R865 drain_right.t0 drain_right.n19 52.3082
R866 drain_right.t2 drain_right.n96 52.3082
R867 drain_right.n66 drain_right.n64 47.0369
R868 drain_right.n141 drain_right.n140 46.5369
R869 drain_right drain_right.n70 29.6888
R870 drain_right.n45 drain_right.n10 13.1884
R871 drain_right.n121 drain_right.n86 13.1884
R872 drain_right.n41 drain_right.n40 12.8005
R873 drain_right.n46 drain_right.n8 12.8005
R874 drain_right.n122 drain_right.n84 12.8005
R875 drain_right.n117 drain_right.n88 12.8005
R876 drain_right.n39 drain_right.n12 12.0247
R877 drain_right.n50 drain_right.n49 12.0247
R878 drain_right.n126 drain_right.n125 12.0247
R879 drain_right.n116 drain_right.n89 12.0247
R880 drain_right.n36 drain_right.n35 11.249
R881 drain_right.n53 drain_right.n6 11.249
R882 drain_right.n129 drain_right.n82 11.249
R883 drain_right.n113 drain_right.n112 11.249
R884 drain_right.n32 drain_right.n14 10.4732
R885 drain_right.n54 drain_right.n4 10.4732
R886 drain_right.n130 drain_right.n80 10.4732
R887 drain_right.n109 drain_right.n91 10.4732
R888 drain_right.n21 drain_right.n20 10.2747
R889 drain_right.n98 drain_right.n97 10.2747
R890 drain_right.n31 drain_right.n16 9.69747
R891 drain_right.n58 drain_right.n57 9.69747
R892 drain_right.n134 drain_right.n133 9.69747
R893 drain_right.n108 drain_right.n93 9.69747
R894 drain_right.n64 drain_right.n63 9.45567
R895 drain_right.n140 drain_right.n139 9.45567
R896 drain_right.n63 drain_right.n62 9.3005
R897 drain_right.n2 drain_right.n1 9.3005
R898 drain_right.n57 drain_right.n56 9.3005
R899 drain_right.n55 drain_right.n54 9.3005
R900 drain_right.n6 drain_right.n5 9.3005
R901 drain_right.n49 drain_right.n48 9.3005
R902 drain_right.n47 drain_right.n46 9.3005
R903 drain_right.n23 drain_right.n22 9.3005
R904 drain_right.n18 drain_right.n17 9.3005
R905 drain_right.n29 drain_right.n28 9.3005
R906 drain_right.n31 drain_right.n30 9.3005
R907 drain_right.n14 drain_right.n13 9.3005
R908 drain_right.n37 drain_right.n36 9.3005
R909 drain_right.n39 drain_right.n38 9.3005
R910 drain_right.n40 drain_right.n9 9.3005
R911 drain_right.n100 drain_right.n99 9.3005
R912 drain_right.n95 drain_right.n94 9.3005
R913 drain_right.n106 drain_right.n105 9.3005
R914 drain_right.n108 drain_right.n107 9.3005
R915 drain_right.n91 drain_right.n90 9.3005
R916 drain_right.n114 drain_right.n113 9.3005
R917 drain_right.n116 drain_right.n115 9.3005
R918 drain_right.n88 drain_right.n85 9.3005
R919 drain_right.n139 drain_right.n138 9.3005
R920 drain_right.n78 drain_right.n77 9.3005
R921 drain_right.n133 drain_right.n132 9.3005
R922 drain_right.n131 drain_right.n130 9.3005
R923 drain_right.n82 drain_right.n81 9.3005
R924 drain_right.n125 drain_right.n124 9.3005
R925 drain_right.n123 drain_right.n122 9.3005
R926 drain_right.n28 drain_right.n27 8.92171
R927 drain_right.n61 drain_right.n2 8.92171
R928 drain_right.n137 drain_right.n78 8.92171
R929 drain_right.n105 drain_right.n104 8.92171
R930 drain_right.n24 drain_right.n18 8.14595
R931 drain_right.n62 drain_right.n0 8.14595
R932 drain_right.n138 drain_right.n76 8.14595
R933 drain_right.n101 drain_right.n95 8.14595
R934 drain_right.n23 drain_right.n20 7.3702
R935 drain_right.n100 drain_right.n97 7.3702
R936 drain_right drain_right.n141 5.90322
R937 drain_right.n24 drain_right.n23 5.81868
R938 drain_right.n64 drain_right.n0 5.81868
R939 drain_right.n140 drain_right.n76 5.81868
R940 drain_right.n101 drain_right.n100 5.81868
R941 drain_right.n27 drain_right.n18 5.04292
R942 drain_right.n62 drain_right.n61 5.04292
R943 drain_right.n138 drain_right.n137 5.04292
R944 drain_right.n104 drain_right.n95 5.04292
R945 drain_right.n28 drain_right.n16 4.26717
R946 drain_right.n58 drain_right.n2 4.26717
R947 drain_right.n134 drain_right.n78 4.26717
R948 drain_right.n105 drain_right.n93 4.26717
R949 drain_right.n32 drain_right.n31 3.49141
R950 drain_right.n57 drain_right.n4 3.49141
R951 drain_right.n133 drain_right.n80 3.49141
R952 drain_right.n109 drain_right.n108 3.49141
R953 drain_right.n22 drain_right.n21 2.84303
R954 drain_right.n99 drain_right.n98 2.84303
R955 drain_right.n35 drain_right.n14 2.71565
R956 drain_right.n54 drain_right.n53 2.71565
R957 drain_right.n130 drain_right.n129 2.71565
R958 drain_right.n112 drain_right.n91 2.71565
R959 drain_right.n36 drain_right.n12 1.93989
R960 drain_right.n50 drain_right.n6 1.93989
R961 drain_right.n126 drain_right.n82 1.93989
R962 drain_right.n113 drain_right.n89 1.93989
R963 drain_right.n67 drain_right.t1 1.6505
R964 drain_right.n67 drain_right.t5 1.6505
R965 drain_right.n68 drain_right.t6 1.6505
R966 drain_right.n68 drain_right.t10 1.6505
R967 drain_right.n65 drain_right.t11 1.6505
R968 drain_right.n65 drain_right.t4 1.6505
R969 drain_right.n71 drain_right.t12 1.6505
R970 drain_right.n71 drain_right.t7 1.6505
R971 drain_right.n72 drain_right.t13 1.6505
R972 drain_right.n72 drain_right.t8 1.6505
R973 drain_right.n74 drain_right.t9 1.6505
R974 drain_right.n74 drain_right.t3 1.6505
R975 drain_right.n41 drain_right.n39 1.16414
R976 drain_right.n49 drain_right.n8 1.16414
R977 drain_right.n125 drain_right.n84 1.16414
R978 drain_right.n117 drain_right.n116 1.16414
R979 drain_right.n141 drain_right.n75 0.5005
R980 drain_right.n75 drain_right.n73 0.5005
R981 drain_right.n40 drain_right.n10 0.388379
R982 drain_right.n46 drain_right.n45 0.388379
R983 drain_right.n122 drain_right.n121 0.388379
R984 drain_right.n88 drain_right.n86 0.388379
R985 drain_right.n70 drain_right.n66 0.320154
R986 drain_right.n22 drain_right.n17 0.155672
R987 drain_right.n29 drain_right.n17 0.155672
R988 drain_right.n30 drain_right.n29 0.155672
R989 drain_right.n30 drain_right.n13 0.155672
R990 drain_right.n37 drain_right.n13 0.155672
R991 drain_right.n38 drain_right.n37 0.155672
R992 drain_right.n38 drain_right.n9 0.155672
R993 drain_right.n47 drain_right.n9 0.155672
R994 drain_right.n48 drain_right.n47 0.155672
R995 drain_right.n48 drain_right.n5 0.155672
R996 drain_right.n55 drain_right.n5 0.155672
R997 drain_right.n56 drain_right.n55 0.155672
R998 drain_right.n56 drain_right.n1 0.155672
R999 drain_right.n63 drain_right.n1 0.155672
R1000 drain_right.n139 drain_right.n77 0.155672
R1001 drain_right.n132 drain_right.n77 0.155672
R1002 drain_right.n132 drain_right.n131 0.155672
R1003 drain_right.n131 drain_right.n81 0.155672
R1004 drain_right.n124 drain_right.n81 0.155672
R1005 drain_right.n124 drain_right.n123 0.155672
R1006 drain_right.n123 drain_right.n85 0.155672
R1007 drain_right.n115 drain_right.n85 0.155672
R1008 drain_right.n115 drain_right.n114 0.155672
R1009 drain_right.n114 drain_right.n90 0.155672
R1010 drain_right.n107 drain_right.n90 0.155672
R1011 drain_right.n107 drain_right.n106 0.155672
R1012 drain_right.n106 drain_right.n94 0.155672
R1013 drain_right.n99 drain_right.n94 0.155672
R1014 drain_right.n70 drain_right.n69 0.070154
C0 minus drain_right 4.63424f
C1 source drain_right 30.406399f
C2 drain_left minus 0.171605f
C3 drain_left source 30.4176f
C4 source minus 4.25538f
C5 drain_right plus 0.314992f
C6 drain_left plus 4.78968f
C7 drain_left drain_right 0.841057f
C8 minus plus 5.2062f
C9 source plus 4.2701f
C10 drain_right a_n1644_n3288# 7.42719f
C11 drain_left a_n1644_n3288# 7.70168f
C12 source a_n1644_n3288# 6.123137f
C13 minus a_n1644_n3288# 6.38646f
C14 plus a_n1644_n3288# 8.40721f
C15 drain_right.n0 a_n1644_n3288# 0.043036f
C16 drain_right.n1 a_n1644_n3288# 0.032489f
C17 drain_right.n2 a_n1644_n3288# 0.017458f
C18 drain_right.n3 a_n1644_n3288# 0.041265f
C19 drain_right.n4 a_n1644_n3288# 0.018485f
C20 drain_right.n5 a_n1644_n3288# 0.032489f
C21 drain_right.n6 a_n1644_n3288# 0.017458f
C22 drain_right.n7 a_n1644_n3288# 0.041265f
C23 drain_right.n8 a_n1644_n3288# 0.018485f
C24 drain_right.n9 a_n1644_n3288# 0.032489f
C25 drain_right.n10 a_n1644_n3288# 0.017972f
C26 drain_right.n11 a_n1644_n3288# 0.041265f
C27 drain_right.n12 a_n1644_n3288# 0.018485f
C28 drain_right.n13 a_n1644_n3288# 0.032489f
C29 drain_right.n14 a_n1644_n3288# 0.017458f
C30 drain_right.n15 a_n1644_n3288# 0.041265f
C31 drain_right.n16 a_n1644_n3288# 0.018485f
C32 drain_right.n17 a_n1644_n3288# 0.032489f
C33 drain_right.n18 a_n1644_n3288# 0.017458f
C34 drain_right.n19 a_n1644_n3288# 0.030949f
C35 drain_right.n20 a_n1644_n3288# 0.029171f
C36 drain_right.t0 a_n1644_n3288# 0.069694f
C37 drain_right.n21 a_n1644_n3288# 0.234244f
C38 drain_right.n22 a_n1644_n3288# 1.63903f
C39 drain_right.n23 a_n1644_n3288# 0.017458f
C40 drain_right.n24 a_n1644_n3288# 0.018485f
C41 drain_right.n25 a_n1644_n3288# 0.041265f
C42 drain_right.n26 a_n1644_n3288# 0.041265f
C43 drain_right.n27 a_n1644_n3288# 0.018485f
C44 drain_right.n28 a_n1644_n3288# 0.017458f
C45 drain_right.n29 a_n1644_n3288# 0.032489f
C46 drain_right.n30 a_n1644_n3288# 0.032489f
C47 drain_right.n31 a_n1644_n3288# 0.017458f
C48 drain_right.n32 a_n1644_n3288# 0.018485f
C49 drain_right.n33 a_n1644_n3288# 0.041265f
C50 drain_right.n34 a_n1644_n3288# 0.041265f
C51 drain_right.n35 a_n1644_n3288# 0.018485f
C52 drain_right.n36 a_n1644_n3288# 0.017458f
C53 drain_right.n37 a_n1644_n3288# 0.032489f
C54 drain_right.n38 a_n1644_n3288# 0.032489f
C55 drain_right.n39 a_n1644_n3288# 0.017458f
C56 drain_right.n40 a_n1644_n3288# 0.017458f
C57 drain_right.n41 a_n1644_n3288# 0.018485f
C58 drain_right.n42 a_n1644_n3288# 0.041265f
C59 drain_right.n43 a_n1644_n3288# 0.041265f
C60 drain_right.n44 a_n1644_n3288# 0.041265f
C61 drain_right.n45 a_n1644_n3288# 0.017972f
C62 drain_right.n46 a_n1644_n3288# 0.017458f
C63 drain_right.n47 a_n1644_n3288# 0.032489f
C64 drain_right.n48 a_n1644_n3288# 0.032489f
C65 drain_right.n49 a_n1644_n3288# 0.017458f
C66 drain_right.n50 a_n1644_n3288# 0.018485f
C67 drain_right.n51 a_n1644_n3288# 0.041265f
C68 drain_right.n52 a_n1644_n3288# 0.041265f
C69 drain_right.n53 a_n1644_n3288# 0.018485f
C70 drain_right.n54 a_n1644_n3288# 0.017458f
C71 drain_right.n55 a_n1644_n3288# 0.032489f
C72 drain_right.n56 a_n1644_n3288# 0.032489f
C73 drain_right.n57 a_n1644_n3288# 0.017458f
C74 drain_right.n58 a_n1644_n3288# 0.018485f
C75 drain_right.n59 a_n1644_n3288# 0.041265f
C76 drain_right.n60 a_n1644_n3288# 0.084681f
C77 drain_right.n61 a_n1644_n3288# 0.018485f
C78 drain_right.n62 a_n1644_n3288# 0.017458f
C79 drain_right.n63 a_n1644_n3288# 0.069772f
C80 drain_right.n64 a_n1644_n3288# 0.070403f
C81 drain_right.t11 a_n1644_n3288# 0.308089f
C82 drain_right.t4 a_n1644_n3288# 0.308089f
C83 drain_right.n65 a_n1644_n3288# 2.74152f
C84 drain_right.n66 a_n1644_n3288# 0.471502f
C85 drain_right.t1 a_n1644_n3288# 0.308089f
C86 drain_right.t5 a_n1644_n3288# 0.308089f
C87 drain_right.n67 a_n1644_n3288# 2.74477f
C88 drain_right.t6 a_n1644_n3288# 0.308089f
C89 drain_right.t10 a_n1644_n3288# 0.308089f
C90 drain_right.n68 a_n1644_n3288# 2.74152f
C91 drain_right.n69 a_n1644_n3288# 0.730311f
C92 drain_right.n70 a_n1644_n3288# 1.44575f
C93 drain_right.t12 a_n1644_n3288# 0.308089f
C94 drain_right.t7 a_n1644_n3288# 0.308089f
C95 drain_right.n71 a_n1644_n3288# 2.74477f
C96 drain_right.t13 a_n1644_n3288# 0.308089f
C97 drain_right.t8 a_n1644_n3288# 0.308089f
C98 drain_right.n72 a_n1644_n3288# 2.74153f
C99 drain_right.n73 a_n1644_n3288# 0.764538f
C100 drain_right.t9 a_n1644_n3288# 0.308089f
C101 drain_right.t3 a_n1644_n3288# 0.308089f
C102 drain_right.n74 a_n1644_n3288# 2.74153f
C103 drain_right.n75 a_n1644_n3288# 0.377346f
C104 drain_right.n76 a_n1644_n3288# 0.043036f
C105 drain_right.n77 a_n1644_n3288# 0.032489f
C106 drain_right.n78 a_n1644_n3288# 0.017458f
C107 drain_right.n79 a_n1644_n3288# 0.041265f
C108 drain_right.n80 a_n1644_n3288# 0.018485f
C109 drain_right.n81 a_n1644_n3288# 0.032489f
C110 drain_right.n82 a_n1644_n3288# 0.017458f
C111 drain_right.n83 a_n1644_n3288# 0.041265f
C112 drain_right.n84 a_n1644_n3288# 0.018485f
C113 drain_right.n85 a_n1644_n3288# 0.032489f
C114 drain_right.n86 a_n1644_n3288# 0.017972f
C115 drain_right.n87 a_n1644_n3288# 0.041265f
C116 drain_right.n88 a_n1644_n3288# 0.017458f
C117 drain_right.n89 a_n1644_n3288# 0.018485f
C118 drain_right.n90 a_n1644_n3288# 0.032489f
C119 drain_right.n91 a_n1644_n3288# 0.017458f
C120 drain_right.n92 a_n1644_n3288# 0.041265f
C121 drain_right.n93 a_n1644_n3288# 0.018485f
C122 drain_right.n94 a_n1644_n3288# 0.032489f
C123 drain_right.n95 a_n1644_n3288# 0.017458f
C124 drain_right.n96 a_n1644_n3288# 0.030949f
C125 drain_right.n97 a_n1644_n3288# 0.029171f
C126 drain_right.t2 a_n1644_n3288# 0.069694f
C127 drain_right.n98 a_n1644_n3288# 0.234244f
C128 drain_right.n99 a_n1644_n3288# 1.63903f
C129 drain_right.n100 a_n1644_n3288# 0.017458f
C130 drain_right.n101 a_n1644_n3288# 0.018485f
C131 drain_right.n102 a_n1644_n3288# 0.041265f
C132 drain_right.n103 a_n1644_n3288# 0.041265f
C133 drain_right.n104 a_n1644_n3288# 0.018485f
C134 drain_right.n105 a_n1644_n3288# 0.017458f
C135 drain_right.n106 a_n1644_n3288# 0.032489f
C136 drain_right.n107 a_n1644_n3288# 0.032489f
C137 drain_right.n108 a_n1644_n3288# 0.017458f
C138 drain_right.n109 a_n1644_n3288# 0.018485f
C139 drain_right.n110 a_n1644_n3288# 0.041265f
C140 drain_right.n111 a_n1644_n3288# 0.041265f
C141 drain_right.n112 a_n1644_n3288# 0.018485f
C142 drain_right.n113 a_n1644_n3288# 0.017458f
C143 drain_right.n114 a_n1644_n3288# 0.032489f
C144 drain_right.n115 a_n1644_n3288# 0.032489f
C145 drain_right.n116 a_n1644_n3288# 0.017458f
C146 drain_right.n117 a_n1644_n3288# 0.018485f
C147 drain_right.n118 a_n1644_n3288# 0.041265f
C148 drain_right.n119 a_n1644_n3288# 0.041265f
C149 drain_right.n120 a_n1644_n3288# 0.041265f
C150 drain_right.n121 a_n1644_n3288# 0.017972f
C151 drain_right.n122 a_n1644_n3288# 0.017458f
C152 drain_right.n123 a_n1644_n3288# 0.032489f
C153 drain_right.n124 a_n1644_n3288# 0.032489f
C154 drain_right.n125 a_n1644_n3288# 0.017458f
C155 drain_right.n126 a_n1644_n3288# 0.018485f
C156 drain_right.n127 a_n1644_n3288# 0.041265f
C157 drain_right.n128 a_n1644_n3288# 0.041265f
C158 drain_right.n129 a_n1644_n3288# 0.018485f
C159 drain_right.n130 a_n1644_n3288# 0.017458f
C160 drain_right.n131 a_n1644_n3288# 0.032489f
C161 drain_right.n132 a_n1644_n3288# 0.032489f
C162 drain_right.n133 a_n1644_n3288# 0.017458f
C163 drain_right.n134 a_n1644_n3288# 0.018485f
C164 drain_right.n135 a_n1644_n3288# 0.041265f
C165 drain_right.n136 a_n1644_n3288# 0.084681f
C166 drain_right.n137 a_n1644_n3288# 0.018485f
C167 drain_right.n138 a_n1644_n3288# 0.017458f
C168 drain_right.n139 a_n1644_n3288# 0.069772f
C169 drain_right.n140 a_n1644_n3288# 0.069214f
C170 drain_right.n141 a_n1644_n3288# 0.379416f
C171 minus.n0 a_n1644_n3288# 0.052933f
C172 minus.t11 a_n1644_n3288# 0.453536f
C173 minus.t4 a_n1644_n3288# 0.448735f
C174 minus.t10 a_n1644_n3288# 0.448735f
C175 minus.t0 a_n1644_n3288# 0.448735f
C176 minus.n1 a_n1644_n3288# 0.19829f
C177 minus.n2 a_n1644_n3288# 0.113301f
C178 minus.t5 a_n1644_n3288# 0.448735f
C179 minus.t1 a_n1644_n3288# 0.448735f
C180 minus.t6 a_n1644_n3288# 0.453536f
C181 minus.n3 a_n1644_n3288# 0.195844f
C182 minus.n4 a_n1644_n3288# 0.18073f
C183 minus.n5 a_n1644_n3288# 0.02017f
C184 minus.n6 a_n1644_n3288# 0.18073f
C185 minus.n7 a_n1644_n3288# 0.02017f
C186 minus.n8 a_n1644_n3288# 0.052933f
C187 minus.n9 a_n1644_n3288# 0.052933f
C188 minus.n10 a_n1644_n3288# 0.052933f
C189 minus.n11 a_n1644_n3288# 0.02017f
C190 minus.n12 a_n1644_n3288# 0.18073f
C191 minus.n13 a_n1644_n3288# 0.02017f
C192 minus.n14 a_n1644_n3288# 0.18073f
C193 minus.n15 a_n1644_n3288# 0.195773f
C194 minus.n16 a_n1644_n3288# 1.79653f
C195 minus.n17 a_n1644_n3288# 0.052933f
C196 minus.t12 a_n1644_n3288# 0.448735f
C197 minus.t3 a_n1644_n3288# 0.448735f
C198 minus.t7 a_n1644_n3288# 0.448735f
C199 minus.n18 a_n1644_n3288# 0.19829f
C200 minus.n19 a_n1644_n3288# 0.113301f
C201 minus.t9 a_n1644_n3288# 0.448735f
C202 minus.t2 a_n1644_n3288# 0.448735f
C203 minus.t13 a_n1644_n3288# 0.453536f
C204 minus.n20 a_n1644_n3288# 0.195844f
C205 minus.n21 a_n1644_n3288# 0.18073f
C206 minus.n22 a_n1644_n3288# 0.02017f
C207 minus.n23 a_n1644_n3288# 0.18073f
C208 minus.n24 a_n1644_n3288# 0.02017f
C209 minus.n25 a_n1644_n3288# 0.052933f
C210 minus.n26 a_n1644_n3288# 0.052933f
C211 minus.n27 a_n1644_n3288# 0.052933f
C212 minus.n28 a_n1644_n3288# 0.02017f
C213 minus.n29 a_n1644_n3288# 0.18073f
C214 minus.n30 a_n1644_n3288# 0.02017f
C215 minus.n31 a_n1644_n3288# 0.18073f
C216 minus.t8 a_n1644_n3288# 0.453536f
C217 minus.n32 a_n1644_n3288# 0.195773f
C218 minus.n33 a_n1644_n3288# 0.339968f
C219 minus.n34 a_n1644_n3288# 2.19017f
C220 source.n0 a_n1644_n3288# 0.044615f
C221 source.n1 a_n1644_n3288# 0.033681f
C222 source.n2 a_n1644_n3288# 0.018099f
C223 source.n3 a_n1644_n3288# 0.042779f
C224 source.n4 a_n1644_n3288# 0.019163f
C225 source.n5 a_n1644_n3288# 0.033681f
C226 source.n6 a_n1644_n3288# 0.018099f
C227 source.n7 a_n1644_n3288# 0.042779f
C228 source.n8 a_n1644_n3288# 0.019163f
C229 source.n9 a_n1644_n3288# 0.033681f
C230 source.n10 a_n1644_n3288# 0.018631f
C231 source.n11 a_n1644_n3288# 0.042779f
C232 source.n12 a_n1644_n3288# 0.018099f
C233 source.n13 a_n1644_n3288# 0.019163f
C234 source.n14 a_n1644_n3288# 0.033681f
C235 source.n15 a_n1644_n3288# 0.018099f
C236 source.n16 a_n1644_n3288# 0.042779f
C237 source.n17 a_n1644_n3288# 0.019163f
C238 source.n18 a_n1644_n3288# 0.033681f
C239 source.n19 a_n1644_n3288# 0.018099f
C240 source.n20 a_n1644_n3288# 0.032084f
C241 source.n21 a_n1644_n3288# 0.030241f
C242 source.t22 a_n1644_n3288# 0.07225f
C243 source.n22 a_n1644_n3288# 0.242835f
C244 source.n23 a_n1644_n3288# 1.69914f
C245 source.n24 a_n1644_n3288# 0.018099f
C246 source.n25 a_n1644_n3288# 0.019163f
C247 source.n26 a_n1644_n3288# 0.042779f
C248 source.n27 a_n1644_n3288# 0.042779f
C249 source.n28 a_n1644_n3288# 0.019163f
C250 source.n29 a_n1644_n3288# 0.018099f
C251 source.n30 a_n1644_n3288# 0.033681f
C252 source.n31 a_n1644_n3288# 0.033681f
C253 source.n32 a_n1644_n3288# 0.018099f
C254 source.n33 a_n1644_n3288# 0.019163f
C255 source.n34 a_n1644_n3288# 0.042779f
C256 source.n35 a_n1644_n3288# 0.042779f
C257 source.n36 a_n1644_n3288# 0.019163f
C258 source.n37 a_n1644_n3288# 0.018099f
C259 source.n38 a_n1644_n3288# 0.033681f
C260 source.n39 a_n1644_n3288# 0.033681f
C261 source.n40 a_n1644_n3288# 0.018099f
C262 source.n41 a_n1644_n3288# 0.019163f
C263 source.n42 a_n1644_n3288# 0.042779f
C264 source.n43 a_n1644_n3288# 0.042779f
C265 source.n44 a_n1644_n3288# 0.042779f
C266 source.n45 a_n1644_n3288# 0.018631f
C267 source.n46 a_n1644_n3288# 0.018099f
C268 source.n47 a_n1644_n3288# 0.033681f
C269 source.n48 a_n1644_n3288# 0.033681f
C270 source.n49 a_n1644_n3288# 0.018099f
C271 source.n50 a_n1644_n3288# 0.019163f
C272 source.n51 a_n1644_n3288# 0.042779f
C273 source.n52 a_n1644_n3288# 0.042779f
C274 source.n53 a_n1644_n3288# 0.019163f
C275 source.n54 a_n1644_n3288# 0.018099f
C276 source.n55 a_n1644_n3288# 0.033681f
C277 source.n56 a_n1644_n3288# 0.033681f
C278 source.n57 a_n1644_n3288# 0.018099f
C279 source.n58 a_n1644_n3288# 0.019163f
C280 source.n59 a_n1644_n3288# 0.042779f
C281 source.n60 a_n1644_n3288# 0.087786f
C282 source.n61 a_n1644_n3288# 0.019163f
C283 source.n62 a_n1644_n3288# 0.018099f
C284 source.n63 a_n1644_n3288# 0.07233f
C285 source.n64 a_n1644_n3288# 0.048449f
C286 source.n65 a_n1644_n3288# 1.34781f
C287 source.t21 a_n1644_n3288# 0.319388f
C288 source.t15 a_n1644_n3288# 0.319388f
C289 source.n66 a_n1644_n3288# 2.73461f
C290 source.n67 a_n1644_n3288# 0.452872f
C291 source.t20 a_n1644_n3288# 0.319388f
C292 source.t27 a_n1644_n3288# 0.319388f
C293 source.n68 a_n1644_n3288# 2.73461f
C294 source.n69 a_n1644_n3288# 0.452872f
C295 source.t24 a_n1644_n3288# 0.319388f
C296 source.t26 a_n1644_n3288# 0.319388f
C297 source.n70 a_n1644_n3288# 2.73461f
C298 source.n71 a_n1644_n3288# 0.476729f
C299 source.n72 a_n1644_n3288# 0.044615f
C300 source.n73 a_n1644_n3288# 0.033681f
C301 source.n74 a_n1644_n3288# 0.018099f
C302 source.n75 a_n1644_n3288# 0.042779f
C303 source.n76 a_n1644_n3288# 0.019163f
C304 source.n77 a_n1644_n3288# 0.033681f
C305 source.n78 a_n1644_n3288# 0.018099f
C306 source.n79 a_n1644_n3288# 0.042779f
C307 source.n80 a_n1644_n3288# 0.019163f
C308 source.n81 a_n1644_n3288# 0.033681f
C309 source.n82 a_n1644_n3288# 0.018631f
C310 source.n83 a_n1644_n3288# 0.042779f
C311 source.n84 a_n1644_n3288# 0.018099f
C312 source.n85 a_n1644_n3288# 0.019163f
C313 source.n86 a_n1644_n3288# 0.033681f
C314 source.n87 a_n1644_n3288# 0.018099f
C315 source.n88 a_n1644_n3288# 0.042779f
C316 source.n89 a_n1644_n3288# 0.019163f
C317 source.n90 a_n1644_n3288# 0.033681f
C318 source.n91 a_n1644_n3288# 0.018099f
C319 source.n92 a_n1644_n3288# 0.032084f
C320 source.n93 a_n1644_n3288# 0.030241f
C321 source.t5 a_n1644_n3288# 0.07225f
C322 source.n94 a_n1644_n3288# 0.242835f
C323 source.n95 a_n1644_n3288# 1.69914f
C324 source.n96 a_n1644_n3288# 0.018099f
C325 source.n97 a_n1644_n3288# 0.019163f
C326 source.n98 a_n1644_n3288# 0.042779f
C327 source.n99 a_n1644_n3288# 0.042779f
C328 source.n100 a_n1644_n3288# 0.019163f
C329 source.n101 a_n1644_n3288# 0.018099f
C330 source.n102 a_n1644_n3288# 0.033681f
C331 source.n103 a_n1644_n3288# 0.033681f
C332 source.n104 a_n1644_n3288# 0.018099f
C333 source.n105 a_n1644_n3288# 0.019163f
C334 source.n106 a_n1644_n3288# 0.042779f
C335 source.n107 a_n1644_n3288# 0.042779f
C336 source.n108 a_n1644_n3288# 0.019163f
C337 source.n109 a_n1644_n3288# 0.018099f
C338 source.n110 a_n1644_n3288# 0.033681f
C339 source.n111 a_n1644_n3288# 0.033681f
C340 source.n112 a_n1644_n3288# 0.018099f
C341 source.n113 a_n1644_n3288# 0.019163f
C342 source.n114 a_n1644_n3288# 0.042779f
C343 source.n115 a_n1644_n3288# 0.042779f
C344 source.n116 a_n1644_n3288# 0.042779f
C345 source.n117 a_n1644_n3288# 0.018631f
C346 source.n118 a_n1644_n3288# 0.018099f
C347 source.n119 a_n1644_n3288# 0.033681f
C348 source.n120 a_n1644_n3288# 0.033681f
C349 source.n121 a_n1644_n3288# 0.018099f
C350 source.n122 a_n1644_n3288# 0.019163f
C351 source.n123 a_n1644_n3288# 0.042779f
C352 source.n124 a_n1644_n3288# 0.042779f
C353 source.n125 a_n1644_n3288# 0.019163f
C354 source.n126 a_n1644_n3288# 0.018099f
C355 source.n127 a_n1644_n3288# 0.033681f
C356 source.n128 a_n1644_n3288# 0.033681f
C357 source.n129 a_n1644_n3288# 0.018099f
C358 source.n130 a_n1644_n3288# 0.019163f
C359 source.n131 a_n1644_n3288# 0.042779f
C360 source.n132 a_n1644_n3288# 0.087786f
C361 source.n133 a_n1644_n3288# 0.019163f
C362 source.n134 a_n1644_n3288# 0.018099f
C363 source.n135 a_n1644_n3288# 0.07233f
C364 source.n136 a_n1644_n3288# 0.048449f
C365 source.n137 a_n1644_n3288# 0.15804f
C366 source.t3 a_n1644_n3288# 0.319388f
C367 source.t0 a_n1644_n3288# 0.319388f
C368 source.n138 a_n1644_n3288# 2.73461f
C369 source.n139 a_n1644_n3288# 0.452872f
C370 source.t10 a_n1644_n3288# 0.319388f
C371 source.t9 a_n1644_n3288# 0.319388f
C372 source.n140 a_n1644_n3288# 2.73461f
C373 source.n141 a_n1644_n3288# 0.452872f
C374 source.t4 a_n1644_n3288# 0.319388f
C375 source.t7 a_n1644_n3288# 0.319388f
C376 source.n142 a_n1644_n3288# 2.73461f
C377 source.n143 a_n1644_n3288# 2.24869f
C378 source.t19 a_n1644_n3288# 0.319388f
C379 source.t17 a_n1644_n3288# 0.319388f
C380 source.n144 a_n1644_n3288# 2.73459f
C381 source.n145 a_n1644_n3288# 2.2487f
C382 source.t25 a_n1644_n3288# 0.319388f
C383 source.t14 a_n1644_n3288# 0.319388f
C384 source.n146 a_n1644_n3288# 2.73459f
C385 source.n147 a_n1644_n3288# 0.452888f
C386 source.t23 a_n1644_n3288# 0.319388f
C387 source.t18 a_n1644_n3288# 0.319388f
C388 source.n148 a_n1644_n3288# 2.73459f
C389 source.n149 a_n1644_n3288# 0.452888f
C390 source.n150 a_n1644_n3288# 0.044615f
C391 source.n151 a_n1644_n3288# 0.033681f
C392 source.n152 a_n1644_n3288# 0.018099f
C393 source.n153 a_n1644_n3288# 0.042779f
C394 source.n154 a_n1644_n3288# 0.019163f
C395 source.n155 a_n1644_n3288# 0.033681f
C396 source.n156 a_n1644_n3288# 0.018099f
C397 source.n157 a_n1644_n3288# 0.042779f
C398 source.n158 a_n1644_n3288# 0.019163f
C399 source.n159 a_n1644_n3288# 0.033681f
C400 source.n160 a_n1644_n3288# 0.018631f
C401 source.n161 a_n1644_n3288# 0.042779f
C402 source.n162 a_n1644_n3288# 0.019163f
C403 source.n163 a_n1644_n3288# 0.033681f
C404 source.n164 a_n1644_n3288# 0.018099f
C405 source.n165 a_n1644_n3288# 0.042779f
C406 source.n166 a_n1644_n3288# 0.019163f
C407 source.n167 a_n1644_n3288# 0.033681f
C408 source.n168 a_n1644_n3288# 0.018099f
C409 source.n169 a_n1644_n3288# 0.032084f
C410 source.n170 a_n1644_n3288# 0.030241f
C411 source.t16 a_n1644_n3288# 0.07225f
C412 source.n171 a_n1644_n3288# 0.242835f
C413 source.n172 a_n1644_n3288# 1.69914f
C414 source.n173 a_n1644_n3288# 0.018099f
C415 source.n174 a_n1644_n3288# 0.019163f
C416 source.n175 a_n1644_n3288# 0.042779f
C417 source.n176 a_n1644_n3288# 0.042779f
C418 source.n177 a_n1644_n3288# 0.019163f
C419 source.n178 a_n1644_n3288# 0.018099f
C420 source.n179 a_n1644_n3288# 0.033681f
C421 source.n180 a_n1644_n3288# 0.033681f
C422 source.n181 a_n1644_n3288# 0.018099f
C423 source.n182 a_n1644_n3288# 0.019163f
C424 source.n183 a_n1644_n3288# 0.042779f
C425 source.n184 a_n1644_n3288# 0.042779f
C426 source.n185 a_n1644_n3288# 0.019163f
C427 source.n186 a_n1644_n3288# 0.018099f
C428 source.n187 a_n1644_n3288# 0.033681f
C429 source.n188 a_n1644_n3288# 0.033681f
C430 source.n189 a_n1644_n3288# 0.018099f
C431 source.n190 a_n1644_n3288# 0.018099f
C432 source.n191 a_n1644_n3288# 0.019163f
C433 source.n192 a_n1644_n3288# 0.042779f
C434 source.n193 a_n1644_n3288# 0.042779f
C435 source.n194 a_n1644_n3288# 0.042779f
C436 source.n195 a_n1644_n3288# 0.018631f
C437 source.n196 a_n1644_n3288# 0.018099f
C438 source.n197 a_n1644_n3288# 0.033681f
C439 source.n198 a_n1644_n3288# 0.033681f
C440 source.n199 a_n1644_n3288# 0.018099f
C441 source.n200 a_n1644_n3288# 0.019163f
C442 source.n201 a_n1644_n3288# 0.042779f
C443 source.n202 a_n1644_n3288# 0.042779f
C444 source.n203 a_n1644_n3288# 0.019163f
C445 source.n204 a_n1644_n3288# 0.018099f
C446 source.n205 a_n1644_n3288# 0.033681f
C447 source.n206 a_n1644_n3288# 0.033681f
C448 source.n207 a_n1644_n3288# 0.018099f
C449 source.n208 a_n1644_n3288# 0.019163f
C450 source.n209 a_n1644_n3288# 0.042779f
C451 source.n210 a_n1644_n3288# 0.087786f
C452 source.n211 a_n1644_n3288# 0.019163f
C453 source.n212 a_n1644_n3288# 0.018099f
C454 source.n213 a_n1644_n3288# 0.07233f
C455 source.n214 a_n1644_n3288# 0.048449f
C456 source.n215 a_n1644_n3288# 0.15804f
C457 source.t13 a_n1644_n3288# 0.319388f
C458 source.t11 a_n1644_n3288# 0.319388f
C459 source.n216 a_n1644_n3288# 2.73459f
C460 source.n217 a_n1644_n3288# 0.476746f
C461 source.t8 a_n1644_n3288# 0.319388f
C462 source.t12 a_n1644_n3288# 0.319388f
C463 source.n218 a_n1644_n3288# 2.73459f
C464 source.n219 a_n1644_n3288# 0.452888f
C465 source.t2 a_n1644_n3288# 0.319388f
C466 source.t1 a_n1644_n3288# 0.319388f
C467 source.n220 a_n1644_n3288# 2.73459f
C468 source.n221 a_n1644_n3288# 0.452888f
C469 source.n222 a_n1644_n3288# 0.044615f
C470 source.n223 a_n1644_n3288# 0.033681f
C471 source.n224 a_n1644_n3288# 0.018099f
C472 source.n225 a_n1644_n3288# 0.042779f
C473 source.n226 a_n1644_n3288# 0.019163f
C474 source.n227 a_n1644_n3288# 0.033681f
C475 source.n228 a_n1644_n3288# 0.018099f
C476 source.n229 a_n1644_n3288# 0.042779f
C477 source.n230 a_n1644_n3288# 0.019163f
C478 source.n231 a_n1644_n3288# 0.033681f
C479 source.n232 a_n1644_n3288# 0.018631f
C480 source.n233 a_n1644_n3288# 0.042779f
C481 source.n234 a_n1644_n3288# 0.019163f
C482 source.n235 a_n1644_n3288# 0.033681f
C483 source.n236 a_n1644_n3288# 0.018099f
C484 source.n237 a_n1644_n3288# 0.042779f
C485 source.n238 a_n1644_n3288# 0.019163f
C486 source.n239 a_n1644_n3288# 0.033681f
C487 source.n240 a_n1644_n3288# 0.018099f
C488 source.n241 a_n1644_n3288# 0.032084f
C489 source.n242 a_n1644_n3288# 0.030241f
C490 source.t6 a_n1644_n3288# 0.07225f
C491 source.n243 a_n1644_n3288# 0.242835f
C492 source.n244 a_n1644_n3288# 1.69914f
C493 source.n245 a_n1644_n3288# 0.018099f
C494 source.n246 a_n1644_n3288# 0.019163f
C495 source.n247 a_n1644_n3288# 0.042779f
C496 source.n248 a_n1644_n3288# 0.042779f
C497 source.n249 a_n1644_n3288# 0.019163f
C498 source.n250 a_n1644_n3288# 0.018099f
C499 source.n251 a_n1644_n3288# 0.033681f
C500 source.n252 a_n1644_n3288# 0.033681f
C501 source.n253 a_n1644_n3288# 0.018099f
C502 source.n254 a_n1644_n3288# 0.019163f
C503 source.n255 a_n1644_n3288# 0.042779f
C504 source.n256 a_n1644_n3288# 0.042779f
C505 source.n257 a_n1644_n3288# 0.019163f
C506 source.n258 a_n1644_n3288# 0.018099f
C507 source.n259 a_n1644_n3288# 0.033681f
C508 source.n260 a_n1644_n3288# 0.033681f
C509 source.n261 a_n1644_n3288# 0.018099f
C510 source.n262 a_n1644_n3288# 0.018099f
C511 source.n263 a_n1644_n3288# 0.019163f
C512 source.n264 a_n1644_n3288# 0.042779f
C513 source.n265 a_n1644_n3288# 0.042779f
C514 source.n266 a_n1644_n3288# 0.042779f
C515 source.n267 a_n1644_n3288# 0.018631f
C516 source.n268 a_n1644_n3288# 0.018099f
C517 source.n269 a_n1644_n3288# 0.033681f
C518 source.n270 a_n1644_n3288# 0.033681f
C519 source.n271 a_n1644_n3288# 0.018099f
C520 source.n272 a_n1644_n3288# 0.019163f
C521 source.n273 a_n1644_n3288# 0.042779f
C522 source.n274 a_n1644_n3288# 0.042779f
C523 source.n275 a_n1644_n3288# 0.019163f
C524 source.n276 a_n1644_n3288# 0.018099f
C525 source.n277 a_n1644_n3288# 0.033681f
C526 source.n278 a_n1644_n3288# 0.033681f
C527 source.n279 a_n1644_n3288# 0.018099f
C528 source.n280 a_n1644_n3288# 0.019163f
C529 source.n281 a_n1644_n3288# 0.042779f
C530 source.n282 a_n1644_n3288# 0.087786f
C531 source.n283 a_n1644_n3288# 0.019163f
C532 source.n284 a_n1644_n3288# 0.018099f
C533 source.n285 a_n1644_n3288# 0.07233f
C534 source.n286 a_n1644_n3288# 0.048449f
C535 source.n287 a_n1644_n3288# 0.317293f
C536 source.n288 a_n1644_n3288# 2.11032f
C537 drain_left.n0 a_n1644_n3288# 0.043126f
C538 drain_left.n1 a_n1644_n3288# 0.032557f
C539 drain_left.n2 a_n1644_n3288# 0.017495f
C540 drain_left.n3 a_n1644_n3288# 0.041351f
C541 drain_left.n4 a_n1644_n3288# 0.018524f
C542 drain_left.n5 a_n1644_n3288# 0.032557f
C543 drain_left.n6 a_n1644_n3288# 0.017495f
C544 drain_left.n7 a_n1644_n3288# 0.041351f
C545 drain_left.n8 a_n1644_n3288# 0.018524f
C546 drain_left.n9 a_n1644_n3288# 0.032557f
C547 drain_left.n10 a_n1644_n3288# 0.018009f
C548 drain_left.n11 a_n1644_n3288# 0.041351f
C549 drain_left.n12 a_n1644_n3288# 0.018524f
C550 drain_left.n13 a_n1644_n3288# 0.032557f
C551 drain_left.n14 a_n1644_n3288# 0.017495f
C552 drain_left.n15 a_n1644_n3288# 0.041351f
C553 drain_left.n16 a_n1644_n3288# 0.018524f
C554 drain_left.n17 a_n1644_n3288# 0.032557f
C555 drain_left.n18 a_n1644_n3288# 0.017495f
C556 drain_left.n19 a_n1644_n3288# 0.031013f
C557 drain_left.n20 a_n1644_n3288# 0.029232f
C558 drain_left.t3 a_n1644_n3288# 0.069839f
C559 drain_left.n21 a_n1644_n3288# 0.234731f
C560 drain_left.n22 a_n1644_n3288# 1.64243f
C561 drain_left.n23 a_n1644_n3288# 0.017495f
C562 drain_left.n24 a_n1644_n3288# 0.018524f
C563 drain_left.n25 a_n1644_n3288# 0.041351f
C564 drain_left.n26 a_n1644_n3288# 0.041351f
C565 drain_left.n27 a_n1644_n3288# 0.018524f
C566 drain_left.n28 a_n1644_n3288# 0.017495f
C567 drain_left.n29 a_n1644_n3288# 0.032557f
C568 drain_left.n30 a_n1644_n3288# 0.032557f
C569 drain_left.n31 a_n1644_n3288# 0.017495f
C570 drain_left.n32 a_n1644_n3288# 0.018524f
C571 drain_left.n33 a_n1644_n3288# 0.041351f
C572 drain_left.n34 a_n1644_n3288# 0.041351f
C573 drain_left.n35 a_n1644_n3288# 0.018524f
C574 drain_left.n36 a_n1644_n3288# 0.017495f
C575 drain_left.n37 a_n1644_n3288# 0.032557f
C576 drain_left.n38 a_n1644_n3288# 0.032557f
C577 drain_left.n39 a_n1644_n3288# 0.017495f
C578 drain_left.n40 a_n1644_n3288# 0.017495f
C579 drain_left.n41 a_n1644_n3288# 0.018524f
C580 drain_left.n42 a_n1644_n3288# 0.041351f
C581 drain_left.n43 a_n1644_n3288# 0.041351f
C582 drain_left.n44 a_n1644_n3288# 0.041351f
C583 drain_left.n45 a_n1644_n3288# 0.018009f
C584 drain_left.n46 a_n1644_n3288# 0.017495f
C585 drain_left.n47 a_n1644_n3288# 0.032557f
C586 drain_left.n48 a_n1644_n3288# 0.032557f
C587 drain_left.n49 a_n1644_n3288# 0.017495f
C588 drain_left.n50 a_n1644_n3288# 0.018524f
C589 drain_left.n51 a_n1644_n3288# 0.041351f
C590 drain_left.n52 a_n1644_n3288# 0.041351f
C591 drain_left.n53 a_n1644_n3288# 0.018524f
C592 drain_left.n54 a_n1644_n3288# 0.017495f
C593 drain_left.n55 a_n1644_n3288# 0.032557f
C594 drain_left.n56 a_n1644_n3288# 0.032557f
C595 drain_left.n57 a_n1644_n3288# 0.017495f
C596 drain_left.n58 a_n1644_n3288# 0.018524f
C597 drain_left.n59 a_n1644_n3288# 0.041351f
C598 drain_left.n60 a_n1644_n3288# 0.084856f
C599 drain_left.n61 a_n1644_n3288# 0.018524f
C600 drain_left.n62 a_n1644_n3288# 0.017495f
C601 drain_left.n63 a_n1644_n3288# 0.069916f
C602 drain_left.n64 a_n1644_n3288# 0.070549f
C603 drain_left.t11 a_n1644_n3288# 0.308728f
C604 drain_left.t12 a_n1644_n3288# 0.308728f
C605 drain_left.n65 a_n1644_n3288# 2.74721f
C606 drain_left.n66 a_n1644_n3288# 0.472481f
C607 drain_left.t9 a_n1644_n3288# 0.308728f
C608 drain_left.t5 a_n1644_n3288# 0.308728f
C609 drain_left.n67 a_n1644_n3288# 2.75046f
C610 drain_left.t0 a_n1644_n3288# 0.308728f
C611 drain_left.t7 a_n1644_n3288# 0.308728f
C612 drain_left.n68 a_n1644_n3288# 2.74721f
C613 drain_left.n69 a_n1644_n3288# 0.731826f
C614 drain_left.n70 a_n1644_n3288# 1.51651f
C615 drain_left.n71 a_n1644_n3288# 0.043126f
C616 drain_left.n72 a_n1644_n3288# 0.032557f
C617 drain_left.n73 a_n1644_n3288# 0.017495f
C618 drain_left.n74 a_n1644_n3288# 0.041351f
C619 drain_left.n75 a_n1644_n3288# 0.018524f
C620 drain_left.n76 a_n1644_n3288# 0.032557f
C621 drain_left.n77 a_n1644_n3288# 0.017495f
C622 drain_left.n78 a_n1644_n3288# 0.041351f
C623 drain_left.n79 a_n1644_n3288# 0.018524f
C624 drain_left.n80 a_n1644_n3288# 0.032557f
C625 drain_left.n81 a_n1644_n3288# 0.018009f
C626 drain_left.n82 a_n1644_n3288# 0.041351f
C627 drain_left.n83 a_n1644_n3288# 0.017495f
C628 drain_left.n84 a_n1644_n3288# 0.018524f
C629 drain_left.n85 a_n1644_n3288# 0.032557f
C630 drain_left.n86 a_n1644_n3288# 0.017495f
C631 drain_left.n87 a_n1644_n3288# 0.041351f
C632 drain_left.n88 a_n1644_n3288# 0.018524f
C633 drain_left.n89 a_n1644_n3288# 0.032557f
C634 drain_left.n90 a_n1644_n3288# 0.017495f
C635 drain_left.n91 a_n1644_n3288# 0.031013f
C636 drain_left.n92 a_n1644_n3288# 0.029232f
C637 drain_left.t8 a_n1644_n3288# 0.069839f
C638 drain_left.n93 a_n1644_n3288# 0.234731f
C639 drain_left.n94 a_n1644_n3288# 1.64243f
C640 drain_left.n95 a_n1644_n3288# 0.017495f
C641 drain_left.n96 a_n1644_n3288# 0.018524f
C642 drain_left.n97 a_n1644_n3288# 0.041351f
C643 drain_left.n98 a_n1644_n3288# 0.041351f
C644 drain_left.n99 a_n1644_n3288# 0.018524f
C645 drain_left.n100 a_n1644_n3288# 0.017495f
C646 drain_left.n101 a_n1644_n3288# 0.032557f
C647 drain_left.n102 a_n1644_n3288# 0.032557f
C648 drain_left.n103 a_n1644_n3288# 0.017495f
C649 drain_left.n104 a_n1644_n3288# 0.018524f
C650 drain_left.n105 a_n1644_n3288# 0.041351f
C651 drain_left.n106 a_n1644_n3288# 0.041351f
C652 drain_left.n107 a_n1644_n3288# 0.018524f
C653 drain_left.n108 a_n1644_n3288# 0.017495f
C654 drain_left.n109 a_n1644_n3288# 0.032557f
C655 drain_left.n110 a_n1644_n3288# 0.032557f
C656 drain_left.n111 a_n1644_n3288# 0.017495f
C657 drain_left.n112 a_n1644_n3288# 0.018524f
C658 drain_left.n113 a_n1644_n3288# 0.041351f
C659 drain_left.n114 a_n1644_n3288# 0.041351f
C660 drain_left.n115 a_n1644_n3288# 0.041351f
C661 drain_left.n116 a_n1644_n3288# 0.018009f
C662 drain_left.n117 a_n1644_n3288# 0.017495f
C663 drain_left.n118 a_n1644_n3288# 0.032557f
C664 drain_left.n119 a_n1644_n3288# 0.032557f
C665 drain_left.n120 a_n1644_n3288# 0.017495f
C666 drain_left.n121 a_n1644_n3288# 0.018524f
C667 drain_left.n122 a_n1644_n3288# 0.041351f
C668 drain_left.n123 a_n1644_n3288# 0.041351f
C669 drain_left.n124 a_n1644_n3288# 0.018524f
C670 drain_left.n125 a_n1644_n3288# 0.017495f
C671 drain_left.n126 a_n1644_n3288# 0.032557f
C672 drain_left.n127 a_n1644_n3288# 0.032557f
C673 drain_left.n128 a_n1644_n3288# 0.017495f
C674 drain_left.n129 a_n1644_n3288# 0.018524f
C675 drain_left.n130 a_n1644_n3288# 0.041351f
C676 drain_left.n131 a_n1644_n3288# 0.084856f
C677 drain_left.n132 a_n1644_n3288# 0.018524f
C678 drain_left.n133 a_n1644_n3288# 0.017495f
C679 drain_left.n134 a_n1644_n3288# 0.069916f
C680 drain_left.n135 a_n1644_n3288# 0.070549f
C681 drain_left.t2 a_n1644_n3288# 0.308728f
C682 drain_left.t1 a_n1644_n3288# 0.308728f
C683 drain_left.n136 a_n1644_n3288# 2.74722f
C684 drain_left.n137 a_n1644_n3288# 0.489027f
C685 drain_left.t4 a_n1644_n3288# 0.308728f
C686 drain_left.t13 a_n1644_n3288# 0.308728f
C687 drain_left.n138 a_n1644_n3288# 2.74722f
C688 drain_left.n139 a_n1644_n3288# 0.378129f
C689 drain_left.t10 a_n1644_n3288# 0.308728f
C690 drain_left.t6 a_n1644_n3288# 0.308728f
C691 drain_left.n140 a_n1644_n3288# 2.74721f
C692 drain_left.n141 a_n1644_n3288# 0.646874f
C693 plus.n0 a_n1644_n3288# 0.054094f
C694 plus.t12 a_n1644_n3288# 0.458581f
C695 plus.t6 a_n1644_n3288# 0.458581f
C696 plus.t0 a_n1644_n3288# 0.458581f
C697 plus.n1 a_n1644_n3288# 0.202641f
C698 plus.n2 a_n1644_n3288# 0.115787f
C699 plus.t7 a_n1644_n3288# 0.458581f
C700 plus.t1 a_n1644_n3288# 0.458581f
C701 plus.t3 a_n1644_n3288# 0.463488f
C702 plus.n3 a_n1644_n3288# 0.200141f
C703 plus.n4 a_n1644_n3288# 0.184696f
C704 plus.n5 a_n1644_n3288# 0.020613f
C705 plus.n6 a_n1644_n3288# 0.184696f
C706 plus.n7 a_n1644_n3288# 0.020613f
C707 plus.n8 a_n1644_n3288# 0.054094f
C708 plus.n9 a_n1644_n3288# 0.054094f
C709 plus.n10 a_n1644_n3288# 0.054094f
C710 plus.n11 a_n1644_n3288# 0.020613f
C711 plus.n12 a_n1644_n3288# 0.184696f
C712 plus.n13 a_n1644_n3288# 0.020613f
C713 plus.n14 a_n1644_n3288# 0.184696f
C714 plus.t5 a_n1644_n3288# 0.463488f
C715 plus.n15 a_n1644_n3288# 0.200069f
C716 plus.n16 a_n1644_n3288# 0.598919f
C717 plus.n17 a_n1644_n3288# 0.054094f
C718 plus.t8 a_n1644_n3288# 0.463488f
C719 plus.t10 a_n1644_n3288# 0.458581f
C720 plus.t2 a_n1644_n3288# 0.458581f
C721 plus.t13 a_n1644_n3288# 0.458581f
C722 plus.n18 a_n1644_n3288# 0.202641f
C723 plus.n19 a_n1644_n3288# 0.115787f
C724 plus.t4 a_n1644_n3288# 0.458581f
C725 plus.t9 a_n1644_n3288# 0.458581f
C726 plus.t11 a_n1644_n3288# 0.463488f
C727 plus.n20 a_n1644_n3288# 0.200141f
C728 plus.n21 a_n1644_n3288# 0.184696f
C729 plus.n22 a_n1644_n3288# 0.020613f
C730 plus.n23 a_n1644_n3288# 0.184696f
C731 plus.n24 a_n1644_n3288# 0.020613f
C732 plus.n25 a_n1644_n3288# 0.054094f
C733 plus.n26 a_n1644_n3288# 0.054094f
C734 plus.n27 a_n1644_n3288# 0.054094f
C735 plus.n28 a_n1644_n3288# 0.020613f
C736 plus.n29 a_n1644_n3288# 0.184696f
C737 plus.n30 a_n1644_n3288# 0.020613f
C738 plus.n31 a_n1644_n3288# 0.184696f
C739 plus.n32 a_n1644_n3288# 0.200069f
C740 plus.n33 a_n1644_n3288# 1.5491f
.ends

