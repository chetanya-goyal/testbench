* NGSPICE file created from diffpair147.ext - technology: sky130A

.subckt diffpair147 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t9 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X1 a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X2 source.t30 plus.t1 drain_left.t0 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 source.t1 minus.t0 drain_right.t15 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X4 source.t7 minus.t1 drain_right.t14 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X5 drain_right.t13 minus.t2 source.t11 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X6 drain_left.t2 plus.t2 source.t29 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X7 source.t28 plus.t3 drain_left.t6 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X8 source.t27 plus.t4 drain_left.t12 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X9 a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X10 a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X11 drain_right.t12 minus.t3 source.t5 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X12 drain_left.t13 plus.t5 source.t26 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 source.t25 plus.t6 drain_left.t4 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X14 drain_right.t11 minus.t4 source.t6 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X15 drain_right.t10 minus.t5 source.t12 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X16 drain_left.t15 plus.t7 source.t24 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X17 drain_right.t9 minus.t6 source.t4 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X18 drain_left.t10 plus.t8 source.t23 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_left.t5 plus.t9 source.t22 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X20 source.t21 plus.t10 drain_left.t7 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X21 drain_left.t14 plus.t11 source.t20 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X22 drain_right.t8 minus.t7 source.t9 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 drain_right.t7 minus.t8 source.t13 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X24 source.t0 minus.t9 drain_right.t6 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X25 drain_left.t11 plus.t12 source.t19 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X26 source.t18 plus.t13 drain_left.t8 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X27 drain_right.t5 minus.t10 source.t2 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X28 source.t3 minus.t11 drain_right.t4 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X29 a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X30 source.t8 minus.t12 drain_right.t3 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X31 source.t15 minus.t13 drain_right.t2 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X32 source.t17 plus.t14 drain_left.t3 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X33 drain_left.t1 plus.t15 source.t16 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X34 source.t14 minus.t14 drain_right.t1 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X35 source.t10 minus.t15 drain_right.t0 a_n2570_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
R0 plus.n9 plus.n8 161.3
R1 plus.n10 plus.n5 161.3
R2 plus.n12 plus.n11 161.3
R3 plus.n13 plus.n4 161.3
R4 plus.n15 plus.n14 161.3
R5 plus.n16 plus.n3 161.3
R6 plus.n18 plus.n17 161.3
R7 plus.n19 plus.n2 161.3
R8 plus.n21 plus.n20 161.3
R9 plus.n22 plus.n1 161.3
R10 plus.n23 plus.n0 161.3
R11 plus.n25 plus.n24 161.3
R12 plus.n35 plus.n34 161.3
R13 plus.n36 plus.n31 161.3
R14 plus.n38 plus.n37 161.3
R15 plus.n39 plus.n30 161.3
R16 plus.n41 plus.n40 161.3
R17 plus.n42 plus.n29 161.3
R18 plus.n44 plus.n43 161.3
R19 plus.n45 plus.n28 161.3
R20 plus.n47 plus.n46 161.3
R21 plus.n48 plus.n27 161.3
R22 plus.n49 plus.n26 161.3
R23 plus.n51 plus.n50 161.3
R24 plus.n7 plus.t4 149.351
R25 plus.n33 plus.t15 149.351
R26 plus.n24 plus.t7 124.977
R27 plus.n22 plus.t0 124.977
R28 plus.n2 plus.t11 124.977
R29 plus.n16 plus.t3 124.977
R30 plus.n4 plus.t9 124.977
R31 plus.n10 plus.t1 124.977
R32 plus.n6 plus.t12 124.977
R33 plus.n50 plus.t13 124.977
R34 plus.n48 plus.t8 124.977
R35 plus.n28 plus.t10 124.977
R36 plus.n42 plus.t5 124.977
R37 plus.n30 plus.t6 124.977
R38 plus.n36 plus.t2 124.977
R39 plus.n32 plus.t14 124.977
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus.n22 plus.n21 32.8641
R45 plus.n9 plus.n6 32.8641
R46 plus.n48 plus.n47 32.8641
R47 plus.n35 plus.n32 32.8641
R48 plus plus.n51 29.1051
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus.n23 plus.n22 10.955
R68 plus.n49 plus.n48 10.955
R69 plus plus.n25 8.51186
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 drain_left.n9 drain_left.n7 101.683
R93 drain_left.n5 drain_left.n3 101.683
R94 drain_left.n2 drain_left.n0 101.683
R95 drain_left.n13 drain_left.n12 100.796
R96 drain_left.n11 drain_left.n10 100.796
R97 drain_left.n9 drain_left.n8 100.796
R98 drain_left.n5 drain_left.n4 100.796
R99 drain_left.n2 drain_left.n1 100.796
R100 drain_left drain_left.n6 25.5629
R101 drain_left.n3 drain_left.t3 9.9005
R102 drain_left.n3 drain_left.t1 9.9005
R103 drain_left.n4 drain_left.t4 9.9005
R104 drain_left.n4 drain_left.t2 9.9005
R105 drain_left.n1 drain_left.t7 9.9005
R106 drain_left.n1 drain_left.t13 9.9005
R107 drain_left.n0 drain_left.t8 9.9005
R108 drain_left.n0 drain_left.t10 9.9005
R109 drain_left.n12 drain_left.t9 9.9005
R110 drain_left.n12 drain_left.t15 9.9005
R111 drain_left.n10 drain_left.t6 9.9005
R112 drain_left.n10 drain_left.t14 9.9005
R113 drain_left.n8 drain_left.t0 9.9005
R114 drain_left.n8 drain_left.t5 9.9005
R115 drain_left.n7 drain_left.t12 9.9005
R116 drain_left.n7 drain_left.t11 9.9005
R117 drain_left drain_left.n13 6.54115
R118 drain_left.n11 drain_left.n9 0.888431
R119 drain_left.n13 drain_left.n11 0.888431
R120 drain_left.n6 drain_left.n5 0.389119
R121 drain_left.n6 drain_left.n2 0.389119
R122 source.n82 source.n80 289.615
R123 source.n68 source.n66 289.615
R124 source.n60 source.n58 289.615
R125 source.n46 source.n44 289.615
R126 source.n2 source.n0 289.615
R127 source.n16 source.n14 289.615
R128 source.n24 source.n22 289.615
R129 source.n38 source.n36 289.615
R130 source.n83 source.n82 185
R131 source.n69 source.n68 185
R132 source.n61 source.n60 185
R133 source.n47 source.n46 185
R134 source.n3 source.n2 185
R135 source.n17 source.n16 185
R136 source.n25 source.n24 185
R137 source.n39 source.n38 185
R138 source.t5 source.n81 167.117
R139 source.t0 source.n67 167.117
R140 source.t16 source.n59 167.117
R141 source.t18 source.n45 167.117
R142 source.t24 source.n1 167.117
R143 source.t27 source.n15 167.117
R144 source.t13 source.n23 167.117
R145 source.t3 source.n37 167.117
R146 source.n9 source.n8 84.1169
R147 source.n11 source.n10 84.1169
R148 source.n13 source.n12 84.1169
R149 source.n31 source.n30 84.1169
R150 source.n33 source.n32 84.1169
R151 source.n35 source.n34 84.1169
R152 source.n79 source.n78 84.1168
R153 source.n77 source.n76 84.1168
R154 source.n75 source.n74 84.1168
R155 source.n57 source.n56 84.1168
R156 source.n55 source.n54 84.1168
R157 source.n53 source.n52 84.1168
R158 source.n82 source.t5 52.3082
R159 source.n68 source.t0 52.3082
R160 source.n60 source.t16 52.3082
R161 source.n46 source.t18 52.3082
R162 source.n2 source.t24 52.3082
R163 source.n16 source.t27 52.3082
R164 source.n24 source.t13 52.3082
R165 source.n38 source.t3 52.3082
R166 source.n87 source.n86 31.4096
R167 source.n73 source.n72 31.4096
R168 source.n65 source.n64 31.4096
R169 source.n51 source.n50 31.4096
R170 source.n7 source.n6 31.4096
R171 source.n21 source.n20 31.4096
R172 source.n29 source.n28 31.4096
R173 source.n43 source.n42 31.4096
R174 source.n51 source.n43 14.5999
R175 source.n78 source.t11 9.9005
R176 source.n78 source.t7 9.9005
R177 source.n76 source.t2 9.9005
R178 source.n76 source.t15 9.9005
R179 source.n74 source.t9 9.9005
R180 source.n74 source.t8 9.9005
R181 source.n56 source.t29 9.9005
R182 source.n56 source.t17 9.9005
R183 source.n54 source.t26 9.9005
R184 source.n54 source.t25 9.9005
R185 source.n52 source.t23 9.9005
R186 source.n52 source.t21 9.9005
R187 source.n8 source.t20 9.9005
R188 source.n8 source.t31 9.9005
R189 source.n10 source.t22 9.9005
R190 source.n10 source.t28 9.9005
R191 source.n12 source.t19 9.9005
R192 source.n12 source.t30 9.9005
R193 source.n30 source.t4 9.9005
R194 source.n30 source.t1 9.9005
R195 source.n32 source.t12 9.9005
R196 source.n32 source.t14 9.9005
R197 source.n34 source.t6 9.9005
R198 source.n34 source.t10 9.9005
R199 source.n83 source.n81 9.71174
R200 source.n69 source.n67 9.71174
R201 source.n61 source.n59 9.71174
R202 source.n47 source.n45 9.71174
R203 source.n3 source.n1 9.71174
R204 source.n17 source.n15 9.71174
R205 source.n25 source.n23 9.71174
R206 source.n39 source.n37 9.71174
R207 source.n86 source.n85 9.45567
R208 source.n72 source.n71 9.45567
R209 source.n64 source.n63 9.45567
R210 source.n50 source.n49 9.45567
R211 source.n6 source.n5 9.45567
R212 source.n20 source.n19 9.45567
R213 source.n28 source.n27 9.45567
R214 source.n42 source.n41 9.45567
R215 source.n85 source.n84 9.3005
R216 source.n71 source.n70 9.3005
R217 source.n63 source.n62 9.3005
R218 source.n49 source.n48 9.3005
R219 source.n5 source.n4 9.3005
R220 source.n19 source.n18 9.3005
R221 source.n27 source.n26 9.3005
R222 source.n41 source.n40 9.3005
R223 source.n88 source.n7 8.893
R224 source.n86 source.n80 8.14595
R225 source.n72 source.n66 8.14595
R226 source.n64 source.n58 8.14595
R227 source.n50 source.n44 8.14595
R228 source.n6 source.n0 8.14595
R229 source.n20 source.n14 8.14595
R230 source.n28 source.n22 8.14595
R231 source.n42 source.n36 8.14595
R232 source.n84 source.n83 7.3702
R233 source.n70 source.n69 7.3702
R234 source.n62 source.n61 7.3702
R235 source.n48 source.n47 7.3702
R236 source.n4 source.n3 7.3702
R237 source.n18 source.n17 7.3702
R238 source.n26 source.n25 7.3702
R239 source.n40 source.n39 7.3702
R240 source.n84 source.n80 5.81868
R241 source.n70 source.n66 5.81868
R242 source.n62 source.n58 5.81868
R243 source.n48 source.n44 5.81868
R244 source.n4 source.n0 5.81868
R245 source.n18 source.n14 5.81868
R246 source.n26 source.n22 5.81868
R247 source.n40 source.n36 5.81868
R248 source.n88 source.n87 5.7074
R249 source.n85 source.n81 3.44771
R250 source.n71 source.n67 3.44771
R251 source.n63 source.n59 3.44771
R252 source.n49 source.n45 3.44771
R253 source.n5 source.n1 3.44771
R254 source.n19 source.n15 3.44771
R255 source.n27 source.n23 3.44771
R256 source.n41 source.n37 3.44771
R257 source.n43 source.n35 0.888431
R258 source.n35 source.n33 0.888431
R259 source.n33 source.n31 0.888431
R260 source.n31 source.n29 0.888431
R261 source.n21 source.n13 0.888431
R262 source.n13 source.n11 0.888431
R263 source.n11 source.n9 0.888431
R264 source.n9 source.n7 0.888431
R265 source.n53 source.n51 0.888431
R266 source.n55 source.n53 0.888431
R267 source.n57 source.n55 0.888431
R268 source.n65 source.n57 0.888431
R269 source.n75 source.n73 0.888431
R270 source.n77 source.n75 0.888431
R271 source.n79 source.n77 0.888431
R272 source.n87 source.n79 0.888431
R273 source.n29 source.n21 0.470328
R274 source.n73 source.n65 0.470328
R275 source source.n88 0.188
R276 minus.n25 minus.n24 161.3
R277 minus.n23 minus.n0 161.3
R278 minus.n22 minus.n21 161.3
R279 minus.n20 minus.n1 161.3
R280 minus.n19 minus.n18 161.3
R281 minus.n17 minus.n2 161.3
R282 minus.n16 minus.n15 161.3
R283 minus.n14 minus.n3 161.3
R284 minus.n13 minus.n12 161.3
R285 minus.n11 minus.n4 161.3
R286 minus.n10 minus.n9 161.3
R287 minus.n8 minus.n5 161.3
R288 minus.n51 minus.n50 161.3
R289 minus.n49 minus.n26 161.3
R290 minus.n48 minus.n47 161.3
R291 minus.n46 minus.n27 161.3
R292 minus.n45 minus.n44 161.3
R293 minus.n43 minus.n28 161.3
R294 minus.n42 minus.n41 161.3
R295 minus.n40 minus.n29 161.3
R296 minus.n39 minus.n38 161.3
R297 minus.n37 minus.n30 161.3
R298 minus.n36 minus.n35 161.3
R299 minus.n34 minus.n31 161.3
R300 minus.n7 minus.t8 149.351
R301 minus.n33 minus.t9 149.351
R302 minus.n6 minus.t0 124.977
R303 minus.n10 minus.t6 124.977
R304 minus.n12 minus.t14 124.977
R305 minus.n16 minus.t5 124.977
R306 minus.n18 minus.t15 124.977
R307 minus.n22 minus.t4 124.977
R308 minus.n24 minus.t11 124.977
R309 minus.n32 minus.t7 124.977
R310 minus.n36 minus.t12 124.977
R311 minus.n38 minus.t10 124.977
R312 minus.n42 minus.t13 124.977
R313 minus.n44 minus.t2 124.977
R314 minus.n48 minus.t1 124.977
R315 minus.n50 minus.t3 124.977
R316 minus.n8 minus.n7 44.9377
R317 minus.n34 minus.n33 44.9377
R318 minus.n24 minus.n23 37.246
R319 minus.n50 minus.n49 37.246
R320 minus.n6 minus.n5 32.8641
R321 minus.n22 minus.n1 32.8641
R322 minus.n32 minus.n31 32.8641
R323 minus.n48 minus.n27 32.8641
R324 minus.n52 minus.n25 31.4361
R325 minus.n11 minus.n10 28.4823
R326 minus.n18 minus.n17 28.4823
R327 minus.n37 minus.n36 28.4823
R328 minus.n44 minus.n43 28.4823
R329 minus.n16 minus.n3 24.1005
R330 minus.n12 minus.n3 24.1005
R331 minus.n38 minus.n29 24.1005
R332 minus.n42 minus.n29 24.1005
R333 minus.n12 minus.n11 19.7187
R334 minus.n17 minus.n16 19.7187
R335 minus.n38 minus.n37 19.7187
R336 minus.n43 minus.n42 19.7187
R337 minus.n7 minus.n6 17.0522
R338 minus.n33 minus.n32 17.0522
R339 minus.n10 minus.n5 15.3369
R340 minus.n18 minus.n1 15.3369
R341 minus.n36 minus.n31 15.3369
R342 minus.n44 minus.n27 15.3369
R343 minus.n23 minus.n22 10.955
R344 minus.n49 minus.n48 10.955
R345 minus.n52 minus.n51 6.6558
R346 minus.n25 minus.n0 0.189894
R347 minus.n21 minus.n0 0.189894
R348 minus.n21 minus.n20 0.189894
R349 minus.n20 minus.n19 0.189894
R350 minus.n19 minus.n2 0.189894
R351 minus.n15 minus.n2 0.189894
R352 minus.n15 minus.n14 0.189894
R353 minus.n14 minus.n13 0.189894
R354 minus.n13 minus.n4 0.189894
R355 minus.n9 minus.n4 0.189894
R356 minus.n9 minus.n8 0.189894
R357 minus.n35 minus.n34 0.189894
R358 minus.n35 minus.n30 0.189894
R359 minus.n39 minus.n30 0.189894
R360 minus.n40 minus.n39 0.189894
R361 minus.n41 minus.n40 0.189894
R362 minus.n41 minus.n28 0.189894
R363 minus.n45 minus.n28 0.189894
R364 minus.n46 minus.n45 0.189894
R365 minus.n47 minus.n46 0.189894
R366 minus.n47 minus.n26 0.189894
R367 minus.n51 minus.n26 0.189894
R368 minus minus.n52 0.188
R369 drain_right.n9 drain_right.n7 101.683
R370 drain_right.n5 drain_right.n3 101.683
R371 drain_right.n2 drain_right.n0 101.683
R372 drain_right.n9 drain_right.n8 100.796
R373 drain_right.n11 drain_right.n10 100.796
R374 drain_right.n13 drain_right.n12 100.796
R375 drain_right.n5 drain_right.n4 100.796
R376 drain_right.n2 drain_right.n1 100.796
R377 drain_right drain_right.n6 25.0096
R378 drain_right.n3 drain_right.t14 9.9005
R379 drain_right.n3 drain_right.t12 9.9005
R380 drain_right.n4 drain_right.t2 9.9005
R381 drain_right.n4 drain_right.t13 9.9005
R382 drain_right.n1 drain_right.t3 9.9005
R383 drain_right.n1 drain_right.t5 9.9005
R384 drain_right.n0 drain_right.t6 9.9005
R385 drain_right.n0 drain_right.t8 9.9005
R386 drain_right.n7 drain_right.t15 9.9005
R387 drain_right.n7 drain_right.t7 9.9005
R388 drain_right.n8 drain_right.t1 9.9005
R389 drain_right.n8 drain_right.t9 9.9005
R390 drain_right.n10 drain_right.t0 9.9005
R391 drain_right.n10 drain_right.t10 9.9005
R392 drain_right.n12 drain_right.t4 9.9005
R393 drain_right.n12 drain_right.t11 9.9005
R394 drain_right drain_right.n13 6.54115
R395 drain_right.n13 drain_right.n11 0.888431
R396 drain_right.n11 drain_right.n9 0.888431
R397 drain_right.n6 drain_right.n5 0.389119
R398 drain_right.n6 drain_right.n2 0.389119
C0 source drain_right 6.18729f
C1 drain_right minus 2.20322f
C2 plus drain_left 2.45776f
C3 source plus 2.79658f
C4 plus minus 4.5062f
C5 plus drain_right 0.417525f
C6 source drain_left 6.18505f
C7 minus drain_left 0.178616f
C8 source minus 2.78262f
C9 drain_right drain_left 1.34352f
C10 drain_right a_n2570_n1288# 4.81776f
C11 drain_left a_n2570_n1288# 5.21034f
C12 source a_n2570_n1288# 3.363547f
C13 minus a_n2570_n1288# 9.425623f
C14 plus a_n2570_n1288# 10.73105f
C15 drain_right.t6 a_n2570_n1288# 0.042088f
C16 drain_right.t8 a_n2570_n1288# 0.042088f
C17 drain_right.n0 a_n2570_n1288# 0.267613f
C18 drain_right.t3 a_n2570_n1288# 0.042088f
C19 drain_right.t5 a_n2570_n1288# 0.042088f
C20 drain_right.n1 a_n2570_n1288# 0.264408f
C21 drain_right.n2 a_n2570_n1288# 0.67868f
C22 drain_right.t14 a_n2570_n1288# 0.042088f
C23 drain_right.t12 a_n2570_n1288# 0.042088f
C24 drain_right.n3 a_n2570_n1288# 0.267613f
C25 drain_right.t2 a_n2570_n1288# 0.042088f
C26 drain_right.t13 a_n2570_n1288# 0.042088f
C27 drain_right.n4 a_n2570_n1288# 0.264408f
C28 drain_right.n5 a_n2570_n1288# 0.67868f
C29 drain_right.n6 a_n2570_n1288# 0.923615f
C30 drain_right.t15 a_n2570_n1288# 0.042088f
C31 drain_right.t7 a_n2570_n1288# 0.042088f
C32 drain_right.n7 a_n2570_n1288# 0.267614f
C33 drain_right.t1 a_n2570_n1288# 0.042088f
C34 drain_right.t9 a_n2570_n1288# 0.042088f
C35 drain_right.n8 a_n2570_n1288# 0.264409f
C36 drain_right.n9 a_n2570_n1288# 0.719934f
C37 drain_right.t0 a_n2570_n1288# 0.042088f
C38 drain_right.t10 a_n2570_n1288# 0.042088f
C39 drain_right.n10 a_n2570_n1288# 0.264409f
C40 drain_right.n11 a_n2570_n1288# 0.356206f
C41 drain_right.t4 a_n2570_n1288# 0.042088f
C42 drain_right.t11 a_n2570_n1288# 0.042088f
C43 drain_right.n12 a_n2570_n1288# 0.264409f
C44 drain_right.n13 a_n2570_n1288# 0.591751f
C45 minus.n0 a_n2570_n1288# 0.043252f
C46 minus.n1 a_n2570_n1288# 0.009815f
C47 minus.t4 a_n2570_n1288# 0.187517f
C48 minus.n2 a_n2570_n1288# 0.043252f
C49 minus.n3 a_n2570_n1288# 0.009815f
C50 minus.t5 a_n2570_n1288# 0.187517f
C51 minus.n4 a_n2570_n1288# 0.043252f
C52 minus.n5 a_n2570_n1288# 0.009815f
C53 minus.t6 a_n2570_n1288# 0.187517f
C54 minus.t8 a_n2570_n1288# 0.208818f
C55 minus.t0 a_n2570_n1288# 0.187517f
C56 minus.n6 a_n2570_n1288# 0.136274f
C57 minus.n7 a_n2570_n1288# 0.112647f
C58 minus.n8 a_n2570_n1288# 0.183033f
C59 minus.n9 a_n2570_n1288# 0.043252f
C60 minus.n10 a_n2570_n1288# 0.130349f
C61 minus.n11 a_n2570_n1288# 0.009815f
C62 minus.t14 a_n2570_n1288# 0.187517f
C63 minus.n12 a_n2570_n1288# 0.130349f
C64 minus.n13 a_n2570_n1288# 0.043252f
C65 minus.n14 a_n2570_n1288# 0.043252f
C66 minus.n15 a_n2570_n1288# 0.043252f
C67 minus.n16 a_n2570_n1288# 0.130349f
C68 minus.n17 a_n2570_n1288# 0.009815f
C69 minus.t15 a_n2570_n1288# 0.187517f
C70 minus.n18 a_n2570_n1288# 0.130349f
C71 minus.n19 a_n2570_n1288# 0.043252f
C72 minus.n20 a_n2570_n1288# 0.043252f
C73 minus.n21 a_n2570_n1288# 0.043252f
C74 minus.n22 a_n2570_n1288# 0.130349f
C75 minus.n23 a_n2570_n1288# 0.009815f
C76 minus.t11 a_n2570_n1288# 0.187517f
C77 minus.n24 a_n2570_n1288# 0.129149f
C78 minus.n25 a_n2570_n1288# 1.22355f
C79 minus.n26 a_n2570_n1288# 0.043252f
C80 minus.n27 a_n2570_n1288# 0.009815f
C81 minus.n28 a_n2570_n1288# 0.043252f
C82 minus.n29 a_n2570_n1288# 0.009815f
C83 minus.n30 a_n2570_n1288# 0.043252f
C84 minus.n31 a_n2570_n1288# 0.009815f
C85 minus.t9 a_n2570_n1288# 0.208818f
C86 minus.t7 a_n2570_n1288# 0.187517f
C87 minus.n32 a_n2570_n1288# 0.136274f
C88 minus.n33 a_n2570_n1288# 0.112647f
C89 minus.n34 a_n2570_n1288# 0.183033f
C90 minus.n35 a_n2570_n1288# 0.043252f
C91 minus.t12 a_n2570_n1288# 0.187517f
C92 minus.n36 a_n2570_n1288# 0.130349f
C93 minus.n37 a_n2570_n1288# 0.009815f
C94 minus.t10 a_n2570_n1288# 0.187517f
C95 minus.n38 a_n2570_n1288# 0.130349f
C96 minus.n39 a_n2570_n1288# 0.043252f
C97 minus.n40 a_n2570_n1288# 0.043252f
C98 minus.n41 a_n2570_n1288# 0.043252f
C99 minus.t13 a_n2570_n1288# 0.187517f
C100 minus.n42 a_n2570_n1288# 0.130349f
C101 minus.n43 a_n2570_n1288# 0.009815f
C102 minus.t2 a_n2570_n1288# 0.187517f
C103 minus.n44 a_n2570_n1288# 0.130349f
C104 minus.n45 a_n2570_n1288# 0.043252f
C105 minus.n46 a_n2570_n1288# 0.043252f
C106 minus.n47 a_n2570_n1288# 0.043252f
C107 minus.t1 a_n2570_n1288# 0.187517f
C108 minus.n48 a_n2570_n1288# 0.130349f
C109 minus.n49 a_n2570_n1288# 0.009815f
C110 minus.t3 a_n2570_n1288# 0.187517f
C111 minus.n50 a_n2570_n1288# 0.129149f
C112 minus.n51 a_n2570_n1288# 0.298534f
C113 minus.n52 a_n2570_n1288# 1.49811f
C114 source.n0 a_n2570_n1288# 0.044625f
C115 source.n1 a_n2570_n1288# 0.098739f
C116 source.t24 a_n2570_n1288# 0.074098f
C117 source.n2 a_n2570_n1288# 0.077277f
C118 source.n3 a_n2570_n1288# 0.024911f
C119 source.n4 a_n2570_n1288# 0.016429f
C120 source.n5 a_n2570_n1288# 0.217644f
C121 source.n6 a_n2570_n1288# 0.048919f
C122 source.n7 a_n2570_n1288# 0.521811f
C123 source.t20 a_n2570_n1288# 0.048321f
C124 source.t31 a_n2570_n1288# 0.048321f
C125 source.n8 a_n2570_n1288# 0.258325f
C126 source.n9 a_n2570_n1288# 0.412654f
C127 source.t22 a_n2570_n1288# 0.048321f
C128 source.t28 a_n2570_n1288# 0.048321f
C129 source.n10 a_n2570_n1288# 0.258325f
C130 source.n11 a_n2570_n1288# 0.412654f
C131 source.t19 a_n2570_n1288# 0.048321f
C132 source.t30 a_n2570_n1288# 0.048321f
C133 source.n12 a_n2570_n1288# 0.258325f
C134 source.n13 a_n2570_n1288# 0.412654f
C135 source.n14 a_n2570_n1288# 0.044625f
C136 source.n15 a_n2570_n1288# 0.098739f
C137 source.t27 a_n2570_n1288# 0.074098f
C138 source.n16 a_n2570_n1288# 0.077277f
C139 source.n17 a_n2570_n1288# 0.024911f
C140 source.n18 a_n2570_n1288# 0.016429f
C141 source.n19 a_n2570_n1288# 0.217644f
C142 source.n20 a_n2570_n1288# 0.048919f
C143 source.n21 a_n2570_n1288# 0.158933f
C144 source.n22 a_n2570_n1288# 0.044625f
C145 source.n23 a_n2570_n1288# 0.098739f
C146 source.t13 a_n2570_n1288# 0.074098f
C147 source.n24 a_n2570_n1288# 0.077277f
C148 source.n25 a_n2570_n1288# 0.024911f
C149 source.n26 a_n2570_n1288# 0.016429f
C150 source.n27 a_n2570_n1288# 0.217644f
C151 source.n28 a_n2570_n1288# 0.048919f
C152 source.n29 a_n2570_n1288# 0.158933f
C153 source.t4 a_n2570_n1288# 0.048321f
C154 source.t1 a_n2570_n1288# 0.048321f
C155 source.n30 a_n2570_n1288# 0.258325f
C156 source.n31 a_n2570_n1288# 0.412654f
C157 source.t12 a_n2570_n1288# 0.048321f
C158 source.t14 a_n2570_n1288# 0.048321f
C159 source.n32 a_n2570_n1288# 0.258325f
C160 source.n33 a_n2570_n1288# 0.412654f
C161 source.t6 a_n2570_n1288# 0.048321f
C162 source.t10 a_n2570_n1288# 0.048321f
C163 source.n34 a_n2570_n1288# 0.258325f
C164 source.n35 a_n2570_n1288# 0.412654f
C165 source.n36 a_n2570_n1288# 0.044625f
C166 source.n37 a_n2570_n1288# 0.098739f
C167 source.t3 a_n2570_n1288# 0.074098f
C168 source.n38 a_n2570_n1288# 0.077277f
C169 source.n39 a_n2570_n1288# 0.024911f
C170 source.n40 a_n2570_n1288# 0.016429f
C171 source.n41 a_n2570_n1288# 0.217644f
C172 source.n42 a_n2570_n1288# 0.048919f
C173 source.n43 a_n2570_n1288# 0.814611f
C174 source.n44 a_n2570_n1288# 0.044625f
C175 source.n45 a_n2570_n1288# 0.098739f
C176 source.t18 a_n2570_n1288# 0.074098f
C177 source.n46 a_n2570_n1288# 0.077277f
C178 source.n47 a_n2570_n1288# 0.024911f
C179 source.n48 a_n2570_n1288# 0.016429f
C180 source.n49 a_n2570_n1288# 0.217644f
C181 source.n50 a_n2570_n1288# 0.048919f
C182 source.n51 a_n2570_n1288# 0.814611f
C183 source.t23 a_n2570_n1288# 0.048321f
C184 source.t21 a_n2570_n1288# 0.048321f
C185 source.n52 a_n2570_n1288# 0.258324f
C186 source.n53 a_n2570_n1288# 0.412656f
C187 source.t26 a_n2570_n1288# 0.048321f
C188 source.t25 a_n2570_n1288# 0.048321f
C189 source.n54 a_n2570_n1288# 0.258324f
C190 source.n55 a_n2570_n1288# 0.412656f
C191 source.t29 a_n2570_n1288# 0.048321f
C192 source.t17 a_n2570_n1288# 0.048321f
C193 source.n56 a_n2570_n1288# 0.258324f
C194 source.n57 a_n2570_n1288# 0.412656f
C195 source.n58 a_n2570_n1288# 0.044625f
C196 source.n59 a_n2570_n1288# 0.098739f
C197 source.t16 a_n2570_n1288# 0.074098f
C198 source.n60 a_n2570_n1288# 0.077277f
C199 source.n61 a_n2570_n1288# 0.024911f
C200 source.n62 a_n2570_n1288# 0.016429f
C201 source.n63 a_n2570_n1288# 0.217644f
C202 source.n64 a_n2570_n1288# 0.048919f
C203 source.n65 a_n2570_n1288# 0.158933f
C204 source.n66 a_n2570_n1288# 0.044625f
C205 source.n67 a_n2570_n1288# 0.098739f
C206 source.t0 a_n2570_n1288# 0.074098f
C207 source.n68 a_n2570_n1288# 0.077277f
C208 source.n69 a_n2570_n1288# 0.024911f
C209 source.n70 a_n2570_n1288# 0.016429f
C210 source.n71 a_n2570_n1288# 0.217644f
C211 source.n72 a_n2570_n1288# 0.048919f
C212 source.n73 a_n2570_n1288# 0.158933f
C213 source.t9 a_n2570_n1288# 0.048321f
C214 source.t8 a_n2570_n1288# 0.048321f
C215 source.n74 a_n2570_n1288# 0.258324f
C216 source.n75 a_n2570_n1288# 0.412656f
C217 source.t2 a_n2570_n1288# 0.048321f
C218 source.t15 a_n2570_n1288# 0.048321f
C219 source.n76 a_n2570_n1288# 0.258324f
C220 source.n77 a_n2570_n1288# 0.412656f
C221 source.t11 a_n2570_n1288# 0.048321f
C222 source.t7 a_n2570_n1288# 0.048321f
C223 source.n78 a_n2570_n1288# 0.258324f
C224 source.n79 a_n2570_n1288# 0.412656f
C225 source.n80 a_n2570_n1288# 0.044625f
C226 source.n81 a_n2570_n1288# 0.098739f
C227 source.t5 a_n2570_n1288# 0.074098f
C228 source.n82 a_n2570_n1288# 0.077277f
C229 source.n83 a_n2570_n1288# 0.024911f
C230 source.n84 a_n2570_n1288# 0.016429f
C231 source.n85 a_n2570_n1288# 0.217644f
C232 source.n86 a_n2570_n1288# 0.048919f
C233 source.n87 a_n2570_n1288# 0.35837f
C234 source.n88 a_n2570_n1288# 0.770787f
C235 drain_left.t8 a_n2570_n1288# 0.043057f
C236 drain_left.t10 a_n2570_n1288# 0.043057f
C237 drain_left.n0 a_n2570_n1288# 0.273775f
C238 drain_left.t7 a_n2570_n1288# 0.043057f
C239 drain_left.t13 a_n2570_n1288# 0.043057f
C240 drain_left.n1 a_n2570_n1288# 0.270497f
C241 drain_left.n2 a_n2570_n1288# 0.694308f
C242 drain_left.t3 a_n2570_n1288# 0.043057f
C243 drain_left.t1 a_n2570_n1288# 0.043057f
C244 drain_left.n3 a_n2570_n1288# 0.273775f
C245 drain_left.t4 a_n2570_n1288# 0.043057f
C246 drain_left.t2 a_n2570_n1288# 0.043057f
C247 drain_left.n4 a_n2570_n1288# 0.270497f
C248 drain_left.n5 a_n2570_n1288# 0.694308f
C249 drain_left.n6 a_n2570_n1288# 0.997886f
C250 drain_left.t12 a_n2570_n1288# 0.043057f
C251 drain_left.t11 a_n2570_n1288# 0.043057f
C252 drain_left.n7 a_n2570_n1288# 0.273776f
C253 drain_left.t0 a_n2570_n1288# 0.043057f
C254 drain_left.t5 a_n2570_n1288# 0.043057f
C255 drain_left.n8 a_n2570_n1288# 0.270498f
C256 drain_left.n9 a_n2570_n1288# 0.736512f
C257 drain_left.t6 a_n2570_n1288# 0.043057f
C258 drain_left.t14 a_n2570_n1288# 0.043057f
C259 drain_left.n10 a_n2570_n1288# 0.270498f
C260 drain_left.n11 a_n2570_n1288# 0.364409f
C261 drain_left.t9 a_n2570_n1288# 0.043057f
C262 drain_left.t15 a_n2570_n1288# 0.043057f
C263 drain_left.n12 a_n2570_n1288# 0.270498f
C264 drain_left.n13 a_n2570_n1288# 0.605377f
C265 plus.n0 a_n2570_n1288# 0.045033f
C266 plus.t7 a_n2570_n1288# 0.195236f
C267 plus.t0 a_n2570_n1288# 0.195236f
C268 plus.n1 a_n2570_n1288# 0.045033f
C269 plus.t11 a_n2570_n1288# 0.195236f
C270 plus.n2 a_n2570_n1288# 0.135715f
C271 plus.n3 a_n2570_n1288# 0.045033f
C272 plus.t3 a_n2570_n1288# 0.195236f
C273 plus.t9 a_n2570_n1288# 0.195236f
C274 plus.n4 a_n2570_n1288# 0.135715f
C275 plus.n5 a_n2570_n1288# 0.045033f
C276 plus.t1 a_n2570_n1288# 0.195236f
C277 plus.t12 a_n2570_n1288# 0.195236f
C278 plus.n6 a_n2570_n1288# 0.141884f
C279 plus.t4 a_n2570_n1288# 0.217414f
C280 plus.n7 a_n2570_n1288# 0.117284f
C281 plus.n8 a_n2570_n1288# 0.190568f
C282 plus.n9 a_n2570_n1288# 0.010219f
C283 plus.n10 a_n2570_n1288# 0.135715f
C284 plus.n11 a_n2570_n1288# 0.010219f
C285 plus.n12 a_n2570_n1288# 0.045033f
C286 plus.n13 a_n2570_n1288# 0.045033f
C287 plus.n14 a_n2570_n1288# 0.045033f
C288 plus.n15 a_n2570_n1288# 0.010219f
C289 plus.n16 a_n2570_n1288# 0.135715f
C290 plus.n17 a_n2570_n1288# 0.010219f
C291 plus.n18 a_n2570_n1288# 0.045033f
C292 plus.n19 a_n2570_n1288# 0.045033f
C293 plus.n20 a_n2570_n1288# 0.045033f
C294 plus.n21 a_n2570_n1288# 0.010219f
C295 plus.n22 a_n2570_n1288# 0.135715f
C296 plus.n23 a_n2570_n1288# 0.010219f
C297 plus.n24 a_n2570_n1288# 0.134466f
C298 plus.n25 a_n2570_n1288# 0.339244f
C299 plus.n26 a_n2570_n1288# 0.045033f
C300 plus.t13 a_n2570_n1288# 0.195236f
C301 plus.n27 a_n2570_n1288# 0.045033f
C302 plus.t8 a_n2570_n1288# 0.195236f
C303 plus.t10 a_n2570_n1288# 0.195236f
C304 plus.n28 a_n2570_n1288# 0.135715f
C305 plus.n29 a_n2570_n1288# 0.045033f
C306 plus.t5 a_n2570_n1288# 0.195236f
C307 plus.t6 a_n2570_n1288# 0.195236f
C308 plus.n30 a_n2570_n1288# 0.135715f
C309 plus.n31 a_n2570_n1288# 0.045033f
C310 plus.t2 a_n2570_n1288# 0.195236f
C311 plus.t14 a_n2570_n1288# 0.195236f
C312 plus.n32 a_n2570_n1288# 0.141884f
C313 plus.t15 a_n2570_n1288# 0.217414f
C314 plus.n33 a_n2570_n1288# 0.117284f
C315 plus.n34 a_n2570_n1288# 0.190568f
C316 plus.n35 a_n2570_n1288# 0.010219f
C317 plus.n36 a_n2570_n1288# 0.135715f
C318 plus.n37 a_n2570_n1288# 0.010219f
C319 plus.n38 a_n2570_n1288# 0.045033f
C320 plus.n39 a_n2570_n1288# 0.045033f
C321 plus.n40 a_n2570_n1288# 0.045033f
C322 plus.n41 a_n2570_n1288# 0.010219f
C323 plus.n42 a_n2570_n1288# 0.135715f
C324 plus.n43 a_n2570_n1288# 0.010219f
C325 plus.n44 a_n2570_n1288# 0.045033f
C326 plus.n45 a_n2570_n1288# 0.045033f
C327 plus.n46 a_n2570_n1288# 0.045033f
C328 plus.n47 a_n2570_n1288# 0.010219f
C329 plus.n48 a_n2570_n1288# 0.135715f
C330 plus.n49 a_n2570_n1288# 0.010219f
C331 plus.n50 a_n2570_n1288# 0.134466f
C332 plus.n51 a_n2570_n1288# 1.21206f
.ends

