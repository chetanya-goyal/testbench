* NGSPICE file created from diffpair208.ext - technology: sky130A

.subckt diffpair208 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t37 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X1 drain_right.t18 minus.t1 source.t33 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X2 source.t6 plus.t0 drain_left.t19 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X3 source.t25 minus.t2 drain_right.t17 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X4 a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X5 source.t32 minus.t3 drain_right.t16 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X6 source.t8 plus.t1 drain_left.t18 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X7 drain_left.t17 plus.t2 source.t39 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X8 source.t38 plus.t3 drain_left.t16 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X9 source.t35 minus.t4 drain_right.t15 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X10 source.t36 minus.t5 drain_right.t14 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X11 drain_right.t13 minus.t6 source.t23 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X12 drain_right.t12 minus.t7 source.t27 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X13 drain_left.t15 plus.t4 source.t9 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X14 drain_right.t11 minus.t8 source.t28 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X15 a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X16 drain_left.t14 plus.t5 source.t7 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X17 drain_right.t10 minus.t9 source.t24 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X18 drain_right.t9 minus.t10 source.t20 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X19 source.t11 plus.t6 drain_left.t13 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X20 source.t14 plus.t7 drain_left.t12 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X21 source.t22 minus.t11 drain_right.t8 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X22 source.t18 minus.t12 drain_right.t7 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X23 source.t0 plus.t8 drain_left.t11 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X24 source.t19 minus.t13 drain_right.t6 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X25 source.t21 minus.t14 drain_right.t5 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X26 source.t16 plus.t9 drain_left.t10 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X27 drain_left.t9 plus.t10 source.t2 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X28 drain_left.t8 plus.t11 source.t10 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X29 drain_right.t4 minus.t15 source.t34 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X30 drain_left.t7 plus.t12 source.t13 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X31 drain_right.t3 minus.t16 source.t30 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X32 source.t31 minus.t17 drain_right.t2 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X33 drain_left.t6 plus.t13 source.t4 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X34 source.t29 minus.t18 drain_right.t1 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X35 drain_left.t5 plus.t14 source.t17 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X36 source.t5 plus.t15 drain_left.t4 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X37 a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X38 drain_left.t3 plus.t16 source.t12 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X39 source.t15 plus.t17 drain_left.t2 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X40 a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X41 drain_right.t0 minus.t19 source.t26 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X42 source.t3 plus.t18 drain_left.t1 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X43 drain_left.t0 plus.t19 source.t1 a_n2542_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
R0 minus.n6 minus.t15 244.149
R1 minus.n34 minus.t5 244.149
R2 minus.n7 minus.t3 223.167
R3 minus.n5 minus.t8 223.167
R4 minus.n13 minus.t18 223.167
R5 minus.n14 minus.t6 223.167
R6 minus.n18 minus.t11 223.167
R7 minus.n19 minus.t0 223.167
R8 minus.n1 minus.t13 223.167
R9 minus.n25 minus.t16 223.167
R10 minus.n26 minus.t4 223.167
R11 minus.n35 minus.t9 223.167
R12 minus.n33 minus.t2 223.167
R13 minus.n41 minus.t7 223.167
R14 minus.n42 minus.t17 223.167
R15 minus.n46 minus.t10 223.167
R16 minus.n47 minus.t14 223.167
R17 minus.n29 minus.t1 223.167
R18 minus.n53 minus.t12 223.167
R19 minus.n54 minus.t19 223.167
R20 minus.n27 minus.n26 161.3
R21 minus.n25 minus.n0 161.3
R22 minus.n24 minus.n23 161.3
R23 minus.n22 minus.n1 161.3
R24 minus.n21 minus.n20 161.3
R25 minus.n19 minus.n2 161.3
R26 minus.n18 minus.n17 161.3
R27 minus.n16 minus.n3 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n4 161.3
R30 minus.n12 minus.n11 161.3
R31 minus.n10 minus.n5 161.3
R32 minus.n9 minus.n8 161.3
R33 minus.n55 minus.n54 161.3
R34 minus.n53 minus.n28 161.3
R35 minus.n52 minus.n51 161.3
R36 minus.n50 minus.n29 161.3
R37 minus.n49 minus.n48 161.3
R38 minus.n47 minus.n30 161.3
R39 minus.n46 minus.n45 161.3
R40 minus.n44 minus.n31 161.3
R41 minus.n43 minus.n42 161.3
R42 minus.n41 minus.n32 161.3
R43 minus.n40 minus.n39 161.3
R44 minus.n38 minus.n33 161.3
R45 minus.n37 minus.n36 161.3
R46 minus.n9 minus.n6 70.4033
R47 minus.n37 minus.n34 70.4033
R48 minus.n14 minus.n13 48.2005
R49 minus.n19 minus.n18 48.2005
R50 minus.n26 minus.n25 48.2005
R51 minus.n42 minus.n41 48.2005
R52 minus.n47 minus.n46 48.2005
R53 minus.n54 minus.n53 48.2005
R54 minus.n12 minus.n5 47.4702
R55 minus.n20 minus.n1 47.4702
R56 minus.n40 minus.n33 47.4702
R57 minus.n48 minus.n29 47.4702
R58 minus.n56 minus.n27 32.0232
R59 minus.n8 minus.n5 25.5611
R60 minus.n24 minus.n1 25.5611
R61 minus.n36 minus.n33 25.5611
R62 minus.n52 minus.n29 25.5611
R63 minus.n18 minus.n3 24.1005
R64 minus.n14 minus.n3 24.1005
R65 minus.n42 minus.n31 24.1005
R66 minus.n46 minus.n31 24.1005
R67 minus.n8 minus.n7 22.6399
R68 minus.n25 minus.n24 22.6399
R69 minus.n36 minus.n35 22.6399
R70 minus.n53 minus.n52 22.6399
R71 minus.n7 minus.n6 20.9576
R72 minus.n35 minus.n34 20.9576
R73 minus.n56 minus.n55 6.59141
R74 minus.n13 minus.n12 0.730803
R75 minus.n20 minus.n19 0.730803
R76 minus.n41 minus.n40 0.730803
R77 minus.n48 minus.n47 0.730803
R78 minus.n27 minus.n0 0.189894
R79 minus.n23 minus.n0 0.189894
R80 minus.n23 minus.n22 0.189894
R81 minus.n22 minus.n21 0.189894
R82 minus.n21 minus.n2 0.189894
R83 minus.n17 minus.n2 0.189894
R84 minus.n17 minus.n16 0.189894
R85 minus.n16 minus.n15 0.189894
R86 minus.n15 minus.n4 0.189894
R87 minus.n11 minus.n4 0.189894
R88 minus.n11 minus.n10 0.189894
R89 minus.n10 minus.n9 0.189894
R90 minus.n38 minus.n37 0.189894
R91 minus.n39 minus.n38 0.189894
R92 minus.n39 minus.n32 0.189894
R93 minus.n43 minus.n32 0.189894
R94 minus.n44 minus.n43 0.189894
R95 minus.n45 minus.n44 0.189894
R96 minus.n45 minus.n30 0.189894
R97 minus.n49 minus.n30 0.189894
R98 minus.n50 minus.n49 0.189894
R99 minus.n51 minus.n50 0.189894
R100 minus.n51 minus.n28 0.189894
R101 minus.n55 minus.n28 0.189894
R102 minus minus.n56 0.188
R103 source.n0 source.t10 69.6943
R104 source.n9 source.t38 69.6943
R105 source.n10 source.t34 69.6943
R106 source.n19 source.t35 69.6943
R107 source.n39 source.t26 69.6942
R108 source.n30 source.t36 69.6942
R109 source.n29 source.t9 69.6942
R110 source.n20 source.t3 69.6942
R111 source.n2 source.n1 63.0943
R112 source.n4 source.n3 63.0943
R113 source.n6 source.n5 63.0943
R114 source.n8 source.n7 63.0943
R115 source.n12 source.n11 63.0943
R116 source.n14 source.n13 63.0943
R117 source.n16 source.n15 63.0943
R118 source.n18 source.n17 63.0943
R119 source.n38 source.n37 63.0942
R120 source.n36 source.n35 63.0942
R121 source.n34 source.n33 63.0942
R122 source.n32 source.n31 63.0942
R123 source.n28 source.n27 63.0942
R124 source.n26 source.n25 63.0942
R125 source.n24 source.n23 63.0942
R126 source.n22 source.n21 63.0942
R127 source.n20 source.n19 15.1851
R128 source.n40 source.n0 9.56437
R129 source.n37 source.t33 6.6005
R130 source.n37 source.t18 6.6005
R131 source.n35 source.t20 6.6005
R132 source.n35 source.t21 6.6005
R133 source.n33 source.t27 6.6005
R134 source.n33 source.t31 6.6005
R135 source.n31 source.t24 6.6005
R136 source.n31 source.t25 6.6005
R137 source.n27 source.t39 6.6005
R138 source.n27 source.t0 6.6005
R139 source.n25 source.t17 6.6005
R140 source.n25 source.t16 6.6005
R141 source.n23 source.t2 6.6005
R142 source.n23 source.t11 6.6005
R143 source.n21 source.t4 6.6005
R144 source.n21 source.t6 6.6005
R145 source.n1 source.t12 6.6005
R146 source.n1 source.t8 6.6005
R147 source.n3 source.t1 6.6005
R148 source.n3 source.t14 6.6005
R149 source.n5 source.t7 6.6005
R150 source.n5 source.t5 6.6005
R151 source.n7 source.t13 6.6005
R152 source.n7 source.t15 6.6005
R153 source.n11 source.t28 6.6005
R154 source.n11 source.t32 6.6005
R155 source.n13 source.t23 6.6005
R156 source.n13 source.t29 6.6005
R157 source.n15 source.t37 6.6005
R158 source.n15 source.t22 6.6005
R159 source.n17 source.t30 6.6005
R160 source.n17 source.t19 6.6005
R161 source.n40 source.n39 5.62119
R162 source.n19 source.n18 0.716017
R163 source.n18 source.n16 0.716017
R164 source.n16 source.n14 0.716017
R165 source.n14 source.n12 0.716017
R166 source.n12 source.n10 0.716017
R167 source.n9 source.n8 0.716017
R168 source.n8 source.n6 0.716017
R169 source.n6 source.n4 0.716017
R170 source.n4 source.n2 0.716017
R171 source.n2 source.n0 0.716017
R172 source.n22 source.n20 0.716017
R173 source.n24 source.n22 0.716017
R174 source.n26 source.n24 0.716017
R175 source.n28 source.n26 0.716017
R176 source.n29 source.n28 0.716017
R177 source.n32 source.n30 0.716017
R178 source.n34 source.n32 0.716017
R179 source.n36 source.n34 0.716017
R180 source.n38 source.n36 0.716017
R181 source.n39 source.n38 0.716017
R182 source.n10 source.n9 0.470328
R183 source.n30 source.n29 0.470328
R184 source source.n40 0.188
R185 drain_right.n10 drain_right.n8 80.4886
R186 drain_right.n6 drain_right.n4 80.4885
R187 drain_right.n2 drain_right.n0 80.4885
R188 drain_right.n10 drain_right.n9 79.7731
R189 drain_right.n12 drain_right.n11 79.7731
R190 drain_right.n14 drain_right.n13 79.7731
R191 drain_right.n16 drain_right.n15 79.7731
R192 drain_right.n7 drain_right.n3 79.773
R193 drain_right.n6 drain_right.n5 79.773
R194 drain_right.n2 drain_right.n1 79.773
R195 drain_right drain_right.n7 25.7198
R196 drain_right.n3 drain_right.t2 6.6005
R197 drain_right.n3 drain_right.t9 6.6005
R198 drain_right.n4 drain_right.t7 6.6005
R199 drain_right.n4 drain_right.t0 6.6005
R200 drain_right.n5 drain_right.t5 6.6005
R201 drain_right.n5 drain_right.t18 6.6005
R202 drain_right.n1 drain_right.t17 6.6005
R203 drain_right.n1 drain_right.t12 6.6005
R204 drain_right.n0 drain_right.t14 6.6005
R205 drain_right.n0 drain_right.t10 6.6005
R206 drain_right.n8 drain_right.t16 6.6005
R207 drain_right.n8 drain_right.t4 6.6005
R208 drain_right.n9 drain_right.t1 6.6005
R209 drain_right.n9 drain_right.t11 6.6005
R210 drain_right.n11 drain_right.t8 6.6005
R211 drain_right.n11 drain_right.t13 6.6005
R212 drain_right.n13 drain_right.t6 6.6005
R213 drain_right.n13 drain_right.t19 6.6005
R214 drain_right.n15 drain_right.t15 6.6005
R215 drain_right.n15 drain_right.t3 6.6005
R216 drain_right drain_right.n16 6.36873
R217 drain_right.n16 drain_right.n14 0.716017
R218 drain_right.n14 drain_right.n12 0.716017
R219 drain_right.n12 drain_right.n10 0.716017
R220 drain_right.n7 drain_right.n6 0.660671
R221 drain_right.n7 drain_right.n2 0.660671
R222 plus.n8 plus.t3 244.149
R223 plus.n36 plus.t4 244.149
R224 plus.n26 plus.t11 223.167
R225 plus.n25 plus.t1 223.167
R226 plus.n1 plus.t16 223.167
R227 plus.n19 plus.t7 223.167
R228 plus.n18 plus.t19 223.167
R229 plus.n4 plus.t15 223.167
R230 plus.n13 plus.t5 223.167
R231 plus.n11 plus.t17 223.167
R232 plus.n7 plus.t12 223.167
R233 plus.n54 plus.t18 223.167
R234 plus.n53 plus.t13 223.167
R235 plus.n29 plus.t0 223.167
R236 plus.n47 plus.t10 223.167
R237 plus.n46 plus.t6 223.167
R238 plus.n32 plus.t14 223.167
R239 plus.n41 plus.t9 223.167
R240 plus.n39 plus.t2 223.167
R241 plus.n35 plus.t8 223.167
R242 plus.n10 plus.n9 161.3
R243 plus.n11 plus.n6 161.3
R244 plus.n12 plus.n5 161.3
R245 plus.n14 plus.n13 161.3
R246 plus.n15 plus.n4 161.3
R247 plus.n17 plus.n16 161.3
R248 plus.n18 plus.n3 161.3
R249 plus.n19 plus.n2 161.3
R250 plus.n21 plus.n20 161.3
R251 plus.n22 plus.n1 161.3
R252 plus.n24 plus.n23 161.3
R253 plus.n25 plus.n0 161.3
R254 plus.n27 plus.n26 161.3
R255 plus.n38 plus.n37 161.3
R256 plus.n39 plus.n34 161.3
R257 plus.n40 plus.n33 161.3
R258 plus.n42 plus.n41 161.3
R259 plus.n43 plus.n32 161.3
R260 plus.n45 plus.n44 161.3
R261 plus.n46 plus.n31 161.3
R262 plus.n47 plus.n30 161.3
R263 plus.n49 plus.n48 161.3
R264 plus.n50 plus.n29 161.3
R265 plus.n52 plus.n51 161.3
R266 plus.n53 plus.n28 161.3
R267 plus.n55 plus.n54 161.3
R268 plus.n9 plus.n8 70.4033
R269 plus.n37 plus.n36 70.4033
R270 plus.n26 plus.n25 48.2005
R271 plus.n19 plus.n18 48.2005
R272 plus.n13 plus.n4 48.2005
R273 plus.n54 plus.n53 48.2005
R274 plus.n47 plus.n46 48.2005
R275 plus.n41 plus.n32 48.2005
R276 plus.n20 plus.n1 47.4702
R277 plus.n12 plus.n11 47.4702
R278 plus.n48 plus.n29 47.4702
R279 plus.n40 plus.n39 47.4702
R280 plus plus.n55 29.3134
R281 plus.n24 plus.n1 25.5611
R282 plus.n11 plus.n10 25.5611
R283 plus.n52 plus.n29 25.5611
R284 plus.n39 plus.n38 25.5611
R285 plus.n17 plus.n4 24.1005
R286 plus.n18 plus.n17 24.1005
R287 plus.n46 plus.n45 24.1005
R288 plus.n45 plus.n32 24.1005
R289 plus.n25 plus.n24 22.6399
R290 plus.n10 plus.n7 22.6399
R291 plus.n53 plus.n52 22.6399
R292 plus.n38 plus.n35 22.6399
R293 plus.n8 plus.n7 20.9576
R294 plus.n36 plus.n35 20.9576
R295 plus plus.n27 8.82626
R296 plus.n20 plus.n19 0.730803
R297 plus.n13 plus.n12 0.730803
R298 plus.n48 plus.n47 0.730803
R299 plus.n41 plus.n40 0.730803
R300 plus.n9 plus.n6 0.189894
R301 plus.n6 plus.n5 0.189894
R302 plus.n14 plus.n5 0.189894
R303 plus.n15 plus.n14 0.189894
R304 plus.n16 plus.n15 0.189894
R305 plus.n16 plus.n3 0.189894
R306 plus.n3 plus.n2 0.189894
R307 plus.n21 plus.n2 0.189894
R308 plus.n22 plus.n21 0.189894
R309 plus.n23 plus.n22 0.189894
R310 plus.n23 plus.n0 0.189894
R311 plus.n27 plus.n0 0.189894
R312 plus.n55 plus.n28 0.189894
R313 plus.n51 plus.n28 0.189894
R314 plus.n51 plus.n50 0.189894
R315 plus.n50 plus.n49 0.189894
R316 plus.n49 plus.n30 0.189894
R317 plus.n31 plus.n30 0.189894
R318 plus.n44 plus.n31 0.189894
R319 plus.n44 plus.n43 0.189894
R320 plus.n43 plus.n42 0.189894
R321 plus.n42 plus.n33 0.189894
R322 plus.n34 plus.n33 0.189894
R323 plus.n37 plus.n34 0.189894
R324 drain_left.n10 drain_left.n8 80.4886
R325 drain_left.n6 drain_left.n4 80.4885
R326 drain_left.n2 drain_left.n0 80.4885
R327 drain_left.n16 drain_left.n15 79.7731
R328 drain_left.n14 drain_left.n13 79.7731
R329 drain_left.n12 drain_left.n11 79.7731
R330 drain_left.n10 drain_left.n9 79.7731
R331 drain_left.n7 drain_left.n3 79.773
R332 drain_left.n6 drain_left.n5 79.773
R333 drain_left.n2 drain_left.n1 79.773
R334 drain_left drain_left.n7 26.273
R335 drain_left.n3 drain_left.t13 6.6005
R336 drain_left.n3 drain_left.t5 6.6005
R337 drain_left.n4 drain_left.t11 6.6005
R338 drain_left.n4 drain_left.t15 6.6005
R339 drain_left.n5 drain_left.t10 6.6005
R340 drain_left.n5 drain_left.t17 6.6005
R341 drain_left.n1 drain_left.t19 6.6005
R342 drain_left.n1 drain_left.t9 6.6005
R343 drain_left.n0 drain_left.t1 6.6005
R344 drain_left.n0 drain_left.t6 6.6005
R345 drain_left.n15 drain_left.t18 6.6005
R346 drain_left.n15 drain_left.t8 6.6005
R347 drain_left.n13 drain_left.t12 6.6005
R348 drain_left.n13 drain_left.t3 6.6005
R349 drain_left.n11 drain_left.t4 6.6005
R350 drain_left.n11 drain_left.t0 6.6005
R351 drain_left.n9 drain_left.t2 6.6005
R352 drain_left.n9 drain_left.t14 6.6005
R353 drain_left.n8 drain_left.t16 6.6005
R354 drain_left.n8 drain_left.t7 6.6005
R355 drain_left drain_left.n16 6.36873
R356 drain_left.n12 drain_left.n10 0.716017
R357 drain_left.n14 drain_left.n12 0.716017
R358 drain_left.n16 drain_left.n14 0.716017
R359 drain_left.n7 drain_left.n6 0.660671
R360 drain_left.n7 drain_left.n2 0.660671
C0 drain_right plus 0.4139f
C1 drain_right drain_left 1.35857f
C2 drain_right source 9.9473f
C3 plus minus 4.66013f
C4 minus drain_left 0.178236f
C5 minus source 3.49562f
C6 plus drain_left 3.29477f
C7 plus source 3.50962f
C8 source drain_left 9.94598f
C9 drain_right minus 3.04308f
C10 drain_right a_n2542_n1488# 5.16873f
C11 drain_left a_n2542_n1488# 5.55402f
C12 source a_n2542_n1488# 3.949537f
C13 minus a_n2542_n1488# 9.377056f
C14 plus a_n2542_n1488# 10.80179f
C15 drain_left.t1 a_n2542_n1488# 0.068382f
C16 drain_left.t6 a_n2542_n1488# 0.068382f
C17 drain_left.n0 a_n2542_n1488# 0.496502f
C18 drain_left.t19 a_n2542_n1488# 0.068382f
C19 drain_left.t9 a_n2542_n1488# 0.068382f
C20 drain_left.n1 a_n2542_n1488# 0.493163f
C21 drain_left.n2 a_n2542_n1488# 0.731956f
C22 drain_left.t13 a_n2542_n1488# 0.068382f
C23 drain_left.t5 a_n2542_n1488# 0.068382f
C24 drain_left.n3 a_n2542_n1488# 0.493163f
C25 drain_left.t11 a_n2542_n1488# 0.068382f
C26 drain_left.t15 a_n2542_n1488# 0.068382f
C27 drain_left.n4 a_n2542_n1488# 0.496502f
C28 drain_left.t10 a_n2542_n1488# 0.068382f
C29 drain_left.t17 a_n2542_n1488# 0.068382f
C30 drain_left.n5 a_n2542_n1488# 0.493163f
C31 drain_left.n6 a_n2542_n1488# 0.731956f
C32 drain_left.n7 a_n2542_n1488# 1.38701f
C33 drain_left.t16 a_n2542_n1488# 0.068382f
C34 drain_left.t7 a_n2542_n1488# 0.068382f
C35 drain_left.n8 a_n2542_n1488# 0.496504f
C36 drain_left.t2 a_n2542_n1488# 0.068382f
C37 drain_left.t14 a_n2542_n1488# 0.068382f
C38 drain_left.n9 a_n2542_n1488# 0.493166f
C39 drain_left.n10 a_n2542_n1488# 0.736083f
C40 drain_left.t4 a_n2542_n1488# 0.068382f
C41 drain_left.t0 a_n2542_n1488# 0.068382f
C42 drain_left.n11 a_n2542_n1488# 0.493166f
C43 drain_left.n12 a_n2542_n1488# 0.363901f
C44 drain_left.t12 a_n2542_n1488# 0.068382f
C45 drain_left.t3 a_n2542_n1488# 0.068382f
C46 drain_left.n13 a_n2542_n1488# 0.493166f
C47 drain_left.n14 a_n2542_n1488# 0.363901f
C48 drain_left.t18 a_n2542_n1488# 0.068382f
C49 drain_left.t8 a_n2542_n1488# 0.068382f
C50 drain_left.n15 a_n2542_n1488# 0.493166f
C51 drain_left.n16 a_n2542_n1488# 0.611718f
C52 plus.n0 a_n2542_n1488# 0.04672f
C53 plus.t11 a_n2542_n1488# 0.210145f
C54 plus.t1 a_n2542_n1488# 0.210145f
C55 plus.t16 a_n2542_n1488# 0.210145f
C56 plus.n1 a_n2542_n1488# 0.130936f
C57 plus.n2 a_n2542_n1488# 0.04672f
C58 plus.t7 a_n2542_n1488# 0.210145f
C59 plus.t19 a_n2542_n1488# 0.210145f
C60 plus.n3 a_n2542_n1488# 0.04672f
C61 plus.t15 a_n2542_n1488# 0.210145f
C62 plus.n4 a_n2542_n1488# 0.130792f
C63 plus.n5 a_n2542_n1488# 0.04672f
C64 plus.t5 a_n2542_n1488# 0.210145f
C65 plus.t17 a_n2542_n1488# 0.210145f
C66 plus.n6 a_n2542_n1488# 0.04672f
C67 plus.t12 a_n2542_n1488# 0.210145f
C68 plus.n7 a_n2542_n1488# 0.130504f
C69 plus.t3 a_n2542_n1488# 0.220982f
C70 plus.n8 a_n2542_n1488# 0.11556f
C71 plus.n9 a_n2542_n1488# 0.15334f
C72 plus.n10 a_n2542_n1488# 0.010602f
C73 plus.n11 a_n2542_n1488# 0.130936f
C74 plus.n12 a_n2542_n1488# 0.010602f
C75 plus.n13 a_n2542_n1488# 0.126183f
C76 plus.n14 a_n2542_n1488# 0.04672f
C77 plus.n15 a_n2542_n1488# 0.04672f
C78 plus.n16 a_n2542_n1488# 0.04672f
C79 plus.n17 a_n2542_n1488# 0.010602f
C80 plus.n18 a_n2542_n1488# 0.130792f
C81 plus.n19 a_n2542_n1488# 0.126183f
C82 plus.n20 a_n2542_n1488# 0.010602f
C83 plus.n21 a_n2542_n1488# 0.04672f
C84 plus.n22 a_n2542_n1488# 0.04672f
C85 plus.n23 a_n2542_n1488# 0.04672f
C86 plus.n24 a_n2542_n1488# 0.010602f
C87 plus.n25 a_n2542_n1488# 0.130504f
C88 plus.n26 a_n2542_n1488# 0.126039f
C89 plus.n27 a_n2542_n1488# 0.359543f
C90 plus.n28 a_n2542_n1488# 0.04672f
C91 plus.t18 a_n2542_n1488# 0.210145f
C92 plus.t13 a_n2542_n1488# 0.210145f
C93 plus.t0 a_n2542_n1488# 0.210145f
C94 plus.n29 a_n2542_n1488# 0.130936f
C95 plus.n30 a_n2542_n1488# 0.04672f
C96 plus.t10 a_n2542_n1488# 0.210145f
C97 plus.n31 a_n2542_n1488# 0.04672f
C98 plus.t6 a_n2542_n1488# 0.210145f
C99 plus.t14 a_n2542_n1488# 0.210145f
C100 plus.n32 a_n2542_n1488# 0.130792f
C101 plus.n33 a_n2542_n1488# 0.04672f
C102 plus.t9 a_n2542_n1488# 0.210145f
C103 plus.n34 a_n2542_n1488# 0.04672f
C104 plus.t2 a_n2542_n1488# 0.210145f
C105 plus.t8 a_n2542_n1488# 0.210145f
C106 plus.n35 a_n2542_n1488# 0.130504f
C107 plus.t4 a_n2542_n1488# 0.220982f
C108 plus.n36 a_n2542_n1488# 0.11556f
C109 plus.n37 a_n2542_n1488# 0.15334f
C110 plus.n38 a_n2542_n1488# 0.010602f
C111 plus.n39 a_n2542_n1488# 0.130936f
C112 plus.n40 a_n2542_n1488# 0.010602f
C113 plus.n41 a_n2542_n1488# 0.126183f
C114 plus.n42 a_n2542_n1488# 0.04672f
C115 plus.n43 a_n2542_n1488# 0.04672f
C116 plus.n44 a_n2542_n1488# 0.04672f
C117 plus.n45 a_n2542_n1488# 0.010602f
C118 plus.n46 a_n2542_n1488# 0.130792f
C119 plus.n47 a_n2542_n1488# 0.126183f
C120 plus.n48 a_n2542_n1488# 0.010602f
C121 plus.n49 a_n2542_n1488# 0.04672f
C122 plus.n50 a_n2542_n1488# 0.04672f
C123 plus.n51 a_n2542_n1488# 0.04672f
C124 plus.n52 a_n2542_n1488# 0.010602f
C125 plus.n53 a_n2542_n1488# 0.130504f
C126 plus.n54 a_n2542_n1488# 0.126039f
C127 plus.n55 a_n2542_n1488# 1.27663f
C128 drain_right.t14 a_n2542_n1488# 0.067404f
C129 drain_right.t10 a_n2542_n1488# 0.067404f
C130 drain_right.n0 a_n2542_n1488# 0.489401f
C131 drain_right.t17 a_n2542_n1488# 0.067404f
C132 drain_right.t12 a_n2542_n1488# 0.067404f
C133 drain_right.n1 a_n2542_n1488# 0.48611f
C134 drain_right.n2 a_n2542_n1488# 0.721488f
C135 drain_right.t2 a_n2542_n1488# 0.067404f
C136 drain_right.t9 a_n2542_n1488# 0.067404f
C137 drain_right.n3 a_n2542_n1488# 0.48611f
C138 drain_right.t7 a_n2542_n1488# 0.067404f
C139 drain_right.t0 a_n2542_n1488# 0.067404f
C140 drain_right.n4 a_n2542_n1488# 0.489401f
C141 drain_right.t5 a_n2542_n1488# 0.067404f
C142 drain_right.t18 a_n2542_n1488# 0.067404f
C143 drain_right.n5 a_n2542_n1488# 0.48611f
C144 drain_right.n6 a_n2542_n1488# 0.721488f
C145 drain_right.n7 a_n2542_n1488# 1.3113f
C146 drain_right.t16 a_n2542_n1488# 0.067404f
C147 drain_right.t4 a_n2542_n1488# 0.067404f
C148 drain_right.n8 a_n2542_n1488# 0.489403f
C149 drain_right.t1 a_n2542_n1488# 0.067404f
C150 drain_right.t11 a_n2542_n1488# 0.067404f
C151 drain_right.n9 a_n2542_n1488# 0.486113f
C152 drain_right.n10 a_n2542_n1488# 0.725556f
C153 drain_right.t8 a_n2542_n1488# 0.067404f
C154 drain_right.t13 a_n2542_n1488# 0.067404f
C155 drain_right.n11 a_n2542_n1488# 0.486113f
C156 drain_right.n12 a_n2542_n1488# 0.358697f
C157 drain_right.t6 a_n2542_n1488# 0.067404f
C158 drain_right.t19 a_n2542_n1488# 0.067404f
C159 drain_right.n13 a_n2542_n1488# 0.486113f
C160 drain_right.n14 a_n2542_n1488# 0.358697f
C161 drain_right.t15 a_n2542_n1488# 0.067404f
C162 drain_right.t3 a_n2542_n1488# 0.067404f
C163 drain_right.n15 a_n2542_n1488# 0.486113f
C164 drain_right.n16 a_n2542_n1488# 0.602969f
C165 source.t10 a_n2542_n1488# 0.585974f
C166 source.n0 a_n2542_n1488# 0.828551f
C167 source.t12 a_n2542_n1488# 0.070567f
C168 source.t8 a_n2542_n1488# 0.070567f
C169 source.n1 a_n2542_n1488# 0.447434f
C170 source.n2 a_n2542_n1488# 0.396559f
C171 source.t1 a_n2542_n1488# 0.070567f
C172 source.t14 a_n2542_n1488# 0.070567f
C173 source.n3 a_n2542_n1488# 0.447434f
C174 source.n4 a_n2542_n1488# 0.396559f
C175 source.t7 a_n2542_n1488# 0.070567f
C176 source.t5 a_n2542_n1488# 0.070567f
C177 source.n5 a_n2542_n1488# 0.447434f
C178 source.n6 a_n2542_n1488# 0.396559f
C179 source.t13 a_n2542_n1488# 0.070567f
C180 source.t15 a_n2542_n1488# 0.070567f
C181 source.n7 a_n2542_n1488# 0.447434f
C182 source.n8 a_n2542_n1488# 0.396559f
C183 source.t38 a_n2542_n1488# 0.585974f
C184 source.n9 a_n2542_n1488# 0.426909f
C185 source.t34 a_n2542_n1488# 0.585974f
C186 source.n10 a_n2542_n1488# 0.426909f
C187 source.t28 a_n2542_n1488# 0.070567f
C188 source.t32 a_n2542_n1488# 0.070567f
C189 source.n11 a_n2542_n1488# 0.447434f
C190 source.n12 a_n2542_n1488# 0.396559f
C191 source.t23 a_n2542_n1488# 0.070567f
C192 source.t29 a_n2542_n1488# 0.070567f
C193 source.n13 a_n2542_n1488# 0.447434f
C194 source.n14 a_n2542_n1488# 0.396559f
C195 source.t37 a_n2542_n1488# 0.070567f
C196 source.t22 a_n2542_n1488# 0.070567f
C197 source.n15 a_n2542_n1488# 0.447434f
C198 source.n16 a_n2542_n1488# 0.396559f
C199 source.t30 a_n2542_n1488# 0.070567f
C200 source.t19 a_n2542_n1488# 0.070567f
C201 source.n17 a_n2542_n1488# 0.447434f
C202 source.n18 a_n2542_n1488# 0.396559f
C203 source.t35 a_n2542_n1488# 0.585974f
C204 source.n19 a_n2542_n1488# 1.14281f
C205 source.t3 a_n2542_n1488# 0.585971f
C206 source.n20 a_n2542_n1488# 1.14282f
C207 source.t4 a_n2542_n1488# 0.070567f
C208 source.t6 a_n2542_n1488# 0.070567f
C209 source.n21 a_n2542_n1488# 0.447431f
C210 source.n22 a_n2542_n1488# 0.396563f
C211 source.t2 a_n2542_n1488# 0.070567f
C212 source.t11 a_n2542_n1488# 0.070567f
C213 source.n23 a_n2542_n1488# 0.447431f
C214 source.n24 a_n2542_n1488# 0.396563f
C215 source.t17 a_n2542_n1488# 0.070567f
C216 source.t16 a_n2542_n1488# 0.070567f
C217 source.n25 a_n2542_n1488# 0.447431f
C218 source.n26 a_n2542_n1488# 0.396563f
C219 source.t39 a_n2542_n1488# 0.070567f
C220 source.t0 a_n2542_n1488# 0.070567f
C221 source.n27 a_n2542_n1488# 0.447431f
C222 source.n28 a_n2542_n1488# 0.396563f
C223 source.t9 a_n2542_n1488# 0.585971f
C224 source.n29 a_n2542_n1488# 0.426912f
C225 source.t36 a_n2542_n1488# 0.585971f
C226 source.n30 a_n2542_n1488# 0.426912f
C227 source.t24 a_n2542_n1488# 0.070567f
C228 source.t25 a_n2542_n1488# 0.070567f
C229 source.n31 a_n2542_n1488# 0.447431f
C230 source.n32 a_n2542_n1488# 0.396563f
C231 source.t27 a_n2542_n1488# 0.070567f
C232 source.t31 a_n2542_n1488# 0.070567f
C233 source.n33 a_n2542_n1488# 0.447431f
C234 source.n34 a_n2542_n1488# 0.396563f
C235 source.t20 a_n2542_n1488# 0.070567f
C236 source.t21 a_n2542_n1488# 0.070567f
C237 source.n35 a_n2542_n1488# 0.447431f
C238 source.n36 a_n2542_n1488# 0.396563f
C239 source.t33 a_n2542_n1488# 0.070567f
C240 source.t18 a_n2542_n1488# 0.070567f
C241 source.n37 a_n2542_n1488# 0.447431f
C242 source.n38 a_n2542_n1488# 0.396563f
C243 source.t26 a_n2542_n1488# 0.585971f
C244 source.n39 a_n2542_n1488# 0.608085f
C245 source.n40 a_n2542_n1488# 0.870166f
C246 minus.n0 a_n2542_n1488# 0.04513f
C247 minus.t13 a_n2542_n1488# 0.202995f
C248 minus.n1 a_n2542_n1488# 0.126481f
C249 minus.n2 a_n2542_n1488# 0.04513f
C250 minus.n3 a_n2542_n1488# 0.010241f
C251 minus.t11 a_n2542_n1488# 0.202995f
C252 minus.n4 a_n2542_n1488# 0.04513f
C253 minus.t8 a_n2542_n1488# 0.202995f
C254 minus.n5 a_n2542_n1488# 0.126481f
C255 minus.t15 a_n2542_n1488# 0.213464f
C256 minus.n6 a_n2542_n1488# 0.111628f
C257 minus.t3 a_n2542_n1488# 0.202995f
C258 minus.n7 a_n2542_n1488# 0.126064f
C259 minus.n8 a_n2542_n1488# 0.010241f
C260 minus.n9 a_n2542_n1488# 0.148123f
C261 minus.n10 a_n2542_n1488# 0.04513f
C262 minus.n11 a_n2542_n1488# 0.04513f
C263 minus.n12 a_n2542_n1488# 0.010241f
C264 minus.t18 a_n2542_n1488# 0.202995f
C265 minus.n13 a_n2542_n1488# 0.12189f
C266 minus.t6 a_n2542_n1488# 0.202995f
C267 minus.n14 a_n2542_n1488# 0.126342f
C268 minus.n15 a_n2542_n1488# 0.04513f
C269 minus.n16 a_n2542_n1488# 0.04513f
C270 minus.n17 a_n2542_n1488# 0.04513f
C271 minus.n18 a_n2542_n1488# 0.126342f
C272 minus.t0 a_n2542_n1488# 0.202995f
C273 minus.n19 a_n2542_n1488# 0.12189f
C274 minus.n20 a_n2542_n1488# 0.010241f
C275 minus.n21 a_n2542_n1488# 0.04513f
C276 minus.n22 a_n2542_n1488# 0.04513f
C277 minus.n23 a_n2542_n1488# 0.04513f
C278 minus.n24 a_n2542_n1488# 0.010241f
C279 minus.t16 a_n2542_n1488# 0.202995f
C280 minus.n25 a_n2542_n1488# 0.126064f
C281 minus.t4 a_n2542_n1488# 0.202995f
C282 minus.n26 a_n2542_n1488# 0.121751f
C283 minus.n27 a_n2542_n1488# 1.31368f
C284 minus.n28 a_n2542_n1488# 0.04513f
C285 minus.t1 a_n2542_n1488# 0.202995f
C286 minus.n29 a_n2542_n1488# 0.126481f
C287 minus.n30 a_n2542_n1488# 0.04513f
C288 minus.n31 a_n2542_n1488# 0.010241f
C289 minus.n32 a_n2542_n1488# 0.04513f
C290 minus.t2 a_n2542_n1488# 0.202995f
C291 minus.n33 a_n2542_n1488# 0.126481f
C292 minus.t5 a_n2542_n1488# 0.213464f
C293 minus.n34 a_n2542_n1488# 0.111628f
C294 minus.t9 a_n2542_n1488# 0.202995f
C295 minus.n35 a_n2542_n1488# 0.126064f
C296 minus.n36 a_n2542_n1488# 0.010241f
C297 minus.n37 a_n2542_n1488# 0.148123f
C298 minus.n38 a_n2542_n1488# 0.04513f
C299 minus.n39 a_n2542_n1488# 0.04513f
C300 minus.n40 a_n2542_n1488# 0.010241f
C301 minus.t7 a_n2542_n1488# 0.202995f
C302 minus.n41 a_n2542_n1488# 0.12189f
C303 minus.t17 a_n2542_n1488# 0.202995f
C304 minus.n42 a_n2542_n1488# 0.126342f
C305 minus.n43 a_n2542_n1488# 0.04513f
C306 minus.n44 a_n2542_n1488# 0.04513f
C307 minus.n45 a_n2542_n1488# 0.04513f
C308 minus.t10 a_n2542_n1488# 0.202995f
C309 minus.n46 a_n2542_n1488# 0.126342f
C310 minus.t14 a_n2542_n1488# 0.202995f
C311 minus.n47 a_n2542_n1488# 0.12189f
C312 minus.n48 a_n2542_n1488# 0.010241f
C313 minus.n49 a_n2542_n1488# 0.04513f
C314 minus.n50 a_n2542_n1488# 0.04513f
C315 minus.n51 a_n2542_n1488# 0.04513f
C316 minus.n52 a_n2542_n1488# 0.010241f
C317 minus.t12 a_n2542_n1488# 0.202995f
C318 minus.n53 a_n2542_n1488# 0.126064f
C319 minus.t19 a_n2542_n1488# 0.202995f
C320 minus.n54 a_n2542_n1488# 0.121751f
C321 minus.n55 a_n2542_n1488# 0.304728f
C322 minus.n56 a_n2542_n1488# 1.60973f
.ends

