* NGSPICE file created from diffpair143.ext - technology: sky130A

.subckt diffpair143 minus drain_right drain_left source plus
X0 a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X1 source.t15 plus.t0 drain_left.t1 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X2 source.t7 minus.t0 drain_right.t7 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 drain_left.t0 plus.t1 source.t14 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X4 source.t13 plus.t2 drain_left.t3 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X5 a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X6 source.t12 plus.t3 drain_left.t2 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X7 drain_right.t6 minus.t1 source.t6 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X8 drain_left.t4 plus.t4 source.t11 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X9 drain_right.t5 minus.t2 source.t3 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X10 drain_right.t4 minus.t3 source.t5 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X11 source.t4 minus.t4 drain_right.t3 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X12 drain_left.t5 plus.t5 source.t10 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X14 a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X15 drain_right.t2 minus.t5 source.t1 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X16 source.t2 minus.t6 drain_right.t1 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X17 source.t9 plus.t6 drain_left.t6 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X18 drain_left.t7 plus.t7 source.t8 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X19 source.t0 minus.t7 drain_right.t0 a_n1746_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
R0 plus.n5 plus.n4 161.3
R1 plus.n6 plus.n1 161.3
R2 plus.n7 plus.n0 161.3
R3 plus.n9 plus.n8 161.3
R4 plus.n15 plus.n14 161.3
R5 plus.n16 plus.n11 161.3
R6 plus.n17 plus.n10 161.3
R7 plus.n19 plus.n18 161.3
R8 plus.n3 plus.t2 147.155
R9 plus.n13 plus.t7 147.155
R10 plus.n8 plus.t4 124.977
R11 plus.n6 plus.t0 124.977
R12 plus.n2 plus.t5 124.977
R13 plus.n18 plus.t3 124.977
R14 plus.n16 plus.t1 124.977
R15 plus.n12 plus.t6 124.977
R16 plus.n4 plus.n3 44.862
R17 plus.n14 plus.n13 44.862
R18 plus.n8 plus.n7 28.4823
R19 plus.n18 plus.n17 28.4823
R20 plus plus.n19 25.9611
R21 plus.n5 plus.n2 24.1005
R22 plus.n6 plus.n5 24.1005
R23 plus.n16 plus.n15 24.1005
R24 plus.n15 plus.n12 24.1005
R25 plus.n7 plus.n6 19.7187
R26 plus.n17 plus.n16 19.7187
R27 plus.n3 plus.n2 19.7081
R28 plus.n13 plus.n12 19.7081
R29 plus plus.n9 8.48914
R30 plus.n4 plus.n1 0.189894
R31 plus.n1 plus.n0 0.189894
R32 plus.n9 plus.n0 0.189894
R33 plus.n19 plus.n10 0.189894
R34 plus.n11 plus.n10 0.189894
R35 plus.n14 plus.n11 0.189894
R36 drain_left.n5 drain_left.n3 101.683
R37 drain_left.n2 drain_left.n1 101.184
R38 drain_left.n2 drain_left.n0 101.184
R39 drain_left.n5 drain_left.n4 100.796
R40 drain_left drain_left.n2 22.8991
R41 drain_left.n1 drain_left.t6 9.9005
R42 drain_left.n1 drain_left.t7 9.9005
R43 drain_left.n0 drain_left.t2 9.9005
R44 drain_left.n0 drain_left.t0 9.9005
R45 drain_left.n4 drain_left.t1 9.9005
R46 drain_left.n4 drain_left.t4 9.9005
R47 drain_left.n3 drain_left.t3 9.9005
R48 drain_left.n3 drain_left.t5 9.9005
R49 drain_left drain_left.n5 6.54115
R50 source.n66 source.n64 289.615
R51 source.n56 source.n54 289.615
R52 source.n48 source.n46 289.615
R53 source.n38 source.n36 289.615
R54 source.n2 source.n0 289.615
R55 source.n12 source.n10 289.615
R56 source.n20 source.n18 289.615
R57 source.n30 source.n28 289.615
R58 source.n67 source.n66 185
R59 source.n57 source.n56 185
R60 source.n49 source.n48 185
R61 source.n39 source.n38 185
R62 source.n3 source.n2 185
R63 source.n13 source.n12 185
R64 source.n21 source.n20 185
R65 source.n31 source.n30 185
R66 source.t1 source.n65 167.117
R67 source.t4 source.n55 167.117
R68 source.t8 source.n47 167.117
R69 source.t12 source.n37 167.117
R70 source.t11 source.n1 167.117
R71 source.t13 source.n11 167.117
R72 source.t5 source.n19 167.117
R73 source.t0 source.n29 167.117
R74 source.n9 source.n8 84.1169
R75 source.n27 source.n26 84.1169
R76 source.n63 source.n62 84.1168
R77 source.n45 source.n44 84.1168
R78 source.n66 source.t1 52.3082
R79 source.n56 source.t4 52.3082
R80 source.n48 source.t8 52.3082
R81 source.n38 source.t12 52.3082
R82 source.n2 source.t11 52.3082
R83 source.n12 source.t13 52.3082
R84 source.n20 source.t5 52.3082
R85 source.n30 source.t0 52.3082
R86 source.n71 source.n70 31.4096
R87 source.n61 source.n60 31.4096
R88 source.n53 source.n52 31.4096
R89 source.n43 source.n42 31.4096
R90 source.n7 source.n6 31.4096
R91 source.n17 source.n16 31.4096
R92 source.n25 source.n24 31.4096
R93 source.n35 source.n34 31.4096
R94 source.n43 source.n35 14.5999
R95 source.n62 source.t3 9.9005
R96 source.n62 source.t2 9.9005
R97 source.n44 source.t14 9.9005
R98 source.n44 source.t9 9.9005
R99 source.n8 source.t10 9.9005
R100 source.n8 source.t15 9.9005
R101 source.n26 source.t6 9.9005
R102 source.n26 source.t7 9.9005
R103 source.n67 source.n65 9.71174
R104 source.n57 source.n55 9.71174
R105 source.n49 source.n47 9.71174
R106 source.n39 source.n37 9.71174
R107 source.n3 source.n1 9.71174
R108 source.n13 source.n11 9.71174
R109 source.n21 source.n19 9.71174
R110 source.n31 source.n29 9.71174
R111 source.n70 source.n69 9.45567
R112 source.n60 source.n59 9.45567
R113 source.n52 source.n51 9.45567
R114 source.n42 source.n41 9.45567
R115 source.n6 source.n5 9.45567
R116 source.n16 source.n15 9.45567
R117 source.n24 source.n23 9.45567
R118 source.n34 source.n33 9.45567
R119 source.n69 source.n68 9.3005
R120 source.n59 source.n58 9.3005
R121 source.n51 source.n50 9.3005
R122 source.n41 source.n40 9.3005
R123 source.n5 source.n4 9.3005
R124 source.n15 source.n14 9.3005
R125 source.n23 source.n22 9.3005
R126 source.n33 source.n32 9.3005
R127 source.n72 source.n7 8.893
R128 source.n70 source.n64 8.14595
R129 source.n60 source.n54 8.14595
R130 source.n52 source.n46 8.14595
R131 source.n42 source.n36 8.14595
R132 source.n6 source.n0 8.14595
R133 source.n16 source.n10 8.14595
R134 source.n24 source.n18 8.14595
R135 source.n34 source.n28 8.14595
R136 source.n68 source.n67 7.3702
R137 source.n58 source.n57 7.3702
R138 source.n50 source.n49 7.3702
R139 source.n40 source.n39 7.3702
R140 source.n4 source.n3 7.3702
R141 source.n14 source.n13 7.3702
R142 source.n22 source.n21 7.3702
R143 source.n32 source.n31 7.3702
R144 source.n68 source.n64 5.81868
R145 source.n58 source.n54 5.81868
R146 source.n50 source.n46 5.81868
R147 source.n40 source.n36 5.81868
R148 source.n4 source.n0 5.81868
R149 source.n14 source.n10 5.81868
R150 source.n22 source.n18 5.81868
R151 source.n32 source.n28 5.81868
R152 source.n72 source.n71 5.7074
R153 source.n69 source.n65 3.44771
R154 source.n59 source.n55 3.44771
R155 source.n51 source.n47 3.44771
R156 source.n41 source.n37 3.44771
R157 source.n5 source.n1 3.44771
R158 source.n15 source.n11 3.44771
R159 source.n23 source.n19 3.44771
R160 source.n33 source.n29 3.44771
R161 source.n35 source.n27 0.888431
R162 source.n27 source.n25 0.888431
R163 source.n17 source.n9 0.888431
R164 source.n9 source.n7 0.888431
R165 source.n45 source.n43 0.888431
R166 source.n53 source.n45 0.888431
R167 source.n63 source.n61 0.888431
R168 source.n71 source.n63 0.888431
R169 source.n25 source.n17 0.470328
R170 source.n61 source.n53 0.470328
R171 source source.n72 0.188
R172 minus.n9 minus.n8 161.3
R173 minus.n7 minus.n0 161.3
R174 minus.n6 minus.n5 161.3
R175 minus.n4 minus.n1 161.3
R176 minus.n19 minus.n18 161.3
R177 minus.n17 minus.n10 161.3
R178 minus.n16 minus.n15 161.3
R179 minus.n14 minus.n11 161.3
R180 minus.n3 minus.t3 147.155
R181 minus.n13 minus.t4 147.155
R182 minus.n2 minus.t0 124.977
R183 minus.n6 minus.t1 124.977
R184 minus.n8 minus.t7 124.977
R185 minus.n12 minus.t2 124.977
R186 minus.n16 minus.t6 124.977
R187 minus.n18 minus.t5 124.977
R188 minus.n4 minus.n3 44.862
R189 minus.n14 minus.n13 44.862
R190 minus.n8 minus.n7 28.4823
R191 minus.n18 minus.n17 28.4823
R192 minus.n20 minus.n9 28.2922
R193 minus.n6 minus.n1 24.1005
R194 minus.n2 minus.n1 24.1005
R195 minus.n12 minus.n11 24.1005
R196 minus.n16 minus.n11 24.1005
R197 minus.n7 minus.n6 19.7187
R198 minus.n17 minus.n16 19.7187
R199 minus.n3 minus.n2 19.7081
R200 minus.n13 minus.n12 19.7081
R201 minus.n20 minus.n19 6.63308
R202 minus.n9 minus.n0 0.189894
R203 minus.n5 minus.n0 0.189894
R204 minus.n5 minus.n4 0.189894
R205 minus.n15 minus.n14 0.189894
R206 minus.n15 minus.n10 0.189894
R207 minus.n19 minus.n10 0.189894
R208 minus minus.n20 0.188
R209 drain_right.n5 drain_right.n3 101.683
R210 drain_right.n2 drain_right.n1 101.184
R211 drain_right.n2 drain_right.n0 101.184
R212 drain_right.n5 drain_right.n4 100.796
R213 drain_right drain_right.n2 22.3458
R214 drain_right.n1 drain_right.t1 9.9005
R215 drain_right.n1 drain_right.t2 9.9005
R216 drain_right.n0 drain_right.t3 9.9005
R217 drain_right.n0 drain_right.t5 9.9005
R218 drain_right.n3 drain_right.t7 9.9005
R219 drain_right.n3 drain_right.t4 9.9005
R220 drain_right.n4 drain_right.t0 9.9005
R221 drain_right.n4 drain_right.t6 9.9005
R222 drain_right drain_right.n5 6.54115
C0 drain_left drain_right 0.821811f
C1 drain_right plus 0.329494f
C2 source minus 1.52017f
C3 drain_left minus 0.176866f
C4 minus plus 3.47516f
C5 drain_right minus 1.25313f
C6 drain_left source 3.6807f
C7 source plus 1.53414f
C8 source drain_right 3.68247f
C9 drain_left plus 1.42194f
C10 drain_right a_n1746_n1288# 3.29499f
C11 drain_left a_n1746_n1288# 3.51005f
C12 source a_n1746_n1288# 3.059775f
C13 minus a_n1746_n1288# 5.946295f
C14 plus a_n1746_n1288# 6.511153f
C15 drain_right.t3 a_n1746_n1288# 0.030393f
C16 drain_right.t5 a_n1746_n1288# 0.030393f
C17 drain_right.n0 a_n1746_n1288# 0.191842f
C18 drain_right.t1 a_n1746_n1288# 0.030393f
C19 drain_right.t2 a_n1746_n1288# 0.030393f
C20 drain_right.n1 a_n1746_n1288# 0.191842f
C21 drain_right.n2 a_n1746_n1288# 0.978797f
C22 drain_right.t7 a_n1746_n1288# 0.030393f
C23 drain_right.t4 a_n1746_n1288# 0.030393f
C24 drain_right.n3 a_n1746_n1288# 0.193254f
C25 drain_right.t0 a_n1746_n1288# 0.030393f
C26 drain_right.t6 a_n1746_n1288# 0.030393f
C27 drain_right.n4 a_n1746_n1288# 0.19094f
C28 drain_right.n5 a_n1746_n1288# 0.689986f
C29 minus.n0 a_n1746_n1288# 0.026429f
C30 minus.n1 a_n1746_n1288# 0.005997f
C31 minus.t1 a_n1746_n1288# 0.114582f
C32 minus.t3 a_n1746_n1288# 0.126566f
C33 minus.t0 a_n1746_n1288# 0.114582f
C34 minus.n2 a_n1746_n1288# 0.082042f
C35 minus.n3 a_n1746_n1288# 0.070098f
C36 minus.n4 a_n1746_n1288# 0.109906f
C37 minus.n5 a_n1746_n1288# 0.026429f
C38 minus.n6 a_n1746_n1288# 0.07965f
C39 minus.n7 a_n1746_n1288# 0.005997f
C40 minus.t7 a_n1746_n1288# 0.114582f
C41 minus.n8 a_n1746_n1288# 0.077939f
C42 minus.n9 a_n1746_n1288# 0.624576f
C43 minus.n10 a_n1746_n1288# 0.026429f
C44 minus.n11 a_n1746_n1288# 0.005997f
C45 minus.t4 a_n1746_n1288# 0.126566f
C46 minus.t2 a_n1746_n1288# 0.114582f
C47 minus.n12 a_n1746_n1288# 0.082042f
C48 minus.n13 a_n1746_n1288# 0.070098f
C49 minus.n14 a_n1746_n1288# 0.109906f
C50 minus.n15 a_n1746_n1288# 0.026429f
C51 minus.t6 a_n1746_n1288# 0.114582f
C52 minus.n16 a_n1746_n1288# 0.07965f
C53 minus.n17 a_n1746_n1288# 0.005997f
C54 minus.t5 a_n1746_n1288# 0.114582f
C55 minus.n18 a_n1746_n1288# 0.077939f
C56 minus.n19 a_n1746_n1288# 0.181023f
C57 minus.n20 a_n1746_n1288# 0.767445f
C58 source.n0 a_n1746_n1288# 0.027846f
C59 source.n1 a_n1746_n1288# 0.061613f
C60 source.t11 a_n1746_n1288# 0.046237f
C61 source.n2 a_n1746_n1288# 0.048221f
C62 source.n3 a_n1746_n1288# 0.015545f
C63 source.n4 a_n1746_n1288# 0.010252f
C64 source.n5 a_n1746_n1288# 0.135809f
C65 source.n6 a_n1746_n1288# 0.030526f
C66 source.n7 a_n1746_n1288# 0.325609f
C67 source.t10 a_n1746_n1288# 0.030152f
C68 source.t15 a_n1746_n1288# 0.030152f
C69 source.n8 a_n1746_n1288# 0.161194f
C70 source.n9 a_n1746_n1288# 0.257495f
C71 source.n10 a_n1746_n1288# 0.027846f
C72 source.n11 a_n1746_n1288# 0.061613f
C73 source.t13 a_n1746_n1288# 0.046237f
C74 source.n12 a_n1746_n1288# 0.048221f
C75 source.n13 a_n1746_n1288# 0.015545f
C76 source.n14 a_n1746_n1288# 0.010252f
C77 source.n15 a_n1746_n1288# 0.135809f
C78 source.n16 a_n1746_n1288# 0.030526f
C79 source.n17 a_n1746_n1288# 0.099174f
C80 source.n18 a_n1746_n1288# 0.027846f
C81 source.n19 a_n1746_n1288# 0.061613f
C82 source.t5 a_n1746_n1288# 0.046237f
C83 source.n20 a_n1746_n1288# 0.048221f
C84 source.n21 a_n1746_n1288# 0.015545f
C85 source.n22 a_n1746_n1288# 0.010252f
C86 source.n23 a_n1746_n1288# 0.135809f
C87 source.n24 a_n1746_n1288# 0.030526f
C88 source.n25 a_n1746_n1288# 0.099174f
C89 source.t6 a_n1746_n1288# 0.030152f
C90 source.t7 a_n1746_n1288# 0.030152f
C91 source.n26 a_n1746_n1288# 0.161194f
C92 source.n27 a_n1746_n1288# 0.257495f
C93 source.n28 a_n1746_n1288# 0.027846f
C94 source.n29 a_n1746_n1288# 0.061613f
C95 source.t0 a_n1746_n1288# 0.046237f
C96 source.n30 a_n1746_n1288# 0.048221f
C97 source.n31 a_n1746_n1288# 0.015545f
C98 source.n32 a_n1746_n1288# 0.010252f
C99 source.n33 a_n1746_n1288# 0.135809f
C100 source.n34 a_n1746_n1288# 0.030526f
C101 source.n35 a_n1746_n1288# 0.508315f
C102 source.n36 a_n1746_n1288# 0.027846f
C103 source.n37 a_n1746_n1288# 0.061613f
C104 source.t12 a_n1746_n1288# 0.046237f
C105 source.n38 a_n1746_n1288# 0.048221f
C106 source.n39 a_n1746_n1288# 0.015545f
C107 source.n40 a_n1746_n1288# 0.010252f
C108 source.n41 a_n1746_n1288# 0.135809f
C109 source.n42 a_n1746_n1288# 0.030526f
C110 source.n43 a_n1746_n1288# 0.508315f
C111 source.t14 a_n1746_n1288# 0.030152f
C112 source.t9 a_n1746_n1288# 0.030152f
C113 source.n44 a_n1746_n1288# 0.161193f
C114 source.n45 a_n1746_n1288# 0.257496f
C115 source.n46 a_n1746_n1288# 0.027846f
C116 source.n47 a_n1746_n1288# 0.061613f
C117 source.t8 a_n1746_n1288# 0.046237f
C118 source.n48 a_n1746_n1288# 0.048221f
C119 source.n49 a_n1746_n1288# 0.015545f
C120 source.n50 a_n1746_n1288# 0.010252f
C121 source.n51 a_n1746_n1288# 0.135809f
C122 source.n52 a_n1746_n1288# 0.030526f
C123 source.n53 a_n1746_n1288# 0.099174f
C124 source.n54 a_n1746_n1288# 0.027846f
C125 source.n55 a_n1746_n1288# 0.061613f
C126 source.t4 a_n1746_n1288# 0.046237f
C127 source.n56 a_n1746_n1288# 0.048221f
C128 source.n57 a_n1746_n1288# 0.015545f
C129 source.n58 a_n1746_n1288# 0.010252f
C130 source.n59 a_n1746_n1288# 0.135809f
C131 source.n60 a_n1746_n1288# 0.030526f
C132 source.n61 a_n1746_n1288# 0.099174f
C133 source.t3 a_n1746_n1288# 0.030152f
C134 source.t2 a_n1746_n1288# 0.030152f
C135 source.n62 a_n1746_n1288# 0.161193f
C136 source.n63 a_n1746_n1288# 0.257496f
C137 source.n64 a_n1746_n1288# 0.027846f
C138 source.n65 a_n1746_n1288# 0.061613f
C139 source.t1 a_n1746_n1288# 0.046237f
C140 source.n66 a_n1746_n1288# 0.048221f
C141 source.n67 a_n1746_n1288# 0.015545f
C142 source.n68 a_n1746_n1288# 0.010252f
C143 source.n69 a_n1746_n1288# 0.135809f
C144 source.n70 a_n1746_n1288# 0.030526f
C145 source.n71 a_n1746_n1288# 0.223622f
C146 source.n72 a_n1746_n1288# 0.480969f
C147 drain_left.t2 a_n1746_n1288# 0.029788f
C148 drain_left.t0 a_n1746_n1288# 0.029788f
C149 drain_left.n0 a_n1746_n1288# 0.188019f
C150 drain_left.t6 a_n1746_n1288# 0.029788f
C151 drain_left.t7 a_n1746_n1288# 0.029788f
C152 drain_left.n1 a_n1746_n1288# 0.188019f
C153 drain_left.n2 a_n1746_n1288# 0.996261f
C154 drain_left.t3 a_n1746_n1288# 0.029788f
C155 drain_left.t5 a_n1746_n1288# 0.029788f
C156 drain_left.n3 a_n1746_n1288# 0.189403f
C157 drain_left.t1 a_n1746_n1288# 0.029788f
C158 drain_left.t4 a_n1746_n1288# 0.029788f
C159 drain_left.n4 a_n1746_n1288# 0.187135f
C160 drain_left.n5 a_n1746_n1288# 0.676237f
C161 plus.n0 a_n1746_n1288# 0.026839f
C162 plus.t4 a_n1746_n1288# 0.116359f
C163 plus.t0 a_n1746_n1288# 0.116359f
C164 plus.n1 a_n1746_n1288# 0.026839f
C165 plus.t5 a_n1746_n1288# 0.116359f
C166 plus.n2 a_n1746_n1288# 0.083314f
C167 plus.t2 a_n1746_n1288# 0.128529f
C168 plus.n3 a_n1746_n1288# 0.071185f
C169 plus.n4 a_n1746_n1288# 0.11161f
C170 plus.n5 a_n1746_n1288# 0.00609f
C171 plus.n6 a_n1746_n1288# 0.080885f
C172 plus.n7 a_n1746_n1288# 0.00609f
C173 plus.n8 a_n1746_n1288# 0.079148f
C174 plus.n9 a_n1746_n1288# 0.20069f
C175 plus.n10 a_n1746_n1288# 0.026839f
C176 plus.t3 a_n1746_n1288# 0.116359f
C177 plus.n11 a_n1746_n1288# 0.026839f
C178 plus.t1 a_n1746_n1288# 0.116359f
C179 plus.t6 a_n1746_n1288# 0.116359f
C180 plus.n12 a_n1746_n1288# 0.083314f
C181 plus.t7 a_n1746_n1288# 0.128529f
C182 plus.n13 a_n1746_n1288# 0.071185f
C183 plus.n14 a_n1746_n1288# 0.11161f
C184 plus.n15 a_n1746_n1288# 0.00609f
C185 plus.n16 a_n1746_n1288# 0.080885f
C186 plus.n17 a_n1746_n1288# 0.00609f
C187 plus.n18 a_n1746_n1288# 0.079148f
C188 plus.n19 a_n1746_n1288# 0.606373f
.ends

