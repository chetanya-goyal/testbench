* NGSPICE file created from diffpair161.ext - technology: sky130A

.subckt diffpair161 minus drain_right drain_left source plus
X0 source minus drain_right a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X1 drain_right minus source a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X2 a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X3 source plus drain_left a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X4 drain_left plus source a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X5 drain_left plus source a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X6 drain_right minus source a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X7 a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X8 source plus drain_left a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X9 a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X10 a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X11 source minus drain_right a_n1106_n1492# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
.ends

