* NGSPICE file created from diffpair149.ext - technology: sky130A

.subckt diffpair149 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t28 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X1 source.t32 plus.t1 drain_left.t22 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X2 a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X3 drain_left.t21 plus.t2 source.t37 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X4 source.t31 plus.t3 drain_left.t20 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X5 source.t35 plus.t4 drain_left.t19 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X6 source.t9 minus.t0 drain_right.t23 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X7 drain_right.t22 minus.t1 source.t8 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X8 source.t46 minus.t2 drain_right.t21 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X9 drain_right.t20 minus.t3 source.t47 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X10 source.t3 minus.t4 drain_right.t19 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X11 drain_left.t18 plus.t5 source.t29 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X12 drain_left.t17 plus.t6 source.t33 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 source.t26 plus.t7 drain_left.t16 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X14 source.t39 plus.t8 drain_left.t15 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X15 drain_right.t18 minus.t5 source.t7 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X16 drain_right.t17 minus.t6 source.t2 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X17 source.t24 plus.t9 drain_left.t14 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X18 source.t12 minus.t7 drain_right.t16 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_right.t15 minus.t8 source.t15 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X20 drain_left.t13 plus.t10 source.t44 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X21 drain_left.t12 plus.t11 source.t40 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X22 source.t27 plus.t12 drain_left.t11 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 drain_right.t14 minus.t9 source.t6 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X24 drain_right.t13 minus.t10 source.t11 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X25 drain_left.t10 plus.t13 source.t41 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X26 drain_right.t12 minus.t11 source.t14 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X27 drain_left.t9 plus.t14 source.t43 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X28 drain_left.t8 plus.t15 source.t30 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X29 source.t34 plus.t16 drain_left.t7 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X30 source.t36 plus.t17 drain_left.t6 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X31 drain_left.t5 plus.t18 source.t23 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X32 drain_right.t11 minus.t12 source.t5 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X33 drain_right.t10 minus.t13 source.t19 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X34 a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X35 source.t1 minus.t14 drain_right.t9 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X36 drain_left.t4 plus.t19 source.t22 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X37 source.t4 minus.t15 drain_right.t8 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X38 source.t13 minus.t16 drain_right.t7 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X39 a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X40 source.t45 plus.t20 drain_left.t3 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X41 drain_right.t6 minus.t17 source.t16 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X42 source.t0 minus.t18 drain_right.t5 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X43 source.t20 minus.t19 drain_right.t4 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X44 drain_right.t3 minus.t20 source.t10 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X45 source.t18 minus.t21 drain_right.t2 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X46 source.t42 plus.t21 drain_left.t2 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X47 drain_left.t1 plus.t22 source.t38 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X48 source.t21 minus.t22 drain_right.t1 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X49 source.t17 minus.t23 drain_right.t0 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X50 source.t25 plus.t23 drain_left.t0 a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X51 a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# a_n3394_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
R0 plus.n13 plus.n12 161.3
R1 plus.n14 plus.n9 161.3
R2 plus.n16 plus.n15 161.3
R3 plus.n17 plus.n8 161.3
R4 plus.n19 plus.n18 161.3
R5 plus.n20 plus.n7 161.3
R6 plus.n22 plus.n21 161.3
R7 plus.n23 plus.n6 161.3
R8 plus.n25 plus.n24 161.3
R9 plus.n26 plus.n5 161.3
R10 plus.n28 plus.n27 161.3
R11 plus.n29 plus.n4 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n3 161.3
R14 plus.n34 plus.n33 161.3
R15 plus.n35 plus.n2 161.3
R16 plus.n37 plus.n36 161.3
R17 plus.n38 plus.n1 161.3
R18 plus.n39 plus.n0 161.3
R19 plus.n41 plus.n40 161.3
R20 plus.n55 plus.n54 161.3
R21 plus.n56 plus.n51 161.3
R22 plus.n58 plus.n57 161.3
R23 plus.n59 plus.n50 161.3
R24 plus.n61 plus.n60 161.3
R25 plus.n62 plus.n49 161.3
R26 plus.n64 plus.n63 161.3
R27 plus.n65 plus.n48 161.3
R28 plus.n67 plus.n66 161.3
R29 plus.n68 plus.n47 161.3
R30 plus.n70 plus.n69 161.3
R31 plus.n71 plus.n46 161.3
R32 plus.n73 plus.n72 161.3
R33 plus.n74 plus.n45 161.3
R34 plus.n76 plus.n75 161.3
R35 plus.n77 plus.n44 161.3
R36 plus.n79 plus.n78 161.3
R37 plus.n80 plus.n43 161.3
R38 plus.n81 plus.n42 161.3
R39 plus.n83 plus.n82 161.3
R40 plus.n11 plus.t8 151.334
R41 plus.n53 plus.t22 151.334
R42 plus.n40 plus.t2 124.977
R43 plus.n38 plus.t17 124.977
R44 plus.n2 plus.t6 124.977
R45 plus.n32 plus.t23 124.977
R46 plus.n4 plus.t13 124.977
R47 plus.n26 plus.t3 124.977
R48 plus.n6 plus.t18 124.977
R49 plus.n20 plus.t7 124.977
R50 plus.n8 plus.t15 124.977
R51 plus.n14 plus.t4 124.977
R52 plus.n10 plus.t19 124.977
R53 plus.n82 plus.t9 124.977
R54 plus.n80 plus.t10 124.977
R55 plus.n44 plus.t1 124.977
R56 plus.n74 plus.t0 124.977
R57 plus.n46 plus.t20 124.977
R58 plus.n68 plus.t14 124.977
R59 plus.n48 plus.t16 124.977
R60 plus.n62 plus.t11 124.977
R61 plus.n50 plus.t12 124.977
R62 plus.n56 plus.t5 124.977
R63 plus.n52 plus.t21 124.977
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus.n33 plus.n2 37.246
R73 plus.n15 plus.n14 37.246
R74 plus.n75 plus.n44 37.246
R75 plus.n57 plus.n56 37.246
R76 plus.n32 plus.n31 32.8641
R77 plus.n19 plus.n8 32.8641
R78 plus.n74 plus.n73 32.8641
R79 plus.n61 plus.n50 32.8641
R80 plus plus.n83 32.249
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus.n31 plus.n4 15.3369
R94 plus.n20 plus.n19 15.3369
R95 plus.n73 plus.n46 15.3369
R96 plus.n62 plus.n61 15.3369
R97 plus.n11 plus.n10 14.1472
R98 plus.n53 plus.n52 14.1472
R99 plus.n33 plus.n32 10.955
R100 plus.n15 plus.n8 10.955
R101 plus.n75 plus.n74 10.955
R102 plus.n57 plus.n50 10.955
R103 plus plus.n41 8.53459
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 source.n98 source.n96 289.615
R149 source.n80 source.n78 289.615
R150 source.n72 source.n70 289.615
R151 source.n54 source.n52 289.615
R152 source.n2 source.n0 289.615
R153 source.n20 source.n18 289.615
R154 source.n28 source.n26 289.615
R155 source.n46 source.n44 289.615
R156 source.n99 source.n98 185
R157 source.n81 source.n80 185
R158 source.n73 source.n72 185
R159 source.n55 source.n54 185
R160 source.n3 source.n2 185
R161 source.n21 source.n20 185
R162 source.n29 source.n28 185
R163 source.n47 source.n46 185
R164 source.t8 source.n97 167.117
R165 source.t1 source.n79 167.117
R166 source.t38 source.n71 167.117
R167 source.t24 source.n53 167.117
R168 source.t37 source.n1 167.117
R169 source.t39 source.n19 167.117
R170 source.t19 source.n27 167.117
R171 source.t4 source.n45 167.117
R172 source.n9 source.n8 84.1169
R173 source.n11 source.n10 84.1169
R174 source.n13 source.n12 84.1169
R175 source.n15 source.n14 84.1169
R176 source.n17 source.n16 84.1169
R177 source.n35 source.n34 84.1169
R178 source.n37 source.n36 84.1169
R179 source.n39 source.n38 84.1169
R180 source.n41 source.n40 84.1169
R181 source.n43 source.n42 84.1169
R182 source.n95 source.n94 84.1168
R183 source.n93 source.n92 84.1168
R184 source.n91 source.n90 84.1168
R185 source.n89 source.n88 84.1168
R186 source.n87 source.n86 84.1168
R187 source.n69 source.n68 84.1168
R188 source.n67 source.n66 84.1168
R189 source.n65 source.n64 84.1168
R190 source.n63 source.n62 84.1168
R191 source.n61 source.n60 84.1168
R192 source.n98 source.t8 52.3082
R193 source.n80 source.t1 52.3082
R194 source.n72 source.t38 52.3082
R195 source.n54 source.t24 52.3082
R196 source.n2 source.t37 52.3082
R197 source.n20 source.t39 52.3082
R198 source.n28 source.t19 52.3082
R199 source.n46 source.t4 52.3082
R200 source.n103 source.n102 31.4096
R201 source.n85 source.n84 31.4096
R202 source.n77 source.n76 31.4096
R203 source.n59 source.n58 31.4096
R204 source.n7 source.n6 31.4096
R205 source.n25 source.n24 31.4096
R206 source.n33 source.n32 31.4096
R207 source.n51 source.n50 31.4096
R208 source.n59 source.n51 14.5999
R209 source.n94 source.t10 9.9005
R210 source.n94 source.t3 9.9005
R211 source.n92 source.t15 9.9005
R212 source.n92 source.t12 9.9005
R213 source.n90 source.t47 9.9005
R214 source.n90 source.t46 9.9005
R215 source.n88 source.t16 9.9005
R216 source.n88 source.t18 9.9005
R217 source.n86 source.t5 9.9005
R218 source.n86 source.t20 9.9005
R219 source.n68 source.t29 9.9005
R220 source.n68 source.t42 9.9005
R221 source.n66 source.t40 9.9005
R222 source.n66 source.t27 9.9005
R223 source.n64 source.t43 9.9005
R224 source.n64 source.t34 9.9005
R225 source.n62 source.t28 9.9005
R226 source.n62 source.t45 9.9005
R227 source.n60 source.t44 9.9005
R228 source.n60 source.t32 9.9005
R229 source.n8 source.t33 9.9005
R230 source.n8 source.t36 9.9005
R231 source.n10 source.t41 9.9005
R232 source.n10 source.t25 9.9005
R233 source.n12 source.t23 9.9005
R234 source.n12 source.t31 9.9005
R235 source.n14 source.t30 9.9005
R236 source.n14 source.t26 9.9005
R237 source.n16 source.t22 9.9005
R238 source.n16 source.t35 9.9005
R239 source.n34 source.t14 9.9005
R240 source.n34 source.t9 9.9005
R241 source.n36 source.t11 9.9005
R242 source.n36 source.t21 9.9005
R243 source.n38 source.t6 9.9005
R244 source.n38 source.t17 9.9005
R245 source.n40 source.t2 9.9005
R246 source.n40 source.t0 9.9005
R247 source.n42 source.t7 9.9005
R248 source.n42 source.t13 9.9005
R249 source.n99 source.n97 9.71174
R250 source.n81 source.n79 9.71174
R251 source.n73 source.n71 9.71174
R252 source.n55 source.n53 9.71174
R253 source.n3 source.n1 9.71174
R254 source.n21 source.n19 9.71174
R255 source.n29 source.n27 9.71174
R256 source.n47 source.n45 9.71174
R257 source.n102 source.n101 9.45567
R258 source.n84 source.n83 9.45567
R259 source.n76 source.n75 9.45567
R260 source.n58 source.n57 9.45567
R261 source.n6 source.n5 9.45567
R262 source.n24 source.n23 9.45567
R263 source.n32 source.n31 9.45567
R264 source.n50 source.n49 9.45567
R265 source.n101 source.n100 9.3005
R266 source.n83 source.n82 9.3005
R267 source.n75 source.n74 9.3005
R268 source.n57 source.n56 9.3005
R269 source.n5 source.n4 9.3005
R270 source.n23 source.n22 9.3005
R271 source.n31 source.n30 9.3005
R272 source.n49 source.n48 9.3005
R273 source.n104 source.n7 8.893
R274 source.n102 source.n96 8.14595
R275 source.n84 source.n78 8.14595
R276 source.n76 source.n70 8.14595
R277 source.n58 source.n52 8.14595
R278 source.n6 source.n0 8.14595
R279 source.n24 source.n18 8.14595
R280 source.n32 source.n26 8.14595
R281 source.n50 source.n44 8.14595
R282 source.n100 source.n99 7.3702
R283 source.n82 source.n81 7.3702
R284 source.n74 source.n73 7.3702
R285 source.n56 source.n55 7.3702
R286 source.n4 source.n3 7.3702
R287 source.n22 source.n21 7.3702
R288 source.n30 source.n29 7.3702
R289 source.n48 source.n47 7.3702
R290 source.n100 source.n96 5.81868
R291 source.n82 source.n78 5.81868
R292 source.n74 source.n70 5.81868
R293 source.n56 source.n52 5.81868
R294 source.n4 source.n0 5.81868
R295 source.n22 source.n18 5.81868
R296 source.n30 source.n26 5.81868
R297 source.n48 source.n44 5.81868
R298 source.n104 source.n103 5.7074
R299 source.n101 source.n97 3.44771
R300 source.n83 source.n79 3.44771
R301 source.n75 source.n71 3.44771
R302 source.n57 source.n53 3.44771
R303 source.n5 source.n1 3.44771
R304 source.n23 source.n19 3.44771
R305 source.n31 source.n27 3.44771
R306 source.n49 source.n45 3.44771
R307 source.n51 source.n43 0.888431
R308 source.n43 source.n41 0.888431
R309 source.n41 source.n39 0.888431
R310 source.n39 source.n37 0.888431
R311 source.n37 source.n35 0.888431
R312 source.n35 source.n33 0.888431
R313 source.n25 source.n17 0.888431
R314 source.n17 source.n15 0.888431
R315 source.n15 source.n13 0.888431
R316 source.n13 source.n11 0.888431
R317 source.n11 source.n9 0.888431
R318 source.n9 source.n7 0.888431
R319 source.n61 source.n59 0.888431
R320 source.n63 source.n61 0.888431
R321 source.n65 source.n63 0.888431
R322 source.n67 source.n65 0.888431
R323 source.n69 source.n67 0.888431
R324 source.n77 source.n69 0.888431
R325 source.n87 source.n85 0.888431
R326 source.n89 source.n87 0.888431
R327 source.n91 source.n89 0.888431
R328 source.n93 source.n91 0.888431
R329 source.n95 source.n93 0.888431
R330 source.n103 source.n95 0.888431
R331 source.n33 source.n25 0.470328
R332 source.n85 source.n77 0.470328
R333 source source.n104 0.188
R334 drain_left.n13 drain_left.n11 101.683
R335 drain_left.n7 drain_left.n5 101.683
R336 drain_left.n2 drain_left.n0 101.683
R337 drain_left.n21 drain_left.n20 100.796
R338 drain_left.n19 drain_left.n18 100.796
R339 drain_left.n17 drain_left.n16 100.796
R340 drain_left.n15 drain_left.n14 100.796
R341 drain_left.n13 drain_left.n12 100.796
R342 drain_left.n7 drain_left.n6 100.796
R343 drain_left.n9 drain_left.n8 100.796
R344 drain_left.n4 drain_left.n3 100.796
R345 drain_left.n2 drain_left.n1 100.796
R346 drain_left drain_left.n10 28.2267
R347 drain_left.n5 drain_left.t2 9.9005
R348 drain_left.n5 drain_left.t1 9.9005
R349 drain_left.n6 drain_left.t11 9.9005
R350 drain_left.n6 drain_left.t18 9.9005
R351 drain_left.n8 drain_left.t7 9.9005
R352 drain_left.n8 drain_left.t12 9.9005
R353 drain_left.n3 drain_left.t3 9.9005
R354 drain_left.n3 drain_left.t9 9.9005
R355 drain_left.n1 drain_left.t22 9.9005
R356 drain_left.n1 drain_left.t23 9.9005
R357 drain_left.n0 drain_left.t14 9.9005
R358 drain_left.n0 drain_left.t13 9.9005
R359 drain_left.n20 drain_left.t6 9.9005
R360 drain_left.n20 drain_left.t21 9.9005
R361 drain_left.n18 drain_left.t0 9.9005
R362 drain_left.n18 drain_left.t17 9.9005
R363 drain_left.n16 drain_left.t20 9.9005
R364 drain_left.n16 drain_left.t10 9.9005
R365 drain_left.n14 drain_left.t16 9.9005
R366 drain_left.n14 drain_left.t5 9.9005
R367 drain_left.n12 drain_left.t19 9.9005
R368 drain_left.n12 drain_left.t8 9.9005
R369 drain_left.n11 drain_left.t15 9.9005
R370 drain_left.n11 drain_left.t4 9.9005
R371 drain_left drain_left.n21 6.54115
R372 drain_left.n9 drain_left.n7 0.888431
R373 drain_left.n4 drain_left.n2 0.888431
R374 drain_left.n15 drain_left.n13 0.888431
R375 drain_left.n17 drain_left.n15 0.888431
R376 drain_left.n19 drain_left.n17 0.888431
R377 drain_left.n21 drain_left.n19 0.888431
R378 drain_left.n10 drain_left.n9 0.389119
R379 drain_left.n10 drain_left.n4 0.389119
R380 minus.n41 minus.n40 161.3
R381 minus.n39 minus.n0 161.3
R382 minus.n38 minus.n37 161.3
R383 minus.n36 minus.n1 161.3
R384 minus.n35 minus.n34 161.3
R385 minus.n33 minus.n2 161.3
R386 minus.n32 minus.n31 161.3
R387 minus.n30 minus.n3 161.3
R388 minus.n29 minus.n28 161.3
R389 minus.n27 minus.n4 161.3
R390 minus.n26 minus.n25 161.3
R391 minus.n24 minus.n5 161.3
R392 minus.n23 minus.n22 161.3
R393 minus.n21 minus.n6 161.3
R394 minus.n20 minus.n19 161.3
R395 minus.n18 minus.n7 161.3
R396 minus.n17 minus.n16 161.3
R397 minus.n15 minus.n8 161.3
R398 minus.n14 minus.n13 161.3
R399 minus.n12 minus.n9 161.3
R400 minus.n83 minus.n82 161.3
R401 minus.n81 minus.n42 161.3
R402 minus.n80 minus.n79 161.3
R403 minus.n78 minus.n43 161.3
R404 minus.n77 minus.n76 161.3
R405 minus.n75 minus.n44 161.3
R406 minus.n74 minus.n73 161.3
R407 minus.n72 minus.n45 161.3
R408 minus.n71 minus.n70 161.3
R409 minus.n69 minus.n46 161.3
R410 minus.n68 minus.n67 161.3
R411 minus.n66 minus.n47 161.3
R412 minus.n65 minus.n64 161.3
R413 minus.n63 minus.n48 161.3
R414 minus.n62 minus.n61 161.3
R415 minus.n60 minus.n49 161.3
R416 minus.n59 minus.n58 161.3
R417 minus.n57 minus.n50 161.3
R418 minus.n56 minus.n55 161.3
R419 minus.n54 minus.n51 161.3
R420 minus.n11 minus.t13 151.334
R421 minus.n53 minus.t14 151.334
R422 minus.n10 minus.t0 124.977
R423 minus.n14 minus.t11 124.977
R424 minus.n16 minus.t22 124.977
R425 minus.n20 minus.t10 124.977
R426 minus.n22 minus.t23 124.977
R427 minus.n26 minus.t9 124.977
R428 minus.n28 minus.t18 124.977
R429 minus.n32 minus.t6 124.977
R430 minus.n34 minus.t16 124.977
R431 minus.n38 minus.t5 124.977
R432 minus.n40 minus.t15 124.977
R433 minus.n52 minus.t12 124.977
R434 minus.n56 minus.t19 124.977
R435 minus.n58 minus.t17 124.977
R436 minus.n62 minus.t21 124.977
R437 minus.n64 minus.t3 124.977
R438 minus.n68 minus.t2 124.977
R439 minus.n70 minus.t8 124.977
R440 minus.n74 minus.t7 124.977
R441 minus.n76 minus.t20 124.977
R442 minus.n80 minus.t4 124.977
R443 minus.n82 minus.t1 124.977
R444 minus.n40 minus.n39 46.0096
R445 minus.n82 minus.n81 46.0096
R446 minus.n12 minus.n11 45.0871
R447 minus.n54 minus.n53 45.0871
R448 minus.n10 minus.n9 41.6278
R449 minus.n38 minus.n1 41.6278
R450 minus.n52 minus.n51 41.6278
R451 minus.n80 minus.n43 41.6278
R452 minus.n15 minus.n14 37.246
R453 minus.n34 minus.n33 37.246
R454 minus.n57 minus.n56 37.246
R455 minus.n76 minus.n75 37.246
R456 minus.n84 minus.n41 34.58
R457 minus.n16 minus.n7 32.8641
R458 minus.n32 minus.n3 32.8641
R459 minus.n58 minus.n49 32.8641
R460 minus.n74 minus.n45 32.8641
R461 minus.n21 minus.n20 28.4823
R462 minus.n28 minus.n27 28.4823
R463 minus.n63 minus.n62 28.4823
R464 minus.n70 minus.n69 28.4823
R465 minus.n26 minus.n5 24.1005
R466 minus.n22 minus.n5 24.1005
R467 minus.n64 minus.n47 24.1005
R468 minus.n68 minus.n47 24.1005
R469 minus.n22 minus.n21 19.7187
R470 minus.n27 minus.n26 19.7187
R471 minus.n64 minus.n63 19.7187
R472 minus.n69 minus.n68 19.7187
R473 minus.n20 minus.n7 15.3369
R474 minus.n28 minus.n3 15.3369
R475 minus.n62 minus.n49 15.3369
R476 minus.n70 minus.n45 15.3369
R477 minus.n11 minus.n10 14.1472
R478 minus.n53 minus.n52 14.1472
R479 minus.n16 minus.n15 10.955
R480 minus.n33 minus.n32 10.955
R481 minus.n58 minus.n57 10.955
R482 minus.n75 minus.n74 10.955
R483 minus.n84 minus.n83 6.67853
R484 minus.n14 minus.n9 6.57323
R485 minus.n34 minus.n1 6.57323
R486 minus.n56 minus.n51 6.57323
R487 minus.n76 minus.n43 6.57323
R488 minus.n39 minus.n38 2.19141
R489 minus.n81 minus.n80 2.19141
R490 minus.n41 minus.n0 0.189894
R491 minus.n37 minus.n0 0.189894
R492 minus.n37 minus.n36 0.189894
R493 minus.n36 minus.n35 0.189894
R494 minus.n35 minus.n2 0.189894
R495 minus.n31 minus.n2 0.189894
R496 minus.n31 minus.n30 0.189894
R497 minus.n30 minus.n29 0.189894
R498 minus.n29 minus.n4 0.189894
R499 minus.n25 minus.n4 0.189894
R500 minus.n25 minus.n24 0.189894
R501 minus.n24 minus.n23 0.189894
R502 minus.n23 minus.n6 0.189894
R503 minus.n19 minus.n6 0.189894
R504 minus.n19 minus.n18 0.189894
R505 minus.n18 minus.n17 0.189894
R506 minus.n17 minus.n8 0.189894
R507 minus.n13 minus.n8 0.189894
R508 minus.n13 minus.n12 0.189894
R509 minus.n55 minus.n54 0.189894
R510 minus.n55 minus.n50 0.189894
R511 minus.n59 minus.n50 0.189894
R512 minus.n60 minus.n59 0.189894
R513 minus.n61 minus.n60 0.189894
R514 minus.n61 minus.n48 0.189894
R515 minus.n65 minus.n48 0.189894
R516 minus.n66 minus.n65 0.189894
R517 minus.n67 minus.n66 0.189894
R518 minus.n67 minus.n46 0.189894
R519 minus.n71 minus.n46 0.189894
R520 minus.n72 minus.n71 0.189894
R521 minus.n73 minus.n72 0.189894
R522 minus.n73 minus.n44 0.189894
R523 minus.n77 minus.n44 0.189894
R524 minus.n78 minus.n77 0.189894
R525 minus.n79 minus.n78 0.189894
R526 minus.n79 minus.n42 0.189894
R527 minus.n83 minus.n42 0.189894
R528 minus minus.n84 0.188
R529 drain_right.n13 drain_right.n11 101.683
R530 drain_right.n7 drain_right.n5 101.683
R531 drain_right.n2 drain_right.n0 101.683
R532 drain_right.n13 drain_right.n12 100.796
R533 drain_right.n15 drain_right.n14 100.796
R534 drain_right.n17 drain_right.n16 100.796
R535 drain_right.n19 drain_right.n18 100.796
R536 drain_right.n21 drain_right.n20 100.796
R537 drain_right.n7 drain_right.n6 100.796
R538 drain_right.n9 drain_right.n8 100.796
R539 drain_right.n4 drain_right.n3 100.796
R540 drain_right.n2 drain_right.n1 100.796
R541 drain_right drain_right.n10 27.6734
R542 drain_right.n5 drain_right.t19 9.9005
R543 drain_right.n5 drain_right.t22 9.9005
R544 drain_right.n6 drain_right.t16 9.9005
R545 drain_right.n6 drain_right.t3 9.9005
R546 drain_right.n8 drain_right.t21 9.9005
R547 drain_right.n8 drain_right.t15 9.9005
R548 drain_right.n3 drain_right.t2 9.9005
R549 drain_right.n3 drain_right.t20 9.9005
R550 drain_right.n1 drain_right.t4 9.9005
R551 drain_right.n1 drain_right.t6 9.9005
R552 drain_right.n0 drain_right.t9 9.9005
R553 drain_right.n0 drain_right.t11 9.9005
R554 drain_right.n11 drain_right.t23 9.9005
R555 drain_right.n11 drain_right.t10 9.9005
R556 drain_right.n12 drain_right.t1 9.9005
R557 drain_right.n12 drain_right.t12 9.9005
R558 drain_right.n14 drain_right.t0 9.9005
R559 drain_right.n14 drain_right.t13 9.9005
R560 drain_right.n16 drain_right.t5 9.9005
R561 drain_right.n16 drain_right.t14 9.9005
R562 drain_right.n18 drain_right.t7 9.9005
R563 drain_right.n18 drain_right.t17 9.9005
R564 drain_right.n20 drain_right.t8 9.9005
R565 drain_right.n20 drain_right.t18 9.9005
R566 drain_right drain_right.n21 6.54115
R567 drain_right.n9 drain_right.n7 0.888431
R568 drain_right.n4 drain_right.n2 0.888431
R569 drain_right.n21 drain_right.n19 0.888431
R570 drain_right.n19 drain_right.n17 0.888431
R571 drain_right.n17 drain_right.n15 0.888431
R572 drain_right.n15 drain_right.n13 0.888431
R573 drain_right.n10 drain_right.n9 0.389119
R574 drain_right.n10 drain_right.n4 0.389119
C0 source drain_left 8.688981f
C1 minus plus 5.53723f
C2 minus drain_left 0.180579f
C3 drain_left plus 3.48836f
C4 source drain_right 8.69155f
C5 drain_right minus 3.14809f
C6 source minus 4.03609f
C7 drain_right plus 0.505789f
C8 source plus 4.05005f
C9 drain_right drain_left 1.87044f
C10 drain_right a_n3394_n1288# 5.96745f
C11 drain_left a_n3394_n1288# 6.47274f
C12 source a_n3394_n1288# 3.664865f
C13 minus a_n3394_n1288# 12.890564f
C14 plus a_n3394_n1288# 14.349219f
C15 drain_right.t9 a_n3394_n1288# 0.042534f
C16 drain_right.t11 a_n3394_n1288# 0.042534f
C17 drain_right.n0 a_n3394_n1288# 0.270447f
C18 drain_right.t4 a_n3394_n1288# 0.042534f
C19 drain_right.t6 a_n3394_n1288# 0.042534f
C20 drain_right.n1 a_n3394_n1288# 0.267209f
C21 drain_right.n2 a_n3394_n1288# 0.727563f
C22 drain_right.t2 a_n3394_n1288# 0.042534f
C23 drain_right.t20 a_n3394_n1288# 0.042534f
C24 drain_right.n3 a_n3394_n1288# 0.267209f
C25 drain_right.n4 a_n3394_n1288# 0.318287f
C26 drain_right.t19 a_n3394_n1288# 0.042534f
C27 drain_right.t22 a_n3394_n1288# 0.042534f
C28 drain_right.n5 a_n3394_n1288# 0.270447f
C29 drain_right.t16 a_n3394_n1288# 0.042534f
C30 drain_right.t3 a_n3394_n1288# 0.042534f
C31 drain_right.n6 a_n3394_n1288# 0.267209f
C32 drain_right.n7 a_n3394_n1288# 0.727563f
C33 drain_right.t21 a_n3394_n1288# 0.042534f
C34 drain_right.t15 a_n3394_n1288# 0.042534f
C35 drain_right.n8 a_n3394_n1288# 0.267209f
C36 drain_right.n9 a_n3394_n1288# 0.318287f
C37 drain_right.n10 a_n3394_n1288# 1.15499f
C38 drain_right.t23 a_n3394_n1288# 0.042534f
C39 drain_right.t10 a_n3394_n1288# 0.042534f
C40 drain_right.n11 a_n3394_n1288# 0.270448f
C41 drain_right.t1 a_n3394_n1288# 0.042534f
C42 drain_right.t12 a_n3394_n1288# 0.042534f
C43 drain_right.n12 a_n3394_n1288# 0.26721f
C44 drain_right.n13 a_n3394_n1288# 0.727561f
C45 drain_right.t0 a_n3394_n1288# 0.042534f
C46 drain_right.t13 a_n3394_n1288# 0.042534f
C47 drain_right.n14 a_n3394_n1288# 0.26721f
C48 drain_right.n15 a_n3394_n1288# 0.35998f
C49 drain_right.t5 a_n3394_n1288# 0.042534f
C50 drain_right.t14 a_n3394_n1288# 0.042534f
C51 drain_right.n16 a_n3394_n1288# 0.26721f
C52 drain_right.n17 a_n3394_n1288# 0.35998f
C53 drain_right.t7 a_n3394_n1288# 0.042534f
C54 drain_right.t17 a_n3394_n1288# 0.042534f
C55 drain_right.n18 a_n3394_n1288# 0.26721f
C56 drain_right.n19 a_n3394_n1288# 0.35998f
C57 drain_right.t8 a_n3394_n1288# 0.042534f
C58 drain_right.t18 a_n3394_n1288# 0.042534f
C59 drain_right.n20 a_n3394_n1288# 0.26721f
C60 drain_right.n21 a_n3394_n1288# 0.598019f
C61 minus.n0 a_n3394_n1288# 0.041062f
C62 minus.n1 a_n3394_n1288# 0.009318f
C63 minus.t5 a_n3394_n1288# 0.17802f
C64 minus.n2 a_n3394_n1288# 0.041062f
C65 minus.n3 a_n3394_n1288# 0.009318f
C66 minus.t6 a_n3394_n1288# 0.17802f
C67 minus.n4 a_n3394_n1288# 0.041062f
C68 minus.n5 a_n3394_n1288# 0.009318f
C69 minus.t9 a_n3394_n1288# 0.17802f
C70 minus.n6 a_n3394_n1288# 0.041062f
C71 minus.n7 a_n3394_n1288# 0.009318f
C72 minus.t10 a_n3394_n1288# 0.17802f
C73 minus.n8 a_n3394_n1288# 0.041062f
C74 minus.n9 a_n3394_n1288# 0.009318f
C75 minus.t11 a_n3394_n1288# 0.17802f
C76 minus.t13 a_n3394_n1288# 0.199699f
C77 minus.t0 a_n3394_n1288# 0.17802f
C78 minus.n10 a_n3394_n1288# 0.132151f
C79 minus.n11 a_n3394_n1288# 0.104255f
C80 minus.n12 a_n3394_n1288# 0.176773f
C81 minus.n13 a_n3394_n1288# 0.041062f
C82 minus.n14 a_n3394_n1288# 0.123748f
C83 minus.n15 a_n3394_n1288# 0.009318f
C84 minus.t22 a_n3394_n1288# 0.17802f
C85 minus.n16 a_n3394_n1288# 0.123748f
C86 minus.n17 a_n3394_n1288# 0.041062f
C87 minus.n18 a_n3394_n1288# 0.041062f
C88 minus.n19 a_n3394_n1288# 0.041062f
C89 minus.n20 a_n3394_n1288# 0.123748f
C90 minus.n21 a_n3394_n1288# 0.009318f
C91 minus.t23 a_n3394_n1288# 0.17802f
C92 minus.n22 a_n3394_n1288# 0.123748f
C93 minus.n23 a_n3394_n1288# 0.041062f
C94 minus.n24 a_n3394_n1288# 0.041062f
C95 minus.n25 a_n3394_n1288# 0.041062f
C96 minus.n26 a_n3394_n1288# 0.123748f
C97 minus.n27 a_n3394_n1288# 0.009318f
C98 minus.t18 a_n3394_n1288# 0.17802f
C99 minus.n28 a_n3394_n1288# 0.123748f
C100 minus.n29 a_n3394_n1288# 0.041062f
C101 minus.n30 a_n3394_n1288# 0.041062f
C102 minus.n31 a_n3394_n1288# 0.041062f
C103 minus.n32 a_n3394_n1288# 0.123748f
C104 minus.n33 a_n3394_n1288# 0.009318f
C105 minus.t16 a_n3394_n1288# 0.17802f
C106 minus.n34 a_n3394_n1288# 0.123748f
C107 minus.n35 a_n3394_n1288# 0.041062f
C108 minus.n36 a_n3394_n1288# 0.041062f
C109 minus.n37 a_n3394_n1288# 0.041062f
C110 minus.n38 a_n3394_n1288# 0.123748f
C111 minus.n39 a_n3394_n1288# 0.009318f
C112 minus.t15 a_n3394_n1288# 0.17802f
C113 minus.n40 a_n3394_n1288# 0.124128f
C114 minus.n41 a_n3394_n1288# 1.35624f
C115 minus.n42 a_n3394_n1288# 0.041062f
C116 minus.n43 a_n3394_n1288# 0.009318f
C117 minus.n44 a_n3394_n1288# 0.041062f
C118 minus.n45 a_n3394_n1288# 0.009318f
C119 minus.n46 a_n3394_n1288# 0.041062f
C120 minus.n47 a_n3394_n1288# 0.009318f
C121 minus.n48 a_n3394_n1288# 0.041062f
C122 minus.n49 a_n3394_n1288# 0.009318f
C123 minus.n50 a_n3394_n1288# 0.041062f
C124 minus.n51 a_n3394_n1288# 0.009318f
C125 minus.t14 a_n3394_n1288# 0.199699f
C126 minus.t12 a_n3394_n1288# 0.17802f
C127 minus.n52 a_n3394_n1288# 0.132151f
C128 minus.n53 a_n3394_n1288# 0.104255f
C129 minus.n54 a_n3394_n1288# 0.176773f
C130 minus.n55 a_n3394_n1288# 0.041062f
C131 minus.t19 a_n3394_n1288# 0.17802f
C132 minus.n56 a_n3394_n1288# 0.123748f
C133 minus.n57 a_n3394_n1288# 0.009318f
C134 minus.t17 a_n3394_n1288# 0.17802f
C135 minus.n58 a_n3394_n1288# 0.123748f
C136 minus.n59 a_n3394_n1288# 0.041062f
C137 minus.n60 a_n3394_n1288# 0.041062f
C138 minus.n61 a_n3394_n1288# 0.041062f
C139 minus.t21 a_n3394_n1288# 0.17802f
C140 minus.n62 a_n3394_n1288# 0.123748f
C141 minus.n63 a_n3394_n1288# 0.009318f
C142 minus.t3 a_n3394_n1288# 0.17802f
C143 minus.n64 a_n3394_n1288# 0.123748f
C144 minus.n65 a_n3394_n1288# 0.041062f
C145 minus.n66 a_n3394_n1288# 0.041062f
C146 minus.n67 a_n3394_n1288# 0.041062f
C147 minus.t2 a_n3394_n1288# 0.17802f
C148 minus.n68 a_n3394_n1288# 0.123748f
C149 minus.n69 a_n3394_n1288# 0.009318f
C150 minus.t8 a_n3394_n1288# 0.17802f
C151 minus.n70 a_n3394_n1288# 0.123748f
C152 minus.n71 a_n3394_n1288# 0.041062f
C153 minus.n72 a_n3394_n1288# 0.041062f
C154 minus.n73 a_n3394_n1288# 0.041062f
C155 minus.t7 a_n3394_n1288# 0.17802f
C156 minus.n74 a_n3394_n1288# 0.123748f
C157 minus.n75 a_n3394_n1288# 0.009318f
C158 minus.t20 a_n3394_n1288# 0.17802f
C159 minus.n76 a_n3394_n1288# 0.123748f
C160 minus.n77 a_n3394_n1288# 0.041062f
C161 minus.n78 a_n3394_n1288# 0.041062f
C162 minus.n79 a_n3394_n1288# 0.041062f
C163 minus.t4 a_n3394_n1288# 0.17802f
C164 minus.n80 a_n3394_n1288# 0.123748f
C165 minus.n81 a_n3394_n1288# 0.009318f
C166 minus.t1 a_n3394_n1288# 0.17802f
C167 minus.n82 a_n3394_n1288# 0.124128f
C168 minus.n83 a_n3394_n1288# 0.28558f
C169 minus.n84 a_n3394_n1288# 1.64872f
C170 drain_left.t14 a_n3394_n1288# 0.043586f
C171 drain_left.t13 a_n3394_n1288# 0.043586f
C172 drain_left.n0 a_n3394_n1288# 0.277142f
C173 drain_left.t22 a_n3394_n1288# 0.043586f
C174 drain_left.t23 a_n3394_n1288# 0.043586f
C175 drain_left.n1 a_n3394_n1288# 0.273824f
C176 drain_left.n2 a_n3394_n1288# 0.745574f
C177 drain_left.t3 a_n3394_n1288# 0.043586f
C178 drain_left.t9 a_n3394_n1288# 0.043586f
C179 drain_left.n3 a_n3394_n1288# 0.273824f
C180 drain_left.n4 a_n3394_n1288# 0.326167f
C181 drain_left.t2 a_n3394_n1288# 0.043586f
C182 drain_left.t1 a_n3394_n1288# 0.043586f
C183 drain_left.n5 a_n3394_n1288# 0.277142f
C184 drain_left.t11 a_n3394_n1288# 0.043586f
C185 drain_left.t18 a_n3394_n1288# 0.043586f
C186 drain_left.n6 a_n3394_n1288# 0.273824f
C187 drain_left.n7 a_n3394_n1288# 0.745574f
C188 drain_left.t7 a_n3394_n1288# 0.043586f
C189 drain_left.t12 a_n3394_n1288# 0.043586f
C190 drain_left.n8 a_n3394_n1288# 0.273824f
C191 drain_left.n9 a_n3394_n1288# 0.326167f
C192 drain_left.n10 a_n3394_n1288# 1.23684f
C193 drain_left.t15 a_n3394_n1288# 0.043586f
C194 drain_left.t4 a_n3394_n1288# 0.043586f
C195 drain_left.n11 a_n3394_n1288# 0.277144f
C196 drain_left.t19 a_n3394_n1288# 0.043586f
C197 drain_left.t8 a_n3394_n1288# 0.043586f
C198 drain_left.n12 a_n3394_n1288# 0.273825f
C199 drain_left.n13 a_n3394_n1288# 0.745572f
C200 drain_left.t16 a_n3394_n1288# 0.043586f
C201 drain_left.t5 a_n3394_n1288# 0.043586f
C202 drain_left.n14 a_n3394_n1288# 0.273825f
C203 drain_left.n15 a_n3394_n1288# 0.368891f
C204 drain_left.t20 a_n3394_n1288# 0.043586f
C205 drain_left.t10 a_n3394_n1288# 0.043586f
C206 drain_left.n16 a_n3394_n1288# 0.273825f
C207 drain_left.n17 a_n3394_n1288# 0.368891f
C208 drain_left.t0 a_n3394_n1288# 0.043586f
C209 drain_left.t17 a_n3394_n1288# 0.043586f
C210 drain_left.n18 a_n3394_n1288# 0.273825f
C211 drain_left.n19 a_n3394_n1288# 0.368891f
C212 drain_left.t6 a_n3394_n1288# 0.043586f
C213 drain_left.t21 a_n3394_n1288# 0.043586f
C214 drain_left.n20 a_n3394_n1288# 0.273825f
C215 drain_left.n21 a_n3394_n1288# 0.612823f
C216 source.n0 a_n3394_n1288# 0.047137f
C217 source.n1 a_n3394_n1288# 0.104297f
C218 source.t37 a_n3394_n1288# 0.07827f
C219 source.n2 a_n3394_n1288# 0.081627f
C220 source.n3 a_n3394_n1288# 0.026313f
C221 source.n4 a_n3394_n1288# 0.017354f
C222 source.n5 a_n3394_n1288# 0.229896f
C223 source.n6 a_n3394_n1288# 0.051673f
C224 source.n7 a_n3394_n1288# 0.551187f
C225 source.t33 a_n3394_n1288# 0.051042f
C226 source.t36 a_n3394_n1288# 0.051042f
C227 source.n8 a_n3394_n1288# 0.272868f
C228 source.n9 a_n3394_n1288# 0.435885f
C229 source.t41 a_n3394_n1288# 0.051042f
C230 source.t25 a_n3394_n1288# 0.051042f
C231 source.n10 a_n3394_n1288# 0.272868f
C232 source.n11 a_n3394_n1288# 0.435885f
C233 source.t23 a_n3394_n1288# 0.051042f
C234 source.t31 a_n3394_n1288# 0.051042f
C235 source.n12 a_n3394_n1288# 0.272868f
C236 source.n13 a_n3394_n1288# 0.435885f
C237 source.t30 a_n3394_n1288# 0.051042f
C238 source.t26 a_n3394_n1288# 0.051042f
C239 source.n14 a_n3394_n1288# 0.272868f
C240 source.n15 a_n3394_n1288# 0.435885f
C241 source.t22 a_n3394_n1288# 0.051042f
C242 source.t35 a_n3394_n1288# 0.051042f
C243 source.n16 a_n3394_n1288# 0.272868f
C244 source.n17 a_n3394_n1288# 0.435885f
C245 source.n18 a_n3394_n1288# 0.047137f
C246 source.n19 a_n3394_n1288# 0.104297f
C247 source.t39 a_n3394_n1288# 0.07827f
C248 source.n20 a_n3394_n1288# 0.081627f
C249 source.n21 a_n3394_n1288# 0.026313f
C250 source.n22 a_n3394_n1288# 0.017354f
C251 source.n23 a_n3394_n1288# 0.229896f
C252 source.n24 a_n3394_n1288# 0.051673f
C253 source.n25 a_n3394_n1288# 0.16788f
C254 source.n26 a_n3394_n1288# 0.047137f
C255 source.n27 a_n3394_n1288# 0.104297f
C256 source.t19 a_n3394_n1288# 0.07827f
C257 source.n28 a_n3394_n1288# 0.081627f
C258 source.n29 a_n3394_n1288# 0.026313f
C259 source.n30 a_n3394_n1288# 0.017354f
C260 source.n31 a_n3394_n1288# 0.229896f
C261 source.n32 a_n3394_n1288# 0.051673f
C262 source.n33 a_n3394_n1288# 0.16788f
C263 source.t14 a_n3394_n1288# 0.051042f
C264 source.t9 a_n3394_n1288# 0.051042f
C265 source.n34 a_n3394_n1288# 0.272868f
C266 source.n35 a_n3394_n1288# 0.435885f
C267 source.t11 a_n3394_n1288# 0.051042f
C268 source.t21 a_n3394_n1288# 0.051042f
C269 source.n36 a_n3394_n1288# 0.272868f
C270 source.n37 a_n3394_n1288# 0.435885f
C271 source.t6 a_n3394_n1288# 0.051042f
C272 source.t17 a_n3394_n1288# 0.051042f
C273 source.n38 a_n3394_n1288# 0.272868f
C274 source.n39 a_n3394_n1288# 0.435885f
C275 source.t2 a_n3394_n1288# 0.051042f
C276 source.t0 a_n3394_n1288# 0.051042f
C277 source.n40 a_n3394_n1288# 0.272868f
C278 source.n41 a_n3394_n1288# 0.435885f
C279 source.t7 a_n3394_n1288# 0.051042f
C280 source.t13 a_n3394_n1288# 0.051042f
C281 source.n42 a_n3394_n1288# 0.272868f
C282 source.n43 a_n3394_n1288# 0.435885f
C283 source.n44 a_n3394_n1288# 0.047137f
C284 source.n45 a_n3394_n1288# 0.104297f
C285 source.t4 a_n3394_n1288# 0.07827f
C286 source.n46 a_n3394_n1288# 0.081627f
C287 source.n47 a_n3394_n1288# 0.026313f
C288 source.n48 a_n3394_n1288# 0.017354f
C289 source.n49 a_n3394_n1288# 0.229896f
C290 source.n50 a_n3394_n1288# 0.051673f
C291 source.n51 a_n3394_n1288# 0.860469f
C292 source.n52 a_n3394_n1288# 0.047137f
C293 source.n53 a_n3394_n1288# 0.104297f
C294 source.t24 a_n3394_n1288# 0.07827f
C295 source.n54 a_n3394_n1288# 0.081627f
C296 source.n55 a_n3394_n1288# 0.026313f
C297 source.n56 a_n3394_n1288# 0.017354f
C298 source.n57 a_n3394_n1288# 0.229896f
C299 source.n58 a_n3394_n1288# 0.051673f
C300 source.n59 a_n3394_n1288# 0.860469f
C301 source.t44 a_n3394_n1288# 0.051042f
C302 source.t32 a_n3394_n1288# 0.051042f
C303 source.n60 a_n3394_n1288# 0.272866f
C304 source.n61 a_n3394_n1288# 0.435886f
C305 source.t28 a_n3394_n1288# 0.051042f
C306 source.t45 a_n3394_n1288# 0.051042f
C307 source.n62 a_n3394_n1288# 0.272866f
C308 source.n63 a_n3394_n1288# 0.435886f
C309 source.t43 a_n3394_n1288# 0.051042f
C310 source.t34 a_n3394_n1288# 0.051042f
C311 source.n64 a_n3394_n1288# 0.272866f
C312 source.n65 a_n3394_n1288# 0.435886f
C313 source.t40 a_n3394_n1288# 0.051042f
C314 source.t27 a_n3394_n1288# 0.051042f
C315 source.n66 a_n3394_n1288# 0.272866f
C316 source.n67 a_n3394_n1288# 0.435886f
C317 source.t29 a_n3394_n1288# 0.051042f
C318 source.t42 a_n3394_n1288# 0.051042f
C319 source.n68 a_n3394_n1288# 0.272866f
C320 source.n69 a_n3394_n1288# 0.435886f
C321 source.n70 a_n3394_n1288# 0.047137f
C322 source.n71 a_n3394_n1288# 0.104297f
C323 source.t38 a_n3394_n1288# 0.07827f
C324 source.n72 a_n3394_n1288# 0.081627f
C325 source.n73 a_n3394_n1288# 0.026313f
C326 source.n74 a_n3394_n1288# 0.017354f
C327 source.n75 a_n3394_n1288# 0.229896f
C328 source.n76 a_n3394_n1288# 0.051673f
C329 source.n77 a_n3394_n1288# 0.16788f
C330 source.n78 a_n3394_n1288# 0.047137f
C331 source.n79 a_n3394_n1288# 0.104297f
C332 source.t1 a_n3394_n1288# 0.07827f
C333 source.n80 a_n3394_n1288# 0.081627f
C334 source.n81 a_n3394_n1288# 0.026313f
C335 source.n82 a_n3394_n1288# 0.017354f
C336 source.n83 a_n3394_n1288# 0.229896f
C337 source.n84 a_n3394_n1288# 0.051673f
C338 source.n85 a_n3394_n1288# 0.16788f
C339 source.t5 a_n3394_n1288# 0.051042f
C340 source.t20 a_n3394_n1288# 0.051042f
C341 source.n86 a_n3394_n1288# 0.272866f
C342 source.n87 a_n3394_n1288# 0.435886f
C343 source.t16 a_n3394_n1288# 0.051042f
C344 source.t18 a_n3394_n1288# 0.051042f
C345 source.n88 a_n3394_n1288# 0.272866f
C346 source.n89 a_n3394_n1288# 0.435886f
C347 source.t47 a_n3394_n1288# 0.051042f
C348 source.t46 a_n3394_n1288# 0.051042f
C349 source.n90 a_n3394_n1288# 0.272866f
C350 source.n91 a_n3394_n1288# 0.435886f
C351 source.t15 a_n3394_n1288# 0.051042f
C352 source.t12 a_n3394_n1288# 0.051042f
C353 source.n92 a_n3394_n1288# 0.272866f
C354 source.n93 a_n3394_n1288# 0.435886f
C355 source.t10 a_n3394_n1288# 0.051042f
C356 source.t3 a_n3394_n1288# 0.051042f
C357 source.n94 a_n3394_n1288# 0.272866f
C358 source.n95 a_n3394_n1288# 0.435886f
C359 source.n96 a_n3394_n1288# 0.047137f
C360 source.n97 a_n3394_n1288# 0.104297f
C361 source.t8 a_n3394_n1288# 0.07827f
C362 source.n98 a_n3394_n1288# 0.081627f
C363 source.n99 a_n3394_n1288# 0.026313f
C364 source.n100 a_n3394_n1288# 0.017354f
C365 source.n101 a_n3394_n1288# 0.229896f
C366 source.n102 a_n3394_n1288# 0.051673f
C367 source.n103 a_n3394_n1288# 0.378544f
C368 source.n104 a_n3394_n1288# 0.814179f
C369 plus.n0 a_n3394_n1288# 0.042974f
C370 plus.t2 a_n3394_n1288# 0.186312f
C371 plus.t17 a_n3394_n1288# 0.186312f
C372 plus.n1 a_n3394_n1288# 0.042974f
C373 plus.t6 a_n3394_n1288# 0.186312f
C374 plus.n2 a_n3394_n1288# 0.129512f
C375 plus.n3 a_n3394_n1288# 0.042974f
C376 plus.t23 a_n3394_n1288# 0.186312f
C377 plus.t13 a_n3394_n1288# 0.186312f
C378 plus.n4 a_n3394_n1288# 0.129512f
C379 plus.n5 a_n3394_n1288# 0.042974f
C380 plus.t3 a_n3394_n1288# 0.186312f
C381 plus.t18 a_n3394_n1288# 0.186312f
C382 plus.n6 a_n3394_n1288# 0.129512f
C383 plus.n7 a_n3394_n1288# 0.042974f
C384 plus.t7 a_n3394_n1288# 0.186312f
C385 plus.t15 a_n3394_n1288# 0.186312f
C386 plus.n8 a_n3394_n1288# 0.129512f
C387 plus.n9 a_n3394_n1288# 0.042974f
C388 plus.t4 a_n3394_n1288# 0.186312f
C389 plus.t19 a_n3394_n1288# 0.186312f
C390 plus.n10 a_n3394_n1288# 0.138306f
C391 plus.t8 a_n3394_n1288# 0.209001f
C392 plus.n11 a_n3394_n1288# 0.109111f
C393 plus.n12 a_n3394_n1288# 0.185007f
C394 plus.n13 a_n3394_n1288# 0.009752f
C395 plus.n14 a_n3394_n1288# 0.129512f
C396 plus.n15 a_n3394_n1288# 0.009752f
C397 plus.n16 a_n3394_n1288# 0.042974f
C398 plus.n17 a_n3394_n1288# 0.042974f
C399 plus.n18 a_n3394_n1288# 0.042974f
C400 plus.n19 a_n3394_n1288# 0.009752f
C401 plus.n20 a_n3394_n1288# 0.129512f
C402 plus.n21 a_n3394_n1288# 0.009752f
C403 plus.n22 a_n3394_n1288# 0.042974f
C404 plus.n23 a_n3394_n1288# 0.042974f
C405 plus.n24 a_n3394_n1288# 0.042974f
C406 plus.n25 a_n3394_n1288# 0.009752f
C407 plus.n26 a_n3394_n1288# 0.129512f
C408 plus.n27 a_n3394_n1288# 0.009752f
C409 plus.n28 a_n3394_n1288# 0.042974f
C410 plus.n29 a_n3394_n1288# 0.042974f
C411 plus.n30 a_n3394_n1288# 0.042974f
C412 plus.n31 a_n3394_n1288# 0.009752f
C413 plus.n32 a_n3394_n1288# 0.129512f
C414 plus.n33 a_n3394_n1288# 0.009752f
C415 plus.n34 a_n3394_n1288# 0.042974f
C416 plus.n35 a_n3394_n1288# 0.042974f
C417 plus.n36 a_n3394_n1288# 0.042974f
C418 plus.n37 a_n3394_n1288# 0.009752f
C419 plus.n38 a_n3394_n1288# 0.129512f
C420 plus.n39 a_n3394_n1288# 0.009752f
C421 plus.n40 a_n3394_n1288# 0.129909f
C422 plus.n41 a_n3394_n1288# 0.32613f
C423 plus.n42 a_n3394_n1288# 0.042974f
C424 plus.t9 a_n3394_n1288# 0.186312f
C425 plus.n43 a_n3394_n1288# 0.042974f
C426 plus.t10 a_n3394_n1288# 0.186312f
C427 plus.t1 a_n3394_n1288# 0.186312f
C428 plus.n44 a_n3394_n1288# 0.129512f
C429 plus.n45 a_n3394_n1288# 0.042974f
C430 plus.t0 a_n3394_n1288# 0.186312f
C431 plus.t20 a_n3394_n1288# 0.186312f
C432 plus.n46 a_n3394_n1288# 0.129512f
C433 plus.n47 a_n3394_n1288# 0.042974f
C434 plus.t14 a_n3394_n1288# 0.186312f
C435 plus.t16 a_n3394_n1288# 0.186312f
C436 plus.n48 a_n3394_n1288# 0.129512f
C437 plus.n49 a_n3394_n1288# 0.042974f
C438 plus.t11 a_n3394_n1288# 0.186312f
C439 plus.t12 a_n3394_n1288# 0.186312f
C440 plus.n50 a_n3394_n1288# 0.129512f
C441 plus.n51 a_n3394_n1288# 0.042974f
C442 plus.t5 a_n3394_n1288# 0.186312f
C443 plus.t21 a_n3394_n1288# 0.186312f
C444 plus.n52 a_n3394_n1288# 0.138306f
C445 plus.t22 a_n3394_n1288# 0.209001f
C446 plus.n53 a_n3394_n1288# 0.109111f
C447 plus.n54 a_n3394_n1288# 0.185007f
C448 plus.n55 a_n3394_n1288# 0.009752f
C449 plus.n56 a_n3394_n1288# 0.129512f
C450 plus.n57 a_n3394_n1288# 0.009752f
C451 plus.n58 a_n3394_n1288# 0.042974f
C452 plus.n59 a_n3394_n1288# 0.042974f
C453 plus.n60 a_n3394_n1288# 0.042974f
C454 plus.n61 a_n3394_n1288# 0.009752f
C455 plus.n62 a_n3394_n1288# 0.129512f
C456 plus.n63 a_n3394_n1288# 0.009752f
C457 plus.n64 a_n3394_n1288# 0.042974f
C458 plus.n65 a_n3394_n1288# 0.042974f
C459 plus.n66 a_n3394_n1288# 0.042974f
C460 plus.n67 a_n3394_n1288# 0.009752f
C461 plus.n68 a_n3394_n1288# 0.129512f
C462 plus.n69 a_n3394_n1288# 0.009752f
C463 plus.n70 a_n3394_n1288# 0.042974f
C464 plus.n71 a_n3394_n1288# 0.042974f
C465 plus.n72 a_n3394_n1288# 0.042974f
C466 plus.n73 a_n3394_n1288# 0.009752f
C467 plus.n74 a_n3394_n1288# 0.129512f
C468 plus.n75 a_n3394_n1288# 0.009752f
C469 plus.n76 a_n3394_n1288# 0.042974f
C470 plus.n77 a_n3394_n1288# 0.042974f
C471 plus.n78 a_n3394_n1288# 0.042974f
C472 plus.n79 a_n3394_n1288# 0.009752f
C473 plus.n80 a_n3394_n1288# 0.129512f
C474 plus.n81 a_n3394_n1288# 0.009752f
C475 plus.n82 a_n3394_n1288# 0.129909f
C476 plus.n83 a_n3394_n1288# 1.34907f
.ends

