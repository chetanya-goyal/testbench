* NGSPICE file created from diffpair706.ext - technology: sky130A

.subckt diffpair706 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t22 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X1 source.t7 plus.t0 drain_left.t13 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X2 a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.7
X3 source.t20 minus.t1 drain_right.t12 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X4 drain_left.t12 plus.t1 source.t0 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X5 drain_left.t11 plus.t2 source.t1 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X6 source.t18 minus.t2 drain_right.t11 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X7 drain_right.t10 minus.t3 source.t25 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X8 source.t2 plus.t3 drain_left.t10 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X9 drain_left.t9 plus.t4 source.t6 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X10 drain_left.t8 plus.t5 source.t9 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X11 drain_left.t7 plus.t6 source.t27 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X12 source.t15 minus.t4 drain_right.t9 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X13 drain_right.t8 minus.t5 source.t24 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X14 a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X15 drain_right.t7 minus.t6 source.t17 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X16 drain_right.t6 minus.t7 source.t16 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X17 drain_right.t5 minus.t8 source.t13 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X18 source.t5 plus.t7 drain_left.t6 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X19 source.t4 plus.t8 drain_left.t5 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X20 drain_left.t4 plus.t9 source.t11 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X21 source.t3 plus.t10 drain_left.t3 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X22 a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X23 drain_right.t4 minus.t9 source.t14 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X24 a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X25 source.t8 plus.t11 drain_left.t2 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X26 drain_left.t1 plus.t12 source.t10 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X27 source.t12 minus.t10 drain_right.t3 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X28 drain_right.t2 minus.t11 source.t23 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X29 source.t21 minus.t12 drain_right.t1 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X30 source.t19 minus.t13 drain_right.t0 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X31 drain_left.t0 plus.t13 source.t26 a_n2364_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
R0 minus.n5 minus.t9 940.679
R1 minus.n27 minus.t5 940.679
R2 minus.n6 minus.t2 916.833
R3 minus.n8 minus.t8 916.833
R4 minus.n12 minus.t12 916.833
R5 minus.n14 minus.t7 916.833
R6 minus.n18 minus.t13 916.833
R7 minus.n20 minus.t6 916.833
R8 minus.n28 minus.t4 916.833
R9 minus.n30 minus.t0 916.833
R10 minus.n34 minus.t1 916.833
R11 minus.n36 minus.t3 916.833
R12 minus.n40 minus.t10 916.833
R13 minus.n42 minus.t11 916.833
R14 minus.n21 minus.n20 161.3
R15 minus.n19 minus.n0 161.3
R16 minus.n18 minus.n17 161.3
R17 minus.n16 minus.n1 161.3
R18 minus.n15 minus.n14 161.3
R19 minus.n13 minus.n2 161.3
R20 minus.n12 minus.n11 161.3
R21 minus.n10 minus.n3 161.3
R22 minus.n9 minus.n8 161.3
R23 minus.n7 minus.n4 161.3
R24 minus.n43 minus.n42 161.3
R25 minus.n41 minus.n22 161.3
R26 minus.n40 minus.n39 161.3
R27 minus.n38 minus.n23 161.3
R28 minus.n37 minus.n36 161.3
R29 minus.n35 minus.n24 161.3
R30 minus.n34 minus.n33 161.3
R31 minus.n32 minus.n25 161.3
R32 minus.n31 minus.n30 161.3
R33 minus.n29 minus.n26 161.3
R34 minus.n44 minus.n21 48.0744
R35 minus.n5 minus.n4 44.9119
R36 minus.n27 minus.n26 44.9119
R37 minus.n20 minus.n19 35.055
R38 minus.n42 minus.n41 35.055
R39 minus.n7 minus.n6 30.6732
R40 minus.n18 minus.n1 30.6732
R41 minus.n29 minus.n28 30.6732
R42 minus.n40 minus.n23 30.6732
R43 minus.n8 minus.n3 26.2914
R44 minus.n14 minus.n13 26.2914
R45 minus.n30 minus.n25 26.2914
R46 minus.n36 minus.n35 26.2914
R47 minus.n12 minus.n3 21.9096
R48 minus.n13 minus.n12 21.9096
R49 minus.n34 minus.n25 21.9096
R50 minus.n35 minus.n34 21.9096
R51 minus.n6 minus.n5 17.739
R52 minus.n28 minus.n27 17.739
R53 minus.n8 minus.n7 17.5278
R54 minus.n14 minus.n1 17.5278
R55 minus.n30 minus.n29 17.5278
R56 minus.n36 minus.n23 17.5278
R57 minus.n19 minus.n18 13.146
R58 minus.n41 minus.n40 13.146
R59 minus.n44 minus.n43 6.65012
R60 minus.n21 minus.n0 0.189894
R61 minus.n17 minus.n0 0.189894
R62 minus.n17 minus.n16 0.189894
R63 minus.n16 minus.n15 0.189894
R64 minus.n15 minus.n2 0.189894
R65 minus.n11 minus.n2 0.189894
R66 minus.n11 minus.n10 0.189894
R67 minus.n10 minus.n9 0.189894
R68 minus.n9 minus.n4 0.189894
R69 minus.n31 minus.n26 0.189894
R70 minus.n32 minus.n31 0.189894
R71 minus.n33 minus.n32 0.189894
R72 minus.n33 minus.n24 0.189894
R73 minus.n37 minus.n24 0.189894
R74 minus.n38 minus.n37 0.189894
R75 minus.n39 minus.n38 0.189894
R76 minus.n39 minus.n22 0.189894
R77 minus.n43 minus.n22 0.189894
R78 minus minus.n44 0.188
R79 source.n578 source.n444 289.615
R80 source.n432 source.n298 289.615
R81 source.n134 source.n0 289.615
R82 source.n280 source.n146 289.615
R83 source.n488 source.n487 185
R84 source.n493 source.n492 185
R85 source.n495 source.n494 185
R86 source.n484 source.n483 185
R87 source.n501 source.n500 185
R88 source.n503 source.n502 185
R89 source.n480 source.n479 185
R90 source.n510 source.n509 185
R91 source.n511 source.n478 185
R92 source.n513 source.n512 185
R93 source.n476 source.n475 185
R94 source.n519 source.n518 185
R95 source.n521 source.n520 185
R96 source.n472 source.n471 185
R97 source.n527 source.n526 185
R98 source.n529 source.n528 185
R99 source.n468 source.n467 185
R100 source.n535 source.n534 185
R101 source.n537 source.n536 185
R102 source.n464 source.n463 185
R103 source.n543 source.n542 185
R104 source.n545 source.n544 185
R105 source.n460 source.n459 185
R106 source.n551 source.n550 185
R107 source.n554 source.n553 185
R108 source.n552 source.n456 185
R109 source.n559 source.n455 185
R110 source.n561 source.n560 185
R111 source.n563 source.n562 185
R112 source.n452 source.n451 185
R113 source.n569 source.n568 185
R114 source.n571 source.n570 185
R115 source.n448 source.n447 185
R116 source.n577 source.n576 185
R117 source.n579 source.n578 185
R118 source.n342 source.n341 185
R119 source.n347 source.n346 185
R120 source.n349 source.n348 185
R121 source.n338 source.n337 185
R122 source.n355 source.n354 185
R123 source.n357 source.n356 185
R124 source.n334 source.n333 185
R125 source.n364 source.n363 185
R126 source.n365 source.n332 185
R127 source.n367 source.n366 185
R128 source.n330 source.n329 185
R129 source.n373 source.n372 185
R130 source.n375 source.n374 185
R131 source.n326 source.n325 185
R132 source.n381 source.n380 185
R133 source.n383 source.n382 185
R134 source.n322 source.n321 185
R135 source.n389 source.n388 185
R136 source.n391 source.n390 185
R137 source.n318 source.n317 185
R138 source.n397 source.n396 185
R139 source.n399 source.n398 185
R140 source.n314 source.n313 185
R141 source.n405 source.n404 185
R142 source.n408 source.n407 185
R143 source.n406 source.n310 185
R144 source.n413 source.n309 185
R145 source.n415 source.n414 185
R146 source.n417 source.n416 185
R147 source.n306 source.n305 185
R148 source.n423 source.n422 185
R149 source.n425 source.n424 185
R150 source.n302 source.n301 185
R151 source.n431 source.n430 185
R152 source.n433 source.n432 185
R153 source.n135 source.n134 185
R154 source.n133 source.n132 185
R155 source.n4 source.n3 185
R156 source.n127 source.n126 185
R157 source.n125 source.n124 185
R158 source.n8 source.n7 185
R159 source.n119 source.n118 185
R160 source.n117 source.n116 185
R161 source.n115 source.n11 185
R162 source.n15 source.n12 185
R163 source.n110 source.n109 185
R164 source.n108 source.n107 185
R165 source.n17 source.n16 185
R166 source.n102 source.n101 185
R167 source.n100 source.n99 185
R168 source.n21 source.n20 185
R169 source.n94 source.n93 185
R170 source.n92 source.n91 185
R171 source.n25 source.n24 185
R172 source.n86 source.n85 185
R173 source.n84 source.n83 185
R174 source.n29 source.n28 185
R175 source.n78 source.n77 185
R176 source.n76 source.n75 185
R177 source.n33 source.n32 185
R178 source.n70 source.n69 185
R179 source.n68 source.n35 185
R180 source.n67 source.n66 185
R181 source.n38 source.n36 185
R182 source.n61 source.n60 185
R183 source.n59 source.n58 185
R184 source.n42 source.n41 185
R185 source.n53 source.n52 185
R186 source.n51 source.n50 185
R187 source.n46 source.n45 185
R188 source.n281 source.n280 185
R189 source.n279 source.n278 185
R190 source.n150 source.n149 185
R191 source.n273 source.n272 185
R192 source.n271 source.n270 185
R193 source.n154 source.n153 185
R194 source.n265 source.n264 185
R195 source.n263 source.n262 185
R196 source.n261 source.n157 185
R197 source.n161 source.n158 185
R198 source.n256 source.n255 185
R199 source.n254 source.n253 185
R200 source.n163 source.n162 185
R201 source.n248 source.n247 185
R202 source.n246 source.n245 185
R203 source.n167 source.n166 185
R204 source.n240 source.n239 185
R205 source.n238 source.n237 185
R206 source.n171 source.n170 185
R207 source.n232 source.n231 185
R208 source.n230 source.n229 185
R209 source.n175 source.n174 185
R210 source.n224 source.n223 185
R211 source.n222 source.n221 185
R212 source.n179 source.n178 185
R213 source.n216 source.n215 185
R214 source.n214 source.n181 185
R215 source.n213 source.n212 185
R216 source.n184 source.n182 185
R217 source.n207 source.n206 185
R218 source.n205 source.n204 185
R219 source.n188 source.n187 185
R220 source.n199 source.n198 185
R221 source.n197 source.n196 185
R222 source.n192 source.n191 185
R223 source.n489 source.t23 149.524
R224 source.n343 source.t26 149.524
R225 source.n47 source.t0 149.524
R226 source.n193 source.t14 149.524
R227 source.n493 source.n487 104.615
R228 source.n494 source.n493 104.615
R229 source.n494 source.n483 104.615
R230 source.n501 source.n483 104.615
R231 source.n502 source.n501 104.615
R232 source.n502 source.n479 104.615
R233 source.n510 source.n479 104.615
R234 source.n511 source.n510 104.615
R235 source.n512 source.n511 104.615
R236 source.n512 source.n475 104.615
R237 source.n519 source.n475 104.615
R238 source.n520 source.n519 104.615
R239 source.n520 source.n471 104.615
R240 source.n527 source.n471 104.615
R241 source.n528 source.n527 104.615
R242 source.n528 source.n467 104.615
R243 source.n535 source.n467 104.615
R244 source.n536 source.n535 104.615
R245 source.n536 source.n463 104.615
R246 source.n543 source.n463 104.615
R247 source.n544 source.n543 104.615
R248 source.n544 source.n459 104.615
R249 source.n551 source.n459 104.615
R250 source.n553 source.n551 104.615
R251 source.n553 source.n552 104.615
R252 source.n552 source.n455 104.615
R253 source.n561 source.n455 104.615
R254 source.n562 source.n561 104.615
R255 source.n562 source.n451 104.615
R256 source.n569 source.n451 104.615
R257 source.n570 source.n569 104.615
R258 source.n570 source.n447 104.615
R259 source.n577 source.n447 104.615
R260 source.n578 source.n577 104.615
R261 source.n347 source.n341 104.615
R262 source.n348 source.n347 104.615
R263 source.n348 source.n337 104.615
R264 source.n355 source.n337 104.615
R265 source.n356 source.n355 104.615
R266 source.n356 source.n333 104.615
R267 source.n364 source.n333 104.615
R268 source.n365 source.n364 104.615
R269 source.n366 source.n365 104.615
R270 source.n366 source.n329 104.615
R271 source.n373 source.n329 104.615
R272 source.n374 source.n373 104.615
R273 source.n374 source.n325 104.615
R274 source.n381 source.n325 104.615
R275 source.n382 source.n381 104.615
R276 source.n382 source.n321 104.615
R277 source.n389 source.n321 104.615
R278 source.n390 source.n389 104.615
R279 source.n390 source.n317 104.615
R280 source.n397 source.n317 104.615
R281 source.n398 source.n397 104.615
R282 source.n398 source.n313 104.615
R283 source.n405 source.n313 104.615
R284 source.n407 source.n405 104.615
R285 source.n407 source.n406 104.615
R286 source.n406 source.n309 104.615
R287 source.n415 source.n309 104.615
R288 source.n416 source.n415 104.615
R289 source.n416 source.n305 104.615
R290 source.n423 source.n305 104.615
R291 source.n424 source.n423 104.615
R292 source.n424 source.n301 104.615
R293 source.n431 source.n301 104.615
R294 source.n432 source.n431 104.615
R295 source.n134 source.n133 104.615
R296 source.n133 source.n3 104.615
R297 source.n126 source.n3 104.615
R298 source.n126 source.n125 104.615
R299 source.n125 source.n7 104.615
R300 source.n118 source.n7 104.615
R301 source.n118 source.n117 104.615
R302 source.n117 source.n11 104.615
R303 source.n15 source.n11 104.615
R304 source.n109 source.n15 104.615
R305 source.n109 source.n108 104.615
R306 source.n108 source.n16 104.615
R307 source.n101 source.n16 104.615
R308 source.n101 source.n100 104.615
R309 source.n100 source.n20 104.615
R310 source.n93 source.n20 104.615
R311 source.n93 source.n92 104.615
R312 source.n92 source.n24 104.615
R313 source.n85 source.n24 104.615
R314 source.n85 source.n84 104.615
R315 source.n84 source.n28 104.615
R316 source.n77 source.n28 104.615
R317 source.n77 source.n76 104.615
R318 source.n76 source.n32 104.615
R319 source.n69 source.n32 104.615
R320 source.n69 source.n68 104.615
R321 source.n68 source.n67 104.615
R322 source.n67 source.n36 104.615
R323 source.n60 source.n36 104.615
R324 source.n60 source.n59 104.615
R325 source.n59 source.n41 104.615
R326 source.n52 source.n41 104.615
R327 source.n52 source.n51 104.615
R328 source.n51 source.n45 104.615
R329 source.n280 source.n279 104.615
R330 source.n279 source.n149 104.615
R331 source.n272 source.n149 104.615
R332 source.n272 source.n271 104.615
R333 source.n271 source.n153 104.615
R334 source.n264 source.n153 104.615
R335 source.n264 source.n263 104.615
R336 source.n263 source.n157 104.615
R337 source.n161 source.n157 104.615
R338 source.n255 source.n161 104.615
R339 source.n255 source.n254 104.615
R340 source.n254 source.n162 104.615
R341 source.n247 source.n162 104.615
R342 source.n247 source.n246 104.615
R343 source.n246 source.n166 104.615
R344 source.n239 source.n166 104.615
R345 source.n239 source.n238 104.615
R346 source.n238 source.n170 104.615
R347 source.n231 source.n170 104.615
R348 source.n231 source.n230 104.615
R349 source.n230 source.n174 104.615
R350 source.n223 source.n174 104.615
R351 source.n223 source.n222 104.615
R352 source.n222 source.n178 104.615
R353 source.n215 source.n178 104.615
R354 source.n215 source.n214 104.615
R355 source.n214 source.n213 104.615
R356 source.n213 source.n182 104.615
R357 source.n206 source.n182 104.615
R358 source.n206 source.n205 104.615
R359 source.n205 source.n187 104.615
R360 source.n198 source.n187 104.615
R361 source.n198 source.n197 104.615
R362 source.n197 source.n191 104.615
R363 source.t23 source.n487 52.3082
R364 source.t26 source.n341 52.3082
R365 source.t0 source.n45 52.3082
R366 source.t14 source.n191 52.3082
R367 source.n443 source.n442 42.0366
R368 source.n441 source.n440 42.0366
R369 source.n439 source.n438 42.0366
R370 source.n297 source.n296 42.0366
R371 source.n295 source.n294 42.0366
R372 source.n293 source.n292 42.0366
R373 source.n141 source.n140 42.0366
R374 source.n143 source.n142 42.0366
R375 source.n145 source.n144 42.0366
R376 source.n287 source.n286 42.0366
R377 source.n289 source.n288 42.0366
R378 source.n291 source.n290 42.0366
R379 source.n293 source.n291 32.9121
R380 source.n583 source.n582 30.6338
R381 source.n437 source.n436 30.6338
R382 source.n139 source.n138 30.6338
R383 source.n285 source.n284 30.6338
R384 source.n584 source.n139 26.3172
R385 source.n513 source.n478 13.1884
R386 source.n560 source.n559 13.1884
R387 source.n367 source.n332 13.1884
R388 source.n414 source.n413 13.1884
R389 source.n116 source.n115 13.1884
R390 source.n70 source.n35 13.1884
R391 source.n262 source.n261 13.1884
R392 source.n216 source.n181 13.1884
R393 source.n509 source.n508 12.8005
R394 source.n514 source.n476 12.8005
R395 source.n558 source.n456 12.8005
R396 source.n563 source.n454 12.8005
R397 source.n363 source.n362 12.8005
R398 source.n368 source.n330 12.8005
R399 source.n412 source.n310 12.8005
R400 source.n417 source.n308 12.8005
R401 source.n119 source.n10 12.8005
R402 source.n114 source.n12 12.8005
R403 source.n71 source.n33 12.8005
R404 source.n66 source.n37 12.8005
R405 source.n265 source.n156 12.8005
R406 source.n260 source.n158 12.8005
R407 source.n217 source.n179 12.8005
R408 source.n212 source.n183 12.8005
R409 source.n507 source.n480 12.0247
R410 source.n518 source.n517 12.0247
R411 source.n555 source.n554 12.0247
R412 source.n564 source.n452 12.0247
R413 source.n361 source.n334 12.0247
R414 source.n372 source.n371 12.0247
R415 source.n409 source.n408 12.0247
R416 source.n418 source.n306 12.0247
R417 source.n120 source.n8 12.0247
R418 source.n111 source.n110 12.0247
R419 source.n75 source.n74 12.0247
R420 source.n65 source.n38 12.0247
R421 source.n266 source.n154 12.0247
R422 source.n257 source.n256 12.0247
R423 source.n221 source.n220 12.0247
R424 source.n211 source.n184 12.0247
R425 source.n504 source.n503 11.249
R426 source.n521 source.n474 11.249
R427 source.n550 source.n458 11.249
R428 source.n568 source.n567 11.249
R429 source.n358 source.n357 11.249
R430 source.n375 source.n328 11.249
R431 source.n404 source.n312 11.249
R432 source.n422 source.n421 11.249
R433 source.n124 source.n123 11.249
R434 source.n107 source.n14 11.249
R435 source.n78 source.n31 11.249
R436 source.n62 source.n61 11.249
R437 source.n270 source.n269 11.249
R438 source.n253 source.n160 11.249
R439 source.n224 source.n177 11.249
R440 source.n208 source.n207 11.249
R441 source.n500 source.n482 10.4732
R442 source.n522 source.n472 10.4732
R443 source.n549 source.n460 10.4732
R444 source.n571 source.n450 10.4732
R445 source.n354 source.n336 10.4732
R446 source.n376 source.n326 10.4732
R447 source.n403 source.n314 10.4732
R448 source.n425 source.n304 10.4732
R449 source.n127 source.n6 10.4732
R450 source.n106 source.n17 10.4732
R451 source.n79 source.n29 10.4732
R452 source.n58 source.n40 10.4732
R453 source.n273 source.n152 10.4732
R454 source.n252 source.n163 10.4732
R455 source.n225 source.n175 10.4732
R456 source.n204 source.n186 10.4732
R457 source.n489 source.n488 10.2747
R458 source.n343 source.n342 10.2747
R459 source.n47 source.n46 10.2747
R460 source.n193 source.n192 10.2747
R461 source.n499 source.n484 9.69747
R462 source.n526 source.n525 9.69747
R463 source.n546 source.n545 9.69747
R464 source.n572 source.n448 9.69747
R465 source.n353 source.n338 9.69747
R466 source.n380 source.n379 9.69747
R467 source.n400 source.n399 9.69747
R468 source.n426 source.n302 9.69747
R469 source.n128 source.n4 9.69747
R470 source.n103 source.n102 9.69747
R471 source.n83 source.n82 9.69747
R472 source.n57 source.n42 9.69747
R473 source.n274 source.n150 9.69747
R474 source.n249 source.n248 9.69747
R475 source.n229 source.n228 9.69747
R476 source.n203 source.n188 9.69747
R477 source.n582 source.n581 9.45567
R478 source.n436 source.n435 9.45567
R479 source.n138 source.n137 9.45567
R480 source.n284 source.n283 9.45567
R481 source.n446 source.n445 9.3005
R482 source.n575 source.n574 9.3005
R483 source.n573 source.n572 9.3005
R484 source.n450 source.n449 9.3005
R485 source.n567 source.n566 9.3005
R486 source.n565 source.n564 9.3005
R487 source.n454 source.n453 9.3005
R488 source.n533 source.n532 9.3005
R489 source.n531 source.n530 9.3005
R490 source.n470 source.n469 9.3005
R491 source.n525 source.n524 9.3005
R492 source.n523 source.n522 9.3005
R493 source.n474 source.n473 9.3005
R494 source.n517 source.n516 9.3005
R495 source.n515 source.n514 9.3005
R496 source.n491 source.n490 9.3005
R497 source.n486 source.n485 9.3005
R498 source.n497 source.n496 9.3005
R499 source.n499 source.n498 9.3005
R500 source.n482 source.n481 9.3005
R501 source.n505 source.n504 9.3005
R502 source.n507 source.n506 9.3005
R503 source.n508 source.n477 9.3005
R504 source.n466 source.n465 9.3005
R505 source.n539 source.n538 9.3005
R506 source.n541 source.n540 9.3005
R507 source.n462 source.n461 9.3005
R508 source.n547 source.n546 9.3005
R509 source.n549 source.n548 9.3005
R510 source.n458 source.n457 9.3005
R511 source.n556 source.n555 9.3005
R512 source.n558 source.n557 9.3005
R513 source.n581 source.n580 9.3005
R514 source.n300 source.n299 9.3005
R515 source.n429 source.n428 9.3005
R516 source.n427 source.n426 9.3005
R517 source.n304 source.n303 9.3005
R518 source.n421 source.n420 9.3005
R519 source.n419 source.n418 9.3005
R520 source.n308 source.n307 9.3005
R521 source.n387 source.n386 9.3005
R522 source.n385 source.n384 9.3005
R523 source.n324 source.n323 9.3005
R524 source.n379 source.n378 9.3005
R525 source.n377 source.n376 9.3005
R526 source.n328 source.n327 9.3005
R527 source.n371 source.n370 9.3005
R528 source.n369 source.n368 9.3005
R529 source.n345 source.n344 9.3005
R530 source.n340 source.n339 9.3005
R531 source.n351 source.n350 9.3005
R532 source.n353 source.n352 9.3005
R533 source.n336 source.n335 9.3005
R534 source.n359 source.n358 9.3005
R535 source.n361 source.n360 9.3005
R536 source.n362 source.n331 9.3005
R537 source.n320 source.n319 9.3005
R538 source.n393 source.n392 9.3005
R539 source.n395 source.n394 9.3005
R540 source.n316 source.n315 9.3005
R541 source.n401 source.n400 9.3005
R542 source.n403 source.n402 9.3005
R543 source.n312 source.n311 9.3005
R544 source.n410 source.n409 9.3005
R545 source.n412 source.n411 9.3005
R546 source.n435 source.n434 9.3005
R547 source.n49 source.n48 9.3005
R548 source.n44 source.n43 9.3005
R549 source.n55 source.n54 9.3005
R550 source.n57 source.n56 9.3005
R551 source.n40 source.n39 9.3005
R552 source.n63 source.n62 9.3005
R553 source.n65 source.n64 9.3005
R554 source.n37 source.n34 9.3005
R555 source.n96 source.n95 9.3005
R556 source.n98 source.n97 9.3005
R557 source.n19 source.n18 9.3005
R558 source.n104 source.n103 9.3005
R559 source.n106 source.n105 9.3005
R560 source.n14 source.n13 9.3005
R561 source.n112 source.n111 9.3005
R562 source.n114 source.n113 9.3005
R563 source.n137 source.n136 9.3005
R564 source.n2 source.n1 9.3005
R565 source.n131 source.n130 9.3005
R566 source.n129 source.n128 9.3005
R567 source.n6 source.n5 9.3005
R568 source.n123 source.n122 9.3005
R569 source.n121 source.n120 9.3005
R570 source.n10 source.n9 9.3005
R571 source.n23 source.n22 9.3005
R572 source.n90 source.n89 9.3005
R573 source.n88 source.n87 9.3005
R574 source.n27 source.n26 9.3005
R575 source.n82 source.n81 9.3005
R576 source.n80 source.n79 9.3005
R577 source.n31 source.n30 9.3005
R578 source.n74 source.n73 9.3005
R579 source.n72 source.n71 9.3005
R580 source.n195 source.n194 9.3005
R581 source.n190 source.n189 9.3005
R582 source.n201 source.n200 9.3005
R583 source.n203 source.n202 9.3005
R584 source.n186 source.n185 9.3005
R585 source.n209 source.n208 9.3005
R586 source.n211 source.n210 9.3005
R587 source.n183 source.n180 9.3005
R588 source.n242 source.n241 9.3005
R589 source.n244 source.n243 9.3005
R590 source.n165 source.n164 9.3005
R591 source.n250 source.n249 9.3005
R592 source.n252 source.n251 9.3005
R593 source.n160 source.n159 9.3005
R594 source.n258 source.n257 9.3005
R595 source.n260 source.n259 9.3005
R596 source.n283 source.n282 9.3005
R597 source.n148 source.n147 9.3005
R598 source.n277 source.n276 9.3005
R599 source.n275 source.n274 9.3005
R600 source.n152 source.n151 9.3005
R601 source.n269 source.n268 9.3005
R602 source.n267 source.n266 9.3005
R603 source.n156 source.n155 9.3005
R604 source.n169 source.n168 9.3005
R605 source.n236 source.n235 9.3005
R606 source.n234 source.n233 9.3005
R607 source.n173 source.n172 9.3005
R608 source.n228 source.n227 9.3005
R609 source.n226 source.n225 9.3005
R610 source.n177 source.n176 9.3005
R611 source.n220 source.n219 9.3005
R612 source.n218 source.n217 9.3005
R613 source.n496 source.n495 8.92171
R614 source.n529 source.n470 8.92171
R615 source.n542 source.n462 8.92171
R616 source.n576 source.n575 8.92171
R617 source.n350 source.n349 8.92171
R618 source.n383 source.n324 8.92171
R619 source.n396 source.n316 8.92171
R620 source.n430 source.n429 8.92171
R621 source.n132 source.n131 8.92171
R622 source.n99 source.n19 8.92171
R623 source.n86 source.n27 8.92171
R624 source.n54 source.n53 8.92171
R625 source.n278 source.n277 8.92171
R626 source.n245 source.n165 8.92171
R627 source.n232 source.n173 8.92171
R628 source.n200 source.n199 8.92171
R629 source.n492 source.n486 8.14595
R630 source.n530 source.n468 8.14595
R631 source.n541 source.n464 8.14595
R632 source.n579 source.n446 8.14595
R633 source.n346 source.n340 8.14595
R634 source.n384 source.n322 8.14595
R635 source.n395 source.n318 8.14595
R636 source.n433 source.n300 8.14595
R637 source.n135 source.n2 8.14595
R638 source.n98 source.n21 8.14595
R639 source.n87 source.n25 8.14595
R640 source.n50 source.n44 8.14595
R641 source.n281 source.n148 8.14595
R642 source.n244 source.n167 8.14595
R643 source.n233 source.n171 8.14595
R644 source.n196 source.n190 8.14595
R645 source.n491 source.n488 7.3702
R646 source.n534 source.n533 7.3702
R647 source.n538 source.n537 7.3702
R648 source.n580 source.n444 7.3702
R649 source.n345 source.n342 7.3702
R650 source.n388 source.n387 7.3702
R651 source.n392 source.n391 7.3702
R652 source.n434 source.n298 7.3702
R653 source.n136 source.n0 7.3702
R654 source.n95 source.n94 7.3702
R655 source.n91 source.n90 7.3702
R656 source.n49 source.n46 7.3702
R657 source.n282 source.n146 7.3702
R658 source.n241 source.n240 7.3702
R659 source.n237 source.n236 7.3702
R660 source.n195 source.n192 7.3702
R661 source.n534 source.n466 6.59444
R662 source.n537 source.n466 6.59444
R663 source.n582 source.n444 6.59444
R664 source.n388 source.n320 6.59444
R665 source.n391 source.n320 6.59444
R666 source.n436 source.n298 6.59444
R667 source.n138 source.n0 6.59444
R668 source.n94 source.n23 6.59444
R669 source.n91 source.n23 6.59444
R670 source.n284 source.n146 6.59444
R671 source.n240 source.n169 6.59444
R672 source.n237 source.n169 6.59444
R673 source.n492 source.n491 5.81868
R674 source.n533 source.n468 5.81868
R675 source.n538 source.n464 5.81868
R676 source.n580 source.n579 5.81868
R677 source.n346 source.n345 5.81868
R678 source.n387 source.n322 5.81868
R679 source.n392 source.n318 5.81868
R680 source.n434 source.n433 5.81868
R681 source.n136 source.n135 5.81868
R682 source.n95 source.n21 5.81868
R683 source.n90 source.n25 5.81868
R684 source.n50 source.n49 5.81868
R685 source.n282 source.n281 5.81868
R686 source.n241 source.n167 5.81868
R687 source.n236 source.n171 5.81868
R688 source.n196 source.n195 5.81868
R689 source.n584 source.n583 5.7074
R690 source.n495 source.n486 5.04292
R691 source.n530 source.n529 5.04292
R692 source.n542 source.n541 5.04292
R693 source.n576 source.n446 5.04292
R694 source.n349 source.n340 5.04292
R695 source.n384 source.n383 5.04292
R696 source.n396 source.n395 5.04292
R697 source.n430 source.n300 5.04292
R698 source.n132 source.n2 5.04292
R699 source.n99 source.n98 5.04292
R700 source.n87 source.n86 5.04292
R701 source.n53 source.n44 5.04292
R702 source.n278 source.n148 5.04292
R703 source.n245 source.n244 5.04292
R704 source.n233 source.n232 5.04292
R705 source.n199 source.n190 5.04292
R706 source.n496 source.n484 4.26717
R707 source.n526 source.n470 4.26717
R708 source.n545 source.n462 4.26717
R709 source.n575 source.n448 4.26717
R710 source.n350 source.n338 4.26717
R711 source.n380 source.n324 4.26717
R712 source.n399 source.n316 4.26717
R713 source.n429 source.n302 4.26717
R714 source.n131 source.n4 4.26717
R715 source.n102 source.n19 4.26717
R716 source.n83 source.n27 4.26717
R717 source.n54 source.n42 4.26717
R718 source.n277 source.n150 4.26717
R719 source.n248 source.n165 4.26717
R720 source.n229 source.n173 4.26717
R721 source.n200 source.n188 4.26717
R722 source.n500 source.n499 3.49141
R723 source.n525 source.n472 3.49141
R724 source.n546 source.n460 3.49141
R725 source.n572 source.n571 3.49141
R726 source.n354 source.n353 3.49141
R727 source.n379 source.n326 3.49141
R728 source.n400 source.n314 3.49141
R729 source.n426 source.n425 3.49141
R730 source.n128 source.n127 3.49141
R731 source.n103 source.n17 3.49141
R732 source.n82 source.n29 3.49141
R733 source.n58 source.n57 3.49141
R734 source.n274 source.n273 3.49141
R735 source.n249 source.n163 3.49141
R736 source.n228 source.n175 3.49141
R737 source.n204 source.n203 3.49141
R738 source.n48 source.n47 2.84303
R739 source.n194 source.n193 2.84303
R740 source.n490 source.n489 2.84303
R741 source.n344 source.n343 2.84303
R742 source.n503 source.n482 2.71565
R743 source.n522 source.n521 2.71565
R744 source.n550 source.n549 2.71565
R745 source.n568 source.n450 2.71565
R746 source.n357 source.n336 2.71565
R747 source.n376 source.n375 2.71565
R748 source.n404 source.n403 2.71565
R749 source.n422 source.n304 2.71565
R750 source.n124 source.n6 2.71565
R751 source.n107 source.n106 2.71565
R752 source.n79 source.n78 2.71565
R753 source.n61 source.n40 2.71565
R754 source.n270 source.n152 2.71565
R755 source.n253 source.n252 2.71565
R756 source.n225 source.n224 2.71565
R757 source.n207 source.n186 2.71565
R758 source.n504 source.n480 1.93989
R759 source.n518 source.n474 1.93989
R760 source.n554 source.n458 1.93989
R761 source.n567 source.n452 1.93989
R762 source.n358 source.n334 1.93989
R763 source.n372 source.n328 1.93989
R764 source.n408 source.n312 1.93989
R765 source.n421 source.n306 1.93989
R766 source.n123 source.n8 1.93989
R767 source.n110 source.n14 1.93989
R768 source.n75 source.n31 1.93989
R769 source.n62 source.n38 1.93989
R770 source.n269 source.n154 1.93989
R771 source.n256 source.n160 1.93989
R772 source.n221 source.n177 1.93989
R773 source.n208 source.n184 1.93989
R774 source.n509 source.n507 1.16414
R775 source.n517 source.n476 1.16414
R776 source.n555 source.n456 1.16414
R777 source.n564 source.n563 1.16414
R778 source.n363 source.n361 1.16414
R779 source.n371 source.n330 1.16414
R780 source.n409 source.n310 1.16414
R781 source.n418 source.n417 1.16414
R782 source.n120 source.n119 1.16414
R783 source.n111 source.n12 1.16414
R784 source.n74 source.n33 1.16414
R785 source.n66 source.n65 1.16414
R786 source.n266 source.n265 1.16414
R787 source.n257 source.n158 1.16414
R788 source.n220 source.n179 1.16414
R789 source.n212 source.n211 1.16414
R790 source.n285 source.n145 0.914293
R791 source.n439 source.n437 0.914293
R792 source.n291 source.n289 0.888431
R793 source.n289 source.n287 0.888431
R794 source.n287 source.n285 0.888431
R795 source.n145 source.n143 0.888431
R796 source.n143 source.n141 0.888431
R797 source.n141 source.n139 0.888431
R798 source.n295 source.n293 0.888431
R799 source.n297 source.n295 0.888431
R800 source.n437 source.n297 0.888431
R801 source.n441 source.n439 0.888431
R802 source.n443 source.n441 0.888431
R803 source.n583 source.n443 0.888431
R804 source.n442 source.t25 0.7925
R805 source.n442 source.t12 0.7925
R806 source.n440 source.t22 0.7925
R807 source.n440 source.t20 0.7925
R808 source.n438 source.t24 0.7925
R809 source.n438 source.t15 0.7925
R810 source.n296 source.t10 0.7925
R811 source.n296 source.t7 0.7925
R812 source.n294 source.t11 0.7925
R813 source.n294 source.t5 0.7925
R814 source.n292 source.t27 0.7925
R815 source.n292 source.t2 0.7925
R816 source.n140 source.t6 0.7925
R817 source.n140 source.t3 0.7925
R818 source.n142 source.t1 0.7925
R819 source.n142 source.t4 0.7925
R820 source.n144 source.t9 0.7925
R821 source.n144 source.t8 0.7925
R822 source.n286 source.t13 0.7925
R823 source.n286 source.t18 0.7925
R824 source.n288 source.t16 0.7925
R825 source.n288 source.t21 0.7925
R826 source.n290 source.t17 0.7925
R827 source.n290 source.t19 0.7925
R828 source.n508 source.n478 0.388379
R829 source.n514 source.n513 0.388379
R830 source.n559 source.n558 0.388379
R831 source.n560 source.n454 0.388379
R832 source.n362 source.n332 0.388379
R833 source.n368 source.n367 0.388379
R834 source.n413 source.n412 0.388379
R835 source.n414 source.n308 0.388379
R836 source.n116 source.n10 0.388379
R837 source.n115 source.n114 0.388379
R838 source.n71 source.n70 0.388379
R839 source.n37 source.n35 0.388379
R840 source.n262 source.n156 0.388379
R841 source.n261 source.n260 0.388379
R842 source.n217 source.n216 0.388379
R843 source.n183 source.n181 0.388379
R844 source source.n584 0.188
R845 source.n490 source.n485 0.155672
R846 source.n497 source.n485 0.155672
R847 source.n498 source.n497 0.155672
R848 source.n498 source.n481 0.155672
R849 source.n505 source.n481 0.155672
R850 source.n506 source.n505 0.155672
R851 source.n506 source.n477 0.155672
R852 source.n515 source.n477 0.155672
R853 source.n516 source.n515 0.155672
R854 source.n516 source.n473 0.155672
R855 source.n523 source.n473 0.155672
R856 source.n524 source.n523 0.155672
R857 source.n524 source.n469 0.155672
R858 source.n531 source.n469 0.155672
R859 source.n532 source.n531 0.155672
R860 source.n532 source.n465 0.155672
R861 source.n539 source.n465 0.155672
R862 source.n540 source.n539 0.155672
R863 source.n540 source.n461 0.155672
R864 source.n547 source.n461 0.155672
R865 source.n548 source.n547 0.155672
R866 source.n548 source.n457 0.155672
R867 source.n556 source.n457 0.155672
R868 source.n557 source.n556 0.155672
R869 source.n557 source.n453 0.155672
R870 source.n565 source.n453 0.155672
R871 source.n566 source.n565 0.155672
R872 source.n566 source.n449 0.155672
R873 source.n573 source.n449 0.155672
R874 source.n574 source.n573 0.155672
R875 source.n574 source.n445 0.155672
R876 source.n581 source.n445 0.155672
R877 source.n344 source.n339 0.155672
R878 source.n351 source.n339 0.155672
R879 source.n352 source.n351 0.155672
R880 source.n352 source.n335 0.155672
R881 source.n359 source.n335 0.155672
R882 source.n360 source.n359 0.155672
R883 source.n360 source.n331 0.155672
R884 source.n369 source.n331 0.155672
R885 source.n370 source.n369 0.155672
R886 source.n370 source.n327 0.155672
R887 source.n377 source.n327 0.155672
R888 source.n378 source.n377 0.155672
R889 source.n378 source.n323 0.155672
R890 source.n385 source.n323 0.155672
R891 source.n386 source.n385 0.155672
R892 source.n386 source.n319 0.155672
R893 source.n393 source.n319 0.155672
R894 source.n394 source.n393 0.155672
R895 source.n394 source.n315 0.155672
R896 source.n401 source.n315 0.155672
R897 source.n402 source.n401 0.155672
R898 source.n402 source.n311 0.155672
R899 source.n410 source.n311 0.155672
R900 source.n411 source.n410 0.155672
R901 source.n411 source.n307 0.155672
R902 source.n419 source.n307 0.155672
R903 source.n420 source.n419 0.155672
R904 source.n420 source.n303 0.155672
R905 source.n427 source.n303 0.155672
R906 source.n428 source.n427 0.155672
R907 source.n428 source.n299 0.155672
R908 source.n435 source.n299 0.155672
R909 source.n137 source.n1 0.155672
R910 source.n130 source.n1 0.155672
R911 source.n130 source.n129 0.155672
R912 source.n129 source.n5 0.155672
R913 source.n122 source.n5 0.155672
R914 source.n122 source.n121 0.155672
R915 source.n121 source.n9 0.155672
R916 source.n113 source.n9 0.155672
R917 source.n113 source.n112 0.155672
R918 source.n112 source.n13 0.155672
R919 source.n105 source.n13 0.155672
R920 source.n105 source.n104 0.155672
R921 source.n104 source.n18 0.155672
R922 source.n97 source.n18 0.155672
R923 source.n97 source.n96 0.155672
R924 source.n96 source.n22 0.155672
R925 source.n89 source.n22 0.155672
R926 source.n89 source.n88 0.155672
R927 source.n88 source.n26 0.155672
R928 source.n81 source.n26 0.155672
R929 source.n81 source.n80 0.155672
R930 source.n80 source.n30 0.155672
R931 source.n73 source.n30 0.155672
R932 source.n73 source.n72 0.155672
R933 source.n72 source.n34 0.155672
R934 source.n64 source.n34 0.155672
R935 source.n64 source.n63 0.155672
R936 source.n63 source.n39 0.155672
R937 source.n56 source.n39 0.155672
R938 source.n56 source.n55 0.155672
R939 source.n55 source.n43 0.155672
R940 source.n48 source.n43 0.155672
R941 source.n283 source.n147 0.155672
R942 source.n276 source.n147 0.155672
R943 source.n276 source.n275 0.155672
R944 source.n275 source.n151 0.155672
R945 source.n268 source.n151 0.155672
R946 source.n268 source.n267 0.155672
R947 source.n267 source.n155 0.155672
R948 source.n259 source.n155 0.155672
R949 source.n259 source.n258 0.155672
R950 source.n258 source.n159 0.155672
R951 source.n251 source.n159 0.155672
R952 source.n251 source.n250 0.155672
R953 source.n250 source.n164 0.155672
R954 source.n243 source.n164 0.155672
R955 source.n243 source.n242 0.155672
R956 source.n242 source.n168 0.155672
R957 source.n235 source.n168 0.155672
R958 source.n235 source.n234 0.155672
R959 source.n234 source.n172 0.155672
R960 source.n227 source.n172 0.155672
R961 source.n227 source.n226 0.155672
R962 source.n226 source.n176 0.155672
R963 source.n219 source.n176 0.155672
R964 source.n219 source.n218 0.155672
R965 source.n218 source.n180 0.155672
R966 source.n210 source.n180 0.155672
R967 source.n210 source.n209 0.155672
R968 source.n209 source.n185 0.155672
R969 source.n202 source.n185 0.155672
R970 source.n202 source.n201 0.155672
R971 source.n201 source.n189 0.155672
R972 source.n194 source.n189 0.155672
R973 drain_right.n134 drain_right.n0 289.615
R974 drain_right.n284 drain_right.n150 289.615
R975 drain_right.n44 drain_right.n43 185
R976 drain_right.n49 drain_right.n48 185
R977 drain_right.n51 drain_right.n50 185
R978 drain_right.n40 drain_right.n39 185
R979 drain_right.n57 drain_right.n56 185
R980 drain_right.n59 drain_right.n58 185
R981 drain_right.n36 drain_right.n35 185
R982 drain_right.n66 drain_right.n65 185
R983 drain_right.n67 drain_right.n34 185
R984 drain_right.n69 drain_right.n68 185
R985 drain_right.n32 drain_right.n31 185
R986 drain_right.n75 drain_right.n74 185
R987 drain_right.n77 drain_right.n76 185
R988 drain_right.n28 drain_right.n27 185
R989 drain_right.n83 drain_right.n82 185
R990 drain_right.n85 drain_right.n84 185
R991 drain_right.n24 drain_right.n23 185
R992 drain_right.n91 drain_right.n90 185
R993 drain_right.n93 drain_right.n92 185
R994 drain_right.n20 drain_right.n19 185
R995 drain_right.n99 drain_right.n98 185
R996 drain_right.n101 drain_right.n100 185
R997 drain_right.n16 drain_right.n15 185
R998 drain_right.n107 drain_right.n106 185
R999 drain_right.n110 drain_right.n109 185
R1000 drain_right.n108 drain_right.n12 185
R1001 drain_right.n115 drain_right.n11 185
R1002 drain_right.n117 drain_right.n116 185
R1003 drain_right.n119 drain_right.n118 185
R1004 drain_right.n8 drain_right.n7 185
R1005 drain_right.n125 drain_right.n124 185
R1006 drain_right.n127 drain_right.n126 185
R1007 drain_right.n4 drain_right.n3 185
R1008 drain_right.n133 drain_right.n132 185
R1009 drain_right.n135 drain_right.n134 185
R1010 drain_right.n285 drain_right.n284 185
R1011 drain_right.n283 drain_right.n282 185
R1012 drain_right.n154 drain_right.n153 185
R1013 drain_right.n277 drain_right.n276 185
R1014 drain_right.n275 drain_right.n274 185
R1015 drain_right.n158 drain_right.n157 185
R1016 drain_right.n269 drain_right.n268 185
R1017 drain_right.n267 drain_right.n266 185
R1018 drain_right.n265 drain_right.n161 185
R1019 drain_right.n165 drain_right.n162 185
R1020 drain_right.n260 drain_right.n259 185
R1021 drain_right.n258 drain_right.n257 185
R1022 drain_right.n167 drain_right.n166 185
R1023 drain_right.n252 drain_right.n251 185
R1024 drain_right.n250 drain_right.n249 185
R1025 drain_right.n171 drain_right.n170 185
R1026 drain_right.n244 drain_right.n243 185
R1027 drain_right.n242 drain_right.n241 185
R1028 drain_right.n175 drain_right.n174 185
R1029 drain_right.n236 drain_right.n235 185
R1030 drain_right.n234 drain_right.n233 185
R1031 drain_right.n179 drain_right.n178 185
R1032 drain_right.n228 drain_right.n227 185
R1033 drain_right.n226 drain_right.n225 185
R1034 drain_right.n183 drain_right.n182 185
R1035 drain_right.n220 drain_right.n219 185
R1036 drain_right.n218 drain_right.n185 185
R1037 drain_right.n217 drain_right.n216 185
R1038 drain_right.n188 drain_right.n186 185
R1039 drain_right.n211 drain_right.n210 185
R1040 drain_right.n209 drain_right.n208 185
R1041 drain_right.n192 drain_right.n191 185
R1042 drain_right.n203 drain_right.n202 185
R1043 drain_right.n201 drain_right.n200 185
R1044 drain_right.n196 drain_right.n195 185
R1045 drain_right.n45 drain_right.t8 149.524
R1046 drain_right.n197 drain_right.t7 149.524
R1047 drain_right.n49 drain_right.n43 104.615
R1048 drain_right.n50 drain_right.n49 104.615
R1049 drain_right.n50 drain_right.n39 104.615
R1050 drain_right.n57 drain_right.n39 104.615
R1051 drain_right.n58 drain_right.n57 104.615
R1052 drain_right.n58 drain_right.n35 104.615
R1053 drain_right.n66 drain_right.n35 104.615
R1054 drain_right.n67 drain_right.n66 104.615
R1055 drain_right.n68 drain_right.n67 104.615
R1056 drain_right.n68 drain_right.n31 104.615
R1057 drain_right.n75 drain_right.n31 104.615
R1058 drain_right.n76 drain_right.n75 104.615
R1059 drain_right.n76 drain_right.n27 104.615
R1060 drain_right.n83 drain_right.n27 104.615
R1061 drain_right.n84 drain_right.n83 104.615
R1062 drain_right.n84 drain_right.n23 104.615
R1063 drain_right.n91 drain_right.n23 104.615
R1064 drain_right.n92 drain_right.n91 104.615
R1065 drain_right.n92 drain_right.n19 104.615
R1066 drain_right.n99 drain_right.n19 104.615
R1067 drain_right.n100 drain_right.n99 104.615
R1068 drain_right.n100 drain_right.n15 104.615
R1069 drain_right.n107 drain_right.n15 104.615
R1070 drain_right.n109 drain_right.n107 104.615
R1071 drain_right.n109 drain_right.n108 104.615
R1072 drain_right.n108 drain_right.n11 104.615
R1073 drain_right.n117 drain_right.n11 104.615
R1074 drain_right.n118 drain_right.n117 104.615
R1075 drain_right.n118 drain_right.n7 104.615
R1076 drain_right.n125 drain_right.n7 104.615
R1077 drain_right.n126 drain_right.n125 104.615
R1078 drain_right.n126 drain_right.n3 104.615
R1079 drain_right.n133 drain_right.n3 104.615
R1080 drain_right.n134 drain_right.n133 104.615
R1081 drain_right.n284 drain_right.n283 104.615
R1082 drain_right.n283 drain_right.n153 104.615
R1083 drain_right.n276 drain_right.n153 104.615
R1084 drain_right.n276 drain_right.n275 104.615
R1085 drain_right.n275 drain_right.n157 104.615
R1086 drain_right.n268 drain_right.n157 104.615
R1087 drain_right.n268 drain_right.n267 104.615
R1088 drain_right.n267 drain_right.n161 104.615
R1089 drain_right.n165 drain_right.n161 104.615
R1090 drain_right.n259 drain_right.n165 104.615
R1091 drain_right.n259 drain_right.n258 104.615
R1092 drain_right.n258 drain_right.n166 104.615
R1093 drain_right.n251 drain_right.n166 104.615
R1094 drain_right.n251 drain_right.n250 104.615
R1095 drain_right.n250 drain_right.n170 104.615
R1096 drain_right.n243 drain_right.n170 104.615
R1097 drain_right.n243 drain_right.n242 104.615
R1098 drain_right.n242 drain_right.n174 104.615
R1099 drain_right.n235 drain_right.n174 104.615
R1100 drain_right.n235 drain_right.n234 104.615
R1101 drain_right.n234 drain_right.n178 104.615
R1102 drain_right.n227 drain_right.n178 104.615
R1103 drain_right.n227 drain_right.n226 104.615
R1104 drain_right.n226 drain_right.n182 104.615
R1105 drain_right.n219 drain_right.n182 104.615
R1106 drain_right.n219 drain_right.n218 104.615
R1107 drain_right.n218 drain_right.n217 104.615
R1108 drain_right.n217 drain_right.n186 104.615
R1109 drain_right.n210 drain_right.n186 104.615
R1110 drain_right.n210 drain_right.n209 104.615
R1111 drain_right.n209 drain_right.n191 104.615
R1112 drain_right.n202 drain_right.n191 104.615
R1113 drain_right.n202 drain_right.n201 104.615
R1114 drain_right.n201 drain_right.n195 104.615
R1115 drain_right.n143 drain_right.n141 59.6034
R1116 drain_right.n147 drain_right.n145 59.6032
R1117 drain_right.n143 drain_right.n142 58.7154
R1118 drain_right.n140 drain_right.n139 58.7154
R1119 drain_right.n147 drain_right.n146 58.7154
R1120 drain_right.n149 drain_right.n148 58.7154
R1121 drain_right.t8 drain_right.n43 52.3082
R1122 drain_right.t7 drain_right.n195 52.3082
R1123 drain_right.n140 drain_right.n138 48.2006
R1124 drain_right.n289 drain_right.n288 47.3126
R1125 drain_right drain_right.n144 41.7679
R1126 drain_right.n69 drain_right.n34 13.1884
R1127 drain_right.n116 drain_right.n115 13.1884
R1128 drain_right.n266 drain_right.n265 13.1884
R1129 drain_right.n220 drain_right.n185 13.1884
R1130 drain_right.n65 drain_right.n64 12.8005
R1131 drain_right.n70 drain_right.n32 12.8005
R1132 drain_right.n114 drain_right.n12 12.8005
R1133 drain_right.n119 drain_right.n10 12.8005
R1134 drain_right.n269 drain_right.n160 12.8005
R1135 drain_right.n264 drain_right.n162 12.8005
R1136 drain_right.n221 drain_right.n183 12.8005
R1137 drain_right.n216 drain_right.n187 12.8005
R1138 drain_right.n63 drain_right.n36 12.0247
R1139 drain_right.n74 drain_right.n73 12.0247
R1140 drain_right.n111 drain_right.n110 12.0247
R1141 drain_right.n120 drain_right.n8 12.0247
R1142 drain_right.n270 drain_right.n158 12.0247
R1143 drain_right.n261 drain_right.n260 12.0247
R1144 drain_right.n225 drain_right.n224 12.0247
R1145 drain_right.n215 drain_right.n188 12.0247
R1146 drain_right.n60 drain_right.n59 11.249
R1147 drain_right.n77 drain_right.n30 11.249
R1148 drain_right.n106 drain_right.n14 11.249
R1149 drain_right.n124 drain_right.n123 11.249
R1150 drain_right.n274 drain_right.n273 11.249
R1151 drain_right.n257 drain_right.n164 11.249
R1152 drain_right.n228 drain_right.n181 11.249
R1153 drain_right.n212 drain_right.n211 11.249
R1154 drain_right.n56 drain_right.n38 10.4732
R1155 drain_right.n78 drain_right.n28 10.4732
R1156 drain_right.n105 drain_right.n16 10.4732
R1157 drain_right.n127 drain_right.n6 10.4732
R1158 drain_right.n277 drain_right.n156 10.4732
R1159 drain_right.n256 drain_right.n167 10.4732
R1160 drain_right.n229 drain_right.n179 10.4732
R1161 drain_right.n208 drain_right.n190 10.4732
R1162 drain_right.n45 drain_right.n44 10.2747
R1163 drain_right.n197 drain_right.n196 10.2747
R1164 drain_right.n55 drain_right.n40 9.69747
R1165 drain_right.n82 drain_right.n81 9.69747
R1166 drain_right.n102 drain_right.n101 9.69747
R1167 drain_right.n128 drain_right.n4 9.69747
R1168 drain_right.n278 drain_right.n154 9.69747
R1169 drain_right.n253 drain_right.n252 9.69747
R1170 drain_right.n233 drain_right.n232 9.69747
R1171 drain_right.n207 drain_right.n192 9.69747
R1172 drain_right.n138 drain_right.n137 9.45567
R1173 drain_right.n288 drain_right.n287 9.45567
R1174 drain_right.n2 drain_right.n1 9.3005
R1175 drain_right.n131 drain_right.n130 9.3005
R1176 drain_right.n129 drain_right.n128 9.3005
R1177 drain_right.n6 drain_right.n5 9.3005
R1178 drain_right.n123 drain_right.n122 9.3005
R1179 drain_right.n121 drain_right.n120 9.3005
R1180 drain_right.n10 drain_right.n9 9.3005
R1181 drain_right.n89 drain_right.n88 9.3005
R1182 drain_right.n87 drain_right.n86 9.3005
R1183 drain_right.n26 drain_right.n25 9.3005
R1184 drain_right.n81 drain_right.n80 9.3005
R1185 drain_right.n79 drain_right.n78 9.3005
R1186 drain_right.n30 drain_right.n29 9.3005
R1187 drain_right.n73 drain_right.n72 9.3005
R1188 drain_right.n71 drain_right.n70 9.3005
R1189 drain_right.n47 drain_right.n46 9.3005
R1190 drain_right.n42 drain_right.n41 9.3005
R1191 drain_right.n53 drain_right.n52 9.3005
R1192 drain_right.n55 drain_right.n54 9.3005
R1193 drain_right.n38 drain_right.n37 9.3005
R1194 drain_right.n61 drain_right.n60 9.3005
R1195 drain_right.n63 drain_right.n62 9.3005
R1196 drain_right.n64 drain_right.n33 9.3005
R1197 drain_right.n22 drain_right.n21 9.3005
R1198 drain_right.n95 drain_right.n94 9.3005
R1199 drain_right.n97 drain_right.n96 9.3005
R1200 drain_right.n18 drain_right.n17 9.3005
R1201 drain_right.n103 drain_right.n102 9.3005
R1202 drain_right.n105 drain_right.n104 9.3005
R1203 drain_right.n14 drain_right.n13 9.3005
R1204 drain_right.n112 drain_right.n111 9.3005
R1205 drain_right.n114 drain_right.n113 9.3005
R1206 drain_right.n137 drain_right.n136 9.3005
R1207 drain_right.n199 drain_right.n198 9.3005
R1208 drain_right.n194 drain_right.n193 9.3005
R1209 drain_right.n205 drain_right.n204 9.3005
R1210 drain_right.n207 drain_right.n206 9.3005
R1211 drain_right.n190 drain_right.n189 9.3005
R1212 drain_right.n213 drain_right.n212 9.3005
R1213 drain_right.n215 drain_right.n214 9.3005
R1214 drain_right.n187 drain_right.n184 9.3005
R1215 drain_right.n246 drain_right.n245 9.3005
R1216 drain_right.n248 drain_right.n247 9.3005
R1217 drain_right.n169 drain_right.n168 9.3005
R1218 drain_right.n254 drain_right.n253 9.3005
R1219 drain_right.n256 drain_right.n255 9.3005
R1220 drain_right.n164 drain_right.n163 9.3005
R1221 drain_right.n262 drain_right.n261 9.3005
R1222 drain_right.n264 drain_right.n263 9.3005
R1223 drain_right.n287 drain_right.n286 9.3005
R1224 drain_right.n152 drain_right.n151 9.3005
R1225 drain_right.n281 drain_right.n280 9.3005
R1226 drain_right.n279 drain_right.n278 9.3005
R1227 drain_right.n156 drain_right.n155 9.3005
R1228 drain_right.n273 drain_right.n272 9.3005
R1229 drain_right.n271 drain_right.n270 9.3005
R1230 drain_right.n160 drain_right.n159 9.3005
R1231 drain_right.n173 drain_right.n172 9.3005
R1232 drain_right.n240 drain_right.n239 9.3005
R1233 drain_right.n238 drain_right.n237 9.3005
R1234 drain_right.n177 drain_right.n176 9.3005
R1235 drain_right.n232 drain_right.n231 9.3005
R1236 drain_right.n230 drain_right.n229 9.3005
R1237 drain_right.n181 drain_right.n180 9.3005
R1238 drain_right.n224 drain_right.n223 9.3005
R1239 drain_right.n222 drain_right.n221 9.3005
R1240 drain_right.n52 drain_right.n51 8.92171
R1241 drain_right.n85 drain_right.n26 8.92171
R1242 drain_right.n98 drain_right.n18 8.92171
R1243 drain_right.n132 drain_right.n131 8.92171
R1244 drain_right.n282 drain_right.n281 8.92171
R1245 drain_right.n249 drain_right.n169 8.92171
R1246 drain_right.n236 drain_right.n177 8.92171
R1247 drain_right.n204 drain_right.n203 8.92171
R1248 drain_right.n48 drain_right.n42 8.14595
R1249 drain_right.n86 drain_right.n24 8.14595
R1250 drain_right.n97 drain_right.n20 8.14595
R1251 drain_right.n135 drain_right.n2 8.14595
R1252 drain_right.n285 drain_right.n152 8.14595
R1253 drain_right.n248 drain_right.n171 8.14595
R1254 drain_right.n237 drain_right.n175 8.14595
R1255 drain_right.n200 drain_right.n194 8.14595
R1256 drain_right.n47 drain_right.n44 7.3702
R1257 drain_right.n90 drain_right.n89 7.3702
R1258 drain_right.n94 drain_right.n93 7.3702
R1259 drain_right.n136 drain_right.n0 7.3702
R1260 drain_right.n286 drain_right.n150 7.3702
R1261 drain_right.n245 drain_right.n244 7.3702
R1262 drain_right.n241 drain_right.n240 7.3702
R1263 drain_right.n199 drain_right.n196 7.3702
R1264 drain_right.n90 drain_right.n22 6.59444
R1265 drain_right.n93 drain_right.n22 6.59444
R1266 drain_right.n138 drain_right.n0 6.59444
R1267 drain_right.n288 drain_right.n150 6.59444
R1268 drain_right.n244 drain_right.n173 6.59444
R1269 drain_right.n241 drain_right.n173 6.59444
R1270 drain_right drain_right.n289 6.09718
R1271 drain_right.n48 drain_right.n47 5.81868
R1272 drain_right.n89 drain_right.n24 5.81868
R1273 drain_right.n94 drain_right.n20 5.81868
R1274 drain_right.n136 drain_right.n135 5.81868
R1275 drain_right.n286 drain_right.n285 5.81868
R1276 drain_right.n245 drain_right.n171 5.81868
R1277 drain_right.n240 drain_right.n175 5.81868
R1278 drain_right.n200 drain_right.n199 5.81868
R1279 drain_right.n51 drain_right.n42 5.04292
R1280 drain_right.n86 drain_right.n85 5.04292
R1281 drain_right.n98 drain_right.n97 5.04292
R1282 drain_right.n132 drain_right.n2 5.04292
R1283 drain_right.n282 drain_right.n152 5.04292
R1284 drain_right.n249 drain_right.n248 5.04292
R1285 drain_right.n237 drain_right.n236 5.04292
R1286 drain_right.n203 drain_right.n194 5.04292
R1287 drain_right.n52 drain_right.n40 4.26717
R1288 drain_right.n82 drain_right.n26 4.26717
R1289 drain_right.n101 drain_right.n18 4.26717
R1290 drain_right.n131 drain_right.n4 4.26717
R1291 drain_right.n281 drain_right.n154 4.26717
R1292 drain_right.n252 drain_right.n169 4.26717
R1293 drain_right.n233 drain_right.n177 4.26717
R1294 drain_right.n204 drain_right.n192 4.26717
R1295 drain_right.n56 drain_right.n55 3.49141
R1296 drain_right.n81 drain_right.n28 3.49141
R1297 drain_right.n102 drain_right.n16 3.49141
R1298 drain_right.n128 drain_right.n127 3.49141
R1299 drain_right.n278 drain_right.n277 3.49141
R1300 drain_right.n253 drain_right.n167 3.49141
R1301 drain_right.n232 drain_right.n179 3.49141
R1302 drain_right.n208 drain_right.n207 3.49141
R1303 drain_right.n198 drain_right.n197 2.84303
R1304 drain_right.n46 drain_right.n45 2.84303
R1305 drain_right.n59 drain_right.n38 2.71565
R1306 drain_right.n78 drain_right.n77 2.71565
R1307 drain_right.n106 drain_right.n105 2.71565
R1308 drain_right.n124 drain_right.n6 2.71565
R1309 drain_right.n274 drain_right.n156 2.71565
R1310 drain_right.n257 drain_right.n256 2.71565
R1311 drain_right.n229 drain_right.n228 2.71565
R1312 drain_right.n211 drain_right.n190 2.71565
R1313 drain_right.n60 drain_right.n36 1.93989
R1314 drain_right.n74 drain_right.n30 1.93989
R1315 drain_right.n110 drain_right.n14 1.93989
R1316 drain_right.n123 drain_right.n8 1.93989
R1317 drain_right.n273 drain_right.n158 1.93989
R1318 drain_right.n260 drain_right.n164 1.93989
R1319 drain_right.n225 drain_right.n181 1.93989
R1320 drain_right.n212 drain_right.n188 1.93989
R1321 drain_right.n65 drain_right.n63 1.16414
R1322 drain_right.n73 drain_right.n32 1.16414
R1323 drain_right.n111 drain_right.n12 1.16414
R1324 drain_right.n120 drain_right.n119 1.16414
R1325 drain_right.n270 drain_right.n269 1.16414
R1326 drain_right.n261 drain_right.n162 1.16414
R1327 drain_right.n224 drain_right.n183 1.16414
R1328 drain_right.n216 drain_right.n215 1.16414
R1329 drain_right.n289 drain_right.n149 0.888431
R1330 drain_right.n149 drain_right.n147 0.888431
R1331 drain_right.n141 drain_right.t3 0.7925
R1332 drain_right.n141 drain_right.t2 0.7925
R1333 drain_right.n142 drain_right.t12 0.7925
R1334 drain_right.n142 drain_right.t10 0.7925
R1335 drain_right.n139 drain_right.t9 0.7925
R1336 drain_right.n139 drain_right.t13 0.7925
R1337 drain_right.n145 drain_right.t11 0.7925
R1338 drain_right.n145 drain_right.t4 0.7925
R1339 drain_right.n146 drain_right.t1 0.7925
R1340 drain_right.n146 drain_right.t5 0.7925
R1341 drain_right.n148 drain_right.t0 0.7925
R1342 drain_right.n148 drain_right.t6 0.7925
R1343 drain_right.n144 drain_right.n140 0.611102
R1344 drain_right.n64 drain_right.n34 0.388379
R1345 drain_right.n70 drain_right.n69 0.388379
R1346 drain_right.n115 drain_right.n114 0.388379
R1347 drain_right.n116 drain_right.n10 0.388379
R1348 drain_right.n266 drain_right.n160 0.388379
R1349 drain_right.n265 drain_right.n264 0.388379
R1350 drain_right.n221 drain_right.n220 0.388379
R1351 drain_right.n187 drain_right.n185 0.388379
R1352 drain_right.n144 drain_right.n143 0.167137
R1353 drain_right.n46 drain_right.n41 0.155672
R1354 drain_right.n53 drain_right.n41 0.155672
R1355 drain_right.n54 drain_right.n53 0.155672
R1356 drain_right.n54 drain_right.n37 0.155672
R1357 drain_right.n61 drain_right.n37 0.155672
R1358 drain_right.n62 drain_right.n61 0.155672
R1359 drain_right.n62 drain_right.n33 0.155672
R1360 drain_right.n71 drain_right.n33 0.155672
R1361 drain_right.n72 drain_right.n71 0.155672
R1362 drain_right.n72 drain_right.n29 0.155672
R1363 drain_right.n79 drain_right.n29 0.155672
R1364 drain_right.n80 drain_right.n79 0.155672
R1365 drain_right.n80 drain_right.n25 0.155672
R1366 drain_right.n87 drain_right.n25 0.155672
R1367 drain_right.n88 drain_right.n87 0.155672
R1368 drain_right.n88 drain_right.n21 0.155672
R1369 drain_right.n95 drain_right.n21 0.155672
R1370 drain_right.n96 drain_right.n95 0.155672
R1371 drain_right.n96 drain_right.n17 0.155672
R1372 drain_right.n103 drain_right.n17 0.155672
R1373 drain_right.n104 drain_right.n103 0.155672
R1374 drain_right.n104 drain_right.n13 0.155672
R1375 drain_right.n112 drain_right.n13 0.155672
R1376 drain_right.n113 drain_right.n112 0.155672
R1377 drain_right.n113 drain_right.n9 0.155672
R1378 drain_right.n121 drain_right.n9 0.155672
R1379 drain_right.n122 drain_right.n121 0.155672
R1380 drain_right.n122 drain_right.n5 0.155672
R1381 drain_right.n129 drain_right.n5 0.155672
R1382 drain_right.n130 drain_right.n129 0.155672
R1383 drain_right.n130 drain_right.n1 0.155672
R1384 drain_right.n137 drain_right.n1 0.155672
R1385 drain_right.n287 drain_right.n151 0.155672
R1386 drain_right.n280 drain_right.n151 0.155672
R1387 drain_right.n280 drain_right.n279 0.155672
R1388 drain_right.n279 drain_right.n155 0.155672
R1389 drain_right.n272 drain_right.n155 0.155672
R1390 drain_right.n272 drain_right.n271 0.155672
R1391 drain_right.n271 drain_right.n159 0.155672
R1392 drain_right.n263 drain_right.n159 0.155672
R1393 drain_right.n263 drain_right.n262 0.155672
R1394 drain_right.n262 drain_right.n163 0.155672
R1395 drain_right.n255 drain_right.n163 0.155672
R1396 drain_right.n255 drain_right.n254 0.155672
R1397 drain_right.n254 drain_right.n168 0.155672
R1398 drain_right.n247 drain_right.n168 0.155672
R1399 drain_right.n247 drain_right.n246 0.155672
R1400 drain_right.n246 drain_right.n172 0.155672
R1401 drain_right.n239 drain_right.n172 0.155672
R1402 drain_right.n239 drain_right.n238 0.155672
R1403 drain_right.n238 drain_right.n176 0.155672
R1404 drain_right.n231 drain_right.n176 0.155672
R1405 drain_right.n231 drain_right.n230 0.155672
R1406 drain_right.n230 drain_right.n180 0.155672
R1407 drain_right.n223 drain_right.n180 0.155672
R1408 drain_right.n223 drain_right.n222 0.155672
R1409 drain_right.n222 drain_right.n184 0.155672
R1410 drain_right.n214 drain_right.n184 0.155672
R1411 drain_right.n214 drain_right.n213 0.155672
R1412 drain_right.n213 drain_right.n189 0.155672
R1413 drain_right.n206 drain_right.n189 0.155672
R1414 drain_right.n206 drain_right.n205 0.155672
R1415 drain_right.n205 drain_right.n193 0.155672
R1416 drain_right.n198 drain_right.n193 0.155672
R1417 plus.n5 plus.t5 940.679
R1418 plus.n27 plus.t13 940.679
R1419 plus.n20 plus.t1 916.833
R1420 plus.n18 plus.t10 916.833
R1421 plus.n2 plus.t4 916.833
R1422 plus.n12 plus.t8 916.833
R1423 plus.n4 plus.t2 916.833
R1424 plus.n6 plus.t11 916.833
R1425 plus.n42 plus.t6 916.833
R1426 plus.n40 plus.t3 916.833
R1427 plus.n24 plus.t9 916.833
R1428 plus.n34 plus.t7 916.833
R1429 plus.n26 plus.t12 916.833
R1430 plus.n28 plus.t0 916.833
R1431 plus.n8 plus.n7 161.3
R1432 plus.n9 plus.n4 161.3
R1433 plus.n11 plus.n10 161.3
R1434 plus.n12 plus.n3 161.3
R1435 plus.n14 plus.n13 161.3
R1436 plus.n15 plus.n2 161.3
R1437 plus.n17 plus.n16 161.3
R1438 plus.n18 plus.n1 161.3
R1439 plus.n19 plus.n0 161.3
R1440 plus.n21 plus.n20 161.3
R1441 plus.n30 plus.n29 161.3
R1442 plus.n31 plus.n26 161.3
R1443 plus.n33 plus.n32 161.3
R1444 plus.n34 plus.n25 161.3
R1445 plus.n36 plus.n35 161.3
R1446 plus.n37 plus.n24 161.3
R1447 plus.n39 plus.n38 161.3
R1448 plus.n40 plus.n23 161.3
R1449 plus.n41 plus.n22 161.3
R1450 plus.n43 plus.n42 161.3
R1451 plus.n30 plus.n27 44.9119
R1452 plus.n8 plus.n5 44.9119
R1453 plus plus.n43 37.0312
R1454 plus.n20 plus.n19 35.055
R1455 plus.n42 plus.n41 35.055
R1456 plus.n18 plus.n17 30.6732
R1457 plus.n7 plus.n6 30.6732
R1458 plus.n40 plus.n39 30.6732
R1459 plus.n29 plus.n28 30.6732
R1460 plus.n13 plus.n2 26.2914
R1461 plus.n11 plus.n4 26.2914
R1462 plus.n35 plus.n24 26.2914
R1463 plus.n33 plus.n26 26.2914
R1464 plus.n13 plus.n12 21.9096
R1465 plus.n12 plus.n11 21.9096
R1466 plus.n35 plus.n34 21.9096
R1467 plus.n34 plus.n33 21.9096
R1468 plus.n28 plus.n27 17.739
R1469 plus.n6 plus.n5 17.739
R1470 plus.n17 plus.n2 17.5278
R1471 plus.n7 plus.n4 17.5278
R1472 plus.n39 plus.n24 17.5278
R1473 plus.n29 plus.n26 17.5278
R1474 plus plus.n21 17.2183
R1475 plus.n19 plus.n18 13.146
R1476 plus.n41 plus.n40 13.146
R1477 plus.n9 plus.n8 0.189894
R1478 plus.n10 plus.n9 0.189894
R1479 plus.n10 plus.n3 0.189894
R1480 plus.n14 plus.n3 0.189894
R1481 plus.n15 plus.n14 0.189894
R1482 plus.n16 plus.n15 0.189894
R1483 plus.n16 plus.n1 0.189894
R1484 plus.n1 plus.n0 0.189894
R1485 plus.n21 plus.n0 0.189894
R1486 plus.n43 plus.n22 0.189894
R1487 plus.n23 plus.n22 0.189894
R1488 plus.n38 plus.n23 0.189894
R1489 plus.n38 plus.n37 0.189894
R1490 plus.n37 plus.n36 0.189894
R1491 plus.n36 plus.n25 0.189894
R1492 plus.n32 plus.n25 0.189894
R1493 plus.n32 plus.n31 0.189894
R1494 plus.n31 plus.n30 0.189894
R1495 drain_left.n134 drain_left.n0 289.615
R1496 drain_left.n279 drain_left.n145 289.615
R1497 drain_left.n44 drain_left.n43 185
R1498 drain_left.n49 drain_left.n48 185
R1499 drain_left.n51 drain_left.n50 185
R1500 drain_left.n40 drain_left.n39 185
R1501 drain_left.n57 drain_left.n56 185
R1502 drain_left.n59 drain_left.n58 185
R1503 drain_left.n36 drain_left.n35 185
R1504 drain_left.n66 drain_left.n65 185
R1505 drain_left.n67 drain_left.n34 185
R1506 drain_left.n69 drain_left.n68 185
R1507 drain_left.n32 drain_left.n31 185
R1508 drain_left.n75 drain_left.n74 185
R1509 drain_left.n77 drain_left.n76 185
R1510 drain_left.n28 drain_left.n27 185
R1511 drain_left.n83 drain_left.n82 185
R1512 drain_left.n85 drain_left.n84 185
R1513 drain_left.n24 drain_left.n23 185
R1514 drain_left.n91 drain_left.n90 185
R1515 drain_left.n93 drain_left.n92 185
R1516 drain_left.n20 drain_left.n19 185
R1517 drain_left.n99 drain_left.n98 185
R1518 drain_left.n101 drain_left.n100 185
R1519 drain_left.n16 drain_left.n15 185
R1520 drain_left.n107 drain_left.n106 185
R1521 drain_left.n110 drain_left.n109 185
R1522 drain_left.n108 drain_left.n12 185
R1523 drain_left.n115 drain_left.n11 185
R1524 drain_left.n117 drain_left.n116 185
R1525 drain_left.n119 drain_left.n118 185
R1526 drain_left.n8 drain_left.n7 185
R1527 drain_left.n125 drain_left.n124 185
R1528 drain_left.n127 drain_left.n126 185
R1529 drain_left.n4 drain_left.n3 185
R1530 drain_left.n133 drain_left.n132 185
R1531 drain_left.n135 drain_left.n134 185
R1532 drain_left.n280 drain_left.n279 185
R1533 drain_left.n278 drain_left.n277 185
R1534 drain_left.n149 drain_left.n148 185
R1535 drain_left.n272 drain_left.n271 185
R1536 drain_left.n270 drain_left.n269 185
R1537 drain_left.n153 drain_left.n152 185
R1538 drain_left.n264 drain_left.n263 185
R1539 drain_left.n262 drain_left.n261 185
R1540 drain_left.n260 drain_left.n156 185
R1541 drain_left.n160 drain_left.n157 185
R1542 drain_left.n255 drain_left.n254 185
R1543 drain_left.n253 drain_left.n252 185
R1544 drain_left.n162 drain_left.n161 185
R1545 drain_left.n247 drain_left.n246 185
R1546 drain_left.n245 drain_left.n244 185
R1547 drain_left.n166 drain_left.n165 185
R1548 drain_left.n239 drain_left.n238 185
R1549 drain_left.n237 drain_left.n236 185
R1550 drain_left.n170 drain_left.n169 185
R1551 drain_left.n231 drain_left.n230 185
R1552 drain_left.n229 drain_left.n228 185
R1553 drain_left.n174 drain_left.n173 185
R1554 drain_left.n223 drain_left.n222 185
R1555 drain_left.n221 drain_left.n220 185
R1556 drain_left.n178 drain_left.n177 185
R1557 drain_left.n215 drain_left.n214 185
R1558 drain_left.n213 drain_left.n180 185
R1559 drain_left.n212 drain_left.n211 185
R1560 drain_left.n183 drain_left.n181 185
R1561 drain_left.n206 drain_left.n205 185
R1562 drain_left.n204 drain_left.n203 185
R1563 drain_left.n187 drain_left.n186 185
R1564 drain_left.n198 drain_left.n197 185
R1565 drain_left.n196 drain_left.n195 185
R1566 drain_left.n191 drain_left.n190 185
R1567 drain_left.n45 drain_left.t7 149.524
R1568 drain_left.n192 drain_left.t8 149.524
R1569 drain_left.n49 drain_left.n43 104.615
R1570 drain_left.n50 drain_left.n49 104.615
R1571 drain_left.n50 drain_left.n39 104.615
R1572 drain_left.n57 drain_left.n39 104.615
R1573 drain_left.n58 drain_left.n57 104.615
R1574 drain_left.n58 drain_left.n35 104.615
R1575 drain_left.n66 drain_left.n35 104.615
R1576 drain_left.n67 drain_left.n66 104.615
R1577 drain_left.n68 drain_left.n67 104.615
R1578 drain_left.n68 drain_left.n31 104.615
R1579 drain_left.n75 drain_left.n31 104.615
R1580 drain_left.n76 drain_left.n75 104.615
R1581 drain_left.n76 drain_left.n27 104.615
R1582 drain_left.n83 drain_left.n27 104.615
R1583 drain_left.n84 drain_left.n83 104.615
R1584 drain_left.n84 drain_left.n23 104.615
R1585 drain_left.n91 drain_left.n23 104.615
R1586 drain_left.n92 drain_left.n91 104.615
R1587 drain_left.n92 drain_left.n19 104.615
R1588 drain_left.n99 drain_left.n19 104.615
R1589 drain_left.n100 drain_left.n99 104.615
R1590 drain_left.n100 drain_left.n15 104.615
R1591 drain_left.n107 drain_left.n15 104.615
R1592 drain_left.n109 drain_left.n107 104.615
R1593 drain_left.n109 drain_left.n108 104.615
R1594 drain_left.n108 drain_left.n11 104.615
R1595 drain_left.n117 drain_left.n11 104.615
R1596 drain_left.n118 drain_left.n117 104.615
R1597 drain_left.n118 drain_left.n7 104.615
R1598 drain_left.n125 drain_left.n7 104.615
R1599 drain_left.n126 drain_left.n125 104.615
R1600 drain_left.n126 drain_left.n3 104.615
R1601 drain_left.n133 drain_left.n3 104.615
R1602 drain_left.n134 drain_left.n133 104.615
R1603 drain_left.n279 drain_left.n278 104.615
R1604 drain_left.n278 drain_left.n148 104.615
R1605 drain_left.n271 drain_left.n148 104.615
R1606 drain_left.n271 drain_left.n270 104.615
R1607 drain_left.n270 drain_left.n152 104.615
R1608 drain_left.n263 drain_left.n152 104.615
R1609 drain_left.n263 drain_left.n262 104.615
R1610 drain_left.n262 drain_left.n156 104.615
R1611 drain_left.n160 drain_left.n156 104.615
R1612 drain_left.n254 drain_left.n160 104.615
R1613 drain_left.n254 drain_left.n253 104.615
R1614 drain_left.n253 drain_left.n161 104.615
R1615 drain_left.n246 drain_left.n161 104.615
R1616 drain_left.n246 drain_left.n245 104.615
R1617 drain_left.n245 drain_left.n165 104.615
R1618 drain_left.n238 drain_left.n165 104.615
R1619 drain_left.n238 drain_left.n237 104.615
R1620 drain_left.n237 drain_left.n169 104.615
R1621 drain_left.n230 drain_left.n169 104.615
R1622 drain_left.n230 drain_left.n229 104.615
R1623 drain_left.n229 drain_left.n173 104.615
R1624 drain_left.n222 drain_left.n173 104.615
R1625 drain_left.n222 drain_left.n221 104.615
R1626 drain_left.n221 drain_left.n177 104.615
R1627 drain_left.n214 drain_left.n177 104.615
R1628 drain_left.n214 drain_left.n213 104.615
R1629 drain_left.n213 drain_left.n212 104.615
R1630 drain_left.n212 drain_left.n181 104.615
R1631 drain_left.n205 drain_left.n181 104.615
R1632 drain_left.n205 drain_left.n204 104.615
R1633 drain_left.n204 drain_left.n186 104.615
R1634 drain_left.n197 drain_left.n186 104.615
R1635 drain_left.n197 drain_left.n196 104.615
R1636 drain_left.n196 drain_left.n190 104.615
R1637 drain_left.n143 drain_left.n141 59.6034
R1638 drain_left.n143 drain_left.n142 58.7154
R1639 drain_left.n140 drain_left.n139 58.7154
R1640 drain_left.n287 drain_left.n286 58.7154
R1641 drain_left.n285 drain_left.n284 58.7154
R1642 drain_left.n289 drain_left.n288 58.7153
R1643 drain_left.t7 drain_left.n43 52.3082
R1644 drain_left.t8 drain_left.n190 52.3082
R1645 drain_left.n140 drain_left.n138 48.2006
R1646 drain_left.n285 drain_left.n283 48.2006
R1647 drain_left drain_left.n144 42.3212
R1648 drain_left.n69 drain_left.n34 13.1884
R1649 drain_left.n116 drain_left.n115 13.1884
R1650 drain_left.n261 drain_left.n260 13.1884
R1651 drain_left.n215 drain_left.n180 13.1884
R1652 drain_left.n65 drain_left.n64 12.8005
R1653 drain_left.n70 drain_left.n32 12.8005
R1654 drain_left.n114 drain_left.n12 12.8005
R1655 drain_left.n119 drain_left.n10 12.8005
R1656 drain_left.n264 drain_left.n155 12.8005
R1657 drain_left.n259 drain_left.n157 12.8005
R1658 drain_left.n216 drain_left.n178 12.8005
R1659 drain_left.n211 drain_left.n182 12.8005
R1660 drain_left.n63 drain_left.n36 12.0247
R1661 drain_left.n74 drain_left.n73 12.0247
R1662 drain_left.n111 drain_left.n110 12.0247
R1663 drain_left.n120 drain_left.n8 12.0247
R1664 drain_left.n265 drain_left.n153 12.0247
R1665 drain_left.n256 drain_left.n255 12.0247
R1666 drain_left.n220 drain_left.n219 12.0247
R1667 drain_left.n210 drain_left.n183 12.0247
R1668 drain_left.n60 drain_left.n59 11.249
R1669 drain_left.n77 drain_left.n30 11.249
R1670 drain_left.n106 drain_left.n14 11.249
R1671 drain_left.n124 drain_left.n123 11.249
R1672 drain_left.n269 drain_left.n268 11.249
R1673 drain_left.n252 drain_left.n159 11.249
R1674 drain_left.n223 drain_left.n176 11.249
R1675 drain_left.n207 drain_left.n206 11.249
R1676 drain_left.n56 drain_left.n38 10.4732
R1677 drain_left.n78 drain_left.n28 10.4732
R1678 drain_left.n105 drain_left.n16 10.4732
R1679 drain_left.n127 drain_left.n6 10.4732
R1680 drain_left.n272 drain_left.n151 10.4732
R1681 drain_left.n251 drain_left.n162 10.4732
R1682 drain_left.n224 drain_left.n174 10.4732
R1683 drain_left.n203 drain_left.n185 10.4732
R1684 drain_left.n45 drain_left.n44 10.2747
R1685 drain_left.n192 drain_left.n191 10.2747
R1686 drain_left.n55 drain_left.n40 9.69747
R1687 drain_left.n82 drain_left.n81 9.69747
R1688 drain_left.n102 drain_left.n101 9.69747
R1689 drain_left.n128 drain_left.n4 9.69747
R1690 drain_left.n273 drain_left.n149 9.69747
R1691 drain_left.n248 drain_left.n247 9.69747
R1692 drain_left.n228 drain_left.n227 9.69747
R1693 drain_left.n202 drain_left.n187 9.69747
R1694 drain_left.n138 drain_left.n137 9.45567
R1695 drain_left.n283 drain_left.n282 9.45567
R1696 drain_left.n2 drain_left.n1 9.3005
R1697 drain_left.n131 drain_left.n130 9.3005
R1698 drain_left.n129 drain_left.n128 9.3005
R1699 drain_left.n6 drain_left.n5 9.3005
R1700 drain_left.n123 drain_left.n122 9.3005
R1701 drain_left.n121 drain_left.n120 9.3005
R1702 drain_left.n10 drain_left.n9 9.3005
R1703 drain_left.n89 drain_left.n88 9.3005
R1704 drain_left.n87 drain_left.n86 9.3005
R1705 drain_left.n26 drain_left.n25 9.3005
R1706 drain_left.n81 drain_left.n80 9.3005
R1707 drain_left.n79 drain_left.n78 9.3005
R1708 drain_left.n30 drain_left.n29 9.3005
R1709 drain_left.n73 drain_left.n72 9.3005
R1710 drain_left.n71 drain_left.n70 9.3005
R1711 drain_left.n47 drain_left.n46 9.3005
R1712 drain_left.n42 drain_left.n41 9.3005
R1713 drain_left.n53 drain_left.n52 9.3005
R1714 drain_left.n55 drain_left.n54 9.3005
R1715 drain_left.n38 drain_left.n37 9.3005
R1716 drain_left.n61 drain_left.n60 9.3005
R1717 drain_left.n63 drain_left.n62 9.3005
R1718 drain_left.n64 drain_left.n33 9.3005
R1719 drain_left.n22 drain_left.n21 9.3005
R1720 drain_left.n95 drain_left.n94 9.3005
R1721 drain_left.n97 drain_left.n96 9.3005
R1722 drain_left.n18 drain_left.n17 9.3005
R1723 drain_left.n103 drain_left.n102 9.3005
R1724 drain_left.n105 drain_left.n104 9.3005
R1725 drain_left.n14 drain_left.n13 9.3005
R1726 drain_left.n112 drain_left.n111 9.3005
R1727 drain_left.n114 drain_left.n113 9.3005
R1728 drain_left.n137 drain_left.n136 9.3005
R1729 drain_left.n194 drain_left.n193 9.3005
R1730 drain_left.n189 drain_left.n188 9.3005
R1731 drain_left.n200 drain_left.n199 9.3005
R1732 drain_left.n202 drain_left.n201 9.3005
R1733 drain_left.n185 drain_left.n184 9.3005
R1734 drain_left.n208 drain_left.n207 9.3005
R1735 drain_left.n210 drain_left.n209 9.3005
R1736 drain_left.n182 drain_left.n179 9.3005
R1737 drain_left.n241 drain_left.n240 9.3005
R1738 drain_left.n243 drain_left.n242 9.3005
R1739 drain_left.n164 drain_left.n163 9.3005
R1740 drain_left.n249 drain_left.n248 9.3005
R1741 drain_left.n251 drain_left.n250 9.3005
R1742 drain_left.n159 drain_left.n158 9.3005
R1743 drain_left.n257 drain_left.n256 9.3005
R1744 drain_left.n259 drain_left.n258 9.3005
R1745 drain_left.n282 drain_left.n281 9.3005
R1746 drain_left.n147 drain_left.n146 9.3005
R1747 drain_left.n276 drain_left.n275 9.3005
R1748 drain_left.n274 drain_left.n273 9.3005
R1749 drain_left.n151 drain_left.n150 9.3005
R1750 drain_left.n268 drain_left.n267 9.3005
R1751 drain_left.n266 drain_left.n265 9.3005
R1752 drain_left.n155 drain_left.n154 9.3005
R1753 drain_left.n168 drain_left.n167 9.3005
R1754 drain_left.n235 drain_left.n234 9.3005
R1755 drain_left.n233 drain_left.n232 9.3005
R1756 drain_left.n172 drain_left.n171 9.3005
R1757 drain_left.n227 drain_left.n226 9.3005
R1758 drain_left.n225 drain_left.n224 9.3005
R1759 drain_left.n176 drain_left.n175 9.3005
R1760 drain_left.n219 drain_left.n218 9.3005
R1761 drain_left.n217 drain_left.n216 9.3005
R1762 drain_left.n52 drain_left.n51 8.92171
R1763 drain_left.n85 drain_left.n26 8.92171
R1764 drain_left.n98 drain_left.n18 8.92171
R1765 drain_left.n132 drain_left.n131 8.92171
R1766 drain_left.n277 drain_left.n276 8.92171
R1767 drain_left.n244 drain_left.n164 8.92171
R1768 drain_left.n231 drain_left.n172 8.92171
R1769 drain_left.n199 drain_left.n198 8.92171
R1770 drain_left.n48 drain_left.n42 8.14595
R1771 drain_left.n86 drain_left.n24 8.14595
R1772 drain_left.n97 drain_left.n20 8.14595
R1773 drain_left.n135 drain_left.n2 8.14595
R1774 drain_left.n280 drain_left.n147 8.14595
R1775 drain_left.n243 drain_left.n166 8.14595
R1776 drain_left.n232 drain_left.n170 8.14595
R1777 drain_left.n195 drain_left.n189 8.14595
R1778 drain_left.n47 drain_left.n44 7.3702
R1779 drain_left.n90 drain_left.n89 7.3702
R1780 drain_left.n94 drain_left.n93 7.3702
R1781 drain_left.n136 drain_left.n0 7.3702
R1782 drain_left.n281 drain_left.n145 7.3702
R1783 drain_left.n240 drain_left.n239 7.3702
R1784 drain_left.n236 drain_left.n235 7.3702
R1785 drain_left.n194 drain_left.n191 7.3702
R1786 drain_left.n90 drain_left.n22 6.59444
R1787 drain_left.n93 drain_left.n22 6.59444
R1788 drain_left.n138 drain_left.n0 6.59444
R1789 drain_left.n283 drain_left.n145 6.59444
R1790 drain_left.n239 drain_left.n168 6.59444
R1791 drain_left.n236 drain_left.n168 6.59444
R1792 drain_left drain_left.n289 6.54115
R1793 drain_left.n48 drain_left.n47 5.81868
R1794 drain_left.n89 drain_left.n24 5.81868
R1795 drain_left.n94 drain_left.n20 5.81868
R1796 drain_left.n136 drain_left.n135 5.81868
R1797 drain_left.n281 drain_left.n280 5.81868
R1798 drain_left.n240 drain_left.n166 5.81868
R1799 drain_left.n235 drain_left.n170 5.81868
R1800 drain_left.n195 drain_left.n194 5.81868
R1801 drain_left.n51 drain_left.n42 5.04292
R1802 drain_left.n86 drain_left.n85 5.04292
R1803 drain_left.n98 drain_left.n97 5.04292
R1804 drain_left.n132 drain_left.n2 5.04292
R1805 drain_left.n277 drain_left.n147 5.04292
R1806 drain_left.n244 drain_left.n243 5.04292
R1807 drain_left.n232 drain_left.n231 5.04292
R1808 drain_left.n198 drain_left.n189 5.04292
R1809 drain_left.n52 drain_left.n40 4.26717
R1810 drain_left.n82 drain_left.n26 4.26717
R1811 drain_left.n101 drain_left.n18 4.26717
R1812 drain_left.n131 drain_left.n4 4.26717
R1813 drain_left.n276 drain_left.n149 4.26717
R1814 drain_left.n247 drain_left.n164 4.26717
R1815 drain_left.n228 drain_left.n172 4.26717
R1816 drain_left.n199 drain_left.n187 4.26717
R1817 drain_left.n56 drain_left.n55 3.49141
R1818 drain_left.n81 drain_left.n28 3.49141
R1819 drain_left.n102 drain_left.n16 3.49141
R1820 drain_left.n128 drain_left.n127 3.49141
R1821 drain_left.n273 drain_left.n272 3.49141
R1822 drain_left.n248 drain_left.n162 3.49141
R1823 drain_left.n227 drain_left.n174 3.49141
R1824 drain_left.n203 drain_left.n202 3.49141
R1825 drain_left.n193 drain_left.n192 2.84303
R1826 drain_left.n46 drain_left.n45 2.84303
R1827 drain_left.n59 drain_left.n38 2.71565
R1828 drain_left.n78 drain_left.n77 2.71565
R1829 drain_left.n106 drain_left.n105 2.71565
R1830 drain_left.n124 drain_left.n6 2.71565
R1831 drain_left.n269 drain_left.n151 2.71565
R1832 drain_left.n252 drain_left.n251 2.71565
R1833 drain_left.n224 drain_left.n223 2.71565
R1834 drain_left.n206 drain_left.n185 2.71565
R1835 drain_left.n60 drain_left.n36 1.93989
R1836 drain_left.n74 drain_left.n30 1.93989
R1837 drain_left.n110 drain_left.n14 1.93989
R1838 drain_left.n123 drain_left.n8 1.93989
R1839 drain_left.n268 drain_left.n153 1.93989
R1840 drain_left.n255 drain_left.n159 1.93989
R1841 drain_left.n220 drain_left.n176 1.93989
R1842 drain_left.n207 drain_left.n183 1.93989
R1843 drain_left.n65 drain_left.n63 1.16414
R1844 drain_left.n73 drain_left.n32 1.16414
R1845 drain_left.n111 drain_left.n12 1.16414
R1846 drain_left.n120 drain_left.n119 1.16414
R1847 drain_left.n265 drain_left.n264 1.16414
R1848 drain_left.n256 drain_left.n157 1.16414
R1849 drain_left.n219 drain_left.n178 1.16414
R1850 drain_left.n211 drain_left.n210 1.16414
R1851 drain_left.n287 drain_left.n285 0.888431
R1852 drain_left.n289 drain_left.n287 0.888431
R1853 drain_left.n141 drain_left.t13 0.7925
R1854 drain_left.n141 drain_left.t0 0.7925
R1855 drain_left.n142 drain_left.t6 0.7925
R1856 drain_left.n142 drain_left.t1 0.7925
R1857 drain_left.n139 drain_left.t10 0.7925
R1858 drain_left.n139 drain_left.t4 0.7925
R1859 drain_left.n288 drain_left.t3 0.7925
R1860 drain_left.n288 drain_left.t12 0.7925
R1861 drain_left.n286 drain_left.t5 0.7925
R1862 drain_left.n286 drain_left.t9 0.7925
R1863 drain_left.n284 drain_left.t2 0.7925
R1864 drain_left.n284 drain_left.t11 0.7925
R1865 drain_left.n144 drain_left.n140 0.611102
R1866 drain_left.n64 drain_left.n34 0.388379
R1867 drain_left.n70 drain_left.n69 0.388379
R1868 drain_left.n115 drain_left.n114 0.388379
R1869 drain_left.n116 drain_left.n10 0.388379
R1870 drain_left.n261 drain_left.n155 0.388379
R1871 drain_left.n260 drain_left.n259 0.388379
R1872 drain_left.n216 drain_left.n215 0.388379
R1873 drain_left.n182 drain_left.n180 0.388379
R1874 drain_left.n144 drain_left.n143 0.167137
R1875 drain_left.n46 drain_left.n41 0.155672
R1876 drain_left.n53 drain_left.n41 0.155672
R1877 drain_left.n54 drain_left.n53 0.155672
R1878 drain_left.n54 drain_left.n37 0.155672
R1879 drain_left.n61 drain_left.n37 0.155672
R1880 drain_left.n62 drain_left.n61 0.155672
R1881 drain_left.n62 drain_left.n33 0.155672
R1882 drain_left.n71 drain_left.n33 0.155672
R1883 drain_left.n72 drain_left.n71 0.155672
R1884 drain_left.n72 drain_left.n29 0.155672
R1885 drain_left.n79 drain_left.n29 0.155672
R1886 drain_left.n80 drain_left.n79 0.155672
R1887 drain_left.n80 drain_left.n25 0.155672
R1888 drain_left.n87 drain_left.n25 0.155672
R1889 drain_left.n88 drain_left.n87 0.155672
R1890 drain_left.n88 drain_left.n21 0.155672
R1891 drain_left.n95 drain_left.n21 0.155672
R1892 drain_left.n96 drain_left.n95 0.155672
R1893 drain_left.n96 drain_left.n17 0.155672
R1894 drain_left.n103 drain_left.n17 0.155672
R1895 drain_left.n104 drain_left.n103 0.155672
R1896 drain_left.n104 drain_left.n13 0.155672
R1897 drain_left.n112 drain_left.n13 0.155672
R1898 drain_left.n113 drain_left.n112 0.155672
R1899 drain_left.n113 drain_left.n9 0.155672
R1900 drain_left.n121 drain_left.n9 0.155672
R1901 drain_left.n122 drain_left.n121 0.155672
R1902 drain_left.n122 drain_left.n5 0.155672
R1903 drain_left.n129 drain_left.n5 0.155672
R1904 drain_left.n130 drain_left.n129 0.155672
R1905 drain_left.n130 drain_left.n1 0.155672
R1906 drain_left.n137 drain_left.n1 0.155672
R1907 drain_left.n282 drain_left.n146 0.155672
R1908 drain_left.n275 drain_left.n146 0.155672
R1909 drain_left.n275 drain_left.n274 0.155672
R1910 drain_left.n274 drain_left.n150 0.155672
R1911 drain_left.n267 drain_left.n150 0.155672
R1912 drain_left.n267 drain_left.n266 0.155672
R1913 drain_left.n266 drain_left.n154 0.155672
R1914 drain_left.n258 drain_left.n154 0.155672
R1915 drain_left.n258 drain_left.n257 0.155672
R1916 drain_left.n257 drain_left.n158 0.155672
R1917 drain_left.n250 drain_left.n158 0.155672
R1918 drain_left.n250 drain_left.n249 0.155672
R1919 drain_left.n249 drain_left.n163 0.155672
R1920 drain_left.n242 drain_left.n163 0.155672
R1921 drain_left.n242 drain_left.n241 0.155672
R1922 drain_left.n241 drain_left.n167 0.155672
R1923 drain_left.n234 drain_left.n167 0.155672
R1924 drain_left.n234 drain_left.n233 0.155672
R1925 drain_left.n233 drain_left.n171 0.155672
R1926 drain_left.n226 drain_left.n171 0.155672
R1927 drain_left.n226 drain_left.n225 0.155672
R1928 drain_left.n225 drain_left.n175 0.155672
R1929 drain_left.n218 drain_left.n175 0.155672
R1930 drain_left.n218 drain_left.n217 0.155672
R1931 drain_left.n217 drain_left.n179 0.155672
R1932 drain_left.n209 drain_left.n179 0.155672
R1933 drain_left.n209 drain_left.n208 0.155672
R1934 drain_left.n208 drain_left.n184 0.155672
R1935 drain_left.n201 drain_left.n184 0.155672
R1936 drain_left.n201 drain_left.n200 0.155672
R1937 drain_left.n200 drain_left.n188 0.155672
R1938 drain_left.n193 drain_left.n188 0.155672
C0 minus plus 8.49988f
C1 minus drain_right 18.3027f
C2 minus drain_left 0.172675f
C3 plus drain_right 0.392997f
C4 plus drain_left 18.531f
C5 source minus 17.7545f
C6 drain_right drain_left 1.23802f
C7 source plus 17.7696f
C8 source drain_right 35.3426f
C9 source drain_left 35.3571f
C10 drain_right a_n2364_n5888# 11.097919f
C11 drain_left a_n2364_n5888# 11.452529f
C12 source a_n2364_n5888# 11.392332f
C13 minus a_n2364_n5888# 10.258803f
C14 plus a_n2364_n5888# 12.63372f
C15 drain_left.n0 a_n2364_n5888# 0.034436f
C16 drain_left.n1 a_n2364_n5888# 0.024979f
C17 drain_left.n2 a_n2364_n5888# 0.013423f
C18 drain_left.n3 a_n2364_n5888# 0.031726f
C19 drain_left.n4 a_n2364_n5888# 0.014212f
C20 drain_left.n5 a_n2364_n5888# 0.024979f
C21 drain_left.n6 a_n2364_n5888# 0.013423f
C22 drain_left.n7 a_n2364_n5888# 0.031726f
C23 drain_left.n8 a_n2364_n5888# 0.014212f
C24 drain_left.n9 a_n2364_n5888# 0.024979f
C25 drain_left.n10 a_n2364_n5888# 0.013423f
C26 drain_left.n11 a_n2364_n5888# 0.031726f
C27 drain_left.n12 a_n2364_n5888# 0.014212f
C28 drain_left.n13 a_n2364_n5888# 0.024979f
C29 drain_left.n14 a_n2364_n5888# 0.013423f
C30 drain_left.n15 a_n2364_n5888# 0.031726f
C31 drain_left.n16 a_n2364_n5888# 0.014212f
C32 drain_left.n17 a_n2364_n5888# 0.024979f
C33 drain_left.n18 a_n2364_n5888# 0.013423f
C34 drain_left.n19 a_n2364_n5888# 0.031726f
C35 drain_left.n20 a_n2364_n5888# 0.014212f
C36 drain_left.n21 a_n2364_n5888# 0.024979f
C37 drain_left.n22 a_n2364_n5888# 0.013423f
C38 drain_left.n23 a_n2364_n5888# 0.031726f
C39 drain_left.n24 a_n2364_n5888# 0.014212f
C40 drain_left.n25 a_n2364_n5888# 0.024979f
C41 drain_left.n26 a_n2364_n5888# 0.013423f
C42 drain_left.n27 a_n2364_n5888# 0.031726f
C43 drain_left.n28 a_n2364_n5888# 0.014212f
C44 drain_left.n29 a_n2364_n5888# 0.024979f
C45 drain_left.n30 a_n2364_n5888# 0.013423f
C46 drain_left.n31 a_n2364_n5888# 0.031726f
C47 drain_left.n32 a_n2364_n5888# 0.014212f
C48 drain_left.n33 a_n2364_n5888# 0.024979f
C49 drain_left.n34 a_n2364_n5888# 0.013818f
C50 drain_left.n35 a_n2364_n5888# 0.031726f
C51 drain_left.n36 a_n2364_n5888# 0.014212f
C52 drain_left.n37 a_n2364_n5888# 0.024979f
C53 drain_left.n38 a_n2364_n5888# 0.013423f
C54 drain_left.n39 a_n2364_n5888# 0.031726f
C55 drain_left.n40 a_n2364_n5888# 0.014212f
C56 drain_left.n41 a_n2364_n5888# 0.024979f
C57 drain_left.n42 a_n2364_n5888# 0.013423f
C58 drain_left.n43 a_n2364_n5888# 0.023795f
C59 drain_left.n44 a_n2364_n5888# 0.022428f
C60 drain_left.t7 a_n2364_n5888# 0.055333f
C61 drain_left.n45 a_n2364_n5888# 0.304767f
C62 drain_left.n46 a_n2364_n5888# 2.7045f
C63 drain_left.n47 a_n2364_n5888# 0.013423f
C64 drain_left.n48 a_n2364_n5888# 0.014212f
C65 drain_left.n49 a_n2364_n5888# 0.031726f
C66 drain_left.n50 a_n2364_n5888# 0.031726f
C67 drain_left.n51 a_n2364_n5888# 0.014212f
C68 drain_left.n52 a_n2364_n5888# 0.013423f
C69 drain_left.n53 a_n2364_n5888# 0.024979f
C70 drain_left.n54 a_n2364_n5888# 0.024979f
C71 drain_left.n55 a_n2364_n5888# 0.013423f
C72 drain_left.n56 a_n2364_n5888# 0.014212f
C73 drain_left.n57 a_n2364_n5888# 0.031726f
C74 drain_left.n58 a_n2364_n5888# 0.031726f
C75 drain_left.n59 a_n2364_n5888# 0.014212f
C76 drain_left.n60 a_n2364_n5888# 0.013423f
C77 drain_left.n61 a_n2364_n5888# 0.024979f
C78 drain_left.n62 a_n2364_n5888# 0.024979f
C79 drain_left.n63 a_n2364_n5888# 0.013423f
C80 drain_left.n64 a_n2364_n5888# 0.013423f
C81 drain_left.n65 a_n2364_n5888# 0.014212f
C82 drain_left.n66 a_n2364_n5888# 0.031726f
C83 drain_left.n67 a_n2364_n5888# 0.031726f
C84 drain_left.n68 a_n2364_n5888# 0.031726f
C85 drain_left.n69 a_n2364_n5888# 0.013818f
C86 drain_left.n70 a_n2364_n5888# 0.013423f
C87 drain_left.n71 a_n2364_n5888# 0.024979f
C88 drain_left.n72 a_n2364_n5888# 0.024979f
C89 drain_left.n73 a_n2364_n5888# 0.013423f
C90 drain_left.n74 a_n2364_n5888# 0.014212f
C91 drain_left.n75 a_n2364_n5888# 0.031726f
C92 drain_left.n76 a_n2364_n5888# 0.031726f
C93 drain_left.n77 a_n2364_n5888# 0.014212f
C94 drain_left.n78 a_n2364_n5888# 0.013423f
C95 drain_left.n79 a_n2364_n5888# 0.024979f
C96 drain_left.n80 a_n2364_n5888# 0.024979f
C97 drain_left.n81 a_n2364_n5888# 0.013423f
C98 drain_left.n82 a_n2364_n5888# 0.014212f
C99 drain_left.n83 a_n2364_n5888# 0.031726f
C100 drain_left.n84 a_n2364_n5888# 0.031726f
C101 drain_left.n85 a_n2364_n5888# 0.014212f
C102 drain_left.n86 a_n2364_n5888# 0.013423f
C103 drain_left.n87 a_n2364_n5888# 0.024979f
C104 drain_left.n88 a_n2364_n5888# 0.024979f
C105 drain_left.n89 a_n2364_n5888# 0.013423f
C106 drain_left.n90 a_n2364_n5888# 0.014212f
C107 drain_left.n91 a_n2364_n5888# 0.031726f
C108 drain_left.n92 a_n2364_n5888# 0.031726f
C109 drain_left.n93 a_n2364_n5888# 0.014212f
C110 drain_left.n94 a_n2364_n5888# 0.013423f
C111 drain_left.n95 a_n2364_n5888# 0.024979f
C112 drain_left.n96 a_n2364_n5888# 0.024979f
C113 drain_left.n97 a_n2364_n5888# 0.013423f
C114 drain_left.n98 a_n2364_n5888# 0.014212f
C115 drain_left.n99 a_n2364_n5888# 0.031726f
C116 drain_left.n100 a_n2364_n5888# 0.031726f
C117 drain_left.n101 a_n2364_n5888# 0.014212f
C118 drain_left.n102 a_n2364_n5888# 0.013423f
C119 drain_left.n103 a_n2364_n5888# 0.024979f
C120 drain_left.n104 a_n2364_n5888# 0.024979f
C121 drain_left.n105 a_n2364_n5888# 0.013423f
C122 drain_left.n106 a_n2364_n5888# 0.014212f
C123 drain_left.n107 a_n2364_n5888# 0.031726f
C124 drain_left.n108 a_n2364_n5888# 0.031726f
C125 drain_left.n109 a_n2364_n5888# 0.031726f
C126 drain_left.n110 a_n2364_n5888# 0.014212f
C127 drain_left.n111 a_n2364_n5888# 0.013423f
C128 drain_left.n112 a_n2364_n5888# 0.024979f
C129 drain_left.n113 a_n2364_n5888# 0.024979f
C130 drain_left.n114 a_n2364_n5888# 0.013423f
C131 drain_left.n115 a_n2364_n5888# 0.013818f
C132 drain_left.n116 a_n2364_n5888# 0.013818f
C133 drain_left.n117 a_n2364_n5888# 0.031726f
C134 drain_left.n118 a_n2364_n5888# 0.031726f
C135 drain_left.n119 a_n2364_n5888# 0.014212f
C136 drain_left.n120 a_n2364_n5888# 0.013423f
C137 drain_left.n121 a_n2364_n5888# 0.024979f
C138 drain_left.n122 a_n2364_n5888# 0.024979f
C139 drain_left.n123 a_n2364_n5888# 0.013423f
C140 drain_left.n124 a_n2364_n5888# 0.014212f
C141 drain_left.n125 a_n2364_n5888# 0.031726f
C142 drain_left.n126 a_n2364_n5888# 0.031726f
C143 drain_left.n127 a_n2364_n5888# 0.014212f
C144 drain_left.n128 a_n2364_n5888# 0.013423f
C145 drain_left.n129 a_n2364_n5888# 0.024979f
C146 drain_left.n130 a_n2364_n5888# 0.024979f
C147 drain_left.n131 a_n2364_n5888# 0.013423f
C148 drain_left.n132 a_n2364_n5888# 0.014212f
C149 drain_left.n133 a_n2364_n5888# 0.031726f
C150 drain_left.n134 a_n2364_n5888# 0.06749f
C151 drain_left.n135 a_n2364_n5888# 0.014212f
C152 drain_left.n136 a_n2364_n5888# 0.013423f
C153 drain_left.n137 a_n2364_n5888# 0.055008f
C154 drain_left.n138 a_n2364_n5888# 0.057f
C155 drain_left.t10 a_n2364_n5888# 0.493482f
C156 drain_left.t4 a_n2364_n5888# 0.493482f
C157 drain_left.n139 a_n2364_n5888# 4.54797f
C158 drain_left.n140 a_n2364_n5888# 0.448541f
C159 drain_left.t13 a_n2364_n5888# 0.493482f
C160 drain_left.t0 a_n2364_n5888# 0.493482f
C161 drain_left.n141 a_n2364_n5888# 4.5534f
C162 drain_left.t6 a_n2364_n5888# 0.493482f
C163 drain_left.t1 a_n2364_n5888# 0.493482f
C164 drain_left.n142 a_n2364_n5888# 4.54797f
C165 drain_left.n143 a_n2364_n5888# 0.658221f
C166 drain_left.n144 a_n2364_n5888# 2.19758f
C167 drain_left.n145 a_n2364_n5888# 0.034436f
C168 drain_left.n146 a_n2364_n5888# 0.024979f
C169 drain_left.n147 a_n2364_n5888# 0.013423f
C170 drain_left.n148 a_n2364_n5888# 0.031726f
C171 drain_left.n149 a_n2364_n5888# 0.014212f
C172 drain_left.n150 a_n2364_n5888# 0.024979f
C173 drain_left.n151 a_n2364_n5888# 0.013423f
C174 drain_left.n152 a_n2364_n5888# 0.031726f
C175 drain_left.n153 a_n2364_n5888# 0.014212f
C176 drain_left.n154 a_n2364_n5888# 0.024979f
C177 drain_left.n155 a_n2364_n5888# 0.013423f
C178 drain_left.n156 a_n2364_n5888# 0.031726f
C179 drain_left.n157 a_n2364_n5888# 0.014212f
C180 drain_left.n158 a_n2364_n5888# 0.024979f
C181 drain_left.n159 a_n2364_n5888# 0.013423f
C182 drain_left.n160 a_n2364_n5888# 0.031726f
C183 drain_left.n161 a_n2364_n5888# 0.031726f
C184 drain_left.n162 a_n2364_n5888# 0.014212f
C185 drain_left.n163 a_n2364_n5888# 0.024979f
C186 drain_left.n164 a_n2364_n5888# 0.013423f
C187 drain_left.n165 a_n2364_n5888# 0.031726f
C188 drain_left.n166 a_n2364_n5888# 0.014212f
C189 drain_left.n167 a_n2364_n5888# 0.024979f
C190 drain_left.n168 a_n2364_n5888# 0.013423f
C191 drain_left.n169 a_n2364_n5888# 0.031726f
C192 drain_left.n170 a_n2364_n5888# 0.014212f
C193 drain_left.n171 a_n2364_n5888# 0.024979f
C194 drain_left.n172 a_n2364_n5888# 0.013423f
C195 drain_left.n173 a_n2364_n5888# 0.031726f
C196 drain_left.n174 a_n2364_n5888# 0.014212f
C197 drain_left.n175 a_n2364_n5888# 0.024979f
C198 drain_left.n176 a_n2364_n5888# 0.013423f
C199 drain_left.n177 a_n2364_n5888# 0.031726f
C200 drain_left.n178 a_n2364_n5888# 0.014212f
C201 drain_left.n179 a_n2364_n5888# 0.024979f
C202 drain_left.n180 a_n2364_n5888# 0.013818f
C203 drain_left.n181 a_n2364_n5888# 0.031726f
C204 drain_left.n182 a_n2364_n5888# 0.013423f
C205 drain_left.n183 a_n2364_n5888# 0.014212f
C206 drain_left.n184 a_n2364_n5888# 0.024979f
C207 drain_left.n185 a_n2364_n5888# 0.013423f
C208 drain_left.n186 a_n2364_n5888# 0.031726f
C209 drain_left.n187 a_n2364_n5888# 0.014212f
C210 drain_left.n188 a_n2364_n5888# 0.024979f
C211 drain_left.n189 a_n2364_n5888# 0.013423f
C212 drain_left.n190 a_n2364_n5888# 0.023795f
C213 drain_left.n191 a_n2364_n5888# 0.022428f
C214 drain_left.t8 a_n2364_n5888# 0.055333f
C215 drain_left.n192 a_n2364_n5888# 0.304767f
C216 drain_left.n193 a_n2364_n5888# 2.7045f
C217 drain_left.n194 a_n2364_n5888# 0.013423f
C218 drain_left.n195 a_n2364_n5888# 0.014212f
C219 drain_left.n196 a_n2364_n5888# 0.031726f
C220 drain_left.n197 a_n2364_n5888# 0.031726f
C221 drain_left.n198 a_n2364_n5888# 0.014212f
C222 drain_left.n199 a_n2364_n5888# 0.013423f
C223 drain_left.n200 a_n2364_n5888# 0.024979f
C224 drain_left.n201 a_n2364_n5888# 0.024979f
C225 drain_left.n202 a_n2364_n5888# 0.013423f
C226 drain_left.n203 a_n2364_n5888# 0.014212f
C227 drain_left.n204 a_n2364_n5888# 0.031726f
C228 drain_left.n205 a_n2364_n5888# 0.031726f
C229 drain_left.n206 a_n2364_n5888# 0.014212f
C230 drain_left.n207 a_n2364_n5888# 0.013423f
C231 drain_left.n208 a_n2364_n5888# 0.024979f
C232 drain_left.n209 a_n2364_n5888# 0.024979f
C233 drain_left.n210 a_n2364_n5888# 0.013423f
C234 drain_left.n211 a_n2364_n5888# 0.014212f
C235 drain_left.n212 a_n2364_n5888# 0.031726f
C236 drain_left.n213 a_n2364_n5888# 0.031726f
C237 drain_left.n214 a_n2364_n5888# 0.031726f
C238 drain_left.n215 a_n2364_n5888# 0.013818f
C239 drain_left.n216 a_n2364_n5888# 0.013423f
C240 drain_left.n217 a_n2364_n5888# 0.024979f
C241 drain_left.n218 a_n2364_n5888# 0.024979f
C242 drain_left.n219 a_n2364_n5888# 0.013423f
C243 drain_left.n220 a_n2364_n5888# 0.014212f
C244 drain_left.n221 a_n2364_n5888# 0.031726f
C245 drain_left.n222 a_n2364_n5888# 0.031726f
C246 drain_left.n223 a_n2364_n5888# 0.014212f
C247 drain_left.n224 a_n2364_n5888# 0.013423f
C248 drain_left.n225 a_n2364_n5888# 0.024979f
C249 drain_left.n226 a_n2364_n5888# 0.024979f
C250 drain_left.n227 a_n2364_n5888# 0.013423f
C251 drain_left.n228 a_n2364_n5888# 0.014212f
C252 drain_left.n229 a_n2364_n5888# 0.031726f
C253 drain_left.n230 a_n2364_n5888# 0.031726f
C254 drain_left.n231 a_n2364_n5888# 0.014212f
C255 drain_left.n232 a_n2364_n5888# 0.013423f
C256 drain_left.n233 a_n2364_n5888# 0.024979f
C257 drain_left.n234 a_n2364_n5888# 0.024979f
C258 drain_left.n235 a_n2364_n5888# 0.013423f
C259 drain_left.n236 a_n2364_n5888# 0.014212f
C260 drain_left.n237 a_n2364_n5888# 0.031726f
C261 drain_left.n238 a_n2364_n5888# 0.031726f
C262 drain_left.n239 a_n2364_n5888# 0.014212f
C263 drain_left.n240 a_n2364_n5888# 0.013423f
C264 drain_left.n241 a_n2364_n5888# 0.024979f
C265 drain_left.n242 a_n2364_n5888# 0.024979f
C266 drain_left.n243 a_n2364_n5888# 0.013423f
C267 drain_left.n244 a_n2364_n5888# 0.014212f
C268 drain_left.n245 a_n2364_n5888# 0.031726f
C269 drain_left.n246 a_n2364_n5888# 0.031726f
C270 drain_left.n247 a_n2364_n5888# 0.014212f
C271 drain_left.n248 a_n2364_n5888# 0.013423f
C272 drain_left.n249 a_n2364_n5888# 0.024979f
C273 drain_left.n250 a_n2364_n5888# 0.024979f
C274 drain_left.n251 a_n2364_n5888# 0.013423f
C275 drain_left.n252 a_n2364_n5888# 0.014212f
C276 drain_left.n253 a_n2364_n5888# 0.031726f
C277 drain_left.n254 a_n2364_n5888# 0.031726f
C278 drain_left.n255 a_n2364_n5888# 0.014212f
C279 drain_left.n256 a_n2364_n5888# 0.013423f
C280 drain_left.n257 a_n2364_n5888# 0.024979f
C281 drain_left.n258 a_n2364_n5888# 0.024979f
C282 drain_left.n259 a_n2364_n5888# 0.013423f
C283 drain_left.n260 a_n2364_n5888# 0.013818f
C284 drain_left.n261 a_n2364_n5888# 0.013818f
C285 drain_left.n262 a_n2364_n5888# 0.031726f
C286 drain_left.n263 a_n2364_n5888# 0.031726f
C287 drain_left.n264 a_n2364_n5888# 0.014212f
C288 drain_left.n265 a_n2364_n5888# 0.013423f
C289 drain_left.n266 a_n2364_n5888# 0.024979f
C290 drain_left.n267 a_n2364_n5888# 0.024979f
C291 drain_left.n268 a_n2364_n5888# 0.013423f
C292 drain_left.n269 a_n2364_n5888# 0.014212f
C293 drain_left.n270 a_n2364_n5888# 0.031726f
C294 drain_left.n271 a_n2364_n5888# 0.031726f
C295 drain_left.n272 a_n2364_n5888# 0.014212f
C296 drain_left.n273 a_n2364_n5888# 0.013423f
C297 drain_left.n274 a_n2364_n5888# 0.024979f
C298 drain_left.n275 a_n2364_n5888# 0.024979f
C299 drain_left.n276 a_n2364_n5888# 0.013423f
C300 drain_left.n277 a_n2364_n5888# 0.014212f
C301 drain_left.n278 a_n2364_n5888# 0.031726f
C302 drain_left.n279 a_n2364_n5888# 0.06749f
C303 drain_left.n280 a_n2364_n5888# 0.014212f
C304 drain_left.n281 a_n2364_n5888# 0.013423f
C305 drain_left.n282 a_n2364_n5888# 0.055008f
C306 drain_left.n283 a_n2364_n5888# 0.057f
C307 drain_left.t2 a_n2364_n5888# 0.493482f
C308 drain_left.t11 a_n2364_n5888# 0.493482f
C309 drain_left.n284 a_n2364_n5888# 4.54797f
C310 drain_left.n285 a_n2364_n5888# 0.469913f
C311 drain_left.t5 a_n2364_n5888# 0.493482f
C312 drain_left.t9 a_n2364_n5888# 0.493482f
C313 drain_left.n286 a_n2364_n5888# 4.54797f
C314 drain_left.n287 a_n2364_n5888# 0.354082f
C315 drain_left.t3 a_n2364_n5888# 0.493482f
C316 drain_left.t12 a_n2364_n5888# 0.493482f
C317 drain_left.n288 a_n2364_n5888# 4.54796f
C318 drain_left.n289 a_n2364_n5888# 0.575035f
C319 plus.n0 a_n2364_n5888# 0.040922f
C320 plus.t1 a_n2364_n5888# 2.02379f
C321 plus.t10 a_n2364_n5888# 2.02379f
C322 plus.n1 a_n2364_n5888# 0.040922f
C323 plus.t4 a_n2364_n5888# 2.02379f
C324 plus.n2 a_n2364_n5888# 0.738785f
C325 plus.n3 a_n2364_n5888# 0.040922f
C326 plus.t8 a_n2364_n5888# 2.02379f
C327 plus.t2 a_n2364_n5888# 2.02379f
C328 plus.n4 a_n2364_n5888# 0.738785f
C329 plus.t5 a_n2364_n5888# 2.04252f
C330 plus.n5 a_n2364_n5888# 0.723612f
C331 plus.t11 a_n2364_n5888# 2.02379f
C332 plus.n6 a_n2364_n5888# 0.743854f
C333 plus.n7 a_n2364_n5888# 0.009286f
C334 plus.n8 a_n2364_n5888# 0.172421f
C335 plus.n9 a_n2364_n5888# 0.040922f
C336 plus.n10 a_n2364_n5888# 0.040922f
C337 plus.n11 a_n2364_n5888# 0.009286f
C338 plus.n12 a_n2364_n5888# 0.738785f
C339 plus.n13 a_n2364_n5888# 0.009286f
C340 plus.n14 a_n2364_n5888# 0.040922f
C341 plus.n15 a_n2364_n5888# 0.040922f
C342 plus.n16 a_n2364_n5888# 0.040922f
C343 plus.n17 a_n2364_n5888# 0.009286f
C344 plus.n18 a_n2364_n5888# 0.738785f
C345 plus.n19 a_n2364_n5888# 0.009286f
C346 plus.n20 a_n2364_n5888# 0.737271f
C347 plus.n21 a_n2364_n5888# 0.744266f
C348 plus.n22 a_n2364_n5888# 0.040922f
C349 plus.t6 a_n2364_n5888# 2.02379f
C350 plus.n23 a_n2364_n5888# 0.040922f
C351 plus.t3 a_n2364_n5888# 2.02379f
C352 plus.t9 a_n2364_n5888# 2.02379f
C353 plus.n24 a_n2364_n5888# 0.738785f
C354 plus.n25 a_n2364_n5888# 0.040922f
C355 plus.t7 a_n2364_n5888# 2.02379f
C356 plus.t12 a_n2364_n5888# 2.02379f
C357 plus.n26 a_n2364_n5888# 0.738785f
C358 plus.t13 a_n2364_n5888# 2.04252f
C359 plus.n27 a_n2364_n5888# 0.723612f
C360 plus.t0 a_n2364_n5888# 2.02379f
C361 plus.n28 a_n2364_n5888# 0.743854f
C362 plus.n29 a_n2364_n5888# 0.009286f
C363 plus.n30 a_n2364_n5888# 0.172421f
C364 plus.n31 a_n2364_n5888# 0.040922f
C365 plus.n32 a_n2364_n5888# 0.040922f
C366 plus.n33 a_n2364_n5888# 0.009286f
C367 plus.n34 a_n2364_n5888# 0.738785f
C368 plus.n35 a_n2364_n5888# 0.009286f
C369 plus.n36 a_n2364_n5888# 0.040922f
C370 plus.n37 a_n2364_n5888# 0.040922f
C371 plus.n38 a_n2364_n5888# 0.040922f
C372 plus.n39 a_n2364_n5888# 0.009286f
C373 plus.n40 a_n2364_n5888# 0.738785f
C374 plus.n41 a_n2364_n5888# 0.009286f
C375 plus.n42 a_n2364_n5888# 0.737271f
C376 plus.n43 a_n2364_n5888# 1.70429f
C377 drain_right.n0 a_n2364_n5888# 0.034307f
C378 drain_right.n1 a_n2364_n5888# 0.024885f
C379 drain_right.n2 a_n2364_n5888# 0.013372f
C380 drain_right.n3 a_n2364_n5888# 0.031607f
C381 drain_right.n4 a_n2364_n5888# 0.014159f
C382 drain_right.n5 a_n2364_n5888# 0.024885f
C383 drain_right.n6 a_n2364_n5888# 0.013372f
C384 drain_right.n7 a_n2364_n5888# 0.031607f
C385 drain_right.n8 a_n2364_n5888# 0.014159f
C386 drain_right.n9 a_n2364_n5888# 0.024885f
C387 drain_right.n10 a_n2364_n5888# 0.013372f
C388 drain_right.n11 a_n2364_n5888# 0.031607f
C389 drain_right.n12 a_n2364_n5888# 0.014159f
C390 drain_right.n13 a_n2364_n5888# 0.024885f
C391 drain_right.n14 a_n2364_n5888# 0.013372f
C392 drain_right.n15 a_n2364_n5888# 0.031607f
C393 drain_right.n16 a_n2364_n5888# 0.014159f
C394 drain_right.n17 a_n2364_n5888# 0.024885f
C395 drain_right.n18 a_n2364_n5888# 0.013372f
C396 drain_right.n19 a_n2364_n5888# 0.031607f
C397 drain_right.n20 a_n2364_n5888# 0.014159f
C398 drain_right.n21 a_n2364_n5888# 0.024885f
C399 drain_right.n22 a_n2364_n5888# 0.013372f
C400 drain_right.n23 a_n2364_n5888# 0.031607f
C401 drain_right.n24 a_n2364_n5888# 0.014159f
C402 drain_right.n25 a_n2364_n5888# 0.024885f
C403 drain_right.n26 a_n2364_n5888# 0.013372f
C404 drain_right.n27 a_n2364_n5888# 0.031607f
C405 drain_right.n28 a_n2364_n5888# 0.014159f
C406 drain_right.n29 a_n2364_n5888# 0.024885f
C407 drain_right.n30 a_n2364_n5888# 0.013372f
C408 drain_right.n31 a_n2364_n5888# 0.031607f
C409 drain_right.n32 a_n2364_n5888# 0.014159f
C410 drain_right.n33 a_n2364_n5888# 0.024885f
C411 drain_right.n34 a_n2364_n5888# 0.013765f
C412 drain_right.n35 a_n2364_n5888# 0.031607f
C413 drain_right.n36 a_n2364_n5888# 0.014159f
C414 drain_right.n37 a_n2364_n5888# 0.024885f
C415 drain_right.n38 a_n2364_n5888# 0.013372f
C416 drain_right.n39 a_n2364_n5888# 0.031607f
C417 drain_right.n40 a_n2364_n5888# 0.014159f
C418 drain_right.n41 a_n2364_n5888# 0.024885f
C419 drain_right.n42 a_n2364_n5888# 0.013372f
C420 drain_right.n43 a_n2364_n5888# 0.023705f
C421 drain_right.n44 a_n2364_n5888# 0.022344f
C422 drain_right.t8 a_n2364_n5888# 0.055125f
C423 drain_right.n45 a_n2364_n5888# 0.303621f
C424 drain_right.n46 a_n2364_n5888# 2.69434f
C425 drain_right.n47 a_n2364_n5888# 0.013372f
C426 drain_right.n48 a_n2364_n5888# 0.014159f
C427 drain_right.n49 a_n2364_n5888# 0.031607f
C428 drain_right.n50 a_n2364_n5888# 0.031607f
C429 drain_right.n51 a_n2364_n5888# 0.014159f
C430 drain_right.n52 a_n2364_n5888# 0.013372f
C431 drain_right.n53 a_n2364_n5888# 0.024885f
C432 drain_right.n54 a_n2364_n5888# 0.024885f
C433 drain_right.n55 a_n2364_n5888# 0.013372f
C434 drain_right.n56 a_n2364_n5888# 0.014159f
C435 drain_right.n57 a_n2364_n5888# 0.031607f
C436 drain_right.n58 a_n2364_n5888# 0.031607f
C437 drain_right.n59 a_n2364_n5888# 0.014159f
C438 drain_right.n60 a_n2364_n5888# 0.013372f
C439 drain_right.n61 a_n2364_n5888# 0.024885f
C440 drain_right.n62 a_n2364_n5888# 0.024885f
C441 drain_right.n63 a_n2364_n5888# 0.013372f
C442 drain_right.n64 a_n2364_n5888# 0.013372f
C443 drain_right.n65 a_n2364_n5888# 0.014159f
C444 drain_right.n66 a_n2364_n5888# 0.031607f
C445 drain_right.n67 a_n2364_n5888# 0.031607f
C446 drain_right.n68 a_n2364_n5888# 0.031607f
C447 drain_right.n69 a_n2364_n5888# 0.013765f
C448 drain_right.n70 a_n2364_n5888# 0.013372f
C449 drain_right.n71 a_n2364_n5888# 0.024885f
C450 drain_right.n72 a_n2364_n5888# 0.024885f
C451 drain_right.n73 a_n2364_n5888# 0.013372f
C452 drain_right.n74 a_n2364_n5888# 0.014159f
C453 drain_right.n75 a_n2364_n5888# 0.031607f
C454 drain_right.n76 a_n2364_n5888# 0.031607f
C455 drain_right.n77 a_n2364_n5888# 0.014159f
C456 drain_right.n78 a_n2364_n5888# 0.013372f
C457 drain_right.n79 a_n2364_n5888# 0.024885f
C458 drain_right.n80 a_n2364_n5888# 0.024885f
C459 drain_right.n81 a_n2364_n5888# 0.013372f
C460 drain_right.n82 a_n2364_n5888# 0.014159f
C461 drain_right.n83 a_n2364_n5888# 0.031607f
C462 drain_right.n84 a_n2364_n5888# 0.031607f
C463 drain_right.n85 a_n2364_n5888# 0.014159f
C464 drain_right.n86 a_n2364_n5888# 0.013372f
C465 drain_right.n87 a_n2364_n5888# 0.024885f
C466 drain_right.n88 a_n2364_n5888# 0.024885f
C467 drain_right.n89 a_n2364_n5888# 0.013372f
C468 drain_right.n90 a_n2364_n5888# 0.014159f
C469 drain_right.n91 a_n2364_n5888# 0.031607f
C470 drain_right.n92 a_n2364_n5888# 0.031607f
C471 drain_right.n93 a_n2364_n5888# 0.014159f
C472 drain_right.n94 a_n2364_n5888# 0.013372f
C473 drain_right.n95 a_n2364_n5888# 0.024885f
C474 drain_right.n96 a_n2364_n5888# 0.024885f
C475 drain_right.n97 a_n2364_n5888# 0.013372f
C476 drain_right.n98 a_n2364_n5888# 0.014159f
C477 drain_right.n99 a_n2364_n5888# 0.031607f
C478 drain_right.n100 a_n2364_n5888# 0.031607f
C479 drain_right.n101 a_n2364_n5888# 0.014159f
C480 drain_right.n102 a_n2364_n5888# 0.013372f
C481 drain_right.n103 a_n2364_n5888# 0.024885f
C482 drain_right.n104 a_n2364_n5888# 0.024885f
C483 drain_right.n105 a_n2364_n5888# 0.013372f
C484 drain_right.n106 a_n2364_n5888# 0.014159f
C485 drain_right.n107 a_n2364_n5888# 0.031607f
C486 drain_right.n108 a_n2364_n5888# 0.031607f
C487 drain_right.n109 a_n2364_n5888# 0.031607f
C488 drain_right.n110 a_n2364_n5888# 0.014159f
C489 drain_right.n111 a_n2364_n5888# 0.013372f
C490 drain_right.n112 a_n2364_n5888# 0.024885f
C491 drain_right.n113 a_n2364_n5888# 0.024885f
C492 drain_right.n114 a_n2364_n5888# 0.013372f
C493 drain_right.n115 a_n2364_n5888# 0.013765f
C494 drain_right.n116 a_n2364_n5888# 0.013765f
C495 drain_right.n117 a_n2364_n5888# 0.031607f
C496 drain_right.n118 a_n2364_n5888# 0.031607f
C497 drain_right.n119 a_n2364_n5888# 0.014159f
C498 drain_right.n120 a_n2364_n5888# 0.013372f
C499 drain_right.n121 a_n2364_n5888# 0.024885f
C500 drain_right.n122 a_n2364_n5888# 0.024885f
C501 drain_right.n123 a_n2364_n5888# 0.013372f
C502 drain_right.n124 a_n2364_n5888# 0.014159f
C503 drain_right.n125 a_n2364_n5888# 0.031607f
C504 drain_right.n126 a_n2364_n5888# 0.031607f
C505 drain_right.n127 a_n2364_n5888# 0.014159f
C506 drain_right.n128 a_n2364_n5888# 0.013372f
C507 drain_right.n129 a_n2364_n5888# 0.024885f
C508 drain_right.n130 a_n2364_n5888# 0.024885f
C509 drain_right.n131 a_n2364_n5888# 0.013372f
C510 drain_right.n132 a_n2364_n5888# 0.014159f
C511 drain_right.n133 a_n2364_n5888# 0.031607f
C512 drain_right.n134 a_n2364_n5888# 0.067236f
C513 drain_right.n135 a_n2364_n5888# 0.014159f
C514 drain_right.n136 a_n2364_n5888# 0.013372f
C515 drain_right.n137 a_n2364_n5888# 0.054801f
C516 drain_right.n138 a_n2364_n5888# 0.056785f
C517 drain_right.t9 a_n2364_n5888# 0.491627f
C518 drain_right.t13 a_n2364_n5888# 0.491627f
C519 drain_right.n139 a_n2364_n5888# 4.53087f
C520 drain_right.n140 a_n2364_n5888# 0.446854f
C521 drain_right.t3 a_n2364_n5888# 0.491627f
C522 drain_right.t2 a_n2364_n5888# 0.491627f
C523 drain_right.n141 a_n2364_n5888# 4.53628f
C524 drain_right.t12 a_n2364_n5888# 0.491627f
C525 drain_right.t10 a_n2364_n5888# 0.491627f
C526 drain_right.n142 a_n2364_n5888# 4.53087f
C527 drain_right.n143 a_n2364_n5888# 0.655746f
C528 drain_right.n144 a_n2364_n5888# 2.13805f
C529 drain_right.t11 a_n2364_n5888# 0.491627f
C530 drain_right.t4 a_n2364_n5888# 0.491627f
C531 drain_right.n145 a_n2364_n5888# 4.53626f
C532 drain_right.t1 a_n2364_n5888# 0.491627f
C533 drain_right.t5 a_n2364_n5888# 0.491627f
C534 drain_right.n146 a_n2364_n5888# 4.53087f
C535 drain_right.n147 a_n2364_n5888# 0.71013f
C536 drain_right.t0 a_n2364_n5888# 0.491627f
C537 drain_right.t6 a_n2364_n5888# 0.491627f
C538 drain_right.n148 a_n2364_n5888# 4.53087f
C539 drain_right.n149 a_n2364_n5888# 0.35275f
C540 drain_right.n150 a_n2364_n5888# 0.034307f
C541 drain_right.n151 a_n2364_n5888# 0.024885f
C542 drain_right.n152 a_n2364_n5888# 0.013372f
C543 drain_right.n153 a_n2364_n5888# 0.031607f
C544 drain_right.n154 a_n2364_n5888# 0.014159f
C545 drain_right.n155 a_n2364_n5888# 0.024885f
C546 drain_right.n156 a_n2364_n5888# 0.013372f
C547 drain_right.n157 a_n2364_n5888# 0.031607f
C548 drain_right.n158 a_n2364_n5888# 0.014159f
C549 drain_right.n159 a_n2364_n5888# 0.024885f
C550 drain_right.n160 a_n2364_n5888# 0.013372f
C551 drain_right.n161 a_n2364_n5888# 0.031607f
C552 drain_right.n162 a_n2364_n5888# 0.014159f
C553 drain_right.n163 a_n2364_n5888# 0.024885f
C554 drain_right.n164 a_n2364_n5888# 0.013372f
C555 drain_right.n165 a_n2364_n5888# 0.031607f
C556 drain_right.n166 a_n2364_n5888# 0.031607f
C557 drain_right.n167 a_n2364_n5888# 0.014159f
C558 drain_right.n168 a_n2364_n5888# 0.024885f
C559 drain_right.n169 a_n2364_n5888# 0.013372f
C560 drain_right.n170 a_n2364_n5888# 0.031607f
C561 drain_right.n171 a_n2364_n5888# 0.014159f
C562 drain_right.n172 a_n2364_n5888# 0.024885f
C563 drain_right.n173 a_n2364_n5888# 0.013372f
C564 drain_right.n174 a_n2364_n5888# 0.031607f
C565 drain_right.n175 a_n2364_n5888# 0.014159f
C566 drain_right.n176 a_n2364_n5888# 0.024885f
C567 drain_right.n177 a_n2364_n5888# 0.013372f
C568 drain_right.n178 a_n2364_n5888# 0.031607f
C569 drain_right.n179 a_n2364_n5888# 0.014159f
C570 drain_right.n180 a_n2364_n5888# 0.024885f
C571 drain_right.n181 a_n2364_n5888# 0.013372f
C572 drain_right.n182 a_n2364_n5888# 0.031607f
C573 drain_right.n183 a_n2364_n5888# 0.014159f
C574 drain_right.n184 a_n2364_n5888# 0.024885f
C575 drain_right.n185 a_n2364_n5888# 0.013765f
C576 drain_right.n186 a_n2364_n5888# 0.031607f
C577 drain_right.n187 a_n2364_n5888# 0.013372f
C578 drain_right.n188 a_n2364_n5888# 0.014159f
C579 drain_right.n189 a_n2364_n5888# 0.024885f
C580 drain_right.n190 a_n2364_n5888# 0.013372f
C581 drain_right.n191 a_n2364_n5888# 0.031607f
C582 drain_right.n192 a_n2364_n5888# 0.014159f
C583 drain_right.n193 a_n2364_n5888# 0.024885f
C584 drain_right.n194 a_n2364_n5888# 0.013372f
C585 drain_right.n195 a_n2364_n5888# 0.023705f
C586 drain_right.n196 a_n2364_n5888# 0.022344f
C587 drain_right.t7 a_n2364_n5888# 0.055125f
C588 drain_right.n197 a_n2364_n5888# 0.303621f
C589 drain_right.n198 a_n2364_n5888# 2.69434f
C590 drain_right.n199 a_n2364_n5888# 0.013372f
C591 drain_right.n200 a_n2364_n5888# 0.014159f
C592 drain_right.n201 a_n2364_n5888# 0.031607f
C593 drain_right.n202 a_n2364_n5888# 0.031607f
C594 drain_right.n203 a_n2364_n5888# 0.014159f
C595 drain_right.n204 a_n2364_n5888# 0.013372f
C596 drain_right.n205 a_n2364_n5888# 0.024885f
C597 drain_right.n206 a_n2364_n5888# 0.024885f
C598 drain_right.n207 a_n2364_n5888# 0.013372f
C599 drain_right.n208 a_n2364_n5888# 0.014159f
C600 drain_right.n209 a_n2364_n5888# 0.031607f
C601 drain_right.n210 a_n2364_n5888# 0.031607f
C602 drain_right.n211 a_n2364_n5888# 0.014159f
C603 drain_right.n212 a_n2364_n5888# 0.013372f
C604 drain_right.n213 a_n2364_n5888# 0.024885f
C605 drain_right.n214 a_n2364_n5888# 0.024885f
C606 drain_right.n215 a_n2364_n5888# 0.013372f
C607 drain_right.n216 a_n2364_n5888# 0.014159f
C608 drain_right.n217 a_n2364_n5888# 0.031607f
C609 drain_right.n218 a_n2364_n5888# 0.031607f
C610 drain_right.n219 a_n2364_n5888# 0.031607f
C611 drain_right.n220 a_n2364_n5888# 0.013765f
C612 drain_right.n221 a_n2364_n5888# 0.013372f
C613 drain_right.n222 a_n2364_n5888# 0.024885f
C614 drain_right.n223 a_n2364_n5888# 0.024885f
C615 drain_right.n224 a_n2364_n5888# 0.013372f
C616 drain_right.n225 a_n2364_n5888# 0.014159f
C617 drain_right.n226 a_n2364_n5888# 0.031607f
C618 drain_right.n227 a_n2364_n5888# 0.031607f
C619 drain_right.n228 a_n2364_n5888# 0.014159f
C620 drain_right.n229 a_n2364_n5888# 0.013372f
C621 drain_right.n230 a_n2364_n5888# 0.024885f
C622 drain_right.n231 a_n2364_n5888# 0.024885f
C623 drain_right.n232 a_n2364_n5888# 0.013372f
C624 drain_right.n233 a_n2364_n5888# 0.014159f
C625 drain_right.n234 a_n2364_n5888# 0.031607f
C626 drain_right.n235 a_n2364_n5888# 0.031607f
C627 drain_right.n236 a_n2364_n5888# 0.014159f
C628 drain_right.n237 a_n2364_n5888# 0.013372f
C629 drain_right.n238 a_n2364_n5888# 0.024885f
C630 drain_right.n239 a_n2364_n5888# 0.024885f
C631 drain_right.n240 a_n2364_n5888# 0.013372f
C632 drain_right.n241 a_n2364_n5888# 0.014159f
C633 drain_right.n242 a_n2364_n5888# 0.031607f
C634 drain_right.n243 a_n2364_n5888# 0.031607f
C635 drain_right.n244 a_n2364_n5888# 0.014159f
C636 drain_right.n245 a_n2364_n5888# 0.013372f
C637 drain_right.n246 a_n2364_n5888# 0.024885f
C638 drain_right.n247 a_n2364_n5888# 0.024885f
C639 drain_right.n248 a_n2364_n5888# 0.013372f
C640 drain_right.n249 a_n2364_n5888# 0.014159f
C641 drain_right.n250 a_n2364_n5888# 0.031607f
C642 drain_right.n251 a_n2364_n5888# 0.031607f
C643 drain_right.n252 a_n2364_n5888# 0.014159f
C644 drain_right.n253 a_n2364_n5888# 0.013372f
C645 drain_right.n254 a_n2364_n5888# 0.024885f
C646 drain_right.n255 a_n2364_n5888# 0.024885f
C647 drain_right.n256 a_n2364_n5888# 0.013372f
C648 drain_right.n257 a_n2364_n5888# 0.014159f
C649 drain_right.n258 a_n2364_n5888# 0.031607f
C650 drain_right.n259 a_n2364_n5888# 0.031607f
C651 drain_right.n260 a_n2364_n5888# 0.014159f
C652 drain_right.n261 a_n2364_n5888# 0.013372f
C653 drain_right.n262 a_n2364_n5888# 0.024885f
C654 drain_right.n263 a_n2364_n5888# 0.024885f
C655 drain_right.n264 a_n2364_n5888# 0.013372f
C656 drain_right.n265 a_n2364_n5888# 0.013765f
C657 drain_right.n266 a_n2364_n5888# 0.013765f
C658 drain_right.n267 a_n2364_n5888# 0.031607f
C659 drain_right.n268 a_n2364_n5888# 0.031607f
C660 drain_right.n269 a_n2364_n5888# 0.014159f
C661 drain_right.n270 a_n2364_n5888# 0.013372f
C662 drain_right.n271 a_n2364_n5888# 0.024885f
C663 drain_right.n272 a_n2364_n5888# 0.024885f
C664 drain_right.n273 a_n2364_n5888# 0.013372f
C665 drain_right.n274 a_n2364_n5888# 0.014159f
C666 drain_right.n275 a_n2364_n5888# 0.031607f
C667 drain_right.n276 a_n2364_n5888# 0.031607f
C668 drain_right.n277 a_n2364_n5888# 0.014159f
C669 drain_right.n278 a_n2364_n5888# 0.013372f
C670 drain_right.n279 a_n2364_n5888# 0.024885f
C671 drain_right.n280 a_n2364_n5888# 0.024885f
C672 drain_right.n281 a_n2364_n5888# 0.013372f
C673 drain_right.n282 a_n2364_n5888# 0.014159f
C674 drain_right.n283 a_n2364_n5888# 0.031607f
C675 drain_right.n284 a_n2364_n5888# 0.067236f
C676 drain_right.n285 a_n2364_n5888# 0.014159f
C677 drain_right.n286 a_n2364_n5888# 0.013372f
C678 drain_right.n287 a_n2364_n5888# 0.054801f
C679 drain_right.n288 a_n2364_n5888# 0.054619f
C680 drain_right.n289 a_n2364_n5888# 0.346271f
C681 source.n0 a_n2364_n5888# 0.034996f
C682 source.n1 a_n2364_n5888# 0.025385f
C683 source.n2 a_n2364_n5888# 0.013641f
C684 source.n3 a_n2364_n5888# 0.032242f
C685 source.n4 a_n2364_n5888# 0.014443f
C686 source.n5 a_n2364_n5888# 0.025385f
C687 source.n6 a_n2364_n5888# 0.013641f
C688 source.n7 a_n2364_n5888# 0.032242f
C689 source.n8 a_n2364_n5888# 0.014443f
C690 source.n9 a_n2364_n5888# 0.025385f
C691 source.n10 a_n2364_n5888# 0.013641f
C692 source.n11 a_n2364_n5888# 0.032242f
C693 source.n12 a_n2364_n5888# 0.014443f
C694 source.n13 a_n2364_n5888# 0.025385f
C695 source.n14 a_n2364_n5888# 0.013641f
C696 source.n15 a_n2364_n5888# 0.032242f
C697 source.n16 a_n2364_n5888# 0.032242f
C698 source.n17 a_n2364_n5888# 0.014443f
C699 source.n18 a_n2364_n5888# 0.025385f
C700 source.n19 a_n2364_n5888# 0.013641f
C701 source.n20 a_n2364_n5888# 0.032242f
C702 source.n21 a_n2364_n5888# 0.014443f
C703 source.n22 a_n2364_n5888# 0.025385f
C704 source.n23 a_n2364_n5888# 0.013641f
C705 source.n24 a_n2364_n5888# 0.032242f
C706 source.n25 a_n2364_n5888# 0.014443f
C707 source.n26 a_n2364_n5888# 0.025385f
C708 source.n27 a_n2364_n5888# 0.013641f
C709 source.n28 a_n2364_n5888# 0.032242f
C710 source.n29 a_n2364_n5888# 0.014443f
C711 source.n30 a_n2364_n5888# 0.025385f
C712 source.n31 a_n2364_n5888# 0.013641f
C713 source.n32 a_n2364_n5888# 0.032242f
C714 source.n33 a_n2364_n5888# 0.014443f
C715 source.n34 a_n2364_n5888# 0.025385f
C716 source.n35 a_n2364_n5888# 0.014042f
C717 source.n36 a_n2364_n5888# 0.032242f
C718 source.n37 a_n2364_n5888# 0.013641f
C719 source.n38 a_n2364_n5888# 0.014443f
C720 source.n39 a_n2364_n5888# 0.025385f
C721 source.n40 a_n2364_n5888# 0.013641f
C722 source.n41 a_n2364_n5888# 0.032242f
C723 source.n42 a_n2364_n5888# 0.014443f
C724 source.n43 a_n2364_n5888# 0.025385f
C725 source.n44 a_n2364_n5888# 0.013641f
C726 source.n45 a_n2364_n5888# 0.024182f
C727 source.n46 a_n2364_n5888# 0.022793f
C728 source.t0 a_n2364_n5888# 0.056232f
C729 source.n47 a_n2364_n5888# 0.30972f
C730 source.n48 a_n2364_n5888# 2.74846f
C731 source.n49 a_n2364_n5888# 0.013641f
C732 source.n50 a_n2364_n5888# 0.014443f
C733 source.n51 a_n2364_n5888# 0.032242f
C734 source.n52 a_n2364_n5888# 0.032242f
C735 source.n53 a_n2364_n5888# 0.014443f
C736 source.n54 a_n2364_n5888# 0.013641f
C737 source.n55 a_n2364_n5888# 0.025385f
C738 source.n56 a_n2364_n5888# 0.025385f
C739 source.n57 a_n2364_n5888# 0.013641f
C740 source.n58 a_n2364_n5888# 0.014443f
C741 source.n59 a_n2364_n5888# 0.032242f
C742 source.n60 a_n2364_n5888# 0.032242f
C743 source.n61 a_n2364_n5888# 0.014443f
C744 source.n62 a_n2364_n5888# 0.013641f
C745 source.n63 a_n2364_n5888# 0.025385f
C746 source.n64 a_n2364_n5888# 0.025385f
C747 source.n65 a_n2364_n5888# 0.013641f
C748 source.n66 a_n2364_n5888# 0.014443f
C749 source.n67 a_n2364_n5888# 0.032242f
C750 source.n68 a_n2364_n5888# 0.032242f
C751 source.n69 a_n2364_n5888# 0.032242f
C752 source.n70 a_n2364_n5888# 0.014042f
C753 source.n71 a_n2364_n5888# 0.013641f
C754 source.n72 a_n2364_n5888# 0.025385f
C755 source.n73 a_n2364_n5888# 0.025385f
C756 source.n74 a_n2364_n5888# 0.013641f
C757 source.n75 a_n2364_n5888# 0.014443f
C758 source.n76 a_n2364_n5888# 0.032242f
C759 source.n77 a_n2364_n5888# 0.032242f
C760 source.n78 a_n2364_n5888# 0.014443f
C761 source.n79 a_n2364_n5888# 0.013641f
C762 source.n80 a_n2364_n5888# 0.025385f
C763 source.n81 a_n2364_n5888# 0.025385f
C764 source.n82 a_n2364_n5888# 0.013641f
C765 source.n83 a_n2364_n5888# 0.014443f
C766 source.n84 a_n2364_n5888# 0.032242f
C767 source.n85 a_n2364_n5888# 0.032242f
C768 source.n86 a_n2364_n5888# 0.014443f
C769 source.n87 a_n2364_n5888# 0.013641f
C770 source.n88 a_n2364_n5888# 0.025385f
C771 source.n89 a_n2364_n5888# 0.025385f
C772 source.n90 a_n2364_n5888# 0.013641f
C773 source.n91 a_n2364_n5888# 0.014443f
C774 source.n92 a_n2364_n5888# 0.032242f
C775 source.n93 a_n2364_n5888# 0.032242f
C776 source.n94 a_n2364_n5888# 0.014443f
C777 source.n95 a_n2364_n5888# 0.013641f
C778 source.n96 a_n2364_n5888# 0.025385f
C779 source.n97 a_n2364_n5888# 0.025385f
C780 source.n98 a_n2364_n5888# 0.013641f
C781 source.n99 a_n2364_n5888# 0.014443f
C782 source.n100 a_n2364_n5888# 0.032242f
C783 source.n101 a_n2364_n5888# 0.032242f
C784 source.n102 a_n2364_n5888# 0.014443f
C785 source.n103 a_n2364_n5888# 0.013641f
C786 source.n104 a_n2364_n5888# 0.025385f
C787 source.n105 a_n2364_n5888# 0.025385f
C788 source.n106 a_n2364_n5888# 0.013641f
C789 source.n107 a_n2364_n5888# 0.014443f
C790 source.n108 a_n2364_n5888# 0.032242f
C791 source.n109 a_n2364_n5888# 0.032242f
C792 source.n110 a_n2364_n5888# 0.014443f
C793 source.n111 a_n2364_n5888# 0.013641f
C794 source.n112 a_n2364_n5888# 0.025385f
C795 source.n113 a_n2364_n5888# 0.025385f
C796 source.n114 a_n2364_n5888# 0.013641f
C797 source.n115 a_n2364_n5888# 0.014042f
C798 source.n116 a_n2364_n5888# 0.014042f
C799 source.n117 a_n2364_n5888# 0.032242f
C800 source.n118 a_n2364_n5888# 0.032242f
C801 source.n119 a_n2364_n5888# 0.014443f
C802 source.n120 a_n2364_n5888# 0.013641f
C803 source.n121 a_n2364_n5888# 0.025385f
C804 source.n122 a_n2364_n5888# 0.025385f
C805 source.n123 a_n2364_n5888# 0.013641f
C806 source.n124 a_n2364_n5888# 0.014443f
C807 source.n125 a_n2364_n5888# 0.032242f
C808 source.n126 a_n2364_n5888# 0.032242f
C809 source.n127 a_n2364_n5888# 0.014443f
C810 source.n128 a_n2364_n5888# 0.013641f
C811 source.n129 a_n2364_n5888# 0.025385f
C812 source.n130 a_n2364_n5888# 0.025385f
C813 source.n131 a_n2364_n5888# 0.013641f
C814 source.n132 a_n2364_n5888# 0.014443f
C815 source.n133 a_n2364_n5888# 0.032242f
C816 source.n134 a_n2364_n5888# 0.068587f
C817 source.n135 a_n2364_n5888# 0.014443f
C818 source.n136 a_n2364_n5888# 0.013641f
C819 source.n137 a_n2364_n5888# 0.055902f
C820 source.n138 a_n2364_n5888# 0.038165f
C821 source.n139 a_n2364_n5888# 2.03875f
C822 source.t6 a_n2364_n5888# 0.501503f
C823 source.t3 a_n2364_n5888# 0.501503f
C824 source.n140 a_n2364_n5888# 4.53867f
C825 source.n141 a_n2364_n5888# 0.408554f
C826 source.t1 a_n2364_n5888# 0.501503f
C827 source.t4 a_n2364_n5888# 0.501503f
C828 source.n142 a_n2364_n5888# 4.53867f
C829 source.n143 a_n2364_n5888# 0.408554f
C830 source.t9 a_n2364_n5888# 0.501503f
C831 source.t8 a_n2364_n5888# 0.501503f
C832 source.n144 a_n2364_n5888# 4.53867f
C833 source.n145 a_n2364_n5888# 0.410669f
C834 source.n146 a_n2364_n5888# 0.034996f
C835 source.n147 a_n2364_n5888# 0.025385f
C836 source.n148 a_n2364_n5888# 0.013641f
C837 source.n149 a_n2364_n5888# 0.032242f
C838 source.n150 a_n2364_n5888# 0.014443f
C839 source.n151 a_n2364_n5888# 0.025385f
C840 source.n152 a_n2364_n5888# 0.013641f
C841 source.n153 a_n2364_n5888# 0.032242f
C842 source.n154 a_n2364_n5888# 0.014443f
C843 source.n155 a_n2364_n5888# 0.025385f
C844 source.n156 a_n2364_n5888# 0.013641f
C845 source.n157 a_n2364_n5888# 0.032242f
C846 source.n158 a_n2364_n5888# 0.014443f
C847 source.n159 a_n2364_n5888# 0.025385f
C848 source.n160 a_n2364_n5888# 0.013641f
C849 source.n161 a_n2364_n5888# 0.032242f
C850 source.n162 a_n2364_n5888# 0.032242f
C851 source.n163 a_n2364_n5888# 0.014443f
C852 source.n164 a_n2364_n5888# 0.025385f
C853 source.n165 a_n2364_n5888# 0.013641f
C854 source.n166 a_n2364_n5888# 0.032242f
C855 source.n167 a_n2364_n5888# 0.014443f
C856 source.n168 a_n2364_n5888# 0.025385f
C857 source.n169 a_n2364_n5888# 0.013641f
C858 source.n170 a_n2364_n5888# 0.032242f
C859 source.n171 a_n2364_n5888# 0.014443f
C860 source.n172 a_n2364_n5888# 0.025385f
C861 source.n173 a_n2364_n5888# 0.013641f
C862 source.n174 a_n2364_n5888# 0.032242f
C863 source.n175 a_n2364_n5888# 0.014443f
C864 source.n176 a_n2364_n5888# 0.025385f
C865 source.n177 a_n2364_n5888# 0.013641f
C866 source.n178 a_n2364_n5888# 0.032242f
C867 source.n179 a_n2364_n5888# 0.014443f
C868 source.n180 a_n2364_n5888# 0.025385f
C869 source.n181 a_n2364_n5888# 0.014042f
C870 source.n182 a_n2364_n5888# 0.032242f
C871 source.n183 a_n2364_n5888# 0.013641f
C872 source.n184 a_n2364_n5888# 0.014443f
C873 source.n185 a_n2364_n5888# 0.025385f
C874 source.n186 a_n2364_n5888# 0.013641f
C875 source.n187 a_n2364_n5888# 0.032242f
C876 source.n188 a_n2364_n5888# 0.014443f
C877 source.n189 a_n2364_n5888# 0.025385f
C878 source.n190 a_n2364_n5888# 0.013641f
C879 source.n191 a_n2364_n5888# 0.024182f
C880 source.n192 a_n2364_n5888# 0.022793f
C881 source.t14 a_n2364_n5888# 0.056232f
C882 source.n193 a_n2364_n5888# 0.30972f
C883 source.n194 a_n2364_n5888# 2.74846f
C884 source.n195 a_n2364_n5888# 0.013641f
C885 source.n196 a_n2364_n5888# 0.014443f
C886 source.n197 a_n2364_n5888# 0.032242f
C887 source.n198 a_n2364_n5888# 0.032242f
C888 source.n199 a_n2364_n5888# 0.014443f
C889 source.n200 a_n2364_n5888# 0.013641f
C890 source.n201 a_n2364_n5888# 0.025385f
C891 source.n202 a_n2364_n5888# 0.025385f
C892 source.n203 a_n2364_n5888# 0.013641f
C893 source.n204 a_n2364_n5888# 0.014443f
C894 source.n205 a_n2364_n5888# 0.032242f
C895 source.n206 a_n2364_n5888# 0.032242f
C896 source.n207 a_n2364_n5888# 0.014443f
C897 source.n208 a_n2364_n5888# 0.013641f
C898 source.n209 a_n2364_n5888# 0.025385f
C899 source.n210 a_n2364_n5888# 0.025385f
C900 source.n211 a_n2364_n5888# 0.013641f
C901 source.n212 a_n2364_n5888# 0.014443f
C902 source.n213 a_n2364_n5888# 0.032242f
C903 source.n214 a_n2364_n5888# 0.032242f
C904 source.n215 a_n2364_n5888# 0.032242f
C905 source.n216 a_n2364_n5888# 0.014042f
C906 source.n217 a_n2364_n5888# 0.013641f
C907 source.n218 a_n2364_n5888# 0.025385f
C908 source.n219 a_n2364_n5888# 0.025385f
C909 source.n220 a_n2364_n5888# 0.013641f
C910 source.n221 a_n2364_n5888# 0.014443f
C911 source.n222 a_n2364_n5888# 0.032242f
C912 source.n223 a_n2364_n5888# 0.032242f
C913 source.n224 a_n2364_n5888# 0.014443f
C914 source.n225 a_n2364_n5888# 0.013641f
C915 source.n226 a_n2364_n5888# 0.025385f
C916 source.n227 a_n2364_n5888# 0.025385f
C917 source.n228 a_n2364_n5888# 0.013641f
C918 source.n229 a_n2364_n5888# 0.014443f
C919 source.n230 a_n2364_n5888# 0.032242f
C920 source.n231 a_n2364_n5888# 0.032242f
C921 source.n232 a_n2364_n5888# 0.014443f
C922 source.n233 a_n2364_n5888# 0.013641f
C923 source.n234 a_n2364_n5888# 0.025385f
C924 source.n235 a_n2364_n5888# 0.025385f
C925 source.n236 a_n2364_n5888# 0.013641f
C926 source.n237 a_n2364_n5888# 0.014443f
C927 source.n238 a_n2364_n5888# 0.032242f
C928 source.n239 a_n2364_n5888# 0.032242f
C929 source.n240 a_n2364_n5888# 0.014443f
C930 source.n241 a_n2364_n5888# 0.013641f
C931 source.n242 a_n2364_n5888# 0.025385f
C932 source.n243 a_n2364_n5888# 0.025385f
C933 source.n244 a_n2364_n5888# 0.013641f
C934 source.n245 a_n2364_n5888# 0.014443f
C935 source.n246 a_n2364_n5888# 0.032242f
C936 source.n247 a_n2364_n5888# 0.032242f
C937 source.n248 a_n2364_n5888# 0.014443f
C938 source.n249 a_n2364_n5888# 0.013641f
C939 source.n250 a_n2364_n5888# 0.025385f
C940 source.n251 a_n2364_n5888# 0.025385f
C941 source.n252 a_n2364_n5888# 0.013641f
C942 source.n253 a_n2364_n5888# 0.014443f
C943 source.n254 a_n2364_n5888# 0.032242f
C944 source.n255 a_n2364_n5888# 0.032242f
C945 source.n256 a_n2364_n5888# 0.014443f
C946 source.n257 a_n2364_n5888# 0.013641f
C947 source.n258 a_n2364_n5888# 0.025385f
C948 source.n259 a_n2364_n5888# 0.025385f
C949 source.n260 a_n2364_n5888# 0.013641f
C950 source.n261 a_n2364_n5888# 0.014042f
C951 source.n262 a_n2364_n5888# 0.014042f
C952 source.n263 a_n2364_n5888# 0.032242f
C953 source.n264 a_n2364_n5888# 0.032242f
C954 source.n265 a_n2364_n5888# 0.014443f
C955 source.n266 a_n2364_n5888# 0.013641f
C956 source.n267 a_n2364_n5888# 0.025385f
C957 source.n268 a_n2364_n5888# 0.025385f
C958 source.n269 a_n2364_n5888# 0.013641f
C959 source.n270 a_n2364_n5888# 0.014443f
C960 source.n271 a_n2364_n5888# 0.032242f
C961 source.n272 a_n2364_n5888# 0.032242f
C962 source.n273 a_n2364_n5888# 0.014443f
C963 source.n274 a_n2364_n5888# 0.013641f
C964 source.n275 a_n2364_n5888# 0.025385f
C965 source.n276 a_n2364_n5888# 0.025385f
C966 source.n277 a_n2364_n5888# 0.013641f
C967 source.n278 a_n2364_n5888# 0.014443f
C968 source.n279 a_n2364_n5888# 0.032242f
C969 source.n280 a_n2364_n5888# 0.068587f
C970 source.n281 a_n2364_n5888# 0.014443f
C971 source.n282 a_n2364_n5888# 0.013641f
C972 source.n283 a_n2364_n5888# 0.055902f
C973 source.n284 a_n2364_n5888# 0.038165f
C974 source.n285 a_n2364_n5888# 0.167492f
C975 source.t13 a_n2364_n5888# 0.501503f
C976 source.t18 a_n2364_n5888# 0.501503f
C977 source.n286 a_n2364_n5888# 4.53867f
C978 source.n287 a_n2364_n5888# 0.408554f
C979 source.t16 a_n2364_n5888# 0.501503f
C980 source.t21 a_n2364_n5888# 0.501503f
C981 source.n288 a_n2364_n5888# 4.53867f
C982 source.n289 a_n2364_n5888# 0.408554f
C983 source.t17 a_n2364_n5888# 0.501503f
C984 source.t19 a_n2364_n5888# 0.501503f
C985 source.n290 a_n2364_n5888# 4.53867f
C986 source.n291 a_n2364_n5888# 2.83691f
C987 source.t27 a_n2364_n5888# 0.501503f
C988 source.t2 a_n2364_n5888# 0.501503f
C989 source.n292 a_n2364_n5888# 4.53867f
C990 source.n293 a_n2364_n5888# 2.83691f
C991 source.t11 a_n2364_n5888# 0.501503f
C992 source.t5 a_n2364_n5888# 0.501503f
C993 source.n294 a_n2364_n5888# 4.53867f
C994 source.n295 a_n2364_n5888# 0.408555f
C995 source.t10 a_n2364_n5888# 0.501503f
C996 source.t7 a_n2364_n5888# 0.501503f
C997 source.n296 a_n2364_n5888# 4.53867f
C998 source.n297 a_n2364_n5888# 0.408555f
C999 source.n298 a_n2364_n5888# 0.034996f
C1000 source.n299 a_n2364_n5888# 0.025385f
C1001 source.n300 a_n2364_n5888# 0.013641f
C1002 source.n301 a_n2364_n5888# 0.032242f
C1003 source.n302 a_n2364_n5888# 0.014443f
C1004 source.n303 a_n2364_n5888# 0.025385f
C1005 source.n304 a_n2364_n5888# 0.013641f
C1006 source.n305 a_n2364_n5888# 0.032242f
C1007 source.n306 a_n2364_n5888# 0.014443f
C1008 source.n307 a_n2364_n5888# 0.025385f
C1009 source.n308 a_n2364_n5888# 0.013641f
C1010 source.n309 a_n2364_n5888# 0.032242f
C1011 source.n310 a_n2364_n5888# 0.014443f
C1012 source.n311 a_n2364_n5888# 0.025385f
C1013 source.n312 a_n2364_n5888# 0.013641f
C1014 source.n313 a_n2364_n5888# 0.032242f
C1015 source.n314 a_n2364_n5888# 0.014443f
C1016 source.n315 a_n2364_n5888# 0.025385f
C1017 source.n316 a_n2364_n5888# 0.013641f
C1018 source.n317 a_n2364_n5888# 0.032242f
C1019 source.n318 a_n2364_n5888# 0.014443f
C1020 source.n319 a_n2364_n5888# 0.025385f
C1021 source.n320 a_n2364_n5888# 0.013641f
C1022 source.n321 a_n2364_n5888# 0.032242f
C1023 source.n322 a_n2364_n5888# 0.014443f
C1024 source.n323 a_n2364_n5888# 0.025385f
C1025 source.n324 a_n2364_n5888# 0.013641f
C1026 source.n325 a_n2364_n5888# 0.032242f
C1027 source.n326 a_n2364_n5888# 0.014443f
C1028 source.n327 a_n2364_n5888# 0.025385f
C1029 source.n328 a_n2364_n5888# 0.013641f
C1030 source.n329 a_n2364_n5888# 0.032242f
C1031 source.n330 a_n2364_n5888# 0.014443f
C1032 source.n331 a_n2364_n5888# 0.025385f
C1033 source.n332 a_n2364_n5888# 0.014042f
C1034 source.n333 a_n2364_n5888# 0.032242f
C1035 source.n334 a_n2364_n5888# 0.014443f
C1036 source.n335 a_n2364_n5888# 0.025385f
C1037 source.n336 a_n2364_n5888# 0.013641f
C1038 source.n337 a_n2364_n5888# 0.032242f
C1039 source.n338 a_n2364_n5888# 0.014443f
C1040 source.n339 a_n2364_n5888# 0.025385f
C1041 source.n340 a_n2364_n5888# 0.013641f
C1042 source.n341 a_n2364_n5888# 0.024182f
C1043 source.n342 a_n2364_n5888# 0.022793f
C1044 source.t26 a_n2364_n5888# 0.056232f
C1045 source.n343 a_n2364_n5888# 0.30972f
C1046 source.n344 a_n2364_n5888# 2.74846f
C1047 source.n345 a_n2364_n5888# 0.013641f
C1048 source.n346 a_n2364_n5888# 0.014443f
C1049 source.n347 a_n2364_n5888# 0.032242f
C1050 source.n348 a_n2364_n5888# 0.032242f
C1051 source.n349 a_n2364_n5888# 0.014443f
C1052 source.n350 a_n2364_n5888# 0.013641f
C1053 source.n351 a_n2364_n5888# 0.025385f
C1054 source.n352 a_n2364_n5888# 0.025385f
C1055 source.n353 a_n2364_n5888# 0.013641f
C1056 source.n354 a_n2364_n5888# 0.014443f
C1057 source.n355 a_n2364_n5888# 0.032242f
C1058 source.n356 a_n2364_n5888# 0.032242f
C1059 source.n357 a_n2364_n5888# 0.014443f
C1060 source.n358 a_n2364_n5888# 0.013641f
C1061 source.n359 a_n2364_n5888# 0.025385f
C1062 source.n360 a_n2364_n5888# 0.025385f
C1063 source.n361 a_n2364_n5888# 0.013641f
C1064 source.n362 a_n2364_n5888# 0.013641f
C1065 source.n363 a_n2364_n5888# 0.014443f
C1066 source.n364 a_n2364_n5888# 0.032242f
C1067 source.n365 a_n2364_n5888# 0.032242f
C1068 source.n366 a_n2364_n5888# 0.032242f
C1069 source.n367 a_n2364_n5888# 0.014042f
C1070 source.n368 a_n2364_n5888# 0.013641f
C1071 source.n369 a_n2364_n5888# 0.025385f
C1072 source.n370 a_n2364_n5888# 0.025385f
C1073 source.n371 a_n2364_n5888# 0.013641f
C1074 source.n372 a_n2364_n5888# 0.014443f
C1075 source.n373 a_n2364_n5888# 0.032242f
C1076 source.n374 a_n2364_n5888# 0.032242f
C1077 source.n375 a_n2364_n5888# 0.014443f
C1078 source.n376 a_n2364_n5888# 0.013641f
C1079 source.n377 a_n2364_n5888# 0.025385f
C1080 source.n378 a_n2364_n5888# 0.025385f
C1081 source.n379 a_n2364_n5888# 0.013641f
C1082 source.n380 a_n2364_n5888# 0.014443f
C1083 source.n381 a_n2364_n5888# 0.032242f
C1084 source.n382 a_n2364_n5888# 0.032242f
C1085 source.n383 a_n2364_n5888# 0.014443f
C1086 source.n384 a_n2364_n5888# 0.013641f
C1087 source.n385 a_n2364_n5888# 0.025385f
C1088 source.n386 a_n2364_n5888# 0.025385f
C1089 source.n387 a_n2364_n5888# 0.013641f
C1090 source.n388 a_n2364_n5888# 0.014443f
C1091 source.n389 a_n2364_n5888# 0.032242f
C1092 source.n390 a_n2364_n5888# 0.032242f
C1093 source.n391 a_n2364_n5888# 0.014443f
C1094 source.n392 a_n2364_n5888# 0.013641f
C1095 source.n393 a_n2364_n5888# 0.025385f
C1096 source.n394 a_n2364_n5888# 0.025385f
C1097 source.n395 a_n2364_n5888# 0.013641f
C1098 source.n396 a_n2364_n5888# 0.014443f
C1099 source.n397 a_n2364_n5888# 0.032242f
C1100 source.n398 a_n2364_n5888# 0.032242f
C1101 source.n399 a_n2364_n5888# 0.014443f
C1102 source.n400 a_n2364_n5888# 0.013641f
C1103 source.n401 a_n2364_n5888# 0.025385f
C1104 source.n402 a_n2364_n5888# 0.025385f
C1105 source.n403 a_n2364_n5888# 0.013641f
C1106 source.n404 a_n2364_n5888# 0.014443f
C1107 source.n405 a_n2364_n5888# 0.032242f
C1108 source.n406 a_n2364_n5888# 0.032242f
C1109 source.n407 a_n2364_n5888# 0.032242f
C1110 source.n408 a_n2364_n5888# 0.014443f
C1111 source.n409 a_n2364_n5888# 0.013641f
C1112 source.n410 a_n2364_n5888# 0.025385f
C1113 source.n411 a_n2364_n5888# 0.025385f
C1114 source.n412 a_n2364_n5888# 0.013641f
C1115 source.n413 a_n2364_n5888# 0.014042f
C1116 source.n414 a_n2364_n5888# 0.014042f
C1117 source.n415 a_n2364_n5888# 0.032242f
C1118 source.n416 a_n2364_n5888# 0.032242f
C1119 source.n417 a_n2364_n5888# 0.014443f
C1120 source.n418 a_n2364_n5888# 0.013641f
C1121 source.n419 a_n2364_n5888# 0.025385f
C1122 source.n420 a_n2364_n5888# 0.025385f
C1123 source.n421 a_n2364_n5888# 0.013641f
C1124 source.n422 a_n2364_n5888# 0.014443f
C1125 source.n423 a_n2364_n5888# 0.032242f
C1126 source.n424 a_n2364_n5888# 0.032242f
C1127 source.n425 a_n2364_n5888# 0.014443f
C1128 source.n426 a_n2364_n5888# 0.013641f
C1129 source.n427 a_n2364_n5888# 0.025385f
C1130 source.n428 a_n2364_n5888# 0.025385f
C1131 source.n429 a_n2364_n5888# 0.013641f
C1132 source.n430 a_n2364_n5888# 0.014443f
C1133 source.n431 a_n2364_n5888# 0.032242f
C1134 source.n432 a_n2364_n5888# 0.068587f
C1135 source.n433 a_n2364_n5888# 0.014443f
C1136 source.n434 a_n2364_n5888# 0.013641f
C1137 source.n435 a_n2364_n5888# 0.055902f
C1138 source.n436 a_n2364_n5888# 0.038165f
C1139 source.n437 a_n2364_n5888# 0.167492f
C1140 source.t24 a_n2364_n5888# 0.501503f
C1141 source.t15 a_n2364_n5888# 0.501503f
C1142 source.n438 a_n2364_n5888# 4.53867f
C1143 source.n439 a_n2364_n5888# 0.410671f
C1144 source.t22 a_n2364_n5888# 0.501503f
C1145 source.t20 a_n2364_n5888# 0.501503f
C1146 source.n440 a_n2364_n5888# 4.53867f
C1147 source.n441 a_n2364_n5888# 0.408555f
C1148 source.t25 a_n2364_n5888# 0.501503f
C1149 source.t12 a_n2364_n5888# 0.501503f
C1150 source.n442 a_n2364_n5888# 4.53867f
C1151 source.n443 a_n2364_n5888# 0.408555f
C1152 source.n444 a_n2364_n5888# 0.034996f
C1153 source.n445 a_n2364_n5888# 0.025385f
C1154 source.n446 a_n2364_n5888# 0.013641f
C1155 source.n447 a_n2364_n5888# 0.032242f
C1156 source.n448 a_n2364_n5888# 0.014443f
C1157 source.n449 a_n2364_n5888# 0.025385f
C1158 source.n450 a_n2364_n5888# 0.013641f
C1159 source.n451 a_n2364_n5888# 0.032242f
C1160 source.n452 a_n2364_n5888# 0.014443f
C1161 source.n453 a_n2364_n5888# 0.025385f
C1162 source.n454 a_n2364_n5888# 0.013641f
C1163 source.n455 a_n2364_n5888# 0.032242f
C1164 source.n456 a_n2364_n5888# 0.014443f
C1165 source.n457 a_n2364_n5888# 0.025385f
C1166 source.n458 a_n2364_n5888# 0.013641f
C1167 source.n459 a_n2364_n5888# 0.032242f
C1168 source.n460 a_n2364_n5888# 0.014443f
C1169 source.n461 a_n2364_n5888# 0.025385f
C1170 source.n462 a_n2364_n5888# 0.013641f
C1171 source.n463 a_n2364_n5888# 0.032242f
C1172 source.n464 a_n2364_n5888# 0.014443f
C1173 source.n465 a_n2364_n5888# 0.025385f
C1174 source.n466 a_n2364_n5888# 0.013641f
C1175 source.n467 a_n2364_n5888# 0.032242f
C1176 source.n468 a_n2364_n5888# 0.014443f
C1177 source.n469 a_n2364_n5888# 0.025385f
C1178 source.n470 a_n2364_n5888# 0.013641f
C1179 source.n471 a_n2364_n5888# 0.032242f
C1180 source.n472 a_n2364_n5888# 0.014443f
C1181 source.n473 a_n2364_n5888# 0.025385f
C1182 source.n474 a_n2364_n5888# 0.013641f
C1183 source.n475 a_n2364_n5888# 0.032242f
C1184 source.n476 a_n2364_n5888# 0.014443f
C1185 source.n477 a_n2364_n5888# 0.025385f
C1186 source.n478 a_n2364_n5888# 0.014042f
C1187 source.n479 a_n2364_n5888# 0.032242f
C1188 source.n480 a_n2364_n5888# 0.014443f
C1189 source.n481 a_n2364_n5888# 0.025385f
C1190 source.n482 a_n2364_n5888# 0.013641f
C1191 source.n483 a_n2364_n5888# 0.032242f
C1192 source.n484 a_n2364_n5888# 0.014443f
C1193 source.n485 a_n2364_n5888# 0.025385f
C1194 source.n486 a_n2364_n5888# 0.013641f
C1195 source.n487 a_n2364_n5888# 0.024182f
C1196 source.n488 a_n2364_n5888# 0.022793f
C1197 source.t23 a_n2364_n5888# 0.056232f
C1198 source.n489 a_n2364_n5888# 0.30972f
C1199 source.n490 a_n2364_n5888# 2.74846f
C1200 source.n491 a_n2364_n5888# 0.013641f
C1201 source.n492 a_n2364_n5888# 0.014443f
C1202 source.n493 a_n2364_n5888# 0.032242f
C1203 source.n494 a_n2364_n5888# 0.032242f
C1204 source.n495 a_n2364_n5888# 0.014443f
C1205 source.n496 a_n2364_n5888# 0.013641f
C1206 source.n497 a_n2364_n5888# 0.025385f
C1207 source.n498 a_n2364_n5888# 0.025385f
C1208 source.n499 a_n2364_n5888# 0.013641f
C1209 source.n500 a_n2364_n5888# 0.014443f
C1210 source.n501 a_n2364_n5888# 0.032242f
C1211 source.n502 a_n2364_n5888# 0.032242f
C1212 source.n503 a_n2364_n5888# 0.014443f
C1213 source.n504 a_n2364_n5888# 0.013641f
C1214 source.n505 a_n2364_n5888# 0.025385f
C1215 source.n506 a_n2364_n5888# 0.025385f
C1216 source.n507 a_n2364_n5888# 0.013641f
C1217 source.n508 a_n2364_n5888# 0.013641f
C1218 source.n509 a_n2364_n5888# 0.014443f
C1219 source.n510 a_n2364_n5888# 0.032242f
C1220 source.n511 a_n2364_n5888# 0.032242f
C1221 source.n512 a_n2364_n5888# 0.032242f
C1222 source.n513 a_n2364_n5888# 0.014042f
C1223 source.n514 a_n2364_n5888# 0.013641f
C1224 source.n515 a_n2364_n5888# 0.025385f
C1225 source.n516 a_n2364_n5888# 0.025385f
C1226 source.n517 a_n2364_n5888# 0.013641f
C1227 source.n518 a_n2364_n5888# 0.014443f
C1228 source.n519 a_n2364_n5888# 0.032242f
C1229 source.n520 a_n2364_n5888# 0.032242f
C1230 source.n521 a_n2364_n5888# 0.014443f
C1231 source.n522 a_n2364_n5888# 0.013641f
C1232 source.n523 a_n2364_n5888# 0.025385f
C1233 source.n524 a_n2364_n5888# 0.025385f
C1234 source.n525 a_n2364_n5888# 0.013641f
C1235 source.n526 a_n2364_n5888# 0.014443f
C1236 source.n527 a_n2364_n5888# 0.032242f
C1237 source.n528 a_n2364_n5888# 0.032242f
C1238 source.n529 a_n2364_n5888# 0.014443f
C1239 source.n530 a_n2364_n5888# 0.013641f
C1240 source.n531 a_n2364_n5888# 0.025385f
C1241 source.n532 a_n2364_n5888# 0.025385f
C1242 source.n533 a_n2364_n5888# 0.013641f
C1243 source.n534 a_n2364_n5888# 0.014443f
C1244 source.n535 a_n2364_n5888# 0.032242f
C1245 source.n536 a_n2364_n5888# 0.032242f
C1246 source.n537 a_n2364_n5888# 0.014443f
C1247 source.n538 a_n2364_n5888# 0.013641f
C1248 source.n539 a_n2364_n5888# 0.025385f
C1249 source.n540 a_n2364_n5888# 0.025385f
C1250 source.n541 a_n2364_n5888# 0.013641f
C1251 source.n542 a_n2364_n5888# 0.014443f
C1252 source.n543 a_n2364_n5888# 0.032242f
C1253 source.n544 a_n2364_n5888# 0.032242f
C1254 source.n545 a_n2364_n5888# 0.014443f
C1255 source.n546 a_n2364_n5888# 0.013641f
C1256 source.n547 a_n2364_n5888# 0.025385f
C1257 source.n548 a_n2364_n5888# 0.025385f
C1258 source.n549 a_n2364_n5888# 0.013641f
C1259 source.n550 a_n2364_n5888# 0.014443f
C1260 source.n551 a_n2364_n5888# 0.032242f
C1261 source.n552 a_n2364_n5888# 0.032242f
C1262 source.n553 a_n2364_n5888# 0.032242f
C1263 source.n554 a_n2364_n5888# 0.014443f
C1264 source.n555 a_n2364_n5888# 0.013641f
C1265 source.n556 a_n2364_n5888# 0.025385f
C1266 source.n557 a_n2364_n5888# 0.025385f
C1267 source.n558 a_n2364_n5888# 0.013641f
C1268 source.n559 a_n2364_n5888# 0.014042f
C1269 source.n560 a_n2364_n5888# 0.014042f
C1270 source.n561 a_n2364_n5888# 0.032242f
C1271 source.n562 a_n2364_n5888# 0.032242f
C1272 source.n563 a_n2364_n5888# 0.014443f
C1273 source.n564 a_n2364_n5888# 0.013641f
C1274 source.n565 a_n2364_n5888# 0.025385f
C1275 source.n566 a_n2364_n5888# 0.025385f
C1276 source.n567 a_n2364_n5888# 0.013641f
C1277 source.n568 a_n2364_n5888# 0.014443f
C1278 source.n569 a_n2364_n5888# 0.032242f
C1279 source.n570 a_n2364_n5888# 0.032242f
C1280 source.n571 a_n2364_n5888# 0.014443f
C1281 source.n572 a_n2364_n5888# 0.013641f
C1282 source.n573 a_n2364_n5888# 0.025385f
C1283 source.n574 a_n2364_n5888# 0.025385f
C1284 source.n575 a_n2364_n5888# 0.013641f
C1285 source.n576 a_n2364_n5888# 0.014443f
C1286 source.n577 a_n2364_n5888# 0.032242f
C1287 source.n578 a_n2364_n5888# 0.068587f
C1288 source.n579 a_n2364_n5888# 0.014443f
C1289 source.n580 a_n2364_n5888# 0.013641f
C1290 source.n581 a_n2364_n5888# 0.055902f
C1291 source.n582 a_n2364_n5888# 0.038165f
C1292 source.n583 a_n2364_n5888# 0.296765f
C1293 source.n584 a_n2364_n5888# 2.72475f
C1294 minus.n0 a_n2364_n5888# 0.040664f
C1295 minus.n1 a_n2364_n5888# 0.009227f
C1296 minus.t13 a_n2364_n5888# 2.01104f
C1297 minus.n2 a_n2364_n5888# 0.040664f
C1298 minus.n3 a_n2364_n5888# 0.009227f
C1299 minus.t12 a_n2364_n5888# 2.01104f
C1300 minus.n4 a_n2364_n5888# 0.171335f
C1301 minus.t9 a_n2364_n5888# 2.02965f
C1302 minus.n5 a_n2364_n5888# 0.719053f
C1303 minus.t2 a_n2364_n5888# 2.01104f
C1304 minus.n6 a_n2364_n5888# 0.739168f
C1305 minus.n7 a_n2364_n5888# 0.009227f
C1306 minus.t8 a_n2364_n5888# 2.01104f
C1307 minus.n8 a_n2364_n5888# 0.734131f
C1308 minus.n9 a_n2364_n5888# 0.040664f
C1309 minus.n10 a_n2364_n5888# 0.040664f
C1310 minus.n11 a_n2364_n5888# 0.040664f
C1311 minus.n12 a_n2364_n5888# 0.734131f
C1312 minus.n13 a_n2364_n5888# 0.009227f
C1313 minus.t7 a_n2364_n5888# 2.01104f
C1314 minus.n14 a_n2364_n5888# 0.734131f
C1315 minus.n15 a_n2364_n5888# 0.040664f
C1316 minus.n16 a_n2364_n5888# 0.040664f
C1317 minus.n17 a_n2364_n5888# 0.040664f
C1318 minus.n18 a_n2364_n5888# 0.734131f
C1319 minus.n19 a_n2364_n5888# 0.009227f
C1320 minus.t6 a_n2364_n5888# 2.01104f
C1321 minus.n20 a_n2364_n5888# 0.732626f
C1322 minus.n21 a_n2364_n5888# 2.19027f
C1323 minus.n22 a_n2364_n5888# 0.040664f
C1324 minus.n23 a_n2364_n5888# 0.009227f
C1325 minus.n24 a_n2364_n5888# 0.040664f
C1326 minus.n25 a_n2364_n5888# 0.009227f
C1327 minus.n26 a_n2364_n5888# 0.171335f
C1328 minus.t5 a_n2364_n5888# 2.02965f
C1329 minus.n27 a_n2364_n5888# 0.719053f
C1330 minus.t4 a_n2364_n5888# 2.01104f
C1331 minus.n28 a_n2364_n5888# 0.739168f
C1332 minus.n29 a_n2364_n5888# 0.009227f
C1333 minus.t0 a_n2364_n5888# 2.01104f
C1334 minus.n30 a_n2364_n5888# 0.734131f
C1335 minus.n31 a_n2364_n5888# 0.040664f
C1336 minus.n32 a_n2364_n5888# 0.040664f
C1337 minus.n33 a_n2364_n5888# 0.040664f
C1338 minus.t1 a_n2364_n5888# 2.01104f
C1339 minus.n34 a_n2364_n5888# 0.734131f
C1340 minus.n35 a_n2364_n5888# 0.009227f
C1341 minus.t3 a_n2364_n5888# 2.01104f
C1342 minus.n36 a_n2364_n5888# 0.734131f
C1343 minus.n37 a_n2364_n5888# 0.040664f
C1344 minus.n38 a_n2364_n5888# 0.040664f
C1345 minus.n39 a_n2364_n5888# 0.040664f
C1346 minus.t10 a_n2364_n5888# 2.01104f
C1347 minus.n40 a_n2364_n5888# 0.734131f
C1348 minus.n41 a_n2364_n5888# 0.009227f
C1349 minus.t11 a_n2364_n5888# 2.01104f
C1350 minus.n42 a_n2364_n5888# 0.732626f
C1351 minus.n43 a_n2364_n5888# 0.280132f
C1352 minus.n44 a_n2364_n5888# 2.5708f
.ends

