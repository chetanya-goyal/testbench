* NGSPICE file created from diffpair317.ext - technology: sky130A

.subckt diffpair317 minus drain_right drain_left source plus
X0 a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X1 source.t23 plus.t0 drain_left.t8 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X3 drain_right.t15 minus.t0 source.t25 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X4 drain_left.t7 plus.t1 source.t22 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X5 a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X6 drain_left.t2 plus.t2 source.t21 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X7 drain_left.t1 plus.t3 source.t20 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X8 a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X9 source.t1 minus.t1 drain_right.t14 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X10 source.t4 minus.t2 drain_right.t13 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X11 drain_right.t12 minus.t3 source.t6 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X12 drain_left.t0 plus.t4 source.t19 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X13 source.t30 minus.t4 drain_right.t11 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X14 source.t29 minus.t5 drain_right.t10 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X15 drain_right.t9 minus.t6 source.t24 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X16 source.t31 minus.t7 drain_right.t8 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X17 source.t18 plus.t5 drain_left.t5 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X18 drain_right.t7 minus.t8 source.t27 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X19 source.t28 minus.t9 drain_right.t6 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X20 drain_right.t5 minus.t10 source.t7 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X21 drain_left.t14 plus.t6 source.t17 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X22 source.t2 minus.t11 drain_right.t4 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X23 drain_right.t3 minus.t12 source.t0 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X24 source.t16 plus.t7 drain_left.t12 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X25 source.t15 plus.t8 drain_left.t11 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X26 drain_left.t4 plus.t9 source.t14 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X27 drain_left.t15 plus.t10 source.t13 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X28 source.t26 minus.t13 drain_right.t2 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X29 source.t12 plus.t11 drain_left.t10 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X30 drain_right.t1 minus.t14 source.t5 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X31 source.t11 plus.t12 drain_left.t9 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X32 drain_left.t3 plus.t13 source.t10 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X33 source.t9 plus.t14 drain_left.t6 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X34 drain_right.t0 minus.t15 source.t3 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X35 source.t8 plus.t15 drain_left.t13 a_n2750_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
R0 plus.n7 plus.t14 250.877
R1 plus.n29 plus.t4 250.877
R2 plus.n20 plus.t6 229.855
R3 plus.n18 plus.t7 229.855
R4 plus.n17 plus.t9 229.855
R5 plus.n3 plus.t12 229.855
R6 plus.n11 plus.t10 229.855
R7 plus.n5 plus.t11 229.855
R8 plus.n6 plus.t13 229.855
R9 plus.n42 plus.t8 229.855
R10 plus.n40 plus.t1 229.855
R11 plus.n39 plus.t5 229.855
R12 plus.n25 plus.t3 229.855
R13 plus.n33 plus.t15 229.855
R14 plus.n27 plus.t2 229.855
R15 plus.n28 plus.t0 229.855
R16 plus.n10 plus.n9 161.3
R17 plus.n11 plus.n4 161.3
R18 plus.n13 plus.n12 161.3
R19 plus.n14 plus.n3 161.3
R20 plus.n16 plus.n15 161.3
R21 plus.n19 plus.n0 161.3
R22 plus.n21 plus.n20 161.3
R23 plus.n32 plus.n31 161.3
R24 plus.n33 plus.n26 161.3
R25 plus.n35 plus.n34 161.3
R26 plus.n36 plus.n25 161.3
R27 plus.n38 plus.n37 161.3
R28 plus.n41 plus.n22 161.3
R29 plus.n43 plus.n42 161.3
R30 plus.n8 plus.n5 80.6037
R31 plus.n17 plus.n2 80.6037
R32 plus.n18 plus.n1 80.6037
R33 plus.n30 plus.n27 80.6037
R34 plus.n39 plus.n24 80.6037
R35 plus.n40 plus.n23 80.6037
R36 plus.n18 plus.n17 48.2005
R37 plus.n6 plus.n5 48.2005
R38 plus.n40 plus.n39 48.2005
R39 plus.n28 plus.n27 48.2005
R40 plus.n17 plus.n16 43.0884
R41 plus.n10 plus.n5 43.0884
R42 plus.n39 plus.n38 43.0884
R43 plus.n32 plus.n27 43.0884
R44 plus.n19 plus.n18 40.1672
R45 plus.n41 plus.n40 40.1672
R46 plus.n8 plus.n7 31.6481
R47 plus.n30 plus.n29 31.6481
R48 plus plus.n43 31.3021
R49 plus.n12 plus.n11 24.1005
R50 plus.n12 plus.n3 24.1005
R51 plus.n34 plus.n25 24.1005
R52 plus.n34 plus.n33 24.1005
R53 plus.n7 plus.n6 17.444
R54 plus.n29 plus.n28 17.444
R55 plus plus.n21 10.027
R56 plus.n20 plus.n19 8.03383
R57 plus.n42 plus.n41 8.03383
R58 plus.n16 plus.n3 5.11262
R59 plus.n11 plus.n10 5.11262
R60 plus.n38 plus.n25 5.11262
R61 plus.n33 plus.n32 5.11262
R62 plus.n2 plus.n1 0.380177
R63 plus.n24 plus.n23 0.380177
R64 plus.n9 plus.n8 0.285035
R65 plus.n15 plus.n2 0.285035
R66 plus.n1 plus.n0 0.285035
R67 plus.n23 plus.n22 0.285035
R68 plus.n37 plus.n24 0.285035
R69 plus.n31 plus.n30 0.285035
R70 plus.n9 plus.n4 0.189894
R71 plus.n13 plus.n4 0.189894
R72 plus.n14 plus.n13 0.189894
R73 plus.n15 plus.n14 0.189894
R74 plus.n21 plus.n0 0.189894
R75 plus.n43 plus.n22 0.189894
R76 plus.n37 plus.n36 0.189894
R77 plus.n36 plus.n35 0.189894
R78 plus.n35 plus.n26 0.189894
R79 plus.n31 plus.n26 0.189894
R80 drain_left.n9 drain_left.n7 68.165
R81 drain_left.n5 drain_left.n3 68.1648
R82 drain_left.n2 drain_left.n0 68.1648
R83 drain_left.n11 drain_left.n10 67.1908
R84 drain_left.n9 drain_left.n8 67.1908
R85 drain_left.n13 drain_left.n12 67.1907
R86 drain_left.n5 drain_left.n4 67.1907
R87 drain_left.n2 drain_left.n1 67.1907
R88 drain_left drain_left.n6 29.1535
R89 drain_left drain_left.n13 6.62735
R90 drain_left.n3 drain_left.t8 3.3005
R91 drain_left.n3 drain_left.t0 3.3005
R92 drain_left.n4 drain_left.t13 3.3005
R93 drain_left.n4 drain_left.t2 3.3005
R94 drain_left.n1 drain_left.t5 3.3005
R95 drain_left.n1 drain_left.t1 3.3005
R96 drain_left.n0 drain_left.t11 3.3005
R97 drain_left.n0 drain_left.t7 3.3005
R98 drain_left.n12 drain_left.t12 3.3005
R99 drain_left.n12 drain_left.t14 3.3005
R100 drain_left.n10 drain_left.t9 3.3005
R101 drain_left.n10 drain_left.t4 3.3005
R102 drain_left.n8 drain_left.t10 3.3005
R103 drain_left.n8 drain_left.t15 3.3005
R104 drain_left.n7 drain_left.t6 3.3005
R105 drain_left.n7 drain_left.t3 3.3005
R106 drain_left.n11 drain_left.n9 0.974638
R107 drain_left.n13 drain_left.n11 0.974638
R108 drain_left.n6 drain_left.n5 0.432223
R109 drain_left.n6 drain_left.n2 0.432223
R110 source.n274 source.n248 289.615
R111 source.n236 source.n210 289.615
R112 source.n204 source.n178 289.615
R113 source.n166 source.n140 289.615
R114 source.n26 source.n0 289.615
R115 source.n64 source.n38 289.615
R116 source.n96 source.n70 289.615
R117 source.n134 source.n108 289.615
R118 source.n259 source.n258 185
R119 source.n256 source.n255 185
R120 source.n265 source.n264 185
R121 source.n267 source.n266 185
R122 source.n252 source.n251 185
R123 source.n273 source.n272 185
R124 source.n275 source.n274 185
R125 source.n221 source.n220 185
R126 source.n218 source.n217 185
R127 source.n227 source.n226 185
R128 source.n229 source.n228 185
R129 source.n214 source.n213 185
R130 source.n235 source.n234 185
R131 source.n237 source.n236 185
R132 source.n189 source.n188 185
R133 source.n186 source.n185 185
R134 source.n195 source.n194 185
R135 source.n197 source.n196 185
R136 source.n182 source.n181 185
R137 source.n203 source.n202 185
R138 source.n205 source.n204 185
R139 source.n151 source.n150 185
R140 source.n148 source.n147 185
R141 source.n157 source.n156 185
R142 source.n159 source.n158 185
R143 source.n144 source.n143 185
R144 source.n165 source.n164 185
R145 source.n167 source.n166 185
R146 source.n27 source.n26 185
R147 source.n25 source.n24 185
R148 source.n4 source.n3 185
R149 source.n19 source.n18 185
R150 source.n17 source.n16 185
R151 source.n8 source.n7 185
R152 source.n11 source.n10 185
R153 source.n65 source.n64 185
R154 source.n63 source.n62 185
R155 source.n42 source.n41 185
R156 source.n57 source.n56 185
R157 source.n55 source.n54 185
R158 source.n46 source.n45 185
R159 source.n49 source.n48 185
R160 source.n97 source.n96 185
R161 source.n95 source.n94 185
R162 source.n74 source.n73 185
R163 source.n89 source.n88 185
R164 source.n87 source.n86 185
R165 source.n78 source.n77 185
R166 source.n81 source.n80 185
R167 source.n135 source.n134 185
R168 source.n133 source.n132 185
R169 source.n112 source.n111 185
R170 source.n127 source.n126 185
R171 source.n125 source.n124 185
R172 source.n116 source.n115 185
R173 source.n119 source.n118 185
R174 source.t7 source.n257 147.661
R175 source.t31 source.n219 147.661
R176 source.t19 source.n187 147.661
R177 source.t15 source.n149 147.661
R178 source.t17 source.n9 147.661
R179 source.t9 source.n47 147.661
R180 source.t27 source.n79 147.661
R181 source.t26 source.n117 147.661
R182 source.n258 source.n255 104.615
R183 source.n265 source.n255 104.615
R184 source.n266 source.n265 104.615
R185 source.n266 source.n251 104.615
R186 source.n273 source.n251 104.615
R187 source.n274 source.n273 104.615
R188 source.n220 source.n217 104.615
R189 source.n227 source.n217 104.615
R190 source.n228 source.n227 104.615
R191 source.n228 source.n213 104.615
R192 source.n235 source.n213 104.615
R193 source.n236 source.n235 104.615
R194 source.n188 source.n185 104.615
R195 source.n195 source.n185 104.615
R196 source.n196 source.n195 104.615
R197 source.n196 source.n181 104.615
R198 source.n203 source.n181 104.615
R199 source.n204 source.n203 104.615
R200 source.n150 source.n147 104.615
R201 source.n157 source.n147 104.615
R202 source.n158 source.n157 104.615
R203 source.n158 source.n143 104.615
R204 source.n165 source.n143 104.615
R205 source.n166 source.n165 104.615
R206 source.n26 source.n25 104.615
R207 source.n25 source.n3 104.615
R208 source.n18 source.n3 104.615
R209 source.n18 source.n17 104.615
R210 source.n17 source.n7 104.615
R211 source.n10 source.n7 104.615
R212 source.n64 source.n63 104.615
R213 source.n63 source.n41 104.615
R214 source.n56 source.n41 104.615
R215 source.n56 source.n55 104.615
R216 source.n55 source.n45 104.615
R217 source.n48 source.n45 104.615
R218 source.n96 source.n95 104.615
R219 source.n95 source.n73 104.615
R220 source.n88 source.n73 104.615
R221 source.n88 source.n87 104.615
R222 source.n87 source.n77 104.615
R223 source.n80 source.n77 104.615
R224 source.n134 source.n133 104.615
R225 source.n133 source.n111 104.615
R226 source.n126 source.n111 104.615
R227 source.n126 source.n125 104.615
R228 source.n125 source.n115 104.615
R229 source.n118 source.n115 104.615
R230 source.n258 source.t7 52.3082
R231 source.n220 source.t31 52.3082
R232 source.n188 source.t19 52.3082
R233 source.n150 source.t15 52.3082
R234 source.n10 source.t17 52.3082
R235 source.n48 source.t9 52.3082
R236 source.n80 source.t27 52.3082
R237 source.n118 source.t26 52.3082
R238 source.n33 source.n32 50.512
R239 source.n35 source.n34 50.512
R240 source.n37 source.n36 50.512
R241 source.n103 source.n102 50.512
R242 source.n105 source.n104 50.512
R243 source.n107 source.n106 50.512
R244 source.n247 source.n246 50.5119
R245 source.n245 source.n244 50.5119
R246 source.n243 source.n242 50.5119
R247 source.n177 source.n176 50.5119
R248 source.n175 source.n174 50.5119
R249 source.n173 source.n172 50.5119
R250 source.n279 source.n278 32.1853
R251 source.n241 source.n240 32.1853
R252 source.n209 source.n208 32.1853
R253 source.n171 source.n170 32.1853
R254 source.n31 source.n30 32.1853
R255 source.n69 source.n68 32.1853
R256 source.n101 source.n100 32.1853
R257 source.n139 source.n138 32.1853
R258 source.n171 source.n139 17.7164
R259 source.n259 source.n257 15.6674
R260 source.n221 source.n219 15.6674
R261 source.n189 source.n187 15.6674
R262 source.n151 source.n149 15.6674
R263 source.n11 source.n9 15.6674
R264 source.n49 source.n47 15.6674
R265 source.n81 source.n79 15.6674
R266 source.n119 source.n117 15.6674
R267 source.n260 source.n256 12.8005
R268 source.n222 source.n218 12.8005
R269 source.n190 source.n186 12.8005
R270 source.n152 source.n148 12.8005
R271 source.n12 source.n8 12.8005
R272 source.n50 source.n46 12.8005
R273 source.n82 source.n78 12.8005
R274 source.n120 source.n116 12.8005
R275 source.n264 source.n263 12.0247
R276 source.n226 source.n225 12.0247
R277 source.n194 source.n193 12.0247
R278 source.n156 source.n155 12.0247
R279 source.n16 source.n15 12.0247
R280 source.n54 source.n53 12.0247
R281 source.n86 source.n85 12.0247
R282 source.n124 source.n123 12.0247
R283 source.n280 source.n31 11.9664
R284 source.n267 source.n254 11.249
R285 source.n229 source.n216 11.249
R286 source.n197 source.n184 11.249
R287 source.n159 source.n146 11.249
R288 source.n19 source.n6 11.249
R289 source.n57 source.n44 11.249
R290 source.n89 source.n76 11.249
R291 source.n127 source.n114 11.249
R292 source.n268 source.n252 10.4732
R293 source.n230 source.n214 10.4732
R294 source.n198 source.n182 10.4732
R295 source.n160 source.n144 10.4732
R296 source.n20 source.n4 10.4732
R297 source.n58 source.n42 10.4732
R298 source.n90 source.n74 10.4732
R299 source.n128 source.n112 10.4732
R300 source.n272 source.n271 9.69747
R301 source.n234 source.n233 9.69747
R302 source.n202 source.n201 9.69747
R303 source.n164 source.n163 9.69747
R304 source.n24 source.n23 9.69747
R305 source.n62 source.n61 9.69747
R306 source.n94 source.n93 9.69747
R307 source.n132 source.n131 9.69747
R308 source.n278 source.n277 9.45567
R309 source.n240 source.n239 9.45567
R310 source.n208 source.n207 9.45567
R311 source.n170 source.n169 9.45567
R312 source.n30 source.n29 9.45567
R313 source.n68 source.n67 9.45567
R314 source.n100 source.n99 9.45567
R315 source.n138 source.n137 9.45567
R316 source.n277 source.n276 9.3005
R317 source.n250 source.n249 9.3005
R318 source.n271 source.n270 9.3005
R319 source.n269 source.n268 9.3005
R320 source.n254 source.n253 9.3005
R321 source.n263 source.n262 9.3005
R322 source.n261 source.n260 9.3005
R323 source.n239 source.n238 9.3005
R324 source.n212 source.n211 9.3005
R325 source.n233 source.n232 9.3005
R326 source.n231 source.n230 9.3005
R327 source.n216 source.n215 9.3005
R328 source.n225 source.n224 9.3005
R329 source.n223 source.n222 9.3005
R330 source.n207 source.n206 9.3005
R331 source.n180 source.n179 9.3005
R332 source.n201 source.n200 9.3005
R333 source.n199 source.n198 9.3005
R334 source.n184 source.n183 9.3005
R335 source.n193 source.n192 9.3005
R336 source.n191 source.n190 9.3005
R337 source.n169 source.n168 9.3005
R338 source.n142 source.n141 9.3005
R339 source.n163 source.n162 9.3005
R340 source.n161 source.n160 9.3005
R341 source.n146 source.n145 9.3005
R342 source.n155 source.n154 9.3005
R343 source.n153 source.n152 9.3005
R344 source.n29 source.n28 9.3005
R345 source.n2 source.n1 9.3005
R346 source.n23 source.n22 9.3005
R347 source.n21 source.n20 9.3005
R348 source.n6 source.n5 9.3005
R349 source.n15 source.n14 9.3005
R350 source.n13 source.n12 9.3005
R351 source.n67 source.n66 9.3005
R352 source.n40 source.n39 9.3005
R353 source.n61 source.n60 9.3005
R354 source.n59 source.n58 9.3005
R355 source.n44 source.n43 9.3005
R356 source.n53 source.n52 9.3005
R357 source.n51 source.n50 9.3005
R358 source.n99 source.n98 9.3005
R359 source.n72 source.n71 9.3005
R360 source.n93 source.n92 9.3005
R361 source.n91 source.n90 9.3005
R362 source.n76 source.n75 9.3005
R363 source.n85 source.n84 9.3005
R364 source.n83 source.n82 9.3005
R365 source.n137 source.n136 9.3005
R366 source.n110 source.n109 9.3005
R367 source.n131 source.n130 9.3005
R368 source.n129 source.n128 9.3005
R369 source.n114 source.n113 9.3005
R370 source.n123 source.n122 9.3005
R371 source.n121 source.n120 9.3005
R372 source.n275 source.n250 8.92171
R373 source.n237 source.n212 8.92171
R374 source.n205 source.n180 8.92171
R375 source.n167 source.n142 8.92171
R376 source.n27 source.n2 8.92171
R377 source.n65 source.n40 8.92171
R378 source.n97 source.n72 8.92171
R379 source.n135 source.n110 8.92171
R380 source.n276 source.n248 8.14595
R381 source.n238 source.n210 8.14595
R382 source.n206 source.n178 8.14595
R383 source.n168 source.n140 8.14595
R384 source.n28 source.n0 8.14595
R385 source.n66 source.n38 8.14595
R386 source.n98 source.n70 8.14595
R387 source.n136 source.n108 8.14595
R388 source.n278 source.n248 5.81868
R389 source.n240 source.n210 5.81868
R390 source.n208 source.n178 5.81868
R391 source.n170 source.n140 5.81868
R392 source.n30 source.n0 5.81868
R393 source.n68 source.n38 5.81868
R394 source.n100 source.n70 5.81868
R395 source.n138 source.n108 5.81868
R396 source.n280 source.n279 5.7505
R397 source.n276 source.n275 5.04292
R398 source.n238 source.n237 5.04292
R399 source.n206 source.n205 5.04292
R400 source.n168 source.n167 5.04292
R401 source.n28 source.n27 5.04292
R402 source.n66 source.n65 5.04292
R403 source.n98 source.n97 5.04292
R404 source.n136 source.n135 5.04292
R405 source.n261 source.n257 4.38594
R406 source.n223 source.n219 4.38594
R407 source.n191 source.n187 4.38594
R408 source.n153 source.n149 4.38594
R409 source.n13 source.n9 4.38594
R410 source.n51 source.n47 4.38594
R411 source.n83 source.n79 4.38594
R412 source.n121 source.n117 4.38594
R413 source.n272 source.n250 4.26717
R414 source.n234 source.n212 4.26717
R415 source.n202 source.n180 4.26717
R416 source.n164 source.n142 4.26717
R417 source.n24 source.n2 4.26717
R418 source.n62 source.n40 4.26717
R419 source.n94 source.n72 4.26717
R420 source.n132 source.n110 4.26717
R421 source.n271 source.n252 3.49141
R422 source.n233 source.n214 3.49141
R423 source.n201 source.n182 3.49141
R424 source.n163 source.n144 3.49141
R425 source.n23 source.n4 3.49141
R426 source.n61 source.n42 3.49141
R427 source.n93 source.n74 3.49141
R428 source.n131 source.n112 3.49141
R429 source.n246 source.t5 3.3005
R430 source.n246 source.t1 3.3005
R431 source.n244 source.t3 3.3005
R432 source.n244 source.t30 3.3005
R433 source.n242 source.t25 3.3005
R434 source.n242 source.t4 3.3005
R435 source.n176 source.t21 3.3005
R436 source.n176 source.t23 3.3005
R437 source.n174 source.t20 3.3005
R438 source.n174 source.t8 3.3005
R439 source.n172 source.t22 3.3005
R440 source.n172 source.t18 3.3005
R441 source.n32 source.t14 3.3005
R442 source.n32 source.t16 3.3005
R443 source.n34 source.t13 3.3005
R444 source.n34 source.t11 3.3005
R445 source.n36 source.t10 3.3005
R446 source.n36 source.t12 3.3005
R447 source.n102 source.t6 3.3005
R448 source.n102 source.t29 3.3005
R449 source.n104 source.t0 3.3005
R450 source.n104 source.t2 3.3005
R451 source.n106 source.t24 3.3005
R452 source.n106 source.t28 3.3005
R453 source.n268 source.n267 2.71565
R454 source.n230 source.n229 2.71565
R455 source.n198 source.n197 2.71565
R456 source.n160 source.n159 2.71565
R457 source.n20 source.n19 2.71565
R458 source.n58 source.n57 2.71565
R459 source.n90 source.n89 2.71565
R460 source.n128 source.n127 2.71565
R461 source.n264 source.n254 1.93989
R462 source.n226 source.n216 1.93989
R463 source.n194 source.n184 1.93989
R464 source.n156 source.n146 1.93989
R465 source.n16 source.n6 1.93989
R466 source.n54 source.n44 1.93989
R467 source.n86 source.n76 1.93989
R468 source.n124 source.n114 1.93989
R469 source.n263 source.n256 1.16414
R470 source.n225 source.n218 1.16414
R471 source.n193 source.n186 1.16414
R472 source.n155 source.n148 1.16414
R473 source.n15 source.n8 1.16414
R474 source.n53 source.n46 1.16414
R475 source.n85 source.n78 1.16414
R476 source.n123 source.n116 1.16414
R477 source.n139 source.n107 0.974638
R478 source.n107 source.n105 0.974638
R479 source.n105 source.n103 0.974638
R480 source.n103 source.n101 0.974638
R481 source.n69 source.n37 0.974638
R482 source.n37 source.n35 0.974638
R483 source.n35 source.n33 0.974638
R484 source.n33 source.n31 0.974638
R485 source.n173 source.n171 0.974638
R486 source.n175 source.n173 0.974638
R487 source.n177 source.n175 0.974638
R488 source.n209 source.n177 0.974638
R489 source.n243 source.n241 0.974638
R490 source.n245 source.n243 0.974638
R491 source.n247 source.n245 0.974638
R492 source.n279 source.n247 0.974638
R493 source.n101 source.n69 0.470328
R494 source.n241 source.n209 0.470328
R495 source.n260 source.n259 0.388379
R496 source.n222 source.n221 0.388379
R497 source.n190 source.n189 0.388379
R498 source.n152 source.n151 0.388379
R499 source.n12 source.n11 0.388379
R500 source.n50 source.n49 0.388379
R501 source.n82 source.n81 0.388379
R502 source.n120 source.n119 0.388379
R503 source source.n280 0.188
R504 source.n262 source.n261 0.155672
R505 source.n262 source.n253 0.155672
R506 source.n269 source.n253 0.155672
R507 source.n270 source.n269 0.155672
R508 source.n270 source.n249 0.155672
R509 source.n277 source.n249 0.155672
R510 source.n224 source.n223 0.155672
R511 source.n224 source.n215 0.155672
R512 source.n231 source.n215 0.155672
R513 source.n232 source.n231 0.155672
R514 source.n232 source.n211 0.155672
R515 source.n239 source.n211 0.155672
R516 source.n192 source.n191 0.155672
R517 source.n192 source.n183 0.155672
R518 source.n199 source.n183 0.155672
R519 source.n200 source.n199 0.155672
R520 source.n200 source.n179 0.155672
R521 source.n207 source.n179 0.155672
R522 source.n154 source.n153 0.155672
R523 source.n154 source.n145 0.155672
R524 source.n161 source.n145 0.155672
R525 source.n162 source.n161 0.155672
R526 source.n162 source.n141 0.155672
R527 source.n169 source.n141 0.155672
R528 source.n29 source.n1 0.155672
R529 source.n22 source.n1 0.155672
R530 source.n22 source.n21 0.155672
R531 source.n21 source.n5 0.155672
R532 source.n14 source.n5 0.155672
R533 source.n14 source.n13 0.155672
R534 source.n67 source.n39 0.155672
R535 source.n60 source.n39 0.155672
R536 source.n60 source.n59 0.155672
R537 source.n59 source.n43 0.155672
R538 source.n52 source.n43 0.155672
R539 source.n52 source.n51 0.155672
R540 source.n99 source.n71 0.155672
R541 source.n92 source.n71 0.155672
R542 source.n92 source.n91 0.155672
R543 source.n91 source.n75 0.155672
R544 source.n84 source.n75 0.155672
R545 source.n84 source.n83 0.155672
R546 source.n137 source.n109 0.155672
R547 source.n130 source.n109 0.155672
R548 source.n130 source.n129 0.155672
R549 source.n129 source.n113 0.155672
R550 source.n122 source.n113 0.155672
R551 source.n122 source.n121 0.155672
R552 minus.n5 minus.t8 250.877
R553 minus.n27 minus.t7 250.877
R554 minus.n6 minus.t5 229.855
R555 minus.n7 minus.t3 229.855
R556 minus.n3 minus.t11 229.855
R557 minus.n13 minus.t12 229.855
R558 minus.n1 minus.t9 229.855
R559 minus.n18 minus.t6 229.855
R560 minus.n20 minus.t13 229.855
R561 minus.n28 minus.t0 229.855
R562 minus.n29 minus.t2 229.855
R563 minus.n25 minus.t15 229.855
R564 minus.n35 minus.t4 229.855
R565 minus.n23 minus.t14 229.855
R566 minus.n40 minus.t1 229.855
R567 minus.n42 minus.t10 229.855
R568 minus.n21 minus.n20 161.3
R569 minus.n19 minus.n0 161.3
R570 minus.n15 minus.n14 161.3
R571 minus.n13 minus.n2 161.3
R572 minus.n12 minus.n11 161.3
R573 minus.n10 minus.n3 161.3
R574 minus.n9 minus.n8 161.3
R575 minus.n43 minus.n42 161.3
R576 minus.n41 minus.n22 161.3
R577 minus.n37 minus.n36 161.3
R578 minus.n35 minus.n24 161.3
R579 minus.n34 minus.n33 161.3
R580 minus.n32 minus.n25 161.3
R581 minus.n31 minus.n30 161.3
R582 minus.n18 minus.n17 80.6037
R583 minus.n16 minus.n1 80.6037
R584 minus.n7 minus.n4 80.6037
R585 minus.n40 minus.n39 80.6037
R586 minus.n38 minus.n23 80.6037
R587 minus.n29 minus.n26 80.6037
R588 minus.n7 minus.n6 48.2005
R589 minus.n18 minus.n1 48.2005
R590 minus.n29 minus.n28 48.2005
R591 minus.n40 minus.n23 48.2005
R592 minus.n8 minus.n7 43.0884
R593 minus.n14 minus.n1 43.0884
R594 minus.n30 minus.n29 43.0884
R595 minus.n36 minus.n23 43.0884
R596 minus.n19 minus.n18 40.1672
R597 minus.n41 minus.n40 40.1672
R598 minus.n44 minus.n21 35.1482
R599 minus.n5 minus.n4 31.6481
R600 minus.n27 minus.n26 31.6481
R601 minus.n13 minus.n12 24.1005
R602 minus.n12 minus.n3 24.1005
R603 minus.n34 minus.n25 24.1005
R604 minus.n35 minus.n34 24.1005
R605 minus.n6 minus.n5 17.444
R606 minus.n28 minus.n27 17.444
R607 minus.n20 minus.n19 8.03383
R608 minus.n42 minus.n41 8.03383
R609 minus.n44 minus.n43 6.6558
R610 minus.n8 minus.n3 5.11262
R611 minus.n14 minus.n13 5.11262
R612 minus.n30 minus.n25 5.11262
R613 minus.n36 minus.n35 5.11262
R614 minus.n17 minus.n16 0.380177
R615 minus.n39 minus.n38 0.380177
R616 minus.n17 minus.n0 0.285035
R617 minus.n16 minus.n15 0.285035
R618 minus.n9 minus.n4 0.285035
R619 minus.n31 minus.n26 0.285035
R620 minus.n38 minus.n37 0.285035
R621 minus.n39 minus.n22 0.285035
R622 minus.n21 minus.n0 0.189894
R623 minus.n15 minus.n2 0.189894
R624 minus.n11 minus.n2 0.189894
R625 minus.n11 minus.n10 0.189894
R626 minus.n10 minus.n9 0.189894
R627 minus.n32 minus.n31 0.189894
R628 minus.n33 minus.n32 0.189894
R629 minus.n33 minus.n24 0.189894
R630 minus.n37 minus.n24 0.189894
R631 minus.n43 minus.n22 0.189894
R632 minus minus.n44 0.188
R633 drain_right.n5 drain_right.n3 68.1648
R634 drain_right.n2 drain_right.n0 68.1648
R635 drain_right.n9 drain_right.n7 68.1648
R636 drain_right.n9 drain_right.n8 67.1908
R637 drain_right.n11 drain_right.n10 67.1908
R638 drain_right.n13 drain_right.n12 67.1908
R639 drain_right.n5 drain_right.n4 67.1907
R640 drain_right.n2 drain_right.n1 67.1907
R641 drain_right drain_right.n6 28.6003
R642 drain_right drain_right.n13 6.62735
R643 drain_right.n3 drain_right.t14 3.3005
R644 drain_right.n3 drain_right.t5 3.3005
R645 drain_right.n4 drain_right.t11 3.3005
R646 drain_right.n4 drain_right.t1 3.3005
R647 drain_right.n1 drain_right.t13 3.3005
R648 drain_right.n1 drain_right.t0 3.3005
R649 drain_right.n0 drain_right.t8 3.3005
R650 drain_right.n0 drain_right.t15 3.3005
R651 drain_right.n7 drain_right.t10 3.3005
R652 drain_right.n7 drain_right.t7 3.3005
R653 drain_right.n8 drain_right.t4 3.3005
R654 drain_right.n8 drain_right.t12 3.3005
R655 drain_right.n10 drain_right.t6 3.3005
R656 drain_right.n10 drain_right.t3 3.3005
R657 drain_right.n12 drain_right.t2 3.3005
R658 drain_right.n12 drain_right.t9 3.3005
R659 drain_right.n13 drain_right.n11 0.974638
R660 drain_right.n11 drain_right.n9 0.974638
R661 drain_right.n6 drain_right.n5 0.432223
R662 drain_right.n6 drain_right.n2 0.432223
C0 plus drain_left 6.06606f
C1 drain_left source 11.0903f
C2 drain_left minus 0.173489f
C3 plus drain_right 0.430381f
C4 drain_right source 11.093f
C5 minus drain_right 5.79269f
C6 plus source 6.25099f
C7 plus minus 5.46491f
C8 minus source 6.23698f
C9 drain_left drain_right 1.44945f
C10 drain_right a_n2750_n2088# 5.8041f
C11 drain_left a_n2750_n2088# 6.20058f
C12 source a_n2750_n2088# 5.760413f
C13 minus a_n2750_n2088# 10.488028f
C14 plus a_n2750_n2088# 11.94229f
C15 drain_right.t8 a_n2750_n2088# 0.125155f
C16 drain_right.t15 a_n2750_n2088# 0.125155f
C17 drain_right.n0 a_n2750_n2088# 1.04937f
C18 drain_right.t13 a_n2750_n2088# 0.125155f
C19 drain_right.t0 a_n2750_n2088# 0.125155f
C20 drain_right.n1 a_n2750_n2088# 1.04379f
C21 drain_right.n2 a_n2750_n2088# 0.720236f
C22 drain_right.t14 a_n2750_n2088# 0.125155f
C23 drain_right.t5 a_n2750_n2088# 0.125155f
C24 drain_right.n3 a_n2750_n2088# 1.04937f
C25 drain_right.t11 a_n2750_n2088# 0.125155f
C26 drain_right.t1 a_n2750_n2088# 0.125155f
C27 drain_right.n4 a_n2750_n2088# 1.04379f
C28 drain_right.n5 a_n2750_n2088# 0.720236f
C29 drain_right.n6 a_n2750_n2088# 1.16988f
C30 drain_right.t10 a_n2750_n2088# 0.125155f
C31 drain_right.t7 a_n2750_n2088# 0.125155f
C32 drain_right.n7 a_n2750_n2088# 1.04937f
C33 drain_right.t4 a_n2750_n2088# 0.125155f
C34 drain_right.t12 a_n2750_n2088# 0.125155f
C35 drain_right.n8 a_n2750_n2088# 1.0438f
C36 drain_right.n9 a_n2750_n2088# 0.764948f
C37 drain_right.t6 a_n2750_n2088# 0.125155f
C38 drain_right.t3 a_n2750_n2088# 0.125155f
C39 drain_right.n10 a_n2750_n2088# 1.0438f
C40 drain_right.n11 a_n2750_n2088# 0.379947f
C41 drain_right.t2 a_n2750_n2088# 0.125155f
C42 drain_right.t9 a_n2750_n2088# 0.125155f
C43 drain_right.n12 a_n2750_n2088# 1.0438f
C44 drain_right.n13 a_n2750_n2088# 0.616641f
C45 minus.n0 a_n2750_n2088# 0.052687f
C46 minus.t9 a_n2750_n2088# 0.549732f
C47 minus.n1 a_n2750_n2088# 0.261688f
C48 minus.t6 a_n2750_n2088# 0.549732f
C49 minus.n2 a_n2750_n2088# 0.039485f
C50 minus.t11 a_n2750_n2088# 0.549732f
C51 minus.n3 a_n2750_n2088# 0.250416f
C52 minus.n4 a_n2750_n2088# 0.226464f
C53 minus.t8 a_n2750_n2088# 0.571006f
C54 minus.n5 a_n2750_n2088# 0.236129f
C55 minus.t5 a_n2750_n2088# 0.549732f
C56 minus.n6 a_n2750_n2088# 0.261997f
C57 minus.t3 a_n2750_n2088# 0.549732f
C58 minus.n7 a_n2750_n2088# 0.261688f
C59 minus.n8 a_n2750_n2088# 0.00896f
C60 minus.n9 a_n2750_n2088# 0.052687f
C61 minus.n10 a_n2750_n2088# 0.039485f
C62 minus.n11 a_n2750_n2088# 0.039485f
C63 minus.n12 a_n2750_n2088# 0.00896f
C64 minus.t12 a_n2750_n2088# 0.549732f
C65 minus.n13 a_n2750_n2088# 0.250416f
C66 minus.n14 a_n2750_n2088# 0.00896f
C67 minus.n15 a_n2750_n2088# 0.052687f
C68 minus.n16 a_n2750_n2088# 0.065767f
C69 minus.n17 a_n2750_n2088# 0.065767f
C70 minus.n18 a_n2750_n2088# 0.261201f
C71 minus.n19 a_n2750_n2088# 0.00896f
C72 minus.t13 a_n2750_n2088# 0.549732f
C73 minus.n20 a_n2750_n2088# 0.246886f
C74 minus.n21 a_n2750_n2088# 1.33742f
C75 minus.n22 a_n2750_n2088# 0.052687f
C76 minus.t14 a_n2750_n2088# 0.549732f
C77 minus.n23 a_n2750_n2088# 0.261688f
C78 minus.n24 a_n2750_n2088# 0.039485f
C79 minus.t15 a_n2750_n2088# 0.549732f
C80 minus.n25 a_n2750_n2088# 0.250416f
C81 minus.n26 a_n2750_n2088# 0.226464f
C82 minus.t7 a_n2750_n2088# 0.571006f
C83 minus.n27 a_n2750_n2088# 0.236129f
C84 minus.t0 a_n2750_n2088# 0.549732f
C85 minus.n28 a_n2750_n2088# 0.261997f
C86 minus.t2 a_n2750_n2088# 0.549732f
C87 minus.n29 a_n2750_n2088# 0.261688f
C88 minus.n30 a_n2750_n2088# 0.00896f
C89 minus.n31 a_n2750_n2088# 0.052687f
C90 minus.n32 a_n2750_n2088# 0.039485f
C91 minus.n33 a_n2750_n2088# 0.039485f
C92 minus.n34 a_n2750_n2088# 0.00896f
C93 minus.t4 a_n2750_n2088# 0.549732f
C94 minus.n35 a_n2750_n2088# 0.250416f
C95 minus.n36 a_n2750_n2088# 0.00896f
C96 minus.n37 a_n2750_n2088# 0.052687f
C97 minus.n38 a_n2750_n2088# 0.065767f
C98 minus.n39 a_n2750_n2088# 0.065767f
C99 minus.t1 a_n2750_n2088# 0.549732f
C100 minus.n40 a_n2750_n2088# 0.261201f
C101 minus.n41 a_n2750_n2088# 0.00896f
C102 minus.t10 a_n2750_n2088# 0.549732f
C103 minus.n42 a_n2750_n2088# 0.246886f
C104 minus.n43 a_n2750_n2088# 0.272529f
C105 minus.n44 a_n2750_n2088# 1.62431f
C106 source.n0 a_n2750_n2088# 0.034947f
C107 source.n1 a_n2750_n2088# 0.024863f
C108 source.n2 a_n2750_n2088# 0.01336f
C109 source.n3 a_n2750_n2088# 0.031578f
C110 source.n4 a_n2750_n2088# 0.014146f
C111 source.n5 a_n2750_n2088# 0.024863f
C112 source.n6 a_n2750_n2088# 0.01336f
C113 source.n7 a_n2750_n2088# 0.031578f
C114 source.n8 a_n2750_n2088# 0.014146f
C115 source.n9 a_n2750_n2088# 0.106395f
C116 source.t17 a_n2750_n2088# 0.051469f
C117 source.n10 a_n2750_n2088# 0.023684f
C118 source.n11 a_n2750_n2088# 0.018653f
C119 source.n12 a_n2750_n2088# 0.01336f
C120 source.n13 a_n2750_n2088# 0.591584f
C121 source.n14 a_n2750_n2088# 0.024863f
C122 source.n15 a_n2750_n2088# 0.01336f
C123 source.n16 a_n2750_n2088# 0.014146f
C124 source.n17 a_n2750_n2088# 0.031578f
C125 source.n18 a_n2750_n2088# 0.031578f
C126 source.n19 a_n2750_n2088# 0.014146f
C127 source.n20 a_n2750_n2088# 0.01336f
C128 source.n21 a_n2750_n2088# 0.024863f
C129 source.n22 a_n2750_n2088# 0.024863f
C130 source.n23 a_n2750_n2088# 0.01336f
C131 source.n24 a_n2750_n2088# 0.014146f
C132 source.n25 a_n2750_n2088# 0.031578f
C133 source.n26 a_n2750_n2088# 0.068362f
C134 source.n27 a_n2750_n2088# 0.014146f
C135 source.n28 a_n2750_n2088# 0.01336f
C136 source.n29 a_n2750_n2088# 0.057469f
C137 source.n30 a_n2750_n2088# 0.038251f
C138 source.n31 a_n2750_n2088# 0.661296f
C139 source.t14 a_n2750_n2088# 0.117884f
C140 source.t16 a_n2750_n2088# 0.117884f
C141 source.n32 a_n2750_n2088# 0.918086f
C142 source.n33 a_n2750_n2088# 0.389146f
C143 source.t13 a_n2750_n2088# 0.117884f
C144 source.t11 a_n2750_n2088# 0.117884f
C145 source.n34 a_n2750_n2088# 0.918086f
C146 source.n35 a_n2750_n2088# 0.389146f
C147 source.t10 a_n2750_n2088# 0.117884f
C148 source.t12 a_n2750_n2088# 0.117884f
C149 source.n36 a_n2750_n2088# 0.918086f
C150 source.n37 a_n2750_n2088# 0.389146f
C151 source.n38 a_n2750_n2088# 0.034947f
C152 source.n39 a_n2750_n2088# 0.024863f
C153 source.n40 a_n2750_n2088# 0.01336f
C154 source.n41 a_n2750_n2088# 0.031578f
C155 source.n42 a_n2750_n2088# 0.014146f
C156 source.n43 a_n2750_n2088# 0.024863f
C157 source.n44 a_n2750_n2088# 0.01336f
C158 source.n45 a_n2750_n2088# 0.031578f
C159 source.n46 a_n2750_n2088# 0.014146f
C160 source.n47 a_n2750_n2088# 0.106395f
C161 source.t9 a_n2750_n2088# 0.051469f
C162 source.n48 a_n2750_n2088# 0.023684f
C163 source.n49 a_n2750_n2088# 0.018653f
C164 source.n50 a_n2750_n2088# 0.01336f
C165 source.n51 a_n2750_n2088# 0.591584f
C166 source.n52 a_n2750_n2088# 0.024863f
C167 source.n53 a_n2750_n2088# 0.01336f
C168 source.n54 a_n2750_n2088# 0.014146f
C169 source.n55 a_n2750_n2088# 0.031578f
C170 source.n56 a_n2750_n2088# 0.031578f
C171 source.n57 a_n2750_n2088# 0.014146f
C172 source.n58 a_n2750_n2088# 0.01336f
C173 source.n59 a_n2750_n2088# 0.024863f
C174 source.n60 a_n2750_n2088# 0.024863f
C175 source.n61 a_n2750_n2088# 0.01336f
C176 source.n62 a_n2750_n2088# 0.014146f
C177 source.n63 a_n2750_n2088# 0.031578f
C178 source.n64 a_n2750_n2088# 0.068362f
C179 source.n65 a_n2750_n2088# 0.014146f
C180 source.n66 a_n2750_n2088# 0.01336f
C181 source.n67 a_n2750_n2088# 0.057469f
C182 source.n68 a_n2750_n2088# 0.038251f
C183 source.n69 a_n2750_n2088# 0.136915f
C184 source.n70 a_n2750_n2088# 0.034947f
C185 source.n71 a_n2750_n2088# 0.024863f
C186 source.n72 a_n2750_n2088# 0.01336f
C187 source.n73 a_n2750_n2088# 0.031578f
C188 source.n74 a_n2750_n2088# 0.014146f
C189 source.n75 a_n2750_n2088# 0.024863f
C190 source.n76 a_n2750_n2088# 0.01336f
C191 source.n77 a_n2750_n2088# 0.031578f
C192 source.n78 a_n2750_n2088# 0.014146f
C193 source.n79 a_n2750_n2088# 0.106395f
C194 source.t27 a_n2750_n2088# 0.051469f
C195 source.n80 a_n2750_n2088# 0.023684f
C196 source.n81 a_n2750_n2088# 0.018653f
C197 source.n82 a_n2750_n2088# 0.01336f
C198 source.n83 a_n2750_n2088# 0.591584f
C199 source.n84 a_n2750_n2088# 0.024863f
C200 source.n85 a_n2750_n2088# 0.01336f
C201 source.n86 a_n2750_n2088# 0.014146f
C202 source.n87 a_n2750_n2088# 0.031578f
C203 source.n88 a_n2750_n2088# 0.031578f
C204 source.n89 a_n2750_n2088# 0.014146f
C205 source.n90 a_n2750_n2088# 0.01336f
C206 source.n91 a_n2750_n2088# 0.024863f
C207 source.n92 a_n2750_n2088# 0.024863f
C208 source.n93 a_n2750_n2088# 0.01336f
C209 source.n94 a_n2750_n2088# 0.014146f
C210 source.n95 a_n2750_n2088# 0.031578f
C211 source.n96 a_n2750_n2088# 0.068362f
C212 source.n97 a_n2750_n2088# 0.014146f
C213 source.n98 a_n2750_n2088# 0.01336f
C214 source.n99 a_n2750_n2088# 0.057469f
C215 source.n100 a_n2750_n2088# 0.038251f
C216 source.n101 a_n2750_n2088# 0.136915f
C217 source.t6 a_n2750_n2088# 0.117884f
C218 source.t29 a_n2750_n2088# 0.117884f
C219 source.n102 a_n2750_n2088# 0.918086f
C220 source.n103 a_n2750_n2088# 0.389146f
C221 source.t0 a_n2750_n2088# 0.117884f
C222 source.t2 a_n2750_n2088# 0.117884f
C223 source.n104 a_n2750_n2088# 0.918086f
C224 source.n105 a_n2750_n2088# 0.389146f
C225 source.t24 a_n2750_n2088# 0.117884f
C226 source.t28 a_n2750_n2088# 0.117884f
C227 source.n106 a_n2750_n2088# 0.918086f
C228 source.n107 a_n2750_n2088# 0.389146f
C229 source.n108 a_n2750_n2088# 0.034947f
C230 source.n109 a_n2750_n2088# 0.024863f
C231 source.n110 a_n2750_n2088# 0.01336f
C232 source.n111 a_n2750_n2088# 0.031578f
C233 source.n112 a_n2750_n2088# 0.014146f
C234 source.n113 a_n2750_n2088# 0.024863f
C235 source.n114 a_n2750_n2088# 0.01336f
C236 source.n115 a_n2750_n2088# 0.031578f
C237 source.n116 a_n2750_n2088# 0.014146f
C238 source.n117 a_n2750_n2088# 0.106395f
C239 source.t26 a_n2750_n2088# 0.051469f
C240 source.n118 a_n2750_n2088# 0.023684f
C241 source.n119 a_n2750_n2088# 0.018653f
C242 source.n120 a_n2750_n2088# 0.01336f
C243 source.n121 a_n2750_n2088# 0.591584f
C244 source.n122 a_n2750_n2088# 0.024863f
C245 source.n123 a_n2750_n2088# 0.01336f
C246 source.n124 a_n2750_n2088# 0.014146f
C247 source.n125 a_n2750_n2088# 0.031578f
C248 source.n126 a_n2750_n2088# 0.031578f
C249 source.n127 a_n2750_n2088# 0.014146f
C250 source.n128 a_n2750_n2088# 0.01336f
C251 source.n129 a_n2750_n2088# 0.024863f
C252 source.n130 a_n2750_n2088# 0.024863f
C253 source.n131 a_n2750_n2088# 0.01336f
C254 source.n132 a_n2750_n2088# 0.014146f
C255 source.n133 a_n2750_n2088# 0.031578f
C256 source.n134 a_n2750_n2088# 0.068362f
C257 source.n135 a_n2750_n2088# 0.014146f
C258 source.n136 a_n2750_n2088# 0.01336f
C259 source.n137 a_n2750_n2088# 0.057469f
C260 source.n138 a_n2750_n2088# 0.038251f
C261 source.n139 a_n2750_n2088# 0.991368f
C262 source.n140 a_n2750_n2088# 0.034947f
C263 source.n141 a_n2750_n2088# 0.024863f
C264 source.n142 a_n2750_n2088# 0.01336f
C265 source.n143 a_n2750_n2088# 0.031578f
C266 source.n144 a_n2750_n2088# 0.014146f
C267 source.n145 a_n2750_n2088# 0.024863f
C268 source.n146 a_n2750_n2088# 0.01336f
C269 source.n147 a_n2750_n2088# 0.031578f
C270 source.n148 a_n2750_n2088# 0.014146f
C271 source.n149 a_n2750_n2088# 0.106395f
C272 source.t15 a_n2750_n2088# 0.051469f
C273 source.n150 a_n2750_n2088# 0.023684f
C274 source.n151 a_n2750_n2088# 0.018653f
C275 source.n152 a_n2750_n2088# 0.01336f
C276 source.n153 a_n2750_n2088# 0.591584f
C277 source.n154 a_n2750_n2088# 0.024863f
C278 source.n155 a_n2750_n2088# 0.01336f
C279 source.n156 a_n2750_n2088# 0.014146f
C280 source.n157 a_n2750_n2088# 0.031578f
C281 source.n158 a_n2750_n2088# 0.031578f
C282 source.n159 a_n2750_n2088# 0.014146f
C283 source.n160 a_n2750_n2088# 0.01336f
C284 source.n161 a_n2750_n2088# 0.024863f
C285 source.n162 a_n2750_n2088# 0.024863f
C286 source.n163 a_n2750_n2088# 0.01336f
C287 source.n164 a_n2750_n2088# 0.014146f
C288 source.n165 a_n2750_n2088# 0.031578f
C289 source.n166 a_n2750_n2088# 0.068362f
C290 source.n167 a_n2750_n2088# 0.014146f
C291 source.n168 a_n2750_n2088# 0.01336f
C292 source.n169 a_n2750_n2088# 0.057469f
C293 source.n170 a_n2750_n2088# 0.038251f
C294 source.n171 a_n2750_n2088# 0.991368f
C295 source.t22 a_n2750_n2088# 0.117884f
C296 source.t18 a_n2750_n2088# 0.117884f
C297 source.n172 a_n2750_n2088# 0.91808f
C298 source.n173 a_n2750_n2088# 0.389153f
C299 source.t20 a_n2750_n2088# 0.117884f
C300 source.t8 a_n2750_n2088# 0.117884f
C301 source.n174 a_n2750_n2088# 0.91808f
C302 source.n175 a_n2750_n2088# 0.389153f
C303 source.t21 a_n2750_n2088# 0.117884f
C304 source.t23 a_n2750_n2088# 0.117884f
C305 source.n176 a_n2750_n2088# 0.91808f
C306 source.n177 a_n2750_n2088# 0.389153f
C307 source.n178 a_n2750_n2088# 0.034947f
C308 source.n179 a_n2750_n2088# 0.024863f
C309 source.n180 a_n2750_n2088# 0.01336f
C310 source.n181 a_n2750_n2088# 0.031578f
C311 source.n182 a_n2750_n2088# 0.014146f
C312 source.n183 a_n2750_n2088# 0.024863f
C313 source.n184 a_n2750_n2088# 0.01336f
C314 source.n185 a_n2750_n2088# 0.031578f
C315 source.n186 a_n2750_n2088# 0.014146f
C316 source.n187 a_n2750_n2088# 0.106395f
C317 source.t19 a_n2750_n2088# 0.051469f
C318 source.n188 a_n2750_n2088# 0.023684f
C319 source.n189 a_n2750_n2088# 0.018653f
C320 source.n190 a_n2750_n2088# 0.01336f
C321 source.n191 a_n2750_n2088# 0.591584f
C322 source.n192 a_n2750_n2088# 0.024863f
C323 source.n193 a_n2750_n2088# 0.01336f
C324 source.n194 a_n2750_n2088# 0.014146f
C325 source.n195 a_n2750_n2088# 0.031578f
C326 source.n196 a_n2750_n2088# 0.031578f
C327 source.n197 a_n2750_n2088# 0.014146f
C328 source.n198 a_n2750_n2088# 0.01336f
C329 source.n199 a_n2750_n2088# 0.024863f
C330 source.n200 a_n2750_n2088# 0.024863f
C331 source.n201 a_n2750_n2088# 0.01336f
C332 source.n202 a_n2750_n2088# 0.014146f
C333 source.n203 a_n2750_n2088# 0.031578f
C334 source.n204 a_n2750_n2088# 0.068362f
C335 source.n205 a_n2750_n2088# 0.014146f
C336 source.n206 a_n2750_n2088# 0.01336f
C337 source.n207 a_n2750_n2088# 0.057469f
C338 source.n208 a_n2750_n2088# 0.038251f
C339 source.n209 a_n2750_n2088# 0.136915f
C340 source.n210 a_n2750_n2088# 0.034947f
C341 source.n211 a_n2750_n2088# 0.024863f
C342 source.n212 a_n2750_n2088# 0.01336f
C343 source.n213 a_n2750_n2088# 0.031578f
C344 source.n214 a_n2750_n2088# 0.014146f
C345 source.n215 a_n2750_n2088# 0.024863f
C346 source.n216 a_n2750_n2088# 0.01336f
C347 source.n217 a_n2750_n2088# 0.031578f
C348 source.n218 a_n2750_n2088# 0.014146f
C349 source.n219 a_n2750_n2088# 0.106395f
C350 source.t31 a_n2750_n2088# 0.051469f
C351 source.n220 a_n2750_n2088# 0.023684f
C352 source.n221 a_n2750_n2088# 0.018653f
C353 source.n222 a_n2750_n2088# 0.01336f
C354 source.n223 a_n2750_n2088# 0.591584f
C355 source.n224 a_n2750_n2088# 0.024863f
C356 source.n225 a_n2750_n2088# 0.01336f
C357 source.n226 a_n2750_n2088# 0.014146f
C358 source.n227 a_n2750_n2088# 0.031578f
C359 source.n228 a_n2750_n2088# 0.031578f
C360 source.n229 a_n2750_n2088# 0.014146f
C361 source.n230 a_n2750_n2088# 0.01336f
C362 source.n231 a_n2750_n2088# 0.024863f
C363 source.n232 a_n2750_n2088# 0.024863f
C364 source.n233 a_n2750_n2088# 0.01336f
C365 source.n234 a_n2750_n2088# 0.014146f
C366 source.n235 a_n2750_n2088# 0.031578f
C367 source.n236 a_n2750_n2088# 0.068362f
C368 source.n237 a_n2750_n2088# 0.014146f
C369 source.n238 a_n2750_n2088# 0.01336f
C370 source.n239 a_n2750_n2088# 0.057469f
C371 source.n240 a_n2750_n2088# 0.038251f
C372 source.n241 a_n2750_n2088# 0.136915f
C373 source.t25 a_n2750_n2088# 0.117884f
C374 source.t4 a_n2750_n2088# 0.117884f
C375 source.n242 a_n2750_n2088# 0.91808f
C376 source.n243 a_n2750_n2088# 0.389153f
C377 source.t3 a_n2750_n2088# 0.117884f
C378 source.t30 a_n2750_n2088# 0.117884f
C379 source.n244 a_n2750_n2088# 0.91808f
C380 source.n245 a_n2750_n2088# 0.389153f
C381 source.t5 a_n2750_n2088# 0.117884f
C382 source.t1 a_n2750_n2088# 0.117884f
C383 source.n246 a_n2750_n2088# 0.91808f
C384 source.n247 a_n2750_n2088# 0.389153f
C385 source.n248 a_n2750_n2088# 0.034947f
C386 source.n249 a_n2750_n2088# 0.024863f
C387 source.n250 a_n2750_n2088# 0.01336f
C388 source.n251 a_n2750_n2088# 0.031578f
C389 source.n252 a_n2750_n2088# 0.014146f
C390 source.n253 a_n2750_n2088# 0.024863f
C391 source.n254 a_n2750_n2088# 0.01336f
C392 source.n255 a_n2750_n2088# 0.031578f
C393 source.n256 a_n2750_n2088# 0.014146f
C394 source.n257 a_n2750_n2088# 0.106395f
C395 source.t7 a_n2750_n2088# 0.051469f
C396 source.n258 a_n2750_n2088# 0.023684f
C397 source.n259 a_n2750_n2088# 0.018653f
C398 source.n260 a_n2750_n2088# 0.01336f
C399 source.n261 a_n2750_n2088# 0.591584f
C400 source.n262 a_n2750_n2088# 0.024863f
C401 source.n263 a_n2750_n2088# 0.01336f
C402 source.n264 a_n2750_n2088# 0.014146f
C403 source.n265 a_n2750_n2088# 0.031578f
C404 source.n266 a_n2750_n2088# 0.031578f
C405 source.n267 a_n2750_n2088# 0.014146f
C406 source.n268 a_n2750_n2088# 0.01336f
C407 source.n269 a_n2750_n2088# 0.024863f
C408 source.n270 a_n2750_n2088# 0.024863f
C409 source.n271 a_n2750_n2088# 0.01336f
C410 source.n272 a_n2750_n2088# 0.014146f
C411 source.n273 a_n2750_n2088# 0.031578f
C412 source.n274 a_n2750_n2088# 0.068362f
C413 source.n275 a_n2750_n2088# 0.014146f
C414 source.n276 a_n2750_n2088# 0.01336f
C415 source.n277 a_n2750_n2088# 0.057469f
C416 source.n278 a_n2750_n2088# 0.038251f
C417 source.n279 a_n2750_n2088# 0.304478f
C418 source.n280 a_n2750_n2088# 1.03465f
C419 drain_left.t11 a_n2750_n2088# 0.126603f
C420 drain_left.t7 a_n2750_n2088# 0.126603f
C421 drain_left.n0 a_n2750_n2088# 1.06152f
C422 drain_left.t5 a_n2750_n2088# 0.126603f
C423 drain_left.t1 a_n2750_n2088# 0.126603f
C424 drain_left.n1 a_n2750_n2088# 1.05587f
C425 drain_left.n2 a_n2750_n2088# 0.728569f
C426 drain_left.t8 a_n2750_n2088# 0.126603f
C427 drain_left.t0 a_n2750_n2088# 0.126603f
C428 drain_left.n3 a_n2750_n2088# 1.06152f
C429 drain_left.t13 a_n2750_n2088# 0.126603f
C430 drain_left.t2 a_n2750_n2088# 0.126603f
C431 drain_left.n4 a_n2750_n2088# 1.05587f
C432 drain_left.n5 a_n2750_n2088# 0.728569f
C433 drain_left.n6 a_n2750_n2088# 1.23689f
C434 drain_left.t6 a_n2750_n2088# 0.126603f
C435 drain_left.t3 a_n2750_n2088# 0.126603f
C436 drain_left.n7 a_n2750_n2088# 1.06152f
C437 drain_left.t10 a_n2750_n2088# 0.126603f
C438 drain_left.t15 a_n2750_n2088# 0.126603f
C439 drain_left.n8 a_n2750_n2088# 1.05587f
C440 drain_left.n9 a_n2750_n2088# 0.773794f
C441 drain_left.t9 a_n2750_n2088# 0.126603f
C442 drain_left.t4 a_n2750_n2088# 0.126603f
C443 drain_left.n10 a_n2750_n2088# 1.05587f
C444 drain_left.n11 a_n2750_n2088# 0.384343f
C445 drain_left.t12 a_n2750_n2088# 0.126603f
C446 drain_left.t14 a_n2750_n2088# 0.126603f
C447 drain_left.n12 a_n2750_n2088# 1.05587f
C448 drain_left.n13 a_n2750_n2088# 0.62378f
C449 plus.n0 a_n2750_n2088# 0.054139f
C450 plus.t6 a_n2750_n2088# 0.564875f
C451 plus.t7 a_n2750_n2088# 0.564875f
C452 plus.n1 a_n2750_n2088# 0.067578f
C453 plus.t9 a_n2750_n2088# 0.564875f
C454 plus.n2 a_n2750_n2088# 0.067578f
C455 plus.t12 a_n2750_n2088# 0.564875f
C456 plus.n3 a_n2750_n2088# 0.257314f
C457 plus.n4 a_n2750_n2088# 0.040572f
C458 plus.t10 a_n2750_n2088# 0.564875f
C459 plus.t11 a_n2750_n2088# 0.564875f
C460 plus.n5 a_n2750_n2088# 0.268897f
C461 plus.t13 a_n2750_n2088# 0.564875f
C462 plus.n6 a_n2750_n2088# 0.269214f
C463 plus.t14 a_n2750_n2088# 0.586735f
C464 plus.n7 a_n2750_n2088# 0.242634f
C465 plus.n8 a_n2750_n2088# 0.232702f
C466 plus.n9 a_n2750_n2088# 0.054139f
C467 plus.n10 a_n2750_n2088# 0.009207f
C468 plus.n11 a_n2750_n2088# 0.257314f
C469 plus.n12 a_n2750_n2088# 0.009207f
C470 plus.n13 a_n2750_n2088# 0.040572f
C471 plus.n14 a_n2750_n2088# 0.040572f
C472 plus.n15 a_n2750_n2088# 0.054139f
C473 plus.n16 a_n2750_n2088# 0.009207f
C474 plus.n17 a_n2750_n2088# 0.268897f
C475 plus.n18 a_n2750_n2088# 0.268396f
C476 plus.n19 a_n2750_n2088# 0.009207f
C477 plus.n20 a_n2750_n2088# 0.253686f
C478 plus.n21 a_n2750_n2088# 0.363114f
C479 plus.n22 a_n2750_n2088# 0.054139f
C480 plus.t8 a_n2750_n2088# 0.564875f
C481 plus.n23 a_n2750_n2088# 0.067578f
C482 plus.t1 a_n2750_n2088# 0.564875f
C483 plus.n24 a_n2750_n2088# 0.067578f
C484 plus.t5 a_n2750_n2088# 0.564875f
C485 plus.t3 a_n2750_n2088# 0.564875f
C486 plus.n25 a_n2750_n2088# 0.257314f
C487 plus.n26 a_n2750_n2088# 0.040572f
C488 plus.t15 a_n2750_n2088# 0.564875f
C489 plus.t2 a_n2750_n2088# 0.564875f
C490 plus.n27 a_n2750_n2088# 0.268897f
C491 plus.t0 a_n2750_n2088# 0.564875f
C492 plus.n28 a_n2750_n2088# 0.269214f
C493 plus.t4 a_n2750_n2088# 0.586735f
C494 plus.n29 a_n2750_n2088# 0.242634f
C495 plus.n30 a_n2750_n2088# 0.232702f
C496 plus.n31 a_n2750_n2088# 0.054139f
C497 plus.n32 a_n2750_n2088# 0.009207f
C498 plus.n33 a_n2750_n2088# 0.257314f
C499 plus.n34 a_n2750_n2088# 0.009207f
C500 plus.n35 a_n2750_n2088# 0.040572f
C501 plus.n36 a_n2750_n2088# 0.040572f
C502 plus.n37 a_n2750_n2088# 0.054139f
C503 plus.n38 a_n2750_n2088# 0.009207f
C504 plus.n39 a_n2750_n2088# 0.268897f
C505 plus.n40 a_n2750_n2088# 0.268396f
C506 plus.n41 a_n2750_n2088# 0.009207f
C507 plus.n42 a_n2750_n2088# 0.253686f
C508 plus.n43 a_n2750_n2088# 1.24523f
.ends

