* NGSPICE file created from diffpair550.ext - technology: sky130A

.subckt diffpair550 minus drain_right drain_left source plus
X0 a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X1 drain_right minus source a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.8
X2 drain_left plus source a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.8
X3 drain_left plus source a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.8
X4 a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X5 drain_right minus source a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.8
X6 a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X7 a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# a_n1168_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
.ends

