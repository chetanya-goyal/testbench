* NGSPICE file created from diffpair284.ext - technology: sky130A

.subckt diffpair284 minus drain_right drain_left source plus
X0 a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X1 source.t15 minus.t0 drain_right.t2 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X2 drain_right.t4 minus.t1 source.t14 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X3 source.t13 minus.t2 drain_right.t7 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X4 drain_left.t9 plus.t0 source.t1 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X5 drain_right.t9 minus.t3 source.t12 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X6 drain_right.t6 minus.t4 source.t11 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X7 source.t16 plus.t1 drain_left.t8 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X8 a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X9 drain_left.t7 plus.t2 source.t17 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X10 source.t18 plus.t3 drain_left.t6 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X11 a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X12 drain_right.t1 minus.t5 source.t10 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X13 source.t19 plus.t4 drain_left.t5 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X14 drain_left.t4 plus.t5 source.t0 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X15 source.t5 plus.t6 drain_left.t3 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X16 source.t9 minus.t6 drain_right.t0 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X17 drain_right.t5 minus.t7 source.t8 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X18 source.t7 minus.t8 drain_right.t8 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X19 a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X20 drain_left.t2 plus.t7 source.t2 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X21 drain_right.t3 minus.t9 source.t6 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X22 drain_left.t1 plus.t8 source.t3 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X23 drain_left.t0 plus.t9 source.t4 a_n1712_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
R0 minus.n2 minus.t5 388.748
R1 minus.n14 minus.t7 388.748
R2 minus.n3 minus.t2 367.767
R3 minus.n1 minus.t4 367.767
R4 minus.n9 minus.t8 367.767
R5 minus.n10 minus.t3 367.767
R6 minus.n15 minus.t6 367.767
R7 minus.n13 minus.t1 367.767
R8 minus.n21 minus.t0 367.767
R9 minus.n22 minus.t9 367.767
R10 minus.n11 minus.n10 161.3
R11 minus.n9 minus.n0 161.3
R12 minus.n8 minus.n7 161.3
R13 minus.n6 minus.n1 161.3
R14 minus.n5 minus.n4 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n18 minus.n13 161.3
R19 minus.n17 minus.n16 161.3
R20 minus.n5 minus.n2 70.4033
R21 minus.n17 minus.n14 70.4033
R22 minus.n10 minus.n9 48.2005
R23 minus.n22 minus.n21 48.2005
R24 minus.n4 minus.n1 36.5157
R25 minus.n8 minus.n1 36.5157
R26 minus.n16 minus.n13 36.5157
R27 minus.n20 minus.n13 36.5157
R28 minus.n24 minus.n11 31.1236
R29 minus.n3 minus.n2 20.9576
R30 minus.n15 minus.n14 20.9576
R31 minus.n4 minus.n3 11.6853
R32 minus.n9 minus.n8 11.6853
R33 minus.n16 minus.n15 11.6853
R34 minus.n21 minus.n20 11.6853
R35 minus.n24 minus.n23 6.563
R36 minus.n11 minus.n0 0.189894
R37 minus.n7 minus.n0 0.189894
R38 minus.n7 minus.n6 0.189894
R39 minus.n6 minus.n5 0.189894
R40 minus.n18 minus.n17 0.189894
R41 minus.n19 minus.n18 0.189894
R42 minus.n19 minus.n12 0.189894
R43 minus.n23 minus.n12 0.189894
R44 minus minus.n24 0.188
R45 drain_right.n26 drain_right.n0 289.615
R46 drain_right.n64 drain_right.n38 289.615
R47 drain_right.n11 drain_right.n10 185
R48 drain_right.n8 drain_right.n7 185
R49 drain_right.n17 drain_right.n16 185
R50 drain_right.n19 drain_right.n18 185
R51 drain_right.n4 drain_right.n3 185
R52 drain_right.n25 drain_right.n24 185
R53 drain_right.n27 drain_right.n26 185
R54 drain_right.n65 drain_right.n64 185
R55 drain_right.n63 drain_right.n62 185
R56 drain_right.n42 drain_right.n41 185
R57 drain_right.n57 drain_right.n56 185
R58 drain_right.n55 drain_right.n54 185
R59 drain_right.n46 drain_right.n45 185
R60 drain_right.n49 drain_right.n48 185
R61 drain_right.t5 drain_right.n9 147.661
R62 drain_right.t9 drain_right.n47 147.661
R63 drain_right.n10 drain_right.n7 104.615
R64 drain_right.n17 drain_right.n7 104.615
R65 drain_right.n18 drain_right.n17 104.615
R66 drain_right.n18 drain_right.n3 104.615
R67 drain_right.n25 drain_right.n3 104.615
R68 drain_right.n26 drain_right.n25 104.615
R69 drain_right.n64 drain_right.n63 104.615
R70 drain_right.n63 drain_right.n41 104.615
R71 drain_right.n56 drain_right.n41 104.615
R72 drain_right.n56 drain_right.n55 104.615
R73 drain_right.n55 drain_right.n45 104.615
R74 drain_right.n48 drain_right.n45 104.615
R75 drain_right.n37 drain_right.n35 67.9062
R76 drain_right.n34 drain_right.n33 67.672
R77 drain_right.n37 drain_right.n36 67.1908
R78 drain_right.n32 drain_right.n31 67.1907
R79 drain_right.n10 drain_right.t5 52.3082
R80 drain_right.n48 drain_right.t9 52.3082
R81 drain_right.n32 drain_right.n30 49.5797
R82 drain_right.n69 drain_right.n68 48.8641
R83 drain_right drain_right.n34 25.3093
R84 drain_right.n11 drain_right.n9 15.6674
R85 drain_right.n49 drain_right.n47 15.6674
R86 drain_right.n12 drain_right.n8 12.8005
R87 drain_right.n50 drain_right.n46 12.8005
R88 drain_right.n16 drain_right.n15 12.0247
R89 drain_right.n54 drain_right.n53 12.0247
R90 drain_right.n19 drain_right.n6 11.249
R91 drain_right.n57 drain_right.n44 11.249
R92 drain_right.n20 drain_right.n4 10.4732
R93 drain_right.n58 drain_right.n42 10.4732
R94 drain_right.n24 drain_right.n23 9.69747
R95 drain_right.n62 drain_right.n61 9.69747
R96 drain_right.n30 drain_right.n29 9.45567
R97 drain_right.n68 drain_right.n67 9.45567
R98 drain_right.n29 drain_right.n28 9.3005
R99 drain_right.n2 drain_right.n1 9.3005
R100 drain_right.n23 drain_right.n22 9.3005
R101 drain_right.n21 drain_right.n20 9.3005
R102 drain_right.n6 drain_right.n5 9.3005
R103 drain_right.n15 drain_right.n14 9.3005
R104 drain_right.n13 drain_right.n12 9.3005
R105 drain_right.n67 drain_right.n66 9.3005
R106 drain_right.n40 drain_right.n39 9.3005
R107 drain_right.n61 drain_right.n60 9.3005
R108 drain_right.n59 drain_right.n58 9.3005
R109 drain_right.n44 drain_right.n43 9.3005
R110 drain_right.n53 drain_right.n52 9.3005
R111 drain_right.n51 drain_right.n50 9.3005
R112 drain_right.n27 drain_right.n2 8.92171
R113 drain_right.n65 drain_right.n40 8.92171
R114 drain_right.n28 drain_right.n0 8.14595
R115 drain_right.n66 drain_right.n38 8.14595
R116 drain_right drain_right.n69 6.01097
R117 drain_right.n30 drain_right.n0 5.81868
R118 drain_right.n68 drain_right.n38 5.81868
R119 drain_right.n28 drain_right.n27 5.04292
R120 drain_right.n66 drain_right.n65 5.04292
R121 drain_right.n13 drain_right.n9 4.38594
R122 drain_right.n51 drain_right.n47 4.38594
R123 drain_right.n24 drain_right.n2 4.26717
R124 drain_right.n62 drain_right.n40 4.26717
R125 drain_right.n23 drain_right.n4 3.49141
R126 drain_right.n61 drain_right.n42 3.49141
R127 drain_right.n33 drain_right.t2 3.3005
R128 drain_right.n33 drain_right.t3 3.3005
R129 drain_right.n31 drain_right.t0 3.3005
R130 drain_right.n31 drain_right.t4 3.3005
R131 drain_right.n35 drain_right.t7 3.3005
R132 drain_right.n35 drain_right.t1 3.3005
R133 drain_right.n36 drain_right.t8 3.3005
R134 drain_right.n36 drain_right.t6 3.3005
R135 drain_right.n20 drain_right.n19 2.71565
R136 drain_right.n58 drain_right.n57 2.71565
R137 drain_right.n16 drain_right.n6 1.93989
R138 drain_right.n54 drain_right.n44 1.93989
R139 drain_right.n15 drain_right.n8 1.16414
R140 drain_right.n53 drain_right.n46 1.16414
R141 drain_right.n69 drain_right.n37 0.716017
R142 drain_right.n12 drain_right.n11 0.388379
R143 drain_right.n50 drain_right.n49 0.388379
R144 drain_right.n14 drain_right.n13 0.155672
R145 drain_right.n14 drain_right.n5 0.155672
R146 drain_right.n21 drain_right.n5 0.155672
R147 drain_right.n22 drain_right.n21 0.155672
R148 drain_right.n22 drain_right.n1 0.155672
R149 drain_right.n29 drain_right.n1 0.155672
R150 drain_right.n67 drain_right.n39 0.155672
R151 drain_right.n60 drain_right.n39 0.155672
R152 drain_right.n60 drain_right.n59 0.155672
R153 drain_right.n59 drain_right.n43 0.155672
R154 drain_right.n52 drain_right.n43 0.155672
R155 drain_right.n52 drain_right.n51 0.155672
R156 drain_right.n34 drain_right.n32 0.124033
R157 source.n138 source.n112 289.615
R158 source.n102 source.n76 289.615
R159 source.n26 source.n0 289.615
R160 source.n62 source.n36 289.615
R161 source.n123 source.n122 185
R162 source.n120 source.n119 185
R163 source.n129 source.n128 185
R164 source.n131 source.n130 185
R165 source.n116 source.n115 185
R166 source.n137 source.n136 185
R167 source.n139 source.n138 185
R168 source.n87 source.n86 185
R169 source.n84 source.n83 185
R170 source.n93 source.n92 185
R171 source.n95 source.n94 185
R172 source.n80 source.n79 185
R173 source.n101 source.n100 185
R174 source.n103 source.n102 185
R175 source.n27 source.n26 185
R176 source.n25 source.n24 185
R177 source.n4 source.n3 185
R178 source.n19 source.n18 185
R179 source.n17 source.n16 185
R180 source.n8 source.n7 185
R181 source.n11 source.n10 185
R182 source.n63 source.n62 185
R183 source.n61 source.n60 185
R184 source.n40 source.n39 185
R185 source.n55 source.n54 185
R186 source.n53 source.n52 185
R187 source.n44 source.n43 185
R188 source.n47 source.n46 185
R189 source.t6 source.n121 147.661
R190 source.t17 source.n85 147.661
R191 source.t2 source.n9 147.661
R192 source.t10 source.n45 147.661
R193 source.n122 source.n119 104.615
R194 source.n129 source.n119 104.615
R195 source.n130 source.n129 104.615
R196 source.n130 source.n115 104.615
R197 source.n137 source.n115 104.615
R198 source.n138 source.n137 104.615
R199 source.n86 source.n83 104.615
R200 source.n93 source.n83 104.615
R201 source.n94 source.n93 104.615
R202 source.n94 source.n79 104.615
R203 source.n101 source.n79 104.615
R204 source.n102 source.n101 104.615
R205 source.n26 source.n25 104.615
R206 source.n25 source.n3 104.615
R207 source.n18 source.n3 104.615
R208 source.n18 source.n17 104.615
R209 source.n17 source.n7 104.615
R210 source.n10 source.n7 104.615
R211 source.n62 source.n61 104.615
R212 source.n61 source.n39 104.615
R213 source.n54 source.n39 104.615
R214 source.n54 source.n53 104.615
R215 source.n53 source.n43 104.615
R216 source.n46 source.n43 104.615
R217 source.n122 source.t6 52.3082
R218 source.n86 source.t17 52.3082
R219 source.n10 source.t2 52.3082
R220 source.n46 source.t10 52.3082
R221 source.n33 source.n32 50.512
R222 source.n35 source.n34 50.512
R223 source.n69 source.n68 50.512
R224 source.n71 source.n70 50.512
R225 source.n111 source.n110 50.5119
R226 source.n109 source.n108 50.5119
R227 source.n75 source.n74 50.5119
R228 source.n73 source.n72 50.5119
R229 source.n143 source.n142 32.1853
R230 source.n107 source.n106 32.1853
R231 source.n31 source.n30 32.1853
R232 source.n67 source.n66 32.1853
R233 source.n73 source.n71 18.1733
R234 source.n123 source.n121 15.6674
R235 source.n87 source.n85 15.6674
R236 source.n11 source.n9 15.6674
R237 source.n47 source.n45 15.6674
R238 source.n124 source.n120 12.8005
R239 source.n88 source.n84 12.8005
R240 source.n12 source.n8 12.8005
R241 source.n48 source.n44 12.8005
R242 source.n128 source.n127 12.0247
R243 source.n92 source.n91 12.0247
R244 source.n16 source.n15 12.0247
R245 source.n52 source.n51 12.0247
R246 source.n144 source.n31 11.8371
R247 source.n131 source.n118 11.249
R248 source.n95 source.n82 11.249
R249 source.n19 source.n6 11.249
R250 source.n55 source.n42 11.249
R251 source.n132 source.n116 10.4732
R252 source.n96 source.n80 10.4732
R253 source.n20 source.n4 10.4732
R254 source.n56 source.n40 10.4732
R255 source.n136 source.n135 9.69747
R256 source.n100 source.n99 9.69747
R257 source.n24 source.n23 9.69747
R258 source.n60 source.n59 9.69747
R259 source.n142 source.n141 9.45567
R260 source.n106 source.n105 9.45567
R261 source.n30 source.n29 9.45567
R262 source.n66 source.n65 9.45567
R263 source.n141 source.n140 9.3005
R264 source.n114 source.n113 9.3005
R265 source.n135 source.n134 9.3005
R266 source.n133 source.n132 9.3005
R267 source.n118 source.n117 9.3005
R268 source.n127 source.n126 9.3005
R269 source.n125 source.n124 9.3005
R270 source.n105 source.n104 9.3005
R271 source.n78 source.n77 9.3005
R272 source.n99 source.n98 9.3005
R273 source.n97 source.n96 9.3005
R274 source.n82 source.n81 9.3005
R275 source.n91 source.n90 9.3005
R276 source.n89 source.n88 9.3005
R277 source.n29 source.n28 9.3005
R278 source.n2 source.n1 9.3005
R279 source.n23 source.n22 9.3005
R280 source.n21 source.n20 9.3005
R281 source.n6 source.n5 9.3005
R282 source.n15 source.n14 9.3005
R283 source.n13 source.n12 9.3005
R284 source.n65 source.n64 9.3005
R285 source.n38 source.n37 9.3005
R286 source.n59 source.n58 9.3005
R287 source.n57 source.n56 9.3005
R288 source.n42 source.n41 9.3005
R289 source.n51 source.n50 9.3005
R290 source.n49 source.n48 9.3005
R291 source.n139 source.n114 8.92171
R292 source.n103 source.n78 8.92171
R293 source.n27 source.n2 8.92171
R294 source.n63 source.n38 8.92171
R295 source.n140 source.n112 8.14595
R296 source.n104 source.n76 8.14595
R297 source.n28 source.n0 8.14595
R298 source.n64 source.n36 8.14595
R299 source.n142 source.n112 5.81868
R300 source.n106 source.n76 5.81868
R301 source.n30 source.n0 5.81868
R302 source.n66 source.n36 5.81868
R303 source.n144 source.n143 5.62119
R304 source.n140 source.n139 5.04292
R305 source.n104 source.n103 5.04292
R306 source.n28 source.n27 5.04292
R307 source.n64 source.n63 5.04292
R308 source.n125 source.n121 4.38594
R309 source.n89 source.n85 4.38594
R310 source.n13 source.n9 4.38594
R311 source.n49 source.n45 4.38594
R312 source.n136 source.n114 4.26717
R313 source.n100 source.n78 4.26717
R314 source.n24 source.n2 4.26717
R315 source.n60 source.n38 4.26717
R316 source.n135 source.n116 3.49141
R317 source.n99 source.n80 3.49141
R318 source.n23 source.n4 3.49141
R319 source.n59 source.n40 3.49141
R320 source.n110 source.t14 3.3005
R321 source.n110 source.t15 3.3005
R322 source.n108 source.t8 3.3005
R323 source.n108 source.t9 3.3005
R324 source.n74 source.t4 3.3005
R325 source.n74 source.t18 3.3005
R326 source.n72 source.t0 3.3005
R327 source.n72 source.t19 3.3005
R328 source.n32 source.t3 3.3005
R329 source.n32 source.t16 3.3005
R330 source.n34 source.t1 3.3005
R331 source.n34 source.t5 3.3005
R332 source.n68 source.t11 3.3005
R333 source.n68 source.t13 3.3005
R334 source.n70 source.t12 3.3005
R335 source.n70 source.t7 3.3005
R336 source.n132 source.n131 2.71565
R337 source.n96 source.n95 2.71565
R338 source.n20 source.n19 2.71565
R339 source.n56 source.n55 2.71565
R340 source.n128 source.n118 1.93989
R341 source.n92 source.n82 1.93989
R342 source.n16 source.n6 1.93989
R343 source.n52 source.n42 1.93989
R344 source.n127 source.n120 1.16414
R345 source.n91 source.n84 1.16414
R346 source.n15 source.n8 1.16414
R347 source.n51 source.n44 1.16414
R348 source.n67 source.n35 0.828086
R349 source.n109 source.n107 0.828086
R350 source.n71 source.n69 0.716017
R351 source.n69 source.n67 0.716017
R352 source.n35 source.n33 0.716017
R353 source.n33 source.n31 0.716017
R354 source.n75 source.n73 0.716017
R355 source.n107 source.n75 0.716017
R356 source.n111 source.n109 0.716017
R357 source.n143 source.n111 0.716017
R358 source.n124 source.n123 0.388379
R359 source.n88 source.n87 0.388379
R360 source.n12 source.n11 0.388379
R361 source.n48 source.n47 0.388379
R362 source source.n144 0.188
R363 source.n126 source.n125 0.155672
R364 source.n126 source.n117 0.155672
R365 source.n133 source.n117 0.155672
R366 source.n134 source.n133 0.155672
R367 source.n134 source.n113 0.155672
R368 source.n141 source.n113 0.155672
R369 source.n90 source.n89 0.155672
R370 source.n90 source.n81 0.155672
R371 source.n97 source.n81 0.155672
R372 source.n98 source.n97 0.155672
R373 source.n98 source.n77 0.155672
R374 source.n105 source.n77 0.155672
R375 source.n29 source.n1 0.155672
R376 source.n22 source.n1 0.155672
R377 source.n22 source.n21 0.155672
R378 source.n21 source.n5 0.155672
R379 source.n14 source.n5 0.155672
R380 source.n14 source.n13 0.155672
R381 source.n65 source.n37 0.155672
R382 source.n58 source.n37 0.155672
R383 source.n58 source.n57 0.155672
R384 source.n57 source.n41 0.155672
R385 source.n50 source.n41 0.155672
R386 source.n50 source.n49 0.155672
R387 plus.n2 plus.t0 388.748
R388 plus.n14 plus.t2 388.748
R389 plus.n10 plus.t7 367.767
R390 plus.n9 plus.t1 367.767
R391 plus.n1 plus.t8 367.767
R392 plus.n3 plus.t6 367.767
R393 plus.n22 plus.t5 367.767
R394 plus.n21 plus.t4 367.767
R395 plus.n13 plus.t9 367.767
R396 plus.n15 plus.t3 367.767
R397 plus.n5 plus.n4 161.3
R398 plus.n6 plus.n1 161.3
R399 plus.n8 plus.n7 161.3
R400 plus.n9 plus.n0 161.3
R401 plus.n11 plus.n10 161.3
R402 plus.n17 plus.n16 161.3
R403 plus.n18 plus.n13 161.3
R404 plus.n20 plus.n19 161.3
R405 plus.n21 plus.n12 161.3
R406 plus.n23 plus.n22 161.3
R407 plus.n5 plus.n2 70.4033
R408 plus.n17 plus.n14 70.4033
R409 plus.n10 plus.n9 48.2005
R410 plus.n22 plus.n21 48.2005
R411 plus.n8 plus.n1 36.5157
R412 plus.n4 plus.n1 36.5157
R413 plus.n20 plus.n13 36.5157
R414 plus.n16 plus.n13 36.5157
R415 plus plus.n23 27.2774
R416 plus.n3 plus.n2 20.9576
R417 plus.n15 plus.n14 20.9576
R418 plus.n9 plus.n8 11.6853
R419 plus.n4 plus.n3 11.6853
R420 plus.n21 plus.n20 11.6853
R421 plus.n16 plus.n15 11.6853
R422 plus plus.n11 9.93421
R423 plus.n6 plus.n5 0.189894
R424 plus.n7 plus.n6 0.189894
R425 plus.n7 plus.n0 0.189894
R426 plus.n11 plus.n0 0.189894
R427 plus.n23 plus.n12 0.189894
R428 plus.n19 plus.n12 0.189894
R429 plus.n19 plus.n18 0.189894
R430 plus.n18 plus.n17 0.189894
R431 drain_left.n26 drain_left.n0 289.615
R432 drain_left.n61 drain_left.n35 289.615
R433 drain_left.n11 drain_left.n10 185
R434 drain_left.n8 drain_left.n7 185
R435 drain_left.n17 drain_left.n16 185
R436 drain_left.n19 drain_left.n18 185
R437 drain_left.n4 drain_left.n3 185
R438 drain_left.n25 drain_left.n24 185
R439 drain_left.n27 drain_left.n26 185
R440 drain_left.n62 drain_left.n61 185
R441 drain_left.n60 drain_left.n59 185
R442 drain_left.n39 drain_left.n38 185
R443 drain_left.n54 drain_left.n53 185
R444 drain_left.n52 drain_left.n51 185
R445 drain_left.n43 drain_left.n42 185
R446 drain_left.n46 drain_left.n45 185
R447 drain_left.t4 drain_left.n9 147.661
R448 drain_left.t9 drain_left.n44 147.661
R449 drain_left.n10 drain_left.n7 104.615
R450 drain_left.n17 drain_left.n7 104.615
R451 drain_left.n18 drain_left.n17 104.615
R452 drain_left.n18 drain_left.n3 104.615
R453 drain_left.n25 drain_left.n3 104.615
R454 drain_left.n26 drain_left.n25 104.615
R455 drain_left.n61 drain_left.n60 104.615
R456 drain_left.n60 drain_left.n38 104.615
R457 drain_left.n53 drain_left.n38 104.615
R458 drain_left.n53 drain_left.n52 104.615
R459 drain_left.n52 drain_left.n42 104.615
R460 drain_left.n45 drain_left.n42 104.615
R461 drain_left.n34 drain_left.n33 67.672
R462 drain_left.n67 drain_left.n66 67.1908
R463 drain_left.n69 drain_left.n68 67.1907
R464 drain_left.n32 drain_left.n31 67.1907
R465 drain_left.n10 drain_left.t4 52.3082
R466 drain_left.n45 drain_left.t9 52.3082
R467 drain_left.n32 drain_left.n30 49.5797
R468 drain_left.n67 drain_left.n65 49.5797
R469 drain_left drain_left.n34 25.8626
R470 drain_left.n11 drain_left.n9 15.6674
R471 drain_left.n46 drain_left.n44 15.6674
R472 drain_left.n12 drain_left.n8 12.8005
R473 drain_left.n47 drain_left.n43 12.8005
R474 drain_left.n16 drain_left.n15 12.0247
R475 drain_left.n51 drain_left.n50 12.0247
R476 drain_left.n19 drain_left.n6 11.249
R477 drain_left.n54 drain_left.n41 11.249
R478 drain_left.n20 drain_left.n4 10.4732
R479 drain_left.n55 drain_left.n39 10.4732
R480 drain_left.n24 drain_left.n23 9.69747
R481 drain_left.n59 drain_left.n58 9.69747
R482 drain_left.n30 drain_left.n29 9.45567
R483 drain_left.n65 drain_left.n64 9.45567
R484 drain_left.n29 drain_left.n28 9.3005
R485 drain_left.n2 drain_left.n1 9.3005
R486 drain_left.n23 drain_left.n22 9.3005
R487 drain_left.n21 drain_left.n20 9.3005
R488 drain_left.n6 drain_left.n5 9.3005
R489 drain_left.n15 drain_left.n14 9.3005
R490 drain_left.n13 drain_left.n12 9.3005
R491 drain_left.n64 drain_left.n63 9.3005
R492 drain_left.n37 drain_left.n36 9.3005
R493 drain_left.n58 drain_left.n57 9.3005
R494 drain_left.n56 drain_left.n55 9.3005
R495 drain_left.n41 drain_left.n40 9.3005
R496 drain_left.n50 drain_left.n49 9.3005
R497 drain_left.n48 drain_left.n47 9.3005
R498 drain_left.n27 drain_left.n2 8.92171
R499 drain_left.n62 drain_left.n37 8.92171
R500 drain_left.n28 drain_left.n0 8.14595
R501 drain_left.n63 drain_left.n35 8.14595
R502 drain_left drain_left.n69 6.36873
R503 drain_left.n30 drain_left.n0 5.81868
R504 drain_left.n65 drain_left.n35 5.81868
R505 drain_left.n28 drain_left.n27 5.04292
R506 drain_left.n63 drain_left.n62 5.04292
R507 drain_left.n13 drain_left.n9 4.38594
R508 drain_left.n48 drain_left.n44 4.38594
R509 drain_left.n24 drain_left.n2 4.26717
R510 drain_left.n59 drain_left.n37 4.26717
R511 drain_left.n23 drain_left.n4 3.49141
R512 drain_left.n58 drain_left.n39 3.49141
R513 drain_left.n33 drain_left.t6 3.3005
R514 drain_left.n33 drain_left.t7 3.3005
R515 drain_left.n31 drain_left.t5 3.3005
R516 drain_left.n31 drain_left.t0 3.3005
R517 drain_left.n68 drain_left.t8 3.3005
R518 drain_left.n68 drain_left.t2 3.3005
R519 drain_left.n66 drain_left.t3 3.3005
R520 drain_left.n66 drain_left.t1 3.3005
R521 drain_left.n20 drain_left.n19 2.71565
R522 drain_left.n55 drain_left.n54 2.71565
R523 drain_left.n16 drain_left.n6 1.93989
R524 drain_left.n51 drain_left.n41 1.93989
R525 drain_left.n15 drain_left.n8 1.16414
R526 drain_left.n50 drain_left.n43 1.16414
R527 drain_left.n69 drain_left.n67 0.716017
R528 drain_left.n12 drain_left.n11 0.388379
R529 drain_left.n47 drain_left.n46 0.388379
R530 drain_left.n14 drain_left.n13 0.155672
R531 drain_left.n14 drain_left.n5 0.155672
R532 drain_left.n21 drain_left.n5 0.155672
R533 drain_left.n22 drain_left.n21 0.155672
R534 drain_left.n22 drain_left.n1 0.155672
R535 drain_left.n29 drain_left.n1 0.155672
R536 drain_left.n64 drain_left.n36 0.155672
R537 drain_left.n57 drain_left.n36 0.155672
R538 drain_left.n57 drain_left.n56 0.155672
R539 drain_left.n56 drain_left.n40 0.155672
R540 drain_left.n49 drain_left.n40 0.155672
R541 drain_left.n49 drain_left.n48 0.155672
R542 drain_left.n34 drain_left.n32 0.124033
C0 drain_left minus 0.171781f
C1 plus source 3.01651f
C2 drain_left drain_right 0.845043f
C3 minus plus 4.17137f
C4 plus drain_right 0.321108f
C5 minus source 3.00221f
C6 drain_right source 9.51745f
C7 minus drain_right 2.9785f
C8 drain_left plus 3.14251f
C9 drain_left source 9.521861f
C10 drain_right a_n1712_n2088# 5.10717f
C11 drain_left a_n1712_n2088# 5.3694f
C12 source a_n1712_n2088# 4.048905f
C13 minus a_n1712_n2088# 6.183603f
C14 plus a_n1712_n2088# 7.64996f
C15 drain_left.n0 a_n1712_n2088# 0.036325f
C16 drain_left.n1 a_n1712_n2088# 0.025843f
C17 drain_left.n2 a_n1712_n2088# 0.013887f
C18 drain_left.n3 a_n1712_n2088# 0.032824f
C19 drain_left.n4 a_n1712_n2088# 0.014704f
C20 drain_left.n5 a_n1712_n2088# 0.025843f
C21 drain_left.n6 a_n1712_n2088# 0.013887f
C22 drain_left.n7 a_n1712_n2088# 0.032824f
C23 drain_left.n8 a_n1712_n2088# 0.014704f
C24 drain_left.n9 a_n1712_n2088# 0.11059f
C25 drain_left.t4 a_n1712_n2088# 0.053498f
C26 drain_left.n10 a_n1712_n2088# 0.024618f
C27 drain_left.n11 a_n1712_n2088# 0.019389f
C28 drain_left.n12 a_n1712_n2088# 0.013887f
C29 drain_left.n13 a_n1712_n2088# 0.614912f
C30 drain_left.n14 a_n1712_n2088# 0.025843f
C31 drain_left.n15 a_n1712_n2088# 0.013887f
C32 drain_left.n16 a_n1712_n2088# 0.014704f
C33 drain_left.n17 a_n1712_n2088# 0.032824f
C34 drain_left.n18 a_n1712_n2088# 0.032824f
C35 drain_left.n19 a_n1712_n2088# 0.014704f
C36 drain_left.n20 a_n1712_n2088# 0.013887f
C37 drain_left.n21 a_n1712_n2088# 0.025843f
C38 drain_left.n22 a_n1712_n2088# 0.025843f
C39 drain_left.n23 a_n1712_n2088# 0.013887f
C40 drain_left.n24 a_n1712_n2088# 0.014704f
C41 drain_left.n25 a_n1712_n2088# 0.032824f
C42 drain_left.n26 a_n1712_n2088# 0.071058f
C43 drain_left.n27 a_n1712_n2088# 0.014704f
C44 drain_left.n28 a_n1712_n2088# 0.013887f
C45 drain_left.n29 a_n1712_n2088# 0.059735f
C46 drain_left.n30 a_n1712_n2088# 0.059182f
C47 drain_left.t5 a_n1712_n2088# 0.122532f
C48 drain_left.t0 a_n1712_n2088# 0.122532f
C49 drain_left.n31 a_n1712_n2088# 1.02192f
C50 drain_left.n32 a_n1712_n2088# 0.392239f
C51 drain_left.t6 a_n1712_n2088# 0.122532f
C52 drain_left.t7 a_n1712_n2088# 0.122532f
C53 drain_left.n33 a_n1712_n2088# 1.0242f
C54 drain_left.n34 a_n1712_n2088# 1.22256f
C55 drain_left.n35 a_n1712_n2088# 0.036325f
C56 drain_left.n36 a_n1712_n2088# 0.025843f
C57 drain_left.n37 a_n1712_n2088# 0.013887f
C58 drain_left.n38 a_n1712_n2088# 0.032824f
C59 drain_left.n39 a_n1712_n2088# 0.014704f
C60 drain_left.n40 a_n1712_n2088# 0.025843f
C61 drain_left.n41 a_n1712_n2088# 0.013887f
C62 drain_left.n42 a_n1712_n2088# 0.032824f
C63 drain_left.n43 a_n1712_n2088# 0.014704f
C64 drain_left.n44 a_n1712_n2088# 0.11059f
C65 drain_left.t9 a_n1712_n2088# 0.053498f
C66 drain_left.n45 a_n1712_n2088# 0.024618f
C67 drain_left.n46 a_n1712_n2088# 0.019389f
C68 drain_left.n47 a_n1712_n2088# 0.013887f
C69 drain_left.n48 a_n1712_n2088# 0.614912f
C70 drain_left.n49 a_n1712_n2088# 0.025843f
C71 drain_left.n50 a_n1712_n2088# 0.013887f
C72 drain_left.n51 a_n1712_n2088# 0.014704f
C73 drain_left.n52 a_n1712_n2088# 0.032824f
C74 drain_left.n53 a_n1712_n2088# 0.032824f
C75 drain_left.n54 a_n1712_n2088# 0.014704f
C76 drain_left.n55 a_n1712_n2088# 0.013887f
C77 drain_left.n56 a_n1712_n2088# 0.025843f
C78 drain_left.n57 a_n1712_n2088# 0.025843f
C79 drain_left.n58 a_n1712_n2088# 0.013887f
C80 drain_left.n59 a_n1712_n2088# 0.014704f
C81 drain_left.n60 a_n1712_n2088# 0.032824f
C82 drain_left.n61 a_n1712_n2088# 0.071058f
C83 drain_left.n62 a_n1712_n2088# 0.014704f
C84 drain_left.n63 a_n1712_n2088# 0.013887f
C85 drain_left.n64 a_n1712_n2088# 0.059735f
C86 drain_left.n65 a_n1712_n2088# 0.059182f
C87 drain_left.t3 a_n1712_n2088# 0.122532f
C88 drain_left.t1 a_n1712_n2088# 0.122532f
C89 drain_left.n66 a_n1712_n2088# 1.02192f
C90 drain_left.n67 a_n1712_n2088# 0.43668f
C91 drain_left.t8 a_n1712_n2088# 0.122532f
C92 drain_left.t2 a_n1712_n2088# 0.122532f
C93 drain_left.n68 a_n1712_n2088# 1.02192f
C94 drain_left.n69 a_n1712_n2088# 0.550946f
C95 plus.n0 a_n1712_n2088# 0.049316f
C96 plus.t7 a_n1712_n2088# 0.429129f
C97 plus.t1 a_n1712_n2088# 0.429129f
C98 plus.t8 a_n1712_n2088# 0.429129f
C99 plus.n1 a_n1712_n2088# 0.207314f
C100 plus.t0 a_n1712_n2088# 0.440043f
C101 plus.n2 a_n1712_n2088# 0.191592f
C102 plus.t6 a_n1712_n2088# 0.429129f
C103 plus.n3 a_n1712_n2088# 0.204578f
C104 plus.n4 a_n1712_n2088# 0.011191f
C105 plus.n5 a_n1712_n2088# 0.157316f
C106 plus.n6 a_n1712_n2088# 0.049316f
C107 plus.n7 a_n1712_n2088# 0.049316f
C108 plus.n8 a_n1712_n2088# 0.011191f
C109 plus.n9 a_n1712_n2088# 0.204578f
C110 plus.n10 a_n1712_n2088# 0.202145f
C111 plus.n11 a_n1712_n2088# 0.430202f
C112 plus.n12 a_n1712_n2088# 0.049316f
C113 plus.t5 a_n1712_n2088# 0.429129f
C114 plus.t4 a_n1712_n2088# 0.429129f
C115 plus.t9 a_n1712_n2088# 0.429129f
C116 plus.n13 a_n1712_n2088# 0.207314f
C117 plus.t2 a_n1712_n2088# 0.440043f
C118 plus.n14 a_n1712_n2088# 0.191592f
C119 plus.t3 a_n1712_n2088# 0.429129f
C120 plus.n15 a_n1712_n2088# 0.204578f
C121 plus.n16 a_n1712_n2088# 0.011191f
C122 plus.n17 a_n1712_n2088# 0.157316f
C123 plus.n18 a_n1712_n2088# 0.049316f
C124 plus.n19 a_n1712_n2088# 0.049316f
C125 plus.n20 a_n1712_n2088# 0.011191f
C126 plus.n21 a_n1712_n2088# 0.204578f
C127 plus.n22 a_n1712_n2088# 0.202145f
C128 plus.n23 a_n1712_n2088# 1.23654f
C129 source.n0 a_n1712_n2088# 0.040025f
C130 source.n1 a_n1712_n2088# 0.028476f
C131 source.n2 a_n1712_n2088# 0.015302f
C132 source.n3 a_n1712_n2088# 0.036167f
C133 source.n4 a_n1712_n2088# 0.016202f
C134 source.n5 a_n1712_n2088# 0.028476f
C135 source.n6 a_n1712_n2088# 0.015302f
C136 source.n7 a_n1712_n2088# 0.036167f
C137 source.n8 a_n1712_n2088# 0.016202f
C138 source.n9 a_n1712_n2088# 0.121856f
C139 source.t2 a_n1712_n2088# 0.058948f
C140 source.n10 a_n1712_n2088# 0.027126f
C141 source.n11 a_n1712_n2088# 0.021364f
C142 source.n12 a_n1712_n2088# 0.015302f
C143 source.n13 a_n1712_n2088# 0.677552f
C144 source.n14 a_n1712_n2088# 0.028476f
C145 source.n15 a_n1712_n2088# 0.015302f
C146 source.n16 a_n1712_n2088# 0.016202f
C147 source.n17 a_n1712_n2088# 0.036167f
C148 source.n18 a_n1712_n2088# 0.036167f
C149 source.n19 a_n1712_n2088# 0.016202f
C150 source.n20 a_n1712_n2088# 0.015302f
C151 source.n21 a_n1712_n2088# 0.028476f
C152 source.n22 a_n1712_n2088# 0.028476f
C153 source.n23 a_n1712_n2088# 0.015302f
C154 source.n24 a_n1712_n2088# 0.016202f
C155 source.n25 a_n1712_n2088# 0.036167f
C156 source.n26 a_n1712_n2088# 0.078296f
C157 source.n27 a_n1712_n2088# 0.016202f
C158 source.n28 a_n1712_n2088# 0.015302f
C159 source.n29 a_n1712_n2088# 0.06582f
C160 source.n30 a_n1712_n2088# 0.04381f
C161 source.n31 a_n1712_n2088# 0.716837f
C162 source.t3 a_n1712_n2088# 0.135014f
C163 source.t16 a_n1712_n2088# 0.135014f
C164 source.n32 a_n1712_n2088# 1.0515f
C165 source.n33 a_n1712_n2088# 0.398237f
C166 source.t1 a_n1712_n2088# 0.135014f
C167 source.t5 a_n1712_n2088# 0.135014f
C168 source.n34 a_n1712_n2088# 1.0515f
C169 source.n35 a_n1712_n2088# 0.40852f
C170 source.n36 a_n1712_n2088# 0.040025f
C171 source.n37 a_n1712_n2088# 0.028476f
C172 source.n38 a_n1712_n2088# 0.015302f
C173 source.n39 a_n1712_n2088# 0.036167f
C174 source.n40 a_n1712_n2088# 0.016202f
C175 source.n41 a_n1712_n2088# 0.028476f
C176 source.n42 a_n1712_n2088# 0.015302f
C177 source.n43 a_n1712_n2088# 0.036167f
C178 source.n44 a_n1712_n2088# 0.016202f
C179 source.n45 a_n1712_n2088# 0.121856f
C180 source.t10 a_n1712_n2088# 0.058948f
C181 source.n46 a_n1712_n2088# 0.027126f
C182 source.n47 a_n1712_n2088# 0.021364f
C183 source.n48 a_n1712_n2088# 0.015302f
C184 source.n49 a_n1712_n2088# 0.677552f
C185 source.n50 a_n1712_n2088# 0.028476f
C186 source.n51 a_n1712_n2088# 0.015302f
C187 source.n52 a_n1712_n2088# 0.016202f
C188 source.n53 a_n1712_n2088# 0.036167f
C189 source.n54 a_n1712_n2088# 0.036167f
C190 source.n55 a_n1712_n2088# 0.016202f
C191 source.n56 a_n1712_n2088# 0.015302f
C192 source.n57 a_n1712_n2088# 0.028476f
C193 source.n58 a_n1712_n2088# 0.028476f
C194 source.n59 a_n1712_n2088# 0.015302f
C195 source.n60 a_n1712_n2088# 0.016202f
C196 source.n61 a_n1712_n2088# 0.036167f
C197 source.n62 a_n1712_n2088# 0.078296f
C198 source.n63 a_n1712_n2088# 0.016202f
C199 source.n64 a_n1712_n2088# 0.015302f
C200 source.n65 a_n1712_n2088# 0.06582f
C201 source.n66 a_n1712_n2088# 0.04381f
C202 source.n67 a_n1712_n2088# 0.165908f
C203 source.t11 a_n1712_n2088# 0.135014f
C204 source.t13 a_n1712_n2088# 0.135014f
C205 source.n68 a_n1712_n2088# 1.0515f
C206 source.n69 a_n1712_n2088# 0.398237f
C207 source.t12 a_n1712_n2088# 0.135014f
C208 source.t7 a_n1712_n2088# 0.135014f
C209 source.n70 a_n1712_n2088# 1.0515f
C210 source.n71 a_n1712_n2088# 1.39624f
C211 source.t0 a_n1712_n2088# 0.135014f
C212 source.t19 a_n1712_n2088# 0.135014f
C213 source.n72 a_n1712_n2088# 1.05149f
C214 source.n73 a_n1712_n2088# 1.39625f
C215 source.t4 a_n1712_n2088# 0.135014f
C216 source.t18 a_n1712_n2088# 0.135014f
C217 source.n74 a_n1712_n2088# 1.05149f
C218 source.n75 a_n1712_n2088# 0.398245f
C219 source.n76 a_n1712_n2088# 0.040025f
C220 source.n77 a_n1712_n2088# 0.028476f
C221 source.n78 a_n1712_n2088# 0.015302f
C222 source.n79 a_n1712_n2088# 0.036167f
C223 source.n80 a_n1712_n2088# 0.016202f
C224 source.n81 a_n1712_n2088# 0.028476f
C225 source.n82 a_n1712_n2088# 0.015302f
C226 source.n83 a_n1712_n2088# 0.036167f
C227 source.n84 a_n1712_n2088# 0.016202f
C228 source.n85 a_n1712_n2088# 0.121856f
C229 source.t17 a_n1712_n2088# 0.058948f
C230 source.n86 a_n1712_n2088# 0.027126f
C231 source.n87 a_n1712_n2088# 0.021364f
C232 source.n88 a_n1712_n2088# 0.015302f
C233 source.n89 a_n1712_n2088# 0.677552f
C234 source.n90 a_n1712_n2088# 0.028476f
C235 source.n91 a_n1712_n2088# 0.015302f
C236 source.n92 a_n1712_n2088# 0.016202f
C237 source.n93 a_n1712_n2088# 0.036167f
C238 source.n94 a_n1712_n2088# 0.036167f
C239 source.n95 a_n1712_n2088# 0.016202f
C240 source.n96 a_n1712_n2088# 0.015302f
C241 source.n97 a_n1712_n2088# 0.028476f
C242 source.n98 a_n1712_n2088# 0.028476f
C243 source.n99 a_n1712_n2088# 0.015302f
C244 source.n100 a_n1712_n2088# 0.016202f
C245 source.n101 a_n1712_n2088# 0.036167f
C246 source.n102 a_n1712_n2088# 0.078296f
C247 source.n103 a_n1712_n2088# 0.016202f
C248 source.n104 a_n1712_n2088# 0.015302f
C249 source.n105 a_n1712_n2088# 0.06582f
C250 source.n106 a_n1712_n2088# 0.04381f
C251 source.n107 a_n1712_n2088# 0.165908f
C252 source.t8 a_n1712_n2088# 0.135014f
C253 source.t9 a_n1712_n2088# 0.135014f
C254 source.n108 a_n1712_n2088# 1.05149f
C255 source.n109 a_n1712_n2088# 0.408527f
C256 source.t14 a_n1712_n2088# 0.135014f
C257 source.t15 a_n1712_n2088# 0.135014f
C258 source.n110 a_n1712_n2088# 1.05149f
C259 source.n111 a_n1712_n2088# 0.398245f
C260 source.n112 a_n1712_n2088# 0.040025f
C261 source.n113 a_n1712_n2088# 0.028476f
C262 source.n114 a_n1712_n2088# 0.015302f
C263 source.n115 a_n1712_n2088# 0.036167f
C264 source.n116 a_n1712_n2088# 0.016202f
C265 source.n117 a_n1712_n2088# 0.028476f
C266 source.n118 a_n1712_n2088# 0.015302f
C267 source.n119 a_n1712_n2088# 0.036167f
C268 source.n120 a_n1712_n2088# 0.016202f
C269 source.n121 a_n1712_n2088# 0.121856f
C270 source.t6 a_n1712_n2088# 0.058948f
C271 source.n122 a_n1712_n2088# 0.027126f
C272 source.n123 a_n1712_n2088# 0.021364f
C273 source.n124 a_n1712_n2088# 0.015302f
C274 source.n125 a_n1712_n2088# 0.677552f
C275 source.n126 a_n1712_n2088# 0.028476f
C276 source.n127 a_n1712_n2088# 0.015302f
C277 source.n128 a_n1712_n2088# 0.016202f
C278 source.n129 a_n1712_n2088# 0.036167f
C279 source.n130 a_n1712_n2088# 0.036167f
C280 source.n131 a_n1712_n2088# 0.016202f
C281 source.n132 a_n1712_n2088# 0.015302f
C282 source.n133 a_n1712_n2088# 0.028476f
C283 source.n134 a_n1712_n2088# 0.028476f
C284 source.n135 a_n1712_n2088# 0.015302f
C285 source.n136 a_n1712_n2088# 0.016202f
C286 source.n137 a_n1712_n2088# 0.036167f
C287 source.n138 a_n1712_n2088# 0.078296f
C288 source.n139 a_n1712_n2088# 0.016202f
C289 source.n140 a_n1712_n2088# 0.015302f
C290 source.n141 a_n1712_n2088# 0.06582f
C291 source.n142 a_n1712_n2088# 0.04381f
C292 source.n143 a_n1712_n2088# 0.306399f
C293 source.n144 a_n1712_n2088# 1.17296f
C294 drain_right.n0 a_n1712_n2088# 0.036328f
C295 drain_right.n1 a_n1712_n2088# 0.025845f
C296 drain_right.n2 a_n1712_n2088# 0.013888f
C297 drain_right.n3 a_n1712_n2088# 0.032827f
C298 drain_right.n4 a_n1712_n2088# 0.014705f
C299 drain_right.n5 a_n1712_n2088# 0.025845f
C300 drain_right.n6 a_n1712_n2088# 0.013888f
C301 drain_right.n7 a_n1712_n2088# 0.032827f
C302 drain_right.n8 a_n1712_n2088# 0.014705f
C303 drain_right.n9 a_n1712_n2088# 0.1106f
C304 drain_right.t5 a_n1712_n2088# 0.053503f
C305 drain_right.n10 a_n1712_n2088# 0.02462f
C306 drain_right.n11 a_n1712_n2088# 0.01939f
C307 drain_right.n12 a_n1712_n2088# 0.013888f
C308 drain_right.n13 a_n1712_n2088# 0.614966f
C309 drain_right.n14 a_n1712_n2088# 0.025845f
C310 drain_right.n15 a_n1712_n2088# 0.013888f
C311 drain_right.n16 a_n1712_n2088# 0.014705f
C312 drain_right.n17 a_n1712_n2088# 0.032827f
C313 drain_right.n18 a_n1712_n2088# 0.032827f
C314 drain_right.n19 a_n1712_n2088# 0.014705f
C315 drain_right.n20 a_n1712_n2088# 0.013888f
C316 drain_right.n21 a_n1712_n2088# 0.025845f
C317 drain_right.n22 a_n1712_n2088# 0.025845f
C318 drain_right.n23 a_n1712_n2088# 0.013888f
C319 drain_right.n24 a_n1712_n2088# 0.014705f
C320 drain_right.n25 a_n1712_n2088# 0.032827f
C321 drain_right.n26 a_n1712_n2088# 0.071064f
C322 drain_right.n27 a_n1712_n2088# 0.014705f
C323 drain_right.n28 a_n1712_n2088# 0.013888f
C324 drain_right.n29 a_n1712_n2088# 0.05974f
C325 drain_right.n30 a_n1712_n2088# 0.059187f
C326 drain_right.t0 a_n1712_n2088# 0.122543f
C327 drain_right.t4 a_n1712_n2088# 0.122543f
C328 drain_right.n31 a_n1712_n2088# 1.02201f
C329 drain_right.n32 a_n1712_n2088# 0.392273f
C330 drain_right.t2 a_n1712_n2088# 0.122543f
C331 drain_right.t3 a_n1712_n2088# 0.122543f
C332 drain_right.n33 a_n1712_n2088# 1.02429f
C333 drain_right.n34 a_n1712_n2088# 1.17008f
C334 drain_right.t7 a_n1712_n2088# 0.122543f
C335 drain_right.t1 a_n1712_n2088# 0.122543f
C336 drain_right.n35 a_n1712_n2088# 1.02558f
C337 drain_right.t8 a_n1712_n2088# 0.122543f
C338 drain_right.t6 a_n1712_n2088# 0.122543f
C339 drain_right.n36 a_n1712_n2088# 1.02201f
C340 drain_right.n37 a_n1712_n2088# 0.664722f
C341 drain_right.n38 a_n1712_n2088# 0.036328f
C342 drain_right.n39 a_n1712_n2088# 0.025845f
C343 drain_right.n40 a_n1712_n2088# 0.013888f
C344 drain_right.n41 a_n1712_n2088# 0.032827f
C345 drain_right.n42 a_n1712_n2088# 0.014705f
C346 drain_right.n43 a_n1712_n2088# 0.025845f
C347 drain_right.n44 a_n1712_n2088# 0.013888f
C348 drain_right.n45 a_n1712_n2088# 0.032827f
C349 drain_right.n46 a_n1712_n2088# 0.014705f
C350 drain_right.n47 a_n1712_n2088# 0.1106f
C351 drain_right.t9 a_n1712_n2088# 0.053503f
C352 drain_right.n48 a_n1712_n2088# 0.02462f
C353 drain_right.n49 a_n1712_n2088# 0.01939f
C354 drain_right.n50 a_n1712_n2088# 0.013888f
C355 drain_right.n51 a_n1712_n2088# 0.614966f
C356 drain_right.n52 a_n1712_n2088# 0.025845f
C357 drain_right.n53 a_n1712_n2088# 0.013888f
C358 drain_right.n54 a_n1712_n2088# 0.014705f
C359 drain_right.n55 a_n1712_n2088# 0.032827f
C360 drain_right.n56 a_n1712_n2088# 0.032827f
C361 drain_right.n57 a_n1712_n2088# 0.014705f
C362 drain_right.n58 a_n1712_n2088# 0.013888f
C363 drain_right.n59 a_n1712_n2088# 0.025845f
C364 drain_right.n60 a_n1712_n2088# 0.025845f
C365 drain_right.n61 a_n1712_n2088# 0.013888f
C366 drain_right.n62 a_n1712_n2088# 0.014705f
C367 drain_right.n63 a_n1712_n2088# 0.032827f
C368 drain_right.n64 a_n1712_n2088# 0.071064f
C369 drain_right.n65 a_n1712_n2088# 0.014705f
C370 drain_right.n66 a_n1712_n2088# 0.013888f
C371 drain_right.n67 a_n1712_n2088# 0.05974f
C372 drain_right.n68 a_n1712_n2088# 0.057609f
C373 drain_right.n69 a_n1712_n2088# 0.335983f
C374 minus.n0 a_n1712_n2088# 0.048369f
C375 minus.t4 a_n1712_n2088# 0.420888f
C376 minus.n1 a_n1712_n2088# 0.203333f
C377 minus.t5 a_n1712_n2088# 0.431592f
C378 minus.n2 a_n1712_n2088# 0.187912f
C379 minus.t2 a_n1712_n2088# 0.420888f
C380 minus.n3 a_n1712_n2088# 0.200649f
C381 minus.n4 a_n1712_n2088# 0.010976f
C382 minus.n5 a_n1712_n2088# 0.154295f
C383 minus.n6 a_n1712_n2088# 0.048369f
C384 minus.n7 a_n1712_n2088# 0.048369f
C385 minus.n8 a_n1712_n2088# 0.010976f
C386 minus.t8 a_n1712_n2088# 0.420888f
C387 minus.n9 a_n1712_n2088# 0.200649f
C388 minus.t3 a_n1712_n2088# 0.420888f
C389 minus.n10 a_n1712_n2088# 0.198263f
C390 minus.n11 a_n1712_n2088# 1.34177f
C391 minus.n12 a_n1712_n2088# 0.048369f
C392 minus.t1 a_n1712_n2088# 0.420888f
C393 minus.n13 a_n1712_n2088# 0.203333f
C394 minus.t7 a_n1712_n2088# 0.431592f
C395 minus.n14 a_n1712_n2088# 0.187912f
C396 minus.t6 a_n1712_n2088# 0.420888f
C397 minus.n15 a_n1712_n2088# 0.200649f
C398 minus.n16 a_n1712_n2088# 0.010976f
C399 minus.n17 a_n1712_n2088# 0.154295f
C400 minus.n18 a_n1712_n2088# 0.048369f
C401 minus.n19 a_n1712_n2088# 0.048369f
C402 minus.n20 a_n1712_n2088# 0.010976f
C403 minus.t0 a_n1712_n2088# 0.420888f
C404 minus.n21 a_n1712_n2088# 0.200649f
C405 minus.t9 a_n1712_n2088# 0.420888f
C406 minus.n22 a_n1712_n2088# 0.198263f
C407 minus.n23 a_n1712_n2088# 0.323379f
C408 minus.n24 a_n1712_n2088# 1.64849f
.ends

