* NGSPICE file created from diffpair77.ext - technology: sky130A

.subckt diffpair77 minus drain_right drain_left source plus
X0 a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 source.t30 minus.t0 drain_right.t11 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X3 source.t29 minus.t1 drain_right.t7 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X4 drain_left.t15 plus.t0 source.t6 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X5 drain_left.t14 plus.t1 source.t4 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X6 source.t28 minus.t2 drain_right.t6 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X7 source.t27 minus.t3 drain_right.t12 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_right.t8 minus.t4 source.t26 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X9 drain_left.t13 plus.t2 source.t3 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X10 drain_left.t12 plus.t3 source.t5 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X11 source.t25 minus.t5 drain_right.t2 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X12 drain_right.t15 minus.t6 source.t24 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X13 drain_right.t0 minus.t7 source.t23 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X14 source.t22 minus.t8 drain_right.t13 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X15 drain_left.t11 plus.t4 source.t2 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X16 source.t21 minus.t9 drain_right.t9 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X17 source.t1 plus.t5 drain_left.t10 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_right.t5 minus.t10 source.t20 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X19 source.t0 plus.t6 drain_left.t9 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X20 drain_left.t8 plus.t7 source.t10 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 drain_left.t7 plus.t8 source.t31 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 source.t19 minus.t11 drain_right.t3 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X23 drain_right.t1 minus.t12 source.t18 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X24 drain_right.t4 minus.t13 source.t17 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X25 source.t13 plus.t9 drain_left.t6 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X26 a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X27 a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X28 source.t9 plus.t10 drain_left.t5 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X29 drain_left.t4 plus.t11 source.t8 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X30 drain_right.t14 minus.t14 source.t16 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X31 drain_right.t10 minus.t15 source.t15 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X32 source.t7 plus.t12 drain_left.t3 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X33 source.t14 plus.t13 drain_left.t2 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X34 source.t12 plus.t14 drain_left.t1 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X35 source.t11 plus.t15 drain_left.t0 a_n2750_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n21 minus.n20 161.3
R1 minus.n19 minus.n0 161.3
R2 minus.n15 minus.n14 161.3
R3 minus.n13 minus.n2 161.3
R4 minus.n12 minus.n11 161.3
R5 minus.n10 minus.n3 161.3
R6 minus.n9 minus.n8 161.3
R7 minus.n43 minus.n42 161.3
R8 minus.n41 minus.n22 161.3
R9 minus.n37 minus.n36 161.3
R10 minus.n35 minus.n24 161.3
R11 minus.n34 minus.n33 161.3
R12 minus.n32 minus.n25 161.3
R13 minus.n31 minus.n30 161.3
R14 minus.n5 minus.t7 100.252
R15 minus.n27 minus.t3 100.252
R16 minus.n18 minus.n17 80.6037
R17 minus.n16 minus.n1 80.6037
R18 minus.n7 minus.n4 80.6037
R19 minus.n40 minus.n39 80.6037
R20 minus.n38 minus.n23 80.6037
R21 minus.n29 minus.n26 80.6037
R22 minus.n6 minus.t5 79.2293
R23 minus.n7 minus.t4 79.2293
R24 minus.n3 minus.t9 79.2293
R25 minus.n13 minus.t10 79.2293
R26 minus.n1 minus.t8 79.2293
R27 minus.n18 minus.t6 79.2293
R28 minus.n20 minus.t11 79.2293
R29 minus.n28 minus.t13 79.2293
R30 minus.n29 minus.t2 79.2293
R31 minus.n25 minus.t12 79.2293
R32 minus.n35 minus.t1 79.2293
R33 minus.n23 minus.t14 79.2293
R34 minus.n40 minus.t0 79.2293
R35 minus.n42 minus.t15 79.2293
R36 minus.n7 minus.n6 48.2005
R37 minus.n18 minus.n1 48.2005
R38 minus.n29 minus.n28 48.2005
R39 minus.n40 minus.n23 48.2005
R40 minus.n8 minus.n7 43.0884
R41 minus.n14 minus.n1 43.0884
R42 minus.n30 minus.n29 43.0884
R43 minus.n36 minus.n23 43.0884
R44 minus.n19 minus.n18 40.1672
R45 minus.n41 minus.n40 40.1672
R46 minus.n5 minus.n4 31.6481
R47 minus.n27 minus.n26 31.6481
R48 minus.n44 minus.n21 31.3603
R49 minus.n13 minus.n12 24.1005
R50 minus.n12 minus.n3 24.1005
R51 minus.n34 minus.n25 24.1005
R52 minus.n35 minus.n34 24.1005
R53 minus.n6 minus.n5 17.444
R54 minus.n28 minus.n27 17.444
R55 minus.n20 minus.n19 8.03383
R56 minus.n42 minus.n41 8.03383
R57 minus.n44 minus.n43 6.6558
R58 minus.n8 minus.n3 5.11262
R59 minus.n14 minus.n13 5.11262
R60 minus.n30 minus.n25 5.11262
R61 minus.n36 minus.n35 5.11262
R62 minus.n17 minus.n16 0.380177
R63 minus.n39 minus.n38 0.380177
R64 minus.n17 minus.n0 0.285035
R65 minus.n16 minus.n15 0.285035
R66 minus.n9 minus.n4 0.285035
R67 minus.n31 minus.n26 0.285035
R68 minus.n38 minus.n37 0.285035
R69 minus.n39 minus.n22 0.285035
R70 minus.n21 minus.n0 0.189894
R71 minus.n15 minus.n2 0.189894
R72 minus.n11 minus.n2 0.189894
R73 minus.n11 minus.n10 0.189894
R74 minus.n10 minus.n9 0.189894
R75 minus.n32 minus.n31 0.189894
R76 minus.n33 minus.n32 0.189894
R77 minus.n33 minus.n24 0.189894
R78 minus.n37 minus.n24 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 drain_right.n9 drain_right.n7 241.107
R82 drain_right.n5 drain_right.n3 241.106
R83 drain_right.n2 drain_right.n0 241.106
R84 drain_right.n9 drain_right.n8 240.132
R85 drain_right.n11 drain_right.n10 240.132
R86 drain_right.n13 drain_right.n12 240.132
R87 drain_right.n5 drain_right.n4 240.131
R88 drain_right.n2 drain_right.n1 240.131
R89 drain_right drain_right.n6 24.8124
R90 drain_right.n3 drain_right.t11 19.8005
R91 drain_right.n3 drain_right.t10 19.8005
R92 drain_right.n4 drain_right.t7 19.8005
R93 drain_right.n4 drain_right.t14 19.8005
R94 drain_right.n1 drain_right.t6 19.8005
R95 drain_right.n1 drain_right.t1 19.8005
R96 drain_right.n0 drain_right.t12 19.8005
R97 drain_right.n0 drain_right.t4 19.8005
R98 drain_right.n7 drain_right.t2 19.8005
R99 drain_right.n7 drain_right.t0 19.8005
R100 drain_right.n8 drain_right.t9 19.8005
R101 drain_right.n8 drain_right.t8 19.8005
R102 drain_right.n10 drain_right.t13 19.8005
R103 drain_right.n10 drain_right.t5 19.8005
R104 drain_right.n12 drain_right.t3 19.8005
R105 drain_right.n12 drain_right.t15 19.8005
R106 drain_right drain_right.n13 6.62735
R107 drain_right.n13 drain_right.n11 0.974638
R108 drain_right.n11 drain_right.n9 0.974638
R109 drain_right.n6 drain_right.n5 0.432223
R110 drain_right.n6 drain_right.n2 0.432223
R111 source.n0 source.t2 243.255
R112 source.n7 source.t14 243.255
R113 source.n8 source.t23 243.255
R114 source.n15 source.t19 243.255
R115 source.n31 source.t15 243.254
R116 source.n24 source.t27 243.254
R117 source.n23 source.t3 243.254
R118 source.n16 source.t1 243.254
R119 source.n2 source.n1 223.454
R120 source.n4 source.n3 223.454
R121 source.n6 source.n5 223.454
R122 source.n10 source.n9 223.454
R123 source.n12 source.n11 223.454
R124 source.n14 source.n13 223.454
R125 source.n30 source.n29 223.453
R126 source.n28 source.n27 223.453
R127 source.n26 source.n25 223.453
R128 source.n22 source.n21 223.453
R129 source.n20 source.n19 223.453
R130 source.n18 source.n17 223.453
R131 source.n29 source.t16 19.8005
R132 source.n29 source.t30 19.8005
R133 source.n27 source.t18 19.8005
R134 source.n27 source.t29 19.8005
R135 source.n25 source.t17 19.8005
R136 source.n25 source.t28 19.8005
R137 source.n21 source.t5 19.8005
R138 source.n21 source.t7 19.8005
R139 source.n19 source.t6 19.8005
R140 source.n19 source.t12 19.8005
R141 source.n17 source.t4 19.8005
R142 source.n17 source.t11 19.8005
R143 source.n1 source.t10 19.8005
R144 source.n1 source.t0 19.8005
R145 source.n3 source.t31 19.8005
R146 source.n3 source.t9 19.8005
R147 source.n5 source.t8 19.8005
R148 source.n5 source.t13 19.8005
R149 source.n9 source.t26 19.8005
R150 source.n9 source.t25 19.8005
R151 source.n11 source.t20 19.8005
R152 source.n11 source.t21 19.8005
R153 source.n13 source.t24 19.8005
R154 source.n13 source.t22 19.8005
R155 source.n16 source.n15 13.9285
R156 source.n32 source.n0 8.17853
R157 source.n32 source.n31 5.7505
R158 source.n15 source.n14 0.974638
R159 source.n14 source.n12 0.974638
R160 source.n12 source.n10 0.974638
R161 source.n10 source.n8 0.974638
R162 source.n7 source.n6 0.974638
R163 source.n6 source.n4 0.974638
R164 source.n4 source.n2 0.974638
R165 source.n2 source.n0 0.974638
R166 source.n18 source.n16 0.974638
R167 source.n20 source.n18 0.974638
R168 source.n22 source.n20 0.974638
R169 source.n23 source.n22 0.974638
R170 source.n26 source.n24 0.974638
R171 source.n28 source.n26 0.974638
R172 source.n30 source.n28 0.974638
R173 source.n31 source.n30 0.974638
R174 source.n8 source.n7 0.470328
R175 source.n24 source.n23 0.470328
R176 source source.n32 0.188
R177 plus.n10 plus.n9 161.3
R178 plus.n11 plus.n4 161.3
R179 plus.n13 plus.n12 161.3
R180 plus.n14 plus.n3 161.3
R181 plus.n16 plus.n15 161.3
R182 plus.n19 plus.n0 161.3
R183 plus.n21 plus.n20 161.3
R184 plus.n32 plus.n31 161.3
R185 plus.n33 plus.n26 161.3
R186 plus.n35 plus.n34 161.3
R187 plus.n36 plus.n25 161.3
R188 plus.n38 plus.n37 161.3
R189 plus.n41 plus.n22 161.3
R190 plus.n43 plus.n42 161.3
R191 plus.n7 plus.t13 100.252
R192 plus.n29 plus.t2 100.252
R193 plus.n8 plus.n5 80.6037
R194 plus.n17 plus.n2 80.6037
R195 plus.n18 plus.n1 80.6037
R196 plus.n30 plus.n27 80.6037
R197 plus.n39 plus.n24 80.6037
R198 plus.n40 plus.n23 80.6037
R199 plus.n20 plus.t4 79.2293
R200 plus.n18 plus.t6 79.2293
R201 plus.n17 plus.t7 79.2293
R202 plus.n3 plus.t10 79.2293
R203 plus.n11 plus.t8 79.2293
R204 plus.n5 plus.t9 79.2293
R205 plus.n6 plus.t11 79.2293
R206 plus.n42 plus.t5 79.2293
R207 plus.n40 plus.t1 79.2293
R208 plus.n39 plus.t15 79.2293
R209 plus.n25 plus.t0 79.2293
R210 plus.n33 plus.t14 79.2293
R211 plus.n27 plus.t3 79.2293
R212 plus.n28 plus.t12 79.2293
R213 plus.n18 plus.n17 48.2005
R214 plus.n6 plus.n5 48.2005
R215 plus.n40 plus.n39 48.2005
R216 plus.n28 plus.n27 48.2005
R217 plus.n17 plus.n16 43.0884
R218 plus.n10 plus.n5 43.0884
R219 plus.n39 plus.n38 43.0884
R220 plus.n32 plus.n27 43.0884
R221 plus.n19 plus.n18 40.1672
R222 plus.n41 plus.n40 40.1672
R223 plus.n8 plus.n7 31.6481
R224 plus.n30 plus.n29 31.6481
R225 plus plus.n43 29.4081
R226 plus.n12 plus.n11 24.1005
R227 plus.n12 plus.n3 24.1005
R228 plus.n34 plus.n25 24.1005
R229 plus.n34 plus.n33 24.1005
R230 plus.n7 plus.n6 17.444
R231 plus.n29 plus.n28 17.444
R232 plus plus.n21 8.13308
R233 plus.n20 plus.n19 8.03383
R234 plus.n42 plus.n41 8.03383
R235 plus.n16 plus.n3 5.11262
R236 plus.n11 plus.n10 5.11262
R237 plus.n38 plus.n25 5.11262
R238 plus.n33 plus.n32 5.11262
R239 plus.n2 plus.n1 0.380177
R240 plus.n24 plus.n23 0.380177
R241 plus.n9 plus.n8 0.285035
R242 plus.n15 plus.n2 0.285035
R243 plus.n1 plus.n0 0.285035
R244 plus.n23 plus.n22 0.285035
R245 plus.n37 plus.n24 0.285035
R246 plus.n31 plus.n30 0.285035
R247 plus.n9 plus.n4 0.189894
R248 plus.n13 plus.n4 0.189894
R249 plus.n14 plus.n13 0.189894
R250 plus.n15 plus.n14 0.189894
R251 plus.n21 plus.n0 0.189894
R252 plus.n43 plus.n22 0.189894
R253 plus.n37 plus.n36 0.189894
R254 plus.n36 plus.n35 0.189894
R255 plus.n35 plus.n26 0.189894
R256 plus.n31 plus.n26 0.189894
R257 drain_left.n9 drain_left.n7 241.107
R258 drain_left.n5 drain_left.n3 241.106
R259 drain_left.n2 drain_left.n0 241.106
R260 drain_left.n13 drain_left.n12 240.132
R261 drain_left.n11 drain_left.n10 240.132
R262 drain_left.n9 drain_left.n8 240.132
R263 drain_left.n5 drain_left.n4 240.131
R264 drain_left.n2 drain_left.n1 240.131
R265 drain_left drain_left.n6 25.3656
R266 drain_left.n3 drain_left.t3 19.8005
R267 drain_left.n3 drain_left.t13 19.8005
R268 drain_left.n4 drain_left.t1 19.8005
R269 drain_left.n4 drain_left.t12 19.8005
R270 drain_left.n1 drain_left.t0 19.8005
R271 drain_left.n1 drain_left.t15 19.8005
R272 drain_left.n0 drain_left.t10 19.8005
R273 drain_left.n0 drain_left.t14 19.8005
R274 drain_left.n12 drain_left.t9 19.8005
R275 drain_left.n12 drain_left.t11 19.8005
R276 drain_left.n10 drain_left.t5 19.8005
R277 drain_left.n10 drain_left.t8 19.8005
R278 drain_left.n8 drain_left.t6 19.8005
R279 drain_left.n8 drain_left.t7 19.8005
R280 drain_left.n7 drain_left.t2 19.8005
R281 drain_left.n7 drain_left.t4 19.8005
R282 drain_left drain_left.n13 6.62735
R283 drain_left.n11 drain_left.n9 0.974638
R284 drain_left.n13 drain_left.n11 0.974638
R285 drain_left.n6 drain_left.n5 0.432223
R286 drain_left.n6 drain_left.n2 0.432223
C0 drain_right minus 1.46604f
C1 plus drain_left 1.73916f
C2 plus source 2.25497f
C3 drain_right drain_left 1.4495f
C4 drain_right source 4.88389f
C5 minus drain_left 0.18074f
C6 minus source 2.24111f
C7 source drain_left 4.88114f
C8 drain_right plus 0.43915f
C9 minus plus 4.54859f
C10 drain_right a_n2750_n1088# 4.43945f
C11 drain_left a_n2750_n1088# 4.78121f
C12 source a_n2750_n1088# 2.819126f
C13 minus a_n2750_n1088# 10.092447f
C14 plus a_n2750_n1088# 11.08146f
C15 drain_left.t10 a_n2750_n1088# 0.015578f
C16 drain_left.t14 a_n2750_n1088# 0.015578f
C17 drain_left.n0 a_n2750_n1088# 0.061622f
C18 drain_left.t0 a_n2750_n1088# 0.015578f
C19 drain_left.t15 a_n2750_n1088# 0.015578f
C20 drain_left.n1 a_n2750_n1088# 0.060533f
C21 drain_left.n2 a_n2750_n1088# 0.496688f
C22 drain_left.t3 a_n2750_n1088# 0.015578f
C23 drain_left.t13 a_n2750_n1088# 0.015578f
C24 drain_left.n3 a_n2750_n1088# 0.061622f
C25 drain_left.t1 a_n2750_n1088# 0.015578f
C26 drain_left.t12 a_n2750_n1088# 0.015578f
C27 drain_left.n4 a_n2750_n1088# 0.060533f
C28 drain_left.n5 a_n2750_n1088# 0.496688f
C29 drain_left.n6 a_n2750_n1088# 0.727554f
C30 drain_left.t2 a_n2750_n1088# 0.015578f
C31 drain_left.t4 a_n2750_n1088# 0.015578f
C32 drain_left.n7 a_n2750_n1088# 0.061622f
C33 drain_left.t6 a_n2750_n1088# 0.015578f
C34 drain_left.t7 a_n2750_n1088# 0.015578f
C35 drain_left.n8 a_n2750_n1088# 0.060533f
C36 drain_left.n9 a_n2750_n1088# 0.530084f
C37 drain_left.t5 a_n2750_n1088# 0.015578f
C38 drain_left.t8 a_n2750_n1088# 0.015578f
C39 drain_left.n10 a_n2750_n1088# 0.060533f
C40 drain_left.n11 a_n2750_n1088# 0.261617f
C41 drain_left.t9 a_n2750_n1088# 0.015578f
C42 drain_left.t11 a_n2750_n1088# 0.015578f
C43 drain_left.n12 a_n2750_n1088# 0.060533f
C44 drain_left.n13 a_n2750_n1088# 0.438387f
C45 plus.n0 a_n2750_n1088# 0.047829f
C46 plus.t4 a_n2750_n1088# 0.097236f
C47 plus.t6 a_n2750_n1088# 0.097236f
C48 plus.n1 a_n2750_n1088# 0.059702f
C49 plus.t7 a_n2750_n1088# 0.097236f
C50 plus.n2 a_n2750_n1088# 0.059702f
C51 plus.t10 a_n2750_n1088# 0.097236f
C52 plus.n3 a_n2750_n1088# 0.09339f
C53 plus.n4 a_n2750_n1088# 0.035844f
C54 plus.t8 a_n2750_n1088# 0.097236f
C55 plus.t9 a_n2750_n1088# 0.097236f
C56 plus.n5 a_n2750_n1088# 0.103623f
C57 plus.t11 a_n2750_n1088# 0.097236f
C58 plus.n6 a_n2750_n1088# 0.103904f
C59 plus.t13 a_n2750_n1088# 0.117477f
C60 plus.n7 a_n2750_n1088# 0.079492f
C61 plus.n8 a_n2750_n1088# 0.205581f
C62 plus.n9 a_n2750_n1088# 0.047829f
C63 plus.n10 a_n2750_n1088# 0.008134f
C64 plus.n11 a_n2750_n1088# 0.09339f
C65 plus.n12 a_n2750_n1088# 0.008134f
C66 plus.n13 a_n2750_n1088# 0.035844f
C67 plus.n14 a_n2750_n1088# 0.035844f
C68 plus.n15 a_n2750_n1088# 0.047829f
C69 plus.n16 a_n2750_n1088# 0.008134f
C70 plus.n17 a_n2750_n1088# 0.103623f
C71 plus.n18 a_n2750_n1088# 0.103181f
C72 plus.n19 a_n2750_n1088# 0.008134f
C73 plus.n20 a_n2750_n1088# 0.090185f
C74 plus.n21 a_n2750_n1088# 0.259517f
C75 plus.n22 a_n2750_n1088# 0.047829f
C76 plus.t5 a_n2750_n1088# 0.097236f
C77 plus.n23 a_n2750_n1088# 0.059702f
C78 plus.t1 a_n2750_n1088# 0.097236f
C79 plus.n24 a_n2750_n1088# 0.059702f
C80 plus.t15 a_n2750_n1088# 0.097236f
C81 plus.t0 a_n2750_n1088# 0.097236f
C82 plus.n25 a_n2750_n1088# 0.09339f
C83 plus.n26 a_n2750_n1088# 0.035844f
C84 plus.t14 a_n2750_n1088# 0.097236f
C85 plus.t3 a_n2750_n1088# 0.097236f
C86 plus.n27 a_n2750_n1088# 0.103623f
C87 plus.t12 a_n2750_n1088# 0.097236f
C88 plus.n28 a_n2750_n1088# 0.103904f
C89 plus.t2 a_n2750_n1088# 0.117477f
C90 plus.n29 a_n2750_n1088# 0.079492f
C91 plus.n30 a_n2750_n1088# 0.205581f
C92 plus.n31 a_n2750_n1088# 0.047829f
C93 plus.n32 a_n2750_n1088# 0.008134f
C94 plus.n33 a_n2750_n1088# 0.09339f
C95 plus.n34 a_n2750_n1088# 0.008134f
C96 plus.n35 a_n2750_n1088# 0.035844f
C97 plus.n36 a_n2750_n1088# 0.035844f
C98 plus.n37 a_n2750_n1088# 0.047829f
C99 plus.n38 a_n2750_n1088# 0.008134f
C100 plus.n39 a_n2750_n1088# 0.103623f
C101 plus.n40 a_n2750_n1088# 0.103181f
C102 plus.n41 a_n2750_n1088# 0.008134f
C103 plus.n42 a_n2750_n1088# 0.090185f
C104 plus.n43 a_n2750_n1088# 0.973472f
C105 source.t2 a_n2750_n1088# 0.157438f
C106 source.n0 a_n2750_n1088# 0.764719f
C107 source.t10 a_n2750_n1088# 0.028286f
C108 source.t0 a_n2750_n1088# 0.028286f
C109 source.n1 a_n2750_n1088# 0.091737f
C110 source.n2 a_n2750_n1088# 0.444555f
C111 source.t31 a_n2750_n1088# 0.028286f
C112 source.t9 a_n2750_n1088# 0.028286f
C113 source.n3 a_n2750_n1088# 0.091737f
C114 source.n4 a_n2750_n1088# 0.444555f
C115 source.t8 a_n2750_n1088# 0.028286f
C116 source.t13 a_n2750_n1088# 0.028286f
C117 source.n5 a_n2750_n1088# 0.091737f
C118 source.n6 a_n2750_n1088# 0.444555f
C119 source.t14 a_n2750_n1088# 0.157438f
C120 source.n7 a_n2750_n1088# 0.397832f
C121 source.t23 a_n2750_n1088# 0.157438f
C122 source.n8 a_n2750_n1088# 0.397832f
C123 source.t26 a_n2750_n1088# 0.028286f
C124 source.t25 a_n2750_n1088# 0.028286f
C125 source.n9 a_n2750_n1088# 0.091737f
C126 source.n10 a_n2750_n1088# 0.444555f
C127 source.t20 a_n2750_n1088# 0.028286f
C128 source.t21 a_n2750_n1088# 0.028286f
C129 source.n11 a_n2750_n1088# 0.091737f
C130 source.n12 a_n2750_n1088# 0.444555f
C131 source.t24 a_n2750_n1088# 0.028286f
C132 source.t22 a_n2750_n1088# 0.028286f
C133 source.n13 a_n2750_n1088# 0.091737f
C134 source.n14 a_n2750_n1088# 0.444555f
C135 source.t19 a_n2750_n1088# 0.157438f
C136 source.n15 a_n2750_n1088# 1.06227f
C137 source.t1 a_n2750_n1088# 0.157438f
C138 source.n16 a_n2750_n1088# 1.06227f
C139 source.t4 a_n2750_n1088# 0.028286f
C140 source.t11 a_n2750_n1088# 0.028286f
C141 source.n17 a_n2750_n1088# 0.091737f
C142 source.n18 a_n2750_n1088# 0.444555f
C143 source.t6 a_n2750_n1088# 0.028286f
C144 source.t12 a_n2750_n1088# 0.028286f
C145 source.n19 a_n2750_n1088# 0.091737f
C146 source.n20 a_n2750_n1088# 0.444555f
C147 source.t5 a_n2750_n1088# 0.028286f
C148 source.t7 a_n2750_n1088# 0.028286f
C149 source.n21 a_n2750_n1088# 0.091737f
C150 source.n22 a_n2750_n1088# 0.444555f
C151 source.t3 a_n2750_n1088# 0.157438f
C152 source.n23 a_n2750_n1088# 0.397832f
C153 source.t27 a_n2750_n1088# 0.157438f
C154 source.n24 a_n2750_n1088# 0.397832f
C155 source.t17 a_n2750_n1088# 0.028286f
C156 source.t28 a_n2750_n1088# 0.028286f
C157 source.n25 a_n2750_n1088# 0.091737f
C158 source.n26 a_n2750_n1088# 0.444555f
C159 source.t18 a_n2750_n1088# 0.028286f
C160 source.t29 a_n2750_n1088# 0.028286f
C161 source.n27 a_n2750_n1088# 0.091737f
C162 source.n28 a_n2750_n1088# 0.444555f
C163 source.t16 a_n2750_n1088# 0.028286f
C164 source.t30 a_n2750_n1088# 0.028286f
C165 source.n29 a_n2750_n1088# 0.091737f
C166 source.n30 a_n2750_n1088# 0.444555f
C167 source.t15 a_n2750_n1088# 0.157438f
C168 source.n31 a_n2750_n1088# 0.639074f
C169 source.n32 a_n2750_n1088# 0.746207f
C170 drain_right.t12 a_n2750_n1088# 0.015827f
C171 drain_right.t4 a_n2750_n1088# 0.015827f
C172 drain_right.n0 a_n2750_n1088# 0.062607f
C173 drain_right.t6 a_n2750_n1088# 0.015827f
C174 drain_right.t1 a_n2750_n1088# 0.015827f
C175 drain_right.n1 a_n2750_n1088# 0.061501f
C176 drain_right.n2 a_n2750_n1088# 0.50463f
C177 drain_right.t11 a_n2750_n1088# 0.015827f
C178 drain_right.t10 a_n2750_n1088# 0.015827f
C179 drain_right.n3 a_n2750_n1088# 0.062607f
C180 drain_right.t7 a_n2750_n1088# 0.015827f
C181 drain_right.t14 a_n2750_n1088# 0.015827f
C182 drain_right.n4 a_n2750_n1088# 0.061501f
C183 drain_right.n5 a_n2750_n1088# 0.50463f
C184 drain_right.n6 a_n2750_n1088# 0.700713f
C185 drain_right.t2 a_n2750_n1088# 0.015827f
C186 drain_right.t0 a_n2750_n1088# 0.015827f
C187 drain_right.n7 a_n2750_n1088# 0.062607f
C188 drain_right.t9 a_n2750_n1088# 0.015827f
C189 drain_right.t8 a_n2750_n1088# 0.015827f
C190 drain_right.n8 a_n2750_n1088# 0.061501f
C191 drain_right.n9 a_n2750_n1088# 0.53856f
C192 drain_right.t13 a_n2750_n1088# 0.015827f
C193 drain_right.t5 a_n2750_n1088# 0.015827f
C194 drain_right.n10 a_n2750_n1088# 0.061501f
C195 drain_right.n11 a_n2750_n1088# 0.2658f
C196 drain_right.t3 a_n2750_n1088# 0.015827f
C197 drain_right.t15 a_n2750_n1088# 0.015827f
C198 drain_right.n12 a_n2750_n1088# 0.061501f
C199 drain_right.n13 a_n2750_n1088# 0.445397f
C200 minus.n0 a_n2750_n1088# 0.046629f
C201 minus.t8 a_n2750_n1088# 0.094796f
C202 minus.n1 a_n2750_n1088# 0.101022f
C203 minus.t6 a_n2750_n1088# 0.094796f
C204 minus.n2 a_n2750_n1088# 0.034944f
C205 minus.t9 a_n2750_n1088# 0.094796f
C206 minus.n3 a_n2750_n1088# 0.091046f
C207 minus.n4 a_n2750_n1088# 0.200422f
C208 minus.t7 a_n2750_n1088# 0.114529f
C209 minus.n5 a_n2750_n1088# 0.077497f
C210 minus.t5 a_n2750_n1088# 0.094796f
C211 minus.n6 a_n2750_n1088# 0.101296f
C212 minus.t4 a_n2750_n1088# 0.094796f
C213 minus.n7 a_n2750_n1088# 0.101022f
C214 minus.n8 a_n2750_n1088# 0.00793f
C215 minus.n9 a_n2750_n1088# 0.046629f
C216 minus.n10 a_n2750_n1088# 0.034944f
C217 minus.n11 a_n2750_n1088# 0.034944f
C218 minus.n12 a_n2750_n1088# 0.00793f
C219 minus.t10 a_n2750_n1088# 0.094796f
C220 minus.n13 a_n2750_n1088# 0.091046f
C221 minus.n14 a_n2750_n1088# 0.00793f
C222 minus.n15 a_n2750_n1088# 0.046629f
C223 minus.n16 a_n2750_n1088# 0.058204f
C224 minus.n17 a_n2750_n1088# 0.058204f
C225 minus.n18 a_n2750_n1088# 0.100591f
C226 minus.n19 a_n2750_n1088# 0.00793f
C227 minus.t11 a_n2750_n1088# 0.094796f
C228 minus.n20 a_n2750_n1088# 0.087922f
C229 minus.n21 a_n2750_n1088# 0.98458f
C230 minus.n22 a_n2750_n1088# 0.046629f
C231 minus.t14 a_n2750_n1088# 0.094796f
C232 minus.n23 a_n2750_n1088# 0.101022f
C233 minus.n24 a_n2750_n1088# 0.034944f
C234 minus.t12 a_n2750_n1088# 0.094796f
C235 minus.n25 a_n2750_n1088# 0.091046f
C236 minus.n26 a_n2750_n1088# 0.200422f
C237 minus.t3 a_n2750_n1088# 0.114529f
C238 minus.n27 a_n2750_n1088# 0.077497f
C239 minus.t13 a_n2750_n1088# 0.094796f
C240 minus.n28 a_n2750_n1088# 0.101296f
C241 minus.t2 a_n2750_n1088# 0.094796f
C242 minus.n29 a_n2750_n1088# 0.101022f
C243 minus.n30 a_n2750_n1088# 0.00793f
C244 minus.n31 a_n2750_n1088# 0.046629f
C245 minus.n32 a_n2750_n1088# 0.034944f
C246 minus.n33 a_n2750_n1088# 0.034944f
C247 minus.n34 a_n2750_n1088# 0.00793f
C248 minus.t1 a_n2750_n1088# 0.094796f
C249 minus.n35 a_n2750_n1088# 0.091046f
C250 minus.n36 a_n2750_n1088# 0.00793f
C251 minus.n37 a_n2750_n1088# 0.046629f
C252 minus.n38 a_n2750_n1088# 0.058204f
C253 minus.n39 a_n2750_n1088# 0.058204f
C254 minus.t0 a_n2750_n1088# 0.094796f
C255 minus.n40 a_n2750_n1088# 0.100591f
C256 minus.n41 a_n2750_n1088# 0.00793f
C257 minus.t15 a_n2750_n1088# 0.094796f
C258 minus.n42 a_n2750_n1088# 0.087922f
C259 minus.n43 a_n2750_n1088# 0.241189f
C260 minus.n44 a_n2750_n1088# 1.20567f
.ends

