* NGSPICE file created from diffpair258.ext - technology: sky130A

.subckt diffpair258 minus drain_right drain_left source plus
X0 source.t37 minus.t0 drain_right.t7 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X1 source.t36 minus.t1 drain_right.t5 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 source.t9 plus.t0 drain_left.t19 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X3 drain_right.t18 minus.t2 source.t35 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 drain_right.t16 minus.t3 source.t34 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X5 source.t33 minus.t4 drain_right.t15 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X6 drain_left.t18 plus.t1 source.t12 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X8 source.t15 plus.t2 drain_left.t17 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X9 drain_left.t16 plus.t3 source.t8 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X10 source.t11 plus.t4 drain_left.t15 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X11 source.t16 plus.t5 drain_left.t14 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X12 source.t32 minus.t5 drain_right.t9 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X13 source.t17 plus.t6 drain_left.t13 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X14 source.t31 minus.t6 drain_right.t19 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X15 drain_left.t12 plus.t7 source.t2 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X16 source.t30 minus.t7 drain_right.t11 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X17 drain_left.t11 plus.t8 source.t6 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X18 drain_left.t10 plus.t9 source.t1 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X19 source.t5 plus.t10 drain_left.t9 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X20 drain_left.t8 plus.t11 source.t10 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X21 drain_left.t7 plus.t12 source.t13 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X22 drain_left.t6 plus.t13 source.t14 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X23 drain_right.t12 minus.t8 source.t29 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X24 drain_right.t2 minus.t9 source.t28 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X25 drain_right.t3 minus.t10 source.t27 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X26 source.t7 plus.t14 drain_left.t5 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X27 source.t38 plus.t15 drain_left.t4 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X28 a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X29 source.t39 plus.t16 drain_left.t3 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X30 drain_left.t2 plus.t17 source.t4 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X31 source.t26 minus.t11 drain_right.t1 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X32 source.t25 minus.t12 drain_right.t13 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X33 source.t24 minus.t13 drain_right.t14 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X34 source.t23 minus.t14 drain_right.t8 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X35 drain_right.t6 minus.t15 source.t22 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X36 drain_right.t4 minus.t16 source.t21 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X37 a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X38 drain_right.t17 minus.t17 source.t20 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X39 drain_left.t1 plus.t18 source.t0 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X40 source.t3 plus.t19 drain_left.t0 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X41 a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X42 drain_right.t10 minus.t18 source.t19 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X43 drain_right.t0 minus.t19 source.t18 a_n1882_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n23 minus.t7 935.884
R1 minus.n5 minus.t9 935.884
R2 minus.n48 minus.t15 935.884
R3 minus.n30 minus.t12 935.884
R4 minus.n22 minus.t8 879.65
R5 minus.n20 minus.t14 879.65
R6 minus.n1 minus.t3 879.65
R7 minus.n15 minus.t5 879.65
R8 minus.n13 minus.t10 879.65
R9 minus.n3 minus.t13 879.65
R10 minus.n8 minus.t2 879.65
R11 minus.n6 minus.t6 879.65
R12 minus.n47 minus.t0 879.65
R13 minus.n45 minus.t18 879.65
R14 minus.n26 minus.t1 879.65
R15 minus.n40 minus.t19 879.65
R16 minus.n38 minus.t4 879.65
R17 minus.n28 minus.t16 879.65
R18 minus.n33 minus.t11 879.65
R19 minus.n31 minus.t17 879.65
R20 minus.n5 minus.n4 161.489
R21 minus.n30 minus.n29 161.489
R22 minus.n24 minus.n23 161.3
R23 minus.n21 minus.n0 161.3
R24 minus.n19 minus.n18 161.3
R25 minus.n17 minus.n16 161.3
R26 minus.n14 minus.n2 161.3
R27 minus.n12 minus.n11 161.3
R28 minus.n10 minus.n9 161.3
R29 minus.n7 minus.n4 161.3
R30 minus.n49 minus.n48 161.3
R31 minus.n46 minus.n25 161.3
R32 minus.n44 minus.n43 161.3
R33 minus.n42 minus.n41 161.3
R34 minus.n39 minus.n27 161.3
R35 minus.n37 minus.n36 161.3
R36 minus.n35 minus.n34 161.3
R37 minus.n32 minus.n29 161.3
R38 minus.n22 minus.n21 51.852
R39 minus.n7 minus.n6 51.852
R40 minus.n32 minus.n31 51.852
R41 minus.n47 minus.n46 51.852
R42 minus.n20 minus.n19 47.4702
R43 minus.n9 minus.n8 47.4702
R44 minus.n34 minus.n33 47.4702
R45 minus.n45 minus.n44 47.4702
R46 minus.n16 minus.n1 43.0884
R47 minus.n12 minus.n3 43.0884
R48 minus.n37 minus.n28 43.0884
R49 minus.n41 minus.n26 43.0884
R50 minus.n15 minus.n14 38.7066
R51 minus.n14 minus.n13 38.7066
R52 minus.n39 minus.n38 38.7066
R53 minus.n40 minus.n39 38.7066
R54 minus.n16 minus.n15 34.3247
R55 minus.n13 minus.n12 34.3247
R56 minus.n38 minus.n37 34.3247
R57 minus.n41 minus.n40 34.3247
R58 minus.n50 minus.n24 31.6823
R59 minus.n19 minus.n1 29.9429
R60 minus.n9 minus.n3 29.9429
R61 minus.n34 minus.n28 29.9429
R62 minus.n44 minus.n26 29.9429
R63 minus.n21 minus.n20 25.5611
R64 minus.n8 minus.n7 25.5611
R65 minus.n33 minus.n32 25.5611
R66 minus.n46 minus.n45 25.5611
R67 minus.n23 minus.n22 21.1793
R68 minus.n6 minus.n5 21.1793
R69 minus.n31 minus.n30 21.1793
R70 minus.n48 minus.n47 21.1793
R71 minus.n50 minus.n49 6.47777
R72 minus.n24 minus.n0 0.189894
R73 minus.n18 minus.n0 0.189894
R74 minus.n18 minus.n17 0.189894
R75 minus.n17 minus.n2 0.189894
R76 minus.n11 minus.n2 0.189894
R77 minus.n11 minus.n10 0.189894
R78 minus.n10 minus.n4 0.189894
R79 minus.n35 minus.n29 0.189894
R80 minus.n36 minus.n35 0.189894
R81 minus.n36 minus.n27 0.189894
R82 minus.n42 minus.n27 0.189894
R83 minus.n43 minus.n42 0.189894
R84 minus.n43 minus.n25 0.189894
R85 minus.n49 minus.n25 0.189894
R86 minus minus.n50 0.188
R87 drain_right.n6 drain_right.n4 67.6476
R88 drain_right.n2 drain_right.n0 67.6476
R89 drain_right.n10 drain_right.n8 67.6476
R90 drain_right.n10 drain_right.n9 67.1908
R91 drain_right.n12 drain_right.n11 67.1908
R92 drain_right.n14 drain_right.n13 67.1908
R93 drain_right.n16 drain_right.n15 67.1908
R94 drain_right.n7 drain_right.n3 67.1907
R95 drain_right.n6 drain_right.n5 67.1907
R96 drain_right.n2 drain_right.n1 67.1907
R97 drain_right drain_right.n7 25.9236
R98 drain_right drain_right.n16 6.11011
R99 drain_right.n3 drain_right.t15 3.3005
R100 drain_right.n3 drain_right.t0 3.3005
R101 drain_right.n4 drain_right.t7 3.3005
R102 drain_right.n4 drain_right.t6 3.3005
R103 drain_right.n5 drain_right.t5 3.3005
R104 drain_right.n5 drain_right.t10 3.3005
R105 drain_right.n1 drain_right.t1 3.3005
R106 drain_right.n1 drain_right.t4 3.3005
R107 drain_right.n0 drain_right.t13 3.3005
R108 drain_right.n0 drain_right.t17 3.3005
R109 drain_right.n8 drain_right.t19 3.3005
R110 drain_right.n8 drain_right.t2 3.3005
R111 drain_right.n9 drain_right.t14 3.3005
R112 drain_right.n9 drain_right.t18 3.3005
R113 drain_right.n11 drain_right.t9 3.3005
R114 drain_right.n11 drain_right.t3 3.3005
R115 drain_right.n13 drain_right.t8 3.3005
R116 drain_right.n13 drain_right.t16 3.3005
R117 drain_right.n15 drain_right.t11 3.3005
R118 drain_right.n15 drain_right.t12 3.3005
R119 drain_right.n16 drain_right.n14 0.457397
R120 drain_right.n14 drain_right.n12 0.457397
R121 drain_right.n12 drain_right.n10 0.457397
R122 drain_right.n7 drain_right.n6 0.402051
R123 drain_right.n7 drain_right.n2 0.402051
R124 source.n282 source.n256 289.615
R125 source.n242 source.n216 289.615
R126 source.n210 source.n184 289.615
R127 source.n170 source.n144 289.615
R128 source.n26 source.n0 289.615
R129 source.n66 source.n40 289.615
R130 source.n98 source.n72 289.615
R131 source.n138 source.n112 289.615
R132 source.n267 source.n266 185
R133 source.n264 source.n263 185
R134 source.n273 source.n272 185
R135 source.n275 source.n274 185
R136 source.n260 source.n259 185
R137 source.n281 source.n280 185
R138 source.n283 source.n282 185
R139 source.n227 source.n226 185
R140 source.n224 source.n223 185
R141 source.n233 source.n232 185
R142 source.n235 source.n234 185
R143 source.n220 source.n219 185
R144 source.n241 source.n240 185
R145 source.n243 source.n242 185
R146 source.n195 source.n194 185
R147 source.n192 source.n191 185
R148 source.n201 source.n200 185
R149 source.n203 source.n202 185
R150 source.n188 source.n187 185
R151 source.n209 source.n208 185
R152 source.n211 source.n210 185
R153 source.n155 source.n154 185
R154 source.n152 source.n151 185
R155 source.n161 source.n160 185
R156 source.n163 source.n162 185
R157 source.n148 source.n147 185
R158 source.n169 source.n168 185
R159 source.n171 source.n170 185
R160 source.n27 source.n26 185
R161 source.n25 source.n24 185
R162 source.n4 source.n3 185
R163 source.n19 source.n18 185
R164 source.n17 source.n16 185
R165 source.n8 source.n7 185
R166 source.n11 source.n10 185
R167 source.n67 source.n66 185
R168 source.n65 source.n64 185
R169 source.n44 source.n43 185
R170 source.n59 source.n58 185
R171 source.n57 source.n56 185
R172 source.n48 source.n47 185
R173 source.n51 source.n50 185
R174 source.n99 source.n98 185
R175 source.n97 source.n96 185
R176 source.n76 source.n75 185
R177 source.n91 source.n90 185
R178 source.n89 source.n88 185
R179 source.n80 source.n79 185
R180 source.n83 source.n82 185
R181 source.n139 source.n138 185
R182 source.n137 source.n136 185
R183 source.n116 source.n115 185
R184 source.n131 source.n130 185
R185 source.n129 source.n128 185
R186 source.n120 source.n119 185
R187 source.n123 source.n122 185
R188 source.t22 source.n265 147.661
R189 source.t25 source.n225 147.661
R190 source.t14 source.n193 147.661
R191 source.t9 source.n153 147.661
R192 source.t2 source.n9 147.661
R193 source.t5 source.n49 147.661
R194 source.t28 source.n81 147.661
R195 source.t30 source.n121 147.661
R196 source.n266 source.n263 104.615
R197 source.n273 source.n263 104.615
R198 source.n274 source.n273 104.615
R199 source.n274 source.n259 104.615
R200 source.n281 source.n259 104.615
R201 source.n282 source.n281 104.615
R202 source.n226 source.n223 104.615
R203 source.n233 source.n223 104.615
R204 source.n234 source.n233 104.615
R205 source.n234 source.n219 104.615
R206 source.n241 source.n219 104.615
R207 source.n242 source.n241 104.615
R208 source.n194 source.n191 104.615
R209 source.n201 source.n191 104.615
R210 source.n202 source.n201 104.615
R211 source.n202 source.n187 104.615
R212 source.n209 source.n187 104.615
R213 source.n210 source.n209 104.615
R214 source.n154 source.n151 104.615
R215 source.n161 source.n151 104.615
R216 source.n162 source.n161 104.615
R217 source.n162 source.n147 104.615
R218 source.n169 source.n147 104.615
R219 source.n170 source.n169 104.615
R220 source.n26 source.n25 104.615
R221 source.n25 source.n3 104.615
R222 source.n18 source.n3 104.615
R223 source.n18 source.n17 104.615
R224 source.n17 source.n7 104.615
R225 source.n10 source.n7 104.615
R226 source.n66 source.n65 104.615
R227 source.n65 source.n43 104.615
R228 source.n58 source.n43 104.615
R229 source.n58 source.n57 104.615
R230 source.n57 source.n47 104.615
R231 source.n50 source.n47 104.615
R232 source.n98 source.n97 104.615
R233 source.n97 source.n75 104.615
R234 source.n90 source.n75 104.615
R235 source.n90 source.n89 104.615
R236 source.n89 source.n79 104.615
R237 source.n82 source.n79 104.615
R238 source.n138 source.n137 104.615
R239 source.n137 source.n115 104.615
R240 source.n130 source.n115 104.615
R241 source.n130 source.n129 104.615
R242 source.n129 source.n119 104.615
R243 source.n122 source.n119 104.615
R244 source.n266 source.t22 52.3082
R245 source.n226 source.t25 52.3082
R246 source.n194 source.t14 52.3082
R247 source.n154 source.t9 52.3082
R248 source.n10 source.t2 52.3082
R249 source.n50 source.t5 52.3082
R250 source.n82 source.t28 52.3082
R251 source.n122 source.t30 52.3082
R252 source.n33 source.n32 50.512
R253 source.n35 source.n34 50.512
R254 source.n37 source.n36 50.512
R255 source.n39 source.n38 50.512
R256 source.n105 source.n104 50.512
R257 source.n107 source.n106 50.512
R258 source.n109 source.n108 50.512
R259 source.n111 source.n110 50.512
R260 source.n255 source.n254 50.5119
R261 source.n253 source.n252 50.5119
R262 source.n251 source.n250 50.5119
R263 source.n249 source.n248 50.5119
R264 source.n183 source.n182 50.5119
R265 source.n181 source.n180 50.5119
R266 source.n179 source.n178 50.5119
R267 source.n177 source.n176 50.5119
R268 source.n287 source.n286 32.1853
R269 source.n247 source.n246 32.1853
R270 source.n215 source.n214 32.1853
R271 source.n175 source.n174 32.1853
R272 source.n31 source.n30 32.1853
R273 source.n71 source.n70 32.1853
R274 source.n103 source.n102 32.1853
R275 source.n143 source.n142 32.1853
R276 source.n175 source.n143 17.1992
R277 source.n267 source.n265 15.6674
R278 source.n227 source.n225 15.6674
R279 source.n195 source.n193 15.6674
R280 source.n155 source.n153 15.6674
R281 source.n11 source.n9 15.6674
R282 source.n51 source.n49 15.6674
R283 source.n83 source.n81 15.6674
R284 source.n123 source.n121 15.6674
R285 source.n268 source.n264 12.8005
R286 source.n228 source.n224 12.8005
R287 source.n196 source.n192 12.8005
R288 source.n156 source.n152 12.8005
R289 source.n12 source.n8 12.8005
R290 source.n52 source.n48 12.8005
R291 source.n84 source.n80 12.8005
R292 source.n124 source.n120 12.8005
R293 source.n272 source.n271 12.0247
R294 source.n232 source.n231 12.0247
R295 source.n200 source.n199 12.0247
R296 source.n160 source.n159 12.0247
R297 source.n16 source.n15 12.0247
R298 source.n56 source.n55 12.0247
R299 source.n88 source.n87 12.0247
R300 source.n128 source.n127 12.0247
R301 source.n288 source.n31 11.7078
R302 source.n275 source.n262 11.249
R303 source.n235 source.n222 11.249
R304 source.n203 source.n190 11.249
R305 source.n163 source.n150 11.249
R306 source.n19 source.n6 11.249
R307 source.n59 source.n46 11.249
R308 source.n91 source.n78 11.249
R309 source.n131 source.n118 11.249
R310 source.n276 source.n260 10.4732
R311 source.n236 source.n220 10.4732
R312 source.n204 source.n188 10.4732
R313 source.n164 source.n148 10.4732
R314 source.n20 source.n4 10.4732
R315 source.n60 source.n44 10.4732
R316 source.n92 source.n76 10.4732
R317 source.n132 source.n116 10.4732
R318 source.n280 source.n279 9.69747
R319 source.n240 source.n239 9.69747
R320 source.n208 source.n207 9.69747
R321 source.n168 source.n167 9.69747
R322 source.n24 source.n23 9.69747
R323 source.n64 source.n63 9.69747
R324 source.n96 source.n95 9.69747
R325 source.n136 source.n135 9.69747
R326 source.n286 source.n285 9.45567
R327 source.n246 source.n245 9.45567
R328 source.n214 source.n213 9.45567
R329 source.n174 source.n173 9.45567
R330 source.n30 source.n29 9.45567
R331 source.n70 source.n69 9.45567
R332 source.n102 source.n101 9.45567
R333 source.n142 source.n141 9.45567
R334 source.n285 source.n284 9.3005
R335 source.n258 source.n257 9.3005
R336 source.n279 source.n278 9.3005
R337 source.n277 source.n276 9.3005
R338 source.n262 source.n261 9.3005
R339 source.n271 source.n270 9.3005
R340 source.n269 source.n268 9.3005
R341 source.n245 source.n244 9.3005
R342 source.n218 source.n217 9.3005
R343 source.n239 source.n238 9.3005
R344 source.n237 source.n236 9.3005
R345 source.n222 source.n221 9.3005
R346 source.n231 source.n230 9.3005
R347 source.n229 source.n228 9.3005
R348 source.n213 source.n212 9.3005
R349 source.n186 source.n185 9.3005
R350 source.n207 source.n206 9.3005
R351 source.n205 source.n204 9.3005
R352 source.n190 source.n189 9.3005
R353 source.n199 source.n198 9.3005
R354 source.n197 source.n196 9.3005
R355 source.n173 source.n172 9.3005
R356 source.n146 source.n145 9.3005
R357 source.n167 source.n166 9.3005
R358 source.n165 source.n164 9.3005
R359 source.n150 source.n149 9.3005
R360 source.n159 source.n158 9.3005
R361 source.n157 source.n156 9.3005
R362 source.n29 source.n28 9.3005
R363 source.n2 source.n1 9.3005
R364 source.n23 source.n22 9.3005
R365 source.n21 source.n20 9.3005
R366 source.n6 source.n5 9.3005
R367 source.n15 source.n14 9.3005
R368 source.n13 source.n12 9.3005
R369 source.n69 source.n68 9.3005
R370 source.n42 source.n41 9.3005
R371 source.n63 source.n62 9.3005
R372 source.n61 source.n60 9.3005
R373 source.n46 source.n45 9.3005
R374 source.n55 source.n54 9.3005
R375 source.n53 source.n52 9.3005
R376 source.n101 source.n100 9.3005
R377 source.n74 source.n73 9.3005
R378 source.n95 source.n94 9.3005
R379 source.n93 source.n92 9.3005
R380 source.n78 source.n77 9.3005
R381 source.n87 source.n86 9.3005
R382 source.n85 source.n84 9.3005
R383 source.n141 source.n140 9.3005
R384 source.n114 source.n113 9.3005
R385 source.n135 source.n134 9.3005
R386 source.n133 source.n132 9.3005
R387 source.n118 source.n117 9.3005
R388 source.n127 source.n126 9.3005
R389 source.n125 source.n124 9.3005
R390 source.n283 source.n258 8.92171
R391 source.n243 source.n218 8.92171
R392 source.n211 source.n186 8.92171
R393 source.n171 source.n146 8.92171
R394 source.n27 source.n2 8.92171
R395 source.n67 source.n42 8.92171
R396 source.n99 source.n74 8.92171
R397 source.n139 source.n114 8.92171
R398 source.n284 source.n256 8.14595
R399 source.n244 source.n216 8.14595
R400 source.n212 source.n184 8.14595
R401 source.n172 source.n144 8.14595
R402 source.n28 source.n0 8.14595
R403 source.n68 source.n40 8.14595
R404 source.n100 source.n72 8.14595
R405 source.n140 source.n112 8.14595
R406 source.n286 source.n256 5.81868
R407 source.n246 source.n216 5.81868
R408 source.n214 source.n184 5.81868
R409 source.n174 source.n144 5.81868
R410 source.n30 source.n0 5.81868
R411 source.n70 source.n40 5.81868
R412 source.n102 source.n72 5.81868
R413 source.n142 source.n112 5.81868
R414 source.n288 source.n287 5.49188
R415 source.n284 source.n283 5.04292
R416 source.n244 source.n243 5.04292
R417 source.n212 source.n211 5.04292
R418 source.n172 source.n171 5.04292
R419 source.n28 source.n27 5.04292
R420 source.n68 source.n67 5.04292
R421 source.n100 source.n99 5.04292
R422 source.n140 source.n139 5.04292
R423 source.n269 source.n265 4.38594
R424 source.n229 source.n225 4.38594
R425 source.n197 source.n193 4.38594
R426 source.n157 source.n153 4.38594
R427 source.n13 source.n9 4.38594
R428 source.n53 source.n49 4.38594
R429 source.n85 source.n81 4.38594
R430 source.n125 source.n121 4.38594
R431 source.n280 source.n258 4.26717
R432 source.n240 source.n218 4.26717
R433 source.n208 source.n186 4.26717
R434 source.n168 source.n146 4.26717
R435 source.n24 source.n2 4.26717
R436 source.n64 source.n42 4.26717
R437 source.n96 source.n74 4.26717
R438 source.n136 source.n114 4.26717
R439 source.n279 source.n260 3.49141
R440 source.n239 source.n220 3.49141
R441 source.n207 source.n188 3.49141
R442 source.n167 source.n148 3.49141
R443 source.n23 source.n4 3.49141
R444 source.n63 source.n44 3.49141
R445 source.n95 source.n76 3.49141
R446 source.n135 source.n116 3.49141
R447 source.n254 source.t19 3.3005
R448 source.n254 source.t37 3.3005
R449 source.n252 source.t18 3.3005
R450 source.n252 source.t36 3.3005
R451 source.n250 source.t21 3.3005
R452 source.n250 source.t33 3.3005
R453 source.n248 source.t20 3.3005
R454 source.n248 source.t26 3.3005
R455 source.n182 source.t10 3.3005
R456 source.n182 source.t7 3.3005
R457 source.n180 source.t13 3.3005
R458 source.n180 source.t17 3.3005
R459 source.n178 source.t6 3.3005
R460 source.n178 source.t16 3.3005
R461 source.n176 source.t12 3.3005
R462 source.n176 source.t11 3.3005
R463 source.n32 source.t0 3.3005
R464 source.n32 source.t38 3.3005
R465 source.n34 source.t1 3.3005
R466 source.n34 source.t15 3.3005
R467 source.n36 source.t4 3.3005
R468 source.n36 source.t39 3.3005
R469 source.n38 source.t8 3.3005
R470 source.n38 source.t3 3.3005
R471 source.n104 source.t35 3.3005
R472 source.n104 source.t31 3.3005
R473 source.n106 source.t27 3.3005
R474 source.n106 source.t24 3.3005
R475 source.n108 source.t34 3.3005
R476 source.n108 source.t32 3.3005
R477 source.n110 source.t29 3.3005
R478 source.n110 source.t23 3.3005
R479 source.n276 source.n275 2.71565
R480 source.n236 source.n235 2.71565
R481 source.n204 source.n203 2.71565
R482 source.n164 source.n163 2.71565
R483 source.n20 source.n19 2.71565
R484 source.n60 source.n59 2.71565
R485 source.n92 source.n91 2.71565
R486 source.n132 source.n131 2.71565
R487 source.n272 source.n262 1.93989
R488 source.n232 source.n222 1.93989
R489 source.n200 source.n190 1.93989
R490 source.n160 source.n150 1.93989
R491 source.n16 source.n6 1.93989
R492 source.n56 source.n46 1.93989
R493 source.n88 source.n78 1.93989
R494 source.n128 source.n118 1.93989
R495 source.n271 source.n264 1.16414
R496 source.n231 source.n224 1.16414
R497 source.n199 source.n192 1.16414
R498 source.n159 source.n152 1.16414
R499 source.n15 source.n8 1.16414
R500 source.n55 source.n48 1.16414
R501 source.n87 source.n80 1.16414
R502 source.n127 source.n120 1.16414
R503 source.n103 source.n71 0.470328
R504 source.n247 source.n215 0.470328
R505 source.n143 source.n111 0.457397
R506 source.n111 source.n109 0.457397
R507 source.n109 source.n107 0.457397
R508 source.n107 source.n105 0.457397
R509 source.n105 source.n103 0.457397
R510 source.n71 source.n39 0.457397
R511 source.n39 source.n37 0.457397
R512 source.n37 source.n35 0.457397
R513 source.n35 source.n33 0.457397
R514 source.n33 source.n31 0.457397
R515 source.n177 source.n175 0.457397
R516 source.n179 source.n177 0.457397
R517 source.n181 source.n179 0.457397
R518 source.n183 source.n181 0.457397
R519 source.n215 source.n183 0.457397
R520 source.n249 source.n247 0.457397
R521 source.n251 source.n249 0.457397
R522 source.n253 source.n251 0.457397
R523 source.n255 source.n253 0.457397
R524 source.n287 source.n255 0.457397
R525 source.n268 source.n267 0.388379
R526 source.n228 source.n227 0.388379
R527 source.n196 source.n195 0.388379
R528 source.n156 source.n155 0.388379
R529 source.n12 source.n11 0.388379
R530 source.n52 source.n51 0.388379
R531 source.n84 source.n83 0.388379
R532 source.n124 source.n123 0.388379
R533 source source.n288 0.188
R534 source.n270 source.n269 0.155672
R535 source.n270 source.n261 0.155672
R536 source.n277 source.n261 0.155672
R537 source.n278 source.n277 0.155672
R538 source.n278 source.n257 0.155672
R539 source.n285 source.n257 0.155672
R540 source.n230 source.n229 0.155672
R541 source.n230 source.n221 0.155672
R542 source.n237 source.n221 0.155672
R543 source.n238 source.n237 0.155672
R544 source.n238 source.n217 0.155672
R545 source.n245 source.n217 0.155672
R546 source.n198 source.n197 0.155672
R547 source.n198 source.n189 0.155672
R548 source.n205 source.n189 0.155672
R549 source.n206 source.n205 0.155672
R550 source.n206 source.n185 0.155672
R551 source.n213 source.n185 0.155672
R552 source.n158 source.n157 0.155672
R553 source.n158 source.n149 0.155672
R554 source.n165 source.n149 0.155672
R555 source.n166 source.n165 0.155672
R556 source.n166 source.n145 0.155672
R557 source.n173 source.n145 0.155672
R558 source.n29 source.n1 0.155672
R559 source.n22 source.n1 0.155672
R560 source.n22 source.n21 0.155672
R561 source.n21 source.n5 0.155672
R562 source.n14 source.n5 0.155672
R563 source.n14 source.n13 0.155672
R564 source.n69 source.n41 0.155672
R565 source.n62 source.n41 0.155672
R566 source.n62 source.n61 0.155672
R567 source.n61 source.n45 0.155672
R568 source.n54 source.n45 0.155672
R569 source.n54 source.n53 0.155672
R570 source.n101 source.n73 0.155672
R571 source.n94 source.n73 0.155672
R572 source.n94 source.n93 0.155672
R573 source.n93 source.n77 0.155672
R574 source.n86 source.n77 0.155672
R575 source.n86 source.n85 0.155672
R576 source.n141 source.n113 0.155672
R577 source.n134 source.n113 0.155672
R578 source.n134 source.n133 0.155672
R579 source.n133 source.n117 0.155672
R580 source.n126 source.n117 0.155672
R581 source.n126 source.n125 0.155672
R582 plus.n5 plus.t10 935.884
R583 plus.n23 plus.t7 935.884
R584 plus.n30 plus.t13 935.884
R585 plus.n48 plus.t0 935.884
R586 plus.n6 plus.t3 879.65
R587 plus.n8 plus.t19 879.65
R588 plus.n3 plus.t17 879.65
R589 plus.n13 plus.t16 879.65
R590 plus.n15 plus.t9 879.65
R591 plus.n1 plus.t2 879.65
R592 plus.n20 plus.t18 879.65
R593 plus.n22 plus.t15 879.65
R594 plus.n31 plus.t14 879.65
R595 plus.n33 plus.t11 879.65
R596 plus.n28 plus.t6 879.65
R597 plus.n38 plus.t12 879.65
R598 plus.n40 plus.t5 879.65
R599 plus.n26 plus.t8 879.65
R600 plus.n45 plus.t4 879.65
R601 plus.n47 plus.t1 879.65
R602 plus.n5 plus.n4 161.489
R603 plus.n30 plus.n29 161.489
R604 plus.n7 plus.n4 161.3
R605 plus.n10 plus.n9 161.3
R606 plus.n12 plus.n11 161.3
R607 plus.n14 plus.n2 161.3
R608 plus.n17 plus.n16 161.3
R609 plus.n19 plus.n18 161.3
R610 plus.n21 plus.n0 161.3
R611 plus.n24 plus.n23 161.3
R612 plus.n32 plus.n29 161.3
R613 plus.n35 plus.n34 161.3
R614 plus.n37 plus.n36 161.3
R615 plus.n39 plus.n27 161.3
R616 plus.n42 plus.n41 161.3
R617 plus.n44 plus.n43 161.3
R618 plus.n46 plus.n25 161.3
R619 plus.n49 plus.n48 161.3
R620 plus.n7 plus.n6 51.852
R621 plus.n22 plus.n21 51.852
R622 plus.n47 plus.n46 51.852
R623 plus.n32 plus.n31 51.852
R624 plus.n9 plus.n8 47.4702
R625 plus.n20 plus.n19 47.4702
R626 plus.n45 plus.n44 47.4702
R627 plus.n34 plus.n33 47.4702
R628 plus.n12 plus.n3 43.0884
R629 plus.n16 plus.n1 43.0884
R630 plus.n41 plus.n26 43.0884
R631 plus.n37 plus.n28 43.0884
R632 plus.n14 plus.n13 38.7066
R633 plus.n15 plus.n14 38.7066
R634 plus.n40 plus.n39 38.7066
R635 plus.n39 plus.n38 38.7066
R636 plus.n13 plus.n12 34.3247
R637 plus.n16 plus.n15 34.3247
R638 plus.n41 plus.n40 34.3247
R639 plus.n38 plus.n37 34.3247
R640 plus.n9 plus.n3 29.9429
R641 plus.n19 plus.n1 29.9429
R642 plus.n44 plus.n26 29.9429
R643 plus.n34 plus.n28 29.9429
R644 plus plus.n49 27.8361
R645 plus.n8 plus.n7 25.5611
R646 plus.n21 plus.n20 25.5611
R647 plus.n46 plus.n45 25.5611
R648 plus.n33 plus.n32 25.5611
R649 plus.n6 plus.n5 21.1793
R650 plus.n23 plus.n22 21.1793
R651 plus.n48 plus.n47 21.1793
R652 plus.n31 plus.n30 21.1793
R653 plus plus.n24 9.84898
R654 plus.n10 plus.n4 0.189894
R655 plus.n11 plus.n10 0.189894
R656 plus.n11 plus.n2 0.189894
R657 plus.n17 plus.n2 0.189894
R658 plus.n18 plus.n17 0.189894
R659 plus.n18 plus.n0 0.189894
R660 plus.n24 plus.n0 0.189894
R661 plus.n49 plus.n25 0.189894
R662 plus.n43 plus.n25 0.189894
R663 plus.n43 plus.n42 0.189894
R664 plus.n42 plus.n27 0.189894
R665 plus.n36 plus.n27 0.189894
R666 plus.n36 plus.n35 0.189894
R667 plus.n35 plus.n29 0.189894
R668 drain_left.n10 drain_left.n8 67.6477
R669 drain_left.n6 drain_left.n4 67.6476
R670 drain_left.n2 drain_left.n0 67.6476
R671 drain_left.n14 drain_left.n13 67.1908
R672 drain_left.n12 drain_left.n11 67.1908
R673 drain_left.n10 drain_left.n9 67.1908
R674 drain_left.n16 drain_left.n15 67.1907
R675 drain_left.n7 drain_left.n3 67.1907
R676 drain_left.n6 drain_left.n5 67.1907
R677 drain_left.n2 drain_left.n1 67.1907
R678 drain_left drain_left.n7 26.4768
R679 drain_left drain_left.n16 6.11011
R680 drain_left.n3 drain_left.t14 3.3005
R681 drain_left.n3 drain_left.t7 3.3005
R682 drain_left.n4 drain_left.t5 3.3005
R683 drain_left.n4 drain_left.t6 3.3005
R684 drain_left.n5 drain_left.t13 3.3005
R685 drain_left.n5 drain_left.t8 3.3005
R686 drain_left.n1 drain_left.t15 3.3005
R687 drain_left.n1 drain_left.t11 3.3005
R688 drain_left.n0 drain_left.t19 3.3005
R689 drain_left.n0 drain_left.t18 3.3005
R690 drain_left.n15 drain_left.t4 3.3005
R691 drain_left.n15 drain_left.t12 3.3005
R692 drain_left.n13 drain_left.t17 3.3005
R693 drain_left.n13 drain_left.t1 3.3005
R694 drain_left.n11 drain_left.t3 3.3005
R695 drain_left.n11 drain_left.t10 3.3005
R696 drain_left.n9 drain_left.t0 3.3005
R697 drain_left.n9 drain_left.t2 3.3005
R698 drain_left.n8 drain_left.t9 3.3005
R699 drain_left.n8 drain_left.t16 3.3005
R700 drain_left.n12 drain_left.n10 0.457397
R701 drain_left.n14 drain_left.n12 0.457397
R702 drain_left.n16 drain_left.n14 0.457397
R703 drain_left.n7 drain_left.n6 0.402051
R704 drain_left.n7 drain_left.n2 0.402051
C0 minus drain_left 0.171252f
C1 minus drain_right 2.95061f
C2 minus source 2.89794f
C3 drain_left plus 3.13367f
C4 plus drain_right 0.337271f
C5 drain_left drain_right 0.982035f
C6 source plus 2.91196f
C7 source drain_left 24.1909f
C8 source drain_right 24.1909f
C9 minus plus 4.39056f
C10 drain_right a_n1882_n2088# 5.63585f
C11 drain_left a_n1882_n2088# 5.92877f
C12 source a_n1882_n2088# 5.320182f
C13 minus a_n1882_n2088# 6.840036f
C14 plus a_n1882_n2088# 8.50321f
C15 drain_left.t19 a_n1882_n2088# 0.180092f
C16 drain_left.t18 a_n1882_n2088# 0.180092f
C17 drain_left.n0 a_n1882_n2088# 1.50491f
C18 drain_left.t15 a_n1882_n2088# 0.180092f
C19 drain_left.t11 a_n1882_n2088# 0.180092f
C20 drain_left.n1 a_n1882_n2088# 1.50197f
C21 drain_left.n2 a_n1882_n2088# 0.84802f
C22 drain_left.t14 a_n1882_n2088# 0.180092f
C23 drain_left.t7 a_n1882_n2088# 0.180092f
C24 drain_left.n3 a_n1882_n2088# 1.50197f
C25 drain_left.t5 a_n1882_n2088# 0.180092f
C26 drain_left.t6 a_n1882_n2088# 0.180092f
C27 drain_left.n4 a_n1882_n2088# 1.50491f
C28 drain_left.t13 a_n1882_n2088# 0.180092f
C29 drain_left.t8 a_n1882_n2088# 0.180092f
C30 drain_left.n5 a_n1882_n2088# 1.50197f
C31 drain_left.n6 a_n1882_n2088# 0.84802f
C32 drain_left.n7 a_n1882_n2088# 1.73895f
C33 drain_left.t9 a_n1882_n2088# 0.180092f
C34 drain_left.t16 a_n1882_n2088# 0.180092f
C35 drain_left.n8 a_n1882_n2088# 1.50491f
C36 drain_left.t0 a_n1882_n2088# 0.180092f
C37 drain_left.t2 a_n1882_n2088# 0.180092f
C38 drain_left.n9 a_n1882_n2088# 1.50197f
C39 drain_left.n10 a_n1882_n2088# 0.852587f
C40 drain_left.t3 a_n1882_n2088# 0.180092f
C41 drain_left.t10 a_n1882_n2088# 0.180092f
C42 drain_left.n11 a_n1882_n2088# 1.50197f
C43 drain_left.n12 a_n1882_n2088# 0.420115f
C44 drain_left.t17 a_n1882_n2088# 0.180092f
C45 drain_left.t1 a_n1882_n2088# 0.180092f
C46 drain_left.n13 a_n1882_n2088# 1.50197f
C47 drain_left.n14 a_n1882_n2088# 0.420115f
C48 drain_left.t4 a_n1882_n2088# 0.180092f
C49 drain_left.t12 a_n1882_n2088# 0.180092f
C50 drain_left.n15 a_n1882_n2088# 1.50197f
C51 drain_left.n16 a_n1882_n2088# 0.730976f
C52 plus.n0 a_n1882_n2088# 0.053719f
C53 plus.t15 a_n1882_n2088# 0.183666f
C54 plus.t18 a_n1882_n2088# 0.183666f
C55 plus.t2 a_n1882_n2088# 0.183666f
C56 plus.n1 a_n1882_n2088# 0.089826f
C57 plus.n2 a_n1882_n2088# 0.053719f
C58 plus.t9 a_n1882_n2088# 0.183666f
C59 plus.t16 a_n1882_n2088# 0.183666f
C60 plus.t17 a_n1882_n2088# 0.183666f
C61 plus.n3 a_n1882_n2088# 0.089826f
C62 plus.n4 a_n1882_n2088# 0.122923f
C63 plus.t19 a_n1882_n2088# 0.183666f
C64 plus.t3 a_n1882_n2088# 0.183666f
C65 plus.t10 a_n1882_n2088# 0.189232f
C66 plus.n5 a_n1882_n2088# 0.10597f
C67 plus.n6 a_n1882_n2088# 0.089826f
C68 plus.n7 a_n1882_n2088# 0.018814f
C69 plus.n8 a_n1882_n2088# 0.089826f
C70 plus.n9 a_n1882_n2088# 0.018814f
C71 plus.n10 a_n1882_n2088# 0.053719f
C72 plus.n11 a_n1882_n2088# 0.053719f
C73 plus.n12 a_n1882_n2088# 0.018814f
C74 plus.n13 a_n1882_n2088# 0.089826f
C75 plus.n14 a_n1882_n2088# 0.018814f
C76 plus.n15 a_n1882_n2088# 0.089826f
C77 plus.n16 a_n1882_n2088# 0.018814f
C78 plus.n17 a_n1882_n2088# 0.053719f
C79 plus.n18 a_n1882_n2088# 0.053719f
C80 plus.n19 a_n1882_n2088# 0.018814f
C81 plus.n20 a_n1882_n2088# 0.089826f
C82 plus.n21 a_n1882_n2088# 0.018814f
C83 plus.n22 a_n1882_n2088# 0.089826f
C84 plus.t7 a_n1882_n2088# 0.189232f
C85 plus.n23 a_n1882_n2088# 0.105888f
C86 plus.n24 a_n1882_n2088# 0.457379f
C87 plus.n25 a_n1882_n2088# 0.053719f
C88 plus.t0 a_n1882_n2088# 0.189232f
C89 plus.t1 a_n1882_n2088# 0.183666f
C90 plus.t4 a_n1882_n2088# 0.183666f
C91 plus.t8 a_n1882_n2088# 0.183666f
C92 plus.n26 a_n1882_n2088# 0.089826f
C93 plus.n27 a_n1882_n2088# 0.053719f
C94 plus.t5 a_n1882_n2088# 0.183666f
C95 plus.t12 a_n1882_n2088# 0.183666f
C96 plus.t6 a_n1882_n2088# 0.183666f
C97 plus.n28 a_n1882_n2088# 0.089826f
C98 plus.n29 a_n1882_n2088# 0.122923f
C99 plus.t11 a_n1882_n2088# 0.183666f
C100 plus.t14 a_n1882_n2088# 0.183666f
C101 plus.t13 a_n1882_n2088# 0.189232f
C102 plus.n30 a_n1882_n2088# 0.10597f
C103 plus.n31 a_n1882_n2088# 0.089826f
C104 plus.n32 a_n1882_n2088# 0.018814f
C105 plus.n33 a_n1882_n2088# 0.089826f
C106 plus.n34 a_n1882_n2088# 0.018814f
C107 plus.n35 a_n1882_n2088# 0.053719f
C108 plus.n36 a_n1882_n2088# 0.053719f
C109 plus.n37 a_n1882_n2088# 0.018814f
C110 plus.n38 a_n1882_n2088# 0.089826f
C111 plus.n39 a_n1882_n2088# 0.018814f
C112 plus.n40 a_n1882_n2088# 0.089826f
C113 plus.n41 a_n1882_n2088# 0.018814f
C114 plus.n42 a_n1882_n2088# 0.053719f
C115 plus.n43 a_n1882_n2088# 0.053719f
C116 plus.n44 a_n1882_n2088# 0.018814f
C117 plus.n45 a_n1882_n2088# 0.089826f
C118 plus.n46 a_n1882_n2088# 0.018814f
C119 plus.n47 a_n1882_n2088# 0.089826f
C120 plus.n48 a_n1882_n2088# 0.105888f
C121 plus.n49 a_n1882_n2088# 1.38269f
C122 source.n0 a_n1882_n2088# 0.048506f
C123 source.n1 a_n1882_n2088# 0.03451f
C124 source.n2 a_n1882_n2088# 0.018544f
C125 source.n3 a_n1882_n2088# 0.043831f
C126 source.n4 a_n1882_n2088# 0.019635f
C127 source.n5 a_n1882_n2088# 0.03451f
C128 source.n6 a_n1882_n2088# 0.018544f
C129 source.n7 a_n1882_n2088# 0.043831f
C130 source.n8 a_n1882_n2088# 0.019635f
C131 source.n9 a_n1882_n2088# 0.147677f
C132 source.t2 a_n1882_n2088# 0.071439f
C133 source.n10 a_n1882_n2088# 0.032873f
C134 source.n11 a_n1882_n2088# 0.025891f
C135 source.n12 a_n1882_n2088# 0.018544f
C136 source.n13 a_n1882_n2088# 0.821123f
C137 source.n14 a_n1882_n2088# 0.03451f
C138 source.n15 a_n1882_n2088# 0.018544f
C139 source.n16 a_n1882_n2088# 0.019635f
C140 source.n17 a_n1882_n2088# 0.043831f
C141 source.n18 a_n1882_n2088# 0.043831f
C142 source.n19 a_n1882_n2088# 0.019635f
C143 source.n20 a_n1882_n2088# 0.018544f
C144 source.n21 a_n1882_n2088# 0.03451f
C145 source.n22 a_n1882_n2088# 0.03451f
C146 source.n23 a_n1882_n2088# 0.018544f
C147 source.n24 a_n1882_n2088# 0.019635f
C148 source.n25 a_n1882_n2088# 0.043831f
C149 source.n26 a_n1882_n2088# 0.094887f
C150 source.n27 a_n1882_n2088# 0.019635f
C151 source.n28 a_n1882_n2088# 0.018544f
C152 source.n29 a_n1882_n2088# 0.079767f
C153 source.n30 a_n1882_n2088# 0.053093f
C154 source.n31 a_n1882_n2088# 0.819449f
C155 source.t0 a_n1882_n2088# 0.163623f
C156 source.t38 a_n1882_n2088# 0.163623f
C157 source.n32 a_n1882_n2088# 1.27431f
C158 source.n33 a_n1882_n2088# 0.425107f
C159 source.t1 a_n1882_n2088# 0.163623f
C160 source.t15 a_n1882_n2088# 0.163623f
C161 source.n34 a_n1882_n2088# 1.27431f
C162 source.n35 a_n1882_n2088# 0.425107f
C163 source.t4 a_n1882_n2088# 0.163623f
C164 source.t39 a_n1882_n2088# 0.163623f
C165 source.n36 a_n1882_n2088# 1.27431f
C166 source.n37 a_n1882_n2088# 0.425107f
C167 source.t8 a_n1882_n2088# 0.163623f
C168 source.t3 a_n1882_n2088# 0.163623f
C169 source.n38 a_n1882_n2088# 1.27431f
C170 source.n39 a_n1882_n2088# 0.425107f
C171 source.n40 a_n1882_n2088# 0.048506f
C172 source.n41 a_n1882_n2088# 0.03451f
C173 source.n42 a_n1882_n2088# 0.018544f
C174 source.n43 a_n1882_n2088# 0.043831f
C175 source.n44 a_n1882_n2088# 0.019635f
C176 source.n45 a_n1882_n2088# 0.03451f
C177 source.n46 a_n1882_n2088# 0.018544f
C178 source.n47 a_n1882_n2088# 0.043831f
C179 source.n48 a_n1882_n2088# 0.019635f
C180 source.n49 a_n1882_n2088# 0.147677f
C181 source.t5 a_n1882_n2088# 0.071439f
C182 source.n50 a_n1882_n2088# 0.032873f
C183 source.n51 a_n1882_n2088# 0.025891f
C184 source.n52 a_n1882_n2088# 0.018544f
C185 source.n53 a_n1882_n2088# 0.821123f
C186 source.n54 a_n1882_n2088# 0.03451f
C187 source.n55 a_n1882_n2088# 0.018544f
C188 source.n56 a_n1882_n2088# 0.019635f
C189 source.n57 a_n1882_n2088# 0.043831f
C190 source.n58 a_n1882_n2088# 0.043831f
C191 source.n59 a_n1882_n2088# 0.019635f
C192 source.n60 a_n1882_n2088# 0.018544f
C193 source.n61 a_n1882_n2088# 0.03451f
C194 source.n62 a_n1882_n2088# 0.03451f
C195 source.n63 a_n1882_n2088# 0.018544f
C196 source.n64 a_n1882_n2088# 0.019635f
C197 source.n65 a_n1882_n2088# 0.043831f
C198 source.n66 a_n1882_n2088# 0.094887f
C199 source.n67 a_n1882_n2088# 0.019635f
C200 source.n68 a_n1882_n2088# 0.018544f
C201 source.n69 a_n1882_n2088# 0.079767f
C202 source.n70 a_n1882_n2088# 0.053093f
C203 source.n71 a_n1882_n2088# 0.132523f
C204 source.n72 a_n1882_n2088# 0.048506f
C205 source.n73 a_n1882_n2088# 0.03451f
C206 source.n74 a_n1882_n2088# 0.018544f
C207 source.n75 a_n1882_n2088# 0.043831f
C208 source.n76 a_n1882_n2088# 0.019635f
C209 source.n77 a_n1882_n2088# 0.03451f
C210 source.n78 a_n1882_n2088# 0.018544f
C211 source.n79 a_n1882_n2088# 0.043831f
C212 source.n80 a_n1882_n2088# 0.019635f
C213 source.n81 a_n1882_n2088# 0.147677f
C214 source.t28 a_n1882_n2088# 0.071439f
C215 source.n82 a_n1882_n2088# 0.032873f
C216 source.n83 a_n1882_n2088# 0.025891f
C217 source.n84 a_n1882_n2088# 0.018544f
C218 source.n85 a_n1882_n2088# 0.821123f
C219 source.n86 a_n1882_n2088# 0.03451f
C220 source.n87 a_n1882_n2088# 0.018544f
C221 source.n88 a_n1882_n2088# 0.019635f
C222 source.n89 a_n1882_n2088# 0.043831f
C223 source.n90 a_n1882_n2088# 0.043831f
C224 source.n91 a_n1882_n2088# 0.019635f
C225 source.n92 a_n1882_n2088# 0.018544f
C226 source.n93 a_n1882_n2088# 0.03451f
C227 source.n94 a_n1882_n2088# 0.03451f
C228 source.n95 a_n1882_n2088# 0.018544f
C229 source.n96 a_n1882_n2088# 0.019635f
C230 source.n97 a_n1882_n2088# 0.043831f
C231 source.n98 a_n1882_n2088# 0.094887f
C232 source.n99 a_n1882_n2088# 0.019635f
C233 source.n100 a_n1882_n2088# 0.018544f
C234 source.n101 a_n1882_n2088# 0.079767f
C235 source.n102 a_n1882_n2088# 0.053093f
C236 source.n103 a_n1882_n2088# 0.132523f
C237 source.t35 a_n1882_n2088# 0.163623f
C238 source.t31 a_n1882_n2088# 0.163623f
C239 source.n104 a_n1882_n2088# 1.27431f
C240 source.n105 a_n1882_n2088# 0.425107f
C241 source.t27 a_n1882_n2088# 0.163623f
C242 source.t24 a_n1882_n2088# 0.163623f
C243 source.n106 a_n1882_n2088# 1.27431f
C244 source.n107 a_n1882_n2088# 0.425107f
C245 source.t34 a_n1882_n2088# 0.163623f
C246 source.t32 a_n1882_n2088# 0.163623f
C247 source.n108 a_n1882_n2088# 1.27431f
C248 source.n109 a_n1882_n2088# 0.425107f
C249 source.t29 a_n1882_n2088# 0.163623f
C250 source.t23 a_n1882_n2088# 0.163623f
C251 source.n110 a_n1882_n2088# 1.27431f
C252 source.n111 a_n1882_n2088# 0.425107f
C253 source.n112 a_n1882_n2088# 0.048506f
C254 source.n113 a_n1882_n2088# 0.03451f
C255 source.n114 a_n1882_n2088# 0.018544f
C256 source.n115 a_n1882_n2088# 0.043831f
C257 source.n116 a_n1882_n2088# 0.019635f
C258 source.n117 a_n1882_n2088# 0.03451f
C259 source.n118 a_n1882_n2088# 0.018544f
C260 source.n119 a_n1882_n2088# 0.043831f
C261 source.n120 a_n1882_n2088# 0.019635f
C262 source.n121 a_n1882_n2088# 0.147677f
C263 source.t30 a_n1882_n2088# 0.071439f
C264 source.n122 a_n1882_n2088# 0.032873f
C265 source.n123 a_n1882_n2088# 0.025891f
C266 source.n124 a_n1882_n2088# 0.018544f
C267 source.n125 a_n1882_n2088# 0.821123f
C268 source.n126 a_n1882_n2088# 0.03451f
C269 source.n127 a_n1882_n2088# 0.018544f
C270 source.n128 a_n1882_n2088# 0.019635f
C271 source.n129 a_n1882_n2088# 0.043831f
C272 source.n130 a_n1882_n2088# 0.043831f
C273 source.n131 a_n1882_n2088# 0.019635f
C274 source.n132 a_n1882_n2088# 0.018544f
C275 source.n133 a_n1882_n2088# 0.03451f
C276 source.n134 a_n1882_n2088# 0.03451f
C277 source.n135 a_n1882_n2088# 0.018544f
C278 source.n136 a_n1882_n2088# 0.019635f
C279 source.n137 a_n1882_n2088# 0.043831f
C280 source.n138 a_n1882_n2088# 0.094887f
C281 source.n139 a_n1882_n2088# 0.019635f
C282 source.n140 a_n1882_n2088# 0.018544f
C283 source.n141 a_n1882_n2088# 0.079767f
C284 source.n142 a_n1882_n2088# 0.053093f
C285 source.n143 a_n1882_n2088# 1.261f
C286 source.n144 a_n1882_n2088# 0.048506f
C287 source.n145 a_n1882_n2088# 0.03451f
C288 source.n146 a_n1882_n2088# 0.018544f
C289 source.n147 a_n1882_n2088# 0.043831f
C290 source.n148 a_n1882_n2088# 0.019635f
C291 source.n149 a_n1882_n2088# 0.03451f
C292 source.n150 a_n1882_n2088# 0.018544f
C293 source.n151 a_n1882_n2088# 0.043831f
C294 source.n152 a_n1882_n2088# 0.019635f
C295 source.n153 a_n1882_n2088# 0.147677f
C296 source.t9 a_n1882_n2088# 0.071439f
C297 source.n154 a_n1882_n2088# 0.032873f
C298 source.n155 a_n1882_n2088# 0.025891f
C299 source.n156 a_n1882_n2088# 0.018544f
C300 source.n157 a_n1882_n2088# 0.821123f
C301 source.n158 a_n1882_n2088# 0.03451f
C302 source.n159 a_n1882_n2088# 0.018544f
C303 source.n160 a_n1882_n2088# 0.019635f
C304 source.n161 a_n1882_n2088# 0.043831f
C305 source.n162 a_n1882_n2088# 0.043831f
C306 source.n163 a_n1882_n2088# 0.019635f
C307 source.n164 a_n1882_n2088# 0.018544f
C308 source.n165 a_n1882_n2088# 0.03451f
C309 source.n166 a_n1882_n2088# 0.03451f
C310 source.n167 a_n1882_n2088# 0.018544f
C311 source.n168 a_n1882_n2088# 0.019635f
C312 source.n169 a_n1882_n2088# 0.043831f
C313 source.n170 a_n1882_n2088# 0.094887f
C314 source.n171 a_n1882_n2088# 0.019635f
C315 source.n172 a_n1882_n2088# 0.018544f
C316 source.n173 a_n1882_n2088# 0.079767f
C317 source.n174 a_n1882_n2088# 0.053093f
C318 source.n175 a_n1882_n2088# 1.261f
C319 source.t12 a_n1882_n2088# 0.163623f
C320 source.t11 a_n1882_n2088# 0.163623f
C321 source.n176 a_n1882_n2088# 1.2743f
C322 source.n177 a_n1882_n2088# 0.425115f
C323 source.t6 a_n1882_n2088# 0.163623f
C324 source.t16 a_n1882_n2088# 0.163623f
C325 source.n178 a_n1882_n2088# 1.2743f
C326 source.n179 a_n1882_n2088# 0.425115f
C327 source.t13 a_n1882_n2088# 0.163623f
C328 source.t17 a_n1882_n2088# 0.163623f
C329 source.n180 a_n1882_n2088# 1.2743f
C330 source.n181 a_n1882_n2088# 0.425115f
C331 source.t10 a_n1882_n2088# 0.163623f
C332 source.t7 a_n1882_n2088# 0.163623f
C333 source.n182 a_n1882_n2088# 1.2743f
C334 source.n183 a_n1882_n2088# 0.425115f
C335 source.n184 a_n1882_n2088# 0.048506f
C336 source.n185 a_n1882_n2088# 0.03451f
C337 source.n186 a_n1882_n2088# 0.018544f
C338 source.n187 a_n1882_n2088# 0.043831f
C339 source.n188 a_n1882_n2088# 0.019635f
C340 source.n189 a_n1882_n2088# 0.03451f
C341 source.n190 a_n1882_n2088# 0.018544f
C342 source.n191 a_n1882_n2088# 0.043831f
C343 source.n192 a_n1882_n2088# 0.019635f
C344 source.n193 a_n1882_n2088# 0.147677f
C345 source.t14 a_n1882_n2088# 0.071439f
C346 source.n194 a_n1882_n2088# 0.032873f
C347 source.n195 a_n1882_n2088# 0.025891f
C348 source.n196 a_n1882_n2088# 0.018544f
C349 source.n197 a_n1882_n2088# 0.821123f
C350 source.n198 a_n1882_n2088# 0.03451f
C351 source.n199 a_n1882_n2088# 0.018544f
C352 source.n200 a_n1882_n2088# 0.019635f
C353 source.n201 a_n1882_n2088# 0.043831f
C354 source.n202 a_n1882_n2088# 0.043831f
C355 source.n203 a_n1882_n2088# 0.019635f
C356 source.n204 a_n1882_n2088# 0.018544f
C357 source.n205 a_n1882_n2088# 0.03451f
C358 source.n206 a_n1882_n2088# 0.03451f
C359 source.n207 a_n1882_n2088# 0.018544f
C360 source.n208 a_n1882_n2088# 0.019635f
C361 source.n209 a_n1882_n2088# 0.043831f
C362 source.n210 a_n1882_n2088# 0.094887f
C363 source.n211 a_n1882_n2088# 0.019635f
C364 source.n212 a_n1882_n2088# 0.018544f
C365 source.n213 a_n1882_n2088# 0.079767f
C366 source.n214 a_n1882_n2088# 0.053093f
C367 source.n215 a_n1882_n2088# 0.132523f
C368 source.n216 a_n1882_n2088# 0.048506f
C369 source.n217 a_n1882_n2088# 0.03451f
C370 source.n218 a_n1882_n2088# 0.018544f
C371 source.n219 a_n1882_n2088# 0.043831f
C372 source.n220 a_n1882_n2088# 0.019635f
C373 source.n221 a_n1882_n2088# 0.03451f
C374 source.n222 a_n1882_n2088# 0.018544f
C375 source.n223 a_n1882_n2088# 0.043831f
C376 source.n224 a_n1882_n2088# 0.019635f
C377 source.n225 a_n1882_n2088# 0.147677f
C378 source.t25 a_n1882_n2088# 0.071439f
C379 source.n226 a_n1882_n2088# 0.032873f
C380 source.n227 a_n1882_n2088# 0.025891f
C381 source.n228 a_n1882_n2088# 0.018544f
C382 source.n229 a_n1882_n2088# 0.821123f
C383 source.n230 a_n1882_n2088# 0.03451f
C384 source.n231 a_n1882_n2088# 0.018544f
C385 source.n232 a_n1882_n2088# 0.019635f
C386 source.n233 a_n1882_n2088# 0.043831f
C387 source.n234 a_n1882_n2088# 0.043831f
C388 source.n235 a_n1882_n2088# 0.019635f
C389 source.n236 a_n1882_n2088# 0.018544f
C390 source.n237 a_n1882_n2088# 0.03451f
C391 source.n238 a_n1882_n2088# 0.03451f
C392 source.n239 a_n1882_n2088# 0.018544f
C393 source.n240 a_n1882_n2088# 0.019635f
C394 source.n241 a_n1882_n2088# 0.043831f
C395 source.n242 a_n1882_n2088# 0.094887f
C396 source.n243 a_n1882_n2088# 0.019635f
C397 source.n244 a_n1882_n2088# 0.018544f
C398 source.n245 a_n1882_n2088# 0.079767f
C399 source.n246 a_n1882_n2088# 0.053093f
C400 source.n247 a_n1882_n2088# 0.132523f
C401 source.t20 a_n1882_n2088# 0.163623f
C402 source.t26 a_n1882_n2088# 0.163623f
C403 source.n248 a_n1882_n2088# 1.2743f
C404 source.n249 a_n1882_n2088# 0.425115f
C405 source.t21 a_n1882_n2088# 0.163623f
C406 source.t33 a_n1882_n2088# 0.163623f
C407 source.n250 a_n1882_n2088# 1.2743f
C408 source.n251 a_n1882_n2088# 0.425115f
C409 source.t18 a_n1882_n2088# 0.163623f
C410 source.t36 a_n1882_n2088# 0.163623f
C411 source.n252 a_n1882_n2088# 1.2743f
C412 source.n253 a_n1882_n2088# 0.425115f
C413 source.t19 a_n1882_n2088# 0.163623f
C414 source.t37 a_n1882_n2088# 0.163623f
C415 source.n254 a_n1882_n2088# 1.2743f
C416 source.n255 a_n1882_n2088# 0.425115f
C417 source.n256 a_n1882_n2088# 0.048506f
C418 source.n257 a_n1882_n2088# 0.03451f
C419 source.n258 a_n1882_n2088# 0.018544f
C420 source.n259 a_n1882_n2088# 0.043831f
C421 source.n260 a_n1882_n2088# 0.019635f
C422 source.n261 a_n1882_n2088# 0.03451f
C423 source.n262 a_n1882_n2088# 0.018544f
C424 source.n263 a_n1882_n2088# 0.043831f
C425 source.n264 a_n1882_n2088# 0.019635f
C426 source.n265 a_n1882_n2088# 0.147677f
C427 source.t22 a_n1882_n2088# 0.071439f
C428 source.n266 a_n1882_n2088# 0.032873f
C429 source.n267 a_n1882_n2088# 0.025891f
C430 source.n268 a_n1882_n2088# 0.018544f
C431 source.n269 a_n1882_n2088# 0.821123f
C432 source.n270 a_n1882_n2088# 0.03451f
C433 source.n271 a_n1882_n2088# 0.018544f
C434 source.n272 a_n1882_n2088# 0.019635f
C435 source.n273 a_n1882_n2088# 0.043831f
C436 source.n274 a_n1882_n2088# 0.043831f
C437 source.n275 a_n1882_n2088# 0.019635f
C438 source.n276 a_n1882_n2088# 0.018544f
C439 source.n277 a_n1882_n2088# 0.03451f
C440 source.n278 a_n1882_n2088# 0.03451f
C441 source.n279 a_n1882_n2088# 0.018544f
C442 source.n280 a_n1882_n2088# 0.019635f
C443 source.n281 a_n1882_n2088# 0.043831f
C444 source.n282 a_n1882_n2088# 0.094887f
C445 source.n283 a_n1882_n2088# 0.019635f
C446 source.n284 a_n1882_n2088# 0.018544f
C447 source.n285 a_n1882_n2088# 0.079767f
C448 source.n286 a_n1882_n2088# 0.053093f
C449 source.n287 a_n1882_n2088# 0.319646f
C450 source.n288 a_n1882_n2088# 1.40744f
C451 drain_right.t13 a_n1882_n2088# 0.180414f
C452 drain_right.t17 a_n1882_n2088# 0.180414f
C453 drain_right.n0 a_n1882_n2088# 1.5076f
C454 drain_right.t1 a_n1882_n2088# 0.180414f
C455 drain_right.t4 a_n1882_n2088# 0.180414f
C456 drain_right.n1 a_n1882_n2088# 1.50465f
C457 drain_right.n2 a_n1882_n2088# 0.849538f
C458 drain_right.t15 a_n1882_n2088# 0.180414f
C459 drain_right.t0 a_n1882_n2088# 0.180414f
C460 drain_right.n3 a_n1882_n2088# 1.50465f
C461 drain_right.t7 a_n1882_n2088# 0.180414f
C462 drain_right.t6 a_n1882_n2088# 0.180414f
C463 drain_right.n4 a_n1882_n2088# 1.5076f
C464 drain_right.t5 a_n1882_n2088# 0.180414f
C465 drain_right.t10 a_n1882_n2088# 0.180414f
C466 drain_right.n5 a_n1882_n2088# 1.50465f
C467 drain_right.n6 a_n1882_n2088# 0.849538f
C468 drain_right.n7 a_n1882_n2088# 1.66489f
C469 drain_right.t19 a_n1882_n2088# 0.180414f
C470 drain_right.t2 a_n1882_n2088# 0.180414f
C471 drain_right.n8 a_n1882_n2088# 1.5076f
C472 drain_right.t14 a_n1882_n2088# 0.180414f
C473 drain_right.t18 a_n1882_n2088# 0.180414f
C474 drain_right.n9 a_n1882_n2088# 1.50466f
C475 drain_right.n10 a_n1882_n2088# 0.85412f
C476 drain_right.t9 a_n1882_n2088# 0.180414f
C477 drain_right.t3 a_n1882_n2088# 0.180414f
C478 drain_right.n11 a_n1882_n2088# 1.50466f
C479 drain_right.n12 a_n1882_n2088# 0.420866f
C480 drain_right.t8 a_n1882_n2088# 0.180414f
C481 drain_right.t16 a_n1882_n2088# 0.180414f
C482 drain_right.n13 a_n1882_n2088# 1.50466f
C483 drain_right.n14 a_n1882_n2088# 0.420866f
C484 drain_right.t11 a_n1882_n2088# 0.180414f
C485 drain_right.t12 a_n1882_n2088# 0.180414f
C486 drain_right.n15 a_n1882_n2088# 1.50466f
C487 drain_right.n16 a_n1882_n2088# 0.732277f
C488 minus.n0 a_n1882_n2088# 0.052653f
C489 minus.t7 a_n1882_n2088# 0.185475f
C490 minus.t8 a_n1882_n2088# 0.180019f
C491 minus.t14 a_n1882_n2088# 0.180019f
C492 minus.t3 a_n1882_n2088# 0.180019f
C493 minus.n1 a_n1882_n2088# 0.088042f
C494 minus.n2 a_n1882_n2088# 0.052653f
C495 minus.t5 a_n1882_n2088# 0.180019f
C496 minus.t10 a_n1882_n2088# 0.180019f
C497 minus.t13 a_n1882_n2088# 0.180019f
C498 minus.n3 a_n1882_n2088# 0.088042f
C499 minus.n4 a_n1882_n2088# 0.120483f
C500 minus.t2 a_n1882_n2088# 0.180019f
C501 minus.t6 a_n1882_n2088# 0.180019f
C502 minus.t9 a_n1882_n2088# 0.185475f
C503 minus.n5 a_n1882_n2088# 0.103866f
C504 minus.n6 a_n1882_n2088# 0.088042f
C505 minus.n7 a_n1882_n2088# 0.01844f
C506 minus.n8 a_n1882_n2088# 0.088042f
C507 minus.n9 a_n1882_n2088# 0.01844f
C508 minus.n10 a_n1882_n2088# 0.052653f
C509 minus.n11 a_n1882_n2088# 0.052653f
C510 minus.n12 a_n1882_n2088# 0.01844f
C511 minus.n13 a_n1882_n2088# 0.088042f
C512 minus.n14 a_n1882_n2088# 0.01844f
C513 minus.n15 a_n1882_n2088# 0.088042f
C514 minus.n16 a_n1882_n2088# 0.01844f
C515 minus.n17 a_n1882_n2088# 0.052653f
C516 minus.n18 a_n1882_n2088# 0.052653f
C517 minus.n19 a_n1882_n2088# 0.01844f
C518 minus.n20 a_n1882_n2088# 0.088042f
C519 minus.n21 a_n1882_n2088# 0.01844f
C520 minus.n22 a_n1882_n2088# 0.088042f
C521 minus.n23 a_n1882_n2088# 0.103786f
C522 minus.n24 a_n1882_n2088# 1.50053f
C523 minus.n25 a_n1882_n2088# 0.052653f
C524 minus.t0 a_n1882_n2088# 0.180019f
C525 minus.t18 a_n1882_n2088# 0.180019f
C526 minus.t1 a_n1882_n2088# 0.180019f
C527 minus.n26 a_n1882_n2088# 0.088042f
C528 minus.n27 a_n1882_n2088# 0.052653f
C529 minus.t19 a_n1882_n2088# 0.180019f
C530 minus.t4 a_n1882_n2088# 0.180019f
C531 minus.t16 a_n1882_n2088# 0.180019f
C532 minus.n28 a_n1882_n2088# 0.088042f
C533 minus.n29 a_n1882_n2088# 0.120483f
C534 minus.t11 a_n1882_n2088# 0.180019f
C535 minus.t17 a_n1882_n2088# 0.180019f
C536 minus.t12 a_n1882_n2088# 0.185475f
C537 minus.n30 a_n1882_n2088# 0.103866f
C538 minus.n31 a_n1882_n2088# 0.088042f
C539 minus.n32 a_n1882_n2088# 0.01844f
C540 minus.n33 a_n1882_n2088# 0.088042f
C541 minus.n34 a_n1882_n2088# 0.01844f
C542 minus.n35 a_n1882_n2088# 0.052653f
C543 minus.n36 a_n1882_n2088# 0.052653f
C544 minus.n37 a_n1882_n2088# 0.01844f
C545 minus.n38 a_n1882_n2088# 0.088042f
C546 minus.n39 a_n1882_n2088# 0.01844f
C547 minus.n40 a_n1882_n2088# 0.088042f
C548 minus.n41 a_n1882_n2088# 0.01844f
C549 minus.n42 a_n1882_n2088# 0.052653f
C550 minus.n43 a_n1882_n2088# 0.052653f
C551 minus.n44 a_n1882_n2088# 0.01844f
C552 minus.n45 a_n1882_n2088# 0.088042f
C553 minus.n46 a_n1882_n2088# 0.01844f
C554 minus.n47 a_n1882_n2088# 0.088042f
C555 minus.t15 a_n1882_n2088# 0.185475f
C556 minus.n48 a_n1882_n2088# 0.103786f
C557 minus.n49 a_n1882_n2088# 0.341468f
C558 minus.n50 a_n1882_n2088# 1.84627f
.ends

