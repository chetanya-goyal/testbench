* NGSPICE file created from diffpair63.ext - technology: sky130A

.subckt diffpair63 minus drain_right drain_left source plus
X0 a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X1 source.t15 plus.t0 drain_left.t4 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X2 source.t5 minus.t0 drain_right.t7 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X3 source.t14 plus.t1 drain_left.t2 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X4 drain_right.t6 minus.t1 source.t2 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X5 source.t3 minus.t2 drain_right.t5 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X6 a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X7 drain_right.t4 minus.t3 source.t4 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X8 source.t1 minus.t4 drain_right.t3 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X9 source.t13 plus.t2 drain_left.t1 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X10 drain_right.t2 minus.t5 source.t6 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X11 drain_left.t0 plus.t3 source.t12 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X12 drain_left.t5 plus.t4 source.t11 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X13 drain_right.t1 minus.t6 source.t7 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X14 drain_left.t7 plus.t5 source.t10 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X15 a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X16 drain_left.t6 plus.t6 source.t9 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X17 a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X18 source.t0 minus.t7 drain_right.t0 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X19 source.t8 plus.t7 drain_left.t3 a_n1746_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n5 plus.n4 161.3
R1 plus.n6 plus.n1 161.3
R2 plus.n7 plus.n0 161.3
R3 plus.n9 plus.n8 161.3
R4 plus.n15 plus.n14 161.3
R5 plus.n16 plus.n11 161.3
R6 plus.n17 plus.n10 161.3
R7 plus.n19 plus.n18 161.3
R8 plus.n3 plus.t1 112.725
R9 plus.n13 plus.t3 112.725
R10 plus.n8 plus.t4 90.5476
R11 plus.n6 plus.t0 90.5476
R12 plus.n2 plus.t5 90.5476
R13 plus.n18 plus.t7 90.5476
R14 plus.n16 plus.t6 90.5476
R15 plus.n12 plus.t2 90.5476
R16 plus.n4 plus.n3 44.862
R17 plus.n14 plus.n13 44.862
R18 plus.n8 plus.n7 28.4823
R19 plus.n18 plus.n17 28.4823
R20 plus plus.n19 25.5824
R21 plus.n5 plus.n2 24.1005
R22 plus.n6 plus.n5 24.1005
R23 plus.n16 plus.n15 24.1005
R24 plus.n15 plus.n12 24.1005
R25 plus.n7 plus.n6 19.7187
R26 plus.n17 plus.n16 19.7187
R27 plus.n3 plus.n2 19.7081
R28 plus.n13 plus.n12 19.7081
R29 plus plus.n9 8.11035
R30 plus.n4 plus.n1 0.189894
R31 plus.n1 plus.n0 0.189894
R32 plus.n9 plus.n0 0.189894
R33 plus.n19 plus.n10 0.189894
R34 plus.n11 plus.n10 0.189894
R35 plus.n14 plus.n11 0.189894
R36 drain_left.n5 drain_left.n3 241.02
R37 drain_left.n2 drain_left.n1 240.52
R38 drain_left.n2 drain_left.n0 240.52
R39 drain_left.n5 drain_left.n4 240.132
R40 drain_left drain_left.n2 22.1415
R41 drain_left.n1 drain_left.t1 19.8005
R42 drain_left.n1 drain_left.t0 19.8005
R43 drain_left.n0 drain_left.t3 19.8005
R44 drain_left.n0 drain_left.t6 19.8005
R45 drain_left.n4 drain_left.t4 19.8005
R46 drain_left.n4 drain_left.t5 19.8005
R47 drain_left.n3 drain_left.t2 19.8005
R48 drain_left.n3 drain_left.t7 19.8005
R49 drain_left drain_left.n5 6.54115
R50 source.n0 source.t11 243.255
R51 source.n3 source.t14 243.255
R52 source.n4 source.t7 243.255
R53 source.n7 source.t0 243.255
R54 source.n15 source.t4 243.254
R55 source.n12 source.t3 243.254
R56 source.n11 source.t12 243.254
R57 source.n8 source.t8 243.254
R58 source.n2 source.n1 223.454
R59 source.n6 source.n5 223.454
R60 source.n14 source.n13 223.453
R61 source.n10 source.n9 223.453
R62 source.n13 source.t2 19.8005
R63 source.n13 source.t1 19.8005
R64 source.n9 source.t9 19.8005
R65 source.n9 source.t13 19.8005
R66 source.n1 source.t10 19.8005
R67 source.n1 source.t15 19.8005
R68 source.n5 source.t6 19.8005
R69 source.n5 source.t5 19.8005
R70 source.n8 source.n7 13.8423
R71 source.n16 source.n0 8.13543
R72 source.n16 source.n15 5.7074
R73 source.n7 source.n6 0.888431
R74 source.n6 source.n4 0.888431
R75 source.n3 source.n2 0.888431
R76 source.n2 source.n0 0.888431
R77 source.n10 source.n8 0.888431
R78 source.n11 source.n10 0.888431
R79 source.n14 source.n12 0.888431
R80 source.n15 source.n14 0.888431
R81 source.n4 source.n3 0.470328
R82 source.n12 source.n11 0.470328
R83 source source.n16 0.188
R84 minus.n9 minus.n8 161.3
R85 minus.n7 minus.n0 161.3
R86 minus.n6 minus.n5 161.3
R87 minus.n4 minus.n1 161.3
R88 minus.n19 minus.n18 161.3
R89 minus.n17 minus.n10 161.3
R90 minus.n16 minus.n15 161.3
R91 minus.n14 minus.n11 161.3
R92 minus.n3 minus.t6 112.725
R93 minus.n13 minus.t2 112.725
R94 minus.n2 minus.t0 90.5476
R95 minus.n6 minus.t5 90.5476
R96 minus.n8 minus.t7 90.5476
R97 minus.n12 minus.t1 90.5476
R98 minus.n16 minus.t4 90.5476
R99 minus.n18 minus.t3 90.5476
R100 minus.n4 minus.n3 44.862
R101 minus.n14 minus.n13 44.862
R102 minus.n8 minus.n7 28.4823
R103 minus.n18 minus.n17 28.4823
R104 minus.n20 minus.n9 27.5346
R105 minus.n6 minus.n1 24.1005
R106 minus.n2 minus.n1 24.1005
R107 minus.n12 minus.n11 24.1005
R108 minus.n16 minus.n11 24.1005
R109 minus.n7 minus.n6 19.7187
R110 minus.n17 minus.n16 19.7187
R111 minus.n3 minus.n2 19.7081
R112 minus.n13 minus.n12 19.7081
R113 minus.n20 minus.n19 6.63308
R114 minus.n9 minus.n0 0.189894
R115 minus.n5 minus.n0 0.189894
R116 minus.n5 minus.n4 0.189894
R117 minus.n15 minus.n14 0.189894
R118 minus.n15 minus.n10 0.189894
R119 minus.n19 minus.n10 0.189894
R120 minus minus.n20 0.188
R121 drain_right.n5 drain_right.n3 241.02
R122 drain_right.n2 drain_right.n1 240.52
R123 drain_right.n2 drain_right.n0 240.52
R124 drain_right.n5 drain_right.n4 240.132
R125 drain_right drain_right.n2 21.5883
R126 drain_right.n1 drain_right.t3 19.8005
R127 drain_right.n1 drain_right.t4 19.8005
R128 drain_right.n0 drain_right.t5 19.8005
R129 drain_right.n0 drain_right.t6 19.8005
R130 drain_right.n3 drain_right.t7 19.8005
R131 drain_right.n3 drain_right.t1 19.8005
R132 drain_right.n4 drain_right.t0 19.8005
R133 drain_right.n4 drain_right.t2 19.8005
R134 drain_right drain_right.n5 6.54115
C0 source minus 1.18365f
C1 drain_left source 2.92415f
C2 drain_right source 2.9259f
C3 drain_left minus 0.178127f
C4 source plus 1.19752f
C5 drain_right minus 0.827094f
C6 drain_left drain_right 0.821863f
C7 plus minus 3.29156f
C8 drain_left plus 0.995868f
C9 drain_right plus 0.331171f
C10 drain_right a_n1746_n1088# 3.128152f
C11 drain_left a_n1746_n1088# 3.340498f
C12 source a_n1746_n1088# 2.434475f
C13 minus a_n1746_n1088# 5.847984f
C14 plus a_n1746_n1088# 6.480966f
C15 drain_right.t5 a_n1746_n1088# 0.01531f
C16 drain_right.t6 a_n1746_n1088# 0.01531f
C17 drain_right.n0 a_n1746_n1088# 0.059853f
C18 drain_right.t3 a_n1746_n1088# 0.01531f
C19 drain_right.t4 a_n1746_n1088# 0.01531f
C20 drain_right.n1 a_n1746_n1088# 0.059853f
C21 drain_right.n2 a_n1746_n1088# 0.930863f
C22 drain_right.t7 a_n1746_n1088# 0.01531f
C23 drain_right.t1 a_n1746_n1088# 0.01531f
C24 drain_right.n3 a_n1746_n1088# 0.060427f
C25 drain_right.t0 a_n1746_n1088# 0.01531f
C26 drain_right.t2 a_n1746_n1088# 0.01531f
C27 drain_right.n4 a_n1746_n1088# 0.059491f
C28 drain_right.n5 a_n1746_n1088# 0.670938f
C29 minus.n0 a_n1746_n1088# 0.030265f
C30 minus.n1 a_n1746_n1088# 0.006868f
C31 minus.t5 a_n1746_n1088# 0.071839f
C32 minus.t6 a_n1746_n1088# 0.08586f
C33 minus.t0 a_n1746_n1088# 0.071839f
C34 minus.n2 a_n1746_n1088# 0.074157f
C35 minus.n3 a_n1746_n1088# 0.060183f
C36 minus.n4 a_n1746_n1088# 0.125856f
C37 minus.n5 a_n1746_n1088# 0.030265f
C38 minus.n6 a_n1746_n1088# 0.071419f
C39 minus.n7 a_n1746_n1088# 0.006868f
C40 minus.t7 a_n1746_n1088# 0.071839f
C41 minus.n8 a_n1746_n1088# 0.069459f
C42 minus.n9 a_n1746_n1088# 0.6819f
C43 minus.n10 a_n1746_n1088# 0.030265f
C44 minus.n11 a_n1746_n1088# 0.006868f
C45 minus.t2 a_n1746_n1088# 0.08586f
C46 minus.t1 a_n1746_n1088# 0.071839f
C47 minus.n12 a_n1746_n1088# 0.074157f
C48 minus.n13 a_n1746_n1088# 0.060183f
C49 minus.n14 a_n1746_n1088# 0.125856f
C50 minus.n15 a_n1746_n1088# 0.030265f
C51 minus.t4 a_n1746_n1088# 0.071839f
C52 minus.n16 a_n1746_n1088# 0.071419f
C53 minus.n17 a_n1746_n1088# 0.006868f
C54 minus.t3 a_n1746_n1088# 0.071839f
C55 minus.n18 a_n1746_n1088# 0.069459f
C56 minus.n19 a_n1746_n1088# 0.207293f
C57 minus.n20 a_n1746_n1088# 0.837497f
C58 source.t11 a_n1746_n1088# 0.097576f
C59 source.n0 a_n1746_n1088# 0.462996f
C60 source.t10 a_n1746_n1088# 0.017531f
C61 source.t15 a_n1746_n1088# 0.017531f
C62 source.n1 a_n1746_n1088# 0.056856f
C63 source.n2 a_n1746_n1088# 0.263199f
C64 source.t14 a_n1746_n1088# 0.097576f
C65 source.n3 a_n1746_n1088# 0.240404f
C66 source.t7 a_n1746_n1088# 0.097576f
C67 source.n4 a_n1746_n1088# 0.240404f
C68 source.t6 a_n1746_n1088# 0.017531f
C69 source.t5 a_n1746_n1088# 0.017531f
C70 source.n5 a_n1746_n1088# 0.056856f
C71 source.n6 a_n1746_n1088# 0.263199f
C72 source.t0 a_n1746_n1088# 0.097576f
C73 source.n7 a_n1746_n1088# 0.646044f
C74 source.t8 a_n1746_n1088# 0.097576f
C75 source.n8 a_n1746_n1088# 0.646044f
C76 source.t9 a_n1746_n1088# 0.017531f
C77 source.t13 a_n1746_n1088# 0.017531f
C78 source.n9 a_n1746_n1088# 0.056856f
C79 source.n10 a_n1746_n1088# 0.263199f
C80 source.t12 a_n1746_n1088# 0.097576f
C81 source.n11 a_n1746_n1088# 0.240404f
C82 source.t3 a_n1746_n1088# 0.097576f
C83 source.n12 a_n1746_n1088# 0.240404f
C84 source.t2 a_n1746_n1088# 0.017531f
C85 source.t1 a_n1746_n1088# 0.017531f
C86 source.n13 a_n1746_n1088# 0.056856f
C87 source.n14 a_n1746_n1088# 0.263199f
C88 source.t4 a_n1746_n1088# 0.097576f
C89 source.n15 a_n1746_n1088# 0.385117f
C90 source.n16 a_n1746_n1088# 0.459755f
C91 drain_left.t3 a_n1746_n1088# 0.01492f
C92 drain_left.t6 a_n1746_n1088# 0.01492f
C93 drain_left.n0 a_n1746_n1088# 0.058329f
C94 drain_left.t1 a_n1746_n1088# 0.01492f
C95 drain_left.t0 a_n1746_n1088# 0.01492f
C96 drain_left.n1 a_n1746_n1088# 0.058329f
C97 drain_left.n2 a_n1746_n1088# 0.943678f
C98 drain_left.t2 a_n1746_n1088# 0.01492f
C99 drain_left.t7 a_n1746_n1088# 0.01492f
C100 drain_left.n3 a_n1746_n1088# 0.058888f
C101 drain_left.t4 a_n1746_n1088# 0.01492f
C102 drain_left.t5 a_n1746_n1088# 0.01492f
C103 drain_left.n4 a_n1746_n1088# 0.057976f
C104 drain_left.n5 a_n1746_n1088# 0.65385f
C105 plus.n0 a_n1746_n1088# 0.030837f
C106 plus.t4 a_n1746_n1088# 0.073197f
C107 plus.t0 a_n1746_n1088# 0.073197f
C108 plus.n1 a_n1746_n1088# 0.030837f
C109 plus.t5 a_n1746_n1088# 0.073197f
C110 plus.n2 a_n1746_n1088# 0.075559f
C111 plus.t1 a_n1746_n1088# 0.087482f
C112 plus.n3 a_n1746_n1088# 0.06132f
C113 plus.n4 a_n1746_n1088# 0.128234f
C114 plus.n5 a_n1746_n1088# 0.006997f
C115 plus.n6 a_n1746_n1088# 0.072768f
C116 plus.n7 a_n1746_n1088# 0.006997f
C117 plus.n8 a_n1746_n1088# 0.070772f
C118 plus.n9 a_n1746_n1088# 0.221547f
C119 plus.n10 a_n1746_n1088# 0.030837f
C120 plus.t7 a_n1746_n1088# 0.073197f
C121 plus.n11 a_n1746_n1088# 0.030837f
C122 plus.t6 a_n1746_n1088# 0.073197f
C123 plus.t2 a_n1746_n1088# 0.073197f
C124 plus.n12 a_n1746_n1088# 0.075559f
C125 plus.t3 a_n1746_n1088# 0.087482f
C126 plus.n13 a_n1746_n1088# 0.06132f
C127 plus.n14 a_n1746_n1088# 0.128234f
C128 plus.n15 a_n1746_n1088# 0.006997f
C129 plus.n16 a_n1746_n1088# 0.072768f
C130 plus.n17 a_n1746_n1088# 0.006997f
C131 plus.n18 a_n1746_n1088# 0.070772f
C132 plus.n19 a_n1746_n1088# 0.674757f
.ends

