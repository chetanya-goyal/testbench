* NGSPICE file created from diffpair485.ext - technology: sky130A

.subckt diffpair485 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t12 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X1 a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X2 source.t18 minus.t1 drain_right.t10 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X3 source.t11 plus.t0 drain_left.t11 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X4 a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X5 a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X6 drain_left.t10 plus.t1 source.t6 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X7 source.t22 minus.t2 drain_right.t9 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X8 drain_right.t8 minus.t3 source.t21 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X9 drain_right.t7 minus.t4 source.t20 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X10 source.t3 plus.t2 drain_left.t9 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X11 source.t16 minus.t5 drain_right.t6 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X12 source.t17 minus.t6 drain_right.t5 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X13 source.t4 plus.t3 drain_left.t8 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X14 drain_right.t4 minus.t7 source.t23 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X15 drain_left.t7 plus.t4 source.t7 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X16 drain_left.t6 plus.t5 source.t8 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X17 source.t13 minus.t8 drain_right.t3 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X18 drain_right.t2 minus.t9 source.t14 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X19 drain_left.t5 plus.t6 source.t0 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X20 source.t10 plus.t7 drain_left.t4 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X21 drain_right.t1 minus.t10 source.t15 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X22 drain_left.t3 plus.t8 source.t2 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X23 drain_left.t2 plus.t9 source.t1 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X24 source.t5 plus.t10 drain_left.t1 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X25 a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X26 source.t9 plus.t11 drain_left.t0 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X27 source.t19 minus.t11 drain_right.t0 a_n1626_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
R0 minus.n13 minus.t8 2673.64
R1 minus.n2 minus.t3 2673.64
R2 minus.n28 minus.t10 2673.64
R3 minus.n17 minus.t1 2673.64
R4 minus.n12 minus.t4 2618.87
R5 minus.n10 minus.t5 2618.87
R6 minus.n3 minus.t7 2618.87
R7 minus.n4 minus.t2 2618.87
R8 minus.n27 minus.t6 2618.87
R9 minus.n25 minus.t0 2618.87
R10 minus.n19 minus.t11 2618.87
R11 minus.n18 minus.t9 2618.87
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 62.0763
R27 minus.n5 minus.n3 62.0763
R28 minus.n20 minus.n19 62.0763
R29 minus.n26 minus.n25 62.0763
R30 minus.n13 minus.n12 40.1672
R31 minus.n4 minus.n2 40.1672
R32 minus.n18 minus.n17 40.1672
R33 minus.n28 minus.n27 40.1672
R34 minus.n30 minus.n14 37.5952
R35 minus.n12 minus.n11 32.8641
R36 minus.n5 minus.n4 32.8641
R37 minus.n20 minus.n18 32.8641
R38 minus.n27 minus.n26 32.8641
R39 minus.n10 minus.n9 10.955
R40 minus.n3 minus.n1 10.955
R41 minus.n19 minus.n16 10.955
R42 minus.n25 minus.n24 10.955
R43 minus.n30 minus.n29 6.54217
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 source.n5 source.t4 46.201
R54 source.n6 source.t21 46.201
R55 source.n11 source.t13 46.201
R56 source.n23 source.t15 46.2008
R57 source.n18 source.t18 46.2008
R58 source.n17 source.t7 46.2008
R59 source.n12 source.t11 46.2008
R60 source.n0 source.t2 46.2008
R61 source.n2 source.n1 44.201
R62 source.n4 source.n3 44.201
R63 source.n8 source.n7 44.201
R64 source.n10 source.n9 44.201
R65 source.n22 source.n21 44.2008
R66 source.n20 source.n19 44.2008
R67 source.n16 source.n15 44.2008
R68 source.n14 source.n13 44.2008
R69 source.n12 source.n11 24.1208
R70 source.n24 source.n0 18.5777
R71 source.n24 source.n23 5.5436
R72 source.n21 source.t12 2.0005
R73 source.n21 source.t17 2.0005
R74 source.n19 source.t14 2.0005
R75 source.n19 source.t19 2.0005
R76 source.n15 source.t6 2.0005
R77 source.n15 source.t5 2.0005
R78 source.n13 source.t0 2.0005
R79 source.n13 source.t3 2.0005
R80 source.n1 source.t8 2.0005
R81 source.n1 source.t9 2.0005
R82 source.n3 source.t1 2.0005
R83 source.n3 source.t10 2.0005
R84 source.n7 source.t23 2.0005
R85 source.n7 source.t22 2.0005
R86 source.n9 source.t20 2.0005
R87 source.n9 source.t16 2.0005
R88 source.n11 source.n10 0.560845
R89 source.n10 source.n8 0.560845
R90 source.n8 source.n6 0.560845
R91 source.n5 source.n4 0.560845
R92 source.n4 source.n2 0.560845
R93 source.n2 source.n0 0.560845
R94 source.n14 source.n12 0.560845
R95 source.n16 source.n14 0.560845
R96 source.n17 source.n16 0.560845
R97 source.n20 source.n18 0.560845
R98 source.n22 source.n20 0.560845
R99 source.n23 source.n22 0.560845
R100 source.n6 source.n5 0.470328
R101 source.n18 source.n17 0.470328
R102 source source.n24 0.188
R103 drain_right.n6 drain_right.n4 61.44
R104 drain_right.n3 drain_right.n2 61.3846
R105 drain_right.n3 drain_right.n0 61.3846
R106 drain_right.n6 drain_right.n5 60.8798
R107 drain_right.n8 drain_right.n7 60.8798
R108 drain_right.n3 drain_right.n1 60.8796
R109 drain_right drain_right.n3 31.8883
R110 drain_right drain_right.n8 6.21356
R111 drain_right.n1 drain_right.t0 2.0005
R112 drain_right.n1 drain_right.t11 2.0005
R113 drain_right.n2 drain_right.t5 2.0005
R114 drain_right.n2 drain_right.t1 2.0005
R115 drain_right.n0 drain_right.t10 2.0005
R116 drain_right.n0 drain_right.t2 2.0005
R117 drain_right.n4 drain_right.t9 2.0005
R118 drain_right.n4 drain_right.t8 2.0005
R119 drain_right.n5 drain_right.t6 2.0005
R120 drain_right.n5 drain_right.t4 2.0005
R121 drain_right.n7 drain_right.t3 2.0005
R122 drain_right.n7 drain_right.t7 2.0005
R123 drain_right.n8 drain_right.n6 0.560845
R124 plus.n2 plus.t3 2673.64
R125 plus.n13 plus.t8 2673.64
R126 plus.n17 plus.t4 2673.64
R127 plus.n28 plus.t0 2673.64
R128 plus.n3 plus.t9 2618.87
R129 plus.n4 plus.t7 2618.87
R130 plus.n10 plus.t5 2618.87
R131 plus.n12 plus.t11 2618.87
R132 plus.n19 plus.t10 2618.87
R133 plus.n18 plus.t1 2618.87
R134 plus.n25 plus.t2 2618.87
R135 plus.n27 plus.t6 2618.87
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 62.0763
R151 plus.n11 plus.n10 62.0763
R152 plus.n26 plus.n25 62.0763
R153 plus.n20 plus.n18 62.0763
R154 plus.n3 plus.n2 40.1672
R155 plus.n13 plus.n12 40.1672
R156 plus.n28 plus.n27 40.1672
R157 plus.n19 plus.n17 40.1672
R158 plus.n5 plus.n3 32.8641
R159 plus.n12 plus.n11 32.8641
R160 plus.n27 plus.n26 32.8641
R161 plus.n20 plus.n19 32.8641
R162 plus plus.n29 30.3399
R163 plus plus.n14 13.3225
R164 plus.n4 plus.n1 10.955
R165 plus.n10 plus.n9 10.955
R166 plus.n25 plus.n24 10.955
R167 plus.n18 plus.n16 10.955
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 61.4402
R177 drain_left.n3 drain_left.n2 61.3846
R178 drain_left.n3 drain_left.n0 61.3846
R179 drain_left.n6 drain_left.n5 60.8798
R180 drain_left.n8 drain_left.n7 60.8796
R181 drain_left.n3 drain_left.n1 60.8796
R182 drain_left drain_left.n3 32.4415
R183 drain_left drain_left.n8 6.21356
R184 drain_left.n1 drain_left.t9 2.0005
R185 drain_left.n1 drain_left.t10 2.0005
R186 drain_left.n2 drain_left.t1 2.0005
R187 drain_left.n2 drain_left.t7 2.0005
R188 drain_left.n0 drain_left.t11 2.0005
R189 drain_left.n0 drain_left.t5 2.0005
R190 drain_left.n7 drain_left.t0 2.0005
R191 drain_left.n7 drain_left.t3 2.0005
R192 drain_left.n5 drain_left.t4 2.0005
R193 drain_left.n5 drain_left.t6 2.0005
R194 drain_left.n4 drain_left.t8 2.0005
R195 drain_left.n4 drain_left.t2 2.0005
R196 drain_left.n8 drain_left.n6 0.560845
C0 minus drain_right 3.46892f
C1 plus drain_right 0.309819f
C2 source drain_left 29.428001f
C3 minus plus 5.71929f
C4 source drain_right 29.427801f
C5 source minus 2.79521f
C6 source plus 2.80925f
C7 drain_right drain_left 0.801529f
C8 minus drain_left 0.170585f
C9 plus drain_left 3.62541f
C10 drain_right a_n1626_n3888# 6.26695f
C11 drain_left a_n1626_n3888# 6.50892f
C12 source a_n1626_n3888# 10.312191f
C13 minus a_n1626_n3888# 6.183053f
C14 plus a_n1626_n3888# 8.561231f
C15 drain_left.t11 a_n1626_n3888# 0.505668f
C16 drain_left.t5 a_n1626_n3888# 0.505668f
C17 drain_left.n0 a_n1626_n3888# 3.36328f
C18 drain_left.t9 a_n1626_n3888# 0.505668f
C19 drain_left.t10 a_n1626_n3888# 0.505668f
C20 drain_left.n1 a_n1626_n3888# 3.36048f
C21 drain_left.t1 a_n1626_n3888# 0.505668f
C22 drain_left.t7 a_n1626_n3888# 0.505668f
C23 drain_left.n2 a_n1626_n3888# 3.36328f
C24 drain_left.n3 a_n1626_n3888# 2.47538f
C25 drain_left.t8 a_n1626_n3888# 0.505668f
C26 drain_left.t2 a_n1626_n3888# 0.505668f
C27 drain_left.n4 a_n1626_n3888# 3.36362f
C28 drain_left.t4 a_n1626_n3888# 0.505668f
C29 drain_left.t6 a_n1626_n3888# 0.505668f
C30 drain_left.n5 a_n1626_n3888# 3.36049f
C31 drain_left.n6 a_n1626_n3888# 0.672771f
C32 drain_left.t0 a_n1626_n3888# 0.505668f
C33 drain_left.t3 a_n1626_n3888# 0.505668f
C34 drain_left.n7 a_n1626_n3888# 3.36048f
C35 drain_left.n8 a_n1626_n3888# 0.567422f
C36 plus.n0 a_n1626_n3888# 0.057378f
C37 plus.t11 a_n1626_n3888# 0.364214f
C38 plus.t5 a_n1626_n3888# 0.364214f
C39 plus.n1 a_n1626_n3888# 0.021688f
C40 plus.t3 a_n1626_n3888# 0.36728f
C41 plus.n2 a_n1626_n3888# 0.170985f
C42 plus.t9 a_n1626_n3888# 0.364214f
C43 plus.n3 a_n1626_n3888# 0.148741f
C44 plus.t7 a_n1626_n3888# 0.364214f
C45 plus.n4 a_n1626_n3888# 0.148741f
C46 plus.n5 a_n1626_n3888# 0.024341f
C47 plus.n6 a_n1626_n3888# 0.128823f
C48 plus.n7 a_n1626_n3888# 0.057378f
C49 plus.n8 a_n1626_n3888# 0.057378f
C50 plus.n9 a_n1626_n3888# 0.021688f
C51 plus.n10 a_n1626_n3888# 0.148741f
C52 plus.n11 a_n1626_n3888# 0.024341f
C53 plus.n12 a_n1626_n3888# 0.148741f
C54 plus.t8 a_n1626_n3888# 0.36728f
C55 plus.n13 a_n1626_n3888# 0.170901f
C56 plus.n14 a_n1626_n3888# 0.730775f
C57 plus.n15 a_n1626_n3888# 0.057378f
C58 plus.t0 a_n1626_n3888# 0.36728f
C59 plus.t6 a_n1626_n3888# 0.364214f
C60 plus.t2 a_n1626_n3888# 0.364214f
C61 plus.n16 a_n1626_n3888# 0.021688f
C62 plus.t4 a_n1626_n3888# 0.36728f
C63 plus.n17 a_n1626_n3888# 0.170985f
C64 plus.t1 a_n1626_n3888# 0.364214f
C65 plus.n18 a_n1626_n3888# 0.148741f
C66 plus.t10 a_n1626_n3888# 0.364214f
C67 plus.n19 a_n1626_n3888# 0.148741f
C68 plus.n20 a_n1626_n3888# 0.024341f
C69 plus.n21 a_n1626_n3888# 0.128823f
C70 plus.n22 a_n1626_n3888# 0.057378f
C71 plus.n23 a_n1626_n3888# 0.057378f
C72 plus.n24 a_n1626_n3888# 0.021688f
C73 plus.n25 a_n1626_n3888# 0.148741f
C74 plus.n26 a_n1626_n3888# 0.024341f
C75 plus.n27 a_n1626_n3888# 0.148741f
C76 plus.n28 a_n1626_n3888# 0.170901f
C77 plus.n29 a_n1626_n3888# 1.76786f
C78 drain_right.t10 a_n1626_n3888# 0.505824f
C79 drain_right.t2 a_n1626_n3888# 0.505824f
C80 drain_right.n0 a_n1626_n3888# 3.36432f
C81 drain_right.t0 a_n1626_n3888# 0.505824f
C82 drain_right.t11 a_n1626_n3888# 0.505824f
C83 drain_right.n1 a_n1626_n3888# 3.36152f
C84 drain_right.t5 a_n1626_n3888# 0.505824f
C85 drain_right.t1 a_n1626_n3888# 0.505824f
C86 drain_right.n2 a_n1626_n3888# 3.36432f
C87 drain_right.n3 a_n1626_n3888# 2.4173f
C88 drain_right.t9 a_n1626_n3888# 0.505824f
C89 drain_right.t8 a_n1626_n3888# 0.505824f
C90 drain_right.n4 a_n1626_n3888# 3.36465f
C91 drain_right.t6 a_n1626_n3888# 0.505824f
C92 drain_right.t4 a_n1626_n3888# 0.505824f
C93 drain_right.n5 a_n1626_n3888# 3.36152f
C94 drain_right.n6 a_n1626_n3888# 0.672989f
C95 drain_right.t3 a_n1626_n3888# 0.505824f
C96 drain_right.t7 a_n1626_n3888# 0.505824f
C97 drain_right.n7 a_n1626_n3888# 3.36152f
C98 drain_right.n8 a_n1626_n3888# 0.567586f
C99 source.t2 a_n1626_n3888# 3.21033f
C100 source.n0 a_n1626_n3888# 1.42916f
C101 source.t8 a_n1626_n3888# 0.403181f
C102 source.t9 a_n1626_n3888# 0.403181f
C103 source.n1 a_n1626_n3888# 2.61162f
C104 source.n2 a_n1626_n3888# 0.302193f
C105 source.t1 a_n1626_n3888# 0.403181f
C106 source.t10 a_n1626_n3888# 0.403181f
C107 source.n3 a_n1626_n3888# 2.61162f
C108 source.n4 a_n1626_n3888# 0.302193f
C109 source.t4 a_n1626_n3888# 3.21033f
C110 source.n5 a_n1626_n3888# 0.422664f
C111 source.t21 a_n1626_n3888# 3.21033f
C112 source.n6 a_n1626_n3888# 0.422664f
C113 source.t23 a_n1626_n3888# 0.403181f
C114 source.t22 a_n1626_n3888# 0.403181f
C115 source.n7 a_n1626_n3888# 2.61162f
C116 source.n8 a_n1626_n3888# 0.302193f
C117 source.t20 a_n1626_n3888# 0.403181f
C118 source.t16 a_n1626_n3888# 0.403181f
C119 source.n9 a_n1626_n3888# 2.61162f
C120 source.n10 a_n1626_n3888# 0.302193f
C121 source.t13 a_n1626_n3888# 3.21033f
C122 source.n11 a_n1626_n3888# 1.80288f
C123 source.t11 a_n1626_n3888# 3.21033f
C124 source.n12 a_n1626_n3888# 1.80288f
C125 source.t0 a_n1626_n3888# 0.403181f
C126 source.t3 a_n1626_n3888# 0.403181f
C127 source.n13 a_n1626_n3888# 2.61162f
C128 source.n14 a_n1626_n3888# 0.302196f
C129 source.t6 a_n1626_n3888# 0.403181f
C130 source.t5 a_n1626_n3888# 0.403181f
C131 source.n15 a_n1626_n3888# 2.61162f
C132 source.n16 a_n1626_n3888# 0.302196f
C133 source.t7 a_n1626_n3888# 3.21033f
C134 source.n17 a_n1626_n3888# 0.422668f
C135 source.t18 a_n1626_n3888# 3.21033f
C136 source.n18 a_n1626_n3888# 0.422668f
C137 source.t14 a_n1626_n3888# 0.403181f
C138 source.t19 a_n1626_n3888# 0.403181f
C139 source.n19 a_n1626_n3888# 2.61162f
C140 source.n20 a_n1626_n3888# 0.302196f
C141 source.t12 a_n1626_n3888# 0.403181f
C142 source.t17 a_n1626_n3888# 0.403181f
C143 source.n21 a_n1626_n3888# 2.61162f
C144 source.n22 a_n1626_n3888# 0.302196f
C145 source.t15 a_n1626_n3888# 3.21033f
C146 source.n23 a_n1626_n3888# 0.550389f
C147 source.n24 a_n1626_n3888# 1.64218f
C148 minus.n0 a_n1626_n3888# 0.056364f
C149 minus.t8 a_n1626_n3888# 0.360785f
C150 minus.t4 a_n1626_n3888# 0.357773f
C151 minus.t5 a_n1626_n3888# 0.357773f
C152 minus.n1 a_n1626_n3888# 0.021304f
C153 minus.t3 a_n1626_n3888# 0.360785f
C154 minus.n2 a_n1626_n3888# 0.167961f
C155 minus.t7 a_n1626_n3888# 0.357773f
C156 minus.n3 a_n1626_n3888# 0.146111f
C157 minus.t2 a_n1626_n3888# 0.357773f
C158 minus.n4 a_n1626_n3888# 0.146111f
C159 minus.n5 a_n1626_n3888# 0.02391f
C160 minus.n6 a_n1626_n3888# 0.126545f
C161 minus.n7 a_n1626_n3888# 0.056364f
C162 minus.n8 a_n1626_n3888# 0.056364f
C163 minus.n9 a_n1626_n3888# 0.021304f
C164 minus.n10 a_n1626_n3888# 0.146111f
C165 minus.n11 a_n1626_n3888# 0.02391f
C166 minus.n12 a_n1626_n3888# 0.146111f
C167 minus.n13 a_n1626_n3888# 0.167879f
C168 minus.n14 a_n1626_n3888# 2.11461f
C169 minus.n15 a_n1626_n3888# 0.056364f
C170 minus.t6 a_n1626_n3888# 0.357773f
C171 minus.t0 a_n1626_n3888# 0.357773f
C172 minus.n16 a_n1626_n3888# 0.021304f
C173 minus.t1 a_n1626_n3888# 0.360785f
C174 minus.n17 a_n1626_n3888# 0.167961f
C175 minus.t9 a_n1626_n3888# 0.357773f
C176 minus.n18 a_n1626_n3888# 0.146111f
C177 minus.t11 a_n1626_n3888# 0.357773f
C178 minus.n19 a_n1626_n3888# 0.146111f
C179 minus.n20 a_n1626_n3888# 0.02391f
C180 minus.n21 a_n1626_n3888# 0.126545f
C181 minus.n22 a_n1626_n3888# 0.056364f
C182 minus.n23 a_n1626_n3888# 0.056364f
C183 minus.n24 a_n1626_n3888# 0.021304f
C184 minus.n25 a_n1626_n3888# 0.146111f
C185 minus.n26 a_n1626_n3888# 0.02391f
C186 minus.n27 a_n1626_n3888# 0.146111f
C187 minus.t10 a_n1626_n3888# 0.360785f
C188 minus.n28 a_n1626_n3888# 0.167879f
C189 minus.n29 a_n1626_n3888# 0.374079f
C190 minus.n30 a_n1626_n3888# 2.55628f
.ends

