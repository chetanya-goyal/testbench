* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t19 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 source.t3 minus.t0 drain_right.t19 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X3 source.t13 minus.t1 drain_right.t18 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X4 drain_right.t17 minus.t2 source.t10 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X5 a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X6 source.t18 plus.t1 drain_left.t18 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X7 drain_left.t17 plus.t2 source.t28 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X8 source.t15 minus.t3 drain_right.t16 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X9 drain_left.t16 plus.t3 source.t31 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 source.t20 plus.t4 drain_left.t15 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X12 drain_right.t15 minus.t4 source.t2 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 drain_left.t14 plus.t5 source.t32 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t39 minus.t5 drain_right.t14 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X16 source.t4 minus.t6 drain_right.t13 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_right.t12 minus.t7 source.t6 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X18 drain_right.t11 minus.t8 source.t37 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 source.t17 plus.t6 drain_left.t13 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X20 source.t36 minus.t9 drain_right.t10 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X21 drain_right.t9 minus.t10 source.t8 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X22 drain_right.t8 minus.t11 source.t7 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_right.t7 minus.t12 source.t38 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X24 source.t24 plus.t7 drain_left.t12 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X25 drain_left.t11 plus.t8 source.t34 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X26 source.t35 plus.t9 drain_left.t10 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X27 drain_right.t6 minus.t13 source.t11 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X28 drain_right.t5 minus.t14 source.t0 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X29 source.t14 minus.t15 drain_right.t4 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X30 source.t1 minus.t16 drain_right.t3 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X31 drain_left.t9 plus.t10 source.t25 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X32 source.t9 minus.t17 drain_right.t2 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X33 source.t26 plus.t11 drain_left.t8 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X34 drain_left.t7 plus.t12 source.t27 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X35 drain_left.t6 plus.t13 source.t30 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X36 source.t33 plus.t14 drain_left.t5 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X37 source.t22 plus.t15 drain_left.t4 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X38 source.t12 minus.t18 drain_right.t1 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X39 drain_right.t0 minus.t19 source.t5 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X40 source.t16 plus.t16 drain_left.t3 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X41 drain_left.t2 plus.t17 source.t23 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X42 drain_left.t1 plus.t18 source.t21 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X43 source.t29 plus.t19 drain_left.t0 a_n2146_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 plus.n6 plus.t9 592.277
R1 plus.n27 plus.t13 592.277
R2 plus.n36 plus.t12 592.277
R3 plus.n56 plus.t11 592.277
R4 plus.n5 plus.t18 530.201
R5 plus.n9 plus.t15 530.201
R6 plus.n3 plus.t10 530.201
R7 plus.n15 plus.t19 530.201
R8 plus.n17 plus.t17 530.201
R9 plus.n18 plus.t14 530.201
R10 plus.n24 plus.t8 530.201
R11 plus.n26 plus.t16 530.201
R12 plus.n35 plus.t7 530.201
R13 plus.n39 plus.t3 530.201
R14 plus.n33 plus.t1 530.201
R15 plus.n45 plus.t0 530.201
R16 plus.n47 plus.t6 530.201
R17 plus.n32 plus.t5 530.201
R18 plus.n53 plus.t4 530.201
R19 plus.n55 plus.t2 530.201
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 69.3793
R47 plus.n19 plus.n18 69.3793
R48 plus.n48 plus.n32 69.3793
R49 plus.n44 plus.n33 69.3793
R50 plus.n9 plus.n8 54.7732
R51 plus.n25 plus.n24 54.7732
R52 plus.n54 plus.n53 54.7732
R53 plus.n39 plus.n38 54.7732
R54 plus.n16 plus.n15 47.4702
R55 plus.n17 plus.n16 47.4702
R56 plus.n47 plus.n46 47.4702
R57 plus.n46 plus.n45 47.4702
R58 plus.n8 plus.n5 40.1672
R59 plus.n26 plus.n25 40.1672
R60 plus.n55 plus.n54 40.1672
R61 plus.n38 plus.n35 40.1672
R62 plus.n6 plus.n5 32.8641
R63 plus.n27 plus.n26 32.8641
R64 plus.n56 plus.n55 32.8641
R65 plus.n36 plus.n35 32.8641
R66 plus plus.n57 27.4043
R67 plus.n15 plus.n14 25.5611
R68 plus.n19 plus.n17 25.5611
R69 plus.n48 plus.n47 25.5611
R70 plus.n45 plus.n44 25.5611
R71 plus.n10 plus.n9 18.2581
R72 plus.n24 plus.n23 18.2581
R73 plus.n53 plus.n52 18.2581
R74 plus.n40 plus.n39 18.2581
R75 plus plus.n28 8.41717
R76 plus.n11 plus.n3 3.65202
R77 plus.n18 plus.n1 3.65202
R78 plus.n32 plus.n30 3.65202
R79 plus.n41 plus.n33 3.65202
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n0 source.t30 99.1169
R99 source.n9 source.t35 99.1169
R100 source.n10 source.t6 99.1169
R101 source.n19 source.t12 99.1169
R102 source.n39 source.t10 99.1168
R103 source.n30 source.t13 99.1168
R104 source.n29 source.t27 99.1168
R105 source.n20 source.t26 99.1168
R106 source.n2 source.n1 84.1169
R107 source.n4 source.n3 84.1169
R108 source.n6 source.n5 84.1169
R109 source.n8 source.n7 84.1169
R110 source.n12 source.n11 84.1169
R111 source.n14 source.n13 84.1169
R112 source.n16 source.n15 84.1169
R113 source.n18 source.n17 84.1169
R114 source.n38 source.n37 84.1168
R115 source.n36 source.n35 84.1168
R116 source.n34 source.n33 84.1168
R117 source.n32 source.n31 84.1168
R118 source.n28 source.n27 84.1168
R119 source.n26 source.n25 84.1168
R120 source.n24 source.n23 84.1168
R121 source.n22 source.n21 84.1168
R122 source.n37 source.t8 15.0005
R123 source.n37 source.t15 15.0005
R124 source.n35 source.t5 15.0005
R125 source.n35 source.t1 15.0005
R126 source.n33 source.t2 15.0005
R127 source.n33 source.t3 15.0005
R128 source.n31 source.t38 15.0005
R129 source.n31 source.t4 15.0005
R130 source.n27 source.t31 15.0005
R131 source.n27 source.t24 15.0005
R132 source.n25 source.t19 15.0005
R133 source.n25 source.t18 15.0005
R134 source.n23 source.t32 15.0005
R135 source.n23 source.t17 15.0005
R136 source.n21 source.t28 15.0005
R137 source.n21 source.t20 15.0005
R138 source.n1 source.t34 15.0005
R139 source.n1 source.t16 15.0005
R140 source.n3 source.t23 15.0005
R141 source.n3 source.t33 15.0005
R142 source.n5 source.t25 15.0005
R143 source.n5 source.t29 15.0005
R144 source.n7 source.t21 15.0005
R145 source.n7 source.t22 15.0005
R146 source.n11 source.t11 15.0005
R147 source.n11 source.t39 15.0005
R148 source.n13 source.t37 15.0005
R149 source.n13 source.t36 15.0005
R150 source.n15 source.t0 15.0005
R151 source.n15 source.t9 15.0005
R152 source.n17 source.t7 15.0005
R153 source.n17 source.t14 15.0005
R154 source.n20 source.n19 14.2723
R155 source.n40 source.n0 8.72921
R156 source.n40 source.n39 5.5436
R157 source.n19 source.n18 0.560845
R158 source.n18 source.n16 0.560845
R159 source.n16 source.n14 0.560845
R160 source.n14 source.n12 0.560845
R161 source.n12 source.n10 0.560845
R162 source.n9 source.n8 0.560845
R163 source.n8 source.n6 0.560845
R164 source.n6 source.n4 0.560845
R165 source.n4 source.n2 0.560845
R166 source.n2 source.n0 0.560845
R167 source.n22 source.n20 0.560845
R168 source.n24 source.n22 0.560845
R169 source.n26 source.n24 0.560845
R170 source.n28 source.n26 0.560845
R171 source.n29 source.n28 0.560845
R172 source.n32 source.n30 0.560845
R173 source.n34 source.n32 0.560845
R174 source.n36 source.n34 0.560845
R175 source.n38 source.n36 0.560845
R176 source.n39 source.n38 0.560845
R177 source.n10 source.n9 0.470328
R178 source.n30 source.n29 0.470328
R179 source source.n40 0.188
R180 drain_left.n10 drain_left.n8 101.356
R181 drain_left.n6 drain_left.n4 101.356
R182 drain_left.n2 drain_left.n0 101.356
R183 drain_left.n16 drain_left.n15 100.796
R184 drain_left.n14 drain_left.n13 100.796
R185 drain_left.n12 drain_left.n11 100.796
R186 drain_left.n10 drain_left.n9 100.796
R187 drain_left.n7 drain_left.n3 100.796
R188 drain_left.n6 drain_left.n5 100.796
R189 drain_left.n2 drain_left.n1 100.796
R190 drain_left drain_left.n7 24.2741
R191 drain_left.n3 drain_left.t13 15.0005
R192 drain_left.n3 drain_left.t19 15.0005
R193 drain_left.n4 drain_left.t12 15.0005
R194 drain_left.n4 drain_left.t7 15.0005
R195 drain_left.n5 drain_left.t18 15.0005
R196 drain_left.n5 drain_left.t16 15.0005
R197 drain_left.n1 drain_left.t15 15.0005
R198 drain_left.n1 drain_left.t14 15.0005
R199 drain_left.n0 drain_left.t8 15.0005
R200 drain_left.n0 drain_left.t17 15.0005
R201 drain_left.n15 drain_left.t3 15.0005
R202 drain_left.n15 drain_left.t6 15.0005
R203 drain_left.n13 drain_left.t5 15.0005
R204 drain_left.n13 drain_left.t11 15.0005
R205 drain_left.n11 drain_left.t0 15.0005
R206 drain_left.n11 drain_left.t2 15.0005
R207 drain_left.n9 drain_left.t4 15.0005
R208 drain_left.n9 drain_left.t9 15.0005
R209 drain_left.n8 drain_left.t10 15.0005
R210 drain_left.n8 drain_left.t1 15.0005
R211 drain_left drain_left.n16 6.21356
R212 drain_left.n12 drain_left.n10 0.560845
R213 drain_left.n14 drain_left.n12 0.560845
R214 drain_left.n16 drain_left.n14 0.560845
R215 drain_left.n7 drain_left.n6 0.505499
R216 drain_left.n7 drain_left.n2 0.505499
R217 minus.n27 minus.t18 592.277
R218 minus.n7 minus.t7 592.277
R219 minus.n56 minus.t2 592.277
R220 minus.n35 minus.t1 592.277
R221 minus.n26 minus.t11 530.201
R222 minus.n24 minus.t15 530.201
R223 minus.n3 minus.t14 530.201
R224 minus.n18 minus.t17 530.201
R225 minus.n16 minus.t8 530.201
R226 minus.n4 minus.t9 530.201
R227 minus.n10 minus.t13 530.201
R228 minus.n6 minus.t5 530.201
R229 minus.n55 minus.t3 530.201
R230 minus.n53 minus.t10 530.201
R231 minus.n47 minus.t16 530.201
R232 minus.n46 minus.t19 530.201
R233 minus.n44 minus.t0 530.201
R234 minus.n32 minus.t4 530.201
R235 minus.n38 minus.t6 530.201
R236 minus.n34 minus.t12 530.201
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 69.3793
R264 minus.n15 minus.n4 69.3793
R265 minus.n43 minus.n32 69.3793
R266 minus.n48 minus.n47 69.3793
R267 minus.n25 minus.n24 54.7732
R268 minus.n10 minus.n9 54.7732
R269 minus.n38 minus.n37 54.7732
R270 minus.n54 minus.n53 54.7732
R271 minus.n18 minus.n17 47.4702
R272 minus.n17 minus.n16 47.4702
R273 minus.n45 minus.n44 47.4702
R274 minus.n46 minus.n45 47.4702
R275 minus.n26 minus.n25 40.1672
R276 minus.n9 minus.n6 40.1672
R277 minus.n37 minus.n34 40.1672
R278 minus.n55 minus.n54 40.1672
R279 minus.n27 minus.n26 32.8641
R280 minus.n7 minus.n6 32.8641
R281 minus.n35 minus.n34 32.8641
R282 minus.n56 minus.n55 32.8641
R283 minus.n58 minus.n28 29.7353
R284 minus.n19 minus.n18 25.5611
R285 minus.n16 minus.n15 25.5611
R286 minus.n44 minus.n43 25.5611
R287 minus.n48 minus.n46 25.5611
R288 minus.n24 minus.n23 18.2581
R289 minus.n11 minus.n10 18.2581
R290 minus.n39 minus.n38 18.2581
R291 minus.n53 minus.n52 18.2581
R292 minus.n58 minus.n57 6.56111
R293 minus.n3 minus.n1 3.65202
R294 minus.n12 minus.n4 3.65202
R295 minus.n40 minus.n32 3.65202
R296 minus.n47 minus.n30 3.65202
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 101.356
R317 drain_right.n6 drain_right.n4 101.356
R318 drain_right.n2 drain_right.n0 101.356
R319 drain_right.n10 drain_right.n9 100.796
R320 drain_right.n12 drain_right.n11 100.796
R321 drain_right.n14 drain_right.n13 100.796
R322 drain_right.n16 drain_right.n15 100.796
R323 drain_right.n7 drain_right.n3 100.796
R324 drain_right.n6 drain_right.n5 100.796
R325 drain_right.n2 drain_right.n1 100.796
R326 drain_right drain_right.n7 23.7208
R327 drain_right.n3 drain_right.t19 15.0005
R328 drain_right.n3 drain_right.t0 15.0005
R329 drain_right.n4 drain_right.t16 15.0005
R330 drain_right.n4 drain_right.t17 15.0005
R331 drain_right.n5 drain_right.t3 15.0005
R332 drain_right.n5 drain_right.t9 15.0005
R333 drain_right.n1 drain_right.t13 15.0005
R334 drain_right.n1 drain_right.t15 15.0005
R335 drain_right.n0 drain_right.t18 15.0005
R336 drain_right.n0 drain_right.t7 15.0005
R337 drain_right.n8 drain_right.t14 15.0005
R338 drain_right.n8 drain_right.t12 15.0005
R339 drain_right.n9 drain_right.t10 15.0005
R340 drain_right.n9 drain_right.t6 15.0005
R341 drain_right.n11 drain_right.t2 15.0005
R342 drain_right.n11 drain_right.t11 15.0005
R343 drain_right.n13 drain_right.t4 15.0005
R344 drain_right.n13 drain_right.t5 15.0005
R345 drain_right.n15 drain_right.t1 15.0005
R346 drain_right.n15 drain_right.t8 15.0005
R347 drain_right drain_right.n16 6.21356
R348 drain_right.n16 drain_right.n14 0.560845
R349 drain_right.n14 drain_right.n12 0.560845
R350 drain_right.n12 drain_right.n10 0.560845
R351 drain_right.n7 drain_right.n6 0.505499
R352 drain_right.n7 drain_right.n2 0.505499
C0 drain_right source 9.19201f
C1 drain_left plus 1.40472f
C2 drain_left minus 0.177493f
C3 plus minus 3.9694f
C4 drain_left source 9.191509f
C5 plus source 1.36068f
C6 minus source 1.34671f
C7 drain_left drain_right 1.13588f
C8 drain_right plus 0.371711f
C9 drain_right minus 1.19407f
C10 drain_right a_n2146_n1288# 4.28089f
C11 drain_left a_n2146_n1288# 4.57101f
C12 source a_n2146_n1288# 3.345717f
C13 minus a_n2146_n1288# 7.122226f
C14 plus a_n2146_n1288# 7.900694f
C15 drain_right.t18 a_n2146_n1288# 0.059468f
C16 drain_right.t7 a_n2146_n1288# 0.059468f
C17 drain_right.n0 a_n2146_n1288# 0.288616f
C18 drain_right.t13 a_n2146_n1288# 0.059468f
C19 drain_right.t15 a_n2146_n1288# 0.059468f
C20 drain_right.n1 a_n2146_n1288# 0.287014f
C21 drain_right.n2 a_n2146_n1288# 0.564623f
C22 drain_right.t19 a_n2146_n1288# 0.059468f
C23 drain_right.t0 a_n2146_n1288# 0.059468f
C24 drain_right.n3 a_n2146_n1288# 0.287014f
C25 drain_right.t16 a_n2146_n1288# 0.059468f
C26 drain_right.t17 a_n2146_n1288# 0.059468f
C27 drain_right.n4 a_n2146_n1288# 0.288616f
C28 drain_right.t3 a_n2146_n1288# 0.059468f
C29 drain_right.t9 a_n2146_n1288# 0.059468f
C30 drain_right.n5 a_n2146_n1288# 0.287014f
C31 drain_right.n6 a_n2146_n1288# 0.564623f
C32 drain_right.n7 a_n2146_n1288# 0.972476f
C33 drain_right.t14 a_n2146_n1288# 0.059468f
C34 drain_right.t12 a_n2146_n1288# 0.059468f
C35 drain_right.n8 a_n2146_n1288# 0.288617f
C36 drain_right.t10 a_n2146_n1288# 0.059468f
C37 drain_right.t6 a_n2146_n1288# 0.059468f
C38 drain_right.n9 a_n2146_n1288# 0.287015f
C39 drain_right.n10 a_n2146_n1288# 0.56791f
C40 drain_right.t2 a_n2146_n1288# 0.059468f
C41 drain_right.t11 a_n2146_n1288# 0.059468f
C42 drain_right.n11 a_n2146_n1288# 0.287015f
C43 drain_right.n12 a_n2146_n1288# 0.279755f
C44 drain_right.t4 a_n2146_n1288# 0.059468f
C45 drain_right.t5 a_n2146_n1288# 0.059468f
C46 drain_right.n13 a_n2146_n1288# 0.287015f
C47 drain_right.n14 a_n2146_n1288# 0.279755f
C48 drain_right.t1 a_n2146_n1288# 0.059468f
C49 drain_right.t8 a_n2146_n1288# 0.059468f
C50 drain_right.n15 a_n2146_n1288# 0.287015f
C51 drain_right.n16 a_n2146_n1288# 0.487145f
C52 minus.n0 a_n2146_n1288# 0.031379f
C53 minus.t18 a_n2146_n1288# 0.030388f
C54 minus.t11 a_n2146_n1288# 0.027701f
C55 minus.t15 a_n2146_n1288# 0.027701f
C56 minus.n1 a_n2146_n1288# 0.010893f
C57 minus.n2 a_n2146_n1288# 0.031379f
C58 minus.t14 a_n2146_n1288# 0.027701f
C59 minus.n3 a_n2146_n1288# 0.024183f
C60 minus.t17 a_n2146_n1288# 0.027701f
C61 minus.t8 a_n2146_n1288# 0.027701f
C62 minus.t9 a_n2146_n1288# 0.027701f
C63 minus.n4 a_n2146_n1288# 0.024183f
C64 minus.n5 a_n2146_n1288# 0.031379f
C65 minus.t13 a_n2146_n1288# 0.027701f
C66 minus.t5 a_n2146_n1288# 0.027701f
C67 minus.n6 a_n2146_n1288# 0.024183f
C68 minus.t7 a_n2146_n1288# 0.030388f
C69 minus.n7 a_n2146_n1288# 0.036307f
C70 minus.n8 a_n2146_n1288# 0.072384f
C71 minus.n9 a_n2146_n1288# 0.013311f
C72 minus.n10 a_n2146_n1288# 0.024183f
C73 minus.n11 a_n2146_n1288# 0.012828f
C74 minus.n12 a_n2146_n1288# 0.010893f
C75 minus.n13 a_n2146_n1288# 0.031379f
C76 minus.n14 a_n2146_n1288# 0.031379f
C77 minus.n15 a_n2146_n1288# 0.013311f
C78 minus.n16 a_n2146_n1288# 0.024183f
C79 minus.n17 a_n2146_n1288# 0.013311f
C80 minus.n18 a_n2146_n1288# 0.024183f
C81 minus.n19 a_n2146_n1288# 0.013311f
C82 minus.n20 a_n2146_n1288# 0.031379f
C83 minus.n21 a_n2146_n1288# 0.031379f
C84 minus.n22 a_n2146_n1288# 0.031379f
C85 minus.n23 a_n2146_n1288# 0.012828f
C86 minus.n24 a_n2146_n1288# 0.024183f
C87 minus.n25 a_n2146_n1288# 0.013311f
C88 minus.n26 a_n2146_n1288# 0.024183f
C89 minus.n27 a_n2146_n1288# 0.036259f
C90 minus.n28 a_n2146_n1288# 0.805822f
C91 minus.n29 a_n2146_n1288# 0.031379f
C92 minus.t3 a_n2146_n1288# 0.027701f
C93 minus.t10 a_n2146_n1288# 0.027701f
C94 minus.n30 a_n2146_n1288# 0.010893f
C95 minus.n31 a_n2146_n1288# 0.031379f
C96 minus.t19 a_n2146_n1288# 0.027701f
C97 minus.t0 a_n2146_n1288# 0.027701f
C98 minus.t4 a_n2146_n1288# 0.027701f
C99 minus.n32 a_n2146_n1288# 0.024183f
C100 minus.n33 a_n2146_n1288# 0.031379f
C101 minus.t6 a_n2146_n1288# 0.027701f
C102 minus.t12 a_n2146_n1288# 0.027701f
C103 minus.n34 a_n2146_n1288# 0.024183f
C104 minus.t1 a_n2146_n1288# 0.030388f
C105 minus.n35 a_n2146_n1288# 0.036307f
C106 minus.n36 a_n2146_n1288# 0.072384f
C107 minus.n37 a_n2146_n1288# 0.013311f
C108 minus.n38 a_n2146_n1288# 0.024183f
C109 minus.n39 a_n2146_n1288# 0.012828f
C110 minus.n40 a_n2146_n1288# 0.010893f
C111 minus.n41 a_n2146_n1288# 0.031379f
C112 minus.n42 a_n2146_n1288# 0.031379f
C113 minus.n43 a_n2146_n1288# 0.013311f
C114 minus.n44 a_n2146_n1288# 0.024183f
C115 minus.n45 a_n2146_n1288# 0.013311f
C116 minus.n46 a_n2146_n1288# 0.024183f
C117 minus.t16 a_n2146_n1288# 0.027701f
C118 minus.n47 a_n2146_n1288# 0.024183f
C119 minus.n48 a_n2146_n1288# 0.013311f
C120 minus.n49 a_n2146_n1288# 0.031379f
C121 minus.n50 a_n2146_n1288# 0.031379f
C122 minus.n51 a_n2146_n1288# 0.031379f
C123 minus.n52 a_n2146_n1288# 0.012828f
C124 minus.n53 a_n2146_n1288# 0.024183f
C125 minus.n54 a_n2146_n1288# 0.013311f
C126 minus.n55 a_n2146_n1288# 0.024183f
C127 minus.t2 a_n2146_n1288# 0.030388f
C128 minus.n56 a_n2146_n1288# 0.036259f
C129 minus.n57 a_n2146_n1288# 0.209654f
C130 minus.n58 a_n2146_n1288# 0.992251f
C131 drain_left.t8 a_n2146_n1288# 0.058847f
C132 drain_left.t17 a_n2146_n1288# 0.058847f
C133 drain_left.n0 a_n2146_n1288# 0.2856f
C134 drain_left.t15 a_n2146_n1288# 0.058847f
C135 drain_left.t14 a_n2146_n1288# 0.058847f
C136 drain_left.n1 a_n2146_n1288# 0.284015f
C137 drain_left.n2 a_n2146_n1288# 0.558724f
C138 drain_left.t13 a_n2146_n1288# 0.058847f
C139 drain_left.t19 a_n2146_n1288# 0.058847f
C140 drain_left.n3 a_n2146_n1288# 0.284015f
C141 drain_left.t12 a_n2146_n1288# 0.058847f
C142 drain_left.t7 a_n2146_n1288# 0.058847f
C143 drain_left.n4 a_n2146_n1288# 0.2856f
C144 drain_left.t18 a_n2146_n1288# 0.058847f
C145 drain_left.t16 a_n2146_n1288# 0.058847f
C146 drain_left.n5 a_n2146_n1288# 0.284015f
C147 drain_left.n6 a_n2146_n1288# 0.558724f
C148 drain_left.n7 a_n2146_n1288# 1.01031f
C149 drain_left.t10 a_n2146_n1288# 0.058847f
C150 drain_left.t1 a_n2146_n1288# 0.058847f
C151 drain_left.n8 a_n2146_n1288# 0.285601f
C152 drain_left.t4 a_n2146_n1288# 0.058847f
C153 drain_left.t9 a_n2146_n1288# 0.058847f
C154 drain_left.n9 a_n2146_n1288# 0.284016f
C155 drain_left.n10 a_n2146_n1288# 0.561976f
C156 drain_left.t0 a_n2146_n1288# 0.058847f
C157 drain_left.t2 a_n2146_n1288# 0.058847f
C158 drain_left.n11 a_n2146_n1288# 0.284016f
C159 drain_left.n12 a_n2146_n1288# 0.276831f
C160 drain_left.t5 a_n2146_n1288# 0.058847f
C161 drain_left.t11 a_n2146_n1288# 0.058847f
C162 drain_left.n13 a_n2146_n1288# 0.284016f
C163 drain_left.n14 a_n2146_n1288# 0.276831f
C164 drain_left.t3 a_n2146_n1288# 0.058847f
C165 drain_left.t6 a_n2146_n1288# 0.058847f
C166 drain_left.n15 a_n2146_n1288# 0.284016f
C167 drain_left.n16 a_n2146_n1288# 0.482055f
C168 source.t30 a_n2146_n1288# 0.326821f
C169 source.n0 a_n2146_n1288# 0.622913f
C170 source.t34 a_n2146_n1288# 0.062247f
C171 source.t16 a_n2146_n1288# 0.062247f
C172 source.n1 a_n2146_n1288# 0.261957f
C173 source.n2 a_n2146_n1288# 0.295963f
C174 source.t23 a_n2146_n1288# 0.062247f
C175 source.t33 a_n2146_n1288# 0.062247f
C176 source.n3 a_n2146_n1288# 0.261957f
C177 source.n4 a_n2146_n1288# 0.295963f
C178 source.t25 a_n2146_n1288# 0.062247f
C179 source.t29 a_n2146_n1288# 0.062247f
C180 source.n5 a_n2146_n1288# 0.261957f
C181 source.n6 a_n2146_n1288# 0.295963f
C182 source.t21 a_n2146_n1288# 0.062247f
C183 source.t22 a_n2146_n1288# 0.062247f
C184 source.n7 a_n2146_n1288# 0.261957f
C185 source.n8 a_n2146_n1288# 0.295963f
C186 source.t35 a_n2146_n1288# 0.326821f
C187 source.n9 a_n2146_n1288# 0.335561f
C188 source.t6 a_n2146_n1288# 0.326821f
C189 source.n10 a_n2146_n1288# 0.335561f
C190 source.t11 a_n2146_n1288# 0.062247f
C191 source.t39 a_n2146_n1288# 0.062247f
C192 source.n11 a_n2146_n1288# 0.261957f
C193 source.n12 a_n2146_n1288# 0.295963f
C194 source.t37 a_n2146_n1288# 0.062247f
C195 source.t36 a_n2146_n1288# 0.062247f
C196 source.n13 a_n2146_n1288# 0.261957f
C197 source.n14 a_n2146_n1288# 0.295963f
C198 source.t0 a_n2146_n1288# 0.062247f
C199 source.t9 a_n2146_n1288# 0.062247f
C200 source.n15 a_n2146_n1288# 0.261957f
C201 source.n16 a_n2146_n1288# 0.295963f
C202 source.t7 a_n2146_n1288# 0.062247f
C203 source.t14 a_n2146_n1288# 0.062247f
C204 source.n17 a_n2146_n1288# 0.261957f
C205 source.n18 a_n2146_n1288# 0.295963f
C206 source.t12 a_n2146_n1288# 0.326821f
C207 source.n19 a_n2146_n1288# 0.865581f
C208 source.t26 a_n2146_n1288# 0.32682f
C209 source.n20 a_n2146_n1288# 0.865583f
C210 source.t28 a_n2146_n1288# 0.062247f
C211 source.t20 a_n2146_n1288# 0.062247f
C212 source.n21 a_n2146_n1288# 0.261955f
C213 source.n22 a_n2146_n1288# 0.295964f
C214 source.t32 a_n2146_n1288# 0.062247f
C215 source.t17 a_n2146_n1288# 0.062247f
C216 source.n23 a_n2146_n1288# 0.261955f
C217 source.n24 a_n2146_n1288# 0.295964f
C218 source.t19 a_n2146_n1288# 0.062247f
C219 source.t18 a_n2146_n1288# 0.062247f
C220 source.n25 a_n2146_n1288# 0.261955f
C221 source.n26 a_n2146_n1288# 0.295964f
C222 source.t31 a_n2146_n1288# 0.062247f
C223 source.t24 a_n2146_n1288# 0.062247f
C224 source.n27 a_n2146_n1288# 0.261955f
C225 source.n28 a_n2146_n1288# 0.295964f
C226 source.t27 a_n2146_n1288# 0.32682f
C227 source.n29 a_n2146_n1288# 0.335562f
C228 source.t13 a_n2146_n1288# 0.32682f
C229 source.n30 a_n2146_n1288# 0.335562f
C230 source.t38 a_n2146_n1288# 0.062247f
C231 source.t4 a_n2146_n1288# 0.062247f
C232 source.n31 a_n2146_n1288# 0.261955f
C233 source.n32 a_n2146_n1288# 0.295964f
C234 source.t2 a_n2146_n1288# 0.062247f
C235 source.t3 a_n2146_n1288# 0.062247f
C236 source.n33 a_n2146_n1288# 0.261955f
C237 source.n34 a_n2146_n1288# 0.295964f
C238 source.t5 a_n2146_n1288# 0.062247f
C239 source.t1 a_n2146_n1288# 0.062247f
C240 source.n35 a_n2146_n1288# 0.261955f
C241 source.n36 a_n2146_n1288# 0.295964f
C242 source.t8 a_n2146_n1288# 0.062247f
C243 source.t15 a_n2146_n1288# 0.062247f
C244 source.n37 a_n2146_n1288# 0.261955f
C245 source.n38 a_n2146_n1288# 0.295964f
C246 source.t10 a_n2146_n1288# 0.32682f
C247 source.n39 a_n2146_n1288# 0.483453f
C248 source.n40 a_n2146_n1288# 0.643287f
C249 plus.n0 a_n2146_n1288# 0.031885f
C250 plus.t16 a_n2146_n1288# 0.028148f
C251 plus.t8 a_n2146_n1288# 0.028148f
C252 plus.n1 a_n2146_n1288# 0.011069f
C253 plus.n2 a_n2146_n1288# 0.031885f
C254 plus.t17 a_n2146_n1288# 0.028148f
C255 plus.t19 a_n2146_n1288# 0.028148f
C256 plus.t10 a_n2146_n1288# 0.028148f
C257 plus.n3 a_n2146_n1288# 0.024573f
C258 plus.n4 a_n2146_n1288# 0.031885f
C259 plus.t15 a_n2146_n1288# 0.028148f
C260 plus.t18 a_n2146_n1288# 0.028148f
C261 plus.n5 a_n2146_n1288# 0.024573f
C262 plus.t9 a_n2146_n1288# 0.030878f
C263 plus.n6 a_n2146_n1288# 0.036893f
C264 plus.n7 a_n2146_n1288# 0.073551f
C265 plus.n8 a_n2146_n1288# 0.013526f
C266 plus.n9 a_n2146_n1288# 0.024573f
C267 plus.n10 a_n2146_n1288# 0.013035f
C268 plus.n11 a_n2146_n1288# 0.011069f
C269 plus.n12 a_n2146_n1288# 0.031885f
C270 plus.n13 a_n2146_n1288# 0.031885f
C271 plus.n14 a_n2146_n1288# 0.013526f
C272 plus.n15 a_n2146_n1288# 0.024573f
C273 plus.n16 a_n2146_n1288# 0.013526f
C274 plus.n17 a_n2146_n1288# 0.024573f
C275 plus.t14 a_n2146_n1288# 0.028148f
C276 plus.n18 a_n2146_n1288# 0.024573f
C277 plus.n19 a_n2146_n1288# 0.013526f
C278 plus.n20 a_n2146_n1288# 0.031885f
C279 plus.n21 a_n2146_n1288# 0.031885f
C280 plus.n22 a_n2146_n1288# 0.031885f
C281 plus.n23 a_n2146_n1288# 0.013035f
C282 plus.n24 a_n2146_n1288# 0.024573f
C283 plus.n25 a_n2146_n1288# 0.013526f
C284 plus.n26 a_n2146_n1288# 0.024573f
C285 plus.t13 a_n2146_n1288# 0.030878f
C286 plus.n27 a_n2146_n1288# 0.036844f
C287 plus.n28 a_n2146_n1288# 0.232768f
C288 plus.n29 a_n2146_n1288# 0.031885f
C289 plus.t11 a_n2146_n1288# 0.030878f
C290 plus.t2 a_n2146_n1288# 0.028148f
C291 plus.t4 a_n2146_n1288# 0.028148f
C292 plus.n30 a_n2146_n1288# 0.011069f
C293 plus.n31 a_n2146_n1288# 0.031885f
C294 plus.t5 a_n2146_n1288# 0.028148f
C295 plus.n32 a_n2146_n1288# 0.024573f
C296 plus.t6 a_n2146_n1288# 0.028148f
C297 plus.t0 a_n2146_n1288# 0.028148f
C298 plus.t1 a_n2146_n1288# 0.028148f
C299 plus.n33 a_n2146_n1288# 0.024573f
C300 plus.n34 a_n2146_n1288# 0.031885f
C301 plus.t3 a_n2146_n1288# 0.028148f
C302 plus.t7 a_n2146_n1288# 0.028148f
C303 plus.n35 a_n2146_n1288# 0.024573f
C304 plus.t12 a_n2146_n1288# 0.030878f
C305 plus.n36 a_n2146_n1288# 0.036893f
C306 plus.n37 a_n2146_n1288# 0.073551f
C307 plus.n38 a_n2146_n1288# 0.013526f
C308 plus.n39 a_n2146_n1288# 0.024573f
C309 plus.n40 a_n2146_n1288# 0.013035f
C310 plus.n41 a_n2146_n1288# 0.011069f
C311 plus.n42 a_n2146_n1288# 0.031885f
C312 plus.n43 a_n2146_n1288# 0.031885f
C313 plus.n44 a_n2146_n1288# 0.013526f
C314 plus.n45 a_n2146_n1288# 0.024573f
C315 plus.n46 a_n2146_n1288# 0.013526f
C316 plus.n47 a_n2146_n1288# 0.024573f
C317 plus.n48 a_n2146_n1288# 0.013526f
C318 plus.n49 a_n2146_n1288# 0.031885f
C319 plus.n50 a_n2146_n1288# 0.031885f
C320 plus.n51 a_n2146_n1288# 0.031885f
C321 plus.n52 a_n2146_n1288# 0.013035f
C322 plus.n53 a_n2146_n1288# 0.024573f
C323 plus.n54 a_n2146_n1288# 0.013526f
C324 plus.n55 a_n2146_n1288# 0.024573f
C325 plus.n56 a_n2146_n1288# 0.036844f
C326 plus.n57 a_n2146_n1288# 0.780238f
.ends

