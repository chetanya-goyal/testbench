* NGSPICE file created from diffpair277.ext - technology: sky130A

.subckt diffpair277 minus drain_right drain_left source plus
X0 source.t31 minus.t0 drain_right.t4 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t30 minus.t1 drain_right.t11 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X2 drain_left.t15 plus.t0 source.t0 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X3 source.t29 minus.t2 drain_right.t7 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X4 drain_right.t6 minus.t3 source.t28 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X5 a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X6 source.t14 plus.t1 drain_left.t14 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 source.t2 plus.t2 drain_left.t13 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X8 source.t9 plus.t3 drain_left.t12 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X9 source.t11 plus.t4 drain_left.t11 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X11 drain_right.t12 minus.t4 source.t27 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X12 drain_right.t0 minus.t5 source.t26 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X13 drain_right.t2 minus.t6 source.t25 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 drain_right.t13 minus.t7 source.t24 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X15 source.t6 plus.t5 drain_left.t10 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X16 drain_right.t10 minus.t8 source.t23 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X17 source.t15 plus.t6 drain_left.t9 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X18 drain_left.t8 plus.t7 source.t7 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X19 drain_left.t7 plus.t8 source.t10 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X20 drain_left.t6 plus.t9 source.t12 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X21 source.t22 minus.t9 drain_right.t9 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X22 drain_right.t5 minus.t10 source.t21 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X23 drain_left.t5 plus.t10 source.t4 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X24 a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X25 source.t20 minus.t11 drain_right.t3 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X26 source.t19 minus.t12 drain_right.t1 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X27 source.t1 plus.t11 drain_left.t4 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X28 drain_right.t8 minus.t13 source.t18 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X29 drain_left.t3 plus.t12 source.t3 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X30 drain_left.t2 plus.t13 source.t5 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X31 source.t17 minus.t14 drain_right.t15 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X32 source.t16 minus.t15 drain_right.t14 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X33 source.t13 plus.t14 drain_left.t1 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X34 a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X35 drain_left.t0 plus.t15 source.t8 a_n1850_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n21 minus.t15 616.376
R1 minus.n5 minus.t10 616.376
R2 minus.n44 minus.t7 616.376
R3 minus.n28 minus.t12 616.376
R4 minus.n20 minus.t4 586.433
R5 minus.n1 minus.t2 586.433
R6 minus.n14 minus.t13 586.433
R7 minus.n12 minus.t9 586.433
R8 minus.n3 minus.t3 586.433
R9 minus.n6 minus.t14 586.433
R10 minus.n43 minus.t0 586.433
R11 minus.n24 minus.t8 586.433
R12 minus.n37 minus.t1 586.433
R13 minus.n35 minus.t5 586.433
R14 minus.n26 minus.t11 586.433
R15 minus.n29 minus.t6 586.433
R16 minus.n5 minus.n4 161.489
R17 minus.n28 minus.n27 161.489
R18 minus.n22 minus.n21 161.3
R19 minus.n19 minus.n0 161.3
R20 minus.n18 minus.n17 161.3
R21 minus.n16 minus.n15 161.3
R22 minus.n13 minus.n2 161.3
R23 minus.n11 minus.n10 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n45 minus.n44 161.3
R27 minus.n42 minus.n23 161.3
R28 minus.n41 minus.n40 161.3
R29 minus.n39 minus.n38 161.3
R30 minus.n36 minus.n25 161.3
R31 minus.n34 minus.n33 161.3
R32 minus.n32 minus.n31 161.3
R33 minus.n30 minus.n27 161.3
R34 minus.n19 minus.n18 73.0308
R35 minus.n8 minus.n7 73.0308
R36 minus.n31 minus.n30 73.0308
R37 minus.n42 minus.n41 73.0308
R38 minus.n15 minus.n1 64.9975
R39 minus.n11 minus.n3 64.9975
R40 minus.n34 minus.n26 64.9975
R41 minus.n38 minus.n24 64.9975
R42 minus.n21 minus.n20 62.0763
R43 minus.n6 minus.n5 62.0763
R44 minus.n29 minus.n28 62.0763
R45 minus.n44 minus.n43 62.0763
R46 minus.n14 minus.n13 46.0096
R47 minus.n13 minus.n12 46.0096
R48 minus.n36 minus.n35 46.0096
R49 minus.n37 minus.n36 46.0096
R50 minus.n46 minus.n22 31.5497
R51 minus.n15 minus.n14 27.0217
R52 minus.n12 minus.n11 27.0217
R53 minus.n35 minus.n34 27.0217
R54 minus.n38 minus.n37 27.0217
R55 minus.n20 minus.n19 10.955
R56 minus.n7 minus.n6 10.955
R57 minus.n30 minus.n29 10.955
R58 minus.n43 minus.n42 10.955
R59 minus.n18 minus.n1 8.03383
R60 minus.n8 minus.n3 8.03383
R61 minus.n31 minus.n26 8.03383
R62 minus.n41 minus.n24 8.03383
R63 minus.n46 minus.n45 6.46641
R64 minus.n22 minus.n0 0.189894
R65 minus.n17 minus.n0 0.189894
R66 minus.n17 minus.n16 0.189894
R67 minus.n16 minus.n2 0.189894
R68 minus.n10 minus.n2 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n32 minus.n27 0.189894
R72 minus.n33 minus.n32 0.189894
R73 minus.n33 minus.n25 0.189894
R74 minus.n39 minus.n25 0.189894
R75 minus.n40 minus.n39 0.189894
R76 minus.n40 minus.n23 0.189894
R77 minus.n45 minus.n23 0.189894
R78 minus minus.n46 0.188
R79 drain_right.n5 drain_right.n3 67.7338
R80 drain_right.n2 drain_right.n0 67.7338
R81 drain_right.n9 drain_right.n7 67.7338
R82 drain_right.n9 drain_right.n8 67.1908
R83 drain_right.n11 drain_right.n10 67.1908
R84 drain_right.n13 drain_right.n12 67.1908
R85 drain_right.n5 drain_right.n4 67.1907
R86 drain_right.n2 drain_right.n1 67.1907
R87 drain_right drain_right.n6 25.7986
R88 drain_right drain_right.n13 6.19632
R89 drain_right.n3 drain_right.t4 3.3005
R90 drain_right.n3 drain_right.t13 3.3005
R91 drain_right.n4 drain_right.t11 3.3005
R92 drain_right.n4 drain_right.t10 3.3005
R93 drain_right.n1 drain_right.t3 3.3005
R94 drain_right.n1 drain_right.t0 3.3005
R95 drain_right.n0 drain_right.t1 3.3005
R96 drain_right.n0 drain_right.t2 3.3005
R97 drain_right.n7 drain_right.t15 3.3005
R98 drain_right.n7 drain_right.t5 3.3005
R99 drain_right.n8 drain_right.t9 3.3005
R100 drain_right.n8 drain_right.t6 3.3005
R101 drain_right.n10 drain_right.t7 3.3005
R102 drain_right.n10 drain_right.t8 3.3005
R103 drain_right.n12 drain_right.t14 3.3005
R104 drain_right.n12 drain_right.t12 3.3005
R105 drain_right.n13 drain_right.n11 0.543603
R106 drain_right.n11 drain_right.n9 0.543603
R107 drain_right.n6 drain_right.n5 0.216706
R108 drain_right.n6 drain_right.n2 0.216706
R109 source.n274 source.n248 289.615
R110 source.n236 source.n210 289.615
R111 source.n204 source.n178 289.615
R112 source.n166 source.n140 289.615
R113 source.n26 source.n0 289.615
R114 source.n64 source.n38 289.615
R115 source.n96 source.n70 289.615
R116 source.n134 source.n108 289.615
R117 source.n259 source.n258 185
R118 source.n256 source.n255 185
R119 source.n265 source.n264 185
R120 source.n267 source.n266 185
R121 source.n252 source.n251 185
R122 source.n273 source.n272 185
R123 source.n275 source.n274 185
R124 source.n221 source.n220 185
R125 source.n218 source.n217 185
R126 source.n227 source.n226 185
R127 source.n229 source.n228 185
R128 source.n214 source.n213 185
R129 source.n235 source.n234 185
R130 source.n237 source.n236 185
R131 source.n189 source.n188 185
R132 source.n186 source.n185 185
R133 source.n195 source.n194 185
R134 source.n197 source.n196 185
R135 source.n182 source.n181 185
R136 source.n203 source.n202 185
R137 source.n205 source.n204 185
R138 source.n151 source.n150 185
R139 source.n148 source.n147 185
R140 source.n157 source.n156 185
R141 source.n159 source.n158 185
R142 source.n144 source.n143 185
R143 source.n165 source.n164 185
R144 source.n167 source.n166 185
R145 source.n27 source.n26 185
R146 source.n25 source.n24 185
R147 source.n4 source.n3 185
R148 source.n19 source.n18 185
R149 source.n17 source.n16 185
R150 source.n8 source.n7 185
R151 source.n11 source.n10 185
R152 source.n65 source.n64 185
R153 source.n63 source.n62 185
R154 source.n42 source.n41 185
R155 source.n57 source.n56 185
R156 source.n55 source.n54 185
R157 source.n46 source.n45 185
R158 source.n49 source.n48 185
R159 source.n97 source.n96 185
R160 source.n95 source.n94 185
R161 source.n74 source.n73 185
R162 source.n89 source.n88 185
R163 source.n87 source.n86 185
R164 source.n78 source.n77 185
R165 source.n81 source.n80 185
R166 source.n135 source.n134 185
R167 source.n133 source.n132 185
R168 source.n112 source.n111 185
R169 source.n127 source.n126 185
R170 source.n125 source.n124 185
R171 source.n116 source.n115 185
R172 source.n119 source.n118 185
R173 source.t24 source.n257 147.661
R174 source.t19 source.n219 147.661
R175 source.t10 source.n187 147.661
R176 source.t6 source.n149 147.661
R177 source.t0 source.n9 147.661
R178 source.t2 source.n47 147.661
R179 source.t21 source.n79 147.661
R180 source.t16 source.n117 147.661
R181 source.n258 source.n255 104.615
R182 source.n265 source.n255 104.615
R183 source.n266 source.n265 104.615
R184 source.n266 source.n251 104.615
R185 source.n273 source.n251 104.615
R186 source.n274 source.n273 104.615
R187 source.n220 source.n217 104.615
R188 source.n227 source.n217 104.615
R189 source.n228 source.n227 104.615
R190 source.n228 source.n213 104.615
R191 source.n235 source.n213 104.615
R192 source.n236 source.n235 104.615
R193 source.n188 source.n185 104.615
R194 source.n195 source.n185 104.615
R195 source.n196 source.n195 104.615
R196 source.n196 source.n181 104.615
R197 source.n203 source.n181 104.615
R198 source.n204 source.n203 104.615
R199 source.n150 source.n147 104.615
R200 source.n157 source.n147 104.615
R201 source.n158 source.n157 104.615
R202 source.n158 source.n143 104.615
R203 source.n165 source.n143 104.615
R204 source.n166 source.n165 104.615
R205 source.n26 source.n25 104.615
R206 source.n25 source.n3 104.615
R207 source.n18 source.n3 104.615
R208 source.n18 source.n17 104.615
R209 source.n17 source.n7 104.615
R210 source.n10 source.n7 104.615
R211 source.n64 source.n63 104.615
R212 source.n63 source.n41 104.615
R213 source.n56 source.n41 104.615
R214 source.n56 source.n55 104.615
R215 source.n55 source.n45 104.615
R216 source.n48 source.n45 104.615
R217 source.n96 source.n95 104.615
R218 source.n95 source.n73 104.615
R219 source.n88 source.n73 104.615
R220 source.n88 source.n87 104.615
R221 source.n87 source.n77 104.615
R222 source.n80 source.n77 104.615
R223 source.n134 source.n133 104.615
R224 source.n133 source.n111 104.615
R225 source.n126 source.n111 104.615
R226 source.n126 source.n125 104.615
R227 source.n125 source.n115 104.615
R228 source.n118 source.n115 104.615
R229 source.n258 source.t24 52.3082
R230 source.n220 source.t19 52.3082
R231 source.n188 source.t10 52.3082
R232 source.n150 source.t6 52.3082
R233 source.n10 source.t0 52.3082
R234 source.n48 source.t2 52.3082
R235 source.n80 source.t21 52.3082
R236 source.n118 source.t16 52.3082
R237 source.n33 source.n32 50.512
R238 source.n35 source.n34 50.512
R239 source.n37 source.n36 50.512
R240 source.n103 source.n102 50.512
R241 source.n105 source.n104 50.512
R242 source.n107 source.n106 50.512
R243 source.n247 source.n246 50.5119
R244 source.n245 source.n244 50.5119
R245 source.n243 source.n242 50.5119
R246 source.n177 source.n176 50.5119
R247 source.n175 source.n174 50.5119
R248 source.n173 source.n172 50.5119
R249 source.n279 source.n278 32.1853
R250 source.n241 source.n240 32.1853
R251 source.n209 source.n208 32.1853
R252 source.n171 source.n170 32.1853
R253 source.n31 source.n30 32.1853
R254 source.n69 source.n68 32.1853
R255 source.n101 source.n100 32.1853
R256 source.n139 source.n138 32.1853
R257 source.n171 source.n139 17.2854
R258 source.n259 source.n257 15.6674
R259 source.n221 source.n219 15.6674
R260 source.n189 source.n187 15.6674
R261 source.n151 source.n149 15.6674
R262 source.n11 source.n9 15.6674
R263 source.n49 source.n47 15.6674
R264 source.n81 source.n79 15.6674
R265 source.n119 source.n117 15.6674
R266 source.n260 source.n256 12.8005
R267 source.n222 source.n218 12.8005
R268 source.n190 source.n186 12.8005
R269 source.n152 source.n148 12.8005
R270 source.n12 source.n8 12.8005
R271 source.n50 source.n46 12.8005
R272 source.n82 source.n78 12.8005
R273 source.n120 source.n116 12.8005
R274 source.n264 source.n263 12.0247
R275 source.n226 source.n225 12.0247
R276 source.n194 source.n193 12.0247
R277 source.n156 source.n155 12.0247
R278 source.n16 source.n15 12.0247
R279 source.n54 source.n53 12.0247
R280 source.n86 source.n85 12.0247
R281 source.n124 source.n123 12.0247
R282 source.n280 source.n31 11.7509
R283 source.n267 source.n254 11.249
R284 source.n229 source.n216 11.249
R285 source.n197 source.n184 11.249
R286 source.n159 source.n146 11.249
R287 source.n19 source.n6 11.249
R288 source.n57 source.n44 11.249
R289 source.n89 source.n76 11.249
R290 source.n127 source.n114 11.249
R291 source.n268 source.n252 10.4732
R292 source.n230 source.n214 10.4732
R293 source.n198 source.n182 10.4732
R294 source.n160 source.n144 10.4732
R295 source.n20 source.n4 10.4732
R296 source.n58 source.n42 10.4732
R297 source.n90 source.n74 10.4732
R298 source.n128 source.n112 10.4732
R299 source.n272 source.n271 9.69747
R300 source.n234 source.n233 9.69747
R301 source.n202 source.n201 9.69747
R302 source.n164 source.n163 9.69747
R303 source.n24 source.n23 9.69747
R304 source.n62 source.n61 9.69747
R305 source.n94 source.n93 9.69747
R306 source.n132 source.n131 9.69747
R307 source.n278 source.n277 9.45567
R308 source.n240 source.n239 9.45567
R309 source.n208 source.n207 9.45567
R310 source.n170 source.n169 9.45567
R311 source.n30 source.n29 9.45567
R312 source.n68 source.n67 9.45567
R313 source.n100 source.n99 9.45567
R314 source.n138 source.n137 9.45567
R315 source.n277 source.n276 9.3005
R316 source.n250 source.n249 9.3005
R317 source.n271 source.n270 9.3005
R318 source.n269 source.n268 9.3005
R319 source.n254 source.n253 9.3005
R320 source.n263 source.n262 9.3005
R321 source.n261 source.n260 9.3005
R322 source.n239 source.n238 9.3005
R323 source.n212 source.n211 9.3005
R324 source.n233 source.n232 9.3005
R325 source.n231 source.n230 9.3005
R326 source.n216 source.n215 9.3005
R327 source.n225 source.n224 9.3005
R328 source.n223 source.n222 9.3005
R329 source.n207 source.n206 9.3005
R330 source.n180 source.n179 9.3005
R331 source.n201 source.n200 9.3005
R332 source.n199 source.n198 9.3005
R333 source.n184 source.n183 9.3005
R334 source.n193 source.n192 9.3005
R335 source.n191 source.n190 9.3005
R336 source.n169 source.n168 9.3005
R337 source.n142 source.n141 9.3005
R338 source.n163 source.n162 9.3005
R339 source.n161 source.n160 9.3005
R340 source.n146 source.n145 9.3005
R341 source.n155 source.n154 9.3005
R342 source.n153 source.n152 9.3005
R343 source.n29 source.n28 9.3005
R344 source.n2 source.n1 9.3005
R345 source.n23 source.n22 9.3005
R346 source.n21 source.n20 9.3005
R347 source.n6 source.n5 9.3005
R348 source.n15 source.n14 9.3005
R349 source.n13 source.n12 9.3005
R350 source.n67 source.n66 9.3005
R351 source.n40 source.n39 9.3005
R352 source.n61 source.n60 9.3005
R353 source.n59 source.n58 9.3005
R354 source.n44 source.n43 9.3005
R355 source.n53 source.n52 9.3005
R356 source.n51 source.n50 9.3005
R357 source.n99 source.n98 9.3005
R358 source.n72 source.n71 9.3005
R359 source.n93 source.n92 9.3005
R360 source.n91 source.n90 9.3005
R361 source.n76 source.n75 9.3005
R362 source.n85 source.n84 9.3005
R363 source.n83 source.n82 9.3005
R364 source.n137 source.n136 9.3005
R365 source.n110 source.n109 9.3005
R366 source.n131 source.n130 9.3005
R367 source.n129 source.n128 9.3005
R368 source.n114 source.n113 9.3005
R369 source.n123 source.n122 9.3005
R370 source.n121 source.n120 9.3005
R371 source.n275 source.n250 8.92171
R372 source.n237 source.n212 8.92171
R373 source.n205 source.n180 8.92171
R374 source.n167 source.n142 8.92171
R375 source.n27 source.n2 8.92171
R376 source.n65 source.n40 8.92171
R377 source.n97 source.n72 8.92171
R378 source.n135 source.n110 8.92171
R379 source.n276 source.n248 8.14595
R380 source.n238 source.n210 8.14595
R381 source.n206 source.n178 8.14595
R382 source.n168 source.n140 8.14595
R383 source.n28 source.n0 8.14595
R384 source.n66 source.n38 8.14595
R385 source.n98 source.n70 8.14595
R386 source.n136 source.n108 8.14595
R387 source.n278 source.n248 5.81868
R388 source.n240 source.n210 5.81868
R389 source.n208 source.n178 5.81868
R390 source.n170 source.n140 5.81868
R391 source.n30 source.n0 5.81868
R392 source.n68 source.n38 5.81868
R393 source.n100 source.n70 5.81868
R394 source.n138 source.n108 5.81868
R395 source.n280 source.n279 5.53498
R396 source.n276 source.n275 5.04292
R397 source.n238 source.n237 5.04292
R398 source.n206 source.n205 5.04292
R399 source.n168 source.n167 5.04292
R400 source.n28 source.n27 5.04292
R401 source.n66 source.n65 5.04292
R402 source.n98 source.n97 5.04292
R403 source.n136 source.n135 5.04292
R404 source.n261 source.n257 4.38594
R405 source.n223 source.n219 4.38594
R406 source.n191 source.n187 4.38594
R407 source.n153 source.n149 4.38594
R408 source.n13 source.n9 4.38594
R409 source.n51 source.n47 4.38594
R410 source.n83 source.n79 4.38594
R411 source.n121 source.n117 4.38594
R412 source.n272 source.n250 4.26717
R413 source.n234 source.n212 4.26717
R414 source.n202 source.n180 4.26717
R415 source.n164 source.n142 4.26717
R416 source.n24 source.n2 4.26717
R417 source.n62 source.n40 4.26717
R418 source.n94 source.n72 4.26717
R419 source.n132 source.n110 4.26717
R420 source.n271 source.n252 3.49141
R421 source.n233 source.n214 3.49141
R422 source.n201 source.n182 3.49141
R423 source.n163 source.n144 3.49141
R424 source.n23 source.n4 3.49141
R425 source.n61 source.n42 3.49141
R426 source.n93 source.n74 3.49141
R427 source.n131 source.n112 3.49141
R428 source.n246 source.t23 3.3005
R429 source.n246 source.t31 3.3005
R430 source.n244 source.t26 3.3005
R431 source.n244 source.t30 3.3005
R432 source.n242 source.t25 3.3005
R433 source.n242 source.t20 3.3005
R434 source.n176 source.t12 3.3005
R435 source.n176 source.t14 3.3005
R436 source.n174 source.t3 3.3005
R437 source.n174 source.t9 3.3005
R438 source.n172 source.t5 3.3005
R439 source.n172 source.t11 3.3005
R440 source.n32 source.t4 3.3005
R441 source.n32 source.t13 3.3005
R442 source.n34 source.t8 3.3005
R443 source.n34 source.t15 3.3005
R444 source.n36 source.t7 3.3005
R445 source.n36 source.t1 3.3005
R446 source.n102 source.t28 3.3005
R447 source.n102 source.t17 3.3005
R448 source.n104 source.t18 3.3005
R449 source.n104 source.t22 3.3005
R450 source.n106 source.t27 3.3005
R451 source.n106 source.t29 3.3005
R452 source.n268 source.n267 2.71565
R453 source.n230 source.n229 2.71565
R454 source.n198 source.n197 2.71565
R455 source.n160 source.n159 2.71565
R456 source.n20 source.n19 2.71565
R457 source.n58 source.n57 2.71565
R458 source.n90 source.n89 2.71565
R459 source.n128 source.n127 2.71565
R460 source.n264 source.n254 1.93989
R461 source.n226 source.n216 1.93989
R462 source.n194 source.n184 1.93989
R463 source.n156 source.n146 1.93989
R464 source.n16 source.n6 1.93989
R465 source.n54 source.n44 1.93989
R466 source.n86 source.n76 1.93989
R467 source.n124 source.n114 1.93989
R468 source.n263 source.n256 1.16414
R469 source.n225 source.n218 1.16414
R470 source.n193 source.n186 1.16414
R471 source.n155 source.n148 1.16414
R472 source.n15 source.n8 1.16414
R473 source.n53 source.n46 1.16414
R474 source.n85 source.n78 1.16414
R475 source.n123 source.n116 1.16414
R476 source.n139 source.n107 0.543603
R477 source.n107 source.n105 0.543603
R478 source.n105 source.n103 0.543603
R479 source.n103 source.n101 0.543603
R480 source.n69 source.n37 0.543603
R481 source.n37 source.n35 0.543603
R482 source.n35 source.n33 0.543603
R483 source.n33 source.n31 0.543603
R484 source.n173 source.n171 0.543603
R485 source.n175 source.n173 0.543603
R486 source.n177 source.n175 0.543603
R487 source.n209 source.n177 0.543603
R488 source.n243 source.n241 0.543603
R489 source.n245 source.n243 0.543603
R490 source.n247 source.n245 0.543603
R491 source.n279 source.n247 0.543603
R492 source.n101 source.n69 0.470328
R493 source.n241 source.n209 0.470328
R494 source.n260 source.n259 0.388379
R495 source.n222 source.n221 0.388379
R496 source.n190 source.n189 0.388379
R497 source.n152 source.n151 0.388379
R498 source.n12 source.n11 0.388379
R499 source.n50 source.n49 0.388379
R500 source.n82 source.n81 0.388379
R501 source.n120 source.n119 0.388379
R502 source source.n280 0.188
R503 source.n262 source.n261 0.155672
R504 source.n262 source.n253 0.155672
R505 source.n269 source.n253 0.155672
R506 source.n270 source.n269 0.155672
R507 source.n270 source.n249 0.155672
R508 source.n277 source.n249 0.155672
R509 source.n224 source.n223 0.155672
R510 source.n224 source.n215 0.155672
R511 source.n231 source.n215 0.155672
R512 source.n232 source.n231 0.155672
R513 source.n232 source.n211 0.155672
R514 source.n239 source.n211 0.155672
R515 source.n192 source.n191 0.155672
R516 source.n192 source.n183 0.155672
R517 source.n199 source.n183 0.155672
R518 source.n200 source.n199 0.155672
R519 source.n200 source.n179 0.155672
R520 source.n207 source.n179 0.155672
R521 source.n154 source.n153 0.155672
R522 source.n154 source.n145 0.155672
R523 source.n161 source.n145 0.155672
R524 source.n162 source.n161 0.155672
R525 source.n162 source.n141 0.155672
R526 source.n169 source.n141 0.155672
R527 source.n29 source.n1 0.155672
R528 source.n22 source.n1 0.155672
R529 source.n22 source.n21 0.155672
R530 source.n21 source.n5 0.155672
R531 source.n14 source.n5 0.155672
R532 source.n14 source.n13 0.155672
R533 source.n67 source.n39 0.155672
R534 source.n60 source.n39 0.155672
R535 source.n60 source.n59 0.155672
R536 source.n59 source.n43 0.155672
R537 source.n52 source.n43 0.155672
R538 source.n52 source.n51 0.155672
R539 source.n99 source.n71 0.155672
R540 source.n92 source.n71 0.155672
R541 source.n92 source.n91 0.155672
R542 source.n91 source.n75 0.155672
R543 source.n84 source.n75 0.155672
R544 source.n84 source.n83 0.155672
R545 source.n137 source.n109 0.155672
R546 source.n130 source.n109 0.155672
R547 source.n130 source.n129 0.155672
R548 source.n129 source.n113 0.155672
R549 source.n122 source.n113 0.155672
R550 source.n122 source.n121 0.155672
R551 plus.n5 plus.t2 616.376
R552 plus.n21 plus.t0 616.376
R553 plus.n28 plus.t8 616.376
R554 plus.n44 plus.t5 616.376
R555 plus.n6 plus.t7 586.433
R556 plus.n3 plus.t11 586.433
R557 plus.n12 plus.t15 586.433
R558 plus.n14 plus.t6 586.433
R559 plus.n1 plus.t10 586.433
R560 plus.n20 plus.t14 586.433
R561 plus.n29 plus.t1 586.433
R562 plus.n26 plus.t9 586.433
R563 plus.n35 plus.t3 586.433
R564 plus.n37 plus.t12 586.433
R565 plus.n24 plus.t4 586.433
R566 plus.n43 plus.t13 586.433
R567 plus.n5 plus.n4 161.489
R568 plus.n28 plus.n27 161.489
R569 plus.n7 plus.n4 161.3
R570 plus.n9 plus.n8 161.3
R571 plus.n11 plus.n10 161.3
R572 plus.n13 plus.n2 161.3
R573 plus.n16 plus.n15 161.3
R574 plus.n18 plus.n17 161.3
R575 plus.n19 plus.n0 161.3
R576 plus.n22 plus.n21 161.3
R577 plus.n30 plus.n27 161.3
R578 plus.n32 plus.n31 161.3
R579 plus.n34 plus.n33 161.3
R580 plus.n36 plus.n25 161.3
R581 plus.n39 plus.n38 161.3
R582 plus.n41 plus.n40 161.3
R583 plus.n42 plus.n23 161.3
R584 plus.n45 plus.n44 161.3
R585 plus.n8 plus.n7 73.0308
R586 plus.n19 plus.n18 73.0308
R587 plus.n42 plus.n41 73.0308
R588 plus.n31 plus.n30 73.0308
R589 plus.n11 plus.n3 64.9975
R590 plus.n15 plus.n1 64.9975
R591 plus.n38 plus.n24 64.9975
R592 plus.n34 plus.n26 64.9975
R593 plus.n6 plus.n5 62.0763
R594 plus.n21 plus.n20 62.0763
R595 plus.n44 plus.n43 62.0763
R596 plus.n29 plus.n28 62.0763
R597 plus.n13 plus.n12 46.0096
R598 plus.n14 plus.n13 46.0096
R599 plus.n37 plus.n36 46.0096
R600 plus.n36 plus.n35 46.0096
R601 plus plus.n45 27.7036
R602 plus.n12 plus.n11 27.0217
R603 plus.n15 plus.n14 27.0217
R604 plus.n38 plus.n37 27.0217
R605 plus.n35 plus.n34 27.0217
R606 plus.n7 plus.n6 10.955
R607 plus.n20 plus.n19 10.955
R608 plus.n43 plus.n42 10.955
R609 plus.n30 plus.n29 10.955
R610 plus plus.n22 9.83762
R611 plus.n8 plus.n3 8.03383
R612 plus.n18 plus.n1 8.03383
R613 plus.n41 plus.n24 8.03383
R614 plus.n31 plus.n26 8.03383
R615 plus.n9 plus.n4 0.189894
R616 plus.n10 plus.n9 0.189894
R617 plus.n10 plus.n2 0.189894
R618 plus.n16 plus.n2 0.189894
R619 plus.n17 plus.n16 0.189894
R620 plus.n17 plus.n0 0.189894
R621 plus.n22 plus.n0 0.189894
R622 plus.n45 plus.n23 0.189894
R623 plus.n40 plus.n23 0.189894
R624 plus.n40 plus.n39 0.189894
R625 plus.n39 plus.n25 0.189894
R626 plus.n33 plus.n25 0.189894
R627 plus.n33 plus.n32 0.189894
R628 plus.n32 plus.n27 0.189894
R629 drain_left.n9 drain_left.n7 67.7339
R630 drain_left.n5 drain_left.n3 67.7338
R631 drain_left.n2 drain_left.n0 67.7338
R632 drain_left.n11 drain_left.n10 67.1908
R633 drain_left.n9 drain_left.n8 67.1908
R634 drain_left.n13 drain_left.n12 67.1907
R635 drain_left.n5 drain_left.n4 67.1907
R636 drain_left.n2 drain_left.n1 67.1907
R637 drain_left drain_left.n6 26.3518
R638 drain_left drain_left.n13 6.19632
R639 drain_left.n3 drain_left.t14 3.3005
R640 drain_left.n3 drain_left.t7 3.3005
R641 drain_left.n4 drain_left.t12 3.3005
R642 drain_left.n4 drain_left.t6 3.3005
R643 drain_left.n1 drain_left.t11 3.3005
R644 drain_left.n1 drain_left.t3 3.3005
R645 drain_left.n0 drain_left.t10 3.3005
R646 drain_left.n0 drain_left.t2 3.3005
R647 drain_left.n12 drain_left.t1 3.3005
R648 drain_left.n12 drain_left.t15 3.3005
R649 drain_left.n10 drain_left.t9 3.3005
R650 drain_left.n10 drain_left.t5 3.3005
R651 drain_left.n8 drain_left.t4 3.3005
R652 drain_left.n8 drain_left.t0 3.3005
R653 drain_left.n7 drain_left.t13 3.3005
R654 drain_left.n7 drain_left.t8 3.3005
R655 drain_left.n11 drain_left.n9 0.543603
R656 drain_left.n13 drain_left.n11 0.543603
R657 drain_left.n6 drain_left.n5 0.216706
R658 drain_left.n6 drain_left.n2 0.216706
C0 drain_left drain_right 0.948737f
C1 plus source 3.22402f
C2 minus drain_right 3.20734f
C3 plus drain_left 3.38704f
C4 drain_left source 16.659399f
C5 plus minus 4.35198f
C6 minus source 3.21f
C7 minus drain_left 0.171647f
C8 plus drain_right 0.334364f
C9 source drain_right 16.6596f
C10 drain_right a_n1850_n2088# 5.221429f
C11 drain_left a_n1850_n2088# 5.51257f
C12 source a_n1850_n2088# 5.341278f
C13 minus a_n1850_n2088# 6.756336f
C14 plus a_n1850_n2088# 8.35171f
C15 drain_left.t10 a_n1850_n2088# 0.158181f
C16 drain_left.t2 a_n1850_n2088# 0.158181f
C17 drain_left.n0 a_n1850_n2088# 1.32244f
C18 drain_left.t11 a_n1850_n2088# 0.158181f
C19 drain_left.t3 a_n1850_n2088# 0.158181f
C20 drain_left.n1 a_n1850_n2088# 1.31923f
C21 drain_left.n2 a_n1850_n2088# 0.753742f
C22 drain_left.t14 a_n1850_n2088# 0.158181f
C23 drain_left.t7 a_n1850_n2088# 0.158181f
C24 drain_left.n3 a_n1850_n2088# 1.32244f
C25 drain_left.t12 a_n1850_n2088# 0.158181f
C26 drain_left.t6 a_n1850_n2088# 0.158181f
C27 drain_left.n4 a_n1850_n2088# 1.31923f
C28 drain_left.n5 a_n1850_n2088# 0.753742f
C29 drain_left.n6 a_n1850_n2088# 1.20031f
C30 drain_left.t13 a_n1850_n2088# 0.158181f
C31 drain_left.t8 a_n1850_n2088# 0.158181f
C32 drain_left.n7 a_n1850_n2088# 1.32245f
C33 drain_left.t4 a_n1850_n2088# 0.158181f
C34 drain_left.t0 a_n1850_n2088# 0.158181f
C35 drain_left.n8 a_n1850_n2088# 1.31923f
C36 drain_left.n9 a_n1850_n2088# 0.785293f
C37 drain_left.t9 a_n1850_n2088# 0.158181f
C38 drain_left.t5 a_n1850_n2088# 0.158181f
C39 drain_left.n10 a_n1850_n2088# 1.31923f
C40 drain_left.n11 a_n1850_n2088# 0.387535f
C41 drain_left.t1 a_n1850_n2088# 0.158181f
C42 drain_left.t15 a_n1850_n2088# 0.158181f
C43 drain_left.n12 a_n1850_n2088# 1.31923f
C44 drain_left.n13 a_n1850_n2088# 0.665232f
C45 plus.n0 a_n1850_n2088# 0.052058f
C46 plus.t14 a_n1850_n2088# 0.266982f
C47 plus.t10 a_n1850_n2088# 0.266982f
C48 plus.n1 a_n1850_n2088# 0.122549f
C49 plus.n2 a_n1850_n2088# 0.052058f
C50 plus.t6 a_n1850_n2088# 0.266982f
C51 plus.t15 a_n1850_n2088# 0.266982f
C52 plus.t11 a_n1850_n2088# 0.266982f
C53 plus.n3 a_n1850_n2088# 0.122549f
C54 plus.n4 a_n1850_n2088# 0.110788f
C55 plus.t7 a_n1850_n2088# 0.266982f
C56 plus.t2 a_n1850_n2088# 0.272943f
C57 plus.n5 a_n1850_n2088# 0.13826f
C58 plus.n6 a_n1850_n2088# 0.122549f
C59 plus.n7 a_n1850_n2088# 0.019677f
C60 plus.n8 a_n1850_n2088# 0.019035f
C61 plus.n9 a_n1850_n2088# 0.052058f
C62 plus.n10 a_n1850_n2088# 0.052058f
C63 plus.n11 a_n1850_n2088# 0.021442f
C64 plus.n12 a_n1850_n2088# 0.122549f
C65 plus.n13 a_n1850_n2088# 0.021442f
C66 plus.n14 a_n1850_n2088# 0.122549f
C67 plus.n15 a_n1850_n2088# 0.021442f
C68 plus.n16 a_n1850_n2088# 0.052058f
C69 plus.n17 a_n1850_n2088# 0.052058f
C70 plus.n18 a_n1850_n2088# 0.019035f
C71 plus.n19 a_n1850_n2088# 0.019677f
C72 plus.n20 a_n1850_n2088# 0.122549f
C73 plus.t0 a_n1850_n2088# 0.272943f
C74 plus.n21 a_n1850_n2088# 0.138191f
C75 plus.n22 a_n1850_n2088# 0.441783f
C76 plus.n23 a_n1850_n2088# 0.052058f
C77 plus.t5 a_n1850_n2088# 0.272943f
C78 plus.t13 a_n1850_n2088# 0.266982f
C79 plus.t4 a_n1850_n2088# 0.266982f
C80 plus.n24 a_n1850_n2088# 0.122549f
C81 plus.n25 a_n1850_n2088# 0.052058f
C82 plus.t12 a_n1850_n2088# 0.266982f
C83 plus.t3 a_n1850_n2088# 0.266982f
C84 plus.t9 a_n1850_n2088# 0.266982f
C85 plus.n26 a_n1850_n2088# 0.122549f
C86 plus.n27 a_n1850_n2088# 0.110788f
C87 plus.t1 a_n1850_n2088# 0.266982f
C88 plus.t8 a_n1850_n2088# 0.272943f
C89 plus.n28 a_n1850_n2088# 0.13826f
C90 plus.n29 a_n1850_n2088# 0.122549f
C91 plus.n30 a_n1850_n2088# 0.019677f
C92 plus.n31 a_n1850_n2088# 0.019035f
C93 plus.n32 a_n1850_n2088# 0.052058f
C94 plus.n33 a_n1850_n2088# 0.052058f
C95 plus.n34 a_n1850_n2088# 0.021442f
C96 plus.n35 a_n1850_n2088# 0.122549f
C97 plus.n36 a_n1850_n2088# 0.021442f
C98 plus.n37 a_n1850_n2088# 0.122549f
C99 plus.n38 a_n1850_n2088# 0.021442f
C100 plus.n39 a_n1850_n2088# 0.052058f
C101 plus.n40 a_n1850_n2088# 0.052058f
C102 plus.n41 a_n1850_n2088# 0.019035f
C103 plus.n42 a_n1850_n2088# 0.019677f
C104 plus.n43 a_n1850_n2088# 0.122549f
C105 plus.n44 a_n1850_n2088# 0.138191f
C106 plus.n45 a_n1850_n2088# 1.33003f
C107 source.n0 a_n1850_n2088# 0.041572f
C108 source.n1 a_n1850_n2088# 0.029577f
C109 source.n2 a_n1850_n2088# 0.015893f
C110 source.n3 a_n1850_n2088# 0.037565f
C111 source.n4 a_n1850_n2088# 0.016828f
C112 source.n5 a_n1850_n2088# 0.029577f
C113 source.n6 a_n1850_n2088# 0.015893f
C114 source.n7 a_n1850_n2088# 0.037565f
C115 source.n8 a_n1850_n2088# 0.016828f
C116 source.n9 a_n1850_n2088# 0.126566f
C117 source.t0 a_n1850_n2088# 0.061227f
C118 source.n10 a_n1850_n2088# 0.028174f
C119 source.n11 a_n1850_n2088# 0.02219f
C120 source.n12 a_n1850_n2088# 0.015893f
C121 source.n13 a_n1850_n2088# 0.703743f
C122 source.n14 a_n1850_n2088# 0.029577f
C123 source.n15 a_n1850_n2088# 0.015893f
C124 source.n16 a_n1850_n2088# 0.016828f
C125 source.n17 a_n1850_n2088# 0.037565f
C126 source.n18 a_n1850_n2088# 0.037565f
C127 source.n19 a_n1850_n2088# 0.016828f
C128 source.n20 a_n1850_n2088# 0.015893f
C129 source.n21 a_n1850_n2088# 0.029577f
C130 source.n22 a_n1850_n2088# 0.029577f
C131 source.n23 a_n1850_n2088# 0.015893f
C132 source.n24 a_n1850_n2088# 0.016828f
C133 source.n25 a_n1850_n2088# 0.037565f
C134 source.n26 a_n1850_n2088# 0.081323f
C135 source.n27 a_n1850_n2088# 0.016828f
C136 source.n28 a_n1850_n2088# 0.015893f
C137 source.n29 a_n1850_n2088# 0.068365f
C138 source.n30 a_n1850_n2088# 0.045503f
C139 source.n31 a_n1850_n2088# 0.716401f
C140 source.t4 a_n1850_n2088# 0.140233f
C141 source.t13 a_n1850_n2088# 0.140233f
C142 source.n32 a_n1850_n2088# 1.09215f
C143 source.n33 a_n1850_n2088# 0.380768f
C144 source.t8 a_n1850_n2088# 0.140233f
C145 source.t15 a_n1850_n2088# 0.140233f
C146 source.n34 a_n1850_n2088# 1.09215f
C147 source.n35 a_n1850_n2088# 0.380768f
C148 source.t7 a_n1850_n2088# 0.140233f
C149 source.t1 a_n1850_n2088# 0.140233f
C150 source.n36 a_n1850_n2088# 1.09215f
C151 source.n37 a_n1850_n2088# 0.380768f
C152 source.n38 a_n1850_n2088# 0.041572f
C153 source.n39 a_n1850_n2088# 0.029577f
C154 source.n40 a_n1850_n2088# 0.015893f
C155 source.n41 a_n1850_n2088# 0.037565f
C156 source.n42 a_n1850_n2088# 0.016828f
C157 source.n43 a_n1850_n2088# 0.029577f
C158 source.n44 a_n1850_n2088# 0.015893f
C159 source.n45 a_n1850_n2088# 0.037565f
C160 source.n46 a_n1850_n2088# 0.016828f
C161 source.n47 a_n1850_n2088# 0.126566f
C162 source.t2 a_n1850_n2088# 0.061227f
C163 source.n48 a_n1850_n2088# 0.028174f
C164 source.n49 a_n1850_n2088# 0.02219f
C165 source.n50 a_n1850_n2088# 0.015893f
C166 source.n51 a_n1850_n2088# 0.703743f
C167 source.n52 a_n1850_n2088# 0.029577f
C168 source.n53 a_n1850_n2088# 0.015893f
C169 source.n54 a_n1850_n2088# 0.016828f
C170 source.n55 a_n1850_n2088# 0.037565f
C171 source.n56 a_n1850_n2088# 0.037565f
C172 source.n57 a_n1850_n2088# 0.016828f
C173 source.n58 a_n1850_n2088# 0.015893f
C174 source.n59 a_n1850_n2088# 0.029577f
C175 source.n60 a_n1850_n2088# 0.029577f
C176 source.n61 a_n1850_n2088# 0.015893f
C177 source.n62 a_n1850_n2088# 0.016828f
C178 source.n63 a_n1850_n2088# 0.037565f
C179 source.n64 a_n1850_n2088# 0.081323f
C180 source.n65 a_n1850_n2088# 0.016828f
C181 source.n66 a_n1850_n2088# 0.015893f
C182 source.n67 a_n1850_n2088# 0.068365f
C183 source.n68 a_n1850_n2088# 0.045503f
C184 source.n69 a_n1850_n2088# 0.121795f
C185 source.n70 a_n1850_n2088# 0.041572f
C186 source.n71 a_n1850_n2088# 0.029577f
C187 source.n72 a_n1850_n2088# 0.015893f
C188 source.n73 a_n1850_n2088# 0.037565f
C189 source.n74 a_n1850_n2088# 0.016828f
C190 source.n75 a_n1850_n2088# 0.029577f
C191 source.n76 a_n1850_n2088# 0.015893f
C192 source.n77 a_n1850_n2088# 0.037565f
C193 source.n78 a_n1850_n2088# 0.016828f
C194 source.n79 a_n1850_n2088# 0.126566f
C195 source.t21 a_n1850_n2088# 0.061227f
C196 source.n80 a_n1850_n2088# 0.028174f
C197 source.n81 a_n1850_n2088# 0.02219f
C198 source.n82 a_n1850_n2088# 0.015893f
C199 source.n83 a_n1850_n2088# 0.703743f
C200 source.n84 a_n1850_n2088# 0.029577f
C201 source.n85 a_n1850_n2088# 0.015893f
C202 source.n86 a_n1850_n2088# 0.016828f
C203 source.n87 a_n1850_n2088# 0.037565f
C204 source.n88 a_n1850_n2088# 0.037565f
C205 source.n89 a_n1850_n2088# 0.016828f
C206 source.n90 a_n1850_n2088# 0.015893f
C207 source.n91 a_n1850_n2088# 0.029577f
C208 source.n92 a_n1850_n2088# 0.029577f
C209 source.n93 a_n1850_n2088# 0.015893f
C210 source.n94 a_n1850_n2088# 0.016828f
C211 source.n95 a_n1850_n2088# 0.037565f
C212 source.n96 a_n1850_n2088# 0.081323f
C213 source.n97 a_n1850_n2088# 0.016828f
C214 source.n98 a_n1850_n2088# 0.015893f
C215 source.n99 a_n1850_n2088# 0.068365f
C216 source.n100 a_n1850_n2088# 0.045503f
C217 source.n101 a_n1850_n2088# 0.121795f
C218 source.t28 a_n1850_n2088# 0.140233f
C219 source.t17 a_n1850_n2088# 0.140233f
C220 source.n102 a_n1850_n2088# 1.09215f
C221 source.n103 a_n1850_n2088# 0.380768f
C222 source.t18 a_n1850_n2088# 0.140233f
C223 source.t22 a_n1850_n2088# 0.140233f
C224 source.n104 a_n1850_n2088# 1.09215f
C225 source.n105 a_n1850_n2088# 0.380768f
C226 source.t27 a_n1850_n2088# 0.140233f
C227 source.t29 a_n1850_n2088# 0.140233f
C228 source.n106 a_n1850_n2088# 1.09215f
C229 source.n107 a_n1850_n2088# 0.380768f
C230 source.n108 a_n1850_n2088# 0.041572f
C231 source.n109 a_n1850_n2088# 0.029577f
C232 source.n110 a_n1850_n2088# 0.015893f
C233 source.n111 a_n1850_n2088# 0.037565f
C234 source.n112 a_n1850_n2088# 0.016828f
C235 source.n113 a_n1850_n2088# 0.029577f
C236 source.n114 a_n1850_n2088# 0.015893f
C237 source.n115 a_n1850_n2088# 0.037565f
C238 source.n116 a_n1850_n2088# 0.016828f
C239 source.n117 a_n1850_n2088# 0.126566f
C240 source.t16 a_n1850_n2088# 0.061227f
C241 source.n118 a_n1850_n2088# 0.028174f
C242 source.n119 a_n1850_n2088# 0.02219f
C243 source.n120 a_n1850_n2088# 0.015893f
C244 source.n121 a_n1850_n2088# 0.703743f
C245 source.n122 a_n1850_n2088# 0.029577f
C246 source.n123 a_n1850_n2088# 0.015893f
C247 source.n124 a_n1850_n2088# 0.016828f
C248 source.n125 a_n1850_n2088# 0.037565f
C249 source.n126 a_n1850_n2088# 0.037565f
C250 source.n127 a_n1850_n2088# 0.016828f
C251 source.n128 a_n1850_n2088# 0.015893f
C252 source.n129 a_n1850_n2088# 0.029577f
C253 source.n130 a_n1850_n2088# 0.029577f
C254 source.n131 a_n1850_n2088# 0.015893f
C255 source.n132 a_n1850_n2088# 0.016828f
C256 source.n133 a_n1850_n2088# 0.037565f
C257 source.n134 a_n1850_n2088# 0.081323f
C258 source.n135 a_n1850_n2088# 0.016828f
C259 source.n136 a_n1850_n2088# 0.015893f
C260 source.n137 a_n1850_n2088# 0.068365f
C261 source.n138 a_n1850_n2088# 0.045503f
C262 source.n139 a_n1850_n2088# 1.09717f
C263 source.n140 a_n1850_n2088# 0.041572f
C264 source.n141 a_n1850_n2088# 0.029577f
C265 source.n142 a_n1850_n2088# 0.015893f
C266 source.n143 a_n1850_n2088# 0.037565f
C267 source.n144 a_n1850_n2088# 0.016828f
C268 source.n145 a_n1850_n2088# 0.029577f
C269 source.n146 a_n1850_n2088# 0.015893f
C270 source.n147 a_n1850_n2088# 0.037565f
C271 source.n148 a_n1850_n2088# 0.016828f
C272 source.n149 a_n1850_n2088# 0.126566f
C273 source.t6 a_n1850_n2088# 0.061227f
C274 source.n150 a_n1850_n2088# 0.028174f
C275 source.n151 a_n1850_n2088# 0.02219f
C276 source.n152 a_n1850_n2088# 0.015893f
C277 source.n153 a_n1850_n2088# 0.703743f
C278 source.n154 a_n1850_n2088# 0.029577f
C279 source.n155 a_n1850_n2088# 0.015893f
C280 source.n156 a_n1850_n2088# 0.016828f
C281 source.n157 a_n1850_n2088# 0.037565f
C282 source.n158 a_n1850_n2088# 0.037565f
C283 source.n159 a_n1850_n2088# 0.016828f
C284 source.n160 a_n1850_n2088# 0.015893f
C285 source.n161 a_n1850_n2088# 0.029577f
C286 source.n162 a_n1850_n2088# 0.029577f
C287 source.n163 a_n1850_n2088# 0.015893f
C288 source.n164 a_n1850_n2088# 0.016828f
C289 source.n165 a_n1850_n2088# 0.037565f
C290 source.n166 a_n1850_n2088# 0.081323f
C291 source.n167 a_n1850_n2088# 0.016828f
C292 source.n168 a_n1850_n2088# 0.015893f
C293 source.n169 a_n1850_n2088# 0.068365f
C294 source.n170 a_n1850_n2088# 0.045503f
C295 source.n171 a_n1850_n2088# 1.09717f
C296 source.t5 a_n1850_n2088# 0.140233f
C297 source.t11 a_n1850_n2088# 0.140233f
C298 source.n172 a_n1850_n2088# 1.09214f
C299 source.n173 a_n1850_n2088# 0.380776f
C300 source.t3 a_n1850_n2088# 0.140233f
C301 source.t9 a_n1850_n2088# 0.140233f
C302 source.n174 a_n1850_n2088# 1.09214f
C303 source.n175 a_n1850_n2088# 0.380776f
C304 source.t12 a_n1850_n2088# 0.140233f
C305 source.t14 a_n1850_n2088# 0.140233f
C306 source.n176 a_n1850_n2088# 1.09214f
C307 source.n177 a_n1850_n2088# 0.380776f
C308 source.n178 a_n1850_n2088# 0.041572f
C309 source.n179 a_n1850_n2088# 0.029577f
C310 source.n180 a_n1850_n2088# 0.015893f
C311 source.n181 a_n1850_n2088# 0.037565f
C312 source.n182 a_n1850_n2088# 0.016828f
C313 source.n183 a_n1850_n2088# 0.029577f
C314 source.n184 a_n1850_n2088# 0.015893f
C315 source.n185 a_n1850_n2088# 0.037565f
C316 source.n186 a_n1850_n2088# 0.016828f
C317 source.n187 a_n1850_n2088# 0.126566f
C318 source.t10 a_n1850_n2088# 0.061227f
C319 source.n188 a_n1850_n2088# 0.028174f
C320 source.n189 a_n1850_n2088# 0.02219f
C321 source.n190 a_n1850_n2088# 0.015893f
C322 source.n191 a_n1850_n2088# 0.703743f
C323 source.n192 a_n1850_n2088# 0.029577f
C324 source.n193 a_n1850_n2088# 0.015893f
C325 source.n194 a_n1850_n2088# 0.016828f
C326 source.n195 a_n1850_n2088# 0.037565f
C327 source.n196 a_n1850_n2088# 0.037565f
C328 source.n197 a_n1850_n2088# 0.016828f
C329 source.n198 a_n1850_n2088# 0.015893f
C330 source.n199 a_n1850_n2088# 0.029577f
C331 source.n200 a_n1850_n2088# 0.029577f
C332 source.n201 a_n1850_n2088# 0.015893f
C333 source.n202 a_n1850_n2088# 0.016828f
C334 source.n203 a_n1850_n2088# 0.037565f
C335 source.n204 a_n1850_n2088# 0.081323f
C336 source.n205 a_n1850_n2088# 0.016828f
C337 source.n206 a_n1850_n2088# 0.015893f
C338 source.n207 a_n1850_n2088# 0.068365f
C339 source.n208 a_n1850_n2088# 0.045503f
C340 source.n209 a_n1850_n2088# 0.121795f
C341 source.n210 a_n1850_n2088# 0.041572f
C342 source.n211 a_n1850_n2088# 0.029577f
C343 source.n212 a_n1850_n2088# 0.015893f
C344 source.n213 a_n1850_n2088# 0.037565f
C345 source.n214 a_n1850_n2088# 0.016828f
C346 source.n215 a_n1850_n2088# 0.029577f
C347 source.n216 a_n1850_n2088# 0.015893f
C348 source.n217 a_n1850_n2088# 0.037565f
C349 source.n218 a_n1850_n2088# 0.016828f
C350 source.n219 a_n1850_n2088# 0.126566f
C351 source.t19 a_n1850_n2088# 0.061227f
C352 source.n220 a_n1850_n2088# 0.028174f
C353 source.n221 a_n1850_n2088# 0.02219f
C354 source.n222 a_n1850_n2088# 0.015893f
C355 source.n223 a_n1850_n2088# 0.703743f
C356 source.n224 a_n1850_n2088# 0.029577f
C357 source.n225 a_n1850_n2088# 0.015893f
C358 source.n226 a_n1850_n2088# 0.016828f
C359 source.n227 a_n1850_n2088# 0.037565f
C360 source.n228 a_n1850_n2088# 0.037565f
C361 source.n229 a_n1850_n2088# 0.016828f
C362 source.n230 a_n1850_n2088# 0.015893f
C363 source.n231 a_n1850_n2088# 0.029577f
C364 source.n232 a_n1850_n2088# 0.029577f
C365 source.n233 a_n1850_n2088# 0.015893f
C366 source.n234 a_n1850_n2088# 0.016828f
C367 source.n235 a_n1850_n2088# 0.037565f
C368 source.n236 a_n1850_n2088# 0.081323f
C369 source.n237 a_n1850_n2088# 0.016828f
C370 source.n238 a_n1850_n2088# 0.015893f
C371 source.n239 a_n1850_n2088# 0.068365f
C372 source.n240 a_n1850_n2088# 0.045503f
C373 source.n241 a_n1850_n2088# 0.121795f
C374 source.t25 a_n1850_n2088# 0.140233f
C375 source.t20 a_n1850_n2088# 0.140233f
C376 source.n242 a_n1850_n2088# 1.09214f
C377 source.n243 a_n1850_n2088# 0.380776f
C378 source.t26 a_n1850_n2088# 0.140233f
C379 source.t30 a_n1850_n2088# 0.140233f
C380 source.n244 a_n1850_n2088# 1.09214f
C381 source.n245 a_n1850_n2088# 0.380776f
C382 source.t23 a_n1850_n2088# 0.140233f
C383 source.t31 a_n1850_n2088# 0.140233f
C384 source.n246 a_n1850_n2088# 1.09214f
C385 source.n247 a_n1850_n2088# 0.380776f
C386 source.n248 a_n1850_n2088# 0.041572f
C387 source.n249 a_n1850_n2088# 0.029577f
C388 source.n250 a_n1850_n2088# 0.015893f
C389 source.n251 a_n1850_n2088# 0.037565f
C390 source.n252 a_n1850_n2088# 0.016828f
C391 source.n253 a_n1850_n2088# 0.029577f
C392 source.n254 a_n1850_n2088# 0.015893f
C393 source.n255 a_n1850_n2088# 0.037565f
C394 source.n256 a_n1850_n2088# 0.016828f
C395 source.n257 a_n1850_n2088# 0.126566f
C396 source.t24 a_n1850_n2088# 0.061227f
C397 source.n258 a_n1850_n2088# 0.028174f
C398 source.n259 a_n1850_n2088# 0.02219f
C399 source.n260 a_n1850_n2088# 0.015893f
C400 source.n261 a_n1850_n2088# 0.703743f
C401 source.n262 a_n1850_n2088# 0.029577f
C402 source.n263 a_n1850_n2088# 0.015893f
C403 source.n264 a_n1850_n2088# 0.016828f
C404 source.n265 a_n1850_n2088# 0.037565f
C405 source.n266 a_n1850_n2088# 0.037565f
C406 source.n267 a_n1850_n2088# 0.016828f
C407 source.n268 a_n1850_n2088# 0.015893f
C408 source.n269 a_n1850_n2088# 0.029577f
C409 source.n270 a_n1850_n2088# 0.029577f
C410 source.n271 a_n1850_n2088# 0.015893f
C411 source.n272 a_n1850_n2088# 0.016828f
C412 source.n273 a_n1850_n2088# 0.037565f
C413 source.n274 a_n1850_n2088# 0.081323f
C414 source.n275 a_n1850_n2088# 0.016828f
C415 source.n276 a_n1850_n2088# 0.015893f
C416 source.n277 a_n1850_n2088# 0.068365f
C417 source.n278 a_n1850_n2088# 0.045503f
C418 source.n279 a_n1850_n2088# 0.288754f
C419 source.n280 a_n1850_n2088# 1.21022f
C420 drain_right.t1 a_n1850_n2088# 0.15763f
C421 drain_right.t2 a_n1850_n2088# 0.15763f
C422 drain_right.n0 a_n1850_n2088# 1.31784f
C423 drain_right.t3 a_n1850_n2088# 0.15763f
C424 drain_right.t0 a_n1850_n2088# 0.15763f
C425 drain_right.n1 a_n1850_n2088# 1.31464f
C426 drain_right.n2 a_n1850_n2088# 0.751119f
C427 drain_right.t4 a_n1850_n2088# 0.15763f
C428 drain_right.t13 a_n1850_n2088# 0.15763f
C429 drain_right.n3 a_n1850_n2088# 1.31784f
C430 drain_right.t11 a_n1850_n2088# 0.15763f
C431 drain_right.t10 a_n1850_n2088# 0.15763f
C432 drain_right.n4 a_n1850_n2088# 1.31464f
C433 drain_right.n5 a_n1850_n2088# 0.751119f
C434 drain_right.n6 a_n1850_n2088# 1.12866f
C435 drain_right.t15 a_n1850_n2088# 0.15763f
C436 drain_right.t5 a_n1850_n2088# 0.15763f
C437 drain_right.n7 a_n1850_n2088# 1.31784f
C438 drain_right.t9 a_n1850_n2088# 0.15763f
C439 drain_right.t6 a_n1850_n2088# 0.15763f
C440 drain_right.n8 a_n1850_n2088# 1.31464f
C441 drain_right.n9 a_n1850_n2088# 0.782566f
C442 drain_right.t7 a_n1850_n2088# 0.15763f
C443 drain_right.t8 a_n1850_n2088# 0.15763f
C444 drain_right.n10 a_n1850_n2088# 1.31464f
C445 drain_right.n11 a_n1850_n2088# 0.386187f
C446 drain_right.t14 a_n1850_n2088# 0.15763f
C447 drain_right.t12 a_n1850_n2088# 0.15763f
C448 drain_right.n12 a_n1850_n2088# 1.31464f
C449 drain_right.n13 a_n1850_n2088# 0.66291f
C450 minus.n0 a_n1850_n2088# 0.050627f
C451 minus.t15 a_n1850_n2088# 0.26544f
C452 minus.t4 a_n1850_n2088# 0.259643f
C453 minus.t2 a_n1850_n2088# 0.259643f
C454 minus.n1 a_n1850_n2088# 0.11918f
C455 minus.n2 a_n1850_n2088# 0.050627f
C456 minus.t13 a_n1850_n2088# 0.259643f
C457 minus.t9 a_n1850_n2088# 0.259643f
C458 minus.t3 a_n1850_n2088# 0.259643f
C459 minus.n3 a_n1850_n2088# 0.11918f
C460 minus.n4 a_n1850_n2088# 0.107743f
C461 minus.t14 a_n1850_n2088# 0.259643f
C462 minus.t10 a_n1850_n2088# 0.26544f
C463 minus.n5 a_n1850_n2088# 0.134459f
C464 minus.n6 a_n1850_n2088# 0.11918f
C465 minus.n7 a_n1850_n2088# 0.019136f
C466 minus.n8 a_n1850_n2088# 0.018512f
C467 minus.n9 a_n1850_n2088# 0.050627f
C468 minus.n10 a_n1850_n2088# 0.050627f
C469 minus.n11 a_n1850_n2088# 0.020853f
C470 minus.n12 a_n1850_n2088# 0.11918f
C471 minus.n13 a_n1850_n2088# 0.020853f
C472 minus.n14 a_n1850_n2088# 0.11918f
C473 minus.n15 a_n1850_n2088# 0.020853f
C474 minus.n16 a_n1850_n2088# 0.050627f
C475 minus.n17 a_n1850_n2088# 0.050627f
C476 minus.n18 a_n1850_n2088# 0.018512f
C477 minus.n19 a_n1850_n2088# 0.019136f
C478 minus.n20 a_n1850_n2088# 0.11918f
C479 minus.n21 a_n1850_n2088# 0.134392f
C480 minus.n22 a_n1850_n2088# 1.43227f
C481 minus.n23 a_n1850_n2088# 0.050627f
C482 minus.t0 a_n1850_n2088# 0.259643f
C483 minus.t8 a_n1850_n2088# 0.259643f
C484 minus.n24 a_n1850_n2088# 0.11918f
C485 minus.n25 a_n1850_n2088# 0.050627f
C486 minus.t1 a_n1850_n2088# 0.259643f
C487 minus.t5 a_n1850_n2088# 0.259643f
C488 minus.t11 a_n1850_n2088# 0.259643f
C489 minus.n26 a_n1850_n2088# 0.11918f
C490 minus.n27 a_n1850_n2088# 0.107743f
C491 minus.t6 a_n1850_n2088# 0.259643f
C492 minus.t12 a_n1850_n2088# 0.26544f
C493 minus.n28 a_n1850_n2088# 0.134459f
C494 minus.n29 a_n1850_n2088# 0.11918f
C495 minus.n30 a_n1850_n2088# 0.019136f
C496 minus.n31 a_n1850_n2088# 0.018512f
C497 minus.n32 a_n1850_n2088# 0.050627f
C498 minus.n33 a_n1850_n2088# 0.050627f
C499 minus.n34 a_n1850_n2088# 0.020853f
C500 minus.n35 a_n1850_n2088# 0.11918f
C501 minus.n36 a_n1850_n2088# 0.020853f
C502 minus.n37 a_n1850_n2088# 0.11918f
C503 minus.n38 a_n1850_n2088# 0.020853f
C504 minus.n39 a_n1850_n2088# 0.050627f
C505 minus.n40 a_n1850_n2088# 0.050627f
C506 minus.n41 a_n1850_n2088# 0.018512f
C507 minus.n42 a_n1850_n2088# 0.019136f
C508 minus.n43 a_n1850_n2088# 0.11918f
C509 minus.t7 a_n1850_n2088# 0.26544f
C510 minus.n44 a_n1850_n2088# 0.134392f
C511 minus.n45 a_n1850_n2088# 0.326976f
C512 minus.n46 a_n1850_n2088# 1.76345f
.ends

