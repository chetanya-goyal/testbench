* NGSPICE file created from diffpair440.ext - technology: sky130A

.subckt diffpair440 minus drain_right drain_left source plus
X0 drain_right minus source a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X1 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.5
X2 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X3 drain_left plus source a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X4 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X5 drain_right minus source a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X6 drain_left plus source a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.5
X7 a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# a_n1048_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
.ends

