* NGSPICE file created from diffpair535.ext - technology: sky130A

.subckt diffpair535 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t12 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X1 drain_left.t11 plus.t0 source.t4 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X2 source.t6 plus.t1 drain_left.t10 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X3 drain_left.t9 plus.t2 source.t2 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X4 drain_right.t10 minus.t1 source.t11 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X5 drain_right.t9 minus.t2 source.t19 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X6 source.t16 minus.t3 drain_right.t8 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X7 drain_left.t8 plus.t3 source.t20 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X8 source.t10 minus.t4 drain_right.t7 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X9 drain_right.t6 minus.t5 source.t17 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X10 source.t21 plus.t4 drain_left.t7 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X11 source.t22 plus.t5 drain_left.t6 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X12 source.t8 minus.t6 drain_right.t5 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X13 drain_right.t4 minus.t7 source.t14 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X14 source.t18 minus.t8 drain_right.t3 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X15 source.t23 plus.t6 drain_left.t5 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X16 drain_left.t4 plus.t7 source.t1 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X17 source.t15 minus.t9 drain_right.t2 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X18 source.t0 plus.t8 drain_left.t3 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X19 drain_right.t1 minus.t10 source.t13 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.6
X20 a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.6
X21 a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X22 drain_left.t2 plus.t9 source.t3 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
X23 source.t5 plus.t10 drain_left.t1 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X24 a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X25 source.t9 minus.t11 drain_right.t0 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.6
X26 a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X27 drain_left.t0 plus.t11 source.t7 a_n2018_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.6
R0 minus.n2 minus.t10 693.032
R1 minus.n14 minus.t11 693.032
R2 minus.n3 minus.t9 667.972
R3 minus.n4 minus.t7 667.972
R4 minus.n1 minus.t6 667.972
R5 minus.n8 minus.t2 667.972
R6 minus.n10 minus.t3 667.972
R7 minus.n15 minus.t5 667.972
R8 minus.n16 minus.t8 667.972
R9 minus.n13 minus.t0 667.972
R10 minus.n20 minus.t4 667.972
R11 minus.n22 minus.t1 667.972
R12 minus.n11 minus.n10 161.3
R13 minus.n9 minus.n0 161.3
R14 minus.n8 minus.n7 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n6 minus.n1 80.6037
R19 minus.n5 minus.n4 80.6037
R20 minus.n18 minus.n13 80.6037
R21 minus.n17 minus.n16 80.6037
R22 minus.n4 minus.n3 48.2005
R23 minus.n4 minus.n1 48.2005
R24 minus.n8 minus.n1 48.2005
R25 minus.n16 minus.n15 48.2005
R26 minus.n16 minus.n13 48.2005
R27 minus.n20 minus.n13 48.2005
R28 minus.n5 minus.n2 45.0744
R29 minus.n17 minus.n14 45.0744
R30 minus.n10 minus.n9 40.1672
R31 minus.n22 minus.n21 40.1672
R32 minus.n24 minus.n11 39.1255
R33 minus.n3 minus.n2 16.1124
R34 minus.n15 minus.n14 16.1124
R35 minus.n9 minus.n8 8.03383
R36 minus.n21 minus.n20 8.03383
R37 minus.n24 minus.n23 6.58762
R38 minus.n6 minus.n5 0.380177
R39 minus.n18 minus.n17 0.380177
R40 minus.n7 minus.n6 0.285035
R41 minus.n19 minus.n18 0.285035
R42 minus.n11 minus.n0 0.189894
R43 minus.n7 minus.n0 0.189894
R44 minus.n19 minus.n12 0.189894
R45 minus.n23 minus.n12 0.189894
R46 minus minus.n24 0.188
R47 source.n5 source.t5 45.521
R48 source.n6 source.t13 45.521
R49 source.n11 source.t16 45.521
R50 source.n23 source.t11 45.5208
R51 source.n18 source.t9 45.5208
R52 source.n17 source.t4 45.5208
R53 source.n12 source.t21 45.5208
R54 source.n0 source.t2 45.5208
R55 source.n2 source.n1 44.201
R56 source.n4 source.n3 44.201
R57 source.n8 source.n7 44.201
R58 source.n10 source.n9 44.201
R59 source.n22 source.n21 44.2008
R60 source.n20 source.n19 44.2008
R61 source.n16 source.n15 44.2008
R62 source.n14 source.n13 44.2008
R63 source.n12 source.n11 24.3622
R64 source.n24 source.n0 18.6984
R65 source.n24 source.n23 5.66429
R66 source.n21 source.t12 1.3205
R67 source.n21 source.t10 1.3205
R68 source.n19 source.t17 1.3205
R69 source.n19 source.t18 1.3205
R70 source.n15 source.t7 1.3205
R71 source.n15 source.t23 1.3205
R72 source.n13 source.t20 1.3205
R73 source.n13 source.t6 1.3205
R74 source.n1 source.t1 1.3205
R75 source.n1 source.t22 1.3205
R76 source.n3 source.t3 1.3205
R77 source.n3 source.t0 1.3205
R78 source.n7 source.t14 1.3205
R79 source.n7 source.t15 1.3205
R80 source.n9 source.t19 1.3205
R81 source.n9 source.t8 1.3205
R82 source.n11 source.n10 0.802224
R83 source.n10 source.n8 0.802224
R84 source.n8 source.n6 0.802224
R85 source.n5 source.n4 0.802224
R86 source.n4 source.n2 0.802224
R87 source.n2 source.n0 0.802224
R88 source.n14 source.n12 0.802224
R89 source.n16 source.n14 0.802224
R90 source.n17 source.n16 0.802224
R91 source.n20 source.n18 0.802224
R92 source.n22 source.n20 0.802224
R93 source.n23 source.n22 0.802224
R94 source.n6 source.n5 0.470328
R95 source.n18 source.n17 0.470328
R96 source source.n24 0.188
R97 drain_right.n6 drain_right.n4 61.6814
R98 drain_right.n3 drain_right.n2 61.6259
R99 drain_right.n3 drain_right.n0 61.6259
R100 drain_right.n6 drain_right.n5 60.8798
R101 drain_right.n8 drain_right.n7 60.8798
R102 drain_right.n3 drain_right.n1 60.8796
R103 drain_right drain_right.n3 33.0952
R104 drain_right drain_right.n8 6.45494
R105 drain_right.n1 drain_right.t3 1.3205
R106 drain_right.n1 drain_right.t11 1.3205
R107 drain_right.n2 drain_right.t7 1.3205
R108 drain_right.n2 drain_right.t10 1.3205
R109 drain_right.n0 drain_right.t0 1.3205
R110 drain_right.n0 drain_right.t6 1.3205
R111 drain_right.n4 drain_right.t2 1.3205
R112 drain_right.n4 drain_right.t1 1.3205
R113 drain_right.n5 drain_right.t5 1.3205
R114 drain_right.n5 drain_right.t4 1.3205
R115 drain_right.n7 drain_right.t8 1.3205
R116 drain_right.n7 drain_right.t9 1.3205
R117 drain_right.n8 drain_right.n6 0.802224
R118 plus.n4 plus.t10 693.032
R119 plus.n16 plus.t0 693.032
R120 plus.n10 plus.t2 667.972
R121 plus.n8 plus.t5 667.972
R122 plus.n7 plus.t7 667.972
R123 plus.n6 plus.t8 667.972
R124 plus.n5 plus.t9 667.972
R125 plus.n22 plus.t4 667.972
R126 plus.n20 plus.t3 667.972
R127 plus.n19 plus.t1 667.972
R128 plus.n18 plus.t11 667.972
R129 plus.n17 plus.t6 667.972
R130 plus.n8 plus.n1 161.3
R131 plus.n9 plus.n0 161.3
R132 plus.n11 plus.n10 161.3
R133 plus.n20 plus.n13 161.3
R134 plus.n21 plus.n12 161.3
R135 plus.n23 plus.n22 161.3
R136 plus.n6 plus.n3 80.6037
R137 plus.n7 plus.n2 80.6037
R138 plus.n18 plus.n15 80.6037
R139 plus.n19 plus.n14 80.6037
R140 plus.n8 plus.n7 48.2005
R141 plus.n7 plus.n6 48.2005
R142 plus.n6 plus.n5 48.2005
R143 plus.n20 plus.n19 48.2005
R144 plus.n19 plus.n18 48.2005
R145 plus.n18 plus.n17 48.2005
R146 plus.n4 plus.n3 45.0744
R147 plus.n16 plus.n15 45.0744
R148 plus.n10 plus.n9 40.1672
R149 plus.n22 plus.n21 40.1672
R150 plus plus.n23 31.8702
R151 plus.n5 plus.n4 16.1124
R152 plus.n17 plus.n16 16.1124
R153 plus plus.n11 13.3679
R154 plus.n9 plus.n8 8.03383
R155 plus.n21 plus.n20 8.03383
R156 plus.n3 plus.n2 0.380177
R157 plus.n15 plus.n14 0.380177
R158 plus.n2 plus.n1 0.285035
R159 plus.n14 plus.n13 0.285035
R160 plus.n1 plus.n0 0.189894
R161 plus.n11 plus.n0 0.189894
R162 plus.n23 plus.n12 0.189894
R163 plus.n13 plus.n12 0.189894
R164 drain_left.n6 drain_left.n4 61.6815
R165 drain_left.n3 drain_left.n2 61.6259
R166 drain_left.n3 drain_left.n0 61.6259
R167 drain_left.n6 drain_left.n5 60.8798
R168 drain_left.n8 drain_left.n7 60.8796
R169 drain_left.n3 drain_left.n1 60.8796
R170 drain_left drain_left.n3 33.6484
R171 drain_left drain_left.n8 6.45494
R172 drain_left.n1 drain_left.t10 1.3205
R173 drain_left.n1 drain_left.t0 1.3205
R174 drain_left.n2 drain_left.t5 1.3205
R175 drain_left.n2 drain_left.t11 1.3205
R176 drain_left.n0 drain_left.t7 1.3205
R177 drain_left.n0 drain_left.t8 1.3205
R178 drain_left.n7 drain_left.t6 1.3205
R179 drain_left.n7 drain_left.t9 1.3205
R180 drain_left.n5 drain_left.t3 1.3205
R181 drain_left.n5 drain_left.t4 1.3205
R182 drain_left.n4 drain_left.t1 1.3205
R183 drain_left.n4 drain_left.t2 1.3205
R184 drain_left.n8 drain_left.n6 0.802224
C0 drain_left drain_right 1.01253f
C1 source drain_right 20.223999f
C2 minus plus 6.21958f
C3 minus drain_left 0.17204f
C4 minus source 8.6368f
C5 plus drain_left 9.10987f
C6 source plus 8.65084f
C7 minus drain_right 8.9127f
C8 source drain_left 20.2225f
C9 plus drain_right 0.352374f
C10 drain_right a_n2018_n3888# 6.70528f
C11 drain_left a_n2018_n3888# 7.00048f
C12 source a_n2018_n3888# 10.688194f
C13 minus a_n2018_n3888# 8.13307f
C14 plus a_n2018_n3888# 10.06222f
C15 drain_left.t7 a_n2018_n3888# 0.332862f
C16 drain_left.t8 a_n2018_n3888# 0.332862f
C17 drain_left.n0 a_n2018_n3888# 3.01331f
C18 drain_left.t10 a_n2018_n3888# 0.332862f
C19 drain_left.t0 a_n2018_n3888# 0.332862f
C20 drain_left.n1 a_n2018_n3888# 3.00868f
C21 drain_left.t5 a_n2018_n3888# 0.332862f
C22 drain_left.t11 a_n2018_n3888# 0.332862f
C23 drain_left.n2 a_n2018_n3888# 3.01331f
C24 drain_left.n3 a_n2018_n3888# 2.70536f
C25 drain_left.t1 a_n2018_n3888# 0.332862f
C26 drain_left.t2 a_n2018_n3888# 0.332862f
C27 drain_left.n4 a_n2018_n3888# 3.0137f
C28 drain_left.t3 a_n2018_n3888# 0.332862f
C29 drain_left.t4 a_n2018_n3888# 0.332862f
C30 drain_left.n5 a_n2018_n3888# 3.00868f
C31 drain_left.n6 a_n2018_n3888# 0.756466f
C32 drain_left.t6 a_n2018_n3888# 0.332862f
C33 drain_left.t9 a_n2018_n3888# 0.332862f
C34 drain_left.n7 a_n2018_n3888# 3.00867f
C35 drain_left.n8 a_n2018_n3888# 0.619967f
C36 plus.n0 a_n2018_n3888# 0.044501f
C37 plus.t2 a_n2018_n3888# 1.13813f
C38 plus.t5 a_n2018_n3888# 1.13813f
C39 plus.n1 a_n2018_n3888# 0.059381f
C40 plus.t7 a_n2018_n3888# 1.13813f
C41 plus.n2 a_n2018_n3888# 0.074122f
C42 plus.t8 a_n2018_n3888# 1.13813f
C43 plus.n3 a_n2018_n3888# 0.228074f
C44 plus.t9 a_n2018_n3888# 1.13813f
C45 plus.t10 a_n2018_n3888# 1.15407f
C46 plus.n4 a_n2018_n3888# 0.428328f
C47 plus.n5 a_n2018_n3888# 0.449828f
C48 plus.n6 a_n2018_n3888# 0.451453f
C49 plus.n7 a_n2018_n3888# 0.451453f
C50 plus.n8 a_n2018_n3888# 0.442864f
C51 plus.n9 a_n2018_n3888# 0.010098f
C52 plus.n10 a_n2018_n3888# 0.439846f
C53 plus.n11 a_n2018_n3888# 0.57152f
C54 plus.n12 a_n2018_n3888# 0.044501f
C55 plus.t4 a_n2018_n3888# 1.13813f
C56 plus.n13 a_n2018_n3888# 0.059381f
C57 plus.t3 a_n2018_n3888# 1.13813f
C58 plus.n14 a_n2018_n3888# 0.074122f
C59 plus.t1 a_n2018_n3888# 1.13813f
C60 plus.n15 a_n2018_n3888# 0.228074f
C61 plus.t11 a_n2018_n3888# 1.13813f
C62 plus.t0 a_n2018_n3888# 1.15407f
C63 plus.n16 a_n2018_n3888# 0.428328f
C64 plus.t6 a_n2018_n3888# 1.13813f
C65 plus.n17 a_n2018_n3888# 0.449828f
C66 plus.n18 a_n2018_n3888# 0.451453f
C67 plus.n19 a_n2018_n3888# 0.451453f
C68 plus.n20 a_n2018_n3888# 0.442864f
C69 plus.n21 a_n2018_n3888# 0.010098f
C70 plus.n22 a_n2018_n3888# 0.439846f
C71 plus.n23 a_n2018_n3888# 1.46523f
C72 drain_right.t0 a_n2018_n3888# 0.331834f
C73 drain_right.t6 a_n2018_n3888# 0.331834f
C74 drain_right.n0 a_n2018_n3888# 3.004f
C75 drain_right.t3 a_n2018_n3888# 0.331834f
C76 drain_right.t11 a_n2018_n3888# 0.331834f
C77 drain_right.n1 a_n2018_n3888# 2.99939f
C78 drain_right.t7 a_n2018_n3888# 0.331834f
C79 drain_right.t10 a_n2018_n3888# 0.331834f
C80 drain_right.n2 a_n2018_n3888# 3.004f
C81 drain_right.n3 a_n2018_n3888# 2.6389f
C82 drain_right.t2 a_n2018_n3888# 0.331834f
C83 drain_right.t1 a_n2018_n3888# 0.331834f
C84 drain_right.n4 a_n2018_n3888# 3.00439f
C85 drain_right.t5 a_n2018_n3888# 0.331834f
C86 drain_right.t4 a_n2018_n3888# 0.331834f
C87 drain_right.n5 a_n2018_n3888# 2.99939f
C88 drain_right.n6 a_n2018_n3888# 0.75414f
C89 drain_right.t8 a_n2018_n3888# 0.331834f
C90 drain_right.t9 a_n2018_n3888# 0.331834f
C91 drain_right.n7 a_n2018_n3888# 2.99939f
C92 drain_right.n8 a_n2018_n3888# 0.618042f
C93 source.t2 a_n2018_n3888# 2.95093f
C94 source.n0 a_n2018_n3888# 1.39666f
C95 source.t1 a_n2018_n3888# 0.26332f
C96 source.t22 a_n2018_n3888# 0.26332f
C97 source.n1 a_n2018_n3888# 2.31305f
C98 source.n2 a_n2018_n3888# 0.333593f
C99 source.t3 a_n2018_n3888# 0.26332f
C100 source.t0 a_n2018_n3888# 0.26332f
C101 source.n3 a_n2018_n3888# 2.31305f
C102 source.n4 a_n2018_n3888# 0.333593f
C103 source.t5 a_n2018_n3888# 2.95093f
C104 source.n5 a_n2018_n3888# 0.390098f
C105 source.t13 a_n2018_n3888# 2.95093f
C106 source.n6 a_n2018_n3888# 0.390098f
C107 source.t14 a_n2018_n3888# 0.26332f
C108 source.t15 a_n2018_n3888# 0.26332f
C109 source.n7 a_n2018_n3888# 2.31305f
C110 source.n8 a_n2018_n3888# 0.333593f
C111 source.t19 a_n2018_n3888# 0.26332f
C112 source.t8 a_n2018_n3888# 0.26332f
C113 source.n9 a_n2018_n3888# 2.31305f
C114 source.n10 a_n2018_n3888# 0.333593f
C115 source.t16 a_n2018_n3888# 2.95093f
C116 source.n11 a_n2018_n3888# 1.77317f
C117 source.t21 a_n2018_n3888# 2.95093f
C118 source.n12 a_n2018_n3888# 1.77318f
C119 source.t20 a_n2018_n3888# 0.26332f
C120 source.t6 a_n2018_n3888# 0.26332f
C121 source.n13 a_n2018_n3888# 2.31305f
C122 source.n14 a_n2018_n3888# 0.333596f
C123 source.t7 a_n2018_n3888# 0.26332f
C124 source.t23 a_n2018_n3888# 0.26332f
C125 source.n15 a_n2018_n3888# 2.31305f
C126 source.n16 a_n2018_n3888# 0.333596f
C127 source.t4 a_n2018_n3888# 2.95093f
C128 source.n17 a_n2018_n3888# 0.390101f
C129 source.t9 a_n2018_n3888# 2.95093f
C130 source.n18 a_n2018_n3888# 0.390101f
C131 source.t17 a_n2018_n3888# 0.26332f
C132 source.t18 a_n2018_n3888# 0.26332f
C133 source.n19 a_n2018_n3888# 2.31305f
C134 source.n20 a_n2018_n3888# 0.333596f
C135 source.t12 a_n2018_n3888# 0.26332f
C136 source.t10 a_n2018_n3888# 0.26332f
C137 source.n21 a_n2018_n3888# 2.31305f
C138 source.n22 a_n2018_n3888# 0.333596f
C139 source.t11 a_n2018_n3888# 2.95093f
C140 source.n23 a_n2018_n3888# 0.530173f
C141 source.n24 a_n2018_n3888# 1.63532f
C142 minus.n0 a_n2018_n3888# 0.043781f
C143 minus.t6 a_n2018_n3888# 1.1197f
C144 minus.n1 a_n2018_n3888# 0.444145f
C145 minus.t2 a_n2018_n3888# 1.1197f
C146 minus.t10 a_n2018_n3888# 1.13539f
C147 minus.n2 a_n2018_n3888# 0.421394f
C148 minus.t9 a_n2018_n3888# 1.1197f
C149 minus.n3 a_n2018_n3888# 0.442546f
C150 minus.t7 a_n2018_n3888# 1.1197f
C151 minus.n4 a_n2018_n3888# 0.444145f
C152 minus.n5 a_n2018_n3888# 0.224382f
C153 minus.n6 a_n2018_n3888# 0.072922f
C154 minus.n7 a_n2018_n3888# 0.05842f
C155 minus.n8 a_n2018_n3888# 0.435694f
C156 minus.n9 a_n2018_n3888# 0.009935f
C157 minus.t3 a_n2018_n3888# 1.1197f
C158 minus.n10 a_n2018_n3888# 0.432725f
C159 minus.n11 a_n2018_n3888# 1.74692f
C160 minus.n12 a_n2018_n3888# 0.043781f
C161 minus.t0 a_n2018_n3888# 1.1197f
C162 minus.n13 a_n2018_n3888# 0.444145f
C163 minus.t11 a_n2018_n3888# 1.13539f
C164 minus.n14 a_n2018_n3888# 0.421394f
C165 minus.t5 a_n2018_n3888# 1.1197f
C166 minus.n15 a_n2018_n3888# 0.442546f
C167 minus.t8 a_n2018_n3888# 1.1197f
C168 minus.n16 a_n2018_n3888# 0.444145f
C169 minus.n17 a_n2018_n3888# 0.224382f
C170 minus.n18 a_n2018_n3888# 0.072922f
C171 minus.n19 a_n2018_n3888# 0.05842f
C172 minus.t4 a_n2018_n3888# 1.1197f
C173 minus.n20 a_n2018_n3888# 0.435694f
C174 minus.n21 a_n2018_n3888# 0.009935f
C175 minus.t1 a_n2018_n3888# 1.1197f
C176 minus.n22 a_n2018_n3888# 0.432725f
C177 minus.n23 a_n2018_n3888# 0.295227f
C178 minus.n24 a_n2018_n3888# 2.10113f
.ends

