* NGSPICE file created from diffpair708.ext - technology: sky130A

.subckt diffpair708 minus drain_right drain_left source plus
X0 source.t38 minus.t0 drain_right.t10 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X1 source.t9 plus.t0 drain_left.t19 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X2 drain_right.t9 minus.t1 source.t37 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X3 source.t17 plus.t1 drain_left.t18 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X4 source.t0 plus.t2 drain_left.t17 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X5 source.t36 minus.t2 drain_right.t8 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X6 source.t35 minus.t3 drain_right.t13 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X7 a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.7
X8 drain_left.t16 plus.t3 source.t16 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X9 source.t3 plus.t4 drain_left.t15 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X10 source.t18 plus.t5 drain_left.t14 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X11 source.t5 plus.t6 drain_left.t13 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X12 drain_left.t12 plus.t7 source.t10 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X13 drain_right.t12 minus.t4 source.t34 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X14 source.t33 minus.t5 drain_right.t11 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X15 drain_right.t5 minus.t6 source.t32 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X16 a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X17 drain_right.t4 minus.t7 source.t31 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X18 drain_right.t3 minus.t8 source.t30 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X19 drain_right.t2 minus.t9 source.t29 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X20 drain_left.t11 plus.t8 source.t4 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X21 drain_right.t1 minus.t10 source.t28 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X22 source.t39 plus.t9 drain_left.t10 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X23 drain_left.t9 plus.t10 source.t12 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X24 drain_left.t8 plus.t11 source.t15 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X25 drain_left.t7 plus.t12 source.t6 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X26 drain_right.t0 minus.t11 source.t27 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
X27 drain_left.t6 plus.t13 source.t13 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X28 a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X29 source.t26 minus.t12 drain_right.t19 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X30 drain_right.t18 minus.t13 source.t25 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X31 a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.7
X32 drain_left.t5 plus.t14 source.t14 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X33 source.t24 minus.t14 drain_right.t17 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X34 source.t2 plus.t15 drain_left.t4 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.7
X35 drain_left.t3 plus.t16 source.t7 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X36 source.t23 minus.t15 drain_right.t16 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X37 drain_right.t15 minus.t16 source.t22 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X38 source.t21 minus.t17 drain_right.t14 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X39 source.t20 minus.t18 drain_right.t7 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X40 source.t19 minus.t19 drain_right.t6 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X41 source.t1 plus.t17 drain_left.t2 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X42 source.t11 plus.t18 drain_left.t1 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.7
X43 drain_left.t0 plus.t19 source.t8 a_n2982_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.7
R0 minus.n9 minus.t11 942.226
R1 minus.n43 minus.t5 942.226
R2 minus.n8 minus.t2 916.833
R3 minus.n12 minus.t10 916.833
R4 minus.n14 minus.t18 916.833
R5 minus.n18 minus.t9 916.833
R6 minus.n20 minus.t19 916.833
R7 minus.n24 minus.t8 916.833
R8 minus.n26 minus.t15 916.833
R9 minus.n30 minus.t6 916.833
R10 minus.n32 minus.t14 916.833
R11 minus.n42 minus.t4 916.833
R12 minus.n46 minus.t0 916.833
R13 minus.n48 minus.t1 916.833
R14 minus.n52 minus.t3 916.833
R15 minus.n54 minus.t16 916.833
R16 minus.n58 minus.t17 916.833
R17 minus.n60 minus.t13 916.833
R18 minus.n64 minus.t12 916.833
R19 minus.n66 minus.t7 916.833
R20 minus.n33 minus.n32 161.3
R21 minus.n31 minus.n0 161.3
R22 minus.n30 minus.n29 161.3
R23 minus.n28 minus.n1 161.3
R24 minus.n27 minus.n26 161.3
R25 minus.n25 minus.n2 161.3
R26 minus.n24 minus.n23 161.3
R27 minus.n22 minus.n3 161.3
R28 minus.n21 minus.n20 161.3
R29 minus.n19 minus.n4 161.3
R30 minus.n18 minus.n17 161.3
R31 minus.n16 minus.n5 161.3
R32 minus.n15 minus.n14 161.3
R33 minus.n13 minus.n6 161.3
R34 minus.n12 minus.n11 161.3
R35 minus.n10 minus.n7 161.3
R36 minus.n67 minus.n66 161.3
R37 minus.n65 minus.n34 161.3
R38 minus.n64 minus.n63 161.3
R39 minus.n62 minus.n35 161.3
R40 minus.n61 minus.n60 161.3
R41 minus.n59 minus.n36 161.3
R42 minus.n58 minus.n57 161.3
R43 minus.n56 minus.n37 161.3
R44 minus.n55 minus.n54 161.3
R45 minus.n53 minus.n38 161.3
R46 minus.n52 minus.n51 161.3
R47 minus.n50 minus.n39 161.3
R48 minus.n49 minus.n48 161.3
R49 minus.n47 minus.n40 161.3
R50 minus.n46 minus.n45 161.3
R51 minus.n44 minus.n41 161.3
R52 minus.n68 minus.n33 50.4323
R53 minus.n10 minus.n9 45.0031
R54 minus.n44 minus.n43 45.0031
R55 minus.n32 minus.n31 41.6278
R56 minus.n66 minus.n65 41.6278
R57 minus.n8 minus.n7 37.246
R58 minus.n30 minus.n1 37.246
R59 minus.n42 minus.n41 37.246
R60 minus.n64 minus.n35 37.246
R61 minus.n13 minus.n12 32.8641
R62 minus.n26 minus.n25 32.8641
R63 minus.n47 minus.n46 32.8641
R64 minus.n60 minus.n59 32.8641
R65 minus.n14 minus.n5 28.4823
R66 minus.n24 minus.n3 28.4823
R67 minus.n48 minus.n39 28.4823
R68 minus.n58 minus.n37 28.4823
R69 minus.n20 minus.n19 24.1005
R70 minus.n19 minus.n18 24.1005
R71 minus.n53 minus.n52 24.1005
R72 minus.n54 minus.n53 24.1005
R73 minus.n18 minus.n5 19.7187
R74 minus.n20 minus.n3 19.7187
R75 minus.n52 minus.n39 19.7187
R76 minus.n54 minus.n37 19.7187
R77 minus.n9 minus.n8 15.6319
R78 minus.n43 minus.n42 15.6319
R79 minus.n14 minus.n13 15.3369
R80 minus.n25 minus.n24 15.3369
R81 minus.n48 minus.n47 15.3369
R82 minus.n59 minus.n58 15.3369
R83 minus.n12 minus.n7 10.955
R84 minus.n26 minus.n1 10.955
R85 minus.n46 minus.n41 10.955
R86 minus.n60 minus.n35 10.955
R87 minus.n68 minus.n67 6.66717
R88 minus.n31 minus.n30 6.57323
R89 minus.n65 minus.n64 6.57323
R90 minus.n33 minus.n0 0.189894
R91 minus.n29 minus.n0 0.189894
R92 minus.n29 minus.n28 0.189894
R93 minus.n28 minus.n27 0.189894
R94 minus.n27 minus.n2 0.189894
R95 minus.n23 minus.n2 0.189894
R96 minus.n23 minus.n22 0.189894
R97 minus.n22 minus.n21 0.189894
R98 minus.n21 minus.n4 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n17 minus.n16 0.189894
R101 minus.n16 minus.n15 0.189894
R102 minus.n15 minus.n6 0.189894
R103 minus.n11 minus.n6 0.189894
R104 minus.n11 minus.n10 0.189894
R105 minus.n45 minus.n44 0.189894
R106 minus.n45 minus.n40 0.189894
R107 minus.n49 minus.n40 0.189894
R108 minus.n50 minus.n49 0.189894
R109 minus.n51 minus.n50 0.189894
R110 minus.n51 minus.n38 0.189894
R111 minus.n55 minus.n38 0.189894
R112 minus.n56 minus.n55 0.189894
R113 minus.n57 minus.n56 0.189894
R114 minus.n57 minus.n36 0.189894
R115 minus.n61 minus.n36 0.189894
R116 minus.n62 minus.n61 0.189894
R117 minus.n63 minus.n62 0.189894
R118 minus.n63 minus.n34 0.189894
R119 minus.n67 minus.n34 0.189894
R120 minus minus.n68 0.188
R121 drain_right.n6 drain_right.n4 59.6034
R122 drain_right.n2 drain_right.n0 59.6034
R123 drain_right.n10 drain_right.n8 59.6032
R124 drain_right.n7 drain_right.n3 58.7154
R125 drain_right.n6 drain_right.n5 58.7154
R126 drain_right.n2 drain_right.n1 58.7154
R127 drain_right.n10 drain_right.n9 58.7154
R128 drain_right.n12 drain_right.n11 58.7154
R129 drain_right.n14 drain_right.n13 58.7154
R130 drain_right.n16 drain_right.n15 58.7154
R131 drain_right drain_right.n7 43.7658
R132 drain_right drain_right.n16 6.54115
R133 drain_right.n16 drain_right.n14 0.888431
R134 drain_right.n14 drain_right.n12 0.888431
R135 drain_right.n12 drain_right.n10 0.888431
R136 drain_right.n7 drain_right.n6 0.833085
R137 drain_right.n7 drain_right.n2 0.833085
R138 drain_right.n3 drain_right.t13 0.7925
R139 drain_right.n3 drain_right.t15 0.7925
R140 drain_right.n4 drain_right.t19 0.7925
R141 drain_right.n4 drain_right.t4 0.7925
R142 drain_right.n5 drain_right.t14 0.7925
R143 drain_right.n5 drain_right.t18 0.7925
R144 drain_right.n1 drain_right.t10 0.7925
R145 drain_right.n1 drain_right.t9 0.7925
R146 drain_right.n0 drain_right.t11 0.7925
R147 drain_right.n0 drain_right.t12 0.7925
R148 drain_right.n8 drain_right.t8 0.7925
R149 drain_right.n8 drain_right.t0 0.7925
R150 drain_right.n9 drain_right.t7 0.7925
R151 drain_right.n9 drain_right.t1 0.7925
R152 drain_right.n11 drain_right.t6 0.7925
R153 drain_right.n11 drain_right.t2 0.7925
R154 drain_right.n13 drain_right.t16 0.7925
R155 drain_right.n13 drain_right.t3 0.7925
R156 drain_right.n15 drain_right.t17 0.7925
R157 drain_right.n15 drain_right.t5 0.7925
R158 source.n1146 source.n1012 289.615
R159 source.n998 source.n864 289.615
R160 source.n858 source.n724 289.615
R161 source.n710 source.n576 289.615
R162 source.n134 source.n0 289.615
R163 source.n282 source.n148 289.615
R164 source.n422 source.n288 289.615
R165 source.n570 source.n436 289.615
R166 source.n1056 source.n1055 185
R167 source.n1061 source.n1060 185
R168 source.n1063 source.n1062 185
R169 source.n1052 source.n1051 185
R170 source.n1069 source.n1068 185
R171 source.n1071 source.n1070 185
R172 source.n1048 source.n1047 185
R173 source.n1078 source.n1077 185
R174 source.n1079 source.n1046 185
R175 source.n1081 source.n1080 185
R176 source.n1044 source.n1043 185
R177 source.n1087 source.n1086 185
R178 source.n1089 source.n1088 185
R179 source.n1040 source.n1039 185
R180 source.n1095 source.n1094 185
R181 source.n1097 source.n1096 185
R182 source.n1036 source.n1035 185
R183 source.n1103 source.n1102 185
R184 source.n1105 source.n1104 185
R185 source.n1032 source.n1031 185
R186 source.n1111 source.n1110 185
R187 source.n1113 source.n1112 185
R188 source.n1028 source.n1027 185
R189 source.n1119 source.n1118 185
R190 source.n1122 source.n1121 185
R191 source.n1120 source.n1024 185
R192 source.n1127 source.n1023 185
R193 source.n1129 source.n1128 185
R194 source.n1131 source.n1130 185
R195 source.n1020 source.n1019 185
R196 source.n1137 source.n1136 185
R197 source.n1139 source.n1138 185
R198 source.n1016 source.n1015 185
R199 source.n1145 source.n1144 185
R200 source.n1147 source.n1146 185
R201 source.n908 source.n907 185
R202 source.n913 source.n912 185
R203 source.n915 source.n914 185
R204 source.n904 source.n903 185
R205 source.n921 source.n920 185
R206 source.n923 source.n922 185
R207 source.n900 source.n899 185
R208 source.n930 source.n929 185
R209 source.n931 source.n898 185
R210 source.n933 source.n932 185
R211 source.n896 source.n895 185
R212 source.n939 source.n938 185
R213 source.n941 source.n940 185
R214 source.n892 source.n891 185
R215 source.n947 source.n946 185
R216 source.n949 source.n948 185
R217 source.n888 source.n887 185
R218 source.n955 source.n954 185
R219 source.n957 source.n956 185
R220 source.n884 source.n883 185
R221 source.n963 source.n962 185
R222 source.n965 source.n964 185
R223 source.n880 source.n879 185
R224 source.n971 source.n970 185
R225 source.n974 source.n973 185
R226 source.n972 source.n876 185
R227 source.n979 source.n875 185
R228 source.n981 source.n980 185
R229 source.n983 source.n982 185
R230 source.n872 source.n871 185
R231 source.n989 source.n988 185
R232 source.n991 source.n990 185
R233 source.n868 source.n867 185
R234 source.n997 source.n996 185
R235 source.n999 source.n998 185
R236 source.n768 source.n767 185
R237 source.n773 source.n772 185
R238 source.n775 source.n774 185
R239 source.n764 source.n763 185
R240 source.n781 source.n780 185
R241 source.n783 source.n782 185
R242 source.n760 source.n759 185
R243 source.n790 source.n789 185
R244 source.n791 source.n758 185
R245 source.n793 source.n792 185
R246 source.n756 source.n755 185
R247 source.n799 source.n798 185
R248 source.n801 source.n800 185
R249 source.n752 source.n751 185
R250 source.n807 source.n806 185
R251 source.n809 source.n808 185
R252 source.n748 source.n747 185
R253 source.n815 source.n814 185
R254 source.n817 source.n816 185
R255 source.n744 source.n743 185
R256 source.n823 source.n822 185
R257 source.n825 source.n824 185
R258 source.n740 source.n739 185
R259 source.n831 source.n830 185
R260 source.n834 source.n833 185
R261 source.n832 source.n736 185
R262 source.n839 source.n735 185
R263 source.n841 source.n840 185
R264 source.n843 source.n842 185
R265 source.n732 source.n731 185
R266 source.n849 source.n848 185
R267 source.n851 source.n850 185
R268 source.n728 source.n727 185
R269 source.n857 source.n856 185
R270 source.n859 source.n858 185
R271 source.n620 source.n619 185
R272 source.n625 source.n624 185
R273 source.n627 source.n626 185
R274 source.n616 source.n615 185
R275 source.n633 source.n632 185
R276 source.n635 source.n634 185
R277 source.n612 source.n611 185
R278 source.n642 source.n641 185
R279 source.n643 source.n610 185
R280 source.n645 source.n644 185
R281 source.n608 source.n607 185
R282 source.n651 source.n650 185
R283 source.n653 source.n652 185
R284 source.n604 source.n603 185
R285 source.n659 source.n658 185
R286 source.n661 source.n660 185
R287 source.n600 source.n599 185
R288 source.n667 source.n666 185
R289 source.n669 source.n668 185
R290 source.n596 source.n595 185
R291 source.n675 source.n674 185
R292 source.n677 source.n676 185
R293 source.n592 source.n591 185
R294 source.n683 source.n682 185
R295 source.n686 source.n685 185
R296 source.n684 source.n588 185
R297 source.n691 source.n587 185
R298 source.n693 source.n692 185
R299 source.n695 source.n694 185
R300 source.n584 source.n583 185
R301 source.n701 source.n700 185
R302 source.n703 source.n702 185
R303 source.n580 source.n579 185
R304 source.n709 source.n708 185
R305 source.n711 source.n710 185
R306 source.n135 source.n134 185
R307 source.n133 source.n132 185
R308 source.n4 source.n3 185
R309 source.n127 source.n126 185
R310 source.n125 source.n124 185
R311 source.n8 source.n7 185
R312 source.n119 source.n118 185
R313 source.n117 source.n116 185
R314 source.n115 source.n11 185
R315 source.n15 source.n12 185
R316 source.n110 source.n109 185
R317 source.n108 source.n107 185
R318 source.n17 source.n16 185
R319 source.n102 source.n101 185
R320 source.n100 source.n99 185
R321 source.n21 source.n20 185
R322 source.n94 source.n93 185
R323 source.n92 source.n91 185
R324 source.n25 source.n24 185
R325 source.n86 source.n85 185
R326 source.n84 source.n83 185
R327 source.n29 source.n28 185
R328 source.n78 source.n77 185
R329 source.n76 source.n75 185
R330 source.n33 source.n32 185
R331 source.n70 source.n69 185
R332 source.n68 source.n35 185
R333 source.n67 source.n66 185
R334 source.n38 source.n36 185
R335 source.n61 source.n60 185
R336 source.n59 source.n58 185
R337 source.n42 source.n41 185
R338 source.n53 source.n52 185
R339 source.n51 source.n50 185
R340 source.n46 source.n45 185
R341 source.n283 source.n282 185
R342 source.n281 source.n280 185
R343 source.n152 source.n151 185
R344 source.n275 source.n274 185
R345 source.n273 source.n272 185
R346 source.n156 source.n155 185
R347 source.n267 source.n266 185
R348 source.n265 source.n264 185
R349 source.n263 source.n159 185
R350 source.n163 source.n160 185
R351 source.n258 source.n257 185
R352 source.n256 source.n255 185
R353 source.n165 source.n164 185
R354 source.n250 source.n249 185
R355 source.n248 source.n247 185
R356 source.n169 source.n168 185
R357 source.n242 source.n241 185
R358 source.n240 source.n239 185
R359 source.n173 source.n172 185
R360 source.n234 source.n233 185
R361 source.n232 source.n231 185
R362 source.n177 source.n176 185
R363 source.n226 source.n225 185
R364 source.n224 source.n223 185
R365 source.n181 source.n180 185
R366 source.n218 source.n217 185
R367 source.n216 source.n183 185
R368 source.n215 source.n214 185
R369 source.n186 source.n184 185
R370 source.n209 source.n208 185
R371 source.n207 source.n206 185
R372 source.n190 source.n189 185
R373 source.n201 source.n200 185
R374 source.n199 source.n198 185
R375 source.n194 source.n193 185
R376 source.n423 source.n422 185
R377 source.n421 source.n420 185
R378 source.n292 source.n291 185
R379 source.n415 source.n414 185
R380 source.n413 source.n412 185
R381 source.n296 source.n295 185
R382 source.n407 source.n406 185
R383 source.n405 source.n404 185
R384 source.n403 source.n299 185
R385 source.n303 source.n300 185
R386 source.n398 source.n397 185
R387 source.n396 source.n395 185
R388 source.n305 source.n304 185
R389 source.n390 source.n389 185
R390 source.n388 source.n387 185
R391 source.n309 source.n308 185
R392 source.n382 source.n381 185
R393 source.n380 source.n379 185
R394 source.n313 source.n312 185
R395 source.n374 source.n373 185
R396 source.n372 source.n371 185
R397 source.n317 source.n316 185
R398 source.n366 source.n365 185
R399 source.n364 source.n363 185
R400 source.n321 source.n320 185
R401 source.n358 source.n357 185
R402 source.n356 source.n323 185
R403 source.n355 source.n354 185
R404 source.n326 source.n324 185
R405 source.n349 source.n348 185
R406 source.n347 source.n346 185
R407 source.n330 source.n329 185
R408 source.n341 source.n340 185
R409 source.n339 source.n338 185
R410 source.n334 source.n333 185
R411 source.n571 source.n570 185
R412 source.n569 source.n568 185
R413 source.n440 source.n439 185
R414 source.n563 source.n562 185
R415 source.n561 source.n560 185
R416 source.n444 source.n443 185
R417 source.n555 source.n554 185
R418 source.n553 source.n552 185
R419 source.n551 source.n447 185
R420 source.n451 source.n448 185
R421 source.n546 source.n545 185
R422 source.n544 source.n543 185
R423 source.n453 source.n452 185
R424 source.n538 source.n537 185
R425 source.n536 source.n535 185
R426 source.n457 source.n456 185
R427 source.n530 source.n529 185
R428 source.n528 source.n527 185
R429 source.n461 source.n460 185
R430 source.n522 source.n521 185
R431 source.n520 source.n519 185
R432 source.n465 source.n464 185
R433 source.n514 source.n513 185
R434 source.n512 source.n511 185
R435 source.n469 source.n468 185
R436 source.n506 source.n505 185
R437 source.n504 source.n471 185
R438 source.n503 source.n502 185
R439 source.n474 source.n472 185
R440 source.n497 source.n496 185
R441 source.n495 source.n494 185
R442 source.n478 source.n477 185
R443 source.n489 source.n488 185
R444 source.n487 source.n486 185
R445 source.n482 source.n481 185
R446 source.n1057 source.t31 149.524
R447 source.n909 source.t33 149.524
R448 source.n769 source.t8 149.524
R449 source.n621 source.t2 149.524
R450 source.n47 source.t16 149.524
R451 source.n195 source.t5 149.524
R452 source.n335 source.t27 149.524
R453 source.n483 source.t24 149.524
R454 source.n1061 source.n1055 104.615
R455 source.n1062 source.n1061 104.615
R456 source.n1062 source.n1051 104.615
R457 source.n1069 source.n1051 104.615
R458 source.n1070 source.n1069 104.615
R459 source.n1070 source.n1047 104.615
R460 source.n1078 source.n1047 104.615
R461 source.n1079 source.n1078 104.615
R462 source.n1080 source.n1079 104.615
R463 source.n1080 source.n1043 104.615
R464 source.n1087 source.n1043 104.615
R465 source.n1088 source.n1087 104.615
R466 source.n1088 source.n1039 104.615
R467 source.n1095 source.n1039 104.615
R468 source.n1096 source.n1095 104.615
R469 source.n1096 source.n1035 104.615
R470 source.n1103 source.n1035 104.615
R471 source.n1104 source.n1103 104.615
R472 source.n1104 source.n1031 104.615
R473 source.n1111 source.n1031 104.615
R474 source.n1112 source.n1111 104.615
R475 source.n1112 source.n1027 104.615
R476 source.n1119 source.n1027 104.615
R477 source.n1121 source.n1119 104.615
R478 source.n1121 source.n1120 104.615
R479 source.n1120 source.n1023 104.615
R480 source.n1129 source.n1023 104.615
R481 source.n1130 source.n1129 104.615
R482 source.n1130 source.n1019 104.615
R483 source.n1137 source.n1019 104.615
R484 source.n1138 source.n1137 104.615
R485 source.n1138 source.n1015 104.615
R486 source.n1145 source.n1015 104.615
R487 source.n1146 source.n1145 104.615
R488 source.n913 source.n907 104.615
R489 source.n914 source.n913 104.615
R490 source.n914 source.n903 104.615
R491 source.n921 source.n903 104.615
R492 source.n922 source.n921 104.615
R493 source.n922 source.n899 104.615
R494 source.n930 source.n899 104.615
R495 source.n931 source.n930 104.615
R496 source.n932 source.n931 104.615
R497 source.n932 source.n895 104.615
R498 source.n939 source.n895 104.615
R499 source.n940 source.n939 104.615
R500 source.n940 source.n891 104.615
R501 source.n947 source.n891 104.615
R502 source.n948 source.n947 104.615
R503 source.n948 source.n887 104.615
R504 source.n955 source.n887 104.615
R505 source.n956 source.n955 104.615
R506 source.n956 source.n883 104.615
R507 source.n963 source.n883 104.615
R508 source.n964 source.n963 104.615
R509 source.n964 source.n879 104.615
R510 source.n971 source.n879 104.615
R511 source.n973 source.n971 104.615
R512 source.n973 source.n972 104.615
R513 source.n972 source.n875 104.615
R514 source.n981 source.n875 104.615
R515 source.n982 source.n981 104.615
R516 source.n982 source.n871 104.615
R517 source.n989 source.n871 104.615
R518 source.n990 source.n989 104.615
R519 source.n990 source.n867 104.615
R520 source.n997 source.n867 104.615
R521 source.n998 source.n997 104.615
R522 source.n773 source.n767 104.615
R523 source.n774 source.n773 104.615
R524 source.n774 source.n763 104.615
R525 source.n781 source.n763 104.615
R526 source.n782 source.n781 104.615
R527 source.n782 source.n759 104.615
R528 source.n790 source.n759 104.615
R529 source.n791 source.n790 104.615
R530 source.n792 source.n791 104.615
R531 source.n792 source.n755 104.615
R532 source.n799 source.n755 104.615
R533 source.n800 source.n799 104.615
R534 source.n800 source.n751 104.615
R535 source.n807 source.n751 104.615
R536 source.n808 source.n807 104.615
R537 source.n808 source.n747 104.615
R538 source.n815 source.n747 104.615
R539 source.n816 source.n815 104.615
R540 source.n816 source.n743 104.615
R541 source.n823 source.n743 104.615
R542 source.n824 source.n823 104.615
R543 source.n824 source.n739 104.615
R544 source.n831 source.n739 104.615
R545 source.n833 source.n831 104.615
R546 source.n833 source.n832 104.615
R547 source.n832 source.n735 104.615
R548 source.n841 source.n735 104.615
R549 source.n842 source.n841 104.615
R550 source.n842 source.n731 104.615
R551 source.n849 source.n731 104.615
R552 source.n850 source.n849 104.615
R553 source.n850 source.n727 104.615
R554 source.n857 source.n727 104.615
R555 source.n858 source.n857 104.615
R556 source.n625 source.n619 104.615
R557 source.n626 source.n625 104.615
R558 source.n626 source.n615 104.615
R559 source.n633 source.n615 104.615
R560 source.n634 source.n633 104.615
R561 source.n634 source.n611 104.615
R562 source.n642 source.n611 104.615
R563 source.n643 source.n642 104.615
R564 source.n644 source.n643 104.615
R565 source.n644 source.n607 104.615
R566 source.n651 source.n607 104.615
R567 source.n652 source.n651 104.615
R568 source.n652 source.n603 104.615
R569 source.n659 source.n603 104.615
R570 source.n660 source.n659 104.615
R571 source.n660 source.n599 104.615
R572 source.n667 source.n599 104.615
R573 source.n668 source.n667 104.615
R574 source.n668 source.n595 104.615
R575 source.n675 source.n595 104.615
R576 source.n676 source.n675 104.615
R577 source.n676 source.n591 104.615
R578 source.n683 source.n591 104.615
R579 source.n685 source.n683 104.615
R580 source.n685 source.n684 104.615
R581 source.n684 source.n587 104.615
R582 source.n693 source.n587 104.615
R583 source.n694 source.n693 104.615
R584 source.n694 source.n583 104.615
R585 source.n701 source.n583 104.615
R586 source.n702 source.n701 104.615
R587 source.n702 source.n579 104.615
R588 source.n709 source.n579 104.615
R589 source.n710 source.n709 104.615
R590 source.n134 source.n133 104.615
R591 source.n133 source.n3 104.615
R592 source.n126 source.n3 104.615
R593 source.n126 source.n125 104.615
R594 source.n125 source.n7 104.615
R595 source.n118 source.n7 104.615
R596 source.n118 source.n117 104.615
R597 source.n117 source.n11 104.615
R598 source.n15 source.n11 104.615
R599 source.n109 source.n15 104.615
R600 source.n109 source.n108 104.615
R601 source.n108 source.n16 104.615
R602 source.n101 source.n16 104.615
R603 source.n101 source.n100 104.615
R604 source.n100 source.n20 104.615
R605 source.n93 source.n20 104.615
R606 source.n93 source.n92 104.615
R607 source.n92 source.n24 104.615
R608 source.n85 source.n24 104.615
R609 source.n85 source.n84 104.615
R610 source.n84 source.n28 104.615
R611 source.n77 source.n28 104.615
R612 source.n77 source.n76 104.615
R613 source.n76 source.n32 104.615
R614 source.n69 source.n32 104.615
R615 source.n69 source.n68 104.615
R616 source.n68 source.n67 104.615
R617 source.n67 source.n36 104.615
R618 source.n60 source.n36 104.615
R619 source.n60 source.n59 104.615
R620 source.n59 source.n41 104.615
R621 source.n52 source.n41 104.615
R622 source.n52 source.n51 104.615
R623 source.n51 source.n45 104.615
R624 source.n282 source.n281 104.615
R625 source.n281 source.n151 104.615
R626 source.n274 source.n151 104.615
R627 source.n274 source.n273 104.615
R628 source.n273 source.n155 104.615
R629 source.n266 source.n155 104.615
R630 source.n266 source.n265 104.615
R631 source.n265 source.n159 104.615
R632 source.n163 source.n159 104.615
R633 source.n257 source.n163 104.615
R634 source.n257 source.n256 104.615
R635 source.n256 source.n164 104.615
R636 source.n249 source.n164 104.615
R637 source.n249 source.n248 104.615
R638 source.n248 source.n168 104.615
R639 source.n241 source.n168 104.615
R640 source.n241 source.n240 104.615
R641 source.n240 source.n172 104.615
R642 source.n233 source.n172 104.615
R643 source.n233 source.n232 104.615
R644 source.n232 source.n176 104.615
R645 source.n225 source.n176 104.615
R646 source.n225 source.n224 104.615
R647 source.n224 source.n180 104.615
R648 source.n217 source.n180 104.615
R649 source.n217 source.n216 104.615
R650 source.n216 source.n215 104.615
R651 source.n215 source.n184 104.615
R652 source.n208 source.n184 104.615
R653 source.n208 source.n207 104.615
R654 source.n207 source.n189 104.615
R655 source.n200 source.n189 104.615
R656 source.n200 source.n199 104.615
R657 source.n199 source.n193 104.615
R658 source.n422 source.n421 104.615
R659 source.n421 source.n291 104.615
R660 source.n414 source.n291 104.615
R661 source.n414 source.n413 104.615
R662 source.n413 source.n295 104.615
R663 source.n406 source.n295 104.615
R664 source.n406 source.n405 104.615
R665 source.n405 source.n299 104.615
R666 source.n303 source.n299 104.615
R667 source.n397 source.n303 104.615
R668 source.n397 source.n396 104.615
R669 source.n396 source.n304 104.615
R670 source.n389 source.n304 104.615
R671 source.n389 source.n388 104.615
R672 source.n388 source.n308 104.615
R673 source.n381 source.n308 104.615
R674 source.n381 source.n380 104.615
R675 source.n380 source.n312 104.615
R676 source.n373 source.n312 104.615
R677 source.n373 source.n372 104.615
R678 source.n372 source.n316 104.615
R679 source.n365 source.n316 104.615
R680 source.n365 source.n364 104.615
R681 source.n364 source.n320 104.615
R682 source.n357 source.n320 104.615
R683 source.n357 source.n356 104.615
R684 source.n356 source.n355 104.615
R685 source.n355 source.n324 104.615
R686 source.n348 source.n324 104.615
R687 source.n348 source.n347 104.615
R688 source.n347 source.n329 104.615
R689 source.n340 source.n329 104.615
R690 source.n340 source.n339 104.615
R691 source.n339 source.n333 104.615
R692 source.n570 source.n569 104.615
R693 source.n569 source.n439 104.615
R694 source.n562 source.n439 104.615
R695 source.n562 source.n561 104.615
R696 source.n561 source.n443 104.615
R697 source.n554 source.n443 104.615
R698 source.n554 source.n553 104.615
R699 source.n553 source.n447 104.615
R700 source.n451 source.n447 104.615
R701 source.n545 source.n451 104.615
R702 source.n545 source.n544 104.615
R703 source.n544 source.n452 104.615
R704 source.n537 source.n452 104.615
R705 source.n537 source.n536 104.615
R706 source.n536 source.n456 104.615
R707 source.n529 source.n456 104.615
R708 source.n529 source.n528 104.615
R709 source.n528 source.n460 104.615
R710 source.n521 source.n460 104.615
R711 source.n521 source.n520 104.615
R712 source.n520 source.n464 104.615
R713 source.n513 source.n464 104.615
R714 source.n513 source.n512 104.615
R715 source.n512 source.n468 104.615
R716 source.n505 source.n468 104.615
R717 source.n505 source.n504 104.615
R718 source.n504 source.n503 104.615
R719 source.n503 source.n472 104.615
R720 source.n496 source.n472 104.615
R721 source.n496 source.n495 104.615
R722 source.n495 source.n477 104.615
R723 source.n488 source.n477 104.615
R724 source.n488 source.n487 104.615
R725 source.n487 source.n481 104.615
R726 source.t31 source.n1055 52.3082
R727 source.t33 source.n907 52.3082
R728 source.t8 source.n767 52.3082
R729 source.t2 source.n619 52.3082
R730 source.t16 source.n45 52.3082
R731 source.t5 source.n193 52.3082
R732 source.t27 source.n333 52.3082
R733 source.t24 source.n481 52.3082
R734 source.n1011 source.n1010 42.0366
R735 source.n1009 source.n1008 42.0366
R736 source.n1007 source.n1006 42.0366
R737 source.n1005 source.n1004 42.0366
R738 source.n723 source.n722 42.0366
R739 source.n721 source.n720 42.0366
R740 source.n719 source.n718 42.0366
R741 source.n717 source.n716 42.0366
R742 source.n141 source.n140 42.0366
R743 source.n143 source.n142 42.0366
R744 source.n145 source.n144 42.0366
R745 source.n147 source.n146 42.0366
R746 source.n429 source.n428 42.0366
R747 source.n431 source.n430 42.0366
R748 source.n433 source.n432 42.0366
R749 source.n435 source.n434 42.0366
R750 source.n715 source.n575 32.0241
R751 source.n1151 source.n1150 30.6338
R752 source.n1003 source.n1002 30.6338
R753 source.n863 source.n862 30.6338
R754 source.n715 source.n714 30.6338
R755 source.n139 source.n138 30.6338
R756 source.n287 source.n286 30.6338
R757 source.n427 source.n426 30.6338
R758 source.n575 source.n574 30.6338
R759 source.n1152 source.n139 26.3172
R760 source.n1081 source.n1046 13.1884
R761 source.n1128 source.n1127 13.1884
R762 source.n933 source.n898 13.1884
R763 source.n980 source.n979 13.1884
R764 source.n793 source.n758 13.1884
R765 source.n840 source.n839 13.1884
R766 source.n645 source.n610 13.1884
R767 source.n692 source.n691 13.1884
R768 source.n116 source.n115 13.1884
R769 source.n70 source.n35 13.1884
R770 source.n264 source.n263 13.1884
R771 source.n218 source.n183 13.1884
R772 source.n404 source.n403 13.1884
R773 source.n358 source.n323 13.1884
R774 source.n552 source.n551 13.1884
R775 source.n506 source.n471 13.1884
R776 source.n1077 source.n1076 12.8005
R777 source.n1082 source.n1044 12.8005
R778 source.n1126 source.n1024 12.8005
R779 source.n1131 source.n1022 12.8005
R780 source.n929 source.n928 12.8005
R781 source.n934 source.n896 12.8005
R782 source.n978 source.n876 12.8005
R783 source.n983 source.n874 12.8005
R784 source.n789 source.n788 12.8005
R785 source.n794 source.n756 12.8005
R786 source.n838 source.n736 12.8005
R787 source.n843 source.n734 12.8005
R788 source.n641 source.n640 12.8005
R789 source.n646 source.n608 12.8005
R790 source.n690 source.n588 12.8005
R791 source.n695 source.n586 12.8005
R792 source.n119 source.n10 12.8005
R793 source.n114 source.n12 12.8005
R794 source.n71 source.n33 12.8005
R795 source.n66 source.n37 12.8005
R796 source.n267 source.n158 12.8005
R797 source.n262 source.n160 12.8005
R798 source.n219 source.n181 12.8005
R799 source.n214 source.n185 12.8005
R800 source.n407 source.n298 12.8005
R801 source.n402 source.n300 12.8005
R802 source.n359 source.n321 12.8005
R803 source.n354 source.n325 12.8005
R804 source.n555 source.n446 12.8005
R805 source.n550 source.n448 12.8005
R806 source.n507 source.n469 12.8005
R807 source.n502 source.n473 12.8005
R808 source.n1075 source.n1048 12.0247
R809 source.n1086 source.n1085 12.0247
R810 source.n1123 source.n1122 12.0247
R811 source.n1132 source.n1020 12.0247
R812 source.n927 source.n900 12.0247
R813 source.n938 source.n937 12.0247
R814 source.n975 source.n974 12.0247
R815 source.n984 source.n872 12.0247
R816 source.n787 source.n760 12.0247
R817 source.n798 source.n797 12.0247
R818 source.n835 source.n834 12.0247
R819 source.n844 source.n732 12.0247
R820 source.n639 source.n612 12.0247
R821 source.n650 source.n649 12.0247
R822 source.n687 source.n686 12.0247
R823 source.n696 source.n584 12.0247
R824 source.n120 source.n8 12.0247
R825 source.n111 source.n110 12.0247
R826 source.n75 source.n74 12.0247
R827 source.n65 source.n38 12.0247
R828 source.n268 source.n156 12.0247
R829 source.n259 source.n258 12.0247
R830 source.n223 source.n222 12.0247
R831 source.n213 source.n186 12.0247
R832 source.n408 source.n296 12.0247
R833 source.n399 source.n398 12.0247
R834 source.n363 source.n362 12.0247
R835 source.n353 source.n326 12.0247
R836 source.n556 source.n444 12.0247
R837 source.n547 source.n546 12.0247
R838 source.n511 source.n510 12.0247
R839 source.n501 source.n474 12.0247
R840 source.n1072 source.n1071 11.249
R841 source.n1089 source.n1042 11.249
R842 source.n1118 source.n1026 11.249
R843 source.n1136 source.n1135 11.249
R844 source.n924 source.n923 11.249
R845 source.n941 source.n894 11.249
R846 source.n970 source.n878 11.249
R847 source.n988 source.n987 11.249
R848 source.n784 source.n783 11.249
R849 source.n801 source.n754 11.249
R850 source.n830 source.n738 11.249
R851 source.n848 source.n847 11.249
R852 source.n636 source.n635 11.249
R853 source.n653 source.n606 11.249
R854 source.n682 source.n590 11.249
R855 source.n700 source.n699 11.249
R856 source.n124 source.n123 11.249
R857 source.n107 source.n14 11.249
R858 source.n78 source.n31 11.249
R859 source.n62 source.n61 11.249
R860 source.n272 source.n271 11.249
R861 source.n255 source.n162 11.249
R862 source.n226 source.n179 11.249
R863 source.n210 source.n209 11.249
R864 source.n412 source.n411 11.249
R865 source.n395 source.n302 11.249
R866 source.n366 source.n319 11.249
R867 source.n350 source.n349 11.249
R868 source.n560 source.n559 11.249
R869 source.n543 source.n450 11.249
R870 source.n514 source.n467 11.249
R871 source.n498 source.n497 11.249
R872 source.n1068 source.n1050 10.4732
R873 source.n1090 source.n1040 10.4732
R874 source.n1117 source.n1028 10.4732
R875 source.n1139 source.n1018 10.4732
R876 source.n920 source.n902 10.4732
R877 source.n942 source.n892 10.4732
R878 source.n969 source.n880 10.4732
R879 source.n991 source.n870 10.4732
R880 source.n780 source.n762 10.4732
R881 source.n802 source.n752 10.4732
R882 source.n829 source.n740 10.4732
R883 source.n851 source.n730 10.4732
R884 source.n632 source.n614 10.4732
R885 source.n654 source.n604 10.4732
R886 source.n681 source.n592 10.4732
R887 source.n703 source.n582 10.4732
R888 source.n127 source.n6 10.4732
R889 source.n106 source.n17 10.4732
R890 source.n79 source.n29 10.4732
R891 source.n58 source.n40 10.4732
R892 source.n275 source.n154 10.4732
R893 source.n254 source.n165 10.4732
R894 source.n227 source.n177 10.4732
R895 source.n206 source.n188 10.4732
R896 source.n415 source.n294 10.4732
R897 source.n394 source.n305 10.4732
R898 source.n367 source.n317 10.4732
R899 source.n346 source.n328 10.4732
R900 source.n563 source.n442 10.4732
R901 source.n542 source.n453 10.4732
R902 source.n515 source.n465 10.4732
R903 source.n494 source.n476 10.4732
R904 source.n1057 source.n1056 10.2747
R905 source.n909 source.n908 10.2747
R906 source.n769 source.n768 10.2747
R907 source.n621 source.n620 10.2747
R908 source.n47 source.n46 10.2747
R909 source.n195 source.n194 10.2747
R910 source.n335 source.n334 10.2747
R911 source.n483 source.n482 10.2747
R912 source.n1067 source.n1052 9.69747
R913 source.n1094 source.n1093 9.69747
R914 source.n1114 source.n1113 9.69747
R915 source.n1140 source.n1016 9.69747
R916 source.n919 source.n904 9.69747
R917 source.n946 source.n945 9.69747
R918 source.n966 source.n965 9.69747
R919 source.n992 source.n868 9.69747
R920 source.n779 source.n764 9.69747
R921 source.n806 source.n805 9.69747
R922 source.n826 source.n825 9.69747
R923 source.n852 source.n728 9.69747
R924 source.n631 source.n616 9.69747
R925 source.n658 source.n657 9.69747
R926 source.n678 source.n677 9.69747
R927 source.n704 source.n580 9.69747
R928 source.n128 source.n4 9.69747
R929 source.n103 source.n102 9.69747
R930 source.n83 source.n82 9.69747
R931 source.n57 source.n42 9.69747
R932 source.n276 source.n152 9.69747
R933 source.n251 source.n250 9.69747
R934 source.n231 source.n230 9.69747
R935 source.n205 source.n190 9.69747
R936 source.n416 source.n292 9.69747
R937 source.n391 source.n390 9.69747
R938 source.n371 source.n370 9.69747
R939 source.n345 source.n330 9.69747
R940 source.n564 source.n440 9.69747
R941 source.n539 source.n538 9.69747
R942 source.n519 source.n518 9.69747
R943 source.n493 source.n478 9.69747
R944 source.n1150 source.n1149 9.45567
R945 source.n1002 source.n1001 9.45567
R946 source.n862 source.n861 9.45567
R947 source.n714 source.n713 9.45567
R948 source.n138 source.n137 9.45567
R949 source.n286 source.n285 9.45567
R950 source.n426 source.n425 9.45567
R951 source.n574 source.n573 9.45567
R952 source.n1014 source.n1013 9.3005
R953 source.n1143 source.n1142 9.3005
R954 source.n1141 source.n1140 9.3005
R955 source.n1018 source.n1017 9.3005
R956 source.n1135 source.n1134 9.3005
R957 source.n1133 source.n1132 9.3005
R958 source.n1022 source.n1021 9.3005
R959 source.n1101 source.n1100 9.3005
R960 source.n1099 source.n1098 9.3005
R961 source.n1038 source.n1037 9.3005
R962 source.n1093 source.n1092 9.3005
R963 source.n1091 source.n1090 9.3005
R964 source.n1042 source.n1041 9.3005
R965 source.n1085 source.n1084 9.3005
R966 source.n1083 source.n1082 9.3005
R967 source.n1059 source.n1058 9.3005
R968 source.n1054 source.n1053 9.3005
R969 source.n1065 source.n1064 9.3005
R970 source.n1067 source.n1066 9.3005
R971 source.n1050 source.n1049 9.3005
R972 source.n1073 source.n1072 9.3005
R973 source.n1075 source.n1074 9.3005
R974 source.n1076 source.n1045 9.3005
R975 source.n1034 source.n1033 9.3005
R976 source.n1107 source.n1106 9.3005
R977 source.n1109 source.n1108 9.3005
R978 source.n1030 source.n1029 9.3005
R979 source.n1115 source.n1114 9.3005
R980 source.n1117 source.n1116 9.3005
R981 source.n1026 source.n1025 9.3005
R982 source.n1124 source.n1123 9.3005
R983 source.n1126 source.n1125 9.3005
R984 source.n1149 source.n1148 9.3005
R985 source.n866 source.n865 9.3005
R986 source.n995 source.n994 9.3005
R987 source.n993 source.n992 9.3005
R988 source.n870 source.n869 9.3005
R989 source.n987 source.n986 9.3005
R990 source.n985 source.n984 9.3005
R991 source.n874 source.n873 9.3005
R992 source.n953 source.n952 9.3005
R993 source.n951 source.n950 9.3005
R994 source.n890 source.n889 9.3005
R995 source.n945 source.n944 9.3005
R996 source.n943 source.n942 9.3005
R997 source.n894 source.n893 9.3005
R998 source.n937 source.n936 9.3005
R999 source.n935 source.n934 9.3005
R1000 source.n911 source.n910 9.3005
R1001 source.n906 source.n905 9.3005
R1002 source.n917 source.n916 9.3005
R1003 source.n919 source.n918 9.3005
R1004 source.n902 source.n901 9.3005
R1005 source.n925 source.n924 9.3005
R1006 source.n927 source.n926 9.3005
R1007 source.n928 source.n897 9.3005
R1008 source.n886 source.n885 9.3005
R1009 source.n959 source.n958 9.3005
R1010 source.n961 source.n960 9.3005
R1011 source.n882 source.n881 9.3005
R1012 source.n967 source.n966 9.3005
R1013 source.n969 source.n968 9.3005
R1014 source.n878 source.n877 9.3005
R1015 source.n976 source.n975 9.3005
R1016 source.n978 source.n977 9.3005
R1017 source.n1001 source.n1000 9.3005
R1018 source.n726 source.n725 9.3005
R1019 source.n855 source.n854 9.3005
R1020 source.n853 source.n852 9.3005
R1021 source.n730 source.n729 9.3005
R1022 source.n847 source.n846 9.3005
R1023 source.n845 source.n844 9.3005
R1024 source.n734 source.n733 9.3005
R1025 source.n813 source.n812 9.3005
R1026 source.n811 source.n810 9.3005
R1027 source.n750 source.n749 9.3005
R1028 source.n805 source.n804 9.3005
R1029 source.n803 source.n802 9.3005
R1030 source.n754 source.n753 9.3005
R1031 source.n797 source.n796 9.3005
R1032 source.n795 source.n794 9.3005
R1033 source.n771 source.n770 9.3005
R1034 source.n766 source.n765 9.3005
R1035 source.n777 source.n776 9.3005
R1036 source.n779 source.n778 9.3005
R1037 source.n762 source.n761 9.3005
R1038 source.n785 source.n784 9.3005
R1039 source.n787 source.n786 9.3005
R1040 source.n788 source.n757 9.3005
R1041 source.n746 source.n745 9.3005
R1042 source.n819 source.n818 9.3005
R1043 source.n821 source.n820 9.3005
R1044 source.n742 source.n741 9.3005
R1045 source.n827 source.n826 9.3005
R1046 source.n829 source.n828 9.3005
R1047 source.n738 source.n737 9.3005
R1048 source.n836 source.n835 9.3005
R1049 source.n838 source.n837 9.3005
R1050 source.n861 source.n860 9.3005
R1051 source.n578 source.n577 9.3005
R1052 source.n707 source.n706 9.3005
R1053 source.n705 source.n704 9.3005
R1054 source.n582 source.n581 9.3005
R1055 source.n699 source.n698 9.3005
R1056 source.n697 source.n696 9.3005
R1057 source.n586 source.n585 9.3005
R1058 source.n665 source.n664 9.3005
R1059 source.n663 source.n662 9.3005
R1060 source.n602 source.n601 9.3005
R1061 source.n657 source.n656 9.3005
R1062 source.n655 source.n654 9.3005
R1063 source.n606 source.n605 9.3005
R1064 source.n649 source.n648 9.3005
R1065 source.n647 source.n646 9.3005
R1066 source.n623 source.n622 9.3005
R1067 source.n618 source.n617 9.3005
R1068 source.n629 source.n628 9.3005
R1069 source.n631 source.n630 9.3005
R1070 source.n614 source.n613 9.3005
R1071 source.n637 source.n636 9.3005
R1072 source.n639 source.n638 9.3005
R1073 source.n640 source.n609 9.3005
R1074 source.n598 source.n597 9.3005
R1075 source.n671 source.n670 9.3005
R1076 source.n673 source.n672 9.3005
R1077 source.n594 source.n593 9.3005
R1078 source.n679 source.n678 9.3005
R1079 source.n681 source.n680 9.3005
R1080 source.n590 source.n589 9.3005
R1081 source.n688 source.n687 9.3005
R1082 source.n690 source.n689 9.3005
R1083 source.n713 source.n712 9.3005
R1084 source.n49 source.n48 9.3005
R1085 source.n44 source.n43 9.3005
R1086 source.n55 source.n54 9.3005
R1087 source.n57 source.n56 9.3005
R1088 source.n40 source.n39 9.3005
R1089 source.n63 source.n62 9.3005
R1090 source.n65 source.n64 9.3005
R1091 source.n37 source.n34 9.3005
R1092 source.n96 source.n95 9.3005
R1093 source.n98 source.n97 9.3005
R1094 source.n19 source.n18 9.3005
R1095 source.n104 source.n103 9.3005
R1096 source.n106 source.n105 9.3005
R1097 source.n14 source.n13 9.3005
R1098 source.n112 source.n111 9.3005
R1099 source.n114 source.n113 9.3005
R1100 source.n137 source.n136 9.3005
R1101 source.n2 source.n1 9.3005
R1102 source.n131 source.n130 9.3005
R1103 source.n129 source.n128 9.3005
R1104 source.n6 source.n5 9.3005
R1105 source.n123 source.n122 9.3005
R1106 source.n121 source.n120 9.3005
R1107 source.n10 source.n9 9.3005
R1108 source.n23 source.n22 9.3005
R1109 source.n90 source.n89 9.3005
R1110 source.n88 source.n87 9.3005
R1111 source.n27 source.n26 9.3005
R1112 source.n82 source.n81 9.3005
R1113 source.n80 source.n79 9.3005
R1114 source.n31 source.n30 9.3005
R1115 source.n74 source.n73 9.3005
R1116 source.n72 source.n71 9.3005
R1117 source.n197 source.n196 9.3005
R1118 source.n192 source.n191 9.3005
R1119 source.n203 source.n202 9.3005
R1120 source.n205 source.n204 9.3005
R1121 source.n188 source.n187 9.3005
R1122 source.n211 source.n210 9.3005
R1123 source.n213 source.n212 9.3005
R1124 source.n185 source.n182 9.3005
R1125 source.n244 source.n243 9.3005
R1126 source.n246 source.n245 9.3005
R1127 source.n167 source.n166 9.3005
R1128 source.n252 source.n251 9.3005
R1129 source.n254 source.n253 9.3005
R1130 source.n162 source.n161 9.3005
R1131 source.n260 source.n259 9.3005
R1132 source.n262 source.n261 9.3005
R1133 source.n285 source.n284 9.3005
R1134 source.n150 source.n149 9.3005
R1135 source.n279 source.n278 9.3005
R1136 source.n277 source.n276 9.3005
R1137 source.n154 source.n153 9.3005
R1138 source.n271 source.n270 9.3005
R1139 source.n269 source.n268 9.3005
R1140 source.n158 source.n157 9.3005
R1141 source.n171 source.n170 9.3005
R1142 source.n238 source.n237 9.3005
R1143 source.n236 source.n235 9.3005
R1144 source.n175 source.n174 9.3005
R1145 source.n230 source.n229 9.3005
R1146 source.n228 source.n227 9.3005
R1147 source.n179 source.n178 9.3005
R1148 source.n222 source.n221 9.3005
R1149 source.n220 source.n219 9.3005
R1150 source.n337 source.n336 9.3005
R1151 source.n332 source.n331 9.3005
R1152 source.n343 source.n342 9.3005
R1153 source.n345 source.n344 9.3005
R1154 source.n328 source.n327 9.3005
R1155 source.n351 source.n350 9.3005
R1156 source.n353 source.n352 9.3005
R1157 source.n325 source.n322 9.3005
R1158 source.n384 source.n383 9.3005
R1159 source.n386 source.n385 9.3005
R1160 source.n307 source.n306 9.3005
R1161 source.n392 source.n391 9.3005
R1162 source.n394 source.n393 9.3005
R1163 source.n302 source.n301 9.3005
R1164 source.n400 source.n399 9.3005
R1165 source.n402 source.n401 9.3005
R1166 source.n425 source.n424 9.3005
R1167 source.n290 source.n289 9.3005
R1168 source.n419 source.n418 9.3005
R1169 source.n417 source.n416 9.3005
R1170 source.n294 source.n293 9.3005
R1171 source.n411 source.n410 9.3005
R1172 source.n409 source.n408 9.3005
R1173 source.n298 source.n297 9.3005
R1174 source.n311 source.n310 9.3005
R1175 source.n378 source.n377 9.3005
R1176 source.n376 source.n375 9.3005
R1177 source.n315 source.n314 9.3005
R1178 source.n370 source.n369 9.3005
R1179 source.n368 source.n367 9.3005
R1180 source.n319 source.n318 9.3005
R1181 source.n362 source.n361 9.3005
R1182 source.n360 source.n359 9.3005
R1183 source.n485 source.n484 9.3005
R1184 source.n480 source.n479 9.3005
R1185 source.n491 source.n490 9.3005
R1186 source.n493 source.n492 9.3005
R1187 source.n476 source.n475 9.3005
R1188 source.n499 source.n498 9.3005
R1189 source.n501 source.n500 9.3005
R1190 source.n473 source.n470 9.3005
R1191 source.n532 source.n531 9.3005
R1192 source.n534 source.n533 9.3005
R1193 source.n455 source.n454 9.3005
R1194 source.n540 source.n539 9.3005
R1195 source.n542 source.n541 9.3005
R1196 source.n450 source.n449 9.3005
R1197 source.n548 source.n547 9.3005
R1198 source.n550 source.n549 9.3005
R1199 source.n573 source.n572 9.3005
R1200 source.n438 source.n437 9.3005
R1201 source.n567 source.n566 9.3005
R1202 source.n565 source.n564 9.3005
R1203 source.n442 source.n441 9.3005
R1204 source.n559 source.n558 9.3005
R1205 source.n557 source.n556 9.3005
R1206 source.n446 source.n445 9.3005
R1207 source.n459 source.n458 9.3005
R1208 source.n526 source.n525 9.3005
R1209 source.n524 source.n523 9.3005
R1210 source.n463 source.n462 9.3005
R1211 source.n518 source.n517 9.3005
R1212 source.n516 source.n515 9.3005
R1213 source.n467 source.n466 9.3005
R1214 source.n510 source.n509 9.3005
R1215 source.n508 source.n507 9.3005
R1216 source.n1064 source.n1063 8.92171
R1217 source.n1097 source.n1038 8.92171
R1218 source.n1110 source.n1030 8.92171
R1219 source.n1144 source.n1143 8.92171
R1220 source.n916 source.n915 8.92171
R1221 source.n949 source.n890 8.92171
R1222 source.n962 source.n882 8.92171
R1223 source.n996 source.n995 8.92171
R1224 source.n776 source.n775 8.92171
R1225 source.n809 source.n750 8.92171
R1226 source.n822 source.n742 8.92171
R1227 source.n856 source.n855 8.92171
R1228 source.n628 source.n627 8.92171
R1229 source.n661 source.n602 8.92171
R1230 source.n674 source.n594 8.92171
R1231 source.n708 source.n707 8.92171
R1232 source.n132 source.n131 8.92171
R1233 source.n99 source.n19 8.92171
R1234 source.n86 source.n27 8.92171
R1235 source.n54 source.n53 8.92171
R1236 source.n280 source.n279 8.92171
R1237 source.n247 source.n167 8.92171
R1238 source.n234 source.n175 8.92171
R1239 source.n202 source.n201 8.92171
R1240 source.n420 source.n419 8.92171
R1241 source.n387 source.n307 8.92171
R1242 source.n374 source.n315 8.92171
R1243 source.n342 source.n341 8.92171
R1244 source.n568 source.n567 8.92171
R1245 source.n535 source.n455 8.92171
R1246 source.n522 source.n463 8.92171
R1247 source.n490 source.n489 8.92171
R1248 source.n1060 source.n1054 8.14595
R1249 source.n1098 source.n1036 8.14595
R1250 source.n1109 source.n1032 8.14595
R1251 source.n1147 source.n1014 8.14595
R1252 source.n912 source.n906 8.14595
R1253 source.n950 source.n888 8.14595
R1254 source.n961 source.n884 8.14595
R1255 source.n999 source.n866 8.14595
R1256 source.n772 source.n766 8.14595
R1257 source.n810 source.n748 8.14595
R1258 source.n821 source.n744 8.14595
R1259 source.n859 source.n726 8.14595
R1260 source.n624 source.n618 8.14595
R1261 source.n662 source.n600 8.14595
R1262 source.n673 source.n596 8.14595
R1263 source.n711 source.n578 8.14595
R1264 source.n135 source.n2 8.14595
R1265 source.n98 source.n21 8.14595
R1266 source.n87 source.n25 8.14595
R1267 source.n50 source.n44 8.14595
R1268 source.n283 source.n150 8.14595
R1269 source.n246 source.n169 8.14595
R1270 source.n235 source.n173 8.14595
R1271 source.n198 source.n192 8.14595
R1272 source.n423 source.n290 8.14595
R1273 source.n386 source.n309 8.14595
R1274 source.n375 source.n313 8.14595
R1275 source.n338 source.n332 8.14595
R1276 source.n571 source.n438 8.14595
R1277 source.n534 source.n457 8.14595
R1278 source.n523 source.n461 8.14595
R1279 source.n486 source.n480 8.14595
R1280 source.n1059 source.n1056 7.3702
R1281 source.n1102 source.n1101 7.3702
R1282 source.n1106 source.n1105 7.3702
R1283 source.n1148 source.n1012 7.3702
R1284 source.n911 source.n908 7.3702
R1285 source.n954 source.n953 7.3702
R1286 source.n958 source.n957 7.3702
R1287 source.n1000 source.n864 7.3702
R1288 source.n771 source.n768 7.3702
R1289 source.n814 source.n813 7.3702
R1290 source.n818 source.n817 7.3702
R1291 source.n860 source.n724 7.3702
R1292 source.n623 source.n620 7.3702
R1293 source.n666 source.n665 7.3702
R1294 source.n670 source.n669 7.3702
R1295 source.n712 source.n576 7.3702
R1296 source.n136 source.n0 7.3702
R1297 source.n95 source.n94 7.3702
R1298 source.n91 source.n90 7.3702
R1299 source.n49 source.n46 7.3702
R1300 source.n284 source.n148 7.3702
R1301 source.n243 source.n242 7.3702
R1302 source.n239 source.n238 7.3702
R1303 source.n197 source.n194 7.3702
R1304 source.n424 source.n288 7.3702
R1305 source.n383 source.n382 7.3702
R1306 source.n379 source.n378 7.3702
R1307 source.n337 source.n334 7.3702
R1308 source.n572 source.n436 7.3702
R1309 source.n531 source.n530 7.3702
R1310 source.n527 source.n526 7.3702
R1311 source.n485 source.n482 7.3702
R1312 source.n1102 source.n1034 6.59444
R1313 source.n1105 source.n1034 6.59444
R1314 source.n1150 source.n1012 6.59444
R1315 source.n954 source.n886 6.59444
R1316 source.n957 source.n886 6.59444
R1317 source.n1002 source.n864 6.59444
R1318 source.n814 source.n746 6.59444
R1319 source.n817 source.n746 6.59444
R1320 source.n862 source.n724 6.59444
R1321 source.n666 source.n598 6.59444
R1322 source.n669 source.n598 6.59444
R1323 source.n714 source.n576 6.59444
R1324 source.n138 source.n0 6.59444
R1325 source.n94 source.n23 6.59444
R1326 source.n91 source.n23 6.59444
R1327 source.n286 source.n148 6.59444
R1328 source.n242 source.n171 6.59444
R1329 source.n239 source.n171 6.59444
R1330 source.n426 source.n288 6.59444
R1331 source.n382 source.n311 6.59444
R1332 source.n379 source.n311 6.59444
R1333 source.n574 source.n436 6.59444
R1334 source.n530 source.n459 6.59444
R1335 source.n527 source.n459 6.59444
R1336 source.n1060 source.n1059 5.81868
R1337 source.n1101 source.n1036 5.81868
R1338 source.n1106 source.n1032 5.81868
R1339 source.n1148 source.n1147 5.81868
R1340 source.n912 source.n911 5.81868
R1341 source.n953 source.n888 5.81868
R1342 source.n958 source.n884 5.81868
R1343 source.n1000 source.n999 5.81868
R1344 source.n772 source.n771 5.81868
R1345 source.n813 source.n748 5.81868
R1346 source.n818 source.n744 5.81868
R1347 source.n860 source.n859 5.81868
R1348 source.n624 source.n623 5.81868
R1349 source.n665 source.n600 5.81868
R1350 source.n670 source.n596 5.81868
R1351 source.n712 source.n711 5.81868
R1352 source.n136 source.n135 5.81868
R1353 source.n95 source.n21 5.81868
R1354 source.n90 source.n25 5.81868
R1355 source.n50 source.n49 5.81868
R1356 source.n284 source.n283 5.81868
R1357 source.n243 source.n169 5.81868
R1358 source.n238 source.n173 5.81868
R1359 source.n198 source.n197 5.81868
R1360 source.n424 source.n423 5.81868
R1361 source.n383 source.n309 5.81868
R1362 source.n378 source.n313 5.81868
R1363 source.n338 source.n337 5.81868
R1364 source.n572 source.n571 5.81868
R1365 source.n531 source.n457 5.81868
R1366 source.n526 source.n461 5.81868
R1367 source.n486 source.n485 5.81868
R1368 source.n1152 source.n1151 5.7074
R1369 source.n1063 source.n1054 5.04292
R1370 source.n1098 source.n1097 5.04292
R1371 source.n1110 source.n1109 5.04292
R1372 source.n1144 source.n1014 5.04292
R1373 source.n915 source.n906 5.04292
R1374 source.n950 source.n949 5.04292
R1375 source.n962 source.n961 5.04292
R1376 source.n996 source.n866 5.04292
R1377 source.n775 source.n766 5.04292
R1378 source.n810 source.n809 5.04292
R1379 source.n822 source.n821 5.04292
R1380 source.n856 source.n726 5.04292
R1381 source.n627 source.n618 5.04292
R1382 source.n662 source.n661 5.04292
R1383 source.n674 source.n673 5.04292
R1384 source.n708 source.n578 5.04292
R1385 source.n132 source.n2 5.04292
R1386 source.n99 source.n98 5.04292
R1387 source.n87 source.n86 5.04292
R1388 source.n53 source.n44 5.04292
R1389 source.n280 source.n150 5.04292
R1390 source.n247 source.n246 5.04292
R1391 source.n235 source.n234 5.04292
R1392 source.n201 source.n192 5.04292
R1393 source.n420 source.n290 5.04292
R1394 source.n387 source.n386 5.04292
R1395 source.n375 source.n374 5.04292
R1396 source.n341 source.n332 5.04292
R1397 source.n568 source.n438 5.04292
R1398 source.n535 source.n534 5.04292
R1399 source.n523 source.n522 5.04292
R1400 source.n489 source.n480 5.04292
R1401 source.n1064 source.n1052 4.26717
R1402 source.n1094 source.n1038 4.26717
R1403 source.n1113 source.n1030 4.26717
R1404 source.n1143 source.n1016 4.26717
R1405 source.n916 source.n904 4.26717
R1406 source.n946 source.n890 4.26717
R1407 source.n965 source.n882 4.26717
R1408 source.n995 source.n868 4.26717
R1409 source.n776 source.n764 4.26717
R1410 source.n806 source.n750 4.26717
R1411 source.n825 source.n742 4.26717
R1412 source.n855 source.n728 4.26717
R1413 source.n628 source.n616 4.26717
R1414 source.n658 source.n602 4.26717
R1415 source.n677 source.n594 4.26717
R1416 source.n707 source.n580 4.26717
R1417 source.n131 source.n4 4.26717
R1418 source.n102 source.n19 4.26717
R1419 source.n83 source.n27 4.26717
R1420 source.n54 source.n42 4.26717
R1421 source.n279 source.n152 4.26717
R1422 source.n250 source.n167 4.26717
R1423 source.n231 source.n175 4.26717
R1424 source.n202 source.n190 4.26717
R1425 source.n419 source.n292 4.26717
R1426 source.n390 source.n307 4.26717
R1427 source.n371 source.n315 4.26717
R1428 source.n342 source.n330 4.26717
R1429 source.n567 source.n440 4.26717
R1430 source.n538 source.n455 4.26717
R1431 source.n519 source.n463 4.26717
R1432 source.n490 source.n478 4.26717
R1433 source.n1068 source.n1067 3.49141
R1434 source.n1093 source.n1040 3.49141
R1435 source.n1114 source.n1028 3.49141
R1436 source.n1140 source.n1139 3.49141
R1437 source.n920 source.n919 3.49141
R1438 source.n945 source.n892 3.49141
R1439 source.n966 source.n880 3.49141
R1440 source.n992 source.n991 3.49141
R1441 source.n780 source.n779 3.49141
R1442 source.n805 source.n752 3.49141
R1443 source.n826 source.n740 3.49141
R1444 source.n852 source.n851 3.49141
R1445 source.n632 source.n631 3.49141
R1446 source.n657 source.n604 3.49141
R1447 source.n678 source.n592 3.49141
R1448 source.n704 source.n703 3.49141
R1449 source.n128 source.n127 3.49141
R1450 source.n103 source.n17 3.49141
R1451 source.n82 source.n29 3.49141
R1452 source.n58 source.n57 3.49141
R1453 source.n276 source.n275 3.49141
R1454 source.n251 source.n165 3.49141
R1455 source.n230 source.n177 3.49141
R1456 source.n206 source.n205 3.49141
R1457 source.n416 source.n415 3.49141
R1458 source.n391 source.n305 3.49141
R1459 source.n370 source.n317 3.49141
R1460 source.n346 source.n345 3.49141
R1461 source.n564 source.n563 3.49141
R1462 source.n539 source.n453 3.49141
R1463 source.n518 source.n465 3.49141
R1464 source.n494 source.n493 3.49141
R1465 source.n48 source.n47 2.84303
R1466 source.n196 source.n195 2.84303
R1467 source.n336 source.n335 2.84303
R1468 source.n484 source.n483 2.84303
R1469 source.n1058 source.n1057 2.84303
R1470 source.n910 source.n909 2.84303
R1471 source.n770 source.n769 2.84303
R1472 source.n622 source.n621 2.84303
R1473 source.n1071 source.n1050 2.71565
R1474 source.n1090 source.n1089 2.71565
R1475 source.n1118 source.n1117 2.71565
R1476 source.n1136 source.n1018 2.71565
R1477 source.n923 source.n902 2.71565
R1478 source.n942 source.n941 2.71565
R1479 source.n970 source.n969 2.71565
R1480 source.n988 source.n870 2.71565
R1481 source.n783 source.n762 2.71565
R1482 source.n802 source.n801 2.71565
R1483 source.n830 source.n829 2.71565
R1484 source.n848 source.n730 2.71565
R1485 source.n635 source.n614 2.71565
R1486 source.n654 source.n653 2.71565
R1487 source.n682 source.n681 2.71565
R1488 source.n700 source.n582 2.71565
R1489 source.n124 source.n6 2.71565
R1490 source.n107 source.n106 2.71565
R1491 source.n79 source.n78 2.71565
R1492 source.n61 source.n40 2.71565
R1493 source.n272 source.n154 2.71565
R1494 source.n255 source.n254 2.71565
R1495 source.n227 source.n226 2.71565
R1496 source.n209 source.n188 2.71565
R1497 source.n412 source.n294 2.71565
R1498 source.n395 source.n394 2.71565
R1499 source.n367 source.n366 2.71565
R1500 source.n349 source.n328 2.71565
R1501 source.n560 source.n442 2.71565
R1502 source.n543 source.n542 2.71565
R1503 source.n515 source.n514 2.71565
R1504 source.n497 source.n476 2.71565
R1505 source.n1072 source.n1048 1.93989
R1506 source.n1086 source.n1042 1.93989
R1507 source.n1122 source.n1026 1.93989
R1508 source.n1135 source.n1020 1.93989
R1509 source.n924 source.n900 1.93989
R1510 source.n938 source.n894 1.93989
R1511 source.n974 source.n878 1.93989
R1512 source.n987 source.n872 1.93989
R1513 source.n784 source.n760 1.93989
R1514 source.n798 source.n754 1.93989
R1515 source.n834 source.n738 1.93989
R1516 source.n847 source.n732 1.93989
R1517 source.n636 source.n612 1.93989
R1518 source.n650 source.n606 1.93989
R1519 source.n686 source.n590 1.93989
R1520 source.n699 source.n584 1.93989
R1521 source.n123 source.n8 1.93989
R1522 source.n110 source.n14 1.93989
R1523 source.n75 source.n31 1.93989
R1524 source.n62 source.n38 1.93989
R1525 source.n271 source.n156 1.93989
R1526 source.n258 source.n162 1.93989
R1527 source.n223 source.n179 1.93989
R1528 source.n210 source.n186 1.93989
R1529 source.n411 source.n296 1.93989
R1530 source.n398 source.n302 1.93989
R1531 source.n363 source.n319 1.93989
R1532 source.n350 source.n326 1.93989
R1533 source.n559 source.n444 1.93989
R1534 source.n546 source.n450 1.93989
R1535 source.n511 source.n467 1.93989
R1536 source.n498 source.n474 1.93989
R1537 source.n1077 source.n1075 1.16414
R1538 source.n1085 source.n1044 1.16414
R1539 source.n1123 source.n1024 1.16414
R1540 source.n1132 source.n1131 1.16414
R1541 source.n929 source.n927 1.16414
R1542 source.n937 source.n896 1.16414
R1543 source.n975 source.n876 1.16414
R1544 source.n984 source.n983 1.16414
R1545 source.n789 source.n787 1.16414
R1546 source.n797 source.n756 1.16414
R1547 source.n835 source.n736 1.16414
R1548 source.n844 source.n843 1.16414
R1549 source.n641 source.n639 1.16414
R1550 source.n649 source.n608 1.16414
R1551 source.n687 source.n588 1.16414
R1552 source.n696 source.n695 1.16414
R1553 source.n120 source.n119 1.16414
R1554 source.n111 source.n12 1.16414
R1555 source.n74 source.n33 1.16414
R1556 source.n66 source.n65 1.16414
R1557 source.n268 source.n267 1.16414
R1558 source.n259 source.n160 1.16414
R1559 source.n222 source.n181 1.16414
R1560 source.n214 source.n213 1.16414
R1561 source.n408 source.n407 1.16414
R1562 source.n399 source.n300 1.16414
R1563 source.n362 source.n321 1.16414
R1564 source.n354 source.n353 1.16414
R1565 source.n556 source.n555 1.16414
R1566 source.n547 source.n448 1.16414
R1567 source.n510 source.n469 1.16414
R1568 source.n502 source.n501 1.16414
R1569 source.n575 source.n435 0.888431
R1570 source.n435 source.n433 0.888431
R1571 source.n433 source.n431 0.888431
R1572 source.n431 source.n429 0.888431
R1573 source.n429 source.n427 0.888431
R1574 source.n287 source.n147 0.888431
R1575 source.n147 source.n145 0.888431
R1576 source.n145 source.n143 0.888431
R1577 source.n143 source.n141 0.888431
R1578 source.n141 source.n139 0.888431
R1579 source.n717 source.n715 0.888431
R1580 source.n719 source.n717 0.888431
R1581 source.n721 source.n719 0.888431
R1582 source.n723 source.n721 0.888431
R1583 source.n863 source.n723 0.888431
R1584 source.n1005 source.n1003 0.888431
R1585 source.n1007 source.n1005 0.888431
R1586 source.n1009 source.n1007 0.888431
R1587 source.n1011 source.n1009 0.888431
R1588 source.n1151 source.n1011 0.888431
R1589 source.n1010 source.t25 0.7925
R1590 source.n1010 source.t26 0.7925
R1591 source.n1008 source.t22 0.7925
R1592 source.n1008 source.t21 0.7925
R1593 source.n1006 source.t37 0.7925
R1594 source.n1006 source.t35 0.7925
R1595 source.n1004 source.t34 0.7925
R1596 source.n1004 source.t38 0.7925
R1597 source.n722 source.t7 0.7925
R1598 source.n722 source.t9 0.7925
R1599 source.n720 source.t15 0.7925
R1600 source.n720 source.t39 0.7925
R1601 source.n718 source.t10 0.7925
R1602 source.n718 source.t3 0.7925
R1603 source.n716 source.t14 0.7925
R1604 source.n716 source.t1 0.7925
R1605 source.n140 source.t4 0.7925
R1606 source.n140 source.t11 0.7925
R1607 source.n142 source.t6 0.7925
R1608 source.n142 source.t17 0.7925
R1609 source.n144 source.t12 0.7925
R1610 source.n144 source.t18 0.7925
R1611 source.n146 source.t13 0.7925
R1612 source.n146 source.t0 0.7925
R1613 source.n428 source.t28 0.7925
R1614 source.n428 source.t36 0.7925
R1615 source.n430 source.t29 0.7925
R1616 source.n430 source.t20 0.7925
R1617 source.n432 source.t30 0.7925
R1618 source.n432 source.t19 0.7925
R1619 source.n434 source.t32 0.7925
R1620 source.n434 source.t23 0.7925
R1621 source.n427 source.n287 0.470328
R1622 source.n1003 source.n863 0.470328
R1623 source.n1076 source.n1046 0.388379
R1624 source.n1082 source.n1081 0.388379
R1625 source.n1127 source.n1126 0.388379
R1626 source.n1128 source.n1022 0.388379
R1627 source.n928 source.n898 0.388379
R1628 source.n934 source.n933 0.388379
R1629 source.n979 source.n978 0.388379
R1630 source.n980 source.n874 0.388379
R1631 source.n788 source.n758 0.388379
R1632 source.n794 source.n793 0.388379
R1633 source.n839 source.n838 0.388379
R1634 source.n840 source.n734 0.388379
R1635 source.n640 source.n610 0.388379
R1636 source.n646 source.n645 0.388379
R1637 source.n691 source.n690 0.388379
R1638 source.n692 source.n586 0.388379
R1639 source.n116 source.n10 0.388379
R1640 source.n115 source.n114 0.388379
R1641 source.n71 source.n70 0.388379
R1642 source.n37 source.n35 0.388379
R1643 source.n264 source.n158 0.388379
R1644 source.n263 source.n262 0.388379
R1645 source.n219 source.n218 0.388379
R1646 source.n185 source.n183 0.388379
R1647 source.n404 source.n298 0.388379
R1648 source.n403 source.n402 0.388379
R1649 source.n359 source.n358 0.388379
R1650 source.n325 source.n323 0.388379
R1651 source.n552 source.n446 0.388379
R1652 source.n551 source.n550 0.388379
R1653 source.n507 source.n506 0.388379
R1654 source.n473 source.n471 0.388379
R1655 source source.n1152 0.188
R1656 source.n1058 source.n1053 0.155672
R1657 source.n1065 source.n1053 0.155672
R1658 source.n1066 source.n1065 0.155672
R1659 source.n1066 source.n1049 0.155672
R1660 source.n1073 source.n1049 0.155672
R1661 source.n1074 source.n1073 0.155672
R1662 source.n1074 source.n1045 0.155672
R1663 source.n1083 source.n1045 0.155672
R1664 source.n1084 source.n1083 0.155672
R1665 source.n1084 source.n1041 0.155672
R1666 source.n1091 source.n1041 0.155672
R1667 source.n1092 source.n1091 0.155672
R1668 source.n1092 source.n1037 0.155672
R1669 source.n1099 source.n1037 0.155672
R1670 source.n1100 source.n1099 0.155672
R1671 source.n1100 source.n1033 0.155672
R1672 source.n1107 source.n1033 0.155672
R1673 source.n1108 source.n1107 0.155672
R1674 source.n1108 source.n1029 0.155672
R1675 source.n1115 source.n1029 0.155672
R1676 source.n1116 source.n1115 0.155672
R1677 source.n1116 source.n1025 0.155672
R1678 source.n1124 source.n1025 0.155672
R1679 source.n1125 source.n1124 0.155672
R1680 source.n1125 source.n1021 0.155672
R1681 source.n1133 source.n1021 0.155672
R1682 source.n1134 source.n1133 0.155672
R1683 source.n1134 source.n1017 0.155672
R1684 source.n1141 source.n1017 0.155672
R1685 source.n1142 source.n1141 0.155672
R1686 source.n1142 source.n1013 0.155672
R1687 source.n1149 source.n1013 0.155672
R1688 source.n910 source.n905 0.155672
R1689 source.n917 source.n905 0.155672
R1690 source.n918 source.n917 0.155672
R1691 source.n918 source.n901 0.155672
R1692 source.n925 source.n901 0.155672
R1693 source.n926 source.n925 0.155672
R1694 source.n926 source.n897 0.155672
R1695 source.n935 source.n897 0.155672
R1696 source.n936 source.n935 0.155672
R1697 source.n936 source.n893 0.155672
R1698 source.n943 source.n893 0.155672
R1699 source.n944 source.n943 0.155672
R1700 source.n944 source.n889 0.155672
R1701 source.n951 source.n889 0.155672
R1702 source.n952 source.n951 0.155672
R1703 source.n952 source.n885 0.155672
R1704 source.n959 source.n885 0.155672
R1705 source.n960 source.n959 0.155672
R1706 source.n960 source.n881 0.155672
R1707 source.n967 source.n881 0.155672
R1708 source.n968 source.n967 0.155672
R1709 source.n968 source.n877 0.155672
R1710 source.n976 source.n877 0.155672
R1711 source.n977 source.n976 0.155672
R1712 source.n977 source.n873 0.155672
R1713 source.n985 source.n873 0.155672
R1714 source.n986 source.n985 0.155672
R1715 source.n986 source.n869 0.155672
R1716 source.n993 source.n869 0.155672
R1717 source.n994 source.n993 0.155672
R1718 source.n994 source.n865 0.155672
R1719 source.n1001 source.n865 0.155672
R1720 source.n770 source.n765 0.155672
R1721 source.n777 source.n765 0.155672
R1722 source.n778 source.n777 0.155672
R1723 source.n778 source.n761 0.155672
R1724 source.n785 source.n761 0.155672
R1725 source.n786 source.n785 0.155672
R1726 source.n786 source.n757 0.155672
R1727 source.n795 source.n757 0.155672
R1728 source.n796 source.n795 0.155672
R1729 source.n796 source.n753 0.155672
R1730 source.n803 source.n753 0.155672
R1731 source.n804 source.n803 0.155672
R1732 source.n804 source.n749 0.155672
R1733 source.n811 source.n749 0.155672
R1734 source.n812 source.n811 0.155672
R1735 source.n812 source.n745 0.155672
R1736 source.n819 source.n745 0.155672
R1737 source.n820 source.n819 0.155672
R1738 source.n820 source.n741 0.155672
R1739 source.n827 source.n741 0.155672
R1740 source.n828 source.n827 0.155672
R1741 source.n828 source.n737 0.155672
R1742 source.n836 source.n737 0.155672
R1743 source.n837 source.n836 0.155672
R1744 source.n837 source.n733 0.155672
R1745 source.n845 source.n733 0.155672
R1746 source.n846 source.n845 0.155672
R1747 source.n846 source.n729 0.155672
R1748 source.n853 source.n729 0.155672
R1749 source.n854 source.n853 0.155672
R1750 source.n854 source.n725 0.155672
R1751 source.n861 source.n725 0.155672
R1752 source.n622 source.n617 0.155672
R1753 source.n629 source.n617 0.155672
R1754 source.n630 source.n629 0.155672
R1755 source.n630 source.n613 0.155672
R1756 source.n637 source.n613 0.155672
R1757 source.n638 source.n637 0.155672
R1758 source.n638 source.n609 0.155672
R1759 source.n647 source.n609 0.155672
R1760 source.n648 source.n647 0.155672
R1761 source.n648 source.n605 0.155672
R1762 source.n655 source.n605 0.155672
R1763 source.n656 source.n655 0.155672
R1764 source.n656 source.n601 0.155672
R1765 source.n663 source.n601 0.155672
R1766 source.n664 source.n663 0.155672
R1767 source.n664 source.n597 0.155672
R1768 source.n671 source.n597 0.155672
R1769 source.n672 source.n671 0.155672
R1770 source.n672 source.n593 0.155672
R1771 source.n679 source.n593 0.155672
R1772 source.n680 source.n679 0.155672
R1773 source.n680 source.n589 0.155672
R1774 source.n688 source.n589 0.155672
R1775 source.n689 source.n688 0.155672
R1776 source.n689 source.n585 0.155672
R1777 source.n697 source.n585 0.155672
R1778 source.n698 source.n697 0.155672
R1779 source.n698 source.n581 0.155672
R1780 source.n705 source.n581 0.155672
R1781 source.n706 source.n705 0.155672
R1782 source.n706 source.n577 0.155672
R1783 source.n713 source.n577 0.155672
R1784 source.n137 source.n1 0.155672
R1785 source.n130 source.n1 0.155672
R1786 source.n130 source.n129 0.155672
R1787 source.n129 source.n5 0.155672
R1788 source.n122 source.n5 0.155672
R1789 source.n122 source.n121 0.155672
R1790 source.n121 source.n9 0.155672
R1791 source.n113 source.n9 0.155672
R1792 source.n113 source.n112 0.155672
R1793 source.n112 source.n13 0.155672
R1794 source.n105 source.n13 0.155672
R1795 source.n105 source.n104 0.155672
R1796 source.n104 source.n18 0.155672
R1797 source.n97 source.n18 0.155672
R1798 source.n97 source.n96 0.155672
R1799 source.n96 source.n22 0.155672
R1800 source.n89 source.n22 0.155672
R1801 source.n89 source.n88 0.155672
R1802 source.n88 source.n26 0.155672
R1803 source.n81 source.n26 0.155672
R1804 source.n81 source.n80 0.155672
R1805 source.n80 source.n30 0.155672
R1806 source.n73 source.n30 0.155672
R1807 source.n73 source.n72 0.155672
R1808 source.n72 source.n34 0.155672
R1809 source.n64 source.n34 0.155672
R1810 source.n64 source.n63 0.155672
R1811 source.n63 source.n39 0.155672
R1812 source.n56 source.n39 0.155672
R1813 source.n56 source.n55 0.155672
R1814 source.n55 source.n43 0.155672
R1815 source.n48 source.n43 0.155672
R1816 source.n285 source.n149 0.155672
R1817 source.n278 source.n149 0.155672
R1818 source.n278 source.n277 0.155672
R1819 source.n277 source.n153 0.155672
R1820 source.n270 source.n153 0.155672
R1821 source.n270 source.n269 0.155672
R1822 source.n269 source.n157 0.155672
R1823 source.n261 source.n157 0.155672
R1824 source.n261 source.n260 0.155672
R1825 source.n260 source.n161 0.155672
R1826 source.n253 source.n161 0.155672
R1827 source.n253 source.n252 0.155672
R1828 source.n252 source.n166 0.155672
R1829 source.n245 source.n166 0.155672
R1830 source.n245 source.n244 0.155672
R1831 source.n244 source.n170 0.155672
R1832 source.n237 source.n170 0.155672
R1833 source.n237 source.n236 0.155672
R1834 source.n236 source.n174 0.155672
R1835 source.n229 source.n174 0.155672
R1836 source.n229 source.n228 0.155672
R1837 source.n228 source.n178 0.155672
R1838 source.n221 source.n178 0.155672
R1839 source.n221 source.n220 0.155672
R1840 source.n220 source.n182 0.155672
R1841 source.n212 source.n182 0.155672
R1842 source.n212 source.n211 0.155672
R1843 source.n211 source.n187 0.155672
R1844 source.n204 source.n187 0.155672
R1845 source.n204 source.n203 0.155672
R1846 source.n203 source.n191 0.155672
R1847 source.n196 source.n191 0.155672
R1848 source.n425 source.n289 0.155672
R1849 source.n418 source.n289 0.155672
R1850 source.n418 source.n417 0.155672
R1851 source.n417 source.n293 0.155672
R1852 source.n410 source.n293 0.155672
R1853 source.n410 source.n409 0.155672
R1854 source.n409 source.n297 0.155672
R1855 source.n401 source.n297 0.155672
R1856 source.n401 source.n400 0.155672
R1857 source.n400 source.n301 0.155672
R1858 source.n393 source.n301 0.155672
R1859 source.n393 source.n392 0.155672
R1860 source.n392 source.n306 0.155672
R1861 source.n385 source.n306 0.155672
R1862 source.n385 source.n384 0.155672
R1863 source.n384 source.n310 0.155672
R1864 source.n377 source.n310 0.155672
R1865 source.n377 source.n376 0.155672
R1866 source.n376 source.n314 0.155672
R1867 source.n369 source.n314 0.155672
R1868 source.n369 source.n368 0.155672
R1869 source.n368 source.n318 0.155672
R1870 source.n361 source.n318 0.155672
R1871 source.n361 source.n360 0.155672
R1872 source.n360 source.n322 0.155672
R1873 source.n352 source.n322 0.155672
R1874 source.n352 source.n351 0.155672
R1875 source.n351 source.n327 0.155672
R1876 source.n344 source.n327 0.155672
R1877 source.n344 source.n343 0.155672
R1878 source.n343 source.n331 0.155672
R1879 source.n336 source.n331 0.155672
R1880 source.n573 source.n437 0.155672
R1881 source.n566 source.n437 0.155672
R1882 source.n566 source.n565 0.155672
R1883 source.n565 source.n441 0.155672
R1884 source.n558 source.n441 0.155672
R1885 source.n558 source.n557 0.155672
R1886 source.n557 source.n445 0.155672
R1887 source.n549 source.n445 0.155672
R1888 source.n549 source.n548 0.155672
R1889 source.n548 source.n449 0.155672
R1890 source.n541 source.n449 0.155672
R1891 source.n541 source.n540 0.155672
R1892 source.n540 source.n454 0.155672
R1893 source.n533 source.n454 0.155672
R1894 source.n533 source.n532 0.155672
R1895 source.n532 source.n458 0.155672
R1896 source.n525 source.n458 0.155672
R1897 source.n525 source.n524 0.155672
R1898 source.n524 source.n462 0.155672
R1899 source.n517 source.n462 0.155672
R1900 source.n517 source.n516 0.155672
R1901 source.n516 source.n466 0.155672
R1902 source.n509 source.n466 0.155672
R1903 source.n509 source.n508 0.155672
R1904 source.n508 source.n470 0.155672
R1905 source.n500 source.n470 0.155672
R1906 source.n500 source.n499 0.155672
R1907 source.n499 source.n475 0.155672
R1908 source.n492 source.n475 0.155672
R1909 source.n492 source.n491 0.155672
R1910 source.n491 source.n479 0.155672
R1911 source.n484 source.n479 0.155672
R1912 plus.n9 plus.t6 942.226
R1913 plus.n43 plus.t19 942.226
R1914 plus.n32 plus.t3 916.833
R1915 plus.n30 plus.t18 916.833
R1916 plus.n2 plus.t8 916.833
R1917 plus.n24 plus.t1 916.833
R1918 plus.n4 plus.t12 916.833
R1919 plus.n18 plus.t5 916.833
R1920 plus.n6 plus.t10 916.833
R1921 plus.n12 plus.t2 916.833
R1922 plus.n8 plus.t13 916.833
R1923 plus.n66 plus.t15 916.833
R1924 plus.n64 plus.t14 916.833
R1925 plus.n36 plus.t17 916.833
R1926 plus.n58 plus.t7 916.833
R1927 plus.n38 plus.t4 916.833
R1928 plus.n52 plus.t11 916.833
R1929 plus.n40 plus.t9 916.833
R1930 plus.n46 plus.t16 916.833
R1931 plus.n42 plus.t0 916.833
R1932 plus.n11 plus.n10 161.3
R1933 plus.n12 plus.n7 161.3
R1934 plus.n14 plus.n13 161.3
R1935 plus.n15 plus.n6 161.3
R1936 plus.n17 plus.n16 161.3
R1937 plus.n18 plus.n5 161.3
R1938 plus.n20 plus.n19 161.3
R1939 plus.n21 plus.n4 161.3
R1940 plus.n23 plus.n22 161.3
R1941 plus.n24 plus.n3 161.3
R1942 plus.n26 plus.n25 161.3
R1943 plus.n27 plus.n2 161.3
R1944 plus.n29 plus.n28 161.3
R1945 plus.n30 plus.n1 161.3
R1946 plus.n31 plus.n0 161.3
R1947 plus.n33 plus.n32 161.3
R1948 plus.n45 plus.n44 161.3
R1949 plus.n46 plus.n41 161.3
R1950 plus.n48 plus.n47 161.3
R1951 plus.n49 plus.n40 161.3
R1952 plus.n51 plus.n50 161.3
R1953 plus.n52 plus.n39 161.3
R1954 plus.n54 plus.n53 161.3
R1955 plus.n55 plus.n38 161.3
R1956 plus.n57 plus.n56 161.3
R1957 plus.n58 plus.n37 161.3
R1958 plus.n60 plus.n59 161.3
R1959 plus.n61 plus.n36 161.3
R1960 plus.n63 plus.n62 161.3
R1961 plus.n64 plus.n35 161.3
R1962 plus.n65 plus.n34 161.3
R1963 plus.n67 plus.n66 161.3
R1964 plus.n10 plus.n9 45.0031
R1965 plus.n44 plus.n43 45.0031
R1966 plus.n32 plus.n31 41.6278
R1967 plus.n66 plus.n65 41.6278
R1968 plus plus.n67 39.3892
R1969 plus.n30 plus.n29 37.246
R1970 plus.n11 plus.n8 37.246
R1971 plus.n64 plus.n63 37.246
R1972 plus.n45 plus.n42 37.246
R1973 plus.n25 plus.n2 32.8641
R1974 plus.n13 plus.n12 32.8641
R1975 plus.n59 plus.n36 32.8641
R1976 plus.n47 plus.n46 32.8641
R1977 plus.n24 plus.n23 28.4823
R1978 plus.n17 plus.n6 28.4823
R1979 plus.n58 plus.n57 28.4823
R1980 plus.n51 plus.n40 28.4823
R1981 plus.n19 plus.n18 24.1005
R1982 plus.n19 plus.n4 24.1005
R1983 plus.n53 plus.n38 24.1005
R1984 plus.n53 plus.n52 24.1005
R1985 plus.n23 plus.n4 19.7187
R1986 plus.n18 plus.n17 19.7187
R1987 plus.n57 plus.n38 19.7187
R1988 plus.n52 plus.n51 19.7187
R1989 plus plus.n33 17.2353
R1990 plus.n9 plus.n8 15.6319
R1991 plus.n43 plus.n42 15.6319
R1992 plus.n25 plus.n24 15.3369
R1993 plus.n13 plus.n6 15.3369
R1994 plus.n59 plus.n58 15.3369
R1995 plus.n47 plus.n40 15.3369
R1996 plus.n29 plus.n2 10.955
R1997 plus.n12 plus.n11 10.955
R1998 plus.n63 plus.n36 10.955
R1999 plus.n46 plus.n45 10.955
R2000 plus.n31 plus.n30 6.57323
R2001 plus.n65 plus.n64 6.57323
R2002 plus.n10 plus.n7 0.189894
R2003 plus.n14 plus.n7 0.189894
R2004 plus.n15 plus.n14 0.189894
R2005 plus.n16 plus.n15 0.189894
R2006 plus.n16 plus.n5 0.189894
R2007 plus.n20 plus.n5 0.189894
R2008 plus.n21 plus.n20 0.189894
R2009 plus.n22 plus.n21 0.189894
R2010 plus.n22 plus.n3 0.189894
R2011 plus.n26 plus.n3 0.189894
R2012 plus.n27 plus.n26 0.189894
R2013 plus.n28 plus.n27 0.189894
R2014 plus.n28 plus.n1 0.189894
R2015 plus.n1 plus.n0 0.189894
R2016 plus.n33 plus.n0 0.189894
R2017 plus.n67 plus.n34 0.189894
R2018 plus.n35 plus.n34 0.189894
R2019 plus.n62 plus.n35 0.189894
R2020 plus.n62 plus.n61 0.189894
R2021 plus.n61 plus.n60 0.189894
R2022 plus.n60 plus.n37 0.189894
R2023 plus.n56 plus.n37 0.189894
R2024 plus.n56 plus.n55 0.189894
R2025 plus.n55 plus.n54 0.189894
R2026 plus.n54 plus.n39 0.189894
R2027 plus.n50 plus.n39 0.189894
R2028 plus.n50 plus.n49 0.189894
R2029 plus.n49 plus.n48 0.189894
R2030 plus.n48 plus.n41 0.189894
R2031 plus.n44 plus.n41 0.189894
R2032 drain_left.n6 drain_left.n4 59.6034
R2033 drain_left.n2 drain_left.n0 59.6034
R2034 drain_left.n10 drain_left.n8 59.6034
R2035 drain_left.n7 drain_left.n3 58.7154
R2036 drain_left.n6 drain_left.n5 58.7154
R2037 drain_left.n2 drain_left.n1 58.7154
R2038 drain_left.n14 drain_left.n13 58.7154
R2039 drain_left.n12 drain_left.n11 58.7154
R2040 drain_left.n10 drain_left.n9 58.7154
R2041 drain_left.n16 drain_left.n15 58.7153
R2042 drain_left drain_left.n7 44.319
R2043 drain_left drain_left.n16 6.54115
R2044 drain_left.n12 drain_left.n10 0.888431
R2045 drain_left.n14 drain_left.n12 0.888431
R2046 drain_left.n16 drain_left.n14 0.888431
R2047 drain_left.n7 drain_left.n6 0.833085
R2048 drain_left.n7 drain_left.n2 0.833085
R2049 drain_left.n3 drain_left.t15 0.7925
R2050 drain_left.n3 drain_left.t8 0.7925
R2051 drain_left.n4 drain_left.t19 0.7925
R2052 drain_left.n4 drain_left.t0 0.7925
R2053 drain_left.n5 drain_left.t10 0.7925
R2054 drain_left.n5 drain_left.t3 0.7925
R2055 drain_left.n1 drain_left.t2 0.7925
R2056 drain_left.n1 drain_left.t12 0.7925
R2057 drain_left.n0 drain_left.t4 0.7925
R2058 drain_left.n0 drain_left.t5 0.7925
R2059 drain_left.n15 drain_left.t1 0.7925
R2060 drain_left.n15 drain_left.t16 0.7925
R2061 drain_left.n13 drain_left.t18 0.7925
R2062 drain_left.n13 drain_left.t11 0.7925
R2063 drain_left.n11 drain_left.t14 0.7925
R2064 drain_left.n11 drain_left.t7 0.7925
R2065 drain_left.n9 drain_left.t17 0.7925
R2066 drain_left.n9 drain_left.t9 0.7925
R2067 drain_left.n8 drain_left.t13 0.7925
R2068 drain_left.n8 drain_left.t6 0.7925
C0 drain_right source 45.6943f
C1 drain_left drain_right 1.59885f
C2 minus plus 9.272941f
C3 plus source 25.150698f
C4 drain_left plus 25.7833f
C5 plus drain_right 0.454687f
C6 minus source 25.136599f
C7 drain_left minus 0.173554f
C8 drain_left source 45.6919f
C9 minus drain_right 25.4858f
C10 drain_right a_n2982_n5888# 9.66624f
C11 drain_left a_n2982_n5888# 10.08054f
C12 source a_n2982_n5888# 16.690647f
C13 minus a_n2982_n5888# 12.877324f
C14 plus a_n2982_n5888# 15.325709f
C15 drain_left.t4 a_n2982_n5888# 0.539306f
C16 drain_left.t5 a_n2982_n5888# 0.539306f
C17 drain_left.n0 a_n2982_n5888# 4.97621f
C18 drain_left.t2 a_n2982_n5888# 0.539306f
C19 drain_left.t12 a_n2982_n5888# 0.539306f
C20 drain_left.n1 a_n2982_n5888# 4.97029f
C21 drain_left.n2 a_n2982_n5888# 0.774883f
C22 drain_left.t15 a_n2982_n5888# 0.539306f
C23 drain_left.t8 a_n2982_n5888# 0.539306f
C24 drain_left.n3 a_n2982_n5888# 4.97029f
C25 drain_left.t19 a_n2982_n5888# 0.539306f
C26 drain_left.t0 a_n2982_n5888# 0.539306f
C27 drain_left.n4 a_n2982_n5888# 4.97621f
C28 drain_left.t10 a_n2982_n5888# 0.539306f
C29 drain_left.t3 a_n2982_n5888# 0.539306f
C30 drain_left.n5 a_n2982_n5888# 4.97029f
C31 drain_left.n6 a_n2982_n5888# 0.774883f
C32 drain_left.n7 a_n2982_n5888# 2.888f
C33 drain_left.t13 a_n2982_n5888# 0.539306f
C34 drain_left.t6 a_n2982_n5888# 0.539306f
C35 drain_left.n8 a_n2982_n5888# 4.97622f
C36 drain_left.t17 a_n2982_n5888# 0.539306f
C37 drain_left.t9 a_n2982_n5888# 0.539306f
C38 drain_left.n9 a_n2982_n5888# 4.97029f
C39 drain_left.n10 a_n2982_n5888# 0.778988f
C40 drain_left.t14 a_n2982_n5888# 0.539306f
C41 drain_left.t7 a_n2982_n5888# 0.539306f
C42 drain_left.n11 a_n2982_n5888# 4.97029f
C43 drain_left.n12 a_n2982_n5888# 0.386961f
C44 drain_left.t18 a_n2982_n5888# 0.539306f
C45 drain_left.t11 a_n2982_n5888# 0.539306f
C46 drain_left.n13 a_n2982_n5888# 4.97029f
C47 drain_left.n14 a_n2982_n5888# 0.386961f
C48 drain_left.t1 a_n2982_n5888# 0.539306f
C49 drain_left.t16 a_n2982_n5888# 0.539306f
C50 drain_left.n15 a_n2982_n5888# 4.97027f
C51 drain_left.n16 a_n2982_n5888# 0.628431f
C52 plus.n0 a_n2982_n5888# 0.039641f
C53 plus.t3 a_n2982_n5888# 1.96047f
C54 plus.t18 a_n2982_n5888# 1.96047f
C55 plus.n1 a_n2982_n5888# 0.039641f
C56 plus.t8 a_n2982_n5888# 1.96047f
C57 plus.n2 a_n2982_n5888# 0.715669f
C58 plus.n3 a_n2982_n5888# 0.039641f
C59 plus.t1 a_n2982_n5888# 1.96047f
C60 plus.t12 a_n2982_n5888# 1.96047f
C61 plus.n4 a_n2982_n5888# 0.715669f
C62 plus.n5 a_n2982_n5888# 0.039641f
C63 plus.t5 a_n2982_n5888# 1.96047f
C64 plus.t10 a_n2982_n5888# 1.96047f
C65 plus.n6 a_n2982_n5888# 0.715669f
C66 plus.n7 a_n2982_n5888# 0.039641f
C67 plus.t2 a_n2982_n5888# 1.96047f
C68 plus.t13 a_n2982_n5888# 1.96047f
C69 plus.n8 a_n2982_n5888# 0.722299f
C70 plus.t6 a_n2982_n5888# 1.97977f
C71 plus.n9 a_n2982_n5888# 0.699216f
C72 plus.n10 a_n2982_n5888# 0.169205f
C73 plus.n11 a_n2982_n5888# 0.008995f
C74 plus.n12 a_n2982_n5888# 0.715669f
C75 plus.n13 a_n2982_n5888# 0.008995f
C76 plus.n14 a_n2982_n5888# 0.039641f
C77 plus.n15 a_n2982_n5888# 0.039641f
C78 plus.n16 a_n2982_n5888# 0.039641f
C79 plus.n17 a_n2982_n5888# 0.008995f
C80 plus.n18 a_n2982_n5888# 0.715669f
C81 plus.n19 a_n2982_n5888# 0.008995f
C82 plus.n20 a_n2982_n5888# 0.039641f
C83 plus.n21 a_n2982_n5888# 0.039641f
C84 plus.n22 a_n2982_n5888# 0.039641f
C85 plus.n23 a_n2982_n5888# 0.008995f
C86 plus.n24 a_n2982_n5888# 0.715669f
C87 plus.n25 a_n2982_n5888# 0.008995f
C88 plus.n26 a_n2982_n5888# 0.039641f
C89 plus.n27 a_n2982_n5888# 0.039641f
C90 plus.n28 a_n2982_n5888# 0.039641f
C91 plus.n29 a_n2982_n5888# 0.008995f
C92 plus.n30 a_n2982_n5888# 0.715669f
C93 plus.n31 a_n2982_n5888# 0.008995f
C94 plus.n32 a_n2982_n5888# 0.715302f
C95 plus.n33 a_n2982_n5888# 0.722491f
C96 plus.n34 a_n2982_n5888# 0.039641f
C97 plus.t15 a_n2982_n5888# 1.96047f
C98 plus.n35 a_n2982_n5888# 0.039641f
C99 plus.t14 a_n2982_n5888# 1.96047f
C100 plus.t17 a_n2982_n5888# 1.96047f
C101 plus.n36 a_n2982_n5888# 0.715669f
C102 plus.n37 a_n2982_n5888# 0.039641f
C103 plus.t7 a_n2982_n5888# 1.96047f
C104 plus.t4 a_n2982_n5888# 1.96047f
C105 plus.n38 a_n2982_n5888# 0.715669f
C106 plus.n39 a_n2982_n5888# 0.039641f
C107 plus.t11 a_n2982_n5888# 1.96047f
C108 plus.t9 a_n2982_n5888# 1.96047f
C109 plus.n40 a_n2982_n5888# 0.715669f
C110 plus.n41 a_n2982_n5888# 0.039641f
C111 plus.t16 a_n2982_n5888# 1.96047f
C112 plus.t0 a_n2982_n5888# 1.96047f
C113 plus.n42 a_n2982_n5888# 0.722299f
C114 plus.t19 a_n2982_n5888# 1.97977f
C115 plus.n43 a_n2982_n5888# 0.699216f
C116 plus.n44 a_n2982_n5888# 0.169205f
C117 plus.n45 a_n2982_n5888# 0.008995f
C118 plus.n46 a_n2982_n5888# 0.715669f
C119 plus.n47 a_n2982_n5888# 0.008995f
C120 plus.n48 a_n2982_n5888# 0.039641f
C121 plus.n49 a_n2982_n5888# 0.039641f
C122 plus.n50 a_n2982_n5888# 0.039641f
C123 plus.n51 a_n2982_n5888# 0.008995f
C124 plus.n52 a_n2982_n5888# 0.715669f
C125 plus.n53 a_n2982_n5888# 0.008995f
C126 plus.n54 a_n2982_n5888# 0.039641f
C127 plus.n55 a_n2982_n5888# 0.039641f
C128 plus.n56 a_n2982_n5888# 0.039641f
C129 plus.n57 a_n2982_n5888# 0.008995f
C130 plus.n58 a_n2982_n5888# 0.715669f
C131 plus.n59 a_n2982_n5888# 0.008995f
C132 plus.n60 a_n2982_n5888# 0.039641f
C133 plus.n61 a_n2982_n5888# 0.039641f
C134 plus.n62 a_n2982_n5888# 0.039641f
C135 plus.n63 a_n2982_n5888# 0.008995f
C136 plus.n64 a_n2982_n5888# 0.715669f
C137 plus.n65 a_n2982_n5888# 0.008995f
C138 plus.n66 a_n2982_n5888# 0.715302f
C139 plus.n67 a_n2982_n5888# 1.78318f
C140 source.n0 a_n2982_n5888# 0.031979f
C141 source.n1 a_n2982_n5888# 0.023196f
C142 source.n2 a_n2982_n5888# 0.012465f
C143 source.n3 a_n2982_n5888# 0.029462f
C144 source.n4 a_n2982_n5888# 0.013198f
C145 source.n5 a_n2982_n5888# 0.023196f
C146 source.n6 a_n2982_n5888# 0.012465f
C147 source.n7 a_n2982_n5888# 0.029462f
C148 source.n8 a_n2982_n5888# 0.013198f
C149 source.n9 a_n2982_n5888# 0.023196f
C150 source.n10 a_n2982_n5888# 0.012465f
C151 source.n11 a_n2982_n5888# 0.029462f
C152 source.n12 a_n2982_n5888# 0.013198f
C153 source.n13 a_n2982_n5888# 0.023196f
C154 source.n14 a_n2982_n5888# 0.012465f
C155 source.n15 a_n2982_n5888# 0.029462f
C156 source.n16 a_n2982_n5888# 0.029462f
C157 source.n17 a_n2982_n5888# 0.013198f
C158 source.n18 a_n2982_n5888# 0.023196f
C159 source.n19 a_n2982_n5888# 0.012465f
C160 source.n20 a_n2982_n5888# 0.029462f
C161 source.n21 a_n2982_n5888# 0.013198f
C162 source.n22 a_n2982_n5888# 0.023196f
C163 source.n23 a_n2982_n5888# 0.012465f
C164 source.n24 a_n2982_n5888# 0.029462f
C165 source.n25 a_n2982_n5888# 0.013198f
C166 source.n26 a_n2982_n5888# 0.023196f
C167 source.n27 a_n2982_n5888# 0.012465f
C168 source.n28 a_n2982_n5888# 0.029462f
C169 source.n29 a_n2982_n5888# 0.013198f
C170 source.n30 a_n2982_n5888# 0.023196f
C171 source.n31 a_n2982_n5888# 0.012465f
C172 source.n32 a_n2982_n5888# 0.029462f
C173 source.n33 a_n2982_n5888# 0.013198f
C174 source.n34 a_n2982_n5888# 0.023196f
C175 source.n35 a_n2982_n5888# 0.012831f
C176 source.n36 a_n2982_n5888# 0.029462f
C177 source.n37 a_n2982_n5888# 0.012465f
C178 source.n38 a_n2982_n5888# 0.013198f
C179 source.n39 a_n2982_n5888# 0.023196f
C180 source.n40 a_n2982_n5888# 0.012465f
C181 source.n41 a_n2982_n5888# 0.029462f
C182 source.n42 a_n2982_n5888# 0.013198f
C183 source.n43 a_n2982_n5888# 0.023196f
C184 source.n44 a_n2982_n5888# 0.012465f
C185 source.n45 a_n2982_n5888# 0.022097f
C186 source.n46 a_n2982_n5888# 0.020828f
C187 source.t16 a_n2982_n5888# 0.051384f
C188 source.n47 a_n2982_n5888# 0.283016f
C189 source.n48 a_n2982_n5888# 2.51149f
C190 source.n49 a_n2982_n5888# 0.012465f
C191 source.n50 a_n2982_n5888# 0.013198f
C192 source.n51 a_n2982_n5888# 0.029462f
C193 source.n52 a_n2982_n5888# 0.029462f
C194 source.n53 a_n2982_n5888# 0.013198f
C195 source.n54 a_n2982_n5888# 0.012465f
C196 source.n55 a_n2982_n5888# 0.023196f
C197 source.n56 a_n2982_n5888# 0.023196f
C198 source.n57 a_n2982_n5888# 0.012465f
C199 source.n58 a_n2982_n5888# 0.013198f
C200 source.n59 a_n2982_n5888# 0.029462f
C201 source.n60 a_n2982_n5888# 0.029462f
C202 source.n61 a_n2982_n5888# 0.013198f
C203 source.n62 a_n2982_n5888# 0.012465f
C204 source.n63 a_n2982_n5888# 0.023196f
C205 source.n64 a_n2982_n5888# 0.023196f
C206 source.n65 a_n2982_n5888# 0.012465f
C207 source.n66 a_n2982_n5888# 0.013198f
C208 source.n67 a_n2982_n5888# 0.029462f
C209 source.n68 a_n2982_n5888# 0.029462f
C210 source.n69 a_n2982_n5888# 0.029462f
C211 source.n70 a_n2982_n5888# 0.012831f
C212 source.n71 a_n2982_n5888# 0.012465f
C213 source.n72 a_n2982_n5888# 0.023196f
C214 source.n73 a_n2982_n5888# 0.023196f
C215 source.n74 a_n2982_n5888# 0.012465f
C216 source.n75 a_n2982_n5888# 0.013198f
C217 source.n76 a_n2982_n5888# 0.029462f
C218 source.n77 a_n2982_n5888# 0.029462f
C219 source.n78 a_n2982_n5888# 0.013198f
C220 source.n79 a_n2982_n5888# 0.012465f
C221 source.n80 a_n2982_n5888# 0.023196f
C222 source.n81 a_n2982_n5888# 0.023196f
C223 source.n82 a_n2982_n5888# 0.012465f
C224 source.n83 a_n2982_n5888# 0.013198f
C225 source.n84 a_n2982_n5888# 0.029462f
C226 source.n85 a_n2982_n5888# 0.029462f
C227 source.n86 a_n2982_n5888# 0.013198f
C228 source.n87 a_n2982_n5888# 0.012465f
C229 source.n88 a_n2982_n5888# 0.023196f
C230 source.n89 a_n2982_n5888# 0.023196f
C231 source.n90 a_n2982_n5888# 0.012465f
C232 source.n91 a_n2982_n5888# 0.013198f
C233 source.n92 a_n2982_n5888# 0.029462f
C234 source.n93 a_n2982_n5888# 0.029462f
C235 source.n94 a_n2982_n5888# 0.013198f
C236 source.n95 a_n2982_n5888# 0.012465f
C237 source.n96 a_n2982_n5888# 0.023196f
C238 source.n97 a_n2982_n5888# 0.023196f
C239 source.n98 a_n2982_n5888# 0.012465f
C240 source.n99 a_n2982_n5888# 0.013198f
C241 source.n100 a_n2982_n5888# 0.029462f
C242 source.n101 a_n2982_n5888# 0.029462f
C243 source.n102 a_n2982_n5888# 0.013198f
C244 source.n103 a_n2982_n5888# 0.012465f
C245 source.n104 a_n2982_n5888# 0.023196f
C246 source.n105 a_n2982_n5888# 0.023196f
C247 source.n106 a_n2982_n5888# 0.012465f
C248 source.n107 a_n2982_n5888# 0.013198f
C249 source.n108 a_n2982_n5888# 0.029462f
C250 source.n109 a_n2982_n5888# 0.029462f
C251 source.n110 a_n2982_n5888# 0.013198f
C252 source.n111 a_n2982_n5888# 0.012465f
C253 source.n112 a_n2982_n5888# 0.023196f
C254 source.n113 a_n2982_n5888# 0.023196f
C255 source.n114 a_n2982_n5888# 0.012465f
C256 source.n115 a_n2982_n5888# 0.012831f
C257 source.n116 a_n2982_n5888# 0.012831f
C258 source.n117 a_n2982_n5888# 0.029462f
C259 source.n118 a_n2982_n5888# 0.029462f
C260 source.n119 a_n2982_n5888# 0.013198f
C261 source.n120 a_n2982_n5888# 0.012465f
C262 source.n121 a_n2982_n5888# 0.023196f
C263 source.n122 a_n2982_n5888# 0.023196f
C264 source.n123 a_n2982_n5888# 0.012465f
C265 source.n124 a_n2982_n5888# 0.013198f
C266 source.n125 a_n2982_n5888# 0.029462f
C267 source.n126 a_n2982_n5888# 0.029462f
C268 source.n127 a_n2982_n5888# 0.013198f
C269 source.n128 a_n2982_n5888# 0.012465f
C270 source.n129 a_n2982_n5888# 0.023196f
C271 source.n130 a_n2982_n5888# 0.023196f
C272 source.n131 a_n2982_n5888# 0.012465f
C273 source.n132 a_n2982_n5888# 0.013198f
C274 source.n133 a_n2982_n5888# 0.029462f
C275 source.n134 a_n2982_n5888# 0.062674f
C276 source.n135 a_n2982_n5888# 0.013198f
C277 source.n136 a_n2982_n5888# 0.012465f
C278 source.n137 a_n2982_n5888# 0.051082f
C279 source.n138 a_n2982_n5888# 0.034875f
C280 source.n139 a_n2982_n5888# 1.86296f
C281 source.t4 a_n2982_n5888# 0.458263f
C282 source.t11 a_n2982_n5888# 0.458263f
C283 source.n140 a_n2982_n5888# 4.14734f
C284 source.n141 a_n2982_n5888# 0.373328f
C285 source.t6 a_n2982_n5888# 0.458263f
C286 source.t17 a_n2982_n5888# 0.458263f
C287 source.n142 a_n2982_n5888# 4.14734f
C288 source.n143 a_n2982_n5888# 0.373328f
C289 source.t12 a_n2982_n5888# 0.458263f
C290 source.t18 a_n2982_n5888# 0.458263f
C291 source.n144 a_n2982_n5888# 4.14734f
C292 source.n145 a_n2982_n5888# 0.373328f
C293 source.t13 a_n2982_n5888# 0.458263f
C294 source.t0 a_n2982_n5888# 0.458263f
C295 source.n146 a_n2982_n5888# 4.14734f
C296 source.n147 a_n2982_n5888# 0.373328f
C297 source.n148 a_n2982_n5888# 0.031979f
C298 source.n149 a_n2982_n5888# 0.023196f
C299 source.n150 a_n2982_n5888# 0.012465f
C300 source.n151 a_n2982_n5888# 0.029462f
C301 source.n152 a_n2982_n5888# 0.013198f
C302 source.n153 a_n2982_n5888# 0.023196f
C303 source.n154 a_n2982_n5888# 0.012465f
C304 source.n155 a_n2982_n5888# 0.029462f
C305 source.n156 a_n2982_n5888# 0.013198f
C306 source.n157 a_n2982_n5888# 0.023196f
C307 source.n158 a_n2982_n5888# 0.012465f
C308 source.n159 a_n2982_n5888# 0.029462f
C309 source.n160 a_n2982_n5888# 0.013198f
C310 source.n161 a_n2982_n5888# 0.023196f
C311 source.n162 a_n2982_n5888# 0.012465f
C312 source.n163 a_n2982_n5888# 0.029462f
C313 source.n164 a_n2982_n5888# 0.029462f
C314 source.n165 a_n2982_n5888# 0.013198f
C315 source.n166 a_n2982_n5888# 0.023196f
C316 source.n167 a_n2982_n5888# 0.012465f
C317 source.n168 a_n2982_n5888# 0.029462f
C318 source.n169 a_n2982_n5888# 0.013198f
C319 source.n170 a_n2982_n5888# 0.023196f
C320 source.n171 a_n2982_n5888# 0.012465f
C321 source.n172 a_n2982_n5888# 0.029462f
C322 source.n173 a_n2982_n5888# 0.013198f
C323 source.n174 a_n2982_n5888# 0.023196f
C324 source.n175 a_n2982_n5888# 0.012465f
C325 source.n176 a_n2982_n5888# 0.029462f
C326 source.n177 a_n2982_n5888# 0.013198f
C327 source.n178 a_n2982_n5888# 0.023196f
C328 source.n179 a_n2982_n5888# 0.012465f
C329 source.n180 a_n2982_n5888# 0.029462f
C330 source.n181 a_n2982_n5888# 0.013198f
C331 source.n182 a_n2982_n5888# 0.023196f
C332 source.n183 a_n2982_n5888# 0.012831f
C333 source.n184 a_n2982_n5888# 0.029462f
C334 source.n185 a_n2982_n5888# 0.012465f
C335 source.n186 a_n2982_n5888# 0.013198f
C336 source.n187 a_n2982_n5888# 0.023196f
C337 source.n188 a_n2982_n5888# 0.012465f
C338 source.n189 a_n2982_n5888# 0.029462f
C339 source.n190 a_n2982_n5888# 0.013198f
C340 source.n191 a_n2982_n5888# 0.023196f
C341 source.n192 a_n2982_n5888# 0.012465f
C342 source.n193 a_n2982_n5888# 0.022097f
C343 source.n194 a_n2982_n5888# 0.020828f
C344 source.t5 a_n2982_n5888# 0.051384f
C345 source.n195 a_n2982_n5888# 0.283016f
C346 source.n196 a_n2982_n5888# 2.51149f
C347 source.n197 a_n2982_n5888# 0.012465f
C348 source.n198 a_n2982_n5888# 0.013198f
C349 source.n199 a_n2982_n5888# 0.029462f
C350 source.n200 a_n2982_n5888# 0.029462f
C351 source.n201 a_n2982_n5888# 0.013198f
C352 source.n202 a_n2982_n5888# 0.012465f
C353 source.n203 a_n2982_n5888# 0.023196f
C354 source.n204 a_n2982_n5888# 0.023196f
C355 source.n205 a_n2982_n5888# 0.012465f
C356 source.n206 a_n2982_n5888# 0.013198f
C357 source.n207 a_n2982_n5888# 0.029462f
C358 source.n208 a_n2982_n5888# 0.029462f
C359 source.n209 a_n2982_n5888# 0.013198f
C360 source.n210 a_n2982_n5888# 0.012465f
C361 source.n211 a_n2982_n5888# 0.023196f
C362 source.n212 a_n2982_n5888# 0.023196f
C363 source.n213 a_n2982_n5888# 0.012465f
C364 source.n214 a_n2982_n5888# 0.013198f
C365 source.n215 a_n2982_n5888# 0.029462f
C366 source.n216 a_n2982_n5888# 0.029462f
C367 source.n217 a_n2982_n5888# 0.029462f
C368 source.n218 a_n2982_n5888# 0.012831f
C369 source.n219 a_n2982_n5888# 0.012465f
C370 source.n220 a_n2982_n5888# 0.023196f
C371 source.n221 a_n2982_n5888# 0.023196f
C372 source.n222 a_n2982_n5888# 0.012465f
C373 source.n223 a_n2982_n5888# 0.013198f
C374 source.n224 a_n2982_n5888# 0.029462f
C375 source.n225 a_n2982_n5888# 0.029462f
C376 source.n226 a_n2982_n5888# 0.013198f
C377 source.n227 a_n2982_n5888# 0.012465f
C378 source.n228 a_n2982_n5888# 0.023196f
C379 source.n229 a_n2982_n5888# 0.023196f
C380 source.n230 a_n2982_n5888# 0.012465f
C381 source.n231 a_n2982_n5888# 0.013198f
C382 source.n232 a_n2982_n5888# 0.029462f
C383 source.n233 a_n2982_n5888# 0.029462f
C384 source.n234 a_n2982_n5888# 0.013198f
C385 source.n235 a_n2982_n5888# 0.012465f
C386 source.n236 a_n2982_n5888# 0.023196f
C387 source.n237 a_n2982_n5888# 0.023196f
C388 source.n238 a_n2982_n5888# 0.012465f
C389 source.n239 a_n2982_n5888# 0.013198f
C390 source.n240 a_n2982_n5888# 0.029462f
C391 source.n241 a_n2982_n5888# 0.029462f
C392 source.n242 a_n2982_n5888# 0.013198f
C393 source.n243 a_n2982_n5888# 0.012465f
C394 source.n244 a_n2982_n5888# 0.023196f
C395 source.n245 a_n2982_n5888# 0.023196f
C396 source.n246 a_n2982_n5888# 0.012465f
C397 source.n247 a_n2982_n5888# 0.013198f
C398 source.n248 a_n2982_n5888# 0.029462f
C399 source.n249 a_n2982_n5888# 0.029462f
C400 source.n250 a_n2982_n5888# 0.013198f
C401 source.n251 a_n2982_n5888# 0.012465f
C402 source.n252 a_n2982_n5888# 0.023196f
C403 source.n253 a_n2982_n5888# 0.023196f
C404 source.n254 a_n2982_n5888# 0.012465f
C405 source.n255 a_n2982_n5888# 0.013198f
C406 source.n256 a_n2982_n5888# 0.029462f
C407 source.n257 a_n2982_n5888# 0.029462f
C408 source.n258 a_n2982_n5888# 0.013198f
C409 source.n259 a_n2982_n5888# 0.012465f
C410 source.n260 a_n2982_n5888# 0.023196f
C411 source.n261 a_n2982_n5888# 0.023196f
C412 source.n262 a_n2982_n5888# 0.012465f
C413 source.n263 a_n2982_n5888# 0.012831f
C414 source.n264 a_n2982_n5888# 0.012831f
C415 source.n265 a_n2982_n5888# 0.029462f
C416 source.n266 a_n2982_n5888# 0.029462f
C417 source.n267 a_n2982_n5888# 0.013198f
C418 source.n268 a_n2982_n5888# 0.012465f
C419 source.n269 a_n2982_n5888# 0.023196f
C420 source.n270 a_n2982_n5888# 0.023196f
C421 source.n271 a_n2982_n5888# 0.012465f
C422 source.n272 a_n2982_n5888# 0.013198f
C423 source.n273 a_n2982_n5888# 0.029462f
C424 source.n274 a_n2982_n5888# 0.029462f
C425 source.n275 a_n2982_n5888# 0.013198f
C426 source.n276 a_n2982_n5888# 0.012465f
C427 source.n277 a_n2982_n5888# 0.023196f
C428 source.n278 a_n2982_n5888# 0.023196f
C429 source.n279 a_n2982_n5888# 0.012465f
C430 source.n280 a_n2982_n5888# 0.013198f
C431 source.n281 a_n2982_n5888# 0.029462f
C432 source.n282 a_n2982_n5888# 0.062674f
C433 source.n283 a_n2982_n5888# 0.013198f
C434 source.n284 a_n2982_n5888# 0.012465f
C435 source.n285 a_n2982_n5888# 0.051082f
C436 source.n286 a_n2982_n5888# 0.034875f
C437 source.n287 a_n2982_n5888# 0.119867f
C438 source.n288 a_n2982_n5888# 0.031979f
C439 source.n289 a_n2982_n5888# 0.023196f
C440 source.n290 a_n2982_n5888# 0.012465f
C441 source.n291 a_n2982_n5888# 0.029462f
C442 source.n292 a_n2982_n5888# 0.013198f
C443 source.n293 a_n2982_n5888# 0.023196f
C444 source.n294 a_n2982_n5888# 0.012465f
C445 source.n295 a_n2982_n5888# 0.029462f
C446 source.n296 a_n2982_n5888# 0.013198f
C447 source.n297 a_n2982_n5888# 0.023196f
C448 source.n298 a_n2982_n5888# 0.012465f
C449 source.n299 a_n2982_n5888# 0.029462f
C450 source.n300 a_n2982_n5888# 0.013198f
C451 source.n301 a_n2982_n5888# 0.023196f
C452 source.n302 a_n2982_n5888# 0.012465f
C453 source.n303 a_n2982_n5888# 0.029462f
C454 source.n304 a_n2982_n5888# 0.029462f
C455 source.n305 a_n2982_n5888# 0.013198f
C456 source.n306 a_n2982_n5888# 0.023196f
C457 source.n307 a_n2982_n5888# 0.012465f
C458 source.n308 a_n2982_n5888# 0.029462f
C459 source.n309 a_n2982_n5888# 0.013198f
C460 source.n310 a_n2982_n5888# 0.023196f
C461 source.n311 a_n2982_n5888# 0.012465f
C462 source.n312 a_n2982_n5888# 0.029462f
C463 source.n313 a_n2982_n5888# 0.013198f
C464 source.n314 a_n2982_n5888# 0.023196f
C465 source.n315 a_n2982_n5888# 0.012465f
C466 source.n316 a_n2982_n5888# 0.029462f
C467 source.n317 a_n2982_n5888# 0.013198f
C468 source.n318 a_n2982_n5888# 0.023196f
C469 source.n319 a_n2982_n5888# 0.012465f
C470 source.n320 a_n2982_n5888# 0.029462f
C471 source.n321 a_n2982_n5888# 0.013198f
C472 source.n322 a_n2982_n5888# 0.023196f
C473 source.n323 a_n2982_n5888# 0.012831f
C474 source.n324 a_n2982_n5888# 0.029462f
C475 source.n325 a_n2982_n5888# 0.012465f
C476 source.n326 a_n2982_n5888# 0.013198f
C477 source.n327 a_n2982_n5888# 0.023196f
C478 source.n328 a_n2982_n5888# 0.012465f
C479 source.n329 a_n2982_n5888# 0.029462f
C480 source.n330 a_n2982_n5888# 0.013198f
C481 source.n331 a_n2982_n5888# 0.023196f
C482 source.n332 a_n2982_n5888# 0.012465f
C483 source.n333 a_n2982_n5888# 0.022097f
C484 source.n334 a_n2982_n5888# 0.020828f
C485 source.t27 a_n2982_n5888# 0.051384f
C486 source.n335 a_n2982_n5888# 0.283016f
C487 source.n336 a_n2982_n5888# 2.51149f
C488 source.n337 a_n2982_n5888# 0.012465f
C489 source.n338 a_n2982_n5888# 0.013198f
C490 source.n339 a_n2982_n5888# 0.029462f
C491 source.n340 a_n2982_n5888# 0.029462f
C492 source.n341 a_n2982_n5888# 0.013198f
C493 source.n342 a_n2982_n5888# 0.012465f
C494 source.n343 a_n2982_n5888# 0.023196f
C495 source.n344 a_n2982_n5888# 0.023196f
C496 source.n345 a_n2982_n5888# 0.012465f
C497 source.n346 a_n2982_n5888# 0.013198f
C498 source.n347 a_n2982_n5888# 0.029462f
C499 source.n348 a_n2982_n5888# 0.029462f
C500 source.n349 a_n2982_n5888# 0.013198f
C501 source.n350 a_n2982_n5888# 0.012465f
C502 source.n351 a_n2982_n5888# 0.023196f
C503 source.n352 a_n2982_n5888# 0.023196f
C504 source.n353 a_n2982_n5888# 0.012465f
C505 source.n354 a_n2982_n5888# 0.013198f
C506 source.n355 a_n2982_n5888# 0.029462f
C507 source.n356 a_n2982_n5888# 0.029462f
C508 source.n357 a_n2982_n5888# 0.029462f
C509 source.n358 a_n2982_n5888# 0.012831f
C510 source.n359 a_n2982_n5888# 0.012465f
C511 source.n360 a_n2982_n5888# 0.023196f
C512 source.n361 a_n2982_n5888# 0.023196f
C513 source.n362 a_n2982_n5888# 0.012465f
C514 source.n363 a_n2982_n5888# 0.013198f
C515 source.n364 a_n2982_n5888# 0.029462f
C516 source.n365 a_n2982_n5888# 0.029462f
C517 source.n366 a_n2982_n5888# 0.013198f
C518 source.n367 a_n2982_n5888# 0.012465f
C519 source.n368 a_n2982_n5888# 0.023196f
C520 source.n369 a_n2982_n5888# 0.023196f
C521 source.n370 a_n2982_n5888# 0.012465f
C522 source.n371 a_n2982_n5888# 0.013198f
C523 source.n372 a_n2982_n5888# 0.029462f
C524 source.n373 a_n2982_n5888# 0.029462f
C525 source.n374 a_n2982_n5888# 0.013198f
C526 source.n375 a_n2982_n5888# 0.012465f
C527 source.n376 a_n2982_n5888# 0.023196f
C528 source.n377 a_n2982_n5888# 0.023196f
C529 source.n378 a_n2982_n5888# 0.012465f
C530 source.n379 a_n2982_n5888# 0.013198f
C531 source.n380 a_n2982_n5888# 0.029462f
C532 source.n381 a_n2982_n5888# 0.029462f
C533 source.n382 a_n2982_n5888# 0.013198f
C534 source.n383 a_n2982_n5888# 0.012465f
C535 source.n384 a_n2982_n5888# 0.023196f
C536 source.n385 a_n2982_n5888# 0.023196f
C537 source.n386 a_n2982_n5888# 0.012465f
C538 source.n387 a_n2982_n5888# 0.013198f
C539 source.n388 a_n2982_n5888# 0.029462f
C540 source.n389 a_n2982_n5888# 0.029462f
C541 source.n390 a_n2982_n5888# 0.013198f
C542 source.n391 a_n2982_n5888# 0.012465f
C543 source.n392 a_n2982_n5888# 0.023196f
C544 source.n393 a_n2982_n5888# 0.023196f
C545 source.n394 a_n2982_n5888# 0.012465f
C546 source.n395 a_n2982_n5888# 0.013198f
C547 source.n396 a_n2982_n5888# 0.029462f
C548 source.n397 a_n2982_n5888# 0.029462f
C549 source.n398 a_n2982_n5888# 0.013198f
C550 source.n399 a_n2982_n5888# 0.012465f
C551 source.n400 a_n2982_n5888# 0.023196f
C552 source.n401 a_n2982_n5888# 0.023196f
C553 source.n402 a_n2982_n5888# 0.012465f
C554 source.n403 a_n2982_n5888# 0.012831f
C555 source.n404 a_n2982_n5888# 0.012831f
C556 source.n405 a_n2982_n5888# 0.029462f
C557 source.n406 a_n2982_n5888# 0.029462f
C558 source.n407 a_n2982_n5888# 0.013198f
C559 source.n408 a_n2982_n5888# 0.012465f
C560 source.n409 a_n2982_n5888# 0.023196f
C561 source.n410 a_n2982_n5888# 0.023196f
C562 source.n411 a_n2982_n5888# 0.012465f
C563 source.n412 a_n2982_n5888# 0.013198f
C564 source.n413 a_n2982_n5888# 0.029462f
C565 source.n414 a_n2982_n5888# 0.029462f
C566 source.n415 a_n2982_n5888# 0.013198f
C567 source.n416 a_n2982_n5888# 0.012465f
C568 source.n417 a_n2982_n5888# 0.023196f
C569 source.n418 a_n2982_n5888# 0.023196f
C570 source.n419 a_n2982_n5888# 0.012465f
C571 source.n420 a_n2982_n5888# 0.013198f
C572 source.n421 a_n2982_n5888# 0.029462f
C573 source.n422 a_n2982_n5888# 0.062674f
C574 source.n423 a_n2982_n5888# 0.013198f
C575 source.n424 a_n2982_n5888# 0.012465f
C576 source.n425 a_n2982_n5888# 0.051082f
C577 source.n426 a_n2982_n5888# 0.034875f
C578 source.n427 a_n2982_n5888# 0.119867f
C579 source.t28 a_n2982_n5888# 0.458263f
C580 source.t36 a_n2982_n5888# 0.458263f
C581 source.n428 a_n2982_n5888# 4.14734f
C582 source.n429 a_n2982_n5888# 0.373328f
C583 source.t29 a_n2982_n5888# 0.458263f
C584 source.t20 a_n2982_n5888# 0.458263f
C585 source.n430 a_n2982_n5888# 4.14734f
C586 source.n431 a_n2982_n5888# 0.373328f
C587 source.t30 a_n2982_n5888# 0.458263f
C588 source.t19 a_n2982_n5888# 0.458263f
C589 source.n432 a_n2982_n5888# 4.14734f
C590 source.n433 a_n2982_n5888# 0.373328f
C591 source.t32 a_n2982_n5888# 0.458263f
C592 source.t23 a_n2982_n5888# 0.458263f
C593 source.n434 a_n2982_n5888# 4.14734f
C594 source.n435 a_n2982_n5888# 0.373328f
C595 source.n436 a_n2982_n5888# 0.031979f
C596 source.n437 a_n2982_n5888# 0.023196f
C597 source.n438 a_n2982_n5888# 0.012465f
C598 source.n439 a_n2982_n5888# 0.029462f
C599 source.n440 a_n2982_n5888# 0.013198f
C600 source.n441 a_n2982_n5888# 0.023196f
C601 source.n442 a_n2982_n5888# 0.012465f
C602 source.n443 a_n2982_n5888# 0.029462f
C603 source.n444 a_n2982_n5888# 0.013198f
C604 source.n445 a_n2982_n5888# 0.023196f
C605 source.n446 a_n2982_n5888# 0.012465f
C606 source.n447 a_n2982_n5888# 0.029462f
C607 source.n448 a_n2982_n5888# 0.013198f
C608 source.n449 a_n2982_n5888# 0.023196f
C609 source.n450 a_n2982_n5888# 0.012465f
C610 source.n451 a_n2982_n5888# 0.029462f
C611 source.n452 a_n2982_n5888# 0.029462f
C612 source.n453 a_n2982_n5888# 0.013198f
C613 source.n454 a_n2982_n5888# 0.023196f
C614 source.n455 a_n2982_n5888# 0.012465f
C615 source.n456 a_n2982_n5888# 0.029462f
C616 source.n457 a_n2982_n5888# 0.013198f
C617 source.n458 a_n2982_n5888# 0.023196f
C618 source.n459 a_n2982_n5888# 0.012465f
C619 source.n460 a_n2982_n5888# 0.029462f
C620 source.n461 a_n2982_n5888# 0.013198f
C621 source.n462 a_n2982_n5888# 0.023196f
C622 source.n463 a_n2982_n5888# 0.012465f
C623 source.n464 a_n2982_n5888# 0.029462f
C624 source.n465 a_n2982_n5888# 0.013198f
C625 source.n466 a_n2982_n5888# 0.023196f
C626 source.n467 a_n2982_n5888# 0.012465f
C627 source.n468 a_n2982_n5888# 0.029462f
C628 source.n469 a_n2982_n5888# 0.013198f
C629 source.n470 a_n2982_n5888# 0.023196f
C630 source.n471 a_n2982_n5888# 0.012831f
C631 source.n472 a_n2982_n5888# 0.029462f
C632 source.n473 a_n2982_n5888# 0.012465f
C633 source.n474 a_n2982_n5888# 0.013198f
C634 source.n475 a_n2982_n5888# 0.023196f
C635 source.n476 a_n2982_n5888# 0.012465f
C636 source.n477 a_n2982_n5888# 0.029462f
C637 source.n478 a_n2982_n5888# 0.013198f
C638 source.n479 a_n2982_n5888# 0.023196f
C639 source.n480 a_n2982_n5888# 0.012465f
C640 source.n481 a_n2982_n5888# 0.022097f
C641 source.n482 a_n2982_n5888# 0.020828f
C642 source.t24 a_n2982_n5888# 0.051384f
C643 source.n483 a_n2982_n5888# 0.283016f
C644 source.n484 a_n2982_n5888# 2.51149f
C645 source.n485 a_n2982_n5888# 0.012465f
C646 source.n486 a_n2982_n5888# 0.013198f
C647 source.n487 a_n2982_n5888# 0.029462f
C648 source.n488 a_n2982_n5888# 0.029462f
C649 source.n489 a_n2982_n5888# 0.013198f
C650 source.n490 a_n2982_n5888# 0.012465f
C651 source.n491 a_n2982_n5888# 0.023196f
C652 source.n492 a_n2982_n5888# 0.023196f
C653 source.n493 a_n2982_n5888# 0.012465f
C654 source.n494 a_n2982_n5888# 0.013198f
C655 source.n495 a_n2982_n5888# 0.029462f
C656 source.n496 a_n2982_n5888# 0.029462f
C657 source.n497 a_n2982_n5888# 0.013198f
C658 source.n498 a_n2982_n5888# 0.012465f
C659 source.n499 a_n2982_n5888# 0.023196f
C660 source.n500 a_n2982_n5888# 0.023196f
C661 source.n501 a_n2982_n5888# 0.012465f
C662 source.n502 a_n2982_n5888# 0.013198f
C663 source.n503 a_n2982_n5888# 0.029462f
C664 source.n504 a_n2982_n5888# 0.029462f
C665 source.n505 a_n2982_n5888# 0.029462f
C666 source.n506 a_n2982_n5888# 0.012831f
C667 source.n507 a_n2982_n5888# 0.012465f
C668 source.n508 a_n2982_n5888# 0.023196f
C669 source.n509 a_n2982_n5888# 0.023196f
C670 source.n510 a_n2982_n5888# 0.012465f
C671 source.n511 a_n2982_n5888# 0.013198f
C672 source.n512 a_n2982_n5888# 0.029462f
C673 source.n513 a_n2982_n5888# 0.029462f
C674 source.n514 a_n2982_n5888# 0.013198f
C675 source.n515 a_n2982_n5888# 0.012465f
C676 source.n516 a_n2982_n5888# 0.023196f
C677 source.n517 a_n2982_n5888# 0.023196f
C678 source.n518 a_n2982_n5888# 0.012465f
C679 source.n519 a_n2982_n5888# 0.013198f
C680 source.n520 a_n2982_n5888# 0.029462f
C681 source.n521 a_n2982_n5888# 0.029462f
C682 source.n522 a_n2982_n5888# 0.013198f
C683 source.n523 a_n2982_n5888# 0.012465f
C684 source.n524 a_n2982_n5888# 0.023196f
C685 source.n525 a_n2982_n5888# 0.023196f
C686 source.n526 a_n2982_n5888# 0.012465f
C687 source.n527 a_n2982_n5888# 0.013198f
C688 source.n528 a_n2982_n5888# 0.029462f
C689 source.n529 a_n2982_n5888# 0.029462f
C690 source.n530 a_n2982_n5888# 0.013198f
C691 source.n531 a_n2982_n5888# 0.012465f
C692 source.n532 a_n2982_n5888# 0.023196f
C693 source.n533 a_n2982_n5888# 0.023196f
C694 source.n534 a_n2982_n5888# 0.012465f
C695 source.n535 a_n2982_n5888# 0.013198f
C696 source.n536 a_n2982_n5888# 0.029462f
C697 source.n537 a_n2982_n5888# 0.029462f
C698 source.n538 a_n2982_n5888# 0.013198f
C699 source.n539 a_n2982_n5888# 0.012465f
C700 source.n540 a_n2982_n5888# 0.023196f
C701 source.n541 a_n2982_n5888# 0.023196f
C702 source.n542 a_n2982_n5888# 0.012465f
C703 source.n543 a_n2982_n5888# 0.013198f
C704 source.n544 a_n2982_n5888# 0.029462f
C705 source.n545 a_n2982_n5888# 0.029462f
C706 source.n546 a_n2982_n5888# 0.013198f
C707 source.n547 a_n2982_n5888# 0.012465f
C708 source.n548 a_n2982_n5888# 0.023196f
C709 source.n549 a_n2982_n5888# 0.023196f
C710 source.n550 a_n2982_n5888# 0.012465f
C711 source.n551 a_n2982_n5888# 0.012831f
C712 source.n552 a_n2982_n5888# 0.012831f
C713 source.n553 a_n2982_n5888# 0.029462f
C714 source.n554 a_n2982_n5888# 0.029462f
C715 source.n555 a_n2982_n5888# 0.013198f
C716 source.n556 a_n2982_n5888# 0.012465f
C717 source.n557 a_n2982_n5888# 0.023196f
C718 source.n558 a_n2982_n5888# 0.023196f
C719 source.n559 a_n2982_n5888# 0.012465f
C720 source.n560 a_n2982_n5888# 0.013198f
C721 source.n561 a_n2982_n5888# 0.029462f
C722 source.n562 a_n2982_n5888# 0.029462f
C723 source.n563 a_n2982_n5888# 0.013198f
C724 source.n564 a_n2982_n5888# 0.012465f
C725 source.n565 a_n2982_n5888# 0.023196f
C726 source.n566 a_n2982_n5888# 0.023196f
C727 source.n567 a_n2982_n5888# 0.012465f
C728 source.n568 a_n2982_n5888# 0.013198f
C729 source.n569 a_n2982_n5888# 0.029462f
C730 source.n570 a_n2982_n5888# 0.062674f
C731 source.n571 a_n2982_n5888# 0.013198f
C732 source.n572 a_n2982_n5888# 0.012465f
C733 source.n573 a_n2982_n5888# 0.051082f
C734 source.n574 a_n2982_n5888# 0.034875f
C735 source.n575 a_n2982_n5888# 2.30373f
C736 source.n576 a_n2982_n5888# 0.031979f
C737 source.n577 a_n2982_n5888# 0.023196f
C738 source.n578 a_n2982_n5888# 0.012465f
C739 source.n579 a_n2982_n5888# 0.029462f
C740 source.n580 a_n2982_n5888# 0.013198f
C741 source.n581 a_n2982_n5888# 0.023196f
C742 source.n582 a_n2982_n5888# 0.012465f
C743 source.n583 a_n2982_n5888# 0.029462f
C744 source.n584 a_n2982_n5888# 0.013198f
C745 source.n585 a_n2982_n5888# 0.023196f
C746 source.n586 a_n2982_n5888# 0.012465f
C747 source.n587 a_n2982_n5888# 0.029462f
C748 source.n588 a_n2982_n5888# 0.013198f
C749 source.n589 a_n2982_n5888# 0.023196f
C750 source.n590 a_n2982_n5888# 0.012465f
C751 source.n591 a_n2982_n5888# 0.029462f
C752 source.n592 a_n2982_n5888# 0.013198f
C753 source.n593 a_n2982_n5888# 0.023196f
C754 source.n594 a_n2982_n5888# 0.012465f
C755 source.n595 a_n2982_n5888# 0.029462f
C756 source.n596 a_n2982_n5888# 0.013198f
C757 source.n597 a_n2982_n5888# 0.023196f
C758 source.n598 a_n2982_n5888# 0.012465f
C759 source.n599 a_n2982_n5888# 0.029462f
C760 source.n600 a_n2982_n5888# 0.013198f
C761 source.n601 a_n2982_n5888# 0.023196f
C762 source.n602 a_n2982_n5888# 0.012465f
C763 source.n603 a_n2982_n5888# 0.029462f
C764 source.n604 a_n2982_n5888# 0.013198f
C765 source.n605 a_n2982_n5888# 0.023196f
C766 source.n606 a_n2982_n5888# 0.012465f
C767 source.n607 a_n2982_n5888# 0.029462f
C768 source.n608 a_n2982_n5888# 0.013198f
C769 source.n609 a_n2982_n5888# 0.023196f
C770 source.n610 a_n2982_n5888# 0.012831f
C771 source.n611 a_n2982_n5888# 0.029462f
C772 source.n612 a_n2982_n5888# 0.013198f
C773 source.n613 a_n2982_n5888# 0.023196f
C774 source.n614 a_n2982_n5888# 0.012465f
C775 source.n615 a_n2982_n5888# 0.029462f
C776 source.n616 a_n2982_n5888# 0.013198f
C777 source.n617 a_n2982_n5888# 0.023196f
C778 source.n618 a_n2982_n5888# 0.012465f
C779 source.n619 a_n2982_n5888# 0.022097f
C780 source.n620 a_n2982_n5888# 0.020828f
C781 source.t2 a_n2982_n5888# 0.051384f
C782 source.n621 a_n2982_n5888# 0.283016f
C783 source.n622 a_n2982_n5888# 2.51149f
C784 source.n623 a_n2982_n5888# 0.012465f
C785 source.n624 a_n2982_n5888# 0.013198f
C786 source.n625 a_n2982_n5888# 0.029462f
C787 source.n626 a_n2982_n5888# 0.029462f
C788 source.n627 a_n2982_n5888# 0.013198f
C789 source.n628 a_n2982_n5888# 0.012465f
C790 source.n629 a_n2982_n5888# 0.023196f
C791 source.n630 a_n2982_n5888# 0.023196f
C792 source.n631 a_n2982_n5888# 0.012465f
C793 source.n632 a_n2982_n5888# 0.013198f
C794 source.n633 a_n2982_n5888# 0.029462f
C795 source.n634 a_n2982_n5888# 0.029462f
C796 source.n635 a_n2982_n5888# 0.013198f
C797 source.n636 a_n2982_n5888# 0.012465f
C798 source.n637 a_n2982_n5888# 0.023196f
C799 source.n638 a_n2982_n5888# 0.023196f
C800 source.n639 a_n2982_n5888# 0.012465f
C801 source.n640 a_n2982_n5888# 0.012465f
C802 source.n641 a_n2982_n5888# 0.013198f
C803 source.n642 a_n2982_n5888# 0.029462f
C804 source.n643 a_n2982_n5888# 0.029462f
C805 source.n644 a_n2982_n5888# 0.029462f
C806 source.n645 a_n2982_n5888# 0.012831f
C807 source.n646 a_n2982_n5888# 0.012465f
C808 source.n647 a_n2982_n5888# 0.023196f
C809 source.n648 a_n2982_n5888# 0.023196f
C810 source.n649 a_n2982_n5888# 0.012465f
C811 source.n650 a_n2982_n5888# 0.013198f
C812 source.n651 a_n2982_n5888# 0.029462f
C813 source.n652 a_n2982_n5888# 0.029462f
C814 source.n653 a_n2982_n5888# 0.013198f
C815 source.n654 a_n2982_n5888# 0.012465f
C816 source.n655 a_n2982_n5888# 0.023196f
C817 source.n656 a_n2982_n5888# 0.023196f
C818 source.n657 a_n2982_n5888# 0.012465f
C819 source.n658 a_n2982_n5888# 0.013198f
C820 source.n659 a_n2982_n5888# 0.029462f
C821 source.n660 a_n2982_n5888# 0.029462f
C822 source.n661 a_n2982_n5888# 0.013198f
C823 source.n662 a_n2982_n5888# 0.012465f
C824 source.n663 a_n2982_n5888# 0.023196f
C825 source.n664 a_n2982_n5888# 0.023196f
C826 source.n665 a_n2982_n5888# 0.012465f
C827 source.n666 a_n2982_n5888# 0.013198f
C828 source.n667 a_n2982_n5888# 0.029462f
C829 source.n668 a_n2982_n5888# 0.029462f
C830 source.n669 a_n2982_n5888# 0.013198f
C831 source.n670 a_n2982_n5888# 0.012465f
C832 source.n671 a_n2982_n5888# 0.023196f
C833 source.n672 a_n2982_n5888# 0.023196f
C834 source.n673 a_n2982_n5888# 0.012465f
C835 source.n674 a_n2982_n5888# 0.013198f
C836 source.n675 a_n2982_n5888# 0.029462f
C837 source.n676 a_n2982_n5888# 0.029462f
C838 source.n677 a_n2982_n5888# 0.013198f
C839 source.n678 a_n2982_n5888# 0.012465f
C840 source.n679 a_n2982_n5888# 0.023196f
C841 source.n680 a_n2982_n5888# 0.023196f
C842 source.n681 a_n2982_n5888# 0.012465f
C843 source.n682 a_n2982_n5888# 0.013198f
C844 source.n683 a_n2982_n5888# 0.029462f
C845 source.n684 a_n2982_n5888# 0.029462f
C846 source.n685 a_n2982_n5888# 0.029462f
C847 source.n686 a_n2982_n5888# 0.013198f
C848 source.n687 a_n2982_n5888# 0.012465f
C849 source.n688 a_n2982_n5888# 0.023196f
C850 source.n689 a_n2982_n5888# 0.023196f
C851 source.n690 a_n2982_n5888# 0.012465f
C852 source.n691 a_n2982_n5888# 0.012831f
C853 source.n692 a_n2982_n5888# 0.012831f
C854 source.n693 a_n2982_n5888# 0.029462f
C855 source.n694 a_n2982_n5888# 0.029462f
C856 source.n695 a_n2982_n5888# 0.013198f
C857 source.n696 a_n2982_n5888# 0.012465f
C858 source.n697 a_n2982_n5888# 0.023196f
C859 source.n698 a_n2982_n5888# 0.023196f
C860 source.n699 a_n2982_n5888# 0.012465f
C861 source.n700 a_n2982_n5888# 0.013198f
C862 source.n701 a_n2982_n5888# 0.029462f
C863 source.n702 a_n2982_n5888# 0.029462f
C864 source.n703 a_n2982_n5888# 0.013198f
C865 source.n704 a_n2982_n5888# 0.012465f
C866 source.n705 a_n2982_n5888# 0.023196f
C867 source.n706 a_n2982_n5888# 0.023196f
C868 source.n707 a_n2982_n5888# 0.012465f
C869 source.n708 a_n2982_n5888# 0.013198f
C870 source.n709 a_n2982_n5888# 0.029462f
C871 source.n710 a_n2982_n5888# 0.062674f
C872 source.n711 a_n2982_n5888# 0.013198f
C873 source.n712 a_n2982_n5888# 0.012465f
C874 source.n713 a_n2982_n5888# 0.051082f
C875 source.n714 a_n2982_n5888# 0.034875f
C876 source.n715 a_n2982_n5888# 2.30373f
C877 source.t14 a_n2982_n5888# 0.458263f
C878 source.t1 a_n2982_n5888# 0.458263f
C879 source.n716 a_n2982_n5888# 4.14734f
C880 source.n717 a_n2982_n5888# 0.37333f
C881 source.t10 a_n2982_n5888# 0.458263f
C882 source.t3 a_n2982_n5888# 0.458263f
C883 source.n718 a_n2982_n5888# 4.14734f
C884 source.n719 a_n2982_n5888# 0.37333f
C885 source.t15 a_n2982_n5888# 0.458263f
C886 source.t39 a_n2982_n5888# 0.458263f
C887 source.n720 a_n2982_n5888# 4.14734f
C888 source.n721 a_n2982_n5888# 0.37333f
C889 source.t7 a_n2982_n5888# 0.458263f
C890 source.t9 a_n2982_n5888# 0.458263f
C891 source.n722 a_n2982_n5888# 4.14734f
C892 source.n723 a_n2982_n5888# 0.37333f
C893 source.n724 a_n2982_n5888# 0.031979f
C894 source.n725 a_n2982_n5888# 0.023196f
C895 source.n726 a_n2982_n5888# 0.012465f
C896 source.n727 a_n2982_n5888# 0.029462f
C897 source.n728 a_n2982_n5888# 0.013198f
C898 source.n729 a_n2982_n5888# 0.023196f
C899 source.n730 a_n2982_n5888# 0.012465f
C900 source.n731 a_n2982_n5888# 0.029462f
C901 source.n732 a_n2982_n5888# 0.013198f
C902 source.n733 a_n2982_n5888# 0.023196f
C903 source.n734 a_n2982_n5888# 0.012465f
C904 source.n735 a_n2982_n5888# 0.029462f
C905 source.n736 a_n2982_n5888# 0.013198f
C906 source.n737 a_n2982_n5888# 0.023196f
C907 source.n738 a_n2982_n5888# 0.012465f
C908 source.n739 a_n2982_n5888# 0.029462f
C909 source.n740 a_n2982_n5888# 0.013198f
C910 source.n741 a_n2982_n5888# 0.023196f
C911 source.n742 a_n2982_n5888# 0.012465f
C912 source.n743 a_n2982_n5888# 0.029462f
C913 source.n744 a_n2982_n5888# 0.013198f
C914 source.n745 a_n2982_n5888# 0.023196f
C915 source.n746 a_n2982_n5888# 0.012465f
C916 source.n747 a_n2982_n5888# 0.029462f
C917 source.n748 a_n2982_n5888# 0.013198f
C918 source.n749 a_n2982_n5888# 0.023196f
C919 source.n750 a_n2982_n5888# 0.012465f
C920 source.n751 a_n2982_n5888# 0.029462f
C921 source.n752 a_n2982_n5888# 0.013198f
C922 source.n753 a_n2982_n5888# 0.023196f
C923 source.n754 a_n2982_n5888# 0.012465f
C924 source.n755 a_n2982_n5888# 0.029462f
C925 source.n756 a_n2982_n5888# 0.013198f
C926 source.n757 a_n2982_n5888# 0.023196f
C927 source.n758 a_n2982_n5888# 0.012831f
C928 source.n759 a_n2982_n5888# 0.029462f
C929 source.n760 a_n2982_n5888# 0.013198f
C930 source.n761 a_n2982_n5888# 0.023196f
C931 source.n762 a_n2982_n5888# 0.012465f
C932 source.n763 a_n2982_n5888# 0.029462f
C933 source.n764 a_n2982_n5888# 0.013198f
C934 source.n765 a_n2982_n5888# 0.023196f
C935 source.n766 a_n2982_n5888# 0.012465f
C936 source.n767 a_n2982_n5888# 0.022097f
C937 source.n768 a_n2982_n5888# 0.020828f
C938 source.t8 a_n2982_n5888# 0.051384f
C939 source.n769 a_n2982_n5888# 0.283016f
C940 source.n770 a_n2982_n5888# 2.51149f
C941 source.n771 a_n2982_n5888# 0.012465f
C942 source.n772 a_n2982_n5888# 0.013198f
C943 source.n773 a_n2982_n5888# 0.029462f
C944 source.n774 a_n2982_n5888# 0.029462f
C945 source.n775 a_n2982_n5888# 0.013198f
C946 source.n776 a_n2982_n5888# 0.012465f
C947 source.n777 a_n2982_n5888# 0.023196f
C948 source.n778 a_n2982_n5888# 0.023196f
C949 source.n779 a_n2982_n5888# 0.012465f
C950 source.n780 a_n2982_n5888# 0.013198f
C951 source.n781 a_n2982_n5888# 0.029462f
C952 source.n782 a_n2982_n5888# 0.029462f
C953 source.n783 a_n2982_n5888# 0.013198f
C954 source.n784 a_n2982_n5888# 0.012465f
C955 source.n785 a_n2982_n5888# 0.023196f
C956 source.n786 a_n2982_n5888# 0.023196f
C957 source.n787 a_n2982_n5888# 0.012465f
C958 source.n788 a_n2982_n5888# 0.012465f
C959 source.n789 a_n2982_n5888# 0.013198f
C960 source.n790 a_n2982_n5888# 0.029462f
C961 source.n791 a_n2982_n5888# 0.029462f
C962 source.n792 a_n2982_n5888# 0.029462f
C963 source.n793 a_n2982_n5888# 0.012831f
C964 source.n794 a_n2982_n5888# 0.012465f
C965 source.n795 a_n2982_n5888# 0.023196f
C966 source.n796 a_n2982_n5888# 0.023196f
C967 source.n797 a_n2982_n5888# 0.012465f
C968 source.n798 a_n2982_n5888# 0.013198f
C969 source.n799 a_n2982_n5888# 0.029462f
C970 source.n800 a_n2982_n5888# 0.029462f
C971 source.n801 a_n2982_n5888# 0.013198f
C972 source.n802 a_n2982_n5888# 0.012465f
C973 source.n803 a_n2982_n5888# 0.023196f
C974 source.n804 a_n2982_n5888# 0.023196f
C975 source.n805 a_n2982_n5888# 0.012465f
C976 source.n806 a_n2982_n5888# 0.013198f
C977 source.n807 a_n2982_n5888# 0.029462f
C978 source.n808 a_n2982_n5888# 0.029462f
C979 source.n809 a_n2982_n5888# 0.013198f
C980 source.n810 a_n2982_n5888# 0.012465f
C981 source.n811 a_n2982_n5888# 0.023196f
C982 source.n812 a_n2982_n5888# 0.023196f
C983 source.n813 a_n2982_n5888# 0.012465f
C984 source.n814 a_n2982_n5888# 0.013198f
C985 source.n815 a_n2982_n5888# 0.029462f
C986 source.n816 a_n2982_n5888# 0.029462f
C987 source.n817 a_n2982_n5888# 0.013198f
C988 source.n818 a_n2982_n5888# 0.012465f
C989 source.n819 a_n2982_n5888# 0.023196f
C990 source.n820 a_n2982_n5888# 0.023196f
C991 source.n821 a_n2982_n5888# 0.012465f
C992 source.n822 a_n2982_n5888# 0.013198f
C993 source.n823 a_n2982_n5888# 0.029462f
C994 source.n824 a_n2982_n5888# 0.029462f
C995 source.n825 a_n2982_n5888# 0.013198f
C996 source.n826 a_n2982_n5888# 0.012465f
C997 source.n827 a_n2982_n5888# 0.023196f
C998 source.n828 a_n2982_n5888# 0.023196f
C999 source.n829 a_n2982_n5888# 0.012465f
C1000 source.n830 a_n2982_n5888# 0.013198f
C1001 source.n831 a_n2982_n5888# 0.029462f
C1002 source.n832 a_n2982_n5888# 0.029462f
C1003 source.n833 a_n2982_n5888# 0.029462f
C1004 source.n834 a_n2982_n5888# 0.013198f
C1005 source.n835 a_n2982_n5888# 0.012465f
C1006 source.n836 a_n2982_n5888# 0.023196f
C1007 source.n837 a_n2982_n5888# 0.023196f
C1008 source.n838 a_n2982_n5888# 0.012465f
C1009 source.n839 a_n2982_n5888# 0.012831f
C1010 source.n840 a_n2982_n5888# 0.012831f
C1011 source.n841 a_n2982_n5888# 0.029462f
C1012 source.n842 a_n2982_n5888# 0.029462f
C1013 source.n843 a_n2982_n5888# 0.013198f
C1014 source.n844 a_n2982_n5888# 0.012465f
C1015 source.n845 a_n2982_n5888# 0.023196f
C1016 source.n846 a_n2982_n5888# 0.023196f
C1017 source.n847 a_n2982_n5888# 0.012465f
C1018 source.n848 a_n2982_n5888# 0.013198f
C1019 source.n849 a_n2982_n5888# 0.029462f
C1020 source.n850 a_n2982_n5888# 0.029462f
C1021 source.n851 a_n2982_n5888# 0.013198f
C1022 source.n852 a_n2982_n5888# 0.012465f
C1023 source.n853 a_n2982_n5888# 0.023196f
C1024 source.n854 a_n2982_n5888# 0.023196f
C1025 source.n855 a_n2982_n5888# 0.012465f
C1026 source.n856 a_n2982_n5888# 0.013198f
C1027 source.n857 a_n2982_n5888# 0.029462f
C1028 source.n858 a_n2982_n5888# 0.062674f
C1029 source.n859 a_n2982_n5888# 0.013198f
C1030 source.n860 a_n2982_n5888# 0.012465f
C1031 source.n861 a_n2982_n5888# 0.051082f
C1032 source.n862 a_n2982_n5888# 0.034875f
C1033 source.n863 a_n2982_n5888# 0.119867f
C1034 source.n864 a_n2982_n5888# 0.031979f
C1035 source.n865 a_n2982_n5888# 0.023196f
C1036 source.n866 a_n2982_n5888# 0.012465f
C1037 source.n867 a_n2982_n5888# 0.029462f
C1038 source.n868 a_n2982_n5888# 0.013198f
C1039 source.n869 a_n2982_n5888# 0.023196f
C1040 source.n870 a_n2982_n5888# 0.012465f
C1041 source.n871 a_n2982_n5888# 0.029462f
C1042 source.n872 a_n2982_n5888# 0.013198f
C1043 source.n873 a_n2982_n5888# 0.023196f
C1044 source.n874 a_n2982_n5888# 0.012465f
C1045 source.n875 a_n2982_n5888# 0.029462f
C1046 source.n876 a_n2982_n5888# 0.013198f
C1047 source.n877 a_n2982_n5888# 0.023196f
C1048 source.n878 a_n2982_n5888# 0.012465f
C1049 source.n879 a_n2982_n5888# 0.029462f
C1050 source.n880 a_n2982_n5888# 0.013198f
C1051 source.n881 a_n2982_n5888# 0.023196f
C1052 source.n882 a_n2982_n5888# 0.012465f
C1053 source.n883 a_n2982_n5888# 0.029462f
C1054 source.n884 a_n2982_n5888# 0.013198f
C1055 source.n885 a_n2982_n5888# 0.023196f
C1056 source.n886 a_n2982_n5888# 0.012465f
C1057 source.n887 a_n2982_n5888# 0.029462f
C1058 source.n888 a_n2982_n5888# 0.013198f
C1059 source.n889 a_n2982_n5888# 0.023196f
C1060 source.n890 a_n2982_n5888# 0.012465f
C1061 source.n891 a_n2982_n5888# 0.029462f
C1062 source.n892 a_n2982_n5888# 0.013198f
C1063 source.n893 a_n2982_n5888# 0.023196f
C1064 source.n894 a_n2982_n5888# 0.012465f
C1065 source.n895 a_n2982_n5888# 0.029462f
C1066 source.n896 a_n2982_n5888# 0.013198f
C1067 source.n897 a_n2982_n5888# 0.023196f
C1068 source.n898 a_n2982_n5888# 0.012831f
C1069 source.n899 a_n2982_n5888# 0.029462f
C1070 source.n900 a_n2982_n5888# 0.013198f
C1071 source.n901 a_n2982_n5888# 0.023196f
C1072 source.n902 a_n2982_n5888# 0.012465f
C1073 source.n903 a_n2982_n5888# 0.029462f
C1074 source.n904 a_n2982_n5888# 0.013198f
C1075 source.n905 a_n2982_n5888# 0.023196f
C1076 source.n906 a_n2982_n5888# 0.012465f
C1077 source.n907 a_n2982_n5888# 0.022097f
C1078 source.n908 a_n2982_n5888# 0.020828f
C1079 source.t33 a_n2982_n5888# 0.051384f
C1080 source.n909 a_n2982_n5888# 0.283016f
C1081 source.n910 a_n2982_n5888# 2.51149f
C1082 source.n911 a_n2982_n5888# 0.012465f
C1083 source.n912 a_n2982_n5888# 0.013198f
C1084 source.n913 a_n2982_n5888# 0.029462f
C1085 source.n914 a_n2982_n5888# 0.029462f
C1086 source.n915 a_n2982_n5888# 0.013198f
C1087 source.n916 a_n2982_n5888# 0.012465f
C1088 source.n917 a_n2982_n5888# 0.023196f
C1089 source.n918 a_n2982_n5888# 0.023196f
C1090 source.n919 a_n2982_n5888# 0.012465f
C1091 source.n920 a_n2982_n5888# 0.013198f
C1092 source.n921 a_n2982_n5888# 0.029462f
C1093 source.n922 a_n2982_n5888# 0.029462f
C1094 source.n923 a_n2982_n5888# 0.013198f
C1095 source.n924 a_n2982_n5888# 0.012465f
C1096 source.n925 a_n2982_n5888# 0.023196f
C1097 source.n926 a_n2982_n5888# 0.023196f
C1098 source.n927 a_n2982_n5888# 0.012465f
C1099 source.n928 a_n2982_n5888# 0.012465f
C1100 source.n929 a_n2982_n5888# 0.013198f
C1101 source.n930 a_n2982_n5888# 0.029462f
C1102 source.n931 a_n2982_n5888# 0.029462f
C1103 source.n932 a_n2982_n5888# 0.029462f
C1104 source.n933 a_n2982_n5888# 0.012831f
C1105 source.n934 a_n2982_n5888# 0.012465f
C1106 source.n935 a_n2982_n5888# 0.023196f
C1107 source.n936 a_n2982_n5888# 0.023196f
C1108 source.n937 a_n2982_n5888# 0.012465f
C1109 source.n938 a_n2982_n5888# 0.013198f
C1110 source.n939 a_n2982_n5888# 0.029462f
C1111 source.n940 a_n2982_n5888# 0.029462f
C1112 source.n941 a_n2982_n5888# 0.013198f
C1113 source.n942 a_n2982_n5888# 0.012465f
C1114 source.n943 a_n2982_n5888# 0.023196f
C1115 source.n944 a_n2982_n5888# 0.023196f
C1116 source.n945 a_n2982_n5888# 0.012465f
C1117 source.n946 a_n2982_n5888# 0.013198f
C1118 source.n947 a_n2982_n5888# 0.029462f
C1119 source.n948 a_n2982_n5888# 0.029462f
C1120 source.n949 a_n2982_n5888# 0.013198f
C1121 source.n950 a_n2982_n5888# 0.012465f
C1122 source.n951 a_n2982_n5888# 0.023196f
C1123 source.n952 a_n2982_n5888# 0.023196f
C1124 source.n953 a_n2982_n5888# 0.012465f
C1125 source.n954 a_n2982_n5888# 0.013198f
C1126 source.n955 a_n2982_n5888# 0.029462f
C1127 source.n956 a_n2982_n5888# 0.029462f
C1128 source.n957 a_n2982_n5888# 0.013198f
C1129 source.n958 a_n2982_n5888# 0.012465f
C1130 source.n959 a_n2982_n5888# 0.023196f
C1131 source.n960 a_n2982_n5888# 0.023196f
C1132 source.n961 a_n2982_n5888# 0.012465f
C1133 source.n962 a_n2982_n5888# 0.013198f
C1134 source.n963 a_n2982_n5888# 0.029462f
C1135 source.n964 a_n2982_n5888# 0.029462f
C1136 source.n965 a_n2982_n5888# 0.013198f
C1137 source.n966 a_n2982_n5888# 0.012465f
C1138 source.n967 a_n2982_n5888# 0.023196f
C1139 source.n968 a_n2982_n5888# 0.023196f
C1140 source.n969 a_n2982_n5888# 0.012465f
C1141 source.n970 a_n2982_n5888# 0.013198f
C1142 source.n971 a_n2982_n5888# 0.029462f
C1143 source.n972 a_n2982_n5888# 0.029462f
C1144 source.n973 a_n2982_n5888# 0.029462f
C1145 source.n974 a_n2982_n5888# 0.013198f
C1146 source.n975 a_n2982_n5888# 0.012465f
C1147 source.n976 a_n2982_n5888# 0.023196f
C1148 source.n977 a_n2982_n5888# 0.023196f
C1149 source.n978 a_n2982_n5888# 0.012465f
C1150 source.n979 a_n2982_n5888# 0.012831f
C1151 source.n980 a_n2982_n5888# 0.012831f
C1152 source.n981 a_n2982_n5888# 0.029462f
C1153 source.n982 a_n2982_n5888# 0.029462f
C1154 source.n983 a_n2982_n5888# 0.013198f
C1155 source.n984 a_n2982_n5888# 0.012465f
C1156 source.n985 a_n2982_n5888# 0.023196f
C1157 source.n986 a_n2982_n5888# 0.023196f
C1158 source.n987 a_n2982_n5888# 0.012465f
C1159 source.n988 a_n2982_n5888# 0.013198f
C1160 source.n989 a_n2982_n5888# 0.029462f
C1161 source.n990 a_n2982_n5888# 0.029462f
C1162 source.n991 a_n2982_n5888# 0.013198f
C1163 source.n992 a_n2982_n5888# 0.012465f
C1164 source.n993 a_n2982_n5888# 0.023196f
C1165 source.n994 a_n2982_n5888# 0.023196f
C1166 source.n995 a_n2982_n5888# 0.012465f
C1167 source.n996 a_n2982_n5888# 0.013198f
C1168 source.n997 a_n2982_n5888# 0.029462f
C1169 source.n998 a_n2982_n5888# 0.062674f
C1170 source.n999 a_n2982_n5888# 0.013198f
C1171 source.n1000 a_n2982_n5888# 0.012465f
C1172 source.n1001 a_n2982_n5888# 0.051082f
C1173 source.n1002 a_n2982_n5888# 0.034875f
C1174 source.n1003 a_n2982_n5888# 0.119867f
C1175 source.t34 a_n2982_n5888# 0.458263f
C1176 source.t38 a_n2982_n5888# 0.458263f
C1177 source.n1004 a_n2982_n5888# 4.14734f
C1178 source.n1005 a_n2982_n5888# 0.37333f
C1179 source.t37 a_n2982_n5888# 0.458263f
C1180 source.t35 a_n2982_n5888# 0.458263f
C1181 source.n1006 a_n2982_n5888# 4.14734f
C1182 source.n1007 a_n2982_n5888# 0.37333f
C1183 source.t22 a_n2982_n5888# 0.458263f
C1184 source.t21 a_n2982_n5888# 0.458263f
C1185 source.n1008 a_n2982_n5888# 4.14734f
C1186 source.n1009 a_n2982_n5888# 0.37333f
C1187 source.t25 a_n2982_n5888# 0.458263f
C1188 source.t26 a_n2982_n5888# 0.458263f
C1189 source.n1010 a_n2982_n5888# 4.14734f
C1190 source.n1011 a_n2982_n5888# 0.37333f
C1191 source.n1012 a_n2982_n5888# 0.031979f
C1192 source.n1013 a_n2982_n5888# 0.023196f
C1193 source.n1014 a_n2982_n5888# 0.012465f
C1194 source.n1015 a_n2982_n5888# 0.029462f
C1195 source.n1016 a_n2982_n5888# 0.013198f
C1196 source.n1017 a_n2982_n5888# 0.023196f
C1197 source.n1018 a_n2982_n5888# 0.012465f
C1198 source.n1019 a_n2982_n5888# 0.029462f
C1199 source.n1020 a_n2982_n5888# 0.013198f
C1200 source.n1021 a_n2982_n5888# 0.023196f
C1201 source.n1022 a_n2982_n5888# 0.012465f
C1202 source.n1023 a_n2982_n5888# 0.029462f
C1203 source.n1024 a_n2982_n5888# 0.013198f
C1204 source.n1025 a_n2982_n5888# 0.023196f
C1205 source.n1026 a_n2982_n5888# 0.012465f
C1206 source.n1027 a_n2982_n5888# 0.029462f
C1207 source.n1028 a_n2982_n5888# 0.013198f
C1208 source.n1029 a_n2982_n5888# 0.023196f
C1209 source.n1030 a_n2982_n5888# 0.012465f
C1210 source.n1031 a_n2982_n5888# 0.029462f
C1211 source.n1032 a_n2982_n5888# 0.013198f
C1212 source.n1033 a_n2982_n5888# 0.023196f
C1213 source.n1034 a_n2982_n5888# 0.012465f
C1214 source.n1035 a_n2982_n5888# 0.029462f
C1215 source.n1036 a_n2982_n5888# 0.013198f
C1216 source.n1037 a_n2982_n5888# 0.023196f
C1217 source.n1038 a_n2982_n5888# 0.012465f
C1218 source.n1039 a_n2982_n5888# 0.029462f
C1219 source.n1040 a_n2982_n5888# 0.013198f
C1220 source.n1041 a_n2982_n5888# 0.023196f
C1221 source.n1042 a_n2982_n5888# 0.012465f
C1222 source.n1043 a_n2982_n5888# 0.029462f
C1223 source.n1044 a_n2982_n5888# 0.013198f
C1224 source.n1045 a_n2982_n5888# 0.023196f
C1225 source.n1046 a_n2982_n5888# 0.012831f
C1226 source.n1047 a_n2982_n5888# 0.029462f
C1227 source.n1048 a_n2982_n5888# 0.013198f
C1228 source.n1049 a_n2982_n5888# 0.023196f
C1229 source.n1050 a_n2982_n5888# 0.012465f
C1230 source.n1051 a_n2982_n5888# 0.029462f
C1231 source.n1052 a_n2982_n5888# 0.013198f
C1232 source.n1053 a_n2982_n5888# 0.023196f
C1233 source.n1054 a_n2982_n5888# 0.012465f
C1234 source.n1055 a_n2982_n5888# 0.022097f
C1235 source.n1056 a_n2982_n5888# 0.020828f
C1236 source.t31 a_n2982_n5888# 0.051384f
C1237 source.n1057 a_n2982_n5888# 0.283016f
C1238 source.n1058 a_n2982_n5888# 2.51149f
C1239 source.n1059 a_n2982_n5888# 0.012465f
C1240 source.n1060 a_n2982_n5888# 0.013198f
C1241 source.n1061 a_n2982_n5888# 0.029462f
C1242 source.n1062 a_n2982_n5888# 0.029462f
C1243 source.n1063 a_n2982_n5888# 0.013198f
C1244 source.n1064 a_n2982_n5888# 0.012465f
C1245 source.n1065 a_n2982_n5888# 0.023196f
C1246 source.n1066 a_n2982_n5888# 0.023196f
C1247 source.n1067 a_n2982_n5888# 0.012465f
C1248 source.n1068 a_n2982_n5888# 0.013198f
C1249 source.n1069 a_n2982_n5888# 0.029462f
C1250 source.n1070 a_n2982_n5888# 0.029462f
C1251 source.n1071 a_n2982_n5888# 0.013198f
C1252 source.n1072 a_n2982_n5888# 0.012465f
C1253 source.n1073 a_n2982_n5888# 0.023196f
C1254 source.n1074 a_n2982_n5888# 0.023196f
C1255 source.n1075 a_n2982_n5888# 0.012465f
C1256 source.n1076 a_n2982_n5888# 0.012465f
C1257 source.n1077 a_n2982_n5888# 0.013198f
C1258 source.n1078 a_n2982_n5888# 0.029462f
C1259 source.n1079 a_n2982_n5888# 0.029462f
C1260 source.n1080 a_n2982_n5888# 0.029462f
C1261 source.n1081 a_n2982_n5888# 0.012831f
C1262 source.n1082 a_n2982_n5888# 0.012465f
C1263 source.n1083 a_n2982_n5888# 0.023196f
C1264 source.n1084 a_n2982_n5888# 0.023196f
C1265 source.n1085 a_n2982_n5888# 0.012465f
C1266 source.n1086 a_n2982_n5888# 0.013198f
C1267 source.n1087 a_n2982_n5888# 0.029462f
C1268 source.n1088 a_n2982_n5888# 0.029462f
C1269 source.n1089 a_n2982_n5888# 0.013198f
C1270 source.n1090 a_n2982_n5888# 0.012465f
C1271 source.n1091 a_n2982_n5888# 0.023196f
C1272 source.n1092 a_n2982_n5888# 0.023196f
C1273 source.n1093 a_n2982_n5888# 0.012465f
C1274 source.n1094 a_n2982_n5888# 0.013198f
C1275 source.n1095 a_n2982_n5888# 0.029462f
C1276 source.n1096 a_n2982_n5888# 0.029462f
C1277 source.n1097 a_n2982_n5888# 0.013198f
C1278 source.n1098 a_n2982_n5888# 0.012465f
C1279 source.n1099 a_n2982_n5888# 0.023196f
C1280 source.n1100 a_n2982_n5888# 0.023196f
C1281 source.n1101 a_n2982_n5888# 0.012465f
C1282 source.n1102 a_n2982_n5888# 0.013198f
C1283 source.n1103 a_n2982_n5888# 0.029462f
C1284 source.n1104 a_n2982_n5888# 0.029462f
C1285 source.n1105 a_n2982_n5888# 0.013198f
C1286 source.n1106 a_n2982_n5888# 0.012465f
C1287 source.n1107 a_n2982_n5888# 0.023196f
C1288 source.n1108 a_n2982_n5888# 0.023196f
C1289 source.n1109 a_n2982_n5888# 0.012465f
C1290 source.n1110 a_n2982_n5888# 0.013198f
C1291 source.n1111 a_n2982_n5888# 0.029462f
C1292 source.n1112 a_n2982_n5888# 0.029462f
C1293 source.n1113 a_n2982_n5888# 0.013198f
C1294 source.n1114 a_n2982_n5888# 0.012465f
C1295 source.n1115 a_n2982_n5888# 0.023196f
C1296 source.n1116 a_n2982_n5888# 0.023196f
C1297 source.n1117 a_n2982_n5888# 0.012465f
C1298 source.n1118 a_n2982_n5888# 0.013198f
C1299 source.n1119 a_n2982_n5888# 0.029462f
C1300 source.n1120 a_n2982_n5888# 0.029462f
C1301 source.n1121 a_n2982_n5888# 0.029462f
C1302 source.n1122 a_n2982_n5888# 0.013198f
C1303 source.n1123 a_n2982_n5888# 0.012465f
C1304 source.n1124 a_n2982_n5888# 0.023196f
C1305 source.n1125 a_n2982_n5888# 0.023196f
C1306 source.n1126 a_n2982_n5888# 0.012465f
C1307 source.n1127 a_n2982_n5888# 0.012831f
C1308 source.n1128 a_n2982_n5888# 0.012831f
C1309 source.n1129 a_n2982_n5888# 0.029462f
C1310 source.n1130 a_n2982_n5888# 0.029462f
C1311 source.n1131 a_n2982_n5888# 0.013198f
C1312 source.n1132 a_n2982_n5888# 0.012465f
C1313 source.n1133 a_n2982_n5888# 0.023196f
C1314 source.n1134 a_n2982_n5888# 0.023196f
C1315 source.n1135 a_n2982_n5888# 0.012465f
C1316 source.n1136 a_n2982_n5888# 0.013198f
C1317 source.n1137 a_n2982_n5888# 0.029462f
C1318 source.n1138 a_n2982_n5888# 0.029462f
C1319 source.n1139 a_n2982_n5888# 0.013198f
C1320 source.n1140 a_n2982_n5888# 0.012465f
C1321 source.n1141 a_n2982_n5888# 0.023196f
C1322 source.n1142 a_n2982_n5888# 0.023196f
C1323 source.n1143 a_n2982_n5888# 0.012465f
C1324 source.n1144 a_n2982_n5888# 0.013198f
C1325 source.n1145 a_n2982_n5888# 0.029462f
C1326 source.n1146 a_n2982_n5888# 0.062674f
C1327 source.n1147 a_n2982_n5888# 0.013198f
C1328 source.n1148 a_n2982_n5888# 0.012465f
C1329 source.n1149 a_n2982_n5888# 0.051082f
C1330 source.n1150 a_n2982_n5888# 0.034875f
C1331 source.n1151 a_n2982_n5888# 0.271178f
C1332 source.n1152 a_n2982_n5888# 2.48982f
C1333 drain_right.t11 a_n2982_n5888# 0.537846f
C1334 drain_right.t12 a_n2982_n5888# 0.537846f
C1335 drain_right.n0 a_n2982_n5888# 4.96275f
C1336 drain_right.t10 a_n2982_n5888# 0.537846f
C1337 drain_right.t9 a_n2982_n5888# 0.537846f
C1338 drain_right.n1 a_n2982_n5888# 4.95683f
C1339 drain_right.n2 a_n2982_n5888# 0.772786f
C1340 drain_right.t13 a_n2982_n5888# 0.537846f
C1341 drain_right.t15 a_n2982_n5888# 0.537846f
C1342 drain_right.n3 a_n2982_n5888# 4.95683f
C1343 drain_right.t19 a_n2982_n5888# 0.537846f
C1344 drain_right.t4 a_n2982_n5888# 0.537846f
C1345 drain_right.n4 a_n2982_n5888# 4.96275f
C1346 drain_right.t14 a_n2982_n5888# 0.537846f
C1347 drain_right.t18 a_n2982_n5888# 0.537846f
C1348 drain_right.n5 a_n2982_n5888# 4.95683f
C1349 drain_right.n6 a_n2982_n5888# 0.772786f
C1350 drain_right.n7 a_n2982_n5888# 2.8245f
C1351 drain_right.t8 a_n2982_n5888# 0.537846f
C1352 drain_right.t0 a_n2982_n5888# 0.537846f
C1353 drain_right.n8 a_n2982_n5888# 4.96274f
C1354 drain_right.t7 a_n2982_n5888# 0.537846f
C1355 drain_right.t1 a_n2982_n5888# 0.537846f
C1356 drain_right.n9 a_n2982_n5888# 4.95684f
C1357 drain_right.n10 a_n2982_n5888# 0.776892f
C1358 drain_right.t6 a_n2982_n5888# 0.537846f
C1359 drain_right.t2 a_n2982_n5888# 0.537846f
C1360 drain_right.n11 a_n2982_n5888# 4.95684f
C1361 drain_right.n12 a_n2982_n5888# 0.385914f
C1362 drain_right.t16 a_n2982_n5888# 0.537846f
C1363 drain_right.t3 a_n2982_n5888# 0.537846f
C1364 drain_right.n13 a_n2982_n5888# 4.95684f
C1365 drain_right.n14 a_n2982_n5888# 0.385914f
C1366 drain_right.t17 a_n2982_n5888# 0.537846f
C1367 drain_right.t5 a_n2982_n5888# 0.537846f
C1368 drain_right.n15 a_n2982_n5888# 4.95684f
C1369 drain_right.n16 a_n2982_n5888# 0.626718f
C1370 minus.n0 a_n2982_n5888# 0.039326f
C1371 minus.n1 a_n2982_n5888# 0.008924f
C1372 minus.t6 a_n2982_n5888# 1.94488f
C1373 minus.n2 a_n2982_n5888# 0.039326f
C1374 minus.n3 a_n2982_n5888# 0.008924f
C1375 minus.t8 a_n2982_n5888# 1.94488f
C1376 minus.n4 a_n2982_n5888# 0.039326f
C1377 minus.n5 a_n2982_n5888# 0.008924f
C1378 minus.t9 a_n2982_n5888# 1.94488f
C1379 minus.n6 a_n2982_n5888# 0.039326f
C1380 minus.n7 a_n2982_n5888# 0.008924f
C1381 minus.t10 a_n2982_n5888# 1.94488f
C1382 minus.t11 a_n2982_n5888# 1.96402f
C1383 minus.t2 a_n2982_n5888# 1.94488f
C1384 minus.n8 a_n2982_n5888# 0.716555f
C1385 minus.n9 a_n2982_n5888# 0.693656f
C1386 minus.n10 a_n2982_n5888# 0.167859f
C1387 minus.n11 a_n2982_n5888# 0.039326f
C1388 minus.n12 a_n2982_n5888# 0.709977f
C1389 minus.n13 a_n2982_n5888# 0.008924f
C1390 minus.t18 a_n2982_n5888# 1.94488f
C1391 minus.n14 a_n2982_n5888# 0.709977f
C1392 minus.n15 a_n2982_n5888# 0.039326f
C1393 minus.n16 a_n2982_n5888# 0.039326f
C1394 minus.n17 a_n2982_n5888# 0.039326f
C1395 minus.n18 a_n2982_n5888# 0.709977f
C1396 minus.n19 a_n2982_n5888# 0.008924f
C1397 minus.t19 a_n2982_n5888# 1.94488f
C1398 minus.n20 a_n2982_n5888# 0.709977f
C1399 minus.n21 a_n2982_n5888# 0.039326f
C1400 minus.n22 a_n2982_n5888# 0.039326f
C1401 minus.n23 a_n2982_n5888# 0.039326f
C1402 minus.n24 a_n2982_n5888# 0.709977f
C1403 minus.n25 a_n2982_n5888# 0.008924f
C1404 minus.t15 a_n2982_n5888# 1.94488f
C1405 minus.n26 a_n2982_n5888# 0.709977f
C1406 minus.n27 a_n2982_n5888# 0.039326f
C1407 minus.n28 a_n2982_n5888# 0.039326f
C1408 minus.n29 a_n2982_n5888# 0.039326f
C1409 minus.n30 a_n2982_n5888# 0.709977f
C1410 minus.n31 a_n2982_n5888# 0.008924f
C1411 minus.t14 a_n2982_n5888# 1.94488f
C1412 minus.n32 a_n2982_n5888# 0.709614f
C1413 minus.n33 a_n2982_n5888# 2.26429f
C1414 minus.n34 a_n2982_n5888# 0.039326f
C1415 minus.n35 a_n2982_n5888# 0.008924f
C1416 minus.n36 a_n2982_n5888# 0.039326f
C1417 minus.n37 a_n2982_n5888# 0.008924f
C1418 minus.n38 a_n2982_n5888# 0.039326f
C1419 minus.n39 a_n2982_n5888# 0.008924f
C1420 minus.n40 a_n2982_n5888# 0.039326f
C1421 minus.n41 a_n2982_n5888# 0.008924f
C1422 minus.t5 a_n2982_n5888# 1.96402f
C1423 minus.t4 a_n2982_n5888# 1.94488f
C1424 minus.n42 a_n2982_n5888# 0.716555f
C1425 minus.n43 a_n2982_n5888# 0.693656f
C1426 minus.n44 a_n2982_n5888# 0.167859f
C1427 minus.n45 a_n2982_n5888# 0.039326f
C1428 minus.t0 a_n2982_n5888# 1.94488f
C1429 minus.n46 a_n2982_n5888# 0.709977f
C1430 minus.n47 a_n2982_n5888# 0.008924f
C1431 minus.t1 a_n2982_n5888# 1.94488f
C1432 minus.n48 a_n2982_n5888# 0.709977f
C1433 minus.n49 a_n2982_n5888# 0.039326f
C1434 minus.n50 a_n2982_n5888# 0.039326f
C1435 minus.n51 a_n2982_n5888# 0.039326f
C1436 minus.t3 a_n2982_n5888# 1.94488f
C1437 minus.n52 a_n2982_n5888# 0.709977f
C1438 minus.n53 a_n2982_n5888# 0.008924f
C1439 minus.t16 a_n2982_n5888# 1.94488f
C1440 minus.n54 a_n2982_n5888# 0.709977f
C1441 minus.n55 a_n2982_n5888# 0.039326f
C1442 minus.n56 a_n2982_n5888# 0.039326f
C1443 minus.n57 a_n2982_n5888# 0.039326f
C1444 minus.t17 a_n2982_n5888# 1.94488f
C1445 minus.n58 a_n2982_n5888# 0.709977f
C1446 minus.n59 a_n2982_n5888# 0.008924f
C1447 minus.t13 a_n2982_n5888# 1.94488f
C1448 minus.n60 a_n2982_n5888# 0.709977f
C1449 minus.n61 a_n2982_n5888# 0.039326f
C1450 minus.n62 a_n2982_n5888# 0.039326f
C1451 minus.n63 a_n2982_n5888# 0.039326f
C1452 minus.t12 a_n2982_n5888# 1.94488f
C1453 minus.n64 a_n2982_n5888# 0.709977f
C1454 minus.n65 a_n2982_n5888# 0.008924f
C1455 minus.t7 a_n2982_n5888# 1.94488f
C1456 minus.n66 a_n2982_n5888# 0.709614f
C1457 minus.n67 a_n2982_n5888# 0.272471f
C1458 minus.n68 a_n2982_n5888# 2.64262f
.ends

