* NGSPICE file created from diffpair269.ext - technology: sky130A

.subckt diffpair269 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t38 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_left.t22 plus.t1 source.t24 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t21 plus.t2 source.t39 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 source.t43 plus.t3 drain_left.t20 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X4 drain_left.t19 plus.t4 source.t45 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X5 drain_left.t18 plus.t5 source.t41 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X6 source.t11 minus.t0 drain_right.t23 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X7 drain_left.t17 plus.t6 source.t42 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X8 source.t15 minus.t1 drain_right.t22 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X9 drain_right.t21 minus.t2 source.t0 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X11 source.t1 minus.t3 drain_right.t20 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X12 drain_left.t16 plus.t7 source.t44 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X13 source.t25 plus.t8 drain_left.t15 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X14 source.t29 plus.t9 drain_left.t14 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 drain_right.t19 minus.t4 source.t7 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X16 source.t2 minus.t5 drain_right.t18 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X17 drain_right.t17 minus.t6 source.t21 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X18 drain_right.t16 minus.t7 source.t12 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 drain_left.t13 plus.t10 source.t28 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X20 source.t17 minus.t8 drain_right.t15 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X21 a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X22 source.t9 minus.t9 drain_right.t14 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X23 source.t46 plus.t11 drain_left.t12 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X24 drain_left.t11 plus.t12 source.t32 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X25 source.t20 minus.t10 drain_right.t13 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X26 source.t23 minus.t11 drain_right.t12 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X27 source.t16 minus.t12 drain_right.t11 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X28 source.t26 plus.t13 drain_left.t10 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X29 source.t30 plus.t14 drain_left.t9 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X30 source.t33 plus.t15 drain_left.t8 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X31 source.t27 plus.t16 drain_left.t7 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X32 drain_left.t6 plus.t17 source.t40 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X33 drain_right.t10 minus.t13 source.t18 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X34 source.t31 plus.t18 drain_left.t5 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X35 drain_right.t9 minus.t14 source.t8 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X36 source.t14 minus.t15 drain_right.t8 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X37 source.t47 plus.t19 drain_left.t4 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X38 drain_right.t7 minus.t16 source.t19 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X39 source.t34 plus.t20 drain_left.t3 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X40 a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X41 source.t22 minus.t17 drain_right.t6 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X42 a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X43 drain_right.t5 minus.t18 source.t4 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X44 drain_right.t4 minus.t19 source.t10 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X45 drain_left.t2 plus.t21 source.t35 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X46 drain_right.t3 minus.t20 source.t13 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X47 drain_right.t2 minus.t21 source.t5 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X48 drain_right.t1 minus.t22 source.t3 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X49 source.t6 minus.t23 drain_right.t0 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X50 drain_left.t1 plus.t22 source.t36 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X51 source.t37 plus.t23 drain_left.t0 a_n2224_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
R0 plus.n6 plus.t8 731.471
R1 plus.n33 plus.t4 731.471
R2 plus.n42 plus.t17 731.471
R3 plus.n68 plus.t3 731.471
R4 plus.n7 plus.t1 703.721
R5 plus.n8 plus.t16 703.721
R6 plus.n14 plus.t0 703.721
R7 plus.n16 plus.t15 703.721
R8 plus.n3 plus.t22 703.721
R9 plus.n21 plus.t14 703.721
R10 plus.n23 plus.t6 703.721
R11 plus.n24 plus.t19 703.721
R12 plus.n30 plus.t5 703.721
R13 plus.n32 plus.t18 703.721
R14 plus.n44 plus.t11 703.721
R15 plus.n43 plus.t2 703.721
R16 plus.n50 plus.t20 703.721
R17 plus.n52 plus.t21 703.721
R18 plus.n39 plus.t13 703.721
R19 plus.n57 plus.t10 703.721
R20 plus.n59 plus.t23 703.721
R21 plus.n38 plus.t12 703.721
R22 plus.n65 plus.t9 703.721
R23 plus.n67 plus.t7 703.721
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus.n17 plus.n3 30.6732
R75 plus.n22 plus.n21 30.6732
R76 plus.n58 plus.n57 30.6732
R77 plus.n53 plus.n39 30.6732
R78 plus plus.n69 29.0861
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 9.80353
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n290 source.n264 289.615
R119 source.n248 source.n222 289.615
R120 source.n216 source.n190 289.615
R121 source.n174 source.n148 289.615
R122 source.n26 source.n0 289.615
R123 source.n68 source.n42 289.615
R124 source.n100 source.n74 289.615
R125 source.n142 source.n116 289.615
R126 source.n275 source.n274 185
R127 source.n272 source.n271 185
R128 source.n281 source.n280 185
R129 source.n283 source.n282 185
R130 source.n268 source.n267 185
R131 source.n289 source.n288 185
R132 source.n291 source.n290 185
R133 source.n233 source.n232 185
R134 source.n230 source.n229 185
R135 source.n239 source.n238 185
R136 source.n241 source.n240 185
R137 source.n226 source.n225 185
R138 source.n247 source.n246 185
R139 source.n249 source.n248 185
R140 source.n201 source.n200 185
R141 source.n198 source.n197 185
R142 source.n207 source.n206 185
R143 source.n209 source.n208 185
R144 source.n194 source.n193 185
R145 source.n215 source.n214 185
R146 source.n217 source.n216 185
R147 source.n159 source.n158 185
R148 source.n156 source.n155 185
R149 source.n165 source.n164 185
R150 source.n167 source.n166 185
R151 source.n152 source.n151 185
R152 source.n173 source.n172 185
R153 source.n175 source.n174 185
R154 source.n27 source.n26 185
R155 source.n25 source.n24 185
R156 source.n4 source.n3 185
R157 source.n19 source.n18 185
R158 source.n17 source.n16 185
R159 source.n8 source.n7 185
R160 source.n11 source.n10 185
R161 source.n69 source.n68 185
R162 source.n67 source.n66 185
R163 source.n46 source.n45 185
R164 source.n61 source.n60 185
R165 source.n59 source.n58 185
R166 source.n50 source.n49 185
R167 source.n53 source.n52 185
R168 source.n101 source.n100 185
R169 source.n99 source.n98 185
R170 source.n78 source.n77 185
R171 source.n93 source.n92 185
R172 source.n91 source.n90 185
R173 source.n82 source.n81 185
R174 source.n85 source.n84 185
R175 source.n143 source.n142 185
R176 source.n141 source.n140 185
R177 source.n120 source.n119 185
R178 source.n135 source.n134 185
R179 source.n133 source.n132 185
R180 source.n124 source.n123 185
R181 source.n127 source.n126 185
R182 source.t21 source.n273 147.661
R183 source.t14 source.n231 147.661
R184 source.t40 source.n199 147.661
R185 source.t43 source.n157 147.661
R186 source.t45 source.n9 147.661
R187 source.t25 source.n51 147.661
R188 source.t19 source.n83 147.661
R189 source.t22 source.n125 147.661
R190 source.n274 source.n271 104.615
R191 source.n281 source.n271 104.615
R192 source.n282 source.n281 104.615
R193 source.n282 source.n267 104.615
R194 source.n289 source.n267 104.615
R195 source.n290 source.n289 104.615
R196 source.n232 source.n229 104.615
R197 source.n239 source.n229 104.615
R198 source.n240 source.n239 104.615
R199 source.n240 source.n225 104.615
R200 source.n247 source.n225 104.615
R201 source.n248 source.n247 104.615
R202 source.n200 source.n197 104.615
R203 source.n207 source.n197 104.615
R204 source.n208 source.n207 104.615
R205 source.n208 source.n193 104.615
R206 source.n215 source.n193 104.615
R207 source.n216 source.n215 104.615
R208 source.n158 source.n155 104.615
R209 source.n165 source.n155 104.615
R210 source.n166 source.n165 104.615
R211 source.n166 source.n151 104.615
R212 source.n173 source.n151 104.615
R213 source.n174 source.n173 104.615
R214 source.n26 source.n25 104.615
R215 source.n25 source.n3 104.615
R216 source.n18 source.n3 104.615
R217 source.n18 source.n17 104.615
R218 source.n17 source.n7 104.615
R219 source.n10 source.n7 104.615
R220 source.n68 source.n67 104.615
R221 source.n67 source.n45 104.615
R222 source.n60 source.n45 104.615
R223 source.n60 source.n59 104.615
R224 source.n59 source.n49 104.615
R225 source.n52 source.n49 104.615
R226 source.n100 source.n99 104.615
R227 source.n99 source.n77 104.615
R228 source.n92 source.n77 104.615
R229 source.n92 source.n91 104.615
R230 source.n91 source.n81 104.615
R231 source.n84 source.n81 104.615
R232 source.n142 source.n141 104.615
R233 source.n141 source.n119 104.615
R234 source.n134 source.n119 104.615
R235 source.n134 source.n133 104.615
R236 source.n133 source.n123 104.615
R237 source.n126 source.n123 104.615
R238 source.n274 source.t21 52.3082
R239 source.n232 source.t14 52.3082
R240 source.n200 source.t40 52.3082
R241 source.n158 source.t43 52.3082
R242 source.n10 source.t45 52.3082
R243 source.n52 source.t25 52.3082
R244 source.n84 source.t19 52.3082
R245 source.n126 source.t22 52.3082
R246 source.n33 source.n32 50.512
R247 source.n35 source.n34 50.512
R248 source.n37 source.n36 50.512
R249 source.n39 source.n38 50.512
R250 source.n41 source.n40 50.512
R251 source.n107 source.n106 50.512
R252 source.n109 source.n108 50.512
R253 source.n111 source.n110 50.512
R254 source.n113 source.n112 50.512
R255 source.n115 source.n114 50.512
R256 source.n263 source.n262 50.5119
R257 source.n261 source.n260 50.5119
R258 source.n259 source.n258 50.5119
R259 source.n257 source.n256 50.5119
R260 source.n255 source.n254 50.5119
R261 source.n189 source.n188 50.5119
R262 source.n187 source.n186 50.5119
R263 source.n185 source.n184 50.5119
R264 source.n183 source.n182 50.5119
R265 source.n181 source.n180 50.5119
R266 source.n295 source.n294 32.1853
R267 source.n253 source.n252 32.1853
R268 source.n221 source.n220 32.1853
R269 source.n179 source.n178 32.1853
R270 source.n31 source.n30 32.1853
R271 source.n73 source.n72 32.1853
R272 source.n105 source.n104 32.1853
R273 source.n147 source.n146 32.1853
R274 source.n179 source.n147 17.2423
R275 source.n275 source.n273 15.6674
R276 source.n233 source.n231 15.6674
R277 source.n201 source.n199 15.6674
R278 source.n159 source.n157 15.6674
R279 source.n11 source.n9 15.6674
R280 source.n53 source.n51 15.6674
R281 source.n85 source.n83 15.6674
R282 source.n127 source.n125 15.6674
R283 source.n276 source.n272 12.8005
R284 source.n234 source.n230 12.8005
R285 source.n202 source.n198 12.8005
R286 source.n160 source.n156 12.8005
R287 source.n12 source.n8 12.8005
R288 source.n54 source.n50 12.8005
R289 source.n86 source.n82 12.8005
R290 source.n128 source.n124 12.8005
R291 source.n280 source.n279 12.0247
R292 source.n238 source.n237 12.0247
R293 source.n206 source.n205 12.0247
R294 source.n164 source.n163 12.0247
R295 source.n16 source.n15 12.0247
R296 source.n58 source.n57 12.0247
R297 source.n90 source.n89 12.0247
R298 source.n132 source.n131 12.0247
R299 source.n296 source.n31 11.7293
R300 source.n283 source.n270 11.249
R301 source.n241 source.n228 11.249
R302 source.n209 source.n196 11.249
R303 source.n167 source.n154 11.249
R304 source.n19 source.n6 11.249
R305 source.n61 source.n48 11.249
R306 source.n93 source.n80 11.249
R307 source.n135 source.n122 11.249
R308 source.n284 source.n268 10.4732
R309 source.n242 source.n226 10.4732
R310 source.n210 source.n194 10.4732
R311 source.n168 source.n152 10.4732
R312 source.n20 source.n4 10.4732
R313 source.n62 source.n46 10.4732
R314 source.n94 source.n78 10.4732
R315 source.n136 source.n120 10.4732
R316 source.n288 source.n287 9.69747
R317 source.n246 source.n245 9.69747
R318 source.n214 source.n213 9.69747
R319 source.n172 source.n171 9.69747
R320 source.n24 source.n23 9.69747
R321 source.n66 source.n65 9.69747
R322 source.n98 source.n97 9.69747
R323 source.n140 source.n139 9.69747
R324 source.n294 source.n293 9.45567
R325 source.n252 source.n251 9.45567
R326 source.n220 source.n219 9.45567
R327 source.n178 source.n177 9.45567
R328 source.n30 source.n29 9.45567
R329 source.n72 source.n71 9.45567
R330 source.n104 source.n103 9.45567
R331 source.n146 source.n145 9.45567
R332 source.n293 source.n292 9.3005
R333 source.n266 source.n265 9.3005
R334 source.n287 source.n286 9.3005
R335 source.n285 source.n284 9.3005
R336 source.n270 source.n269 9.3005
R337 source.n279 source.n278 9.3005
R338 source.n277 source.n276 9.3005
R339 source.n251 source.n250 9.3005
R340 source.n224 source.n223 9.3005
R341 source.n245 source.n244 9.3005
R342 source.n243 source.n242 9.3005
R343 source.n228 source.n227 9.3005
R344 source.n237 source.n236 9.3005
R345 source.n235 source.n234 9.3005
R346 source.n219 source.n218 9.3005
R347 source.n192 source.n191 9.3005
R348 source.n213 source.n212 9.3005
R349 source.n211 source.n210 9.3005
R350 source.n196 source.n195 9.3005
R351 source.n205 source.n204 9.3005
R352 source.n203 source.n202 9.3005
R353 source.n177 source.n176 9.3005
R354 source.n150 source.n149 9.3005
R355 source.n171 source.n170 9.3005
R356 source.n169 source.n168 9.3005
R357 source.n154 source.n153 9.3005
R358 source.n163 source.n162 9.3005
R359 source.n161 source.n160 9.3005
R360 source.n29 source.n28 9.3005
R361 source.n2 source.n1 9.3005
R362 source.n23 source.n22 9.3005
R363 source.n21 source.n20 9.3005
R364 source.n6 source.n5 9.3005
R365 source.n15 source.n14 9.3005
R366 source.n13 source.n12 9.3005
R367 source.n71 source.n70 9.3005
R368 source.n44 source.n43 9.3005
R369 source.n65 source.n64 9.3005
R370 source.n63 source.n62 9.3005
R371 source.n48 source.n47 9.3005
R372 source.n57 source.n56 9.3005
R373 source.n55 source.n54 9.3005
R374 source.n103 source.n102 9.3005
R375 source.n76 source.n75 9.3005
R376 source.n97 source.n96 9.3005
R377 source.n95 source.n94 9.3005
R378 source.n80 source.n79 9.3005
R379 source.n89 source.n88 9.3005
R380 source.n87 source.n86 9.3005
R381 source.n145 source.n144 9.3005
R382 source.n118 source.n117 9.3005
R383 source.n139 source.n138 9.3005
R384 source.n137 source.n136 9.3005
R385 source.n122 source.n121 9.3005
R386 source.n131 source.n130 9.3005
R387 source.n129 source.n128 9.3005
R388 source.n291 source.n266 8.92171
R389 source.n249 source.n224 8.92171
R390 source.n217 source.n192 8.92171
R391 source.n175 source.n150 8.92171
R392 source.n27 source.n2 8.92171
R393 source.n69 source.n44 8.92171
R394 source.n101 source.n76 8.92171
R395 source.n143 source.n118 8.92171
R396 source.n292 source.n264 8.14595
R397 source.n250 source.n222 8.14595
R398 source.n218 source.n190 8.14595
R399 source.n176 source.n148 8.14595
R400 source.n28 source.n0 8.14595
R401 source.n70 source.n42 8.14595
R402 source.n102 source.n74 8.14595
R403 source.n144 source.n116 8.14595
R404 source.n294 source.n264 5.81868
R405 source.n252 source.n222 5.81868
R406 source.n220 source.n190 5.81868
R407 source.n178 source.n148 5.81868
R408 source.n30 source.n0 5.81868
R409 source.n72 source.n42 5.81868
R410 source.n104 source.n74 5.81868
R411 source.n146 source.n116 5.81868
R412 source.n296 source.n295 5.51343
R413 source.n292 source.n291 5.04292
R414 source.n250 source.n249 5.04292
R415 source.n218 source.n217 5.04292
R416 source.n176 source.n175 5.04292
R417 source.n28 source.n27 5.04292
R418 source.n70 source.n69 5.04292
R419 source.n102 source.n101 5.04292
R420 source.n144 source.n143 5.04292
R421 source.n277 source.n273 4.38594
R422 source.n235 source.n231 4.38594
R423 source.n203 source.n199 4.38594
R424 source.n161 source.n157 4.38594
R425 source.n13 source.n9 4.38594
R426 source.n55 source.n51 4.38594
R427 source.n87 source.n83 4.38594
R428 source.n129 source.n125 4.38594
R429 source.n288 source.n266 4.26717
R430 source.n246 source.n224 4.26717
R431 source.n214 source.n192 4.26717
R432 source.n172 source.n150 4.26717
R433 source.n24 source.n2 4.26717
R434 source.n66 source.n44 4.26717
R435 source.n98 source.n76 4.26717
R436 source.n140 source.n118 4.26717
R437 source.n287 source.n268 3.49141
R438 source.n245 source.n226 3.49141
R439 source.n213 source.n194 3.49141
R440 source.n171 source.n152 3.49141
R441 source.n23 source.n4 3.49141
R442 source.n65 source.n46 3.49141
R443 source.n97 source.n78 3.49141
R444 source.n139 source.n120 3.49141
R445 source.n262 source.t10 3.3005
R446 source.n262 source.t16 3.3005
R447 source.n260 source.t12 3.3005
R448 source.n260 source.t1 3.3005
R449 source.n258 source.t18 3.3005
R450 source.n258 source.t9 3.3005
R451 source.n256 source.t7 3.3005
R452 source.n256 source.t6 3.3005
R453 source.n254 source.t4 3.3005
R454 source.n254 source.t23 3.3005
R455 source.n188 source.t39 3.3005
R456 source.n188 source.t46 3.3005
R457 source.n186 source.t35 3.3005
R458 source.n186 source.t34 3.3005
R459 source.n184 source.t28 3.3005
R460 source.n184 source.t26 3.3005
R461 source.n182 source.t32 3.3005
R462 source.n182 source.t37 3.3005
R463 source.n180 source.t44 3.3005
R464 source.n180 source.t29 3.3005
R465 source.n32 source.t41 3.3005
R466 source.n32 source.t31 3.3005
R467 source.n34 source.t42 3.3005
R468 source.n34 source.t47 3.3005
R469 source.n36 source.t36 3.3005
R470 source.n36 source.t30 3.3005
R471 source.n38 source.t38 3.3005
R472 source.n38 source.t33 3.3005
R473 source.n40 source.t24 3.3005
R474 source.n40 source.t27 3.3005
R475 source.n106 source.t8 3.3005
R476 source.n106 source.t15 3.3005
R477 source.n108 source.t13 3.3005
R478 source.n108 source.t11 3.3005
R479 source.n110 source.t5 3.3005
R480 source.n110 source.t17 3.3005
R481 source.n112 source.t3 3.3005
R482 source.n112 source.t2 3.3005
R483 source.n114 source.t0 3.3005
R484 source.n114 source.t20 3.3005
R485 source.n284 source.n283 2.71565
R486 source.n242 source.n241 2.71565
R487 source.n210 source.n209 2.71565
R488 source.n168 source.n167 2.71565
R489 source.n20 source.n19 2.71565
R490 source.n62 source.n61 2.71565
R491 source.n94 source.n93 2.71565
R492 source.n136 source.n135 2.71565
R493 source.n280 source.n270 1.93989
R494 source.n238 source.n228 1.93989
R495 source.n206 source.n196 1.93989
R496 source.n164 source.n154 1.93989
R497 source.n16 source.n6 1.93989
R498 source.n58 source.n48 1.93989
R499 source.n90 source.n80 1.93989
R500 source.n132 source.n122 1.93989
R501 source.n279 source.n272 1.16414
R502 source.n237 source.n230 1.16414
R503 source.n205 source.n198 1.16414
R504 source.n163 source.n156 1.16414
R505 source.n15 source.n8 1.16414
R506 source.n57 source.n50 1.16414
R507 source.n89 source.n82 1.16414
R508 source.n131 source.n124 1.16414
R509 source.n147 source.n115 0.5005
R510 source.n115 source.n113 0.5005
R511 source.n113 source.n111 0.5005
R512 source.n111 source.n109 0.5005
R513 source.n109 source.n107 0.5005
R514 source.n107 source.n105 0.5005
R515 source.n73 source.n41 0.5005
R516 source.n41 source.n39 0.5005
R517 source.n39 source.n37 0.5005
R518 source.n37 source.n35 0.5005
R519 source.n35 source.n33 0.5005
R520 source.n33 source.n31 0.5005
R521 source.n181 source.n179 0.5005
R522 source.n183 source.n181 0.5005
R523 source.n185 source.n183 0.5005
R524 source.n187 source.n185 0.5005
R525 source.n189 source.n187 0.5005
R526 source.n221 source.n189 0.5005
R527 source.n255 source.n253 0.5005
R528 source.n257 source.n255 0.5005
R529 source.n259 source.n257 0.5005
R530 source.n261 source.n259 0.5005
R531 source.n263 source.n261 0.5005
R532 source.n295 source.n263 0.5005
R533 source.n105 source.n73 0.470328
R534 source.n253 source.n221 0.470328
R535 source.n276 source.n275 0.388379
R536 source.n234 source.n233 0.388379
R537 source.n202 source.n201 0.388379
R538 source.n160 source.n159 0.388379
R539 source.n12 source.n11 0.388379
R540 source.n54 source.n53 0.388379
R541 source.n86 source.n85 0.388379
R542 source.n128 source.n127 0.388379
R543 source source.n296 0.188
R544 source.n278 source.n277 0.155672
R545 source.n278 source.n269 0.155672
R546 source.n285 source.n269 0.155672
R547 source.n286 source.n285 0.155672
R548 source.n286 source.n265 0.155672
R549 source.n293 source.n265 0.155672
R550 source.n236 source.n235 0.155672
R551 source.n236 source.n227 0.155672
R552 source.n243 source.n227 0.155672
R553 source.n244 source.n243 0.155672
R554 source.n244 source.n223 0.155672
R555 source.n251 source.n223 0.155672
R556 source.n204 source.n203 0.155672
R557 source.n204 source.n195 0.155672
R558 source.n211 source.n195 0.155672
R559 source.n212 source.n211 0.155672
R560 source.n212 source.n191 0.155672
R561 source.n219 source.n191 0.155672
R562 source.n162 source.n161 0.155672
R563 source.n162 source.n153 0.155672
R564 source.n169 source.n153 0.155672
R565 source.n170 source.n169 0.155672
R566 source.n170 source.n149 0.155672
R567 source.n177 source.n149 0.155672
R568 source.n29 source.n1 0.155672
R569 source.n22 source.n1 0.155672
R570 source.n22 source.n21 0.155672
R571 source.n21 source.n5 0.155672
R572 source.n14 source.n5 0.155672
R573 source.n14 source.n13 0.155672
R574 source.n71 source.n43 0.155672
R575 source.n64 source.n43 0.155672
R576 source.n64 source.n63 0.155672
R577 source.n63 source.n47 0.155672
R578 source.n56 source.n47 0.155672
R579 source.n56 source.n55 0.155672
R580 source.n103 source.n75 0.155672
R581 source.n96 source.n75 0.155672
R582 source.n96 source.n95 0.155672
R583 source.n95 source.n79 0.155672
R584 source.n88 source.n79 0.155672
R585 source.n88 source.n87 0.155672
R586 source.n145 source.n117 0.155672
R587 source.n138 source.n117 0.155672
R588 source.n138 source.n137 0.155672
R589 source.n137 source.n121 0.155672
R590 source.n130 source.n121 0.155672
R591 source.n130 source.n129 0.155672
R592 drain_left.n13 drain_left.n11 67.6908
R593 drain_left.n7 drain_left.n5 67.6907
R594 drain_left.n2 drain_left.n0 67.6907
R595 drain_left.n19 drain_left.n18 67.1908
R596 drain_left.n17 drain_left.n16 67.1908
R597 drain_left.n15 drain_left.n14 67.1908
R598 drain_left.n13 drain_left.n12 67.1908
R599 drain_left.n21 drain_left.n20 67.1907
R600 drain_left.n7 drain_left.n6 67.1907
R601 drain_left.n9 drain_left.n8 67.1907
R602 drain_left.n4 drain_left.n3 67.1907
R603 drain_left.n2 drain_left.n1 67.1907
R604 drain_left drain_left.n10 27.5716
R605 drain_left drain_left.n21 6.15322
R606 drain_left.n5 drain_left.t12 3.3005
R607 drain_left.n5 drain_left.t6 3.3005
R608 drain_left.n6 drain_left.t3 3.3005
R609 drain_left.n6 drain_left.t21 3.3005
R610 drain_left.n8 drain_left.t10 3.3005
R611 drain_left.n8 drain_left.t2 3.3005
R612 drain_left.n3 drain_left.t0 3.3005
R613 drain_left.n3 drain_left.t13 3.3005
R614 drain_left.n1 drain_left.t14 3.3005
R615 drain_left.n1 drain_left.t11 3.3005
R616 drain_left.n0 drain_left.t20 3.3005
R617 drain_left.n0 drain_left.t16 3.3005
R618 drain_left.n20 drain_left.t5 3.3005
R619 drain_left.n20 drain_left.t19 3.3005
R620 drain_left.n18 drain_left.t4 3.3005
R621 drain_left.n18 drain_left.t18 3.3005
R622 drain_left.n16 drain_left.t9 3.3005
R623 drain_left.n16 drain_left.t17 3.3005
R624 drain_left.n14 drain_left.t8 3.3005
R625 drain_left.n14 drain_left.t1 3.3005
R626 drain_left.n12 drain_left.t7 3.3005
R627 drain_left.n12 drain_left.t23 3.3005
R628 drain_left.n11 drain_left.t15 3.3005
R629 drain_left.n11 drain_left.t22 3.3005
R630 drain_left.n9 drain_left.n7 0.5005
R631 drain_left.n4 drain_left.n2 0.5005
R632 drain_left.n15 drain_left.n13 0.5005
R633 drain_left.n17 drain_left.n15 0.5005
R634 drain_left.n19 drain_left.n17 0.5005
R635 drain_left.n21 drain_left.n19 0.5005
R636 drain_left.n10 drain_left.n9 0.195154
R637 drain_left.n10 drain_left.n4 0.195154
R638 minus.n33 minus.t17 731.471
R639 minus.n7 minus.t16 731.471
R640 minus.n68 minus.t6 731.471
R641 minus.n41 minus.t15 731.471
R642 minus.n32 minus.t2 703.721
R643 minus.n30 minus.t10 703.721
R644 minus.n3 minus.t22 703.721
R645 minus.n24 minus.t5 703.721
R646 minus.n22 minus.t21 703.721
R647 minus.n4 minus.t8 703.721
R648 minus.n17 minus.t20 703.721
R649 minus.n15 minus.t0 703.721
R650 minus.n8 minus.t14 703.721
R651 minus.n9 minus.t1 703.721
R652 minus.n67 minus.t12 703.721
R653 minus.n65 minus.t19 703.721
R654 minus.n59 minus.t3 703.721
R655 minus.n58 minus.t7 703.721
R656 minus.n56 minus.t9 703.721
R657 minus.n38 minus.t13 703.721
R658 minus.n51 minus.t23 703.721
R659 minus.n49 minus.t4 703.721
R660 minus.n43 minus.t11 703.721
R661 minus.n42 minus.t18 703.721
R662 minus.n11 minus.n7 161.489
R663 minus.n45 minus.n41 161.489
R664 minus.n34 minus.n33 161.3
R665 minus.n31 minus.n0 161.3
R666 minus.n29 minus.n28 161.3
R667 minus.n27 minus.n1 161.3
R668 minus.n26 minus.n25 161.3
R669 minus.n23 minus.n2 161.3
R670 minus.n21 minus.n20 161.3
R671 minus.n19 minus.n18 161.3
R672 minus.n16 minus.n5 161.3
R673 minus.n14 minus.n13 161.3
R674 minus.n12 minus.n6 161.3
R675 minus.n11 minus.n10 161.3
R676 minus.n69 minus.n68 161.3
R677 minus.n66 minus.n35 161.3
R678 minus.n64 minus.n63 161.3
R679 minus.n62 minus.n36 161.3
R680 minus.n61 minus.n60 161.3
R681 minus.n57 minus.n37 161.3
R682 minus.n55 minus.n54 161.3
R683 minus.n53 minus.n52 161.3
R684 minus.n50 minus.n39 161.3
R685 minus.n48 minus.n47 161.3
R686 minus.n46 minus.n40 161.3
R687 minus.n45 minus.n44 161.3
R688 minus.n29 minus.n1 73.0308
R689 minus.n14 minus.n6 73.0308
R690 minus.n48 minus.n40 73.0308
R691 minus.n64 minus.n36 73.0308
R692 minus.n31 minus.n30 68.649
R693 minus.n10 minus.n8 68.649
R694 minus.n44 minus.n43 68.649
R695 minus.n66 minus.n65 68.649
R696 minus.n25 minus.n3 65.7278
R697 minus.n16 minus.n15 65.7278
R698 minus.n50 minus.n49 65.7278
R699 minus.n60 minus.n59 65.7278
R700 minus.n33 minus.n32 56.9641
R701 minus.n9 minus.n7 56.9641
R702 minus.n42 minus.n41 56.9641
R703 minus.n68 minus.n67 56.9641
R704 minus.n24 minus.n23 54.0429
R705 minus.n18 minus.n17 54.0429
R706 minus.n52 minus.n51 54.0429
R707 minus.n58 minus.n57 54.0429
R708 minus.n22 minus.n21 42.3581
R709 minus.n21 minus.n4 42.3581
R710 minus.n55 minus.n38 42.3581
R711 minus.n56 minus.n55 42.3581
R712 minus.n70 minus.n34 32.9323
R713 minus.n23 minus.n22 30.6732
R714 minus.n18 minus.n4 30.6732
R715 minus.n52 minus.n38 30.6732
R716 minus.n57 minus.n56 30.6732
R717 minus.n25 minus.n24 18.9884
R718 minus.n17 minus.n16 18.9884
R719 minus.n51 minus.n50 18.9884
R720 minus.n60 minus.n58 18.9884
R721 minus.n32 minus.n31 16.0672
R722 minus.n10 minus.n9 16.0672
R723 minus.n44 minus.n42 16.0672
R724 minus.n67 minus.n66 16.0672
R725 minus.n3 minus.n1 7.30353
R726 minus.n15 minus.n14 7.30353
R727 minus.n49 minus.n48 7.30353
R728 minus.n59 minus.n36 7.30353
R729 minus.n70 minus.n69 6.43232
R730 minus.n30 minus.n29 4.38232
R731 minus.n8 minus.n6 4.38232
R732 minus.n43 minus.n40 4.38232
R733 minus.n65 minus.n64 4.38232
R734 minus.n34 minus.n0 0.189894
R735 minus.n28 minus.n0 0.189894
R736 minus.n28 minus.n27 0.189894
R737 minus.n27 minus.n26 0.189894
R738 minus.n26 minus.n2 0.189894
R739 minus.n20 minus.n2 0.189894
R740 minus.n20 minus.n19 0.189894
R741 minus.n19 minus.n5 0.189894
R742 minus.n13 minus.n5 0.189894
R743 minus.n13 minus.n12 0.189894
R744 minus.n12 minus.n11 0.189894
R745 minus.n46 minus.n45 0.189894
R746 minus.n47 minus.n46 0.189894
R747 minus.n47 minus.n39 0.189894
R748 minus.n53 minus.n39 0.189894
R749 minus.n54 minus.n53 0.189894
R750 minus.n54 minus.n37 0.189894
R751 minus.n61 minus.n37 0.189894
R752 minus.n62 minus.n61 0.189894
R753 minus.n63 minus.n62 0.189894
R754 minus.n63 minus.n35 0.189894
R755 minus.n69 minus.n35 0.189894
R756 minus minus.n70 0.188
R757 drain_right.n13 drain_right.n11 67.6907
R758 drain_right.n7 drain_right.n5 67.6907
R759 drain_right.n2 drain_right.n0 67.6907
R760 drain_right.n13 drain_right.n12 67.1908
R761 drain_right.n15 drain_right.n14 67.1908
R762 drain_right.n17 drain_right.n16 67.1908
R763 drain_right.n19 drain_right.n18 67.1908
R764 drain_right.n21 drain_right.n20 67.1908
R765 drain_right.n7 drain_right.n6 67.1907
R766 drain_right.n9 drain_right.n8 67.1907
R767 drain_right.n4 drain_right.n3 67.1907
R768 drain_right.n2 drain_right.n1 67.1907
R769 drain_right drain_right.n10 27.0184
R770 drain_right drain_right.n21 6.15322
R771 drain_right.n5 drain_right.t11 3.3005
R772 drain_right.n5 drain_right.t17 3.3005
R773 drain_right.n6 drain_right.t20 3.3005
R774 drain_right.n6 drain_right.t4 3.3005
R775 drain_right.n8 drain_right.t14 3.3005
R776 drain_right.n8 drain_right.t16 3.3005
R777 drain_right.n3 drain_right.t0 3.3005
R778 drain_right.n3 drain_right.t10 3.3005
R779 drain_right.n1 drain_right.t12 3.3005
R780 drain_right.n1 drain_right.t19 3.3005
R781 drain_right.n0 drain_right.t8 3.3005
R782 drain_right.n0 drain_right.t5 3.3005
R783 drain_right.n11 drain_right.t22 3.3005
R784 drain_right.n11 drain_right.t7 3.3005
R785 drain_right.n12 drain_right.t23 3.3005
R786 drain_right.n12 drain_right.t9 3.3005
R787 drain_right.n14 drain_right.t15 3.3005
R788 drain_right.n14 drain_right.t3 3.3005
R789 drain_right.n16 drain_right.t18 3.3005
R790 drain_right.n16 drain_right.t2 3.3005
R791 drain_right.n18 drain_right.t13 3.3005
R792 drain_right.n18 drain_right.t1 3.3005
R793 drain_right.n20 drain_right.t6 3.3005
R794 drain_right.n20 drain_right.t21 3.3005
R795 drain_right.n9 drain_right.n7 0.5005
R796 drain_right.n4 drain_right.n2 0.5005
R797 drain_right.n21 drain_right.n19 0.5005
R798 drain_right.n19 drain_right.n17 0.5005
R799 drain_right.n17 drain_right.n15 0.5005
R800 drain_right.n15 drain_right.n13 0.5005
R801 drain_right.n10 drain_right.n9 0.195154
R802 drain_right.n10 drain_right.n4 0.195154
C0 source minus 4.06948f
C1 drain_right plus 0.374075f
C2 minus plus 4.82303f
C3 drain_right drain_left 1.19771f
C4 drain_left minus 0.172313f
C5 source plus 4.0835f
C6 drain_left source 26.14f
C7 drain_left plus 4.22756f
C8 drain_right minus 4.00889f
C9 drain_right source 26.1404f
C10 drain_right a_n2224_n2088# 5.98123f
C11 drain_left a_n2224_n2088# 6.32173f
C12 source a_n2224_n2088# 5.49462f
C13 minus a_n2224_n2088# 8.238338f
C14 plus a_n2224_n2088# 9.91725f
C15 drain_right.t8 a_n2224_n2088# 0.168788f
C16 drain_right.t5 a_n2224_n2088# 0.168788f
C17 drain_right.n0 a_n2224_n2088# 1.41078f
C18 drain_right.t12 a_n2224_n2088# 0.168788f
C19 drain_right.t19 a_n2224_n2088# 0.168788f
C20 drain_right.n1 a_n2224_n2088# 1.40769f
C21 drain_right.n2 a_n2224_n2088# 0.818531f
C22 drain_right.t0 a_n2224_n2088# 0.168788f
C23 drain_right.t10 a_n2224_n2088# 0.168788f
C24 drain_right.n3 a_n2224_n2088# 1.40769f
C25 drain_right.n4 a_n2224_n2088# 0.372855f
C26 drain_right.t11 a_n2224_n2088# 0.168788f
C27 drain_right.t17 a_n2224_n2088# 0.168788f
C28 drain_right.n5 a_n2224_n2088# 1.41078f
C29 drain_right.t20 a_n2224_n2088# 0.168788f
C30 drain_right.t4 a_n2224_n2088# 0.168788f
C31 drain_right.n6 a_n2224_n2088# 1.40769f
C32 drain_right.n7 a_n2224_n2088# 0.818531f
C33 drain_right.t14 a_n2224_n2088# 0.168788f
C34 drain_right.t16 a_n2224_n2088# 0.168788f
C35 drain_right.n8 a_n2224_n2088# 1.40769f
C36 drain_right.n9 a_n2224_n2088# 0.372855f
C37 drain_right.n10 a_n2224_n2088# 1.34018f
C38 drain_right.t22 a_n2224_n2088# 0.168788f
C39 drain_right.t7 a_n2224_n2088# 0.168788f
C40 drain_right.n11 a_n2224_n2088# 1.41078f
C41 drain_right.t23 a_n2224_n2088# 0.168788f
C42 drain_right.t9 a_n2224_n2088# 0.168788f
C43 drain_right.n12 a_n2224_n2088# 1.4077f
C44 drain_right.n13 a_n2224_n2088# 0.818525f
C45 drain_right.t15 a_n2224_n2088# 0.168788f
C46 drain_right.t3 a_n2224_n2088# 0.168788f
C47 drain_right.n14 a_n2224_n2088# 1.4077f
C48 drain_right.n15 a_n2224_n2088# 0.403634f
C49 drain_right.t18 a_n2224_n2088# 0.168788f
C50 drain_right.t2 a_n2224_n2088# 0.168788f
C51 drain_right.n16 a_n2224_n2088# 1.4077f
C52 drain_right.n17 a_n2224_n2088# 0.403634f
C53 drain_right.t13 a_n2224_n2088# 0.168788f
C54 drain_right.t1 a_n2224_n2088# 0.168788f
C55 drain_right.n18 a_n2224_n2088# 1.4077f
C56 drain_right.n19 a_n2224_n2088# 0.403634f
C57 drain_right.t6 a_n2224_n2088# 0.168788f
C58 drain_right.t21 a_n2224_n2088# 0.168788f
C59 drain_right.n20 a_n2224_n2088# 1.4077f
C60 drain_right.n21 a_n2224_n2088# 0.697478f
C61 minus.n0 a_n2224_n2088# 0.049762f
C62 minus.t17 a_n2224_n2088# 0.216401f
C63 minus.t2 a_n2224_n2088# 0.212671f
C64 minus.t10 a_n2224_n2088# 0.212671f
C65 minus.n1 a_n2224_n2088# 0.018042f
C66 minus.n2 a_n2224_n2088# 0.049762f
C67 minus.t22 a_n2224_n2088# 0.212671f
C68 minus.n3 a_n2224_n2088# 0.100176f
C69 minus.t5 a_n2224_n2088# 0.212671f
C70 minus.t21 a_n2224_n2088# 0.212671f
C71 minus.t8 a_n2224_n2088# 0.212671f
C72 minus.n4 a_n2224_n2088# 0.100176f
C73 minus.n5 a_n2224_n2088# 0.049762f
C74 minus.t20 a_n2224_n2088# 0.212671f
C75 minus.t0 a_n2224_n2088# 0.212671f
C76 minus.n6 a_n2224_n2088# 0.017428f
C77 minus.t16 a_n2224_n2088# 0.216401f
C78 minus.n7 a_n2224_n2088# 0.113629f
C79 minus.t14 a_n2224_n2088# 0.212671f
C80 minus.n8 a_n2224_n2088# 0.100176f
C81 minus.t1 a_n2224_n2088# 0.212671f
C82 minus.n9 a_n2224_n2088# 0.100176f
C83 minus.n10 a_n2224_n2088# 0.018962f
C84 minus.n11 a_n2224_n2088# 0.103449f
C85 minus.n12 a_n2224_n2088# 0.049762f
C86 minus.n13 a_n2224_n2088# 0.049762f
C87 minus.n14 a_n2224_n2088# 0.018042f
C88 minus.n15 a_n2224_n2088# 0.100176f
C89 minus.n16 a_n2224_n2088# 0.018962f
C90 minus.n17 a_n2224_n2088# 0.100176f
C91 minus.n18 a_n2224_n2088# 0.018962f
C92 minus.n19 a_n2224_n2088# 0.049762f
C93 minus.n20 a_n2224_n2088# 0.049762f
C94 minus.n21 a_n2224_n2088# 0.018962f
C95 minus.n22 a_n2224_n2088# 0.100176f
C96 minus.n23 a_n2224_n2088# 0.018962f
C97 minus.n24 a_n2224_n2088# 0.100176f
C98 minus.n25 a_n2224_n2088# 0.018962f
C99 minus.n26 a_n2224_n2088# 0.049762f
C100 minus.n27 a_n2224_n2088# 0.049762f
C101 minus.n28 a_n2224_n2088# 0.049762f
C102 minus.n29 a_n2224_n2088# 0.017428f
C103 minus.n30 a_n2224_n2088# 0.100176f
C104 minus.n31 a_n2224_n2088# 0.018962f
C105 minus.n32 a_n2224_n2088# 0.100176f
C106 minus.n33 a_n2224_n2088# 0.113566f
C107 minus.n34 a_n2224_n2088# 1.50963f
C108 minus.n35 a_n2224_n2088# 0.049762f
C109 minus.t12 a_n2224_n2088# 0.212671f
C110 minus.t19 a_n2224_n2088# 0.212671f
C111 minus.n36 a_n2224_n2088# 0.018042f
C112 minus.n37 a_n2224_n2088# 0.049762f
C113 minus.t7 a_n2224_n2088# 0.212671f
C114 minus.t9 a_n2224_n2088# 0.212671f
C115 minus.t13 a_n2224_n2088# 0.212671f
C116 minus.n38 a_n2224_n2088# 0.100176f
C117 minus.n39 a_n2224_n2088# 0.049762f
C118 minus.t23 a_n2224_n2088# 0.212671f
C119 minus.t4 a_n2224_n2088# 0.212671f
C120 minus.n40 a_n2224_n2088# 0.017428f
C121 minus.t15 a_n2224_n2088# 0.216401f
C122 minus.n41 a_n2224_n2088# 0.113629f
C123 minus.t18 a_n2224_n2088# 0.212671f
C124 minus.n42 a_n2224_n2088# 0.100176f
C125 minus.t11 a_n2224_n2088# 0.212671f
C126 minus.n43 a_n2224_n2088# 0.100176f
C127 minus.n44 a_n2224_n2088# 0.018962f
C128 minus.n45 a_n2224_n2088# 0.103449f
C129 minus.n46 a_n2224_n2088# 0.049762f
C130 minus.n47 a_n2224_n2088# 0.049762f
C131 minus.n48 a_n2224_n2088# 0.018042f
C132 minus.n49 a_n2224_n2088# 0.100176f
C133 minus.n50 a_n2224_n2088# 0.018962f
C134 minus.n51 a_n2224_n2088# 0.100176f
C135 minus.n52 a_n2224_n2088# 0.018962f
C136 minus.n53 a_n2224_n2088# 0.049762f
C137 minus.n54 a_n2224_n2088# 0.049762f
C138 minus.n55 a_n2224_n2088# 0.018962f
C139 minus.n56 a_n2224_n2088# 0.100176f
C140 minus.n57 a_n2224_n2088# 0.018962f
C141 minus.n58 a_n2224_n2088# 0.100176f
C142 minus.t3 a_n2224_n2088# 0.212671f
C143 minus.n59 a_n2224_n2088# 0.100176f
C144 minus.n60 a_n2224_n2088# 0.018962f
C145 minus.n61 a_n2224_n2088# 0.049762f
C146 minus.n62 a_n2224_n2088# 0.049762f
C147 minus.n63 a_n2224_n2088# 0.049762f
C148 minus.n64 a_n2224_n2088# 0.017428f
C149 minus.n65 a_n2224_n2088# 0.100176f
C150 minus.n66 a_n2224_n2088# 0.018962f
C151 minus.n67 a_n2224_n2088# 0.100176f
C152 minus.t6 a_n2224_n2088# 0.216401f
C153 minus.n68 a_n2224_n2088# 0.113566f
C154 minus.n69 a_n2224_n2088# 0.31737f
C155 minus.n70 a_n2224_n2088# 1.85392f
C156 drain_left.t20 a_n2224_n2088# 0.169127f
C157 drain_left.t16 a_n2224_n2088# 0.169127f
C158 drain_left.n0 a_n2224_n2088# 1.41361f
C159 drain_left.t14 a_n2224_n2088# 0.169127f
C160 drain_left.t11 a_n2224_n2088# 0.169127f
C161 drain_left.n1 a_n2224_n2088# 1.41052f
C162 drain_left.n2 a_n2224_n2088# 0.820176f
C163 drain_left.t0 a_n2224_n2088# 0.169127f
C164 drain_left.t13 a_n2224_n2088# 0.169127f
C165 drain_left.n3 a_n2224_n2088# 1.41052f
C166 drain_left.n4 a_n2224_n2088# 0.373604f
C167 drain_left.t12 a_n2224_n2088# 0.169127f
C168 drain_left.t6 a_n2224_n2088# 0.169127f
C169 drain_left.n5 a_n2224_n2088# 1.41361f
C170 drain_left.t3 a_n2224_n2088# 0.169127f
C171 drain_left.t21 a_n2224_n2088# 0.169127f
C172 drain_left.n6 a_n2224_n2088# 1.41052f
C173 drain_left.n7 a_n2224_n2088# 0.820176f
C174 drain_left.t10 a_n2224_n2088# 0.169127f
C175 drain_left.t2 a_n2224_n2088# 0.169127f
C176 drain_left.n8 a_n2224_n2088# 1.41052f
C177 drain_left.n9 a_n2224_n2088# 0.373604f
C178 drain_left.n10 a_n2224_n2088# 1.41482f
C179 drain_left.t15 a_n2224_n2088# 0.169127f
C180 drain_left.t22 a_n2224_n2088# 0.169127f
C181 drain_left.n11 a_n2224_n2088# 1.41362f
C182 drain_left.t7 a_n2224_n2088# 0.169127f
C183 drain_left.t23 a_n2224_n2088# 0.169127f
C184 drain_left.n12 a_n2224_n2088# 1.41053f
C185 drain_left.n13 a_n2224_n2088# 0.820162f
C186 drain_left.t8 a_n2224_n2088# 0.169127f
C187 drain_left.t1 a_n2224_n2088# 0.169127f
C188 drain_left.n14 a_n2224_n2088# 1.41053f
C189 drain_left.n15 a_n2224_n2088# 0.404444f
C190 drain_left.t9 a_n2224_n2088# 0.169127f
C191 drain_left.t17 a_n2224_n2088# 0.169127f
C192 drain_left.n16 a_n2224_n2088# 1.41053f
C193 drain_left.n17 a_n2224_n2088# 0.404444f
C194 drain_left.t4 a_n2224_n2088# 0.169127f
C195 drain_left.t18 a_n2224_n2088# 0.169127f
C196 drain_left.n18 a_n2224_n2088# 1.41053f
C197 drain_left.n19 a_n2224_n2088# 0.404444f
C198 drain_left.t5 a_n2224_n2088# 0.169127f
C199 drain_left.t19 a_n2224_n2088# 0.169127f
C200 drain_left.n20 a_n2224_n2088# 1.41052f
C201 drain_left.n21 a_n2224_n2088# 0.698886f
C202 source.n0 a_n2224_n2088# 0.046835f
C203 source.n1 a_n2224_n2088# 0.03332f
C204 source.n2 a_n2224_n2088# 0.017905f
C205 source.n3 a_n2224_n2088# 0.042321f
C206 source.n4 a_n2224_n2088# 0.018958f
C207 source.n5 a_n2224_n2088# 0.03332f
C208 source.n6 a_n2224_n2088# 0.017905f
C209 source.n7 a_n2224_n2088# 0.042321f
C210 source.n8 a_n2224_n2088# 0.018958f
C211 source.n9 a_n2224_n2088# 0.142588f
C212 source.t45 a_n2224_n2088# 0.068977f
C213 source.n10 a_n2224_n2088# 0.03174f
C214 source.n11 a_n2224_n2088# 0.024998f
C215 source.n12 a_n2224_n2088# 0.017905f
C216 source.n13 a_n2224_n2088# 0.792825f
C217 source.n14 a_n2224_n2088# 0.03332f
C218 source.n15 a_n2224_n2088# 0.017905f
C219 source.n16 a_n2224_n2088# 0.018958f
C220 source.n17 a_n2224_n2088# 0.042321f
C221 source.n18 a_n2224_n2088# 0.042321f
C222 source.n19 a_n2224_n2088# 0.018958f
C223 source.n20 a_n2224_n2088# 0.017905f
C224 source.n21 a_n2224_n2088# 0.03332f
C225 source.n22 a_n2224_n2088# 0.03332f
C226 source.n23 a_n2224_n2088# 0.017905f
C227 source.n24 a_n2224_n2088# 0.018958f
C228 source.n25 a_n2224_n2088# 0.042321f
C229 source.n26 a_n2224_n2088# 0.091617f
C230 source.n27 a_n2224_n2088# 0.018958f
C231 source.n28 a_n2224_n2088# 0.017905f
C232 source.n29 a_n2224_n2088# 0.077018f
C233 source.n30 a_n2224_n2088# 0.051263f
C234 source.n31 a_n2224_n2088# 0.799148f
C235 source.t41 a_n2224_n2088# 0.157984f
C236 source.t31 a_n2224_n2088# 0.157984f
C237 source.n32 a_n2224_n2088# 1.23039f
C238 source.n33 a_n2224_n2088# 0.419711f
C239 source.t42 a_n2224_n2088# 0.157984f
C240 source.t47 a_n2224_n2088# 0.157984f
C241 source.n34 a_n2224_n2088# 1.23039f
C242 source.n35 a_n2224_n2088# 0.419711f
C243 source.t36 a_n2224_n2088# 0.157984f
C244 source.t30 a_n2224_n2088# 0.157984f
C245 source.n36 a_n2224_n2088# 1.23039f
C246 source.n37 a_n2224_n2088# 0.419711f
C247 source.t38 a_n2224_n2088# 0.157984f
C248 source.t33 a_n2224_n2088# 0.157984f
C249 source.n38 a_n2224_n2088# 1.23039f
C250 source.n39 a_n2224_n2088# 0.419711f
C251 source.t24 a_n2224_n2088# 0.157984f
C252 source.t27 a_n2224_n2088# 0.157984f
C253 source.n40 a_n2224_n2088# 1.23039f
C254 source.n41 a_n2224_n2088# 0.419711f
C255 source.n42 a_n2224_n2088# 0.046835f
C256 source.n43 a_n2224_n2088# 0.03332f
C257 source.n44 a_n2224_n2088# 0.017905f
C258 source.n45 a_n2224_n2088# 0.042321f
C259 source.n46 a_n2224_n2088# 0.018958f
C260 source.n47 a_n2224_n2088# 0.03332f
C261 source.n48 a_n2224_n2088# 0.017905f
C262 source.n49 a_n2224_n2088# 0.042321f
C263 source.n50 a_n2224_n2088# 0.018958f
C264 source.n51 a_n2224_n2088# 0.142588f
C265 source.t25 a_n2224_n2088# 0.068977f
C266 source.n52 a_n2224_n2088# 0.03174f
C267 source.n53 a_n2224_n2088# 0.024998f
C268 source.n54 a_n2224_n2088# 0.017905f
C269 source.n55 a_n2224_n2088# 0.792825f
C270 source.n56 a_n2224_n2088# 0.03332f
C271 source.n57 a_n2224_n2088# 0.017905f
C272 source.n58 a_n2224_n2088# 0.018958f
C273 source.n59 a_n2224_n2088# 0.042321f
C274 source.n60 a_n2224_n2088# 0.042321f
C275 source.n61 a_n2224_n2088# 0.018958f
C276 source.n62 a_n2224_n2088# 0.017905f
C277 source.n63 a_n2224_n2088# 0.03332f
C278 source.n64 a_n2224_n2088# 0.03332f
C279 source.n65 a_n2224_n2088# 0.017905f
C280 source.n66 a_n2224_n2088# 0.018958f
C281 source.n67 a_n2224_n2088# 0.042321f
C282 source.n68 a_n2224_n2088# 0.091617f
C283 source.n69 a_n2224_n2088# 0.018958f
C284 source.n70 a_n2224_n2088# 0.017905f
C285 source.n71 a_n2224_n2088# 0.077018f
C286 source.n72 a_n2224_n2088# 0.051263f
C287 source.n73 a_n2224_n2088# 0.132584f
C288 source.n74 a_n2224_n2088# 0.046835f
C289 source.n75 a_n2224_n2088# 0.03332f
C290 source.n76 a_n2224_n2088# 0.017905f
C291 source.n77 a_n2224_n2088# 0.042321f
C292 source.n78 a_n2224_n2088# 0.018958f
C293 source.n79 a_n2224_n2088# 0.03332f
C294 source.n80 a_n2224_n2088# 0.017905f
C295 source.n81 a_n2224_n2088# 0.042321f
C296 source.n82 a_n2224_n2088# 0.018958f
C297 source.n83 a_n2224_n2088# 0.142588f
C298 source.t19 a_n2224_n2088# 0.068977f
C299 source.n84 a_n2224_n2088# 0.03174f
C300 source.n85 a_n2224_n2088# 0.024998f
C301 source.n86 a_n2224_n2088# 0.017905f
C302 source.n87 a_n2224_n2088# 0.792825f
C303 source.n88 a_n2224_n2088# 0.03332f
C304 source.n89 a_n2224_n2088# 0.017905f
C305 source.n90 a_n2224_n2088# 0.018958f
C306 source.n91 a_n2224_n2088# 0.042321f
C307 source.n92 a_n2224_n2088# 0.042321f
C308 source.n93 a_n2224_n2088# 0.018958f
C309 source.n94 a_n2224_n2088# 0.017905f
C310 source.n95 a_n2224_n2088# 0.03332f
C311 source.n96 a_n2224_n2088# 0.03332f
C312 source.n97 a_n2224_n2088# 0.017905f
C313 source.n98 a_n2224_n2088# 0.018958f
C314 source.n99 a_n2224_n2088# 0.042321f
C315 source.n100 a_n2224_n2088# 0.091617f
C316 source.n101 a_n2224_n2088# 0.018958f
C317 source.n102 a_n2224_n2088# 0.017905f
C318 source.n103 a_n2224_n2088# 0.077018f
C319 source.n104 a_n2224_n2088# 0.051263f
C320 source.n105 a_n2224_n2088# 0.132584f
C321 source.t8 a_n2224_n2088# 0.157984f
C322 source.t15 a_n2224_n2088# 0.157984f
C323 source.n106 a_n2224_n2088# 1.23039f
C324 source.n107 a_n2224_n2088# 0.419711f
C325 source.t13 a_n2224_n2088# 0.157984f
C326 source.t11 a_n2224_n2088# 0.157984f
C327 source.n108 a_n2224_n2088# 1.23039f
C328 source.n109 a_n2224_n2088# 0.419711f
C329 source.t5 a_n2224_n2088# 0.157984f
C330 source.t17 a_n2224_n2088# 0.157984f
C331 source.n110 a_n2224_n2088# 1.23039f
C332 source.n111 a_n2224_n2088# 0.419711f
C333 source.t3 a_n2224_n2088# 0.157984f
C334 source.t2 a_n2224_n2088# 0.157984f
C335 source.n112 a_n2224_n2088# 1.23039f
C336 source.n113 a_n2224_n2088# 0.419711f
C337 source.t0 a_n2224_n2088# 0.157984f
C338 source.t20 a_n2224_n2088# 0.157984f
C339 source.n114 a_n2224_n2088# 1.23039f
C340 source.n115 a_n2224_n2088# 0.419711f
C341 source.n116 a_n2224_n2088# 0.046835f
C342 source.n117 a_n2224_n2088# 0.03332f
C343 source.n118 a_n2224_n2088# 0.017905f
C344 source.n119 a_n2224_n2088# 0.042321f
C345 source.n120 a_n2224_n2088# 0.018958f
C346 source.n121 a_n2224_n2088# 0.03332f
C347 source.n122 a_n2224_n2088# 0.017905f
C348 source.n123 a_n2224_n2088# 0.042321f
C349 source.n124 a_n2224_n2088# 0.018958f
C350 source.n125 a_n2224_n2088# 0.142588f
C351 source.t22 a_n2224_n2088# 0.068977f
C352 source.n126 a_n2224_n2088# 0.03174f
C353 source.n127 a_n2224_n2088# 0.024998f
C354 source.n128 a_n2224_n2088# 0.017905f
C355 source.n129 a_n2224_n2088# 0.792825f
C356 source.n130 a_n2224_n2088# 0.03332f
C357 source.n131 a_n2224_n2088# 0.017905f
C358 source.n132 a_n2224_n2088# 0.018958f
C359 source.n133 a_n2224_n2088# 0.042321f
C360 source.n134 a_n2224_n2088# 0.042321f
C361 source.n135 a_n2224_n2088# 0.018958f
C362 source.n136 a_n2224_n2088# 0.017905f
C363 source.n137 a_n2224_n2088# 0.03332f
C364 source.n138 a_n2224_n2088# 0.03332f
C365 source.n139 a_n2224_n2088# 0.017905f
C366 source.n140 a_n2224_n2088# 0.018958f
C367 source.n141 a_n2224_n2088# 0.042321f
C368 source.n142 a_n2224_n2088# 0.091617f
C369 source.n143 a_n2224_n2088# 0.018958f
C370 source.n144 a_n2224_n2088# 0.017905f
C371 source.n145 a_n2224_n2088# 0.077018f
C372 source.n146 a_n2224_n2088# 0.051263f
C373 source.n147 a_n2224_n2088# 1.22679f
C374 source.n148 a_n2224_n2088# 0.046835f
C375 source.n149 a_n2224_n2088# 0.03332f
C376 source.n150 a_n2224_n2088# 0.017905f
C377 source.n151 a_n2224_n2088# 0.042321f
C378 source.n152 a_n2224_n2088# 0.018958f
C379 source.n153 a_n2224_n2088# 0.03332f
C380 source.n154 a_n2224_n2088# 0.017905f
C381 source.n155 a_n2224_n2088# 0.042321f
C382 source.n156 a_n2224_n2088# 0.018958f
C383 source.n157 a_n2224_n2088# 0.142588f
C384 source.t43 a_n2224_n2088# 0.068977f
C385 source.n158 a_n2224_n2088# 0.03174f
C386 source.n159 a_n2224_n2088# 0.024998f
C387 source.n160 a_n2224_n2088# 0.017905f
C388 source.n161 a_n2224_n2088# 0.792825f
C389 source.n162 a_n2224_n2088# 0.03332f
C390 source.n163 a_n2224_n2088# 0.017905f
C391 source.n164 a_n2224_n2088# 0.018958f
C392 source.n165 a_n2224_n2088# 0.042321f
C393 source.n166 a_n2224_n2088# 0.042321f
C394 source.n167 a_n2224_n2088# 0.018958f
C395 source.n168 a_n2224_n2088# 0.017905f
C396 source.n169 a_n2224_n2088# 0.03332f
C397 source.n170 a_n2224_n2088# 0.03332f
C398 source.n171 a_n2224_n2088# 0.017905f
C399 source.n172 a_n2224_n2088# 0.018958f
C400 source.n173 a_n2224_n2088# 0.042321f
C401 source.n174 a_n2224_n2088# 0.091617f
C402 source.n175 a_n2224_n2088# 0.018958f
C403 source.n176 a_n2224_n2088# 0.017905f
C404 source.n177 a_n2224_n2088# 0.077018f
C405 source.n178 a_n2224_n2088# 0.051263f
C406 source.n179 a_n2224_n2088# 1.22679f
C407 source.t44 a_n2224_n2088# 0.157984f
C408 source.t29 a_n2224_n2088# 0.157984f
C409 source.n180 a_n2224_n2088# 1.23039f
C410 source.n181 a_n2224_n2088# 0.41972f
C411 source.t32 a_n2224_n2088# 0.157984f
C412 source.t37 a_n2224_n2088# 0.157984f
C413 source.n182 a_n2224_n2088# 1.23039f
C414 source.n183 a_n2224_n2088# 0.41972f
C415 source.t28 a_n2224_n2088# 0.157984f
C416 source.t26 a_n2224_n2088# 0.157984f
C417 source.n184 a_n2224_n2088# 1.23039f
C418 source.n185 a_n2224_n2088# 0.41972f
C419 source.t35 a_n2224_n2088# 0.157984f
C420 source.t34 a_n2224_n2088# 0.157984f
C421 source.n186 a_n2224_n2088# 1.23039f
C422 source.n187 a_n2224_n2088# 0.41972f
C423 source.t39 a_n2224_n2088# 0.157984f
C424 source.t46 a_n2224_n2088# 0.157984f
C425 source.n188 a_n2224_n2088# 1.23039f
C426 source.n189 a_n2224_n2088# 0.41972f
C427 source.n190 a_n2224_n2088# 0.046835f
C428 source.n191 a_n2224_n2088# 0.03332f
C429 source.n192 a_n2224_n2088# 0.017905f
C430 source.n193 a_n2224_n2088# 0.042321f
C431 source.n194 a_n2224_n2088# 0.018958f
C432 source.n195 a_n2224_n2088# 0.03332f
C433 source.n196 a_n2224_n2088# 0.017905f
C434 source.n197 a_n2224_n2088# 0.042321f
C435 source.n198 a_n2224_n2088# 0.018958f
C436 source.n199 a_n2224_n2088# 0.142588f
C437 source.t40 a_n2224_n2088# 0.068977f
C438 source.n200 a_n2224_n2088# 0.03174f
C439 source.n201 a_n2224_n2088# 0.024998f
C440 source.n202 a_n2224_n2088# 0.017905f
C441 source.n203 a_n2224_n2088# 0.792825f
C442 source.n204 a_n2224_n2088# 0.03332f
C443 source.n205 a_n2224_n2088# 0.017905f
C444 source.n206 a_n2224_n2088# 0.018958f
C445 source.n207 a_n2224_n2088# 0.042321f
C446 source.n208 a_n2224_n2088# 0.042321f
C447 source.n209 a_n2224_n2088# 0.018958f
C448 source.n210 a_n2224_n2088# 0.017905f
C449 source.n211 a_n2224_n2088# 0.03332f
C450 source.n212 a_n2224_n2088# 0.03332f
C451 source.n213 a_n2224_n2088# 0.017905f
C452 source.n214 a_n2224_n2088# 0.018958f
C453 source.n215 a_n2224_n2088# 0.042321f
C454 source.n216 a_n2224_n2088# 0.091617f
C455 source.n217 a_n2224_n2088# 0.018958f
C456 source.n218 a_n2224_n2088# 0.017905f
C457 source.n219 a_n2224_n2088# 0.077018f
C458 source.n220 a_n2224_n2088# 0.051263f
C459 source.n221 a_n2224_n2088# 0.132584f
C460 source.n222 a_n2224_n2088# 0.046835f
C461 source.n223 a_n2224_n2088# 0.03332f
C462 source.n224 a_n2224_n2088# 0.017905f
C463 source.n225 a_n2224_n2088# 0.042321f
C464 source.n226 a_n2224_n2088# 0.018958f
C465 source.n227 a_n2224_n2088# 0.03332f
C466 source.n228 a_n2224_n2088# 0.017905f
C467 source.n229 a_n2224_n2088# 0.042321f
C468 source.n230 a_n2224_n2088# 0.018958f
C469 source.n231 a_n2224_n2088# 0.142588f
C470 source.t14 a_n2224_n2088# 0.068977f
C471 source.n232 a_n2224_n2088# 0.03174f
C472 source.n233 a_n2224_n2088# 0.024998f
C473 source.n234 a_n2224_n2088# 0.017905f
C474 source.n235 a_n2224_n2088# 0.792825f
C475 source.n236 a_n2224_n2088# 0.03332f
C476 source.n237 a_n2224_n2088# 0.017905f
C477 source.n238 a_n2224_n2088# 0.018958f
C478 source.n239 a_n2224_n2088# 0.042321f
C479 source.n240 a_n2224_n2088# 0.042321f
C480 source.n241 a_n2224_n2088# 0.018958f
C481 source.n242 a_n2224_n2088# 0.017905f
C482 source.n243 a_n2224_n2088# 0.03332f
C483 source.n244 a_n2224_n2088# 0.03332f
C484 source.n245 a_n2224_n2088# 0.017905f
C485 source.n246 a_n2224_n2088# 0.018958f
C486 source.n247 a_n2224_n2088# 0.042321f
C487 source.n248 a_n2224_n2088# 0.091617f
C488 source.n249 a_n2224_n2088# 0.018958f
C489 source.n250 a_n2224_n2088# 0.017905f
C490 source.n251 a_n2224_n2088# 0.077018f
C491 source.n252 a_n2224_n2088# 0.051263f
C492 source.n253 a_n2224_n2088# 0.132584f
C493 source.t4 a_n2224_n2088# 0.157984f
C494 source.t23 a_n2224_n2088# 0.157984f
C495 source.n254 a_n2224_n2088# 1.23039f
C496 source.n255 a_n2224_n2088# 0.41972f
C497 source.t7 a_n2224_n2088# 0.157984f
C498 source.t6 a_n2224_n2088# 0.157984f
C499 source.n256 a_n2224_n2088# 1.23039f
C500 source.n257 a_n2224_n2088# 0.41972f
C501 source.t18 a_n2224_n2088# 0.157984f
C502 source.t9 a_n2224_n2088# 0.157984f
C503 source.n258 a_n2224_n2088# 1.23039f
C504 source.n259 a_n2224_n2088# 0.41972f
C505 source.t12 a_n2224_n2088# 0.157984f
C506 source.t1 a_n2224_n2088# 0.157984f
C507 source.n260 a_n2224_n2088# 1.23039f
C508 source.n261 a_n2224_n2088# 0.41972f
C509 source.t10 a_n2224_n2088# 0.157984f
C510 source.t16 a_n2224_n2088# 0.157984f
C511 source.n262 a_n2224_n2088# 1.23039f
C512 source.n263 a_n2224_n2088# 0.41972f
C513 source.n264 a_n2224_n2088# 0.046835f
C514 source.n265 a_n2224_n2088# 0.03332f
C515 source.n266 a_n2224_n2088# 0.017905f
C516 source.n267 a_n2224_n2088# 0.042321f
C517 source.n268 a_n2224_n2088# 0.018958f
C518 source.n269 a_n2224_n2088# 0.03332f
C519 source.n270 a_n2224_n2088# 0.017905f
C520 source.n271 a_n2224_n2088# 0.042321f
C521 source.n272 a_n2224_n2088# 0.018958f
C522 source.n273 a_n2224_n2088# 0.142588f
C523 source.t21 a_n2224_n2088# 0.068977f
C524 source.n274 a_n2224_n2088# 0.03174f
C525 source.n275 a_n2224_n2088# 0.024998f
C526 source.n276 a_n2224_n2088# 0.017905f
C527 source.n277 a_n2224_n2088# 0.792825f
C528 source.n278 a_n2224_n2088# 0.03332f
C529 source.n279 a_n2224_n2088# 0.017905f
C530 source.n280 a_n2224_n2088# 0.018958f
C531 source.n281 a_n2224_n2088# 0.042321f
C532 source.n282 a_n2224_n2088# 0.042321f
C533 source.n283 a_n2224_n2088# 0.018958f
C534 source.n284 a_n2224_n2088# 0.017905f
C535 source.n285 a_n2224_n2088# 0.03332f
C536 source.n286 a_n2224_n2088# 0.03332f
C537 source.n287 a_n2224_n2088# 0.017905f
C538 source.n288 a_n2224_n2088# 0.018958f
C539 source.n289 a_n2224_n2088# 0.042321f
C540 source.n290 a_n2224_n2088# 0.091617f
C541 source.n291 a_n2224_n2088# 0.018958f
C542 source.n292 a_n2224_n2088# 0.017905f
C543 source.n293 a_n2224_n2088# 0.077018f
C544 source.n294 a_n2224_n2088# 0.051263f
C545 source.n295 a_n2224_n2088# 0.316972f
C546 source.n296 a_n2224_n2088# 1.36117f
C547 plus.n0 a_n2224_n2088# 0.050931f
C548 plus.t18 a_n2224_n2088# 0.217666f
C549 plus.t5 a_n2224_n2088# 0.217666f
C550 plus.n1 a_n2224_n2088# 0.018465f
C551 plus.n2 a_n2224_n2088# 0.050931f
C552 plus.t6 a_n2224_n2088# 0.217666f
C553 plus.t14 a_n2224_n2088# 0.217666f
C554 plus.t22 a_n2224_n2088# 0.217666f
C555 plus.n3 a_n2224_n2088# 0.102529f
C556 plus.n4 a_n2224_n2088# 0.050931f
C557 plus.t15 a_n2224_n2088# 0.217666f
C558 plus.t0 a_n2224_n2088# 0.217666f
C559 plus.n5 a_n2224_n2088# 0.017837f
C560 plus.t8 a_n2224_n2088# 0.221484f
C561 plus.n6 a_n2224_n2088# 0.116298f
C562 plus.t1 a_n2224_n2088# 0.217666f
C563 plus.n7 a_n2224_n2088# 0.102529f
C564 plus.t16 a_n2224_n2088# 0.217666f
C565 plus.n8 a_n2224_n2088# 0.102529f
C566 plus.n9 a_n2224_n2088# 0.019407f
C567 plus.n10 a_n2224_n2088# 0.105879f
C568 plus.n11 a_n2224_n2088# 0.050931f
C569 plus.n12 a_n2224_n2088# 0.050931f
C570 plus.n13 a_n2224_n2088# 0.018465f
C571 plus.n14 a_n2224_n2088# 0.102529f
C572 plus.n15 a_n2224_n2088# 0.019407f
C573 plus.n16 a_n2224_n2088# 0.102529f
C574 plus.n17 a_n2224_n2088# 0.019407f
C575 plus.n18 a_n2224_n2088# 0.050931f
C576 plus.n19 a_n2224_n2088# 0.050931f
C577 plus.n20 a_n2224_n2088# 0.019407f
C578 plus.n21 a_n2224_n2088# 0.102529f
C579 plus.n22 a_n2224_n2088# 0.019407f
C580 plus.n23 a_n2224_n2088# 0.102529f
C581 plus.t19 a_n2224_n2088# 0.217666f
C582 plus.n24 a_n2224_n2088# 0.102529f
C583 plus.n25 a_n2224_n2088# 0.019407f
C584 plus.n26 a_n2224_n2088# 0.050931f
C585 plus.n27 a_n2224_n2088# 0.050931f
C586 plus.n28 a_n2224_n2088# 0.050931f
C587 plus.n29 a_n2224_n2088# 0.017837f
C588 plus.n30 a_n2224_n2088# 0.102529f
C589 plus.n31 a_n2224_n2088# 0.019407f
C590 plus.n32 a_n2224_n2088# 0.102529f
C591 plus.t4 a_n2224_n2088# 0.221484f
C592 plus.n33 a_n2224_n2088# 0.116234f
C593 plus.n34 a_n2224_n2088# 0.427932f
C594 plus.n35 a_n2224_n2088# 0.050931f
C595 plus.t3 a_n2224_n2088# 0.221484f
C596 plus.t7 a_n2224_n2088# 0.217666f
C597 plus.t9 a_n2224_n2088# 0.217666f
C598 plus.n36 a_n2224_n2088# 0.018465f
C599 plus.n37 a_n2224_n2088# 0.050931f
C600 plus.t12 a_n2224_n2088# 0.217666f
C601 plus.n38 a_n2224_n2088# 0.102529f
C602 plus.t23 a_n2224_n2088# 0.217666f
C603 plus.t10 a_n2224_n2088# 0.217666f
C604 plus.t13 a_n2224_n2088# 0.217666f
C605 plus.n39 a_n2224_n2088# 0.102529f
C606 plus.n40 a_n2224_n2088# 0.050931f
C607 plus.t21 a_n2224_n2088# 0.217666f
C608 plus.t20 a_n2224_n2088# 0.217666f
C609 plus.n41 a_n2224_n2088# 0.017837f
C610 plus.t17 a_n2224_n2088# 0.221484f
C611 plus.n42 a_n2224_n2088# 0.116298f
C612 plus.t2 a_n2224_n2088# 0.217666f
C613 plus.n43 a_n2224_n2088# 0.102529f
C614 plus.t11 a_n2224_n2088# 0.217666f
C615 plus.n44 a_n2224_n2088# 0.102529f
C616 plus.n45 a_n2224_n2088# 0.019407f
C617 plus.n46 a_n2224_n2088# 0.105879f
C618 plus.n47 a_n2224_n2088# 0.050931f
C619 plus.n48 a_n2224_n2088# 0.050931f
C620 plus.n49 a_n2224_n2088# 0.018465f
C621 plus.n50 a_n2224_n2088# 0.102529f
C622 plus.n51 a_n2224_n2088# 0.019407f
C623 plus.n52 a_n2224_n2088# 0.102529f
C624 plus.n53 a_n2224_n2088# 0.019407f
C625 plus.n54 a_n2224_n2088# 0.050931f
C626 plus.n55 a_n2224_n2088# 0.050931f
C627 plus.n56 a_n2224_n2088# 0.019407f
C628 plus.n57 a_n2224_n2088# 0.102529f
C629 plus.n58 a_n2224_n2088# 0.019407f
C630 plus.n59 a_n2224_n2088# 0.102529f
C631 plus.n60 a_n2224_n2088# 0.019407f
C632 plus.n61 a_n2224_n2088# 0.050931f
C633 plus.n62 a_n2224_n2088# 0.050931f
C634 plus.n63 a_n2224_n2088# 0.050931f
C635 plus.n64 a_n2224_n2088# 0.017837f
C636 plus.n65 a_n2224_n2088# 0.102529f
C637 plus.n66 a_n2224_n2088# 0.019407f
C638 plus.n67 a_n2224_n2088# 0.102529f
C639 plus.n68 a_n2224_n2088# 0.116234f
C640 plus.n69 a_n2224_n2088# 1.39556f
.ends

