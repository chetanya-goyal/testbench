* NGSPICE file created from diffpair251.ext - technology: sky130A

.subckt diffpair251 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t7 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X1 source.t0 plus.t0 drain_left.t3 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X2 a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X3 a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X4 source.t6 minus.t1 drain_right.t2 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X5 drain_right.t1 minus.t2 source.t5 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X6 a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X7 drain_left.t2 plus.t1 source.t1 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X8 source.t4 minus.t3 drain_right.t0 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X9 a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X10 source.t3 plus.t2 drain_left.t1 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X11 drain_left.t0 plus.t3 source.t2 a_n1034_n2092# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
R0 minus.n0 minus.t3 918.356
R1 minus.n0 minus.t0 918.356
R2 minus.n1 minus.t2 918.356
R3 minus.n1 minus.t1 918.356
R4 minus.n2 minus.n0 189.739
R5 minus.n2 minus.n1 167.732
R6 minus minus.n2 0.188
R7 source.n250 source.n224 289.615
R8 source.n218 source.n192 289.615
R9 source.n186 source.n160 289.615
R10 source.n154 source.n128 289.615
R11 source.n26 source.n0 289.615
R12 source.n58 source.n32 289.615
R13 source.n90 source.n64 289.615
R14 source.n122 source.n96 289.615
R15 source.n235 source.n234 185
R16 source.n232 source.n231 185
R17 source.n241 source.n240 185
R18 source.n243 source.n242 185
R19 source.n228 source.n227 185
R20 source.n249 source.n248 185
R21 source.n251 source.n250 185
R22 source.n203 source.n202 185
R23 source.n200 source.n199 185
R24 source.n209 source.n208 185
R25 source.n211 source.n210 185
R26 source.n196 source.n195 185
R27 source.n217 source.n216 185
R28 source.n219 source.n218 185
R29 source.n171 source.n170 185
R30 source.n168 source.n167 185
R31 source.n177 source.n176 185
R32 source.n179 source.n178 185
R33 source.n164 source.n163 185
R34 source.n185 source.n184 185
R35 source.n187 source.n186 185
R36 source.n139 source.n138 185
R37 source.n136 source.n135 185
R38 source.n145 source.n144 185
R39 source.n147 source.n146 185
R40 source.n132 source.n131 185
R41 source.n153 source.n152 185
R42 source.n155 source.n154 185
R43 source.n27 source.n26 185
R44 source.n25 source.n24 185
R45 source.n4 source.n3 185
R46 source.n19 source.n18 185
R47 source.n17 source.n16 185
R48 source.n8 source.n7 185
R49 source.n11 source.n10 185
R50 source.n59 source.n58 185
R51 source.n57 source.n56 185
R52 source.n36 source.n35 185
R53 source.n51 source.n50 185
R54 source.n49 source.n48 185
R55 source.n40 source.n39 185
R56 source.n43 source.n42 185
R57 source.n91 source.n90 185
R58 source.n89 source.n88 185
R59 source.n68 source.n67 185
R60 source.n83 source.n82 185
R61 source.n81 source.n80 185
R62 source.n72 source.n71 185
R63 source.n75 source.n74 185
R64 source.n123 source.n122 185
R65 source.n121 source.n120 185
R66 source.n100 source.n99 185
R67 source.n115 source.n114 185
R68 source.n113 source.n112 185
R69 source.n104 source.n103 185
R70 source.n107 source.n106 185
R71 source.t5 source.n233 147.661
R72 source.t6 source.n201 147.661
R73 source.t2 source.n169 147.661
R74 source.t0 source.n137 147.661
R75 source.t1 source.n9 147.661
R76 source.t3 source.n41 147.661
R77 source.t7 source.n73 147.661
R78 source.t4 source.n105 147.661
R79 source.n234 source.n231 104.615
R80 source.n241 source.n231 104.615
R81 source.n242 source.n241 104.615
R82 source.n242 source.n227 104.615
R83 source.n249 source.n227 104.615
R84 source.n250 source.n249 104.615
R85 source.n202 source.n199 104.615
R86 source.n209 source.n199 104.615
R87 source.n210 source.n209 104.615
R88 source.n210 source.n195 104.615
R89 source.n217 source.n195 104.615
R90 source.n218 source.n217 104.615
R91 source.n170 source.n167 104.615
R92 source.n177 source.n167 104.615
R93 source.n178 source.n177 104.615
R94 source.n178 source.n163 104.615
R95 source.n185 source.n163 104.615
R96 source.n186 source.n185 104.615
R97 source.n138 source.n135 104.615
R98 source.n145 source.n135 104.615
R99 source.n146 source.n145 104.615
R100 source.n146 source.n131 104.615
R101 source.n153 source.n131 104.615
R102 source.n154 source.n153 104.615
R103 source.n26 source.n25 104.615
R104 source.n25 source.n3 104.615
R105 source.n18 source.n3 104.615
R106 source.n18 source.n17 104.615
R107 source.n17 source.n7 104.615
R108 source.n10 source.n7 104.615
R109 source.n58 source.n57 104.615
R110 source.n57 source.n35 104.615
R111 source.n50 source.n35 104.615
R112 source.n50 source.n49 104.615
R113 source.n49 source.n39 104.615
R114 source.n42 source.n39 104.615
R115 source.n90 source.n89 104.615
R116 source.n89 source.n67 104.615
R117 source.n82 source.n67 104.615
R118 source.n82 source.n81 104.615
R119 source.n81 source.n71 104.615
R120 source.n74 source.n71 104.615
R121 source.n122 source.n121 104.615
R122 source.n121 source.n99 104.615
R123 source.n114 source.n99 104.615
R124 source.n114 source.n113 104.615
R125 source.n113 source.n103 104.615
R126 source.n106 source.n103 104.615
R127 source.n234 source.t5 52.3082
R128 source.n202 source.t6 52.3082
R129 source.n170 source.t2 52.3082
R130 source.n138 source.t0 52.3082
R131 source.n10 source.t1 52.3082
R132 source.n42 source.t3 52.3082
R133 source.n74 source.t7 52.3082
R134 source.n106 source.t4 52.3082
R135 source.n255 source.n254 32.1853
R136 source.n223 source.n222 32.1853
R137 source.n191 source.n190 32.1853
R138 source.n159 source.n158 32.1853
R139 source.n31 source.n30 32.1853
R140 source.n63 source.n62 32.1853
R141 source.n95 source.n94 32.1853
R142 source.n127 source.n126 32.1853
R143 source.n159 source.n127 17.2143
R144 source.n235 source.n233 15.6674
R145 source.n203 source.n201 15.6674
R146 source.n171 source.n169 15.6674
R147 source.n139 source.n137 15.6674
R148 source.n11 source.n9 15.6674
R149 source.n43 source.n41 15.6674
R150 source.n75 source.n73 15.6674
R151 source.n107 source.n105 15.6674
R152 source.n236 source.n232 12.8005
R153 source.n204 source.n200 12.8005
R154 source.n172 source.n168 12.8005
R155 source.n140 source.n136 12.8005
R156 source.n12 source.n8 12.8005
R157 source.n44 source.n40 12.8005
R158 source.n76 source.n72 12.8005
R159 source.n108 source.n104 12.8005
R160 source.n240 source.n239 12.0247
R161 source.n208 source.n207 12.0247
R162 source.n176 source.n175 12.0247
R163 source.n144 source.n143 12.0247
R164 source.n16 source.n15 12.0247
R165 source.n48 source.n47 12.0247
R166 source.n80 source.n79 12.0247
R167 source.n112 source.n111 12.0247
R168 source.n256 source.n31 11.7229
R169 source.n243 source.n230 11.249
R170 source.n211 source.n198 11.249
R171 source.n179 source.n166 11.249
R172 source.n147 source.n134 11.249
R173 source.n19 source.n6 11.249
R174 source.n51 source.n38 11.249
R175 source.n83 source.n70 11.249
R176 source.n115 source.n102 11.249
R177 source.n244 source.n228 10.4732
R178 source.n212 source.n196 10.4732
R179 source.n180 source.n164 10.4732
R180 source.n148 source.n132 10.4732
R181 source.n20 source.n4 10.4732
R182 source.n52 source.n36 10.4732
R183 source.n84 source.n68 10.4732
R184 source.n116 source.n100 10.4732
R185 source.n248 source.n247 9.69747
R186 source.n216 source.n215 9.69747
R187 source.n184 source.n183 9.69747
R188 source.n152 source.n151 9.69747
R189 source.n24 source.n23 9.69747
R190 source.n56 source.n55 9.69747
R191 source.n88 source.n87 9.69747
R192 source.n120 source.n119 9.69747
R193 source.n254 source.n253 9.45567
R194 source.n222 source.n221 9.45567
R195 source.n190 source.n189 9.45567
R196 source.n158 source.n157 9.45567
R197 source.n30 source.n29 9.45567
R198 source.n62 source.n61 9.45567
R199 source.n94 source.n93 9.45567
R200 source.n126 source.n125 9.45567
R201 source.n253 source.n252 9.3005
R202 source.n226 source.n225 9.3005
R203 source.n247 source.n246 9.3005
R204 source.n245 source.n244 9.3005
R205 source.n230 source.n229 9.3005
R206 source.n239 source.n238 9.3005
R207 source.n237 source.n236 9.3005
R208 source.n221 source.n220 9.3005
R209 source.n194 source.n193 9.3005
R210 source.n215 source.n214 9.3005
R211 source.n213 source.n212 9.3005
R212 source.n198 source.n197 9.3005
R213 source.n207 source.n206 9.3005
R214 source.n205 source.n204 9.3005
R215 source.n189 source.n188 9.3005
R216 source.n162 source.n161 9.3005
R217 source.n183 source.n182 9.3005
R218 source.n181 source.n180 9.3005
R219 source.n166 source.n165 9.3005
R220 source.n175 source.n174 9.3005
R221 source.n173 source.n172 9.3005
R222 source.n157 source.n156 9.3005
R223 source.n130 source.n129 9.3005
R224 source.n151 source.n150 9.3005
R225 source.n149 source.n148 9.3005
R226 source.n134 source.n133 9.3005
R227 source.n143 source.n142 9.3005
R228 source.n141 source.n140 9.3005
R229 source.n29 source.n28 9.3005
R230 source.n2 source.n1 9.3005
R231 source.n23 source.n22 9.3005
R232 source.n21 source.n20 9.3005
R233 source.n6 source.n5 9.3005
R234 source.n15 source.n14 9.3005
R235 source.n13 source.n12 9.3005
R236 source.n61 source.n60 9.3005
R237 source.n34 source.n33 9.3005
R238 source.n55 source.n54 9.3005
R239 source.n53 source.n52 9.3005
R240 source.n38 source.n37 9.3005
R241 source.n47 source.n46 9.3005
R242 source.n45 source.n44 9.3005
R243 source.n93 source.n92 9.3005
R244 source.n66 source.n65 9.3005
R245 source.n87 source.n86 9.3005
R246 source.n85 source.n84 9.3005
R247 source.n70 source.n69 9.3005
R248 source.n79 source.n78 9.3005
R249 source.n77 source.n76 9.3005
R250 source.n125 source.n124 9.3005
R251 source.n98 source.n97 9.3005
R252 source.n119 source.n118 9.3005
R253 source.n117 source.n116 9.3005
R254 source.n102 source.n101 9.3005
R255 source.n111 source.n110 9.3005
R256 source.n109 source.n108 9.3005
R257 source.n251 source.n226 8.92171
R258 source.n219 source.n194 8.92171
R259 source.n187 source.n162 8.92171
R260 source.n155 source.n130 8.92171
R261 source.n27 source.n2 8.92171
R262 source.n59 source.n34 8.92171
R263 source.n91 source.n66 8.92171
R264 source.n123 source.n98 8.92171
R265 source.n252 source.n224 8.14595
R266 source.n220 source.n192 8.14595
R267 source.n188 source.n160 8.14595
R268 source.n156 source.n128 8.14595
R269 source.n28 source.n0 8.14595
R270 source.n60 source.n32 8.14595
R271 source.n92 source.n64 8.14595
R272 source.n124 source.n96 8.14595
R273 source.n254 source.n224 5.81868
R274 source.n222 source.n192 5.81868
R275 source.n190 source.n160 5.81868
R276 source.n158 source.n128 5.81868
R277 source.n30 source.n0 5.81868
R278 source.n62 source.n32 5.81868
R279 source.n94 source.n64 5.81868
R280 source.n126 source.n96 5.81868
R281 source.n256 source.n255 5.49188
R282 source.n252 source.n251 5.04292
R283 source.n220 source.n219 5.04292
R284 source.n188 source.n187 5.04292
R285 source.n156 source.n155 5.04292
R286 source.n28 source.n27 5.04292
R287 source.n60 source.n59 5.04292
R288 source.n92 source.n91 5.04292
R289 source.n124 source.n123 5.04292
R290 source.n237 source.n233 4.38594
R291 source.n205 source.n201 4.38594
R292 source.n173 source.n169 4.38594
R293 source.n141 source.n137 4.38594
R294 source.n13 source.n9 4.38594
R295 source.n45 source.n41 4.38594
R296 source.n77 source.n73 4.38594
R297 source.n109 source.n105 4.38594
R298 source.n248 source.n226 4.26717
R299 source.n216 source.n194 4.26717
R300 source.n184 source.n162 4.26717
R301 source.n152 source.n130 4.26717
R302 source.n24 source.n2 4.26717
R303 source.n56 source.n34 4.26717
R304 source.n88 source.n66 4.26717
R305 source.n120 source.n98 4.26717
R306 source.n247 source.n228 3.49141
R307 source.n215 source.n196 3.49141
R308 source.n183 source.n164 3.49141
R309 source.n151 source.n132 3.49141
R310 source.n23 source.n4 3.49141
R311 source.n55 source.n36 3.49141
R312 source.n87 source.n68 3.49141
R313 source.n119 source.n100 3.49141
R314 source.n244 source.n243 2.71565
R315 source.n212 source.n211 2.71565
R316 source.n180 source.n179 2.71565
R317 source.n148 source.n147 2.71565
R318 source.n20 source.n19 2.71565
R319 source.n52 source.n51 2.71565
R320 source.n84 source.n83 2.71565
R321 source.n116 source.n115 2.71565
R322 source.n240 source.n230 1.93989
R323 source.n208 source.n198 1.93989
R324 source.n176 source.n166 1.93989
R325 source.n144 source.n134 1.93989
R326 source.n16 source.n6 1.93989
R327 source.n48 source.n38 1.93989
R328 source.n80 source.n70 1.93989
R329 source.n112 source.n102 1.93989
R330 source.n239 source.n232 1.16414
R331 source.n207 source.n200 1.16414
R332 source.n175 source.n168 1.16414
R333 source.n143 source.n136 1.16414
R334 source.n15 source.n8 1.16414
R335 source.n47 source.n40 1.16414
R336 source.n79 source.n72 1.16414
R337 source.n111 source.n104 1.16414
R338 source.n95 source.n63 0.470328
R339 source.n223 source.n191 0.470328
R340 source.n127 source.n95 0.457397
R341 source.n63 source.n31 0.457397
R342 source.n191 source.n159 0.457397
R343 source.n255 source.n223 0.457397
R344 source.n236 source.n235 0.388379
R345 source.n204 source.n203 0.388379
R346 source.n172 source.n171 0.388379
R347 source.n140 source.n139 0.388379
R348 source.n12 source.n11 0.388379
R349 source.n44 source.n43 0.388379
R350 source.n76 source.n75 0.388379
R351 source.n108 source.n107 0.388379
R352 source source.n256 0.188
R353 source.n238 source.n237 0.155672
R354 source.n238 source.n229 0.155672
R355 source.n245 source.n229 0.155672
R356 source.n246 source.n245 0.155672
R357 source.n246 source.n225 0.155672
R358 source.n253 source.n225 0.155672
R359 source.n206 source.n205 0.155672
R360 source.n206 source.n197 0.155672
R361 source.n213 source.n197 0.155672
R362 source.n214 source.n213 0.155672
R363 source.n214 source.n193 0.155672
R364 source.n221 source.n193 0.155672
R365 source.n174 source.n173 0.155672
R366 source.n174 source.n165 0.155672
R367 source.n181 source.n165 0.155672
R368 source.n182 source.n181 0.155672
R369 source.n182 source.n161 0.155672
R370 source.n189 source.n161 0.155672
R371 source.n142 source.n141 0.155672
R372 source.n142 source.n133 0.155672
R373 source.n149 source.n133 0.155672
R374 source.n150 source.n149 0.155672
R375 source.n150 source.n129 0.155672
R376 source.n157 source.n129 0.155672
R377 source.n29 source.n1 0.155672
R378 source.n22 source.n1 0.155672
R379 source.n22 source.n21 0.155672
R380 source.n21 source.n5 0.155672
R381 source.n14 source.n5 0.155672
R382 source.n14 source.n13 0.155672
R383 source.n61 source.n33 0.155672
R384 source.n54 source.n33 0.155672
R385 source.n54 source.n53 0.155672
R386 source.n53 source.n37 0.155672
R387 source.n46 source.n37 0.155672
R388 source.n46 source.n45 0.155672
R389 source.n93 source.n65 0.155672
R390 source.n86 source.n65 0.155672
R391 source.n86 source.n85 0.155672
R392 source.n85 source.n69 0.155672
R393 source.n78 source.n69 0.155672
R394 source.n78 source.n77 0.155672
R395 source.n125 source.n97 0.155672
R396 source.n118 source.n97 0.155672
R397 source.n118 source.n117 0.155672
R398 source.n117 source.n101 0.155672
R399 source.n110 source.n101 0.155672
R400 source.n110 source.n109 0.155672
R401 drain_right drain_right.n0 90.3875
R402 drain_right drain_right.n1 73.3003
R403 drain_right.n0 drain_right.t2 3.3005
R404 drain_right.n0 drain_right.t1 3.3005
R405 drain_right.n1 drain_right.t0 3.3005
R406 drain_right.n1 drain_right.t3 3.3005
R407 plus.n0 plus.t2 918.356
R408 plus.n0 plus.t1 918.356
R409 plus.n1 plus.t3 918.356
R410 plus.n1 plus.t0 918.356
R411 plus plus.n1 185.893
R412 plus plus.n0 171.103
R413 drain_left drain_left.n0 90.9407
R414 drain_left drain_left.n1 73.3003
R415 drain_left.n0 drain_left.t3 3.3005
R416 drain_left.n0 drain_left.t0 3.3005
R417 drain_left.n1 drain_left.t1 3.3005
R418 drain_left.n1 drain_left.t2 3.3005
C0 drain_right source 6.20398f
C1 drain_right minus 0.998293f
C2 source minus 0.739162f
C3 drain_left plus 1.093f
C4 drain_right drain_left 0.457115f
C5 source drain_left 6.20603f
C6 drain_right plus 0.248706f
C7 source plus 0.75318f
C8 drain_left minus 0.171239f
C9 plus minus 3.32888f
C10 drain_right a_n1034_n2092# 4.9398f
C11 drain_left a_n1034_n2092# 5.07966f
C12 source a_n1034_n2092# 4.78296f
C13 minus a_n1034_n2092# 3.493806f
C14 plus a_n1034_n2092# 5.62962f
C15 drain_left.t3 a_n1034_n2092# 0.136475f
C16 drain_left.t0 a_n1034_n2092# 0.136475f
C17 drain_left.n0 a_n1034_n2092# 1.38369f
C18 drain_left.t1 a_n1034_n2092# 0.136475f
C19 drain_left.t2 a_n1034_n2092# 0.136475f
C20 drain_left.n1 a_n1034_n2092# 1.18534f
C21 plus.t2 a_n1034_n2092# 0.145279f
C22 plus.t1 a_n1034_n2092# 0.145279f
C23 plus.n0 a_n1034_n2092# 0.166648f
C24 plus.t0 a_n1034_n2092# 0.145279f
C25 plus.t3 a_n1034_n2092# 0.145279f
C26 plus.n1 a_n1034_n2092# 0.265101f
C27 drain_right.t2 a_n1034_n2092# 0.139f
C28 drain_right.t1 a_n1034_n2092# 0.139f
C29 drain_right.n0 a_n1034_n2092# 1.38946f
C30 drain_right.t0 a_n1034_n2092# 0.139f
C31 drain_right.t3 a_n1034_n2092# 0.139f
C32 drain_right.n1 a_n1034_n2092# 1.20727f
C33 source.n0 a_n1034_n2092# 0.027614f
C34 source.n1 a_n1034_n2092# 0.019645f
C35 source.n2 a_n1034_n2092# 0.010557f
C36 source.n3 a_n1034_n2092# 0.024952f
C37 source.n4 a_n1034_n2092# 0.011178f
C38 source.n5 a_n1034_n2092# 0.019645f
C39 source.n6 a_n1034_n2092# 0.010557f
C40 source.n7 a_n1034_n2092# 0.024952f
C41 source.n8 a_n1034_n2092# 0.011178f
C42 source.n9 a_n1034_n2092# 0.084069f
C43 source.t1 a_n1034_n2092# 0.040669f
C44 source.n10 a_n1034_n2092# 0.018714f
C45 source.n11 a_n1034_n2092# 0.014739f
C46 source.n12 a_n1034_n2092# 0.010557f
C47 source.n13 a_n1034_n2092# 0.467445f
C48 source.n14 a_n1034_n2092# 0.019645f
C49 source.n15 a_n1034_n2092# 0.010557f
C50 source.n16 a_n1034_n2092# 0.011178f
C51 source.n17 a_n1034_n2092# 0.024952f
C52 source.n18 a_n1034_n2092# 0.024952f
C53 source.n19 a_n1034_n2092# 0.011178f
C54 source.n20 a_n1034_n2092# 0.010557f
C55 source.n21 a_n1034_n2092# 0.019645f
C56 source.n22 a_n1034_n2092# 0.019645f
C57 source.n23 a_n1034_n2092# 0.010557f
C58 source.n24 a_n1034_n2092# 0.011178f
C59 source.n25 a_n1034_n2092# 0.024952f
C60 source.n26 a_n1034_n2092# 0.054017f
C61 source.n27 a_n1034_n2092# 0.011178f
C62 source.n28 a_n1034_n2092# 0.010557f
C63 source.n29 a_n1034_n2092# 0.04541f
C64 source.n30 a_n1034_n2092# 0.030225f
C65 source.n31 a_n1034_n2092# 0.467477f
C66 source.n32 a_n1034_n2092# 0.027614f
C67 source.n33 a_n1034_n2092# 0.019645f
C68 source.n34 a_n1034_n2092# 0.010557f
C69 source.n35 a_n1034_n2092# 0.024952f
C70 source.n36 a_n1034_n2092# 0.011178f
C71 source.n37 a_n1034_n2092# 0.019645f
C72 source.n38 a_n1034_n2092# 0.010557f
C73 source.n39 a_n1034_n2092# 0.024952f
C74 source.n40 a_n1034_n2092# 0.011178f
C75 source.n41 a_n1034_n2092# 0.084069f
C76 source.t3 a_n1034_n2092# 0.040669f
C77 source.n42 a_n1034_n2092# 0.018714f
C78 source.n43 a_n1034_n2092# 0.014739f
C79 source.n44 a_n1034_n2092# 0.010557f
C80 source.n45 a_n1034_n2092# 0.467445f
C81 source.n46 a_n1034_n2092# 0.019645f
C82 source.n47 a_n1034_n2092# 0.010557f
C83 source.n48 a_n1034_n2092# 0.011178f
C84 source.n49 a_n1034_n2092# 0.024952f
C85 source.n50 a_n1034_n2092# 0.024952f
C86 source.n51 a_n1034_n2092# 0.011178f
C87 source.n52 a_n1034_n2092# 0.010557f
C88 source.n53 a_n1034_n2092# 0.019645f
C89 source.n54 a_n1034_n2092# 0.019645f
C90 source.n55 a_n1034_n2092# 0.010557f
C91 source.n56 a_n1034_n2092# 0.011178f
C92 source.n57 a_n1034_n2092# 0.024952f
C93 source.n58 a_n1034_n2092# 0.054017f
C94 source.n59 a_n1034_n2092# 0.011178f
C95 source.n60 a_n1034_n2092# 0.010557f
C96 source.n61 a_n1034_n2092# 0.04541f
C97 source.n62 a_n1034_n2092# 0.030225f
C98 source.n63 a_n1034_n2092# 0.075442f
C99 source.n64 a_n1034_n2092# 0.027614f
C100 source.n65 a_n1034_n2092# 0.019645f
C101 source.n66 a_n1034_n2092# 0.010557f
C102 source.n67 a_n1034_n2092# 0.024952f
C103 source.n68 a_n1034_n2092# 0.011178f
C104 source.n69 a_n1034_n2092# 0.019645f
C105 source.n70 a_n1034_n2092# 0.010557f
C106 source.n71 a_n1034_n2092# 0.024952f
C107 source.n72 a_n1034_n2092# 0.011178f
C108 source.n73 a_n1034_n2092# 0.084069f
C109 source.t7 a_n1034_n2092# 0.040669f
C110 source.n74 a_n1034_n2092# 0.018714f
C111 source.n75 a_n1034_n2092# 0.014739f
C112 source.n76 a_n1034_n2092# 0.010557f
C113 source.n77 a_n1034_n2092# 0.467445f
C114 source.n78 a_n1034_n2092# 0.019645f
C115 source.n79 a_n1034_n2092# 0.010557f
C116 source.n80 a_n1034_n2092# 0.011178f
C117 source.n81 a_n1034_n2092# 0.024952f
C118 source.n82 a_n1034_n2092# 0.024952f
C119 source.n83 a_n1034_n2092# 0.011178f
C120 source.n84 a_n1034_n2092# 0.010557f
C121 source.n85 a_n1034_n2092# 0.019645f
C122 source.n86 a_n1034_n2092# 0.019645f
C123 source.n87 a_n1034_n2092# 0.010557f
C124 source.n88 a_n1034_n2092# 0.011178f
C125 source.n89 a_n1034_n2092# 0.024952f
C126 source.n90 a_n1034_n2092# 0.054017f
C127 source.n91 a_n1034_n2092# 0.011178f
C128 source.n92 a_n1034_n2092# 0.010557f
C129 source.n93 a_n1034_n2092# 0.04541f
C130 source.n94 a_n1034_n2092# 0.030225f
C131 source.n95 a_n1034_n2092# 0.075442f
C132 source.n96 a_n1034_n2092# 0.027614f
C133 source.n97 a_n1034_n2092# 0.019645f
C134 source.n98 a_n1034_n2092# 0.010557f
C135 source.n99 a_n1034_n2092# 0.024952f
C136 source.n100 a_n1034_n2092# 0.011178f
C137 source.n101 a_n1034_n2092# 0.019645f
C138 source.n102 a_n1034_n2092# 0.010557f
C139 source.n103 a_n1034_n2092# 0.024952f
C140 source.n104 a_n1034_n2092# 0.011178f
C141 source.n105 a_n1034_n2092# 0.084069f
C142 source.t4 a_n1034_n2092# 0.040669f
C143 source.n106 a_n1034_n2092# 0.018714f
C144 source.n107 a_n1034_n2092# 0.014739f
C145 source.n108 a_n1034_n2092# 0.010557f
C146 source.n109 a_n1034_n2092# 0.467445f
C147 source.n110 a_n1034_n2092# 0.019645f
C148 source.n111 a_n1034_n2092# 0.010557f
C149 source.n112 a_n1034_n2092# 0.011178f
C150 source.n113 a_n1034_n2092# 0.024952f
C151 source.n114 a_n1034_n2092# 0.024952f
C152 source.n115 a_n1034_n2092# 0.011178f
C153 source.n116 a_n1034_n2092# 0.010557f
C154 source.n117 a_n1034_n2092# 0.019645f
C155 source.n118 a_n1034_n2092# 0.019645f
C156 source.n119 a_n1034_n2092# 0.010557f
C157 source.n120 a_n1034_n2092# 0.011178f
C158 source.n121 a_n1034_n2092# 0.024952f
C159 source.n122 a_n1034_n2092# 0.054017f
C160 source.n123 a_n1034_n2092# 0.011178f
C161 source.n124 a_n1034_n2092# 0.010557f
C162 source.n125 a_n1034_n2092# 0.04541f
C163 source.n126 a_n1034_n2092# 0.030225f
C164 source.n127 a_n1034_n2092# 0.719096f
C165 source.n128 a_n1034_n2092# 0.027614f
C166 source.n129 a_n1034_n2092# 0.019645f
C167 source.n130 a_n1034_n2092# 0.010557f
C168 source.n131 a_n1034_n2092# 0.024952f
C169 source.n132 a_n1034_n2092# 0.011178f
C170 source.n133 a_n1034_n2092# 0.019645f
C171 source.n134 a_n1034_n2092# 0.010557f
C172 source.n135 a_n1034_n2092# 0.024952f
C173 source.n136 a_n1034_n2092# 0.011178f
C174 source.n137 a_n1034_n2092# 0.084069f
C175 source.t0 a_n1034_n2092# 0.040669f
C176 source.n138 a_n1034_n2092# 0.018714f
C177 source.n139 a_n1034_n2092# 0.014739f
C178 source.n140 a_n1034_n2092# 0.010557f
C179 source.n141 a_n1034_n2092# 0.467445f
C180 source.n142 a_n1034_n2092# 0.019645f
C181 source.n143 a_n1034_n2092# 0.010557f
C182 source.n144 a_n1034_n2092# 0.011178f
C183 source.n145 a_n1034_n2092# 0.024952f
C184 source.n146 a_n1034_n2092# 0.024952f
C185 source.n147 a_n1034_n2092# 0.011178f
C186 source.n148 a_n1034_n2092# 0.010557f
C187 source.n149 a_n1034_n2092# 0.019645f
C188 source.n150 a_n1034_n2092# 0.019645f
C189 source.n151 a_n1034_n2092# 0.010557f
C190 source.n152 a_n1034_n2092# 0.011178f
C191 source.n153 a_n1034_n2092# 0.024952f
C192 source.n154 a_n1034_n2092# 0.054017f
C193 source.n155 a_n1034_n2092# 0.011178f
C194 source.n156 a_n1034_n2092# 0.010557f
C195 source.n157 a_n1034_n2092# 0.04541f
C196 source.n158 a_n1034_n2092# 0.030225f
C197 source.n159 a_n1034_n2092# 0.719096f
C198 source.n160 a_n1034_n2092# 0.027614f
C199 source.n161 a_n1034_n2092# 0.019645f
C200 source.n162 a_n1034_n2092# 0.010557f
C201 source.n163 a_n1034_n2092# 0.024952f
C202 source.n164 a_n1034_n2092# 0.011178f
C203 source.n165 a_n1034_n2092# 0.019645f
C204 source.n166 a_n1034_n2092# 0.010557f
C205 source.n167 a_n1034_n2092# 0.024952f
C206 source.n168 a_n1034_n2092# 0.011178f
C207 source.n169 a_n1034_n2092# 0.084069f
C208 source.t2 a_n1034_n2092# 0.040669f
C209 source.n170 a_n1034_n2092# 0.018714f
C210 source.n171 a_n1034_n2092# 0.014739f
C211 source.n172 a_n1034_n2092# 0.010557f
C212 source.n173 a_n1034_n2092# 0.467445f
C213 source.n174 a_n1034_n2092# 0.019645f
C214 source.n175 a_n1034_n2092# 0.010557f
C215 source.n176 a_n1034_n2092# 0.011178f
C216 source.n177 a_n1034_n2092# 0.024952f
C217 source.n178 a_n1034_n2092# 0.024952f
C218 source.n179 a_n1034_n2092# 0.011178f
C219 source.n180 a_n1034_n2092# 0.010557f
C220 source.n181 a_n1034_n2092# 0.019645f
C221 source.n182 a_n1034_n2092# 0.019645f
C222 source.n183 a_n1034_n2092# 0.010557f
C223 source.n184 a_n1034_n2092# 0.011178f
C224 source.n185 a_n1034_n2092# 0.024952f
C225 source.n186 a_n1034_n2092# 0.054017f
C226 source.n187 a_n1034_n2092# 0.011178f
C227 source.n188 a_n1034_n2092# 0.010557f
C228 source.n189 a_n1034_n2092# 0.04541f
C229 source.n190 a_n1034_n2092# 0.030225f
C230 source.n191 a_n1034_n2092# 0.075442f
C231 source.n192 a_n1034_n2092# 0.027614f
C232 source.n193 a_n1034_n2092# 0.019645f
C233 source.n194 a_n1034_n2092# 0.010557f
C234 source.n195 a_n1034_n2092# 0.024952f
C235 source.n196 a_n1034_n2092# 0.011178f
C236 source.n197 a_n1034_n2092# 0.019645f
C237 source.n198 a_n1034_n2092# 0.010557f
C238 source.n199 a_n1034_n2092# 0.024952f
C239 source.n200 a_n1034_n2092# 0.011178f
C240 source.n201 a_n1034_n2092# 0.084069f
C241 source.t6 a_n1034_n2092# 0.040669f
C242 source.n202 a_n1034_n2092# 0.018714f
C243 source.n203 a_n1034_n2092# 0.014739f
C244 source.n204 a_n1034_n2092# 0.010557f
C245 source.n205 a_n1034_n2092# 0.467445f
C246 source.n206 a_n1034_n2092# 0.019645f
C247 source.n207 a_n1034_n2092# 0.010557f
C248 source.n208 a_n1034_n2092# 0.011178f
C249 source.n209 a_n1034_n2092# 0.024952f
C250 source.n210 a_n1034_n2092# 0.024952f
C251 source.n211 a_n1034_n2092# 0.011178f
C252 source.n212 a_n1034_n2092# 0.010557f
C253 source.n213 a_n1034_n2092# 0.019645f
C254 source.n214 a_n1034_n2092# 0.019645f
C255 source.n215 a_n1034_n2092# 0.010557f
C256 source.n216 a_n1034_n2092# 0.011178f
C257 source.n217 a_n1034_n2092# 0.024952f
C258 source.n218 a_n1034_n2092# 0.054017f
C259 source.n219 a_n1034_n2092# 0.011178f
C260 source.n220 a_n1034_n2092# 0.010557f
C261 source.n221 a_n1034_n2092# 0.04541f
C262 source.n222 a_n1034_n2092# 0.030225f
C263 source.n223 a_n1034_n2092# 0.075442f
C264 source.n224 a_n1034_n2092# 0.027614f
C265 source.n225 a_n1034_n2092# 0.019645f
C266 source.n226 a_n1034_n2092# 0.010557f
C267 source.n227 a_n1034_n2092# 0.024952f
C268 source.n228 a_n1034_n2092# 0.011178f
C269 source.n229 a_n1034_n2092# 0.019645f
C270 source.n230 a_n1034_n2092# 0.010557f
C271 source.n231 a_n1034_n2092# 0.024952f
C272 source.n232 a_n1034_n2092# 0.011178f
C273 source.n233 a_n1034_n2092# 0.084069f
C274 source.t5 a_n1034_n2092# 0.040669f
C275 source.n234 a_n1034_n2092# 0.018714f
C276 source.n235 a_n1034_n2092# 0.014739f
C277 source.n236 a_n1034_n2092# 0.010557f
C278 source.n237 a_n1034_n2092# 0.467445f
C279 source.n238 a_n1034_n2092# 0.019645f
C280 source.n239 a_n1034_n2092# 0.010557f
C281 source.n240 a_n1034_n2092# 0.011178f
C282 source.n241 a_n1034_n2092# 0.024952f
C283 source.n242 a_n1034_n2092# 0.024952f
C284 source.n243 a_n1034_n2092# 0.011178f
C285 source.n244 a_n1034_n2092# 0.010557f
C286 source.n245 a_n1034_n2092# 0.019645f
C287 source.n246 a_n1034_n2092# 0.019645f
C288 source.n247 a_n1034_n2092# 0.010557f
C289 source.n248 a_n1034_n2092# 0.011178f
C290 source.n249 a_n1034_n2092# 0.024952f
C291 source.n250 a_n1034_n2092# 0.054017f
C292 source.n251 a_n1034_n2092# 0.011178f
C293 source.n252 a_n1034_n2092# 0.010557f
C294 source.n253 a_n1034_n2092# 0.04541f
C295 source.n254 a_n1034_n2092# 0.030225f
C296 source.n255 a_n1034_n2092# 0.181966f
C297 source.n256 a_n1034_n2092# 0.802722f
C298 minus.t3 a_n1034_n2092# 0.141663f
C299 minus.t0 a_n1034_n2092# 0.141663f
C300 minus.n0 a_n1034_n2092# 0.28739f
C301 minus.t1 a_n1034_n2092# 0.141663f
C302 minus.t2 a_n1034_n2092# 0.141663f
C303 minus.n1 a_n1034_n2092# 0.152775f
C304 minus.n2 a_n1034_n2092# 2.26651f
.ends

