* NGSPICE file created from diffpair686.ext - technology: sky130A

.subckt diffpair686 minus drain_right drain_left source plus
X0 a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.5
X1 drain_right.t13 minus.t0 source.t27 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.5
X2 a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.5
X3 source.t18 minus.t1 drain_right.t12 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X4 source.t12 plus.t0 drain_left.t13 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X5 drain_left.t12 plus.t1 source.t4 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X6 drain_left.t11 plus.t2 source.t13 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.5
X7 source.t26 minus.t2 drain_right.t11 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X8 drain_right.t10 minus.t3 source.t20 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.5
X9 drain_right.t9 minus.t4 source.t19 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X10 drain_right.t8 minus.t5 source.t15 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X11 drain_right.t7 minus.t6 source.t17 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X12 drain_left.t10 plus.t3 source.t2 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.5
X13 source.t7 plus.t4 drain_left.t9 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X14 a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.5
X15 drain_left.t8 plus.t5 source.t10 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X16 a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.5
X17 drain_left.t7 plus.t6 source.t5 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.5
X18 source.t14 minus.t7 drain_right.t6 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X19 source.t6 plus.t7 drain_left.t6 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X20 source.t24 minus.t8 drain_right.t5 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X21 drain_right.t4 minus.t9 source.t23 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X22 drain_right.t3 minus.t10 source.t22 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.5
X23 source.t9 plus.t8 drain_left.t5 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X24 drain_right.t2 minus.t11 source.t21 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.5
X25 source.t25 minus.t12 drain_right.t1 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X26 source.t16 minus.t13 drain_right.t0 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X27 drain_left.t4 plus.t9 source.t0 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X28 drain_left.t3 plus.t10 source.t8 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X29 source.t11 plus.t11 drain_left.t2 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
X30 drain_left.t1 plus.t12 source.t1 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.5
X31 source.t3 plus.t13 drain_left.t0 a_n2044_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.5
R0 minus.n4 minus.t10 1304.55
R1 minus.n20 minus.t3 1304.55
R2 minus.n3 minus.t1 1283.57
R3 minus.n7 minus.t5 1283.57
R4 minus.n8 minus.t13 1283.57
R5 minus.n1 minus.t4 1283.57
R6 minus.n13 minus.t7 1283.57
R7 minus.n14 minus.t0 1283.57
R8 minus.n19 minus.t2 1283.57
R9 minus.n23 minus.t9 1283.57
R10 minus.n24 minus.t8 1283.57
R11 minus.n17 minus.t6 1283.57
R12 minus.n29 minus.t12 1283.57
R13 minus.n30 minus.t11 1283.57
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n0 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n1 161.3
R18 minus.n7 minus.n2 161.3
R19 minus.n6 minus.n5 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n16 161.3
R22 minus.n28 minus.n27 161.3
R23 minus.n26 minus.n17 161.3
R24 minus.n23 minus.n18 161.3
R25 minus.n22 minus.n21 161.3
R26 minus.n9 minus.n8 80.6037
R27 minus.n25 minus.n24 80.6037
R28 minus.n5 minus.n4 70.4033
R29 minus.n21 minus.n20 70.4033
R30 minus.n8 minus.n7 48.2005
R31 minus.n8 minus.n1 48.2005
R32 minus.n14 minus.n13 48.2005
R33 minus.n24 minus.n23 48.2005
R34 minus.n24 minus.n17 48.2005
R35 minus.n30 minus.n29 48.2005
R36 minus.n32 minus.n15 46.8054
R37 minus.n7 minus.n6 24.8308
R38 minus.n12 minus.n1 24.8308
R39 minus.n23 minus.n22 24.8308
R40 minus.n28 minus.n17 24.8308
R41 minus.n6 minus.n3 23.3702
R42 minus.n13 minus.n12 23.3702
R43 minus.n22 minus.n19 23.3702
R44 minus.n29 minus.n28 23.3702
R45 minus.n4 minus.n3 20.9576
R46 minus.n20 minus.n19 20.9576
R47 minus.n32 minus.n31 6.5933
R48 minus.n10 minus.n9 0.285035
R49 minus.n9 minus.n2 0.285035
R50 minus.n25 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n5 minus.n2 0.189894
R56 minus.n21 minus.n18 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n16 0.189894
R59 minus.n31 minus.n16 0.189894
R60 minus minus.n32 0.188
R61 source.n578 source.n444 289.615
R62 source.n432 source.n298 289.615
R63 source.n134 source.n0 289.615
R64 source.n280 source.n146 289.615
R65 source.n488 source.n487 185
R66 source.n493 source.n492 185
R67 source.n495 source.n494 185
R68 source.n484 source.n483 185
R69 source.n501 source.n500 185
R70 source.n503 source.n502 185
R71 source.n480 source.n479 185
R72 source.n510 source.n509 185
R73 source.n511 source.n478 185
R74 source.n513 source.n512 185
R75 source.n476 source.n475 185
R76 source.n519 source.n518 185
R77 source.n521 source.n520 185
R78 source.n472 source.n471 185
R79 source.n527 source.n526 185
R80 source.n529 source.n528 185
R81 source.n468 source.n467 185
R82 source.n535 source.n534 185
R83 source.n537 source.n536 185
R84 source.n464 source.n463 185
R85 source.n543 source.n542 185
R86 source.n545 source.n544 185
R87 source.n460 source.n459 185
R88 source.n551 source.n550 185
R89 source.n554 source.n553 185
R90 source.n552 source.n456 185
R91 source.n559 source.n455 185
R92 source.n561 source.n560 185
R93 source.n563 source.n562 185
R94 source.n452 source.n451 185
R95 source.n569 source.n568 185
R96 source.n571 source.n570 185
R97 source.n448 source.n447 185
R98 source.n577 source.n576 185
R99 source.n579 source.n578 185
R100 source.n342 source.n341 185
R101 source.n347 source.n346 185
R102 source.n349 source.n348 185
R103 source.n338 source.n337 185
R104 source.n355 source.n354 185
R105 source.n357 source.n356 185
R106 source.n334 source.n333 185
R107 source.n364 source.n363 185
R108 source.n365 source.n332 185
R109 source.n367 source.n366 185
R110 source.n330 source.n329 185
R111 source.n373 source.n372 185
R112 source.n375 source.n374 185
R113 source.n326 source.n325 185
R114 source.n381 source.n380 185
R115 source.n383 source.n382 185
R116 source.n322 source.n321 185
R117 source.n389 source.n388 185
R118 source.n391 source.n390 185
R119 source.n318 source.n317 185
R120 source.n397 source.n396 185
R121 source.n399 source.n398 185
R122 source.n314 source.n313 185
R123 source.n405 source.n404 185
R124 source.n408 source.n407 185
R125 source.n406 source.n310 185
R126 source.n413 source.n309 185
R127 source.n415 source.n414 185
R128 source.n417 source.n416 185
R129 source.n306 source.n305 185
R130 source.n423 source.n422 185
R131 source.n425 source.n424 185
R132 source.n302 source.n301 185
R133 source.n431 source.n430 185
R134 source.n433 source.n432 185
R135 source.n135 source.n134 185
R136 source.n133 source.n132 185
R137 source.n4 source.n3 185
R138 source.n127 source.n126 185
R139 source.n125 source.n124 185
R140 source.n8 source.n7 185
R141 source.n119 source.n118 185
R142 source.n117 source.n116 185
R143 source.n115 source.n11 185
R144 source.n15 source.n12 185
R145 source.n110 source.n109 185
R146 source.n108 source.n107 185
R147 source.n17 source.n16 185
R148 source.n102 source.n101 185
R149 source.n100 source.n99 185
R150 source.n21 source.n20 185
R151 source.n94 source.n93 185
R152 source.n92 source.n91 185
R153 source.n25 source.n24 185
R154 source.n86 source.n85 185
R155 source.n84 source.n83 185
R156 source.n29 source.n28 185
R157 source.n78 source.n77 185
R158 source.n76 source.n75 185
R159 source.n33 source.n32 185
R160 source.n70 source.n69 185
R161 source.n68 source.n35 185
R162 source.n67 source.n66 185
R163 source.n38 source.n36 185
R164 source.n61 source.n60 185
R165 source.n59 source.n58 185
R166 source.n42 source.n41 185
R167 source.n53 source.n52 185
R168 source.n51 source.n50 185
R169 source.n46 source.n45 185
R170 source.n281 source.n280 185
R171 source.n279 source.n278 185
R172 source.n150 source.n149 185
R173 source.n273 source.n272 185
R174 source.n271 source.n270 185
R175 source.n154 source.n153 185
R176 source.n265 source.n264 185
R177 source.n263 source.n262 185
R178 source.n261 source.n157 185
R179 source.n161 source.n158 185
R180 source.n256 source.n255 185
R181 source.n254 source.n253 185
R182 source.n163 source.n162 185
R183 source.n248 source.n247 185
R184 source.n246 source.n245 185
R185 source.n167 source.n166 185
R186 source.n240 source.n239 185
R187 source.n238 source.n237 185
R188 source.n171 source.n170 185
R189 source.n232 source.n231 185
R190 source.n230 source.n229 185
R191 source.n175 source.n174 185
R192 source.n224 source.n223 185
R193 source.n222 source.n221 185
R194 source.n179 source.n178 185
R195 source.n216 source.n215 185
R196 source.n214 source.n181 185
R197 source.n213 source.n212 185
R198 source.n184 source.n182 185
R199 source.n207 source.n206 185
R200 source.n205 source.n204 185
R201 source.n188 source.n187 185
R202 source.n199 source.n198 185
R203 source.n197 source.n196 185
R204 source.n192 source.n191 185
R205 source.n489 source.t21 149.524
R206 source.n343 source.t1 149.524
R207 source.n47 source.t5 149.524
R208 source.n193 source.t22 149.524
R209 source.n493 source.n487 104.615
R210 source.n494 source.n493 104.615
R211 source.n494 source.n483 104.615
R212 source.n501 source.n483 104.615
R213 source.n502 source.n501 104.615
R214 source.n502 source.n479 104.615
R215 source.n510 source.n479 104.615
R216 source.n511 source.n510 104.615
R217 source.n512 source.n511 104.615
R218 source.n512 source.n475 104.615
R219 source.n519 source.n475 104.615
R220 source.n520 source.n519 104.615
R221 source.n520 source.n471 104.615
R222 source.n527 source.n471 104.615
R223 source.n528 source.n527 104.615
R224 source.n528 source.n467 104.615
R225 source.n535 source.n467 104.615
R226 source.n536 source.n535 104.615
R227 source.n536 source.n463 104.615
R228 source.n543 source.n463 104.615
R229 source.n544 source.n543 104.615
R230 source.n544 source.n459 104.615
R231 source.n551 source.n459 104.615
R232 source.n553 source.n551 104.615
R233 source.n553 source.n552 104.615
R234 source.n552 source.n455 104.615
R235 source.n561 source.n455 104.615
R236 source.n562 source.n561 104.615
R237 source.n562 source.n451 104.615
R238 source.n569 source.n451 104.615
R239 source.n570 source.n569 104.615
R240 source.n570 source.n447 104.615
R241 source.n577 source.n447 104.615
R242 source.n578 source.n577 104.615
R243 source.n347 source.n341 104.615
R244 source.n348 source.n347 104.615
R245 source.n348 source.n337 104.615
R246 source.n355 source.n337 104.615
R247 source.n356 source.n355 104.615
R248 source.n356 source.n333 104.615
R249 source.n364 source.n333 104.615
R250 source.n365 source.n364 104.615
R251 source.n366 source.n365 104.615
R252 source.n366 source.n329 104.615
R253 source.n373 source.n329 104.615
R254 source.n374 source.n373 104.615
R255 source.n374 source.n325 104.615
R256 source.n381 source.n325 104.615
R257 source.n382 source.n381 104.615
R258 source.n382 source.n321 104.615
R259 source.n389 source.n321 104.615
R260 source.n390 source.n389 104.615
R261 source.n390 source.n317 104.615
R262 source.n397 source.n317 104.615
R263 source.n398 source.n397 104.615
R264 source.n398 source.n313 104.615
R265 source.n405 source.n313 104.615
R266 source.n407 source.n405 104.615
R267 source.n407 source.n406 104.615
R268 source.n406 source.n309 104.615
R269 source.n415 source.n309 104.615
R270 source.n416 source.n415 104.615
R271 source.n416 source.n305 104.615
R272 source.n423 source.n305 104.615
R273 source.n424 source.n423 104.615
R274 source.n424 source.n301 104.615
R275 source.n431 source.n301 104.615
R276 source.n432 source.n431 104.615
R277 source.n134 source.n133 104.615
R278 source.n133 source.n3 104.615
R279 source.n126 source.n3 104.615
R280 source.n126 source.n125 104.615
R281 source.n125 source.n7 104.615
R282 source.n118 source.n7 104.615
R283 source.n118 source.n117 104.615
R284 source.n117 source.n11 104.615
R285 source.n15 source.n11 104.615
R286 source.n109 source.n15 104.615
R287 source.n109 source.n108 104.615
R288 source.n108 source.n16 104.615
R289 source.n101 source.n16 104.615
R290 source.n101 source.n100 104.615
R291 source.n100 source.n20 104.615
R292 source.n93 source.n20 104.615
R293 source.n93 source.n92 104.615
R294 source.n92 source.n24 104.615
R295 source.n85 source.n24 104.615
R296 source.n85 source.n84 104.615
R297 source.n84 source.n28 104.615
R298 source.n77 source.n28 104.615
R299 source.n77 source.n76 104.615
R300 source.n76 source.n32 104.615
R301 source.n69 source.n32 104.615
R302 source.n69 source.n68 104.615
R303 source.n68 source.n67 104.615
R304 source.n67 source.n36 104.615
R305 source.n60 source.n36 104.615
R306 source.n60 source.n59 104.615
R307 source.n59 source.n41 104.615
R308 source.n52 source.n41 104.615
R309 source.n52 source.n51 104.615
R310 source.n51 source.n45 104.615
R311 source.n280 source.n279 104.615
R312 source.n279 source.n149 104.615
R313 source.n272 source.n149 104.615
R314 source.n272 source.n271 104.615
R315 source.n271 source.n153 104.615
R316 source.n264 source.n153 104.615
R317 source.n264 source.n263 104.615
R318 source.n263 source.n157 104.615
R319 source.n161 source.n157 104.615
R320 source.n255 source.n161 104.615
R321 source.n255 source.n254 104.615
R322 source.n254 source.n162 104.615
R323 source.n247 source.n162 104.615
R324 source.n247 source.n246 104.615
R325 source.n246 source.n166 104.615
R326 source.n239 source.n166 104.615
R327 source.n239 source.n238 104.615
R328 source.n238 source.n170 104.615
R329 source.n231 source.n170 104.615
R330 source.n231 source.n230 104.615
R331 source.n230 source.n174 104.615
R332 source.n223 source.n174 104.615
R333 source.n223 source.n222 104.615
R334 source.n222 source.n178 104.615
R335 source.n215 source.n178 104.615
R336 source.n215 source.n214 104.615
R337 source.n214 source.n213 104.615
R338 source.n213 source.n182 104.615
R339 source.n206 source.n182 104.615
R340 source.n206 source.n205 104.615
R341 source.n205 source.n187 104.615
R342 source.n198 source.n187 104.615
R343 source.n198 source.n197 104.615
R344 source.n197 source.n191 104.615
R345 source.t21 source.n487 52.3082
R346 source.t1 source.n341 52.3082
R347 source.t5 source.n45 52.3082
R348 source.t22 source.n191 52.3082
R349 source.n443 source.n442 42.0366
R350 source.n441 source.n440 42.0366
R351 source.n439 source.n438 42.0366
R352 source.n297 source.n296 42.0366
R353 source.n295 source.n294 42.0366
R354 source.n293 source.n292 42.0366
R355 source.n141 source.n140 42.0366
R356 source.n143 source.n142 42.0366
R357 source.n145 source.n144 42.0366
R358 source.n287 source.n286 42.0366
R359 source.n289 source.n288 42.0366
R360 source.n291 source.n290 42.0366
R361 source.n293 source.n291 32.5672
R362 source.n583 source.n582 30.6338
R363 source.n437 source.n436 30.6338
R364 source.n139 source.n138 30.6338
R365 source.n285 source.n284 30.6338
R366 source.n584 source.n139 26.231
R367 source.n513 source.n478 13.1884
R368 source.n560 source.n559 13.1884
R369 source.n367 source.n332 13.1884
R370 source.n414 source.n413 13.1884
R371 source.n116 source.n115 13.1884
R372 source.n70 source.n35 13.1884
R373 source.n262 source.n261 13.1884
R374 source.n216 source.n181 13.1884
R375 source.n509 source.n508 12.8005
R376 source.n514 source.n476 12.8005
R377 source.n558 source.n456 12.8005
R378 source.n563 source.n454 12.8005
R379 source.n363 source.n362 12.8005
R380 source.n368 source.n330 12.8005
R381 source.n412 source.n310 12.8005
R382 source.n417 source.n308 12.8005
R383 source.n119 source.n10 12.8005
R384 source.n114 source.n12 12.8005
R385 source.n71 source.n33 12.8005
R386 source.n66 source.n37 12.8005
R387 source.n265 source.n156 12.8005
R388 source.n260 source.n158 12.8005
R389 source.n217 source.n179 12.8005
R390 source.n212 source.n183 12.8005
R391 source.n507 source.n480 12.0247
R392 source.n518 source.n517 12.0247
R393 source.n555 source.n554 12.0247
R394 source.n564 source.n452 12.0247
R395 source.n361 source.n334 12.0247
R396 source.n372 source.n371 12.0247
R397 source.n409 source.n408 12.0247
R398 source.n418 source.n306 12.0247
R399 source.n120 source.n8 12.0247
R400 source.n111 source.n110 12.0247
R401 source.n75 source.n74 12.0247
R402 source.n65 source.n38 12.0247
R403 source.n266 source.n154 12.0247
R404 source.n257 source.n256 12.0247
R405 source.n221 source.n220 12.0247
R406 source.n211 source.n184 12.0247
R407 source.n504 source.n503 11.249
R408 source.n521 source.n474 11.249
R409 source.n550 source.n458 11.249
R410 source.n568 source.n567 11.249
R411 source.n358 source.n357 11.249
R412 source.n375 source.n328 11.249
R413 source.n404 source.n312 11.249
R414 source.n422 source.n421 11.249
R415 source.n124 source.n123 11.249
R416 source.n107 source.n14 11.249
R417 source.n78 source.n31 11.249
R418 source.n62 source.n61 11.249
R419 source.n270 source.n269 11.249
R420 source.n253 source.n160 11.249
R421 source.n224 source.n177 11.249
R422 source.n208 source.n207 11.249
R423 source.n500 source.n482 10.4732
R424 source.n522 source.n472 10.4732
R425 source.n549 source.n460 10.4732
R426 source.n571 source.n450 10.4732
R427 source.n354 source.n336 10.4732
R428 source.n376 source.n326 10.4732
R429 source.n403 source.n314 10.4732
R430 source.n425 source.n304 10.4732
R431 source.n127 source.n6 10.4732
R432 source.n106 source.n17 10.4732
R433 source.n79 source.n29 10.4732
R434 source.n58 source.n40 10.4732
R435 source.n273 source.n152 10.4732
R436 source.n252 source.n163 10.4732
R437 source.n225 source.n175 10.4732
R438 source.n204 source.n186 10.4732
R439 source.n489 source.n488 10.2747
R440 source.n343 source.n342 10.2747
R441 source.n47 source.n46 10.2747
R442 source.n193 source.n192 10.2747
R443 source.n499 source.n484 9.69747
R444 source.n526 source.n525 9.69747
R445 source.n546 source.n545 9.69747
R446 source.n572 source.n448 9.69747
R447 source.n353 source.n338 9.69747
R448 source.n380 source.n379 9.69747
R449 source.n400 source.n399 9.69747
R450 source.n426 source.n302 9.69747
R451 source.n128 source.n4 9.69747
R452 source.n103 source.n102 9.69747
R453 source.n83 source.n82 9.69747
R454 source.n57 source.n42 9.69747
R455 source.n274 source.n150 9.69747
R456 source.n249 source.n248 9.69747
R457 source.n229 source.n228 9.69747
R458 source.n203 source.n188 9.69747
R459 source.n582 source.n581 9.45567
R460 source.n436 source.n435 9.45567
R461 source.n138 source.n137 9.45567
R462 source.n284 source.n283 9.45567
R463 source.n446 source.n445 9.3005
R464 source.n575 source.n574 9.3005
R465 source.n573 source.n572 9.3005
R466 source.n450 source.n449 9.3005
R467 source.n567 source.n566 9.3005
R468 source.n565 source.n564 9.3005
R469 source.n454 source.n453 9.3005
R470 source.n533 source.n532 9.3005
R471 source.n531 source.n530 9.3005
R472 source.n470 source.n469 9.3005
R473 source.n525 source.n524 9.3005
R474 source.n523 source.n522 9.3005
R475 source.n474 source.n473 9.3005
R476 source.n517 source.n516 9.3005
R477 source.n515 source.n514 9.3005
R478 source.n491 source.n490 9.3005
R479 source.n486 source.n485 9.3005
R480 source.n497 source.n496 9.3005
R481 source.n499 source.n498 9.3005
R482 source.n482 source.n481 9.3005
R483 source.n505 source.n504 9.3005
R484 source.n507 source.n506 9.3005
R485 source.n508 source.n477 9.3005
R486 source.n466 source.n465 9.3005
R487 source.n539 source.n538 9.3005
R488 source.n541 source.n540 9.3005
R489 source.n462 source.n461 9.3005
R490 source.n547 source.n546 9.3005
R491 source.n549 source.n548 9.3005
R492 source.n458 source.n457 9.3005
R493 source.n556 source.n555 9.3005
R494 source.n558 source.n557 9.3005
R495 source.n581 source.n580 9.3005
R496 source.n300 source.n299 9.3005
R497 source.n429 source.n428 9.3005
R498 source.n427 source.n426 9.3005
R499 source.n304 source.n303 9.3005
R500 source.n421 source.n420 9.3005
R501 source.n419 source.n418 9.3005
R502 source.n308 source.n307 9.3005
R503 source.n387 source.n386 9.3005
R504 source.n385 source.n384 9.3005
R505 source.n324 source.n323 9.3005
R506 source.n379 source.n378 9.3005
R507 source.n377 source.n376 9.3005
R508 source.n328 source.n327 9.3005
R509 source.n371 source.n370 9.3005
R510 source.n369 source.n368 9.3005
R511 source.n345 source.n344 9.3005
R512 source.n340 source.n339 9.3005
R513 source.n351 source.n350 9.3005
R514 source.n353 source.n352 9.3005
R515 source.n336 source.n335 9.3005
R516 source.n359 source.n358 9.3005
R517 source.n361 source.n360 9.3005
R518 source.n362 source.n331 9.3005
R519 source.n320 source.n319 9.3005
R520 source.n393 source.n392 9.3005
R521 source.n395 source.n394 9.3005
R522 source.n316 source.n315 9.3005
R523 source.n401 source.n400 9.3005
R524 source.n403 source.n402 9.3005
R525 source.n312 source.n311 9.3005
R526 source.n410 source.n409 9.3005
R527 source.n412 source.n411 9.3005
R528 source.n435 source.n434 9.3005
R529 source.n49 source.n48 9.3005
R530 source.n44 source.n43 9.3005
R531 source.n55 source.n54 9.3005
R532 source.n57 source.n56 9.3005
R533 source.n40 source.n39 9.3005
R534 source.n63 source.n62 9.3005
R535 source.n65 source.n64 9.3005
R536 source.n37 source.n34 9.3005
R537 source.n96 source.n95 9.3005
R538 source.n98 source.n97 9.3005
R539 source.n19 source.n18 9.3005
R540 source.n104 source.n103 9.3005
R541 source.n106 source.n105 9.3005
R542 source.n14 source.n13 9.3005
R543 source.n112 source.n111 9.3005
R544 source.n114 source.n113 9.3005
R545 source.n137 source.n136 9.3005
R546 source.n2 source.n1 9.3005
R547 source.n131 source.n130 9.3005
R548 source.n129 source.n128 9.3005
R549 source.n6 source.n5 9.3005
R550 source.n123 source.n122 9.3005
R551 source.n121 source.n120 9.3005
R552 source.n10 source.n9 9.3005
R553 source.n23 source.n22 9.3005
R554 source.n90 source.n89 9.3005
R555 source.n88 source.n87 9.3005
R556 source.n27 source.n26 9.3005
R557 source.n82 source.n81 9.3005
R558 source.n80 source.n79 9.3005
R559 source.n31 source.n30 9.3005
R560 source.n74 source.n73 9.3005
R561 source.n72 source.n71 9.3005
R562 source.n195 source.n194 9.3005
R563 source.n190 source.n189 9.3005
R564 source.n201 source.n200 9.3005
R565 source.n203 source.n202 9.3005
R566 source.n186 source.n185 9.3005
R567 source.n209 source.n208 9.3005
R568 source.n211 source.n210 9.3005
R569 source.n183 source.n180 9.3005
R570 source.n242 source.n241 9.3005
R571 source.n244 source.n243 9.3005
R572 source.n165 source.n164 9.3005
R573 source.n250 source.n249 9.3005
R574 source.n252 source.n251 9.3005
R575 source.n160 source.n159 9.3005
R576 source.n258 source.n257 9.3005
R577 source.n260 source.n259 9.3005
R578 source.n283 source.n282 9.3005
R579 source.n148 source.n147 9.3005
R580 source.n277 source.n276 9.3005
R581 source.n275 source.n274 9.3005
R582 source.n152 source.n151 9.3005
R583 source.n269 source.n268 9.3005
R584 source.n267 source.n266 9.3005
R585 source.n156 source.n155 9.3005
R586 source.n169 source.n168 9.3005
R587 source.n236 source.n235 9.3005
R588 source.n234 source.n233 9.3005
R589 source.n173 source.n172 9.3005
R590 source.n228 source.n227 9.3005
R591 source.n226 source.n225 9.3005
R592 source.n177 source.n176 9.3005
R593 source.n220 source.n219 9.3005
R594 source.n218 source.n217 9.3005
R595 source.n496 source.n495 8.92171
R596 source.n529 source.n470 8.92171
R597 source.n542 source.n462 8.92171
R598 source.n576 source.n575 8.92171
R599 source.n350 source.n349 8.92171
R600 source.n383 source.n324 8.92171
R601 source.n396 source.n316 8.92171
R602 source.n430 source.n429 8.92171
R603 source.n132 source.n131 8.92171
R604 source.n99 source.n19 8.92171
R605 source.n86 source.n27 8.92171
R606 source.n54 source.n53 8.92171
R607 source.n278 source.n277 8.92171
R608 source.n245 source.n165 8.92171
R609 source.n232 source.n173 8.92171
R610 source.n200 source.n199 8.92171
R611 source.n492 source.n486 8.14595
R612 source.n530 source.n468 8.14595
R613 source.n541 source.n464 8.14595
R614 source.n579 source.n446 8.14595
R615 source.n346 source.n340 8.14595
R616 source.n384 source.n322 8.14595
R617 source.n395 source.n318 8.14595
R618 source.n433 source.n300 8.14595
R619 source.n135 source.n2 8.14595
R620 source.n98 source.n21 8.14595
R621 source.n87 source.n25 8.14595
R622 source.n50 source.n44 8.14595
R623 source.n281 source.n148 8.14595
R624 source.n244 source.n167 8.14595
R625 source.n233 source.n171 8.14595
R626 source.n196 source.n190 8.14595
R627 source.n491 source.n488 7.3702
R628 source.n534 source.n533 7.3702
R629 source.n538 source.n537 7.3702
R630 source.n580 source.n444 7.3702
R631 source.n345 source.n342 7.3702
R632 source.n388 source.n387 7.3702
R633 source.n392 source.n391 7.3702
R634 source.n434 source.n298 7.3702
R635 source.n136 source.n0 7.3702
R636 source.n95 source.n94 7.3702
R637 source.n91 source.n90 7.3702
R638 source.n49 source.n46 7.3702
R639 source.n282 source.n146 7.3702
R640 source.n241 source.n240 7.3702
R641 source.n237 source.n236 7.3702
R642 source.n195 source.n192 7.3702
R643 source.n534 source.n466 6.59444
R644 source.n537 source.n466 6.59444
R645 source.n582 source.n444 6.59444
R646 source.n388 source.n320 6.59444
R647 source.n391 source.n320 6.59444
R648 source.n436 source.n298 6.59444
R649 source.n138 source.n0 6.59444
R650 source.n94 source.n23 6.59444
R651 source.n91 source.n23 6.59444
R652 source.n284 source.n146 6.59444
R653 source.n240 source.n169 6.59444
R654 source.n237 source.n169 6.59444
R655 source.n492 source.n491 5.81868
R656 source.n533 source.n468 5.81868
R657 source.n538 source.n464 5.81868
R658 source.n580 source.n579 5.81868
R659 source.n346 source.n345 5.81868
R660 source.n387 source.n322 5.81868
R661 source.n392 source.n318 5.81868
R662 source.n434 source.n433 5.81868
R663 source.n136 source.n135 5.81868
R664 source.n95 source.n21 5.81868
R665 source.n90 source.n25 5.81868
R666 source.n50 source.n49 5.81868
R667 source.n282 source.n281 5.81868
R668 source.n241 source.n167 5.81868
R669 source.n236 source.n171 5.81868
R670 source.n196 source.n195 5.81868
R671 source.n584 source.n583 5.62119
R672 source.n495 source.n486 5.04292
R673 source.n530 source.n529 5.04292
R674 source.n542 source.n541 5.04292
R675 source.n576 source.n446 5.04292
R676 source.n349 source.n340 5.04292
R677 source.n384 source.n383 5.04292
R678 source.n396 source.n395 5.04292
R679 source.n430 source.n300 5.04292
R680 source.n132 source.n2 5.04292
R681 source.n99 source.n98 5.04292
R682 source.n87 source.n86 5.04292
R683 source.n53 source.n44 5.04292
R684 source.n278 source.n148 5.04292
R685 source.n245 source.n244 5.04292
R686 source.n233 source.n232 5.04292
R687 source.n199 source.n190 5.04292
R688 source.n496 source.n484 4.26717
R689 source.n526 source.n470 4.26717
R690 source.n545 source.n462 4.26717
R691 source.n575 source.n448 4.26717
R692 source.n350 source.n338 4.26717
R693 source.n380 source.n324 4.26717
R694 source.n399 source.n316 4.26717
R695 source.n429 source.n302 4.26717
R696 source.n131 source.n4 4.26717
R697 source.n102 source.n19 4.26717
R698 source.n83 source.n27 4.26717
R699 source.n54 source.n42 4.26717
R700 source.n277 source.n150 4.26717
R701 source.n248 source.n165 4.26717
R702 source.n229 source.n173 4.26717
R703 source.n200 source.n188 4.26717
R704 source.n500 source.n499 3.49141
R705 source.n525 source.n472 3.49141
R706 source.n546 source.n460 3.49141
R707 source.n572 source.n571 3.49141
R708 source.n354 source.n353 3.49141
R709 source.n379 source.n326 3.49141
R710 source.n400 source.n314 3.49141
R711 source.n426 source.n425 3.49141
R712 source.n128 source.n127 3.49141
R713 source.n103 source.n17 3.49141
R714 source.n82 source.n29 3.49141
R715 source.n58 source.n57 3.49141
R716 source.n274 source.n273 3.49141
R717 source.n249 source.n163 3.49141
R718 source.n228 source.n175 3.49141
R719 source.n204 source.n203 3.49141
R720 source.n48 source.n47 2.84303
R721 source.n194 source.n193 2.84303
R722 source.n490 source.n489 2.84303
R723 source.n344 source.n343 2.84303
R724 source.n503 source.n482 2.71565
R725 source.n522 source.n521 2.71565
R726 source.n550 source.n549 2.71565
R727 source.n568 source.n450 2.71565
R728 source.n357 source.n336 2.71565
R729 source.n376 source.n375 2.71565
R730 source.n404 source.n403 2.71565
R731 source.n422 source.n304 2.71565
R732 source.n124 source.n6 2.71565
R733 source.n107 source.n106 2.71565
R734 source.n79 source.n78 2.71565
R735 source.n61 source.n40 2.71565
R736 source.n270 source.n152 2.71565
R737 source.n253 source.n252 2.71565
R738 source.n225 source.n224 2.71565
R739 source.n207 source.n186 2.71565
R740 source.n504 source.n480 1.93989
R741 source.n518 source.n474 1.93989
R742 source.n554 source.n458 1.93989
R743 source.n567 source.n452 1.93989
R744 source.n358 source.n334 1.93989
R745 source.n372 source.n328 1.93989
R746 source.n408 source.n312 1.93989
R747 source.n421 source.n306 1.93989
R748 source.n123 source.n8 1.93989
R749 source.n110 source.n14 1.93989
R750 source.n75 source.n31 1.93989
R751 source.n62 source.n38 1.93989
R752 source.n269 source.n154 1.93989
R753 source.n256 source.n160 1.93989
R754 source.n221 source.n177 1.93989
R755 source.n208 source.n184 1.93989
R756 source.n509 source.n507 1.16414
R757 source.n517 source.n476 1.16414
R758 source.n555 source.n456 1.16414
R759 source.n564 source.n563 1.16414
R760 source.n363 source.n361 1.16414
R761 source.n371 source.n330 1.16414
R762 source.n409 source.n310 1.16414
R763 source.n418 source.n417 1.16414
R764 source.n120 source.n119 1.16414
R765 source.n111 source.n12 1.16414
R766 source.n74 source.n33 1.16414
R767 source.n66 source.n65 1.16414
R768 source.n266 source.n265 1.16414
R769 source.n257 source.n158 1.16414
R770 source.n220 source.n179 1.16414
R771 source.n212 source.n211 1.16414
R772 source.n285 source.n145 0.828086
R773 source.n439 source.n437 0.828086
R774 source.n442 source.t17 0.7925
R775 source.n442 source.t25 0.7925
R776 source.n440 source.t23 0.7925
R777 source.n440 source.t24 0.7925
R778 source.n438 source.t20 0.7925
R779 source.n438 source.t26 0.7925
R780 source.n296 source.t10 0.7925
R781 source.n296 source.t3 0.7925
R782 source.n294 source.t4 0.7925
R783 source.n294 source.t12 0.7925
R784 source.n292 source.t2 0.7925
R785 source.n292 source.t6 0.7925
R786 source.n140 source.t0 0.7925
R787 source.n140 source.t11 0.7925
R788 source.n142 source.t8 0.7925
R789 source.n142 source.t7 0.7925
R790 source.n144 source.t13 0.7925
R791 source.n144 source.t9 0.7925
R792 source.n286 source.t15 0.7925
R793 source.n286 source.t18 0.7925
R794 source.n288 source.t19 0.7925
R795 source.n288 source.t16 0.7925
R796 source.n290 source.t27 0.7925
R797 source.n290 source.t14 0.7925
R798 source.n291 source.n289 0.716017
R799 source.n289 source.n287 0.716017
R800 source.n287 source.n285 0.716017
R801 source.n145 source.n143 0.716017
R802 source.n143 source.n141 0.716017
R803 source.n141 source.n139 0.716017
R804 source.n295 source.n293 0.716017
R805 source.n297 source.n295 0.716017
R806 source.n437 source.n297 0.716017
R807 source.n441 source.n439 0.716017
R808 source.n443 source.n441 0.716017
R809 source.n583 source.n443 0.716017
R810 source.n508 source.n478 0.388379
R811 source.n514 source.n513 0.388379
R812 source.n559 source.n558 0.388379
R813 source.n560 source.n454 0.388379
R814 source.n362 source.n332 0.388379
R815 source.n368 source.n367 0.388379
R816 source.n413 source.n412 0.388379
R817 source.n414 source.n308 0.388379
R818 source.n116 source.n10 0.388379
R819 source.n115 source.n114 0.388379
R820 source.n71 source.n70 0.388379
R821 source.n37 source.n35 0.388379
R822 source.n262 source.n156 0.388379
R823 source.n261 source.n260 0.388379
R824 source.n217 source.n216 0.388379
R825 source.n183 source.n181 0.388379
R826 source source.n584 0.188
R827 source.n490 source.n485 0.155672
R828 source.n497 source.n485 0.155672
R829 source.n498 source.n497 0.155672
R830 source.n498 source.n481 0.155672
R831 source.n505 source.n481 0.155672
R832 source.n506 source.n505 0.155672
R833 source.n506 source.n477 0.155672
R834 source.n515 source.n477 0.155672
R835 source.n516 source.n515 0.155672
R836 source.n516 source.n473 0.155672
R837 source.n523 source.n473 0.155672
R838 source.n524 source.n523 0.155672
R839 source.n524 source.n469 0.155672
R840 source.n531 source.n469 0.155672
R841 source.n532 source.n531 0.155672
R842 source.n532 source.n465 0.155672
R843 source.n539 source.n465 0.155672
R844 source.n540 source.n539 0.155672
R845 source.n540 source.n461 0.155672
R846 source.n547 source.n461 0.155672
R847 source.n548 source.n547 0.155672
R848 source.n548 source.n457 0.155672
R849 source.n556 source.n457 0.155672
R850 source.n557 source.n556 0.155672
R851 source.n557 source.n453 0.155672
R852 source.n565 source.n453 0.155672
R853 source.n566 source.n565 0.155672
R854 source.n566 source.n449 0.155672
R855 source.n573 source.n449 0.155672
R856 source.n574 source.n573 0.155672
R857 source.n574 source.n445 0.155672
R858 source.n581 source.n445 0.155672
R859 source.n344 source.n339 0.155672
R860 source.n351 source.n339 0.155672
R861 source.n352 source.n351 0.155672
R862 source.n352 source.n335 0.155672
R863 source.n359 source.n335 0.155672
R864 source.n360 source.n359 0.155672
R865 source.n360 source.n331 0.155672
R866 source.n369 source.n331 0.155672
R867 source.n370 source.n369 0.155672
R868 source.n370 source.n327 0.155672
R869 source.n377 source.n327 0.155672
R870 source.n378 source.n377 0.155672
R871 source.n378 source.n323 0.155672
R872 source.n385 source.n323 0.155672
R873 source.n386 source.n385 0.155672
R874 source.n386 source.n319 0.155672
R875 source.n393 source.n319 0.155672
R876 source.n394 source.n393 0.155672
R877 source.n394 source.n315 0.155672
R878 source.n401 source.n315 0.155672
R879 source.n402 source.n401 0.155672
R880 source.n402 source.n311 0.155672
R881 source.n410 source.n311 0.155672
R882 source.n411 source.n410 0.155672
R883 source.n411 source.n307 0.155672
R884 source.n419 source.n307 0.155672
R885 source.n420 source.n419 0.155672
R886 source.n420 source.n303 0.155672
R887 source.n427 source.n303 0.155672
R888 source.n428 source.n427 0.155672
R889 source.n428 source.n299 0.155672
R890 source.n435 source.n299 0.155672
R891 source.n137 source.n1 0.155672
R892 source.n130 source.n1 0.155672
R893 source.n130 source.n129 0.155672
R894 source.n129 source.n5 0.155672
R895 source.n122 source.n5 0.155672
R896 source.n122 source.n121 0.155672
R897 source.n121 source.n9 0.155672
R898 source.n113 source.n9 0.155672
R899 source.n113 source.n112 0.155672
R900 source.n112 source.n13 0.155672
R901 source.n105 source.n13 0.155672
R902 source.n105 source.n104 0.155672
R903 source.n104 source.n18 0.155672
R904 source.n97 source.n18 0.155672
R905 source.n97 source.n96 0.155672
R906 source.n96 source.n22 0.155672
R907 source.n89 source.n22 0.155672
R908 source.n89 source.n88 0.155672
R909 source.n88 source.n26 0.155672
R910 source.n81 source.n26 0.155672
R911 source.n81 source.n80 0.155672
R912 source.n80 source.n30 0.155672
R913 source.n73 source.n30 0.155672
R914 source.n73 source.n72 0.155672
R915 source.n72 source.n34 0.155672
R916 source.n64 source.n34 0.155672
R917 source.n64 source.n63 0.155672
R918 source.n63 source.n39 0.155672
R919 source.n56 source.n39 0.155672
R920 source.n56 source.n55 0.155672
R921 source.n55 source.n43 0.155672
R922 source.n48 source.n43 0.155672
R923 source.n283 source.n147 0.155672
R924 source.n276 source.n147 0.155672
R925 source.n276 source.n275 0.155672
R926 source.n275 source.n151 0.155672
R927 source.n268 source.n151 0.155672
R928 source.n268 source.n267 0.155672
R929 source.n267 source.n155 0.155672
R930 source.n259 source.n155 0.155672
R931 source.n259 source.n258 0.155672
R932 source.n258 source.n159 0.155672
R933 source.n251 source.n159 0.155672
R934 source.n251 source.n250 0.155672
R935 source.n250 source.n164 0.155672
R936 source.n243 source.n164 0.155672
R937 source.n243 source.n242 0.155672
R938 source.n242 source.n168 0.155672
R939 source.n235 source.n168 0.155672
R940 source.n235 source.n234 0.155672
R941 source.n234 source.n172 0.155672
R942 source.n227 source.n172 0.155672
R943 source.n227 source.n226 0.155672
R944 source.n226 source.n176 0.155672
R945 source.n219 source.n176 0.155672
R946 source.n219 source.n218 0.155672
R947 source.n218 source.n180 0.155672
R948 source.n210 source.n180 0.155672
R949 source.n210 source.n209 0.155672
R950 source.n209 source.n185 0.155672
R951 source.n202 source.n185 0.155672
R952 source.n202 source.n201 0.155672
R953 source.n201 source.n189 0.155672
R954 source.n194 source.n189 0.155672
R955 drain_right.n134 drain_right.n0 289.615
R956 drain_right.n284 drain_right.n150 289.615
R957 drain_right.n44 drain_right.n43 185
R958 drain_right.n49 drain_right.n48 185
R959 drain_right.n51 drain_right.n50 185
R960 drain_right.n40 drain_right.n39 185
R961 drain_right.n57 drain_right.n56 185
R962 drain_right.n59 drain_right.n58 185
R963 drain_right.n36 drain_right.n35 185
R964 drain_right.n66 drain_right.n65 185
R965 drain_right.n67 drain_right.n34 185
R966 drain_right.n69 drain_right.n68 185
R967 drain_right.n32 drain_right.n31 185
R968 drain_right.n75 drain_right.n74 185
R969 drain_right.n77 drain_right.n76 185
R970 drain_right.n28 drain_right.n27 185
R971 drain_right.n83 drain_right.n82 185
R972 drain_right.n85 drain_right.n84 185
R973 drain_right.n24 drain_right.n23 185
R974 drain_right.n91 drain_right.n90 185
R975 drain_right.n93 drain_right.n92 185
R976 drain_right.n20 drain_right.n19 185
R977 drain_right.n99 drain_right.n98 185
R978 drain_right.n101 drain_right.n100 185
R979 drain_right.n16 drain_right.n15 185
R980 drain_right.n107 drain_right.n106 185
R981 drain_right.n110 drain_right.n109 185
R982 drain_right.n108 drain_right.n12 185
R983 drain_right.n115 drain_right.n11 185
R984 drain_right.n117 drain_right.n116 185
R985 drain_right.n119 drain_right.n118 185
R986 drain_right.n8 drain_right.n7 185
R987 drain_right.n125 drain_right.n124 185
R988 drain_right.n127 drain_right.n126 185
R989 drain_right.n4 drain_right.n3 185
R990 drain_right.n133 drain_right.n132 185
R991 drain_right.n135 drain_right.n134 185
R992 drain_right.n285 drain_right.n284 185
R993 drain_right.n283 drain_right.n282 185
R994 drain_right.n154 drain_right.n153 185
R995 drain_right.n277 drain_right.n276 185
R996 drain_right.n275 drain_right.n274 185
R997 drain_right.n158 drain_right.n157 185
R998 drain_right.n269 drain_right.n268 185
R999 drain_right.n267 drain_right.n266 185
R1000 drain_right.n265 drain_right.n161 185
R1001 drain_right.n165 drain_right.n162 185
R1002 drain_right.n260 drain_right.n259 185
R1003 drain_right.n258 drain_right.n257 185
R1004 drain_right.n167 drain_right.n166 185
R1005 drain_right.n252 drain_right.n251 185
R1006 drain_right.n250 drain_right.n249 185
R1007 drain_right.n171 drain_right.n170 185
R1008 drain_right.n244 drain_right.n243 185
R1009 drain_right.n242 drain_right.n241 185
R1010 drain_right.n175 drain_right.n174 185
R1011 drain_right.n236 drain_right.n235 185
R1012 drain_right.n234 drain_right.n233 185
R1013 drain_right.n179 drain_right.n178 185
R1014 drain_right.n228 drain_right.n227 185
R1015 drain_right.n226 drain_right.n225 185
R1016 drain_right.n183 drain_right.n182 185
R1017 drain_right.n220 drain_right.n219 185
R1018 drain_right.n218 drain_right.n185 185
R1019 drain_right.n217 drain_right.n216 185
R1020 drain_right.n188 drain_right.n186 185
R1021 drain_right.n211 drain_right.n210 185
R1022 drain_right.n209 drain_right.n208 185
R1023 drain_right.n192 drain_right.n191 185
R1024 drain_right.n203 drain_right.n202 185
R1025 drain_right.n201 drain_right.n200 185
R1026 drain_right.n196 drain_right.n195 185
R1027 drain_right.n45 drain_right.t10 149.524
R1028 drain_right.n197 drain_right.t13 149.524
R1029 drain_right.n49 drain_right.n43 104.615
R1030 drain_right.n50 drain_right.n49 104.615
R1031 drain_right.n50 drain_right.n39 104.615
R1032 drain_right.n57 drain_right.n39 104.615
R1033 drain_right.n58 drain_right.n57 104.615
R1034 drain_right.n58 drain_right.n35 104.615
R1035 drain_right.n66 drain_right.n35 104.615
R1036 drain_right.n67 drain_right.n66 104.615
R1037 drain_right.n68 drain_right.n67 104.615
R1038 drain_right.n68 drain_right.n31 104.615
R1039 drain_right.n75 drain_right.n31 104.615
R1040 drain_right.n76 drain_right.n75 104.615
R1041 drain_right.n76 drain_right.n27 104.615
R1042 drain_right.n83 drain_right.n27 104.615
R1043 drain_right.n84 drain_right.n83 104.615
R1044 drain_right.n84 drain_right.n23 104.615
R1045 drain_right.n91 drain_right.n23 104.615
R1046 drain_right.n92 drain_right.n91 104.615
R1047 drain_right.n92 drain_right.n19 104.615
R1048 drain_right.n99 drain_right.n19 104.615
R1049 drain_right.n100 drain_right.n99 104.615
R1050 drain_right.n100 drain_right.n15 104.615
R1051 drain_right.n107 drain_right.n15 104.615
R1052 drain_right.n109 drain_right.n107 104.615
R1053 drain_right.n109 drain_right.n108 104.615
R1054 drain_right.n108 drain_right.n11 104.615
R1055 drain_right.n117 drain_right.n11 104.615
R1056 drain_right.n118 drain_right.n117 104.615
R1057 drain_right.n118 drain_right.n7 104.615
R1058 drain_right.n125 drain_right.n7 104.615
R1059 drain_right.n126 drain_right.n125 104.615
R1060 drain_right.n126 drain_right.n3 104.615
R1061 drain_right.n133 drain_right.n3 104.615
R1062 drain_right.n134 drain_right.n133 104.615
R1063 drain_right.n284 drain_right.n283 104.615
R1064 drain_right.n283 drain_right.n153 104.615
R1065 drain_right.n276 drain_right.n153 104.615
R1066 drain_right.n276 drain_right.n275 104.615
R1067 drain_right.n275 drain_right.n157 104.615
R1068 drain_right.n268 drain_right.n157 104.615
R1069 drain_right.n268 drain_right.n267 104.615
R1070 drain_right.n267 drain_right.n161 104.615
R1071 drain_right.n165 drain_right.n161 104.615
R1072 drain_right.n259 drain_right.n165 104.615
R1073 drain_right.n259 drain_right.n258 104.615
R1074 drain_right.n258 drain_right.n166 104.615
R1075 drain_right.n251 drain_right.n166 104.615
R1076 drain_right.n251 drain_right.n250 104.615
R1077 drain_right.n250 drain_right.n170 104.615
R1078 drain_right.n243 drain_right.n170 104.615
R1079 drain_right.n243 drain_right.n242 104.615
R1080 drain_right.n242 drain_right.n174 104.615
R1081 drain_right.n235 drain_right.n174 104.615
R1082 drain_right.n235 drain_right.n234 104.615
R1083 drain_right.n234 drain_right.n178 104.615
R1084 drain_right.n227 drain_right.n178 104.615
R1085 drain_right.n227 drain_right.n226 104.615
R1086 drain_right.n226 drain_right.n182 104.615
R1087 drain_right.n219 drain_right.n182 104.615
R1088 drain_right.n219 drain_right.n218 104.615
R1089 drain_right.n218 drain_right.n217 104.615
R1090 drain_right.n217 drain_right.n186 104.615
R1091 drain_right.n210 drain_right.n186 104.615
R1092 drain_right.n210 drain_right.n209 104.615
R1093 drain_right.n209 drain_right.n191 104.615
R1094 drain_right.n202 drain_right.n191 104.615
R1095 drain_right.n202 drain_right.n201 104.615
R1096 drain_right.n201 drain_right.n195 104.615
R1097 drain_right.n143 drain_right.n141 59.431
R1098 drain_right.n147 drain_right.n145 59.4308
R1099 drain_right.n143 drain_right.n142 58.7154
R1100 drain_right.n140 drain_right.n139 58.7154
R1101 drain_right.n147 drain_right.n146 58.7154
R1102 drain_right.n149 drain_right.n148 58.7154
R1103 drain_right.t10 drain_right.n43 52.3082
R1104 drain_right.t13 drain_right.n195 52.3082
R1105 drain_right.n140 drain_right.n138 48.0281
R1106 drain_right.n289 drain_right.n288 47.3126
R1107 drain_right drain_right.n144 40.7766
R1108 drain_right.n69 drain_right.n34 13.1884
R1109 drain_right.n116 drain_right.n115 13.1884
R1110 drain_right.n266 drain_right.n265 13.1884
R1111 drain_right.n220 drain_right.n185 13.1884
R1112 drain_right.n65 drain_right.n64 12.8005
R1113 drain_right.n70 drain_right.n32 12.8005
R1114 drain_right.n114 drain_right.n12 12.8005
R1115 drain_right.n119 drain_right.n10 12.8005
R1116 drain_right.n269 drain_right.n160 12.8005
R1117 drain_right.n264 drain_right.n162 12.8005
R1118 drain_right.n221 drain_right.n183 12.8005
R1119 drain_right.n216 drain_right.n187 12.8005
R1120 drain_right.n63 drain_right.n36 12.0247
R1121 drain_right.n74 drain_right.n73 12.0247
R1122 drain_right.n111 drain_right.n110 12.0247
R1123 drain_right.n120 drain_right.n8 12.0247
R1124 drain_right.n270 drain_right.n158 12.0247
R1125 drain_right.n261 drain_right.n260 12.0247
R1126 drain_right.n225 drain_right.n224 12.0247
R1127 drain_right.n215 drain_right.n188 12.0247
R1128 drain_right.n60 drain_right.n59 11.249
R1129 drain_right.n77 drain_right.n30 11.249
R1130 drain_right.n106 drain_right.n14 11.249
R1131 drain_right.n124 drain_right.n123 11.249
R1132 drain_right.n274 drain_right.n273 11.249
R1133 drain_right.n257 drain_right.n164 11.249
R1134 drain_right.n228 drain_right.n181 11.249
R1135 drain_right.n212 drain_right.n211 11.249
R1136 drain_right.n56 drain_right.n38 10.4732
R1137 drain_right.n78 drain_right.n28 10.4732
R1138 drain_right.n105 drain_right.n16 10.4732
R1139 drain_right.n127 drain_right.n6 10.4732
R1140 drain_right.n277 drain_right.n156 10.4732
R1141 drain_right.n256 drain_right.n167 10.4732
R1142 drain_right.n229 drain_right.n179 10.4732
R1143 drain_right.n208 drain_right.n190 10.4732
R1144 drain_right.n45 drain_right.n44 10.2747
R1145 drain_right.n197 drain_right.n196 10.2747
R1146 drain_right.n55 drain_right.n40 9.69747
R1147 drain_right.n82 drain_right.n81 9.69747
R1148 drain_right.n102 drain_right.n101 9.69747
R1149 drain_right.n128 drain_right.n4 9.69747
R1150 drain_right.n278 drain_right.n154 9.69747
R1151 drain_right.n253 drain_right.n252 9.69747
R1152 drain_right.n233 drain_right.n232 9.69747
R1153 drain_right.n207 drain_right.n192 9.69747
R1154 drain_right.n138 drain_right.n137 9.45567
R1155 drain_right.n288 drain_right.n287 9.45567
R1156 drain_right.n2 drain_right.n1 9.3005
R1157 drain_right.n131 drain_right.n130 9.3005
R1158 drain_right.n129 drain_right.n128 9.3005
R1159 drain_right.n6 drain_right.n5 9.3005
R1160 drain_right.n123 drain_right.n122 9.3005
R1161 drain_right.n121 drain_right.n120 9.3005
R1162 drain_right.n10 drain_right.n9 9.3005
R1163 drain_right.n89 drain_right.n88 9.3005
R1164 drain_right.n87 drain_right.n86 9.3005
R1165 drain_right.n26 drain_right.n25 9.3005
R1166 drain_right.n81 drain_right.n80 9.3005
R1167 drain_right.n79 drain_right.n78 9.3005
R1168 drain_right.n30 drain_right.n29 9.3005
R1169 drain_right.n73 drain_right.n72 9.3005
R1170 drain_right.n71 drain_right.n70 9.3005
R1171 drain_right.n47 drain_right.n46 9.3005
R1172 drain_right.n42 drain_right.n41 9.3005
R1173 drain_right.n53 drain_right.n52 9.3005
R1174 drain_right.n55 drain_right.n54 9.3005
R1175 drain_right.n38 drain_right.n37 9.3005
R1176 drain_right.n61 drain_right.n60 9.3005
R1177 drain_right.n63 drain_right.n62 9.3005
R1178 drain_right.n64 drain_right.n33 9.3005
R1179 drain_right.n22 drain_right.n21 9.3005
R1180 drain_right.n95 drain_right.n94 9.3005
R1181 drain_right.n97 drain_right.n96 9.3005
R1182 drain_right.n18 drain_right.n17 9.3005
R1183 drain_right.n103 drain_right.n102 9.3005
R1184 drain_right.n105 drain_right.n104 9.3005
R1185 drain_right.n14 drain_right.n13 9.3005
R1186 drain_right.n112 drain_right.n111 9.3005
R1187 drain_right.n114 drain_right.n113 9.3005
R1188 drain_right.n137 drain_right.n136 9.3005
R1189 drain_right.n199 drain_right.n198 9.3005
R1190 drain_right.n194 drain_right.n193 9.3005
R1191 drain_right.n205 drain_right.n204 9.3005
R1192 drain_right.n207 drain_right.n206 9.3005
R1193 drain_right.n190 drain_right.n189 9.3005
R1194 drain_right.n213 drain_right.n212 9.3005
R1195 drain_right.n215 drain_right.n214 9.3005
R1196 drain_right.n187 drain_right.n184 9.3005
R1197 drain_right.n246 drain_right.n245 9.3005
R1198 drain_right.n248 drain_right.n247 9.3005
R1199 drain_right.n169 drain_right.n168 9.3005
R1200 drain_right.n254 drain_right.n253 9.3005
R1201 drain_right.n256 drain_right.n255 9.3005
R1202 drain_right.n164 drain_right.n163 9.3005
R1203 drain_right.n262 drain_right.n261 9.3005
R1204 drain_right.n264 drain_right.n263 9.3005
R1205 drain_right.n287 drain_right.n286 9.3005
R1206 drain_right.n152 drain_right.n151 9.3005
R1207 drain_right.n281 drain_right.n280 9.3005
R1208 drain_right.n279 drain_right.n278 9.3005
R1209 drain_right.n156 drain_right.n155 9.3005
R1210 drain_right.n273 drain_right.n272 9.3005
R1211 drain_right.n271 drain_right.n270 9.3005
R1212 drain_right.n160 drain_right.n159 9.3005
R1213 drain_right.n173 drain_right.n172 9.3005
R1214 drain_right.n240 drain_right.n239 9.3005
R1215 drain_right.n238 drain_right.n237 9.3005
R1216 drain_right.n177 drain_right.n176 9.3005
R1217 drain_right.n232 drain_right.n231 9.3005
R1218 drain_right.n230 drain_right.n229 9.3005
R1219 drain_right.n181 drain_right.n180 9.3005
R1220 drain_right.n224 drain_right.n223 9.3005
R1221 drain_right.n222 drain_right.n221 9.3005
R1222 drain_right.n52 drain_right.n51 8.92171
R1223 drain_right.n85 drain_right.n26 8.92171
R1224 drain_right.n98 drain_right.n18 8.92171
R1225 drain_right.n132 drain_right.n131 8.92171
R1226 drain_right.n282 drain_right.n281 8.92171
R1227 drain_right.n249 drain_right.n169 8.92171
R1228 drain_right.n236 drain_right.n177 8.92171
R1229 drain_right.n204 drain_right.n203 8.92171
R1230 drain_right.n48 drain_right.n42 8.14595
R1231 drain_right.n86 drain_right.n24 8.14595
R1232 drain_right.n97 drain_right.n20 8.14595
R1233 drain_right.n135 drain_right.n2 8.14595
R1234 drain_right.n285 drain_right.n152 8.14595
R1235 drain_right.n248 drain_right.n171 8.14595
R1236 drain_right.n237 drain_right.n175 8.14595
R1237 drain_right.n200 drain_right.n194 8.14595
R1238 drain_right.n47 drain_right.n44 7.3702
R1239 drain_right.n90 drain_right.n89 7.3702
R1240 drain_right.n94 drain_right.n93 7.3702
R1241 drain_right.n136 drain_right.n0 7.3702
R1242 drain_right.n286 drain_right.n150 7.3702
R1243 drain_right.n245 drain_right.n244 7.3702
R1244 drain_right.n241 drain_right.n240 7.3702
R1245 drain_right.n199 drain_right.n196 7.3702
R1246 drain_right.n90 drain_right.n22 6.59444
R1247 drain_right.n93 drain_right.n22 6.59444
R1248 drain_right.n138 drain_right.n0 6.59444
R1249 drain_right.n288 drain_right.n150 6.59444
R1250 drain_right.n244 drain_right.n173 6.59444
R1251 drain_right.n241 drain_right.n173 6.59444
R1252 drain_right drain_right.n289 6.01097
R1253 drain_right.n48 drain_right.n47 5.81868
R1254 drain_right.n89 drain_right.n24 5.81868
R1255 drain_right.n94 drain_right.n20 5.81868
R1256 drain_right.n136 drain_right.n135 5.81868
R1257 drain_right.n286 drain_right.n285 5.81868
R1258 drain_right.n245 drain_right.n171 5.81868
R1259 drain_right.n240 drain_right.n175 5.81868
R1260 drain_right.n200 drain_right.n199 5.81868
R1261 drain_right.n51 drain_right.n42 5.04292
R1262 drain_right.n86 drain_right.n85 5.04292
R1263 drain_right.n98 drain_right.n97 5.04292
R1264 drain_right.n132 drain_right.n2 5.04292
R1265 drain_right.n282 drain_right.n152 5.04292
R1266 drain_right.n249 drain_right.n248 5.04292
R1267 drain_right.n237 drain_right.n236 5.04292
R1268 drain_right.n203 drain_right.n194 5.04292
R1269 drain_right.n52 drain_right.n40 4.26717
R1270 drain_right.n82 drain_right.n26 4.26717
R1271 drain_right.n101 drain_right.n18 4.26717
R1272 drain_right.n131 drain_right.n4 4.26717
R1273 drain_right.n281 drain_right.n154 4.26717
R1274 drain_right.n252 drain_right.n169 4.26717
R1275 drain_right.n233 drain_right.n177 4.26717
R1276 drain_right.n204 drain_right.n192 4.26717
R1277 drain_right.n56 drain_right.n55 3.49141
R1278 drain_right.n81 drain_right.n28 3.49141
R1279 drain_right.n102 drain_right.n16 3.49141
R1280 drain_right.n128 drain_right.n127 3.49141
R1281 drain_right.n278 drain_right.n277 3.49141
R1282 drain_right.n253 drain_right.n167 3.49141
R1283 drain_right.n232 drain_right.n179 3.49141
R1284 drain_right.n208 drain_right.n207 3.49141
R1285 drain_right.n198 drain_right.n197 2.84303
R1286 drain_right.n46 drain_right.n45 2.84303
R1287 drain_right.n59 drain_right.n38 2.71565
R1288 drain_right.n78 drain_right.n77 2.71565
R1289 drain_right.n106 drain_right.n105 2.71565
R1290 drain_right.n124 drain_right.n6 2.71565
R1291 drain_right.n274 drain_right.n156 2.71565
R1292 drain_right.n257 drain_right.n256 2.71565
R1293 drain_right.n229 drain_right.n228 2.71565
R1294 drain_right.n211 drain_right.n190 2.71565
R1295 drain_right.n60 drain_right.n36 1.93989
R1296 drain_right.n74 drain_right.n30 1.93989
R1297 drain_right.n110 drain_right.n14 1.93989
R1298 drain_right.n123 drain_right.n8 1.93989
R1299 drain_right.n273 drain_right.n158 1.93989
R1300 drain_right.n260 drain_right.n164 1.93989
R1301 drain_right.n225 drain_right.n181 1.93989
R1302 drain_right.n212 drain_right.n188 1.93989
R1303 drain_right.n65 drain_right.n63 1.16414
R1304 drain_right.n73 drain_right.n32 1.16414
R1305 drain_right.n111 drain_right.n12 1.16414
R1306 drain_right.n120 drain_right.n119 1.16414
R1307 drain_right.n270 drain_right.n269 1.16414
R1308 drain_right.n261 drain_right.n162 1.16414
R1309 drain_right.n224 drain_right.n183 1.16414
R1310 drain_right.n216 drain_right.n215 1.16414
R1311 drain_right.n141 drain_right.t1 0.7925
R1312 drain_right.n141 drain_right.t2 0.7925
R1313 drain_right.n142 drain_right.t5 0.7925
R1314 drain_right.n142 drain_right.t7 0.7925
R1315 drain_right.n139 drain_right.t11 0.7925
R1316 drain_right.n139 drain_right.t4 0.7925
R1317 drain_right.n145 drain_right.t12 0.7925
R1318 drain_right.n145 drain_right.t3 0.7925
R1319 drain_right.n146 drain_right.t0 0.7925
R1320 drain_right.n146 drain_right.t8 0.7925
R1321 drain_right.n148 drain_right.t6 0.7925
R1322 drain_right.n148 drain_right.t9 0.7925
R1323 drain_right.n289 drain_right.n149 0.716017
R1324 drain_right.n149 drain_right.n147 0.716017
R1325 drain_right.n144 drain_right.n140 0.481792
R1326 drain_right.n64 drain_right.n34 0.388379
R1327 drain_right.n70 drain_right.n69 0.388379
R1328 drain_right.n115 drain_right.n114 0.388379
R1329 drain_right.n116 drain_right.n10 0.388379
R1330 drain_right.n266 drain_right.n160 0.388379
R1331 drain_right.n265 drain_right.n264 0.388379
R1332 drain_right.n221 drain_right.n220 0.388379
R1333 drain_right.n187 drain_right.n185 0.388379
R1334 drain_right.n46 drain_right.n41 0.155672
R1335 drain_right.n53 drain_right.n41 0.155672
R1336 drain_right.n54 drain_right.n53 0.155672
R1337 drain_right.n54 drain_right.n37 0.155672
R1338 drain_right.n61 drain_right.n37 0.155672
R1339 drain_right.n62 drain_right.n61 0.155672
R1340 drain_right.n62 drain_right.n33 0.155672
R1341 drain_right.n71 drain_right.n33 0.155672
R1342 drain_right.n72 drain_right.n71 0.155672
R1343 drain_right.n72 drain_right.n29 0.155672
R1344 drain_right.n79 drain_right.n29 0.155672
R1345 drain_right.n80 drain_right.n79 0.155672
R1346 drain_right.n80 drain_right.n25 0.155672
R1347 drain_right.n87 drain_right.n25 0.155672
R1348 drain_right.n88 drain_right.n87 0.155672
R1349 drain_right.n88 drain_right.n21 0.155672
R1350 drain_right.n95 drain_right.n21 0.155672
R1351 drain_right.n96 drain_right.n95 0.155672
R1352 drain_right.n96 drain_right.n17 0.155672
R1353 drain_right.n103 drain_right.n17 0.155672
R1354 drain_right.n104 drain_right.n103 0.155672
R1355 drain_right.n104 drain_right.n13 0.155672
R1356 drain_right.n112 drain_right.n13 0.155672
R1357 drain_right.n113 drain_right.n112 0.155672
R1358 drain_right.n113 drain_right.n9 0.155672
R1359 drain_right.n121 drain_right.n9 0.155672
R1360 drain_right.n122 drain_right.n121 0.155672
R1361 drain_right.n122 drain_right.n5 0.155672
R1362 drain_right.n129 drain_right.n5 0.155672
R1363 drain_right.n130 drain_right.n129 0.155672
R1364 drain_right.n130 drain_right.n1 0.155672
R1365 drain_right.n137 drain_right.n1 0.155672
R1366 drain_right.n287 drain_right.n151 0.155672
R1367 drain_right.n280 drain_right.n151 0.155672
R1368 drain_right.n280 drain_right.n279 0.155672
R1369 drain_right.n279 drain_right.n155 0.155672
R1370 drain_right.n272 drain_right.n155 0.155672
R1371 drain_right.n272 drain_right.n271 0.155672
R1372 drain_right.n271 drain_right.n159 0.155672
R1373 drain_right.n263 drain_right.n159 0.155672
R1374 drain_right.n263 drain_right.n262 0.155672
R1375 drain_right.n262 drain_right.n163 0.155672
R1376 drain_right.n255 drain_right.n163 0.155672
R1377 drain_right.n255 drain_right.n254 0.155672
R1378 drain_right.n254 drain_right.n168 0.155672
R1379 drain_right.n247 drain_right.n168 0.155672
R1380 drain_right.n247 drain_right.n246 0.155672
R1381 drain_right.n246 drain_right.n172 0.155672
R1382 drain_right.n239 drain_right.n172 0.155672
R1383 drain_right.n239 drain_right.n238 0.155672
R1384 drain_right.n238 drain_right.n176 0.155672
R1385 drain_right.n231 drain_right.n176 0.155672
R1386 drain_right.n231 drain_right.n230 0.155672
R1387 drain_right.n230 drain_right.n180 0.155672
R1388 drain_right.n223 drain_right.n180 0.155672
R1389 drain_right.n223 drain_right.n222 0.155672
R1390 drain_right.n222 drain_right.n184 0.155672
R1391 drain_right.n214 drain_right.n184 0.155672
R1392 drain_right.n214 drain_right.n213 0.155672
R1393 drain_right.n213 drain_right.n189 0.155672
R1394 drain_right.n206 drain_right.n189 0.155672
R1395 drain_right.n206 drain_right.n205 0.155672
R1396 drain_right.n205 drain_right.n193 0.155672
R1397 drain_right.n198 drain_right.n193 0.155672
R1398 drain_right.n144 drain_right.n143 0.124033
R1399 plus.n4 plus.t2 1304.55
R1400 plus.n20 plus.t12 1304.55
R1401 plus.n14 plus.t6 1283.57
R1402 plus.n13 plus.t11 1283.57
R1403 plus.n1 plus.t9 1283.57
R1404 plus.n8 plus.t4 1283.57
R1405 plus.n7 plus.t10 1283.57
R1406 plus.n3 plus.t8 1283.57
R1407 plus.n30 plus.t3 1283.57
R1408 plus.n29 plus.t7 1283.57
R1409 plus.n17 plus.t1 1283.57
R1410 plus.n24 plus.t0 1283.57
R1411 plus.n23 plus.t5 1283.57
R1412 plus.n19 plus.t13 1283.57
R1413 plus.n6 plus.n5 161.3
R1414 plus.n7 plus.n2 161.3
R1415 plus.n10 plus.n1 161.3
R1416 plus.n12 plus.n11 161.3
R1417 plus.n13 plus.n0 161.3
R1418 plus.n15 plus.n14 161.3
R1419 plus.n22 plus.n21 161.3
R1420 plus.n23 plus.n18 161.3
R1421 plus.n26 plus.n17 161.3
R1422 plus.n28 plus.n27 161.3
R1423 plus.n29 plus.n16 161.3
R1424 plus.n31 plus.n30 161.3
R1425 plus.n9 plus.n8 80.6037
R1426 plus.n25 plus.n24 80.6037
R1427 plus.n5 plus.n4 70.4033
R1428 plus.n21 plus.n20 70.4033
R1429 plus.n14 plus.n13 48.2005
R1430 plus.n8 plus.n1 48.2005
R1431 plus.n8 plus.n7 48.2005
R1432 plus.n30 plus.n29 48.2005
R1433 plus.n24 plus.n17 48.2005
R1434 plus.n24 plus.n23 48.2005
R1435 plus plus.n31 35.7623
R1436 plus.n12 plus.n1 24.8308
R1437 plus.n7 plus.n6 24.8308
R1438 plus.n28 plus.n17 24.8308
R1439 plus.n23 plus.n22 24.8308
R1440 plus.n13 plus.n12 23.3702
R1441 plus.n6 plus.n3 23.3702
R1442 plus.n29 plus.n28 23.3702
R1443 plus.n22 plus.n19 23.3702
R1444 plus.n4 plus.n3 20.9576
R1445 plus.n20 plus.n19 20.9576
R1446 plus plus.n15 17.1615
R1447 plus.n9 plus.n2 0.285035
R1448 plus.n10 plus.n9 0.285035
R1449 plus.n26 plus.n25 0.285035
R1450 plus.n25 plus.n18 0.285035
R1451 plus.n5 plus.n2 0.189894
R1452 plus.n11 plus.n10 0.189894
R1453 plus.n11 plus.n0 0.189894
R1454 plus.n15 plus.n0 0.189894
R1455 plus.n31 plus.n16 0.189894
R1456 plus.n27 plus.n16 0.189894
R1457 plus.n27 plus.n26 0.189894
R1458 plus.n21 plus.n18 0.189894
R1459 drain_left.n134 drain_left.n0 289.615
R1460 drain_left.n279 drain_left.n145 289.615
R1461 drain_left.n44 drain_left.n43 185
R1462 drain_left.n49 drain_left.n48 185
R1463 drain_left.n51 drain_left.n50 185
R1464 drain_left.n40 drain_left.n39 185
R1465 drain_left.n57 drain_left.n56 185
R1466 drain_left.n59 drain_left.n58 185
R1467 drain_left.n36 drain_left.n35 185
R1468 drain_left.n66 drain_left.n65 185
R1469 drain_left.n67 drain_left.n34 185
R1470 drain_left.n69 drain_left.n68 185
R1471 drain_left.n32 drain_left.n31 185
R1472 drain_left.n75 drain_left.n74 185
R1473 drain_left.n77 drain_left.n76 185
R1474 drain_left.n28 drain_left.n27 185
R1475 drain_left.n83 drain_left.n82 185
R1476 drain_left.n85 drain_left.n84 185
R1477 drain_left.n24 drain_left.n23 185
R1478 drain_left.n91 drain_left.n90 185
R1479 drain_left.n93 drain_left.n92 185
R1480 drain_left.n20 drain_left.n19 185
R1481 drain_left.n99 drain_left.n98 185
R1482 drain_left.n101 drain_left.n100 185
R1483 drain_left.n16 drain_left.n15 185
R1484 drain_left.n107 drain_left.n106 185
R1485 drain_left.n110 drain_left.n109 185
R1486 drain_left.n108 drain_left.n12 185
R1487 drain_left.n115 drain_left.n11 185
R1488 drain_left.n117 drain_left.n116 185
R1489 drain_left.n119 drain_left.n118 185
R1490 drain_left.n8 drain_left.n7 185
R1491 drain_left.n125 drain_left.n124 185
R1492 drain_left.n127 drain_left.n126 185
R1493 drain_left.n4 drain_left.n3 185
R1494 drain_left.n133 drain_left.n132 185
R1495 drain_left.n135 drain_left.n134 185
R1496 drain_left.n280 drain_left.n279 185
R1497 drain_left.n278 drain_left.n277 185
R1498 drain_left.n149 drain_left.n148 185
R1499 drain_left.n272 drain_left.n271 185
R1500 drain_left.n270 drain_left.n269 185
R1501 drain_left.n153 drain_left.n152 185
R1502 drain_left.n264 drain_left.n263 185
R1503 drain_left.n262 drain_left.n261 185
R1504 drain_left.n260 drain_left.n156 185
R1505 drain_left.n160 drain_left.n157 185
R1506 drain_left.n255 drain_left.n254 185
R1507 drain_left.n253 drain_left.n252 185
R1508 drain_left.n162 drain_left.n161 185
R1509 drain_left.n247 drain_left.n246 185
R1510 drain_left.n245 drain_left.n244 185
R1511 drain_left.n166 drain_left.n165 185
R1512 drain_left.n239 drain_left.n238 185
R1513 drain_left.n237 drain_left.n236 185
R1514 drain_left.n170 drain_left.n169 185
R1515 drain_left.n231 drain_left.n230 185
R1516 drain_left.n229 drain_left.n228 185
R1517 drain_left.n174 drain_left.n173 185
R1518 drain_left.n223 drain_left.n222 185
R1519 drain_left.n221 drain_left.n220 185
R1520 drain_left.n178 drain_left.n177 185
R1521 drain_left.n215 drain_left.n214 185
R1522 drain_left.n213 drain_left.n180 185
R1523 drain_left.n212 drain_left.n211 185
R1524 drain_left.n183 drain_left.n181 185
R1525 drain_left.n206 drain_left.n205 185
R1526 drain_left.n204 drain_left.n203 185
R1527 drain_left.n187 drain_left.n186 185
R1528 drain_left.n198 drain_left.n197 185
R1529 drain_left.n196 drain_left.n195 185
R1530 drain_left.n191 drain_left.n190 185
R1531 drain_left.n45 drain_left.t10 149.524
R1532 drain_left.n192 drain_left.t11 149.524
R1533 drain_left.n49 drain_left.n43 104.615
R1534 drain_left.n50 drain_left.n49 104.615
R1535 drain_left.n50 drain_left.n39 104.615
R1536 drain_left.n57 drain_left.n39 104.615
R1537 drain_left.n58 drain_left.n57 104.615
R1538 drain_left.n58 drain_left.n35 104.615
R1539 drain_left.n66 drain_left.n35 104.615
R1540 drain_left.n67 drain_left.n66 104.615
R1541 drain_left.n68 drain_left.n67 104.615
R1542 drain_left.n68 drain_left.n31 104.615
R1543 drain_left.n75 drain_left.n31 104.615
R1544 drain_left.n76 drain_left.n75 104.615
R1545 drain_left.n76 drain_left.n27 104.615
R1546 drain_left.n83 drain_left.n27 104.615
R1547 drain_left.n84 drain_left.n83 104.615
R1548 drain_left.n84 drain_left.n23 104.615
R1549 drain_left.n91 drain_left.n23 104.615
R1550 drain_left.n92 drain_left.n91 104.615
R1551 drain_left.n92 drain_left.n19 104.615
R1552 drain_left.n99 drain_left.n19 104.615
R1553 drain_left.n100 drain_left.n99 104.615
R1554 drain_left.n100 drain_left.n15 104.615
R1555 drain_left.n107 drain_left.n15 104.615
R1556 drain_left.n109 drain_left.n107 104.615
R1557 drain_left.n109 drain_left.n108 104.615
R1558 drain_left.n108 drain_left.n11 104.615
R1559 drain_left.n117 drain_left.n11 104.615
R1560 drain_left.n118 drain_left.n117 104.615
R1561 drain_left.n118 drain_left.n7 104.615
R1562 drain_left.n125 drain_left.n7 104.615
R1563 drain_left.n126 drain_left.n125 104.615
R1564 drain_left.n126 drain_left.n3 104.615
R1565 drain_left.n133 drain_left.n3 104.615
R1566 drain_left.n134 drain_left.n133 104.615
R1567 drain_left.n279 drain_left.n278 104.615
R1568 drain_left.n278 drain_left.n148 104.615
R1569 drain_left.n271 drain_left.n148 104.615
R1570 drain_left.n271 drain_left.n270 104.615
R1571 drain_left.n270 drain_left.n152 104.615
R1572 drain_left.n263 drain_left.n152 104.615
R1573 drain_left.n263 drain_left.n262 104.615
R1574 drain_left.n262 drain_left.n156 104.615
R1575 drain_left.n160 drain_left.n156 104.615
R1576 drain_left.n254 drain_left.n160 104.615
R1577 drain_left.n254 drain_left.n253 104.615
R1578 drain_left.n253 drain_left.n161 104.615
R1579 drain_left.n246 drain_left.n161 104.615
R1580 drain_left.n246 drain_left.n245 104.615
R1581 drain_left.n245 drain_left.n165 104.615
R1582 drain_left.n238 drain_left.n165 104.615
R1583 drain_left.n238 drain_left.n237 104.615
R1584 drain_left.n237 drain_left.n169 104.615
R1585 drain_left.n230 drain_left.n169 104.615
R1586 drain_left.n230 drain_left.n229 104.615
R1587 drain_left.n229 drain_left.n173 104.615
R1588 drain_left.n222 drain_left.n173 104.615
R1589 drain_left.n222 drain_left.n221 104.615
R1590 drain_left.n221 drain_left.n177 104.615
R1591 drain_left.n214 drain_left.n177 104.615
R1592 drain_left.n214 drain_left.n213 104.615
R1593 drain_left.n213 drain_left.n212 104.615
R1594 drain_left.n212 drain_left.n181 104.615
R1595 drain_left.n205 drain_left.n181 104.615
R1596 drain_left.n205 drain_left.n204 104.615
R1597 drain_left.n204 drain_left.n186 104.615
R1598 drain_left.n197 drain_left.n186 104.615
R1599 drain_left.n197 drain_left.n196 104.615
R1600 drain_left.n196 drain_left.n190 104.615
R1601 drain_left.n143 drain_left.n141 59.431
R1602 drain_left.n143 drain_left.n142 58.7154
R1603 drain_left.n140 drain_left.n139 58.7154
R1604 drain_left.n287 drain_left.n286 58.7154
R1605 drain_left.n285 drain_left.n284 58.7154
R1606 drain_left.n289 drain_left.n288 58.7153
R1607 drain_left.t10 drain_left.n43 52.3082
R1608 drain_left.t11 drain_left.n190 52.3082
R1609 drain_left.n140 drain_left.n138 48.0281
R1610 drain_left.n285 drain_left.n283 48.0281
R1611 drain_left drain_left.n144 41.3298
R1612 drain_left.n69 drain_left.n34 13.1884
R1613 drain_left.n116 drain_left.n115 13.1884
R1614 drain_left.n261 drain_left.n260 13.1884
R1615 drain_left.n215 drain_left.n180 13.1884
R1616 drain_left.n65 drain_left.n64 12.8005
R1617 drain_left.n70 drain_left.n32 12.8005
R1618 drain_left.n114 drain_left.n12 12.8005
R1619 drain_left.n119 drain_left.n10 12.8005
R1620 drain_left.n264 drain_left.n155 12.8005
R1621 drain_left.n259 drain_left.n157 12.8005
R1622 drain_left.n216 drain_left.n178 12.8005
R1623 drain_left.n211 drain_left.n182 12.8005
R1624 drain_left.n63 drain_left.n36 12.0247
R1625 drain_left.n74 drain_left.n73 12.0247
R1626 drain_left.n111 drain_left.n110 12.0247
R1627 drain_left.n120 drain_left.n8 12.0247
R1628 drain_left.n265 drain_left.n153 12.0247
R1629 drain_left.n256 drain_left.n255 12.0247
R1630 drain_left.n220 drain_left.n219 12.0247
R1631 drain_left.n210 drain_left.n183 12.0247
R1632 drain_left.n60 drain_left.n59 11.249
R1633 drain_left.n77 drain_left.n30 11.249
R1634 drain_left.n106 drain_left.n14 11.249
R1635 drain_left.n124 drain_left.n123 11.249
R1636 drain_left.n269 drain_left.n268 11.249
R1637 drain_left.n252 drain_left.n159 11.249
R1638 drain_left.n223 drain_left.n176 11.249
R1639 drain_left.n207 drain_left.n206 11.249
R1640 drain_left.n56 drain_left.n38 10.4732
R1641 drain_left.n78 drain_left.n28 10.4732
R1642 drain_left.n105 drain_left.n16 10.4732
R1643 drain_left.n127 drain_left.n6 10.4732
R1644 drain_left.n272 drain_left.n151 10.4732
R1645 drain_left.n251 drain_left.n162 10.4732
R1646 drain_left.n224 drain_left.n174 10.4732
R1647 drain_left.n203 drain_left.n185 10.4732
R1648 drain_left.n45 drain_left.n44 10.2747
R1649 drain_left.n192 drain_left.n191 10.2747
R1650 drain_left.n55 drain_left.n40 9.69747
R1651 drain_left.n82 drain_left.n81 9.69747
R1652 drain_left.n102 drain_left.n101 9.69747
R1653 drain_left.n128 drain_left.n4 9.69747
R1654 drain_left.n273 drain_left.n149 9.69747
R1655 drain_left.n248 drain_left.n247 9.69747
R1656 drain_left.n228 drain_left.n227 9.69747
R1657 drain_left.n202 drain_left.n187 9.69747
R1658 drain_left.n138 drain_left.n137 9.45567
R1659 drain_left.n283 drain_left.n282 9.45567
R1660 drain_left.n2 drain_left.n1 9.3005
R1661 drain_left.n131 drain_left.n130 9.3005
R1662 drain_left.n129 drain_left.n128 9.3005
R1663 drain_left.n6 drain_left.n5 9.3005
R1664 drain_left.n123 drain_left.n122 9.3005
R1665 drain_left.n121 drain_left.n120 9.3005
R1666 drain_left.n10 drain_left.n9 9.3005
R1667 drain_left.n89 drain_left.n88 9.3005
R1668 drain_left.n87 drain_left.n86 9.3005
R1669 drain_left.n26 drain_left.n25 9.3005
R1670 drain_left.n81 drain_left.n80 9.3005
R1671 drain_left.n79 drain_left.n78 9.3005
R1672 drain_left.n30 drain_left.n29 9.3005
R1673 drain_left.n73 drain_left.n72 9.3005
R1674 drain_left.n71 drain_left.n70 9.3005
R1675 drain_left.n47 drain_left.n46 9.3005
R1676 drain_left.n42 drain_left.n41 9.3005
R1677 drain_left.n53 drain_left.n52 9.3005
R1678 drain_left.n55 drain_left.n54 9.3005
R1679 drain_left.n38 drain_left.n37 9.3005
R1680 drain_left.n61 drain_left.n60 9.3005
R1681 drain_left.n63 drain_left.n62 9.3005
R1682 drain_left.n64 drain_left.n33 9.3005
R1683 drain_left.n22 drain_left.n21 9.3005
R1684 drain_left.n95 drain_left.n94 9.3005
R1685 drain_left.n97 drain_left.n96 9.3005
R1686 drain_left.n18 drain_left.n17 9.3005
R1687 drain_left.n103 drain_left.n102 9.3005
R1688 drain_left.n105 drain_left.n104 9.3005
R1689 drain_left.n14 drain_left.n13 9.3005
R1690 drain_left.n112 drain_left.n111 9.3005
R1691 drain_left.n114 drain_left.n113 9.3005
R1692 drain_left.n137 drain_left.n136 9.3005
R1693 drain_left.n194 drain_left.n193 9.3005
R1694 drain_left.n189 drain_left.n188 9.3005
R1695 drain_left.n200 drain_left.n199 9.3005
R1696 drain_left.n202 drain_left.n201 9.3005
R1697 drain_left.n185 drain_left.n184 9.3005
R1698 drain_left.n208 drain_left.n207 9.3005
R1699 drain_left.n210 drain_left.n209 9.3005
R1700 drain_left.n182 drain_left.n179 9.3005
R1701 drain_left.n241 drain_left.n240 9.3005
R1702 drain_left.n243 drain_left.n242 9.3005
R1703 drain_left.n164 drain_left.n163 9.3005
R1704 drain_left.n249 drain_left.n248 9.3005
R1705 drain_left.n251 drain_left.n250 9.3005
R1706 drain_left.n159 drain_left.n158 9.3005
R1707 drain_left.n257 drain_left.n256 9.3005
R1708 drain_left.n259 drain_left.n258 9.3005
R1709 drain_left.n282 drain_left.n281 9.3005
R1710 drain_left.n147 drain_left.n146 9.3005
R1711 drain_left.n276 drain_left.n275 9.3005
R1712 drain_left.n274 drain_left.n273 9.3005
R1713 drain_left.n151 drain_left.n150 9.3005
R1714 drain_left.n268 drain_left.n267 9.3005
R1715 drain_left.n266 drain_left.n265 9.3005
R1716 drain_left.n155 drain_left.n154 9.3005
R1717 drain_left.n168 drain_left.n167 9.3005
R1718 drain_left.n235 drain_left.n234 9.3005
R1719 drain_left.n233 drain_left.n232 9.3005
R1720 drain_left.n172 drain_left.n171 9.3005
R1721 drain_left.n227 drain_left.n226 9.3005
R1722 drain_left.n225 drain_left.n224 9.3005
R1723 drain_left.n176 drain_left.n175 9.3005
R1724 drain_left.n219 drain_left.n218 9.3005
R1725 drain_left.n217 drain_left.n216 9.3005
R1726 drain_left.n52 drain_left.n51 8.92171
R1727 drain_left.n85 drain_left.n26 8.92171
R1728 drain_left.n98 drain_left.n18 8.92171
R1729 drain_left.n132 drain_left.n131 8.92171
R1730 drain_left.n277 drain_left.n276 8.92171
R1731 drain_left.n244 drain_left.n164 8.92171
R1732 drain_left.n231 drain_left.n172 8.92171
R1733 drain_left.n199 drain_left.n198 8.92171
R1734 drain_left.n48 drain_left.n42 8.14595
R1735 drain_left.n86 drain_left.n24 8.14595
R1736 drain_left.n97 drain_left.n20 8.14595
R1737 drain_left.n135 drain_left.n2 8.14595
R1738 drain_left.n280 drain_left.n147 8.14595
R1739 drain_left.n243 drain_left.n166 8.14595
R1740 drain_left.n232 drain_left.n170 8.14595
R1741 drain_left.n195 drain_left.n189 8.14595
R1742 drain_left.n47 drain_left.n44 7.3702
R1743 drain_left.n90 drain_left.n89 7.3702
R1744 drain_left.n94 drain_left.n93 7.3702
R1745 drain_left.n136 drain_left.n0 7.3702
R1746 drain_left.n281 drain_left.n145 7.3702
R1747 drain_left.n240 drain_left.n239 7.3702
R1748 drain_left.n236 drain_left.n235 7.3702
R1749 drain_left.n194 drain_left.n191 7.3702
R1750 drain_left.n90 drain_left.n22 6.59444
R1751 drain_left.n93 drain_left.n22 6.59444
R1752 drain_left.n138 drain_left.n0 6.59444
R1753 drain_left.n283 drain_left.n145 6.59444
R1754 drain_left.n239 drain_left.n168 6.59444
R1755 drain_left.n236 drain_left.n168 6.59444
R1756 drain_left drain_left.n289 6.36873
R1757 drain_left.n48 drain_left.n47 5.81868
R1758 drain_left.n89 drain_left.n24 5.81868
R1759 drain_left.n94 drain_left.n20 5.81868
R1760 drain_left.n136 drain_left.n135 5.81868
R1761 drain_left.n281 drain_left.n280 5.81868
R1762 drain_left.n240 drain_left.n166 5.81868
R1763 drain_left.n235 drain_left.n170 5.81868
R1764 drain_left.n195 drain_left.n194 5.81868
R1765 drain_left.n51 drain_left.n42 5.04292
R1766 drain_left.n86 drain_left.n85 5.04292
R1767 drain_left.n98 drain_left.n97 5.04292
R1768 drain_left.n132 drain_left.n2 5.04292
R1769 drain_left.n277 drain_left.n147 5.04292
R1770 drain_left.n244 drain_left.n243 5.04292
R1771 drain_left.n232 drain_left.n231 5.04292
R1772 drain_left.n198 drain_left.n189 5.04292
R1773 drain_left.n52 drain_left.n40 4.26717
R1774 drain_left.n82 drain_left.n26 4.26717
R1775 drain_left.n101 drain_left.n18 4.26717
R1776 drain_left.n131 drain_left.n4 4.26717
R1777 drain_left.n276 drain_left.n149 4.26717
R1778 drain_left.n247 drain_left.n164 4.26717
R1779 drain_left.n228 drain_left.n172 4.26717
R1780 drain_left.n199 drain_left.n187 4.26717
R1781 drain_left.n56 drain_left.n55 3.49141
R1782 drain_left.n81 drain_left.n28 3.49141
R1783 drain_left.n102 drain_left.n16 3.49141
R1784 drain_left.n128 drain_left.n127 3.49141
R1785 drain_left.n273 drain_left.n272 3.49141
R1786 drain_left.n248 drain_left.n162 3.49141
R1787 drain_left.n227 drain_left.n174 3.49141
R1788 drain_left.n203 drain_left.n202 3.49141
R1789 drain_left.n193 drain_left.n192 2.84303
R1790 drain_left.n46 drain_left.n45 2.84303
R1791 drain_left.n59 drain_left.n38 2.71565
R1792 drain_left.n78 drain_left.n77 2.71565
R1793 drain_left.n106 drain_left.n105 2.71565
R1794 drain_left.n124 drain_left.n6 2.71565
R1795 drain_left.n269 drain_left.n151 2.71565
R1796 drain_left.n252 drain_left.n251 2.71565
R1797 drain_left.n224 drain_left.n223 2.71565
R1798 drain_left.n206 drain_left.n185 2.71565
R1799 drain_left.n60 drain_left.n36 1.93989
R1800 drain_left.n74 drain_left.n30 1.93989
R1801 drain_left.n110 drain_left.n14 1.93989
R1802 drain_left.n123 drain_left.n8 1.93989
R1803 drain_left.n268 drain_left.n153 1.93989
R1804 drain_left.n255 drain_left.n159 1.93989
R1805 drain_left.n220 drain_left.n176 1.93989
R1806 drain_left.n207 drain_left.n183 1.93989
R1807 drain_left.n65 drain_left.n63 1.16414
R1808 drain_left.n73 drain_left.n32 1.16414
R1809 drain_left.n111 drain_left.n12 1.16414
R1810 drain_left.n120 drain_left.n119 1.16414
R1811 drain_left.n265 drain_left.n264 1.16414
R1812 drain_left.n256 drain_left.n157 1.16414
R1813 drain_left.n219 drain_left.n178 1.16414
R1814 drain_left.n211 drain_left.n210 1.16414
R1815 drain_left.n141 drain_left.t0 0.7925
R1816 drain_left.n141 drain_left.t1 0.7925
R1817 drain_left.n142 drain_left.t13 0.7925
R1818 drain_left.n142 drain_left.t8 0.7925
R1819 drain_left.n139 drain_left.t6 0.7925
R1820 drain_left.n139 drain_left.t12 0.7925
R1821 drain_left.n288 drain_left.t2 0.7925
R1822 drain_left.n288 drain_left.t7 0.7925
R1823 drain_left.n286 drain_left.t9 0.7925
R1824 drain_left.n286 drain_left.t4 0.7925
R1825 drain_left.n284 drain_left.t5 0.7925
R1826 drain_left.n284 drain_left.t3 0.7925
R1827 drain_left.n287 drain_left.n285 0.716017
R1828 drain_left.n289 drain_left.n287 0.716017
R1829 drain_left.n144 drain_left.n140 0.481792
R1830 drain_left.n64 drain_left.n34 0.388379
R1831 drain_left.n70 drain_left.n69 0.388379
R1832 drain_left.n115 drain_left.n114 0.388379
R1833 drain_left.n116 drain_left.n10 0.388379
R1834 drain_left.n261 drain_left.n155 0.388379
R1835 drain_left.n260 drain_left.n259 0.388379
R1836 drain_left.n216 drain_left.n215 0.388379
R1837 drain_left.n182 drain_left.n180 0.388379
R1838 drain_left.n46 drain_left.n41 0.155672
R1839 drain_left.n53 drain_left.n41 0.155672
R1840 drain_left.n54 drain_left.n53 0.155672
R1841 drain_left.n54 drain_left.n37 0.155672
R1842 drain_left.n61 drain_left.n37 0.155672
R1843 drain_left.n62 drain_left.n61 0.155672
R1844 drain_left.n62 drain_left.n33 0.155672
R1845 drain_left.n71 drain_left.n33 0.155672
R1846 drain_left.n72 drain_left.n71 0.155672
R1847 drain_left.n72 drain_left.n29 0.155672
R1848 drain_left.n79 drain_left.n29 0.155672
R1849 drain_left.n80 drain_left.n79 0.155672
R1850 drain_left.n80 drain_left.n25 0.155672
R1851 drain_left.n87 drain_left.n25 0.155672
R1852 drain_left.n88 drain_left.n87 0.155672
R1853 drain_left.n88 drain_left.n21 0.155672
R1854 drain_left.n95 drain_left.n21 0.155672
R1855 drain_left.n96 drain_left.n95 0.155672
R1856 drain_left.n96 drain_left.n17 0.155672
R1857 drain_left.n103 drain_left.n17 0.155672
R1858 drain_left.n104 drain_left.n103 0.155672
R1859 drain_left.n104 drain_left.n13 0.155672
R1860 drain_left.n112 drain_left.n13 0.155672
R1861 drain_left.n113 drain_left.n112 0.155672
R1862 drain_left.n113 drain_left.n9 0.155672
R1863 drain_left.n121 drain_left.n9 0.155672
R1864 drain_left.n122 drain_left.n121 0.155672
R1865 drain_left.n122 drain_left.n5 0.155672
R1866 drain_left.n129 drain_left.n5 0.155672
R1867 drain_left.n130 drain_left.n129 0.155672
R1868 drain_left.n130 drain_left.n1 0.155672
R1869 drain_left.n137 drain_left.n1 0.155672
R1870 drain_left.n282 drain_left.n146 0.155672
R1871 drain_left.n275 drain_left.n146 0.155672
R1872 drain_left.n275 drain_left.n274 0.155672
R1873 drain_left.n274 drain_left.n150 0.155672
R1874 drain_left.n267 drain_left.n150 0.155672
R1875 drain_left.n267 drain_left.n266 0.155672
R1876 drain_left.n266 drain_left.n154 0.155672
R1877 drain_left.n258 drain_left.n154 0.155672
R1878 drain_left.n258 drain_left.n257 0.155672
R1879 drain_left.n257 drain_left.n158 0.155672
R1880 drain_left.n250 drain_left.n158 0.155672
R1881 drain_left.n250 drain_left.n249 0.155672
R1882 drain_left.n249 drain_left.n163 0.155672
R1883 drain_left.n242 drain_left.n163 0.155672
R1884 drain_left.n242 drain_left.n241 0.155672
R1885 drain_left.n241 drain_left.n167 0.155672
R1886 drain_left.n234 drain_left.n167 0.155672
R1887 drain_left.n234 drain_left.n233 0.155672
R1888 drain_left.n233 drain_left.n171 0.155672
R1889 drain_left.n226 drain_left.n171 0.155672
R1890 drain_left.n226 drain_left.n225 0.155672
R1891 drain_left.n225 drain_left.n175 0.155672
R1892 drain_left.n218 drain_left.n175 0.155672
R1893 drain_left.n218 drain_left.n217 0.155672
R1894 drain_left.n217 drain_left.n179 0.155672
R1895 drain_left.n209 drain_left.n179 0.155672
R1896 drain_left.n209 drain_left.n208 0.155672
R1897 drain_left.n208 drain_left.n184 0.155672
R1898 drain_left.n201 drain_left.n184 0.155672
R1899 drain_left.n201 drain_left.n200 0.155672
R1900 drain_left.n200 drain_left.n188 0.155672
R1901 drain_left.n193 drain_left.n188 0.155672
R1902 drain_left.n144 drain_left.n143 0.124033
C0 plus drain_right 0.359555f
C1 minus drain_left 0.172393f
C2 source drain_left 42.500603f
C3 minus drain_right 14.9189f
C4 minus plus 8.103241f
C5 source drain_right 42.482998f
C6 source plus 14.250599f
C7 minus source 14.2354f
C8 drain_left drain_right 1.06395f
C9 drain_left plus 15.113501f
C10 drain_right a_n2044_n5888# 11.02172f
C11 drain_left a_n2044_n5888# 11.333529f
C12 source a_n2044_n5888# 11.044921f
C13 minus a_n2044_n5888# 8.91586f
C14 plus a_n2044_n5888# 11.506802f
C15 drain_left.n0 a_n2044_n5888# 0.037053f
C16 drain_left.n1 a_n2044_n5888# 0.026877f
C17 drain_left.n2 a_n2044_n5888# 0.014443f
C18 drain_left.n3 a_n2044_n5888# 0.034137f
C19 drain_left.n4 a_n2044_n5888# 0.015292f
C20 drain_left.n5 a_n2044_n5888# 0.026877f
C21 drain_left.n6 a_n2044_n5888# 0.014443f
C22 drain_left.n7 a_n2044_n5888# 0.034137f
C23 drain_left.n8 a_n2044_n5888# 0.015292f
C24 drain_left.n9 a_n2044_n5888# 0.026877f
C25 drain_left.n10 a_n2044_n5888# 0.014443f
C26 drain_left.n11 a_n2044_n5888# 0.034137f
C27 drain_left.n12 a_n2044_n5888# 0.015292f
C28 drain_left.n13 a_n2044_n5888# 0.026877f
C29 drain_left.n14 a_n2044_n5888# 0.014443f
C30 drain_left.n15 a_n2044_n5888# 0.034137f
C31 drain_left.n16 a_n2044_n5888# 0.015292f
C32 drain_left.n17 a_n2044_n5888# 0.026877f
C33 drain_left.n18 a_n2044_n5888# 0.014443f
C34 drain_left.n19 a_n2044_n5888# 0.034137f
C35 drain_left.n20 a_n2044_n5888# 0.015292f
C36 drain_left.n21 a_n2044_n5888# 0.026877f
C37 drain_left.n22 a_n2044_n5888# 0.014443f
C38 drain_left.n23 a_n2044_n5888# 0.034137f
C39 drain_left.n24 a_n2044_n5888# 0.015292f
C40 drain_left.n25 a_n2044_n5888# 0.026877f
C41 drain_left.n26 a_n2044_n5888# 0.014443f
C42 drain_left.n27 a_n2044_n5888# 0.034137f
C43 drain_left.n28 a_n2044_n5888# 0.015292f
C44 drain_left.n29 a_n2044_n5888# 0.026877f
C45 drain_left.n30 a_n2044_n5888# 0.014443f
C46 drain_left.n31 a_n2044_n5888# 0.034137f
C47 drain_left.n32 a_n2044_n5888# 0.015292f
C48 drain_left.n33 a_n2044_n5888# 0.026877f
C49 drain_left.n34 a_n2044_n5888# 0.014867f
C50 drain_left.n35 a_n2044_n5888# 0.034137f
C51 drain_left.n36 a_n2044_n5888# 0.015292f
C52 drain_left.n37 a_n2044_n5888# 0.026877f
C53 drain_left.n38 a_n2044_n5888# 0.014443f
C54 drain_left.n39 a_n2044_n5888# 0.034137f
C55 drain_left.n40 a_n2044_n5888# 0.015292f
C56 drain_left.n41 a_n2044_n5888# 0.026877f
C57 drain_left.n42 a_n2044_n5888# 0.014443f
C58 drain_left.n43 a_n2044_n5888# 0.025603f
C59 drain_left.n44 a_n2044_n5888# 0.024132f
C60 drain_left.t10 a_n2044_n5888# 0.059537f
C61 drain_left.n45 a_n2044_n5888# 0.327925f
C62 drain_left.n46 a_n2044_n5888# 2.91001f
C63 drain_left.n47 a_n2044_n5888# 0.014443f
C64 drain_left.n48 a_n2044_n5888# 0.015292f
C65 drain_left.n49 a_n2044_n5888# 0.034137f
C66 drain_left.n50 a_n2044_n5888# 0.034137f
C67 drain_left.n51 a_n2044_n5888# 0.015292f
C68 drain_left.n52 a_n2044_n5888# 0.014443f
C69 drain_left.n53 a_n2044_n5888# 0.026877f
C70 drain_left.n54 a_n2044_n5888# 0.026877f
C71 drain_left.n55 a_n2044_n5888# 0.014443f
C72 drain_left.n56 a_n2044_n5888# 0.015292f
C73 drain_left.n57 a_n2044_n5888# 0.034137f
C74 drain_left.n58 a_n2044_n5888# 0.034137f
C75 drain_left.n59 a_n2044_n5888# 0.015292f
C76 drain_left.n60 a_n2044_n5888# 0.014443f
C77 drain_left.n61 a_n2044_n5888# 0.026877f
C78 drain_left.n62 a_n2044_n5888# 0.026877f
C79 drain_left.n63 a_n2044_n5888# 0.014443f
C80 drain_left.n64 a_n2044_n5888# 0.014443f
C81 drain_left.n65 a_n2044_n5888# 0.015292f
C82 drain_left.n66 a_n2044_n5888# 0.034137f
C83 drain_left.n67 a_n2044_n5888# 0.034137f
C84 drain_left.n68 a_n2044_n5888# 0.034137f
C85 drain_left.n69 a_n2044_n5888# 0.014867f
C86 drain_left.n70 a_n2044_n5888# 0.014443f
C87 drain_left.n71 a_n2044_n5888# 0.026877f
C88 drain_left.n72 a_n2044_n5888# 0.026877f
C89 drain_left.n73 a_n2044_n5888# 0.014443f
C90 drain_left.n74 a_n2044_n5888# 0.015292f
C91 drain_left.n75 a_n2044_n5888# 0.034137f
C92 drain_left.n76 a_n2044_n5888# 0.034137f
C93 drain_left.n77 a_n2044_n5888# 0.015292f
C94 drain_left.n78 a_n2044_n5888# 0.014443f
C95 drain_left.n79 a_n2044_n5888# 0.026877f
C96 drain_left.n80 a_n2044_n5888# 0.026877f
C97 drain_left.n81 a_n2044_n5888# 0.014443f
C98 drain_left.n82 a_n2044_n5888# 0.015292f
C99 drain_left.n83 a_n2044_n5888# 0.034137f
C100 drain_left.n84 a_n2044_n5888# 0.034137f
C101 drain_left.n85 a_n2044_n5888# 0.015292f
C102 drain_left.n86 a_n2044_n5888# 0.014443f
C103 drain_left.n87 a_n2044_n5888# 0.026877f
C104 drain_left.n88 a_n2044_n5888# 0.026877f
C105 drain_left.n89 a_n2044_n5888# 0.014443f
C106 drain_left.n90 a_n2044_n5888# 0.015292f
C107 drain_left.n91 a_n2044_n5888# 0.034137f
C108 drain_left.n92 a_n2044_n5888# 0.034137f
C109 drain_left.n93 a_n2044_n5888# 0.015292f
C110 drain_left.n94 a_n2044_n5888# 0.014443f
C111 drain_left.n95 a_n2044_n5888# 0.026877f
C112 drain_left.n96 a_n2044_n5888# 0.026877f
C113 drain_left.n97 a_n2044_n5888# 0.014443f
C114 drain_left.n98 a_n2044_n5888# 0.015292f
C115 drain_left.n99 a_n2044_n5888# 0.034137f
C116 drain_left.n100 a_n2044_n5888# 0.034137f
C117 drain_left.n101 a_n2044_n5888# 0.015292f
C118 drain_left.n102 a_n2044_n5888# 0.014443f
C119 drain_left.n103 a_n2044_n5888# 0.026877f
C120 drain_left.n104 a_n2044_n5888# 0.026877f
C121 drain_left.n105 a_n2044_n5888# 0.014443f
C122 drain_left.n106 a_n2044_n5888# 0.015292f
C123 drain_left.n107 a_n2044_n5888# 0.034137f
C124 drain_left.n108 a_n2044_n5888# 0.034137f
C125 drain_left.n109 a_n2044_n5888# 0.034137f
C126 drain_left.n110 a_n2044_n5888# 0.015292f
C127 drain_left.n111 a_n2044_n5888# 0.014443f
C128 drain_left.n112 a_n2044_n5888# 0.026877f
C129 drain_left.n113 a_n2044_n5888# 0.026877f
C130 drain_left.n114 a_n2044_n5888# 0.014443f
C131 drain_left.n115 a_n2044_n5888# 0.014867f
C132 drain_left.n116 a_n2044_n5888# 0.014867f
C133 drain_left.n117 a_n2044_n5888# 0.034137f
C134 drain_left.n118 a_n2044_n5888# 0.034137f
C135 drain_left.n119 a_n2044_n5888# 0.015292f
C136 drain_left.n120 a_n2044_n5888# 0.014443f
C137 drain_left.n121 a_n2044_n5888# 0.026877f
C138 drain_left.n122 a_n2044_n5888# 0.026877f
C139 drain_left.n123 a_n2044_n5888# 0.014443f
C140 drain_left.n124 a_n2044_n5888# 0.015292f
C141 drain_left.n125 a_n2044_n5888# 0.034137f
C142 drain_left.n126 a_n2044_n5888# 0.034137f
C143 drain_left.n127 a_n2044_n5888# 0.015292f
C144 drain_left.n128 a_n2044_n5888# 0.014443f
C145 drain_left.n129 a_n2044_n5888# 0.026877f
C146 drain_left.n130 a_n2044_n5888# 0.026877f
C147 drain_left.n131 a_n2044_n5888# 0.014443f
C148 drain_left.n132 a_n2044_n5888# 0.015292f
C149 drain_left.n133 a_n2044_n5888# 0.034137f
C150 drain_left.n134 a_n2044_n5888# 0.072619f
C151 drain_left.n135 a_n2044_n5888# 0.015292f
C152 drain_left.n136 a_n2044_n5888# 0.014443f
C153 drain_left.n137 a_n2044_n5888# 0.059188f
C154 drain_left.n138 a_n2044_n5888# 0.060661f
C155 drain_left.t6 a_n2044_n5888# 0.53098f
C156 drain_left.t12 a_n2044_n5888# 0.53098f
C157 drain_left.n139 a_n2044_n5888# 4.89356f
C158 drain_left.n140 a_n2044_n5888# 0.442506f
C159 drain_left.t0 a_n2044_n5888# 0.53098f
C160 drain_left.t1 a_n2044_n5888# 0.53098f
C161 drain_left.n141 a_n2044_n5888# 4.89791f
C162 drain_left.t13 a_n2044_n5888# 0.53098f
C163 drain_left.t8 a_n2044_n5888# 0.53098f
C164 drain_left.n142 a_n2044_n5888# 4.89356f
C165 drain_left.n143 a_n2044_n5888# 0.662493f
C166 drain_left.n144 a_n2044_n5888# 2.26302f
C167 drain_left.n145 a_n2044_n5888# 0.037053f
C168 drain_left.n146 a_n2044_n5888# 0.026877f
C169 drain_left.n147 a_n2044_n5888# 0.014443f
C170 drain_left.n148 a_n2044_n5888# 0.034137f
C171 drain_left.n149 a_n2044_n5888# 0.015292f
C172 drain_left.n150 a_n2044_n5888# 0.026877f
C173 drain_left.n151 a_n2044_n5888# 0.014443f
C174 drain_left.n152 a_n2044_n5888# 0.034137f
C175 drain_left.n153 a_n2044_n5888# 0.015292f
C176 drain_left.n154 a_n2044_n5888# 0.026877f
C177 drain_left.n155 a_n2044_n5888# 0.014443f
C178 drain_left.n156 a_n2044_n5888# 0.034137f
C179 drain_left.n157 a_n2044_n5888# 0.015292f
C180 drain_left.n158 a_n2044_n5888# 0.026877f
C181 drain_left.n159 a_n2044_n5888# 0.014443f
C182 drain_left.n160 a_n2044_n5888# 0.034137f
C183 drain_left.n161 a_n2044_n5888# 0.034137f
C184 drain_left.n162 a_n2044_n5888# 0.015292f
C185 drain_left.n163 a_n2044_n5888# 0.026877f
C186 drain_left.n164 a_n2044_n5888# 0.014443f
C187 drain_left.n165 a_n2044_n5888# 0.034137f
C188 drain_left.n166 a_n2044_n5888# 0.015292f
C189 drain_left.n167 a_n2044_n5888# 0.026877f
C190 drain_left.n168 a_n2044_n5888# 0.014443f
C191 drain_left.n169 a_n2044_n5888# 0.034137f
C192 drain_left.n170 a_n2044_n5888# 0.015292f
C193 drain_left.n171 a_n2044_n5888# 0.026877f
C194 drain_left.n172 a_n2044_n5888# 0.014443f
C195 drain_left.n173 a_n2044_n5888# 0.034137f
C196 drain_left.n174 a_n2044_n5888# 0.015292f
C197 drain_left.n175 a_n2044_n5888# 0.026877f
C198 drain_left.n176 a_n2044_n5888# 0.014443f
C199 drain_left.n177 a_n2044_n5888# 0.034137f
C200 drain_left.n178 a_n2044_n5888# 0.015292f
C201 drain_left.n179 a_n2044_n5888# 0.026877f
C202 drain_left.n180 a_n2044_n5888# 0.014867f
C203 drain_left.n181 a_n2044_n5888# 0.034137f
C204 drain_left.n182 a_n2044_n5888# 0.014443f
C205 drain_left.n183 a_n2044_n5888# 0.015292f
C206 drain_left.n184 a_n2044_n5888# 0.026877f
C207 drain_left.n185 a_n2044_n5888# 0.014443f
C208 drain_left.n186 a_n2044_n5888# 0.034137f
C209 drain_left.n187 a_n2044_n5888# 0.015292f
C210 drain_left.n188 a_n2044_n5888# 0.026877f
C211 drain_left.n189 a_n2044_n5888# 0.014443f
C212 drain_left.n190 a_n2044_n5888# 0.025603f
C213 drain_left.n191 a_n2044_n5888# 0.024132f
C214 drain_left.t11 a_n2044_n5888# 0.059537f
C215 drain_left.n192 a_n2044_n5888# 0.327925f
C216 drain_left.n193 a_n2044_n5888# 2.91001f
C217 drain_left.n194 a_n2044_n5888# 0.014443f
C218 drain_left.n195 a_n2044_n5888# 0.015292f
C219 drain_left.n196 a_n2044_n5888# 0.034137f
C220 drain_left.n197 a_n2044_n5888# 0.034137f
C221 drain_left.n198 a_n2044_n5888# 0.015292f
C222 drain_left.n199 a_n2044_n5888# 0.014443f
C223 drain_left.n200 a_n2044_n5888# 0.026877f
C224 drain_left.n201 a_n2044_n5888# 0.026877f
C225 drain_left.n202 a_n2044_n5888# 0.014443f
C226 drain_left.n203 a_n2044_n5888# 0.015292f
C227 drain_left.n204 a_n2044_n5888# 0.034137f
C228 drain_left.n205 a_n2044_n5888# 0.034137f
C229 drain_left.n206 a_n2044_n5888# 0.015292f
C230 drain_left.n207 a_n2044_n5888# 0.014443f
C231 drain_left.n208 a_n2044_n5888# 0.026877f
C232 drain_left.n209 a_n2044_n5888# 0.026877f
C233 drain_left.n210 a_n2044_n5888# 0.014443f
C234 drain_left.n211 a_n2044_n5888# 0.015292f
C235 drain_left.n212 a_n2044_n5888# 0.034137f
C236 drain_left.n213 a_n2044_n5888# 0.034137f
C237 drain_left.n214 a_n2044_n5888# 0.034137f
C238 drain_left.n215 a_n2044_n5888# 0.014867f
C239 drain_left.n216 a_n2044_n5888# 0.014443f
C240 drain_left.n217 a_n2044_n5888# 0.026877f
C241 drain_left.n218 a_n2044_n5888# 0.026877f
C242 drain_left.n219 a_n2044_n5888# 0.014443f
C243 drain_left.n220 a_n2044_n5888# 0.015292f
C244 drain_left.n221 a_n2044_n5888# 0.034137f
C245 drain_left.n222 a_n2044_n5888# 0.034137f
C246 drain_left.n223 a_n2044_n5888# 0.015292f
C247 drain_left.n224 a_n2044_n5888# 0.014443f
C248 drain_left.n225 a_n2044_n5888# 0.026877f
C249 drain_left.n226 a_n2044_n5888# 0.026877f
C250 drain_left.n227 a_n2044_n5888# 0.014443f
C251 drain_left.n228 a_n2044_n5888# 0.015292f
C252 drain_left.n229 a_n2044_n5888# 0.034137f
C253 drain_left.n230 a_n2044_n5888# 0.034137f
C254 drain_left.n231 a_n2044_n5888# 0.015292f
C255 drain_left.n232 a_n2044_n5888# 0.014443f
C256 drain_left.n233 a_n2044_n5888# 0.026877f
C257 drain_left.n234 a_n2044_n5888# 0.026877f
C258 drain_left.n235 a_n2044_n5888# 0.014443f
C259 drain_left.n236 a_n2044_n5888# 0.015292f
C260 drain_left.n237 a_n2044_n5888# 0.034137f
C261 drain_left.n238 a_n2044_n5888# 0.034137f
C262 drain_left.n239 a_n2044_n5888# 0.015292f
C263 drain_left.n240 a_n2044_n5888# 0.014443f
C264 drain_left.n241 a_n2044_n5888# 0.026877f
C265 drain_left.n242 a_n2044_n5888# 0.026877f
C266 drain_left.n243 a_n2044_n5888# 0.014443f
C267 drain_left.n244 a_n2044_n5888# 0.015292f
C268 drain_left.n245 a_n2044_n5888# 0.034137f
C269 drain_left.n246 a_n2044_n5888# 0.034137f
C270 drain_left.n247 a_n2044_n5888# 0.015292f
C271 drain_left.n248 a_n2044_n5888# 0.014443f
C272 drain_left.n249 a_n2044_n5888# 0.026877f
C273 drain_left.n250 a_n2044_n5888# 0.026877f
C274 drain_left.n251 a_n2044_n5888# 0.014443f
C275 drain_left.n252 a_n2044_n5888# 0.015292f
C276 drain_left.n253 a_n2044_n5888# 0.034137f
C277 drain_left.n254 a_n2044_n5888# 0.034137f
C278 drain_left.n255 a_n2044_n5888# 0.015292f
C279 drain_left.n256 a_n2044_n5888# 0.014443f
C280 drain_left.n257 a_n2044_n5888# 0.026877f
C281 drain_left.n258 a_n2044_n5888# 0.026877f
C282 drain_left.n259 a_n2044_n5888# 0.014443f
C283 drain_left.n260 a_n2044_n5888# 0.014867f
C284 drain_left.n261 a_n2044_n5888# 0.014867f
C285 drain_left.n262 a_n2044_n5888# 0.034137f
C286 drain_left.n263 a_n2044_n5888# 0.034137f
C287 drain_left.n264 a_n2044_n5888# 0.015292f
C288 drain_left.n265 a_n2044_n5888# 0.014443f
C289 drain_left.n266 a_n2044_n5888# 0.026877f
C290 drain_left.n267 a_n2044_n5888# 0.026877f
C291 drain_left.n268 a_n2044_n5888# 0.014443f
C292 drain_left.n269 a_n2044_n5888# 0.015292f
C293 drain_left.n270 a_n2044_n5888# 0.034137f
C294 drain_left.n271 a_n2044_n5888# 0.034137f
C295 drain_left.n272 a_n2044_n5888# 0.015292f
C296 drain_left.n273 a_n2044_n5888# 0.014443f
C297 drain_left.n274 a_n2044_n5888# 0.026877f
C298 drain_left.n275 a_n2044_n5888# 0.026877f
C299 drain_left.n276 a_n2044_n5888# 0.014443f
C300 drain_left.n277 a_n2044_n5888# 0.015292f
C301 drain_left.n278 a_n2044_n5888# 0.034137f
C302 drain_left.n279 a_n2044_n5888# 0.072619f
C303 drain_left.n280 a_n2044_n5888# 0.015292f
C304 drain_left.n281 a_n2044_n5888# 0.014443f
C305 drain_left.n282 a_n2044_n5888# 0.059188f
C306 drain_left.n283 a_n2044_n5888# 0.060661f
C307 drain_left.t5 a_n2044_n5888# 0.53098f
C308 drain_left.t3 a_n2044_n5888# 0.53098f
C309 drain_left.n284 a_n2044_n5888# 4.89356f
C310 drain_left.n285 a_n2044_n5888# 0.461495f
C311 drain_left.t9 a_n2044_n5888# 0.53098f
C312 drain_left.t4 a_n2044_n5888# 0.53098f
C313 drain_left.n286 a_n2044_n5888# 4.89356f
C314 drain_left.n287 a_n2044_n5888# 0.351123f
C315 drain_left.t2 a_n2044_n5888# 0.53098f
C316 drain_left.t7 a_n2044_n5888# 0.53098f
C317 drain_left.n288 a_n2044_n5888# 4.89354f
C318 drain_left.n289 a_n2044_n5888# 0.582049f
C319 plus.n0 a_n2044_n5888# 0.045999f
C320 plus.t6 a_n2044_n5888# 1.62491f
C321 plus.t11 a_n2044_n5888# 1.62491f
C322 plus.t9 a_n2044_n5888# 1.62491f
C323 plus.n1 a_n2044_n5888# 0.601586f
C324 plus.n2 a_n2044_n5888# 0.06138f
C325 plus.t4 a_n2044_n5888# 1.62491f
C326 plus.t10 a_n2044_n5888# 1.62491f
C327 plus.t8 a_n2044_n5888# 1.62491f
C328 plus.n3 a_n2044_n5888# 0.601302f
C329 plus.t2 a_n2044_n5888# 1.63451f
C330 plus.n4 a_n2044_n5888# 0.587519f
C331 plus.n5 a_n2044_n5888# 0.151256f
C332 plus.n6 a_n2044_n5888# 0.010438f
C333 plus.n7 a_n2044_n5888# 0.601586f
C334 plus.n8 a_n2044_n5888# 0.607203f
C335 plus.n9 a_n2044_n5888# 0.061236f
C336 plus.n10 a_n2044_n5888# 0.06138f
C337 plus.n11 a_n2044_n5888# 0.045999f
C338 plus.n12 a_n2044_n5888# 0.010438f
C339 plus.n13 a_n2044_n5888# 0.601302f
C340 plus.n14 a_n2044_n5888# 0.596765f
C341 plus.n15 a_n2044_n5888# 0.830749f
C342 plus.n16 a_n2044_n5888# 0.045999f
C343 plus.t3 a_n2044_n5888# 1.62491f
C344 plus.t7 a_n2044_n5888# 1.62491f
C345 plus.t1 a_n2044_n5888# 1.62491f
C346 plus.n17 a_n2044_n5888# 0.601586f
C347 plus.n18 a_n2044_n5888# 0.06138f
C348 plus.t0 a_n2044_n5888# 1.62491f
C349 plus.t5 a_n2044_n5888# 1.62491f
C350 plus.t13 a_n2044_n5888# 1.62491f
C351 plus.n19 a_n2044_n5888# 0.601302f
C352 plus.t12 a_n2044_n5888# 1.63451f
C353 plus.n20 a_n2044_n5888# 0.587519f
C354 plus.n21 a_n2044_n5888# 0.151256f
C355 plus.n22 a_n2044_n5888# 0.010438f
C356 plus.n23 a_n2044_n5888# 0.601586f
C357 plus.n24 a_n2044_n5888# 0.607203f
C358 plus.n25 a_n2044_n5888# 0.061236f
C359 plus.n26 a_n2044_n5888# 0.06138f
C360 plus.n27 a_n2044_n5888# 0.045999f
C361 plus.n28 a_n2044_n5888# 0.010438f
C362 plus.n29 a_n2044_n5888# 0.601302f
C363 plus.n30 a_n2044_n5888# 0.596765f
C364 plus.n31 a_n2044_n5888# 1.83272f
C365 drain_right.n0 a_n2044_n5888# 0.036992f
C366 drain_right.n1 a_n2044_n5888# 0.026833f
C367 drain_right.n2 a_n2044_n5888# 0.014419f
C368 drain_right.n3 a_n2044_n5888# 0.034081f
C369 drain_right.n4 a_n2044_n5888# 0.015267f
C370 drain_right.n5 a_n2044_n5888# 0.026833f
C371 drain_right.n6 a_n2044_n5888# 0.014419f
C372 drain_right.n7 a_n2044_n5888# 0.034081f
C373 drain_right.n8 a_n2044_n5888# 0.015267f
C374 drain_right.n9 a_n2044_n5888# 0.026833f
C375 drain_right.n10 a_n2044_n5888# 0.014419f
C376 drain_right.n11 a_n2044_n5888# 0.034081f
C377 drain_right.n12 a_n2044_n5888# 0.015267f
C378 drain_right.n13 a_n2044_n5888# 0.026833f
C379 drain_right.n14 a_n2044_n5888# 0.014419f
C380 drain_right.n15 a_n2044_n5888# 0.034081f
C381 drain_right.n16 a_n2044_n5888# 0.015267f
C382 drain_right.n17 a_n2044_n5888# 0.026833f
C383 drain_right.n18 a_n2044_n5888# 0.014419f
C384 drain_right.n19 a_n2044_n5888# 0.034081f
C385 drain_right.n20 a_n2044_n5888# 0.015267f
C386 drain_right.n21 a_n2044_n5888# 0.026833f
C387 drain_right.n22 a_n2044_n5888# 0.014419f
C388 drain_right.n23 a_n2044_n5888# 0.034081f
C389 drain_right.n24 a_n2044_n5888# 0.015267f
C390 drain_right.n25 a_n2044_n5888# 0.026833f
C391 drain_right.n26 a_n2044_n5888# 0.014419f
C392 drain_right.n27 a_n2044_n5888# 0.034081f
C393 drain_right.n28 a_n2044_n5888# 0.015267f
C394 drain_right.n29 a_n2044_n5888# 0.026833f
C395 drain_right.n30 a_n2044_n5888# 0.014419f
C396 drain_right.n31 a_n2044_n5888# 0.034081f
C397 drain_right.n32 a_n2044_n5888# 0.015267f
C398 drain_right.n33 a_n2044_n5888# 0.026833f
C399 drain_right.n34 a_n2044_n5888# 0.014843f
C400 drain_right.n35 a_n2044_n5888# 0.034081f
C401 drain_right.n36 a_n2044_n5888# 0.015267f
C402 drain_right.n37 a_n2044_n5888# 0.026833f
C403 drain_right.n38 a_n2044_n5888# 0.014419f
C404 drain_right.n39 a_n2044_n5888# 0.034081f
C405 drain_right.n40 a_n2044_n5888# 0.015267f
C406 drain_right.n41 a_n2044_n5888# 0.026833f
C407 drain_right.n42 a_n2044_n5888# 0.014419f
C408 drain_right.n43 a_n2044_n5888# 0.025561f
C409 drain_right.n44 a_n2044_n5888# 0.024093f
C410 drain_right.t10 a_n2044_n5888# 0.059439f
C411 drain_right.n45 a_n2044_n5888# 0.327384f
C412 drain_right.n46 a_n2044_n5888# 2.90521f
C413 drain_right.n47 a_n2044_n5888# 0.014419f
C414 drain_right.n48 a_n2044_n5888# 0.015267f
C415 drain_right.n49 a_n2044_n5888# 0.034081f
C416 drain_right.n50 a_n2044_n5888# 0.034081f
C417 drain_right.n51 a_n2044_n5888# 0.015267f
C418 drain_right.n52 a_n2044_n5888# 0.014419f
C419 drain_right.n53 a_n2044_n5888# 0.026833f
C420 drain_right.n54 a_n2044_n5888# 0.026833f
C421 drain_right.n55 a_n2044_n5888# 0.014419f
C422 drain_right.n56 a_n2044_n5888# 0.015267f
C423 drain_right.n57 a_n2044_n5888# 0.034081f
C424 drain_right.n58 a_n2044_n5888# 0.034081f
C425 drain_right.n59 a_n2044_n5888# 0.015267f
C426 drain_right.n60 a_n2044_n5888# 0.014419f
C427 drain_right.n61 a_n2044_n5888# 0.026833f
C428 drain_right.n62 a_n2044_n5888# 0.026833f
C429 drain_right.n63 a_n2044_n5888# 0.014419f
C430 drain_right.n64 a_n2044_n5888# 0.014419f
C431 drain_right.n65 a_n2044_n5888# 0.015267f
C432 drain_right.n66 a_n2044_n5888# 0.034081f
C433 drain_right.n67 a_n2044_n5888# 0.034081f
C434 drain_right.n68 a_n2044_n5888# 0.034081f
C435 drain_right.n69 a_n2044_n5888# 0.014843f
C436 drain_right.n70 a_n2044_n5888# 0.014419f
C437 drain_right.n71 a_n2044_n5888# 0.026833f
C438 drain_right.n72 a_n2044_n5888# 0.026833f
C439 drain_right.n73 a_n2044_n5888# 0.014419f
C440 drain_right.n74 a_n2044_n5888# 0.015267f
C441 drain_right.n75 a_n2044_n5888# 0.034081f
C442 drain_right.n76 a_n2044_n5888# 0.034081f
C443 drain_right.n77 a_n2044_n5888# 0.015267f
C444 drain_right.n78 a_n2044_n5888# 0.014419f
C445 drain_right.n79 a_n2044_n5888# 0.026833f
C446 drain_right.n80 a_n2044_n5888# 0.026833f
C447 drain_right.n81 a_n2044_n5888# 0.014419f
C448 drain_right.n82 a_n2044_n5888# 0.015267f
C449 drain_right.n83 a_n2044_n5888# 0.034081f
C450 drain_right.n84 a_n2044_n5888# 0.034081f
C451 drain_right.n85 a_n2044_n5888# 0.015267f
C452 drain_right.n86 a_n2044_n5888# 0.014419f
C453 drain_right.n87 a_n2044_n5888# 0.026833f
C454 drain_right.n88 a_n2044_n5888# 0.026833f
C455 drain_right.n89 a_n2044_n5888# 0.014419f
C456 drain_right.n90 a_n2044_n5888# 0.015267f
C457 drain_right.n91 a_n2044_n5888# 0.034081f
C458 drain_right.n92 a_n2044_n5888# 0.034081f
C459 drain_right.n93 a_n2044_n5888# 0.015267f
C460 drain_right.n94 a_n2044_n5888# 0.014419f
C461 drain_right.n95 a_n2044_n5888# 0.026833f
C462 drain_right.n96 a_n2044_n5888# 0.026833f
C463 drain_right.n97 a_n2044_n5888# 0.014419f
C464 drain_right.n98 a_n2044_n5888# 0.015267f
C465 drain_right.n99 a_n2044_n5888# 0.034081f
C466 drain_right.n100 a_n2044_n5888# 0.034081f
C467 drain_right.n101 a_n2044_n5888# 0.015267f
C468 drain_right.n102 a_n2044_n5888# 0.014419f
C469 drain_right.n103 a_n2044_n5888# 0.026833f
C470 drain_right.n104 a_n2044_n5888# 0.026833f
C471 drain_right.n105 a_n2044_n5888# 0.014419f
C472 drain_right.n106 a_n2044_n5888# 0.015267f
C473 drain_right.n107 a_n2044_n5888# 0.034081f
C474 drain_right.n108 a_n2044_n5888# 0.034081f
C475 drain_right.n109 a_n2044_n5888# 0.034081f
C476 drain_right.n110 a_n2044_n5888# 0.015267f
C477 drain_right.n111 a_n2044_n5888# 0.014419f
C478 drain_right.n112 a_n2044_n5888# 0.026833f
C479 drain_right.n113 a_n2044_n5888# 0.026833f
C480 drain_right.n114 a_n2044_n5888# 0.014419f
C481 drain_right.n115 a_n2044_n5888# 0.014843f
C482 drain_right.n116 a_n2044_n5888# 0.014843f
C483 drain_right.n117 a_n2044_n5888# 0.034081f
C484 drain_right.n118 a_n2044_n5888# 0.034081f
C485 drain_right.n119 a_n2044_n5888# 0.015267f
C486 drain_right.n120 a_n2044_n5888# 0.014419f
C487 drain_right.n121 a_n2044_n5888# 0.026833f
C488 drain_right.n122 a_n2044_n5888# 0.026833f
C489 drain_right.n123 a_n2044_n5888# 0.014419f
C490 drain_right.n124 a_n2044_n5888# 0.015267f
C491 drain_right.n125 a_n2044_n5888# 0.034081f
C492 drain_right.n126 a_n2044_n5888# 0.034081f
C493 drain_right.n127 a_n2044_n5888# 0.015267f
C494 drain_right.n128 a_n2044_n5888# 0.014419f
C495 drain_right.n129 a_n2044_n5888# 0.026833f
C496 drain_right.n130 a_n2044_n5888# 0.026833f
C497 drain_right.n131 a_n2044_n5888# 0.014419f
C498 drain_right.n132 a_n2044_n5888# 0.015267f
C499 drain_right.n133 a_n2044_n5888# 0.034081f
C500 drain_right.n134 a_n2044_n5888# 0.072499f
C501 drain_right.n135 a_n2044_n5888# 0.015267f
C502 drain_right.n136 a_n2044_n5888# 0.014419f
C503 drain_right.n137 a_n2044_n5888# 0.059091f
C504 drain_right.n138 a_n2044_n5888# 0.060561f
C505 drain_right.t11 a_n2044_n5888# 0.530104f
C506 drain_right.t4 a_n2044_n5888# 0.530104f
C507 drain_right.n139 a_n2044_n5888# 4.88548f
C508 drain_right.n140 a_n2044_n5888# 0.441776f
C509 drain_right.t1 a_n2044_n5888# 0.530104f
C510 drain_right.t2 a_n2044_n5888# 0.530104f
C511 drain_right.n141 a_n2044_n5888# 4.88983f
C512 drain_right.t5 a_n2044_n5888# 0.530104f
C513 drain_right.t7 a_n2044_n5888# 0.530104f
C514 drain_right.n142 a_n2044_n5888# 4.88548f
C515 drain_right.n143 a_n2044_n5888# 0.6614f
C516 drain_right.n144 a_n2044_n5888# 2.20379f
C517 drain_right.t12 a_n2044_n5888# 0.530104f
C518 drain_right.t3 a_n2044_n5888# 0.530104f
C519 drain_right.n145 a_n2044_n5888# 4.88982f
C520 drain_right.t0 a_n2044_n5888# 0.530104f
C521 drain_right.t8 a_n2044_n5888# 0.530104f
C522 drain_right.n146 a_n2044_n5888# 4.88548f
C523 drain_right.n147 a_n2044_n5888# 0.707558f
C524 drain_right.t6 a_n2044_n5888# 0.530104f
C525 drain_right.t9 a_n2044_n5888# 0.530104f
C526 drain_right.n148 a_n2044_n5888# 4.88548f
C527 drain_right.n149 a_n2044_n5888# 0.350544f
C528 drain_right.n150 a_n2044_n5888# 0.036992f
C529 drain_right.n151 a_n2044_n5888# 0.026833f
C530 drain_right.n152 a_n2044_n5888# 0.014419f
C531 drain_right.n153 a_n2044_n5888# 0.034081f
C532 drain_right.n154 a_n2044_n5888# 0.015267f
C533 drain_right.n155 a_n2044_n5888# 0.026833f
C534 drain_right.n156 a_n2044_n5888# 0.014419f
C535 drain_right.n157 a_n2044_n5888# 0.034081f
C536 drain_right.n158 a_n2044_n5888# 0.015267f
C537 drain_right.n159 a_n2044_n5888# 0.026833f
C538 drain_right.n160 a_n2044_n5888# 0.014419f
C539 drain_right.n161 a_n2044_n5888# 0.034081f
C540 drain_right.n162 a_n2044_n5888# 0.015267f
C541 drain_right.n163 a_n2044_n5888# 0.026833f
C542 drain_right.n164 a_n2044_n5888# 0.014419f
C543 drain_right.n165 a_n2044_n5888# 0.034081f
C544 drain_right.n166 a_n2044_n5888# 0.034081f
C545 drain_right.n167 a_n2044_n5888# 0.015267f
C546 drain_right.n168 a_n2044_n5888# 0.026833f
C547 drain_right.n169 a_n2044_n5888# 0.014419f
C548 drain_right.n170 a_n2044_n5888# 0.034081f
C549 drain_right.n171 a_n2044_n5888# 0.015267f
C550 drain_right.n172 a_n2044_n5888# 0.026833f
C551 drain_right.n173 a_n2044_n5888# 0.014419f
C552 drain_right.n174 a_n2044_n5888# 0.034081f
C553 drain_right.n175 a_n2044_n5888# 0.015267f
C554 drain_right.n176 a_n2044_n5888# 0.026833f
C555 drain_right.n177 a_n2044_n5888# 0.014419f
C556 drain_right.n178 a_n2044_n5888# 0.034081f
C557 drain_right.n179 a_n2044_n5888# 0.015267f
C558 drain_right.n180 a_n2044_n5888# 0.026833f
C559 drain_right.n181 a_n2044_n5888# 0.014419f
C560 drain_right.n182 a_n2044_n5888# 0.034081f
C561 drain_right.n183 a_n2044_n5888# 0.015267f
C562 drain_right.n184 a_n2044_n5888# 0.026833f
C563 drain_right.n185 a_n2044_n5888# 0.014843f
C564 drain_right.n186 a_n2044_n5888# 0.034081f
C565 drain_right.n187 a_n2044_n5888# 0.014419f
C566 drain_right.n188 a_n2044_n5888# 0.015267f
C567 drain_right.n189 a_n2044_n5888# 0.026833f
C568 drain_right.n190 a_n2044_n5888# 0.014419f
C569 drain_right.n191 a_n2044_n5888# 0.034081f
C570 drain_right.n192 a_n2044_n5888# 0.015267f
C571 drain_right.n193 a_n2044_n5888# 0.026833f
C572 drain_right.n194 a_n2044_n5888# 0.014419f
C573 drain_right.n195 a_n2044_n5888# 0.025561f
C574 drain_right.n196 a_n2044_n5888# 0.024093f
C575 drain_right.t13 a_n2044_n5888# 0.059439f
C576 drain_right.n197 a_n2044_n5888# 0.327384f
C577 drain_right.n198 a_n2044_n5888# 2.90521f
C578 drain_right.n199 a_n2044_n5888# 0.014419f
C579 drain_right.n200 a_n2044_n5888# 0.015267f
C580 drain_right.n201 a_n2044_n5888# 0.034081f
C581 drain_right.n202 a_n2044_n5888# 0.034081f
C582 drain_right.n203 a_n2044_n5888# 0.015267f
C583 drain_right.n204 a_n2044_n5888# 0.014419f
C584 drain_right.n205 a_n2044_n5888# 0.026833f
C585 drain_right.n206 a_n2044_n5888# 0.026833f
C586 drain_right.n207 a_n2044_n5888# 0.014419f
C587 drain_right.n208 a_n2044_n5888# 0.015267f
C588 drain_right.n209 a_n2044_n5888# 0.034081f
C589 drain_right.n210 a_n2044_n5888# 0.034081f
C590 drain_right.n211 a_n2044_n5888# 0.015267f
C591 drain_right.n212 a_n2044_n5888# 0.014419f
C592 drain_right.n213 a_n2044_n5888# 0.026833f
C593 drain_right.n214 a_n2044_n5888# 0.026833f
C594 drain_right.n215 a_n2044_n5888# 0.014419f
C595 drain_right.n216 a_n2044_n5888# 0.015267f
C596 drain_right.n217 a_n2044_n5888# 0.034081f
C597 drain_right.n218 a_n2044_n5888# 0.034081f
C598 drain_right.n219 a_n2044_n5888# 0.034081f
C599 drain_right.n220 a_n2044_n5888# 0.014843f
C600 drain_right.n221 a_n2044_n5888# 0.014419f
C601 drain_right.n222 a_n2044_n5888# 0.026833f
C602 drain_right.n223 a_n2044_n5888# 0.026833f
C603 drain_right.n224 a_n2044_n5888# 0.014419f
C604 drain_right.n225 a_n2044_n5888# 0.015267f
C605 drain_right.n226 a_n2044_n5888# 0.034081f
C606 drain_right.n227 a_n2044_n5888# 0.034081f
C607 drain_right.n228 a_n2044_n5888# 0.015267f
C608 drain_right.n229 a_n2044_n5888# 0.014419f
C609 drain_right.n230 a_n2044_n5888# 0.026833f
C610 drain_right.n231 a_n2044_n5888# 0.026833f
C611 drain_right.n232 a_n2044_n5888# 0.014419f
C612 drain_right.n233 a_n2044_n5888# 0.015267f
C613 drain_right.n234 a_n2044_n5888# 0.034081f
C614 drain_right.n235 a_n2044_n5888# 0.034081f
C615 drain_right.n236 a_n2044_n5888# 0.015267f
C616 drain_right.n237 a_n2044_n5888# 0.014419f
C617 drain_right.n238 a_n2044_n5888# 0.026833f
C618 drain_right.n239 a_n2044_n5888# 0.026833f
C619 drain_right.n240 a_n2044_n5888# 0.014419f
C620 drain_right.n241 a_n2044_n5888# 0.015267f
C621 drain_right.n242 a_n2044_n5888# 0.034081f
C622 drain_right.n243 a_n2044_n5888# 0.034081f
C623 drain_right.n244 a_n2044_n5888# 0.015267f
C624 drain_right.n245 a_n2044_n5888# 0.014419f
C625 drain_right.n246 a_n2044_n5888# 0.026833f
C626 drain_right.n247 a_n2044_n5888# 0.026833f
C627 drain_right.n248 a_n2044_n5888# 0.014419f
C628 drain_right.n249 a_n2044_n5888# 0.015267f
C629 drain_right.n250 a_n2044_n5888# 0.034081f
C630 drain_right.n251 a_n2044_n5888# 0.034081f
C631 drain_right.n252 a_n2044_n5888# 0.015267f
C632 drain_right.n253 a_n2044_n5888# 0.014419f
C633 drain_right.n254 a_n2044_n5888# 0.026833f
C634 drain_right.n255 a_n2044_n5888# 0.026833f
C635 drain_right.n256 a_n2044_n5888# 0.014419f
C636 drain_right.n257 a_n2044_n5888# 0.015267f
C637 drain_right.n258 a_n2044_n5888# 0.034081f
C638 drain_right.n259 a_n2044_n5888# 0.034081f
C639 drain_right.n260 a_n2044_n5888# 0.015267f
C640 drain_right.n261 a_n2044_n5888# 0.014419f
C641 drain_right.n262 a_n2044_n5888# 0.026833f
C642 drain_right.n263 a_n2044_n5888# 0.026833f
C643 drain_right.n264 a_n2044_n5888# 0.014419f
C644 drain_right.n265 a_n2044_n5888# 0.014843f
C645 drain_right.n266 a_n2044_n5888# 0.014843f
C646 drain_right.n267 a_n2044_n5888# 0.034081f
C647 drain_right.n268 a_n2044_n5888# 0.034081f
C648 drain_right.n269 a_n2044_n5888# 0.015267f
C649 drain_right.n270 a_n2044_n5888# 0.014419f
C650 drain_right.n271 a_n2044_n5888# 0.026833f
C651 drain_right.n272 a_n2044_n5888# 0.026833f
C652 drain_right.n273 a_n2044_n5888# 0.014419f
C653 drain_right.n274 a_n2044_n5888# 0.015267f
C654 drain_right.n275 a_n2044_n5888# 0.034081f
C655 drain_right.n276 a_n2044_n5888# 0.034081f
C656 drain_right.n277 a_n2044_n5888# 0.015267f
C657 drain_right.n278 a_n2044_n5888# 0.014419f
C658 drain_right.n279 a_n2044_n5888# 0.026833f
C659 drain_right.n280 a_n2044_n5888# 0.026833f
C660 drain_right.n281 a_n2044_n5888# 0.014419f
C661 drain_right.n282 a_n2044_n5888# 0.015267f
C662 drain_right.n283 a_n2044_n5888# 0.034081f
C663 drain_right.n284 a_n2044_n5888# 0.072499f
C664 drain_right.n285 a_n2044_n5888# 0.015267f
C665 drain_right.n286 a_n2044_n5888# 0.014419f
C666 drain_right.n287 a_n2044_n5888# 0.059091f
C667 drain_right.n288 a_n2044_n5888# 0.058894f
C668 drain_right.n289 a_n2044_n5888# 0.347143f
C669 source.n0 a_n2044_n5888# 0.037526f
C670 source.n1 a_n2044_n5888# 0.02722f
C671 source.n2 a_n2044_n5888# 0.014627f
C672 source.n3 a_n2044_n5888# 0.034573f
C673 source.n4 a_n2044_n5888# 0.015487f
C674 source.n5 a_n2044_n5888# 0.02722f
C675 source.n6 a_n2044_n5888# 0.014627f
C676 source.n7 a_n2044_n5888# 0.034573f
C677 source.n8 a_n2044_n5888# 0.015487f
C678 source.n9 a_n2044_n5888# 0.02722f
C679 source.n10 a_n2044_n5888# 0.014627f
C680 source.n11 a_n2044_n5888# 0.034573f
C681 source.n12 a_n2044_n5888# 0.015487f
C682 source.n13 a_n2044_n5888# 0.02722f
C683 source.n14 a_n2044_n5888# 0.014627f
C684 source.n15 a_n2044_n5888# 0.034573f
C685 source.n16 a_n2044_n5888# 0.034573f
C686 source.n17 a_n2044_n5888# 0.015487f
C687 source.n18 a_n2044_n5888# 0.02722f
C688 source.n19 a_n2044_n5888# 0.014627f
C689 source.n20 a_n2044_n5888# 0.034573f
C690 source.n21 a_n2044_n5888# 0.015487f
C691 source.n22 a_n2044_n5888# 0.02722f
C692 source.n23 a_n2044_n5888# 0.014627f
C693 source.n24 a_n2044_n5888# 0.034573f
C694 source.n25 a_n2044_n5888# 0.015487f
C695 source.n26 a_n2044_n5888# 0.02722f
C696 source.n27 a_n2044_n5888# 0.014627f
C697 source.n28 a_n2044_n5888# 0.034573f
C698 source.n29 a_n2044_n5888# 0.015487f
C699 source.n30 a_n2044_n5888# 0.02722f
C700 source.n31 a_n2044_n5888# 0.014627f
C701 source.n32 a_n2044_n5888# 0.034573f
C702 source.n33 a_n2044_n5888# 0.015487f
C703 source.n34 a_n2044_n5888# 0.02722f
C704 source.n35 a_n2044_n5888# 0.015057f
C705 source.n36 a_n2044_n5888# 0.034573f
C706 source.n37 a_n2044_n5888# 0.014627f
C707 source.n38 a_n2044_n5888# 0.015487f
C708 source.n39 a_n2044_n5888# 0.02722f
C709 source.n40 a_n2044_n5888# 0.014627f
C710 source.n41 a_n2044_n5888# 0.034573f
C711 source.n42 a_n2044_n5888# 0.015487f
C712 source.n43 a_n2044_n5888# 0.02722f
C713 source.n44 a_n2044_n5888# 0.014627f
C714 source.n45 a_n2044_n5888# 0.025929f
C715 source.n46 a_n2044_n5888# 0.02444f
C716 source.t5 a_n2044_n5888# 0.060297f
C717 source.n47 a_n2044_n5888# 0.332108f
C718 source.n48 a_n2044_n5888# 2.94713f
C719 source.n49 a_n2044_n5888# 0.014627f
C720 source.n50 a_n2044_n5888# 0.015487f
C721 source.n51 a_n2044_n5888# 0.034573f
C722 source.n52 a_n2044_n5888# 0.034573f
C723 source.n53 a_n2044_n5888# 0.015487f
C724 source.n54 a_n2044_n5888# 0.014627f
C725 source.n55 a_n2044_n5888# 0.02722f
C726 source.n56 a_n2044_n5888# 0.02722f
C727 source.n57 a_n2044_n5888# 0.014627f
C728 source.n58 a_n2044_n5888# 0.015487f
C729 source.n59 a_n2044_n5888# 0.034573f
C730 source.n60 a_n2044_n5888# 0.034573f
C731 source.n61 a_n2044_n5888# 0.015487f
C732 source.n62 a_n2044_n5888# 0.014627f
C733 source.n63 a_n2044_n5888# 0.02722f
C734 source.n64 a_n2044_n5888# 0.02722f
C735 source.n65 a_n2044_n5888# 0.014627f
C736 source.n66 a_n2044_n5888# 0.015487f
C737 source.n67 a_n2044_n5888# 0.034573f
C738 source.n68 a_n2044_n5888# 0.034573f
C739 source.n69 a_n2044_n5888# 0.034573f
C740 source.n70 a_n2044_n5888# 0.015057f
C741 source.n71 a_n2044_n5888# 0.014627f
C742 source.n72 a_n2044_n5888# 0.02722f
C743 source.n73 a_n2044_n5888# 0.02722f
C744 source.n74 a_n2044_n5888# 0.014627f
C745 source.n75 a_n2044_n5888# 0.015487f
C746 source.n76 a_n2044_n5888# 0.034573f
C747 source.n77 a_n2044_n5888# 0.034573f
C748 source.n78 a_n2044_n5888# 0.015487f
C749 source.n79 a_n2044_n5888# 0.014627f
C750 source.n80 a_n2044_n5888# 0.02722f
C751 source.n81 a_n2044_n5888# 0.02722f
C752 source.n82 a_n2044_n5888# 0.014627f
C753 source.n83 a_n2044_n5888# 0.015487f
C754 source.n84 a_n2044_n5888# 0.034573f
C755 source.n85 a_n2044_n5888# 0.034573f
C756 source.n86 a_n2044_n5888# 0.015487f
C757 source.n87 a_n2044_n5888# 0.014627f
C758 source.n88 a_n2044_n5888# 0.02722f
C759 source.n89 a_n2044_n5888# 0.02722f
C760 source.n90 a_n2044_n5888# 0.014627f
C761 source.n91 a_n2044_n5888# 0.015487f
C762 source.n92 a_n2044_n5888# 0.034573f
C763 source.n93 a_n2044_n5888# 0.034573f
C764 source.n94 a_n2044_n5888# 0.015487f
C765 source.n95 a_n2044_n5888# 0.014627f
C766 source.n96 a_n2044_n5888# 0.02722f
C767 source.n97 a_n2044_n5888# 0.02722f
C768 source.n98 a_n2044_n5888# 0.014627f
C769 source.n99 a_n2044_n5888# 0.015487f
C770 source.n100 a_n2044_n5888# 0.034573f
C771 source.n101 a_n2044_n5888# 0.034573f
C772 source.n102 a_n2044_n5888# 0.015487f
C773 source.n103 a_n2044_n5888# 0.014627f
C774 source.n104 a_n2044_n5888# 0.02722f
C775 source.n105 a_n2044_n5888# 0.02722f
C776 source.n106 a_n2044_n5888# 0.014627f
C777 source.n107 a_n2044_n5888# 0.015487f
C778 source.n108 a_n2044_n5888# 0.034573f
C779 source.n109 a_n2044_n5888# 0.034573f
C780 source.n110 a_n2044_n5888# 0.015487f
C781 source.n111 a_n2044_n5888# 0.014627f
C782 source.n112 a_n2044_n5888# 0.02722f
C783 source.n113 a_n2044_n5888# 0.02722f
C784 source.n114 a_n2044_n5888# 0.014627f
C785 source.n115 a_n2044_n5888# 0.015057f
C786 source.n116 a_n2044_n5888# 0.015057f
C787 source.n117 a_n2044_n5888# 0.034573f
C788 source.n118 a_n2044_n5888# 0.034573f
C789 source.n119 a_n2044_n5888# 0.015487f
C790 source.n120 a_n2044_n5888# 0.014627f
C791 source.n121 a_n2044_n5888# 0.02722f
C792 source.n122 a_n2044_n5888# 0.02722f
C793 source.n123 a_n2044_n5888# 0.014627f
C794 source.n124 a_n2044_n5888# 0.015487f
C795 source.n125 a_n2044_n5888# 0.034573f
C796 source.n126 a_n2044_n5888# 0.034573f
C797 source.n127 a_n2044_n5888# 0.015487f
C798 source.n128 a_n2044_n5888# 0.014627f
C799 source.n129 a_n2044_n5888# 0.02722f
C800 source.n130 a_n2044_n5888# 0.02722f
C801 source.n131 a_n2044_n5888# 0.014627f
C802 source.n132 a_n2044_n5888# 0.015487f
C803 source.n133 a_n2044_n5888# 0.034573f
C804 source.n134 a_n2044_n5888# 0.073545f
C805 source.n135 a_n2044_n5888# 0.015487f
C806 source.n136 a_n2044_n5888# 0.014627f
C807 source.n137 a_n2044_n5888# 0.059943f
C808 source.n138 a_n2044_n5888# 0.040924f
C809 source.n139 a_n2044_n5888# 2.1627f
C810 source.t0 a_n2044_n5888# 0.537754f
C811 source.t11 a_n2044_n5888# 0.537754f
C812 source.n140 a_n2044_n5888# 4.86675f
C813 source.n141 a_n2044_n5888# 0.407841f
C814 source.t8 a_n2044_n5888# 0.537754f
C815 source.t7 a_n2044_n5888# 0.537754f
C816 source.n142 a_n2044_n5888# 4.86675f
C817 source.n143 a_n2044_n5888# 0.407841f
C818 source.t13 a_n2044_n5888# 0.537754f
C819 source.t9 a_n2044_n5888# 0.537754f
C820 source.n144 a_n2044_n5888# 4.86675f
C821 source.n145 a_n2044_n5888# 0.417671f
C822 source.n146 a_n2044_n5888# 0.037526f
C823 source.n147 a_n2044_n5888# 0.02722f
C824 source.n148 a_n2044_n5888# 0.014627f
C825 source.n149 a_n2044_n5888# 0.034573f
C826 source.n150 a_n2044_n5888# 0.015487f
C827 source.n151 a_n2044_n5888# 0.02722f
C828 source.n152 a_n2044_n5888# 0.014627f
C829 source.n153 a_n2044_n5888# 0.034573f
C830 source.n154 a_n2044_n5888# 0.015487f
C831 source.n155 a_n2044_n5888# 0.02722f
C832 source.n156 a_n2044_n5888# 0.014627f
C833 source.n157 a_n2044_n5888# 0.034573f
C834 source.n158 a_n2044_n5888# 0.015487f
C835 source.n159 a_n2044_n5888# 0.02722f
C836 source.n160 a_n2044_n5888# 0.014627f
C837 source.n161 a_n2044_n5888# 0.034573f
C838 source.n162 a_n2044_n5888# 0.034573f
C839 source.n163 a_n2044_n5888# 0.015487f
C840 source.n164 a_n2044_n5888# 0.02722f
C841 source.n165 a_n2044_n5888# 0.014627f
C842 source.n166 a_n2044_n5888# 0.034573f
C843 source.n167 a_n2044_n5888# 0.015487f
C844 source.n168 a_n2044_n5888# 0.02722f
C845 source.n169 a_n2044_n5888# 0.014627f
C846 source.n170 a_n2044_n5888# 0.034573f
C847 source.n171 a_n2044_n5888# 0.015487f
C848 source.n172 a_n2044_n5888# 0.02722f
C849 source.n173 a_n2044_n5888# 0.014627f
C850 source.n174 a_n2044_n5888# 0.034573f
C851 source.n175 a_n2044_n5888# 0.015487f
C852 source.n176 a_n2044_n5888# 0.02722f
C853 source.n177 a_n2044_n5888# 0.014627f
C854 source.n178 a_n2044_n5888# 0.034573f
C855 source.n179 a_n2044_n5888# 0.015487f
C856 source.n180 a_n2044_n5888# 0.02722f
C857 source.n181 a_n2044_n5888# 0.015057f
C858 source.n182 a_n2044_n5888# 0.034573f
C859 source.n183 a_n2044_n5888# 0.014627f
C860 source.n184 a_n2044_n5888# 0.015487f
C861 source.n185 a_n2044_n5888# 0.02722f
C862 source.n186 a_n2044_n5888# 0.014627f
C863 source.n187 a_n2044_n5888# 0.034573f
C864 source.n188 a_n2044_n5888# 0.015487f
C865 source.n189 a_n2044_n5888# 0.02722f
C866 source.n190 a_n2044_n5888# 0.014627f
C867 source.n191 a_n2044_n5888# 0.025929f
C868 source.n192 a_n2044_n5888# 0.02444f
C869 source.t22 a_n2044_n5888# 0.060297f
C870 source.n193 a_n2044_n5888# 0.332108f
C871 source.n194 a_n2044_n5888# 2.94713f
C872 source.n195 a_n2044_n5888# 0.014627f
C873 source.n196 a_n2044_n5888# 0.015487f
C874 source.n197 a_n2044_n5888# 0.034573f
C875 source.n198 a_n2044_n5888# 0.034573f
C876 source.n199 a_n2044_n5888# 0.015487f
C877 source.n200 a_n2044_n5888# 0.014627f
C878 source.n201 a_n2044_n5888# 0.02722f
C879 source.n202 a_n2044_n5888# 0.02722f
C880 source.n203 a_n2044_n5888# 0.014627f
C881 source.n204 a_n2044_n5888# 0.015487f
C882 source.n205 a_n2044_n5888# 0.034573f
C883 source.n206 a_n2044_n5888# 0.034573f
C884 source.n207 a_n2044_n5888# 0.015487f
C885 source.n208 a_n2044_n5888# 0.014627f
C886 source.n209 a_n2044_n5888# 0.02722f
C887 source.n210 a_n2044_n5888# 0.02722f
C888 source.n211 a_n2044_n5888# 0.014627f
C889 source.n212 a_n2044_n5888# 0.015487f
C890 source.n213 a_n2044_n5888# 0.034573f
C891 source.n214 a_n2044_n5888# 0.034573f
C892 source.n215 a_n2044_n5888# 0.034573f
C893 source.n216 a_n2044_n5888# 0.015057f
C894 source.n217 a_n2044_n5888# 0.014627f
C895 source.n218 a_n2044_n5888# 0.02722f
C896 source.n219 a_n2044_n5888# 0.02722f
C897 source.n220 a_n2044_n5888# 0.014627f
C898 source.n221 a_n2044_n5888# 0.015487f
C899 source.n222 a_n2044_n5888# 0.034573f
C900 source.n223 a_n2044_n5888# 0.034573f
C901 source.n224 a_n2044_n5888# 0.015487f
C902 source.n225 a_n2044_n5888# 0.014627f
C903 source.n226 a_n2044_n5888# 0.02722f
C904 source.n227 a_n2044_n5888# 0.02722f
C905 source.n228 a_n2044_n5888# 0.014627f
C906 source.n229 a_n2044_n5888# 0.015487f
C907 source.n230 a_n2044_n5888# 0.034573f
C908 source.n231 a_n2044_n5888# 0.034573f
C909 source.n232 a_n2044_n5888# 0.015487f
C910 source.n233 a_n2044_n5888# 0.014627f
C911 source.n234 a_n2044_n5888# 0.02722f
C912 source.n235 a_n2044_n5888# 0.02722f
C913 source.n236 a_n2044_n5888# 0.014627f
C914 source.n237 a_n2044_n5888# 0.015487f
C915 source.n238 a_n2044_n5888# 0.034573f
C916 source.n239 a_n2044_n5888# 0.034573f
C917 source.n240 a_n2044_n5888# 0.015487f
C918 source.n241 a_n2044_n5888# 0.014627f
C919 source.n242 a_n2044_n5888# 0.02722f
C920 source.n243 a_n2044_n5888# 0.02722f
C921 source.n244 a_n2044_n5888# 0.014627f
C922 source.n245 a_n2044_n5888# 0.015487f
C923 source.n246 a_n2044_n5888# 0.034573f
C924 source.n247 a_n2044_n5888# 0.034573f
C925 source.n248 a_n2044_n5888# 0.015487f
C926 source.n249 a_n2044_n5888# 0.014627f
C927 source.n250 a_n2044_n5888# 0.02722f
C928 source.n251 a_n2044_n5888# 0.02722f
C929 source.n252 a_n2044_n5888# 0.014627f
C930 source.n253 a_n2044_n5888# 0.015487f
C931 source.n254 a_n2044_n5888# 0.034573f
C932 source.n255 a_n2044_n5888# 0.034573f
C933 source.n256 a_n2044_n5888# 0.015487f
C934 source.n257 a_n2044_n5888# 0.014627f
C935 source.n258 a_n2044_n5888# 0.02722f
C936 source.n259 a_n2044_n5888# 0.02722f
C937 source.n260 a_n2044_n5888# 0.014627f
C938 source.n261 a_n2044_n5888# 0.015057f
C939 source.n262 a_n2044_n5888# 0.015057f
C940 source.n263 a_n2044_n5888# 0.034573f
C941 source.n264 a_n2044_n5888# 0.034573f
C942 source.n265 a_n2044_n5888# 0.015487f
C943 source.n266 a_n2044_n5888# 0.014627f
C944 source.n267 a_n2044_n5888# 0.02722f
C945 source.n268 a_n2044_n5888# 0.02722f
C946 source.n269 a_n2044_n5888# 0.014627f
C947 source.n270 a_n2044_n5888# 0.015487f
C948 source.n271 a_n2044_n5888# 0.034573f
C949 source.n272 a_n2044_n5888# 0.034573f
C950 source.n273 a_n2044_n5888# 0.015487f
C951 source.n274 a_n2044_n5888# 0.014627f
C952 source.n275 a_n2044_n5888# 0.02722f
C953 source.n276 a_n2044_n5888# 0.02722f
C954 source.n277 a_n2044_n5888# 0.014627f
C955 source.n278 a_n2044_n5888# 0.015487f
C956 source.n279 a_n2044_n5888# 0.034573f
C957 source.n280 a_n2044_n5888# 0.073545f
C958 source.n281 a_n2044_n5888# 0.015487f
C959 source.n282 a_n2044_n5888# 0.014627f
C960 source.n283 a_n2044_n5888# 0.059943f
C961 source.n284 a_n2044_n5888# 0.040924f
C962 source.n285 a_n2044_n5888# 0.156916f
C963 source.t15 a_n2044_n5888# 0.537754f
C964 source.t18 a_n2044_n5888# 0.537754f
C965 source.n286 a_n2044_n5888# 4.86675f
C966 source.n287 a_n2044_n5888# 0.407841f
C967 source.t19 a_n2044_n5888# 0.537754f
C968 source.t16 a_n2044_n5888# 0.537754f
C969 source.n288 a_n2044_n5888# 4.86675f
C970 source.n289 a_n2044_n5888# 0.407841f
C971 source.t27 a_n2044_n5888# 0.537754f
C972 source.t14 a_n2044_n5888# 0.537754f
C973 source.n290 a_n2044_n5888# 4.86675f
C974 source.n291 a_n2044_n5888# 2.99661f
C975 source.t2 a_n2044_n5888# 0.537754f
C976 source.t6 a_n2044_n5888# 0.537754f
C977 source.n292 a_n2044_n5888# 4.86675f
C978 source.n293 a_n2044_n5888# 2.99661f
C979 source.t4 a_n2044_n5888# 0.537754f
C980 source.t12 a_n2044_n5888# 0.537754f
C981 source.n294 a_n2044_n5888# 4.86675f
C982 source.n295 a_n2044_n5888# 0.407843f
C983 source.t10 a_n2044_n5888# 0.537754f
C984 source.t3 a_n2044_n5888# 0.537754f
C985 source.n296 a_n2044_n5888# 4.86675f
C986 source.n297 a_n2044_n5888# 0.407843f
C987 source.n298 a_n2044_n5888# 0.037526f
C988 source.n299 a_n2044_n5888# 0.02722f
C989 source.n300 a_n2044_n5888# 0.014627f
C990 source.n301 a_n2044_n5888# 0.034573f
C991 source.n302 a_n2044_n5888# 0.015487f
C992 source.n303 a_n2044_n5888# 0.02722f
C993 source.n304 a_n2044_n5888# 0.014627f
C994 source.n305 a_n2044_n5888# 0.034573f
C995 source.n306 a_n2044_n5888# 0.015487f
C996 source.n307 a_n2044_n5888# 0.02722f
C997 source.n308 a_n2044_n5888# 0.014627f
C998 source.n309 a_n2044_n5888# 0.034573f
C999 source.n310 a_n2044_n5888# 0.015487f
C1000 source.n311 a_n2044_n5888# 0.02722f
C1001 source.n312 a_n2044_n5888# 0.014627f
C1002 source.n313 a_n2044_n5888# 0.034573f
C1003 source.n314 a_n2044_n5888# 0.015487f
C1004 source.n315 a_n2044_n5888# 0.02722f
C1005 source.n316 a_n2044_n5888# 0.014627f
C1006 source.n317 a_n2044_n5888# 0.034573f
C1007 source.n318 a_n2044_n5888# 0.015487f
C1008 source.n319 a_n2044_n5888# 0.02722f
C1009 source.n320 a_n2044_n5888# 0.014627f
C1010 source.n321 a_n2044_n5888# 0.034573f
C1011 source.n322 a_n2044_n5888# 0.015487f
C1012 source.n323 a_n2044_n5888# 0.02722f
C1013 source.n324 a_n2044_n5888# 0.014627f
C1014 source.n325 a_n2044_n5888# 0.034573f
C1015 source.n326 a_n2044_n5888# 0.015487f
C1016 source.n327 a_n2044_n5888# 0.02722f
C1017 source.n328 a_n2044_n5888# 0.014627f
C1018 source.n329 a_n2044_n5888# 0.034573f
C1019 source.n330 a_n2044_n5888# 0.015487f
C1020 source.n331 a_n2044_n5888# 0.02722f
C1021 source.n332 a_n2044_n5888# 0.015057f
C1022 source.n333 a_n2044_n5888# 0.034573f
C1023 source.n334 a_n2044_n5888# 0.015487f
C1024 source.n335 a_n2044_n5888# 0.02722f
C1025 source.n336 a_n2044_n5888# 0.014627f
C1026 source.n337 a_n2044_n5888# 0.034573f
C1027 source.n338 a_n2044_n5888# 0.015487f
C1028 source.n339 a_n2044_n5888# 0.02722f
C1029 source.n340 a_n2044_n5888# 0.014627f
C1030 source.n341 a_n2044_n5888# 0.025929f
C1031 source.n342 a_n2044_n5888# 0.02444f
C1032 source.t1 a_n2044_n5888# 0.060297f
C1033 source.n343 a_n2044_n5888# 0.332108f
C1034 source.n344 a_n2044_n5888# 2.94714f
C1035 source.n345 a_n2044_n5888# 0.014627f
C1036 source.n346 a_n2044_n5888# 0.015487f
C1037 source.n347 a_n2044_n5888# 0.034573f
C1038 source.n348 a_n2044_n5888# 0.034573f
C1039 source.n349 a_n2044_n5888# 0.015487f
C1040 source.n350 a_n2044_n5888# 0.014627f
C1041 source.n351 a_n2044_n5888# 0.02722f
C1042 source.n352 a_n2044_n5888# 0.02722f
C1043 source.n353 a_n2044_n5888# 0.014627f
C1044 source.n354 a_n2044_n5888# 0.015487f
C1045 source.n355 a_n2044_n5888# 0.034573f
C1046 source.n356 a_n2044_n5888# 0.034573f
C1047 source.n357 a_n2044_n5888# 0.015487f
C1048 source.n358 a_n2044_n5888# 0.014627f
C1049 source.n359 a_n2044_n5888# 0.02722f
C1050 source.n360 a_n2044_n5888# 0.02722f
C1051 source.n361 a_n2044_n5888# 0.014627f
C1052 source.n362 a_n2044_n5888# 0.014627f
C1053 source.n363 a_n2044_n5888# 0.015487f
C1054 source.n364 a_n2044_n5888# 0.034573f
C1055 source.n365 a_n2044_n5888# 0.034573f
C1056 source.n366 a_n2044_n5888# 0.034573f
C1057 source.n367 a_n2044_n5888# 0.015057f
C1058 source.n368 a_n2044_n5888# 0.014627f
C1059 source.n369 a_n2044_n5888# 0.02722f
C1060 source.n370 a_n2044_n5888# 0.02722f
C1061 source.n371 a_n2044_n5888# 0.014627f
C1062 source.n372 a_n2044_n5888# 0.015487f
C1063 source.n373 a_n2044_n5888# 0.034573f
C1064 source.n374 a_n2044_n5888# 0.034573f
C1065 source.n375 a_n2044_n5888# 0.015487f
C1066 source.n376 a_n2044_n5888# 0.014627f
C1067 source.n377 a_n2044_n5888# 0.02722f
C1068 source.n378 a_n2044_n5888# 0.02722f
C1069 source.n379 a_n2044_n5888# 0.014627f
C1070 source.n380 a_n2044_n5888# 0.015487f
C1071 source.n381 a_n2044_n5888# 0.034573f
C1072 source.n382 a_n2044_n5888# 0.034573f
C1073 source.n383 a_n2044_n5888# 0.015487f
C1074 source.n384 a_n2044_n5888# 0.014627f
C1075 source.n385 a_n2044_n5888# 0.02722f
C1076 source.n386 a_n2044_n5888# 0.02722f
C1077 source.n387 a_n2044_n5888# 0.014627f
C1078 source.n388 a_n2044_n5888# 0.015487f
C1079 source.n389 a_n2044_n5888# 0.034573f
C1080 source.n390 a_n2044_n5888# 0.034573f
C1081 source.n391 a_n2044_n5888# 0.015487f
C1082 source.n392 a_n2044_n5888# 0.014627f
C1083 source.n393 a_n2044_n5888# 0.02722f
C1084 source.n394 a_n2044_n5888# 0.02722f
C1085 source.n395 a_n2044_n5888# 0.014627f
C1086 source.n396 a_n2044_n5888# 0.015487f
C1087 source.n397 a_n2044_n5888# 0.034573f
C1088 source.n398 a_n2044_n5888# 0.034573f
C1089 source.n399 a_n2044_n5888# 0.015487f
C1090 source.n400 a_n2044_n5888# 0.014627f
C1091 source.n401 a_n2044_n5888# 0.02722f
C1092 source.n402 a_n2044_n5888# 0.02722f
C1093 source.n403 a_n2044_n5888# 0.014627f
C1094 source.n404 a_n2044_n5888# 0.015487f
C1095 source.n405 a_n2044_n5888# 0.034573f
C1096 source.n406 a_n2044_n5888# 0.034573f
C1097 source.n407 a_n2044_n5888# 0.034573f
C1098 source.n408 a_n2044_n5888# 0.015487f
C1099 source.n409 a_n2044_n5888# 0.014627f
C1100 source.n410 a_n2044_n5888# 0.02722f
C1101 source.n411 a_n2044_n5888# 0.02722f
C1102 source.n412 a_n2044_n5888# 0.014627f
C1103 source.n413 a_n2044_n5888# 0.015057f
C1104 source.n414 a_n2044_n5888# 0.015057f
C1105 source.n415 a_n2044_n5888# 0.034573f
C1106 source.n416 a_n2044_n5888# 0.034573f
C1107 source.n417 a_n2044_n5888# 0.015487f
C1108 source.n418 a_n2044_n5888# 0.014627f
C1109 source.n419 a_n2044_n5888# 0.02722f
C1110 source.n420 a_n2044_n5888# 0.02722f
C1111 source.n421 a_n2044_n5888# 0.014627f
C1112 source.n422 a_n2044_n5888# 0.015487f
C1113 source.n423 a_n2044_n5888# 0.034573f
C1114 source.n424 a_n2044_n5888# 0.034573f
C1115 source.n425 a_n2044_n5888# 0.015487f
C1116 source.n426 a_n2044_n5888# 0.014627f
C1117 source.n427 a_n2044_n5888# 0.02722f
C1118 source.n428 a_n2044_n5888# 0.02722f
C1119 source.n429 a_n2044_n5888# 0.014627f
C1120 source.n430 a_n2044_n5888# 0.015487f
C1121 source.n431 a_n2044_n5888# 0.034573f
C1122 source.n432 a_n2044_n5888# 0.073545f
C1123 source.n433 a_n2044_n5888# 0.015487f
C1124 source.n434 a_n2044_n5888# 0.014627f
C1125 source.n435 a_n2044_n5888# 0.059943f
C1126 source.n436 a_n2044_n5888# 0.040924f
C1127 source.n437 a_n2044_n5888# 0.156916f
C1128 source.t20 a_n2044_n5888# 0.537754f
C1129 source.t26 a_n2044_n5888# 0.537754f
C1130 source.n438 a_n2044_n5888# 4.86675f
C1131 source.n439 a_n2044_n5888# 0.417673f
C1132 source.t23 a_n2044_n5888# 0.537754f
C1133 source.t24 a_n2044_n5888# 0.537754f
C1134 source.n440 a_n2044_n5888# 4.86675f
C1135 source.n441 a_n2044_n5888# 0.407843f
C1136 source.t17 a_n2044_n5888# 0.537754f
C1137 source.t25 a_n2044_n5888# 0.537754f
C1138 source.n442 a_n2044_n5888# 4.86675f
C1139 source.n443 a_n2044_n5888# 0.407843f
C1140 source.n444 a_n2044_n5888# 0.037526f
C1141 source.n445 a_n2044_n5888# 0.02722f
C1142 source.n446 a_n2044_n5888# 0.014627f
C1143 source.n447 a_n2044_n5888# 0.034573f
C1144 source.n448 a_n2044_n5888# 0.015487f
C1145 source.n449 a_n2044_n5888# 0.02722f
C1146 source.n450 a_n2044_n5888# 0.014627f
C1147 source.n451 a_n2044_n5888# 0.034573f
C1148 source.n452 a_n2044_n5888# 0.015487f
C1149 source.n453 a_n2044_n5888# 0.02722f
C1150 source.n454 a_n2044_n5888# 0.014627f
C1151 source.n455 a_n2044_n5888# 0.034573f
C1152 source.n456 a_n2044_n5888# 0.015487f
C1153 source.n457 a_n2044_n5888# 0.02722f
C1154 source.n458 a_n2044_n5888# 0.014627f
C1155 source.n459 a_n2044_n5888# 0.034573f
C1156 source.n460 a_n2044_n5888# 0.015487f
C1157 source.n461 a_n2044_n5888# 0.02722f
C1158 source.n462 a_n2044_n5888# 0.014627f
C1159 source.n463 a_n2044_n5888# 0.034573f
C1160 source.n464 a_n2044_n5888# 0.015487f
C1161 source.n465 a_n2044_n5888# 0.02722f
C1162 source.n466 a_n2044_n5888# 0.014627f
C1163 source.n467 a_n2044_n5888# 0.034573f
C1164 source.n468 a_n2044_n5888# 0.015487f
C1165 source.n469 a_n2044_n5888# 0.02722f
C1166 source.n470 a_n2044_n5888# 0.014627f
C1167 source.n471 a_n2044_n5888# 0.034573f
C1168 source.n472 a_n2044_n5888# 0.015487f
C1169 source.n473 a_n2044_n5888# 0.02722f
C1170 source.n474 a_n2044_n5888# 0.014627f
C1171 source.n475 a_n2044_n5888# 0.034573f
C1172 source.n476 a_n2044_n5888# 0.015487f
C1173 source.n477 a_n2044_n5888# 0.02722f
C1174 source.n478 a_n2044_n5888# 0.015057f
C1175 source.n479 a_n2044_n5888# 0.034573f
C1176 source.n480 a_n2044_n5888# 0.015487f
C1177 source.n481 a_n2044_n5888# 0.02722f
C1178 source.n482 a_n2044_n5888# 0.014627f
C1179 source.n483 a_n2044_n5888# 0.034573f
C1180 source.n484 a_n2044_n5888# 0.015487f
C1181 source.n485 a_n2044_n5888# 0.02722f
C1182 source.n486 a_n2044_n5888# 0.014627f
C1183 source.n487 a_n2044_n5888# 0.025929f
C1184 source.n488 a_n2044_n5888# 0.02444f
C1185 source.t21 a_n2044_n5888# 0.060297f
C1186 source.n489 a_n2044_n5888# 0.332108f
C1187 source.n490 a_n2044_n5888# 2.94714f
C1188 source.n491 a_n2044_n5888# 0.014627f
C1189 source.n492 a_n2044_n5888# 0.015487f
C1190 source.n493 a_n2044_n5888# 0.034573f
C1191 source.n494 a_n2044_n5888# 0.034573f
C1192 source.n495 a_n2044_n5888# 0.015487f
C1193 source.n496 a_n2044_n5888# 0.014627f
C1194 source.n497 a_n2044_n5888# 0.02722f
C1195 source.n498 a_n2044_n5888# 0.02722f
C1196 source.n499 a_n2044_n5888# 0.014627f
C1197 source.n500 a_n2044_n5888# 0.015487f
C1198 source.n501 a_n2044_n5888# 0.034573f
C1199 source.n502 a_n2044_n5888# 0.034573f
C1200 source.n503 a_n2044_n5888# 0.015487f
C1201 source.n504 a_n2044_n5888# 0.014627f
C1202 source.n505 a_n2044_n5888# 0.02722f
C1203 source.n506 a_n2044_n5888# 0.02722f
C1204 source.n507 a_n2044_n5888# 0.014627f
C1205 source.n508 a_n2044_n5888# 0.014627f
C1206 source.n509 a_n2044_n5888# 0.015487f
C1207 source.n510 a_n2044_n5888# 0.034573f
C1208 source.n511 a_n2044_n5888# 0.034573f
C1209 source.n512 a_n2044_n5888# 0.034573f
C1210 source.n513 a_n2044_n5888# 0.015057f
C1211 source.n514 a_n2044_n5888# 0.014627f
C1212 source.n515 a_n2044_n5888# 0.02722f
C1213 source.n516 a_n2044_n5888# 0.02722f
C1214 source.n517 a_n2044_n5888# 0.014627f
C1215 source.n518 a_n2044_n5888# 0.015487f
C1216 source.n519 a_n2044_n5888# 0.034573f
C1217 source.n520 a_n2044_n5888# 0.034573f
C1218 source.n521 a_n2044_n5888# 0.015487f
C1219 source.n522 a_n2044_n5888# 0.014627f
C1220 source.n523 a_n2044_n5888# 0.02722f
C1221 source.n524 a_n2044_n5888# 0.02722f
C1222 source.n525 a_n2044_n5888# 0.014627f
C1223 source.n526 a_n2044_n5888# 0.015487f
C1224 source.n527 a_n2044_n5888# 0.034573f
C1225 source.n528 a_n2044_n5888# 0.034573f
C1226 source.n529 a_n2044_n5888# 0.015487f
C1227 source.n530 a_n2044_n5888# 0.014627f
C1228 source.n531 a_n2044_n5888# 0.02722f
C1229 source.n532 a_n2044_n5888# 0.02722f
C1230 source.n533 a_n2044_n5888# 0.014627f
C1231 source.n534 a_n2044_n5888# 0.015487f
C1232 source.n535 a_n2044_n5888# 0.034573f
C1233 source.n536 a_n2044_n5888# 0.034573f
C1234 source.n537 a_n2044_n5888# 0.015487f
C1235 source.n538 a_n2044_n5888# 0.014627f
C1236 source.n539 a_n2044_n5888# 0.02722f
C1237 source.n540 a_n2044_n5888# 0.02722f
C1238 source.n541 a_n2044_n5888# 0.014627f
C1239 source.n542 a_n2044_n5888# 0.015487f
C1240 source.n543 a_n2044_n5888# 0.034573f
C1241 source.n544 a_n2044_n5888# 0.034573f
C1242 source.n545 a_n2044_n5888# 0.015487f
C1243 source.n546 a_n2044_n5888# 0.014627f
C1244 source.n547 a_n2044_n5888# 0.02722f
C1245 source.n548 a_n2044_n5888# 0.02722f
C1246 source.n549 a_n2044_n5888# 0.014627f
C1247 source.n550 a_n2044_n5888# 0.015487f
C1248 source.n551 a_n2044_n5888# 0.034573f
C1249 source.n552 a_n2044_n5888# 0.034573f
C1250 source.n553 a_n2044_n5888# 0.034573f
C1251 source.n554 a_n2044_n5888# 0.015487f
C1252 source.n555 a_n2044_n5888# 0.014627f
C1253 source.n556 a_n2044_n5888# 0.02722f
C1254 source.n557 a_n2044_n5888# 0.02722f
C1255 source.n558 a_n2044_n5888# 0.014627f
C1256 source.n559 a_n2044_n5888# 0.015057f
C1257 source.n560 a_n2044_n5888# 0.015057f
C1258 source.n561 a_n2044_n5888# 0.034573f
C1259 source.n562 a_n2044_n5888# 0.034573f
C1260 source.n563 a_n2044_n5888# 0.015487f
C1261 source.n564 a_n2044_n5888# 0.014627f
C1262 source.n565 a_n2044_n5888# 0.02722f
C1263 source.n566 a_n2044_n5888# 0.02722f
C1264 source.n567 a_n2044_n5888# 0.014627f
C1265 source.n568 a_n2044_n5888# 0.015487f
C1266 source.n569 a_n2044_n5888# 0.034573f
C1267 source.n570 a_n2044_n5888# 0.034573f
C1268 source.n571 a_n2044_n5888# 0.015487f
C1269 source.n572 a_n2044_n5888# 0.014627f
C1270 source.n573 a_n2044_n5888# 0.02722f
C1271 source.n574 a_n2044_n5888# 0.02722f
C1272 source.n575 a_n2044_n5888# 0.014627f
C1273 source.n576 a_n2044_n5888# 0.015487f
C1274 source.n577 a_n2044_n5888# 0.034573f
C1275 source.n578 a_n2044_n5888# 0.073545f
C1276 source.n579 a_n2044_n5888# 0.015487f
C1277 source.n580 a_n2044_n5888# 0.014627f
C1278 source.n581 a_n2044_n5888# 0.059943f
C1279 source.n582 a_n2044_n5888# 0.040924f
C1280 source.n583 a_n2044_n5888# 0.291212f
C1281 source.n584 a_n2044_n5888# 2.91164f
C1282 minus.n0 a_n2044_n5888# 0.045518f
C1283 minus.t4 a_n2044_n5888# 1.60793f
C1284 minus.n1 a_n2044_n5888# 0.595297f
C1285 minus.n2 a_n2044_n5888# 0.060738f
C1286 minus.t1 a_n2044_n5888# 1.60793f
C1287 minus.n3 a_n2044_n5888# 0.595016f
C1288 minus.t10 a_n2044_n5888# 1.61742f
C1289 minus.n4 a_n2044_n5888# 0.581377f
C1290 minus.n5 a_n2044_n5888# 0.149674f
C1291 minus.n6 a_n2044_n5888# 0.010329f
C1292 minus.t5 a_n2044_n5888# 1.60793f
C1293 minus.n7 a_n2044_n5888# 0.595297f
C1294 minus.t13 a_n2044_n5888# 1.60793f
C1295 minus.n8 a_n2044_n5888# 0.600855f
C1296 minus.n9 a_n2044_n5888# 0.060596f
C1297 minus.n10 a_n2044_n5888# 0.060738f
C1298 minus.n11 a_n2044_n5888# 0.045518f
C1299 minus.n12 a_n2044_n5888# 0.010329f
C1300 minus.t7 a_n2044_n5888# 1.60793f
C1301 minus.n13 a_n2044_n5888# 0.595016f
C1302 minus.t0 a_n2044_n5888# 1.60793f
C1303 minus.n14 a_n2044_n5888# 0.590526f
C1304 minus.n15 a_n2044_n5888# 2.35967f
C1305 minus.n16 a_n2044_n5888# 0.045518f
C1306 minus.t6 a_n2044_n5888# 1.60793f
C1307 minus.n17 a_n2044_n5888# 0.595297f
C1308 minus.n18 a_n2044_n5888# 0.060738f
C1309 minus.t2 a_n2044_n5888# 1.60793f
C1310 minus.n19 a_n2044_n5888# 0.595016f
C1311 minus.t3 a_n2044_n5888# 1.61742f
C1312 minus.n20 a_n2044_n5888# 0.581377f
C1313 minus.n21 a_n2044_n5888# 0.149674f
C1314 minus.n22 a_n2044_n5888# 0.010329f
C1315 minus.t9 a_n2044_n5888# 1.60793f
C1316 minus.n23 a_n2044_n5888# 0.595297f
C1317 minus.t8 a_n2044_n5888# 1.60793f
C1318 minus.n24 a_n2044_n5888# 0.600855f
C1319 minus.n25 a_n2044_n5888# 0.060596f
C1320 minus.n26 a_n2044_n5888# 0.060738f
C1321 minus.n27 a_n2044_n5888# 0.045518f
C1322 minus.n28 a_n2044_n5888# 0.010329f
C1323 minus.t12 a_n2044_n5888# 1.60793f
C1324 minus.n29 a_n2044_n5888# 0.595016f
C1325 minus.t11 a_n2044_n5888# 1.60793f
C1326 minus.n30 a_n2044_n5888# 0.590526f
C1327 minus.n31 a_n2044_n5888# 0.307546f
C1328 minus.n32 a_n2044_n5888# 2.7793f
.ends

