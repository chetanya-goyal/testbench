* NGSPICE file created from diffpair31.ext - technology: sky130A

.subckt diffpair31 minus drain_right drain_left source plus
X0 a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X1 drain_right minus source a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X2 source minus drain_right a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X3 source minus drain_right a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X4 a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X5 source plus drain_left a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X6 a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X7 a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X8 source plus drain_left a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X9 drain_right minus source a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X10 drain_left plus source a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X11 drain_left plus source a_n1094_n1092# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
.ends

