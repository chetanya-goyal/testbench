* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t23 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X1 drain_right.t13 minus.t0 source.t11 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X2 drain_right.t12 minus.t1 source.t1 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 source.t17 plus.t1 drain_left.t12 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X4 a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X5 drain_left.t11 plus.t2 source.t16 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X6 source.t5 minus.t2 drain_right.t11 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X7 drain_left.t10 plus.t3 source.t14 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X8 a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X9 source.t7 minus.t3 drain_right.t10 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 drain_right.t9 minus.t4 source.t0 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 drain_right.t8 minus.t5 source.t8 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X12 drain_right.t7 minus.t6 source.t4 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X13 source.t15 plus.t4 drain_left.t9 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t6 minus.t7 drain_right.t6 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 source.t9 minus.t8 drain_right.t5 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 source.t27 plus.t5 drain_left.t8 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_left.t7 plus.t6 source.t18 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X18 drain_right.t4 minus.t9 source.t3 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 drain_right.t3 minus.t10 source.t12 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X20 a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X21 drain_right.t2 minus.t11 source.t13 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X22 source.t24 plus.t7 drain_left.t6 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X23 source.t2 minus.t12 drain_right.t1 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X24 a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X25 drain_left.t5 plus.t8 source.t21 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X26 drain_left.t4 plus.t9 source.t19 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X27 drain_left.t3 plus.t10 source.t25 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X28 source.t10 minus.t13 drain_right.t0 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X29 source.t22 plus.t11 drain_left.t2 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X30 source.t26 plus.t12 drain_left.t1 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X31 drain_left.t0 plus.t13 source.t20 a_n1756_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
R0 plus.n3 plus.t6 595.928
R1 plus.n15 plus.t9 595.928
R2 plus.n20 plus.t8 595.928
R3 plus.n32 plus.t3 595.928
R4 plus.n1 plus.t7 530.201
R5 plus.n4 plus.t12 530.201
R6 plus.n6 plus.t10 530.201
R7 plus.n12 plus.t13 530.201
R8 plus.n14 plus.t11 530.201
R9 plus.n18 plus.t1 530.201
R10 plus.n21 plus.t5 530.201
R11 plus.n23 plus.t2 530.201
R12 plus.n29 plus.t0 530.201
R13 plus.n31 plus.t4 530.201
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 51.1217
R33 plus.n13 plus.n12 51.1217
R34 plus.n30 plus.n29 51.1217
R35 plus.n23 plus.n22 51.1217
R36 plus.n5 plus.n4 43.8187
R37 plus.n14 plus.n13 43.8187
R38 plus.n31 plus.n30 43.8187
R39 plus.n22 plus.n21 43.8187
R40 plus.n4 plus.n3 29.2126
R41 plus.n15 plus.n14 29.2126
R42 plus.n32 plus.n31 29.2126
R43 plus.n21 plus.n20 29.2126
R44 plus plus.n33 25.9365
R45 plus.n7 plus.n6 21.9096
R46 plus.n12 plus.n11 21.9096
R47 plus.n29 plus.n28 21.9096
R48 plus.n24 plus.n23 21.9096
R49 plus plus.n16 8.42664
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 source.n0 source.t19 99.1169
R61 source.n7 source.t8 99.1169
R62 source.n27 source.t13 99.1168
R63 source.n20 source.t21 99.1168
R64 source.n2 source.n1 84.1169
R65 source.n4 source.n3 84.1169
R66 source.n6 source.n5 84.1169
R67 source.n9 source.n8 84.1169
R68 source.n11 source.n10 84.1169
R69 source.n13 source.n12 84.1169
R70 source.n26 source.n25 84.1168
R71 source.n24 source.n23 84.1168
R72 source.n22 source.n21 84.1168
R73 source.n19 source.n18 84.1168
R74 source.n17 source.n16 84.1168
R75 source.n15 source.n14 84.1168
R76 source.n25 source.t11 15.0005
R77 source.n25 source.t10 15.0005
R78 source.n23 source.t0 15.0005
R79 source.n23 source.t5 15.0005
R80 source.n21 source.t1 15.0005
R81 source.n21 source.t9 15.0005
R82 source.n18 source.t16 15.0005
R83 source.n18 source.t27 15.0005
R84 source.n16 source.t23 15.0005
R85 source.n16 source.t17 15.0005
R86 source.n14 source.t14 15.0005
R87 source.n14 source.t15 15.0005
R88 source.n1 source.t20 15.0005
R89 source.n1 source.t22 15.0005
R90 source.n3 source.t25 15.0005
R91 source.n3 source.t24 15.0005
R92 source.n5 source.t18 15.0005
R93 source.n5 source.t26 15.0005
R94 source.n8 source.t3 15.0005
R95 source.n8 source.t7 15.0005
R96 source.n10 source.t4 15.0005
R97 source.n10 source.t6 15.0005
R98 source.n12 source.t12 15.0005
R99 source.n12 source.t2 15.0005
R100 source.n15 source.n13 14.8327
R101 source.n28 source.n0 8.72921
R102 source.n28 source.n27 5.5436
R103 source.n7 source.n6 0.7505
R104 source.n22 source.n20 0.7505
R105 source.n13 source.n11 0.560845
R106 source.n11 source.n9 0.560845
R107 source.n9 source.n7 0.560845
R108 source.n6 source.n4 0.560845
R109 source.n4 source.n2 0.560845
R110 source.n2 source.n0 0.560845
R111 source.n17 source.n15 0.560845
R112 source.n19 source.n17 0.560845
R113 source.n20 source.n19 0.560845
R114 source.n24 source.n22 0.560845
R115 source.n26 source.n24 0.560845
R116 source.n27 source.n26 0.560845
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t7 116.356
R119 drain_left.n1 drain_left.t10 116.356
R120 drain_left.n4 drain_left.n2 101.356
R121 drain_left.n11 drain_left.n10 100.796
R122 drain_left.n9 drain_left.n8 100.796
R123 drain_left.n7 drain_left.n6 100.796
R124 drain_left.n4 drain_left.n3 100.796
R125 drain_left.n1 drain_left.n0 100.796
R126 drain_left drain_left.n5 23.0133
R127 drain_left.n2 drain_left.t8 15.0005
R128 drain_left.n2 drain_left.t5 15.0005
R129 drain_left.n3 drain_left.t12 15.0005
R130 drain_left.n3 drain_left.t11 15.0005
R131 drain_left.n0 drain_left.t9 15.0005
R132 drain_left.n0 drain_left.t13 15.0005
R133 drain_left.n10 drain_left.t2 15.0005
R134 drain_left.n10 drain_left.t4 15.0005
R135 drain_left.n8 drain_left.t6 15.0005
R136 drain_left.n8 drain_left.t0 15.0005
R137 drain_left.n6 drain_left.t1 15.0005
R138 drain_left.n6 drain_left.t3 15.0005
R139 drain_left drain_left.n11 6.21356
R140 drain_left.n9 drain_left.n7 0.560845
R141 drain_left.n11 drain_left.n9 0.560845
R142 drain_left.n5 drain_left.n1 0.365413
R143 drain_left.n5 drain_left.n4 0.0852402
R144 minus.n15 minus.t10 595.928
R145 minus.n3 minus.t5 595.928
R146 minus.n32 minus.t11 595.928
R147 minus.n20 minus.t1 595.928
R148 minus.n1 minus.t7 530.201
R149 minus.n14 minus.t12 530.201
R150 minus.n12 minus.t6 530.201
R151 minus.n6 minus.t9 530.201
R152 minus.n4 minus.t3 530.201
R153 minus.n18 minus.t2 530.201
R154 minus.n31 minus.t13 530.201
R155 minus.n29 minus.t0 530.201
R156 minus.n23 minus.t4 530.201
R157 minus.n21 minus.t8 530.201
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 51.1217
R177 minus.n6 minus.n5 51.1217
R178 minus.n23 minus.n22 51.1217
R179 minus.n30 minus.n29 51.1217
R180 minus.n14 minus.n13 43.8187
R181 minus.n5 minus.n4 43.8187
R182 minus.n22 minus.n21 43.8187
R183 minus.n31 minus.n30 43.8187
R184 minus.n15 minus.n14 29.2126
R185 minus.n4 minus.n3 29.2126
R186 minus.n21 minus.n20 29.2126
R187 minus.n32 minus.n31 29.2126
R188 minus.n34 minus.n16 28.2675
R189 minus.n12 minus.n11 21.9096
R190 minus.n7 minus.n6 21.9096
R191 minus.n24 minus.n23 21.9096
R192 minus.n29 minus.n28 21.9096
R193 minus.n34 minus.n33 6.57058
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t12 116.356
R206 drain_right.n11 drain_right.t3 115.796
R207 drain_right.n8 drain_right.n6 101.356
R208 drain_right.n4 drain_right.n2 101.356
R209 drain_right.n8 drain_right.n7 100.796
R210 drain_right.n10 drain_right.n9 100.796
R211 drain_right.n4 drain_right.n3 100.796
R212 drain_right.n1 drain_right.n0 100.796
R213 drain_right drain_right.n5 22.4601
R214 drain_right.n2 drain_right.t0 15.0005
R215 drain_right.n2 drain_right.t2 15.0005
R216 drain_right.n3 drain_right.t11 15.0005
R217 drain_right.n3 drain_right.t13 15.0005
R218 drain_right.n0 drain_right.t5 15.0005
R219 drain_right.n0 drain_right.t9 15.0005
R220 drain_right.n6 drain_right.t10 15.0005
R221 drain_right.n6 drain_right.t8 15.0005
R222 drain_right.n7 drain_right.t6 15.0005
R223 drain_right.n7 drain_right.t4 15.0005
R224 drain_right.n9 drain_right.t1 15.0005
R225 drain_right.n9 drain_right.t7 15.0005
R226 drain_right drain_right.n11 5.93339
R227 drain_right.n11 drain_right.n10 0.560845
R228 drain_right.n10 drain_right.n8 0.560845
R229 drain_right.n5 drain_right.n1 0.365413
R230 drain_right.n5 drain_right.n4 0.0852402
C0 drain_right minus 0.916312f
C1 drain_right plus 0.331272f
C2 plus minus 3.48017f
C3 drain_right drain_left 0.897561f
C4 drain_right source 7.00753f
C5 minus drain_left 0.177443f
C6 plus drain_left 1.08588f
C7 minus source 1.0168f
C8 plus source 1.03087f
C9 source drain_left 7.00979f
C10 drain_right a_n1756_n1288# 3.90203f
C11 drain_left a_n1756_n1288# 4.15014f
C12 source a_n1756_n1288# 2.634306f
C13 minus a_n1756_n1288# 5.661115f
C14 plus a_n1756_n1288# 6.451344f
C15 drain_right.t12 a_n1756_n1288# 0.328046f
C16 drain_right.t5 a_n1756_n1288# 0.055405f
C17 drain_right.t9 a_n1756_n1288# 0.055405f
C18 drain_right.n0 a_n1756_n1288# 0.267404f
C19 drain_right.n1 a_n1756_n1288# 0.514814f
C20 drain_right.t0 a_n1756_n1288# 0.055405f
C21 drain_right.t2 a_n1756_n1288# 0.055405f
C22 drain_right.n2 a_n1756_n1288# 0.268896f
C23 drain_right.t11 a_n1756_n1288# 0.055405f
C24 drain_right.t13 a_n1756_n1288# 0.055405f
C25 drain_right.n3 a_n1756_n1288# 0.267404f
C26 drain_right.n4 a_n1756_n1288# 0.499982f
C27 drain_right.n5 a_n1756_n1288# 0.592467f
C28 drain_right.t10 a_n1756_n1288# 0.055405f
C29 drain_right.t8 a_n1756_n1288# 0.055405f
C30 drain_right.n6 a_n1756_n1288# 0.268897f
C31 drain_right.t6 a_n1756_n1288# 0.055405f
C32 drain_right.t4 a_n1756_n1288# 0.055405f
C33 drain_right.n7 a_n1756_n1288# 0.267405f
C34 drain_right.n8 a_n1756_n1288# 0.529108f
C35 drain_right.t1 a_n1756_n1288# 0.055405f
C36 drain_right.t7 a_n1756_n1288# 0.055405f
C37 drain_right.n9 a_n1756_n1288# 0.267405f
C38 drain_right.n10 a_n1756_n1288# 0.260641f
C39 drain_right.t3 a_n1756_n1288# 0.326753f
C40 drain_right.n11 a_n1756_n1288# 0.462577f
C41 minus.n0 a_n1756_n1288# 0.034408f
C42 minus.t10 a_n1756_n1288# 0.033534f
C43 minus.t12 a_n1756_n1288# 0.030375f
C44 minus.t6 a_n1756_n1288# 0.030375f
C45 minus.t7 a_n1756_n1288# 0.030375f
C46 minus.n1 a_n1756_n1288# 0.037932f
C47 minus.n2 a_n1756_n1288# 0.080431f
C48 minus.t9 a_n1756_n1288# 0.030375f
C49 minus.t3 a_n1756_n1288# 0.030375f
C50 minus.t5 a_n1756_n1288# 0.033534f
C51 minus.n3 a_n1756_n1288# 0.040131f
C52 minus.n4 a_n1756_n1288# 0.026518f
C53 minus.n5 a_n1756_n1288# 0.014597f
C54 minus.n6 a_n1756_n1288# 0.026518f
C55 minus.n7 a_n1756_n1288# 0.014597f
C56 minus.n8 a_n1756_n1288# 0.034408f
C57 minus.n9 a_n1756_n1288# 0.034408f
C58 minus.n10 a_n1756_n1288# 0.034408f
C59 minus.n11 a_n1756_n1288# 0.014597f
C60 minus.n12 a_n1756_n1288# 0.026518f
C61 minus.n13 a_n1756_n1288# 0.014597f
C62 minus.n14 a_n1756_n1288# 0.026518f
C63 minus.n15 a_n1756_n1288# 0.040077f
C64 minus.n16 a_n1756_n1288# 0.809779f
C65 minus.n17 a_n1756_n1288# 0.034408f
C66 minus.t13 a_n1756_n1288# 0.030375f
C67 minus.t0 a_n1756_n1288# 0.030375f
C68 minus.t2 a_n1756_n1288# 0.030375f
C69 minus.n18 a_n1756_n1288# 0.037932f
C70 minus.n19 a_n1756_n1288# 0.080431f
C71 minus.t4 a_n1756_n1288# 0.030375f
C72 minus.t8 a_n1756_n1288# 0.030375f
C73 minus.t1 a_n1756_n1288# 0.033534f
C74 minus.n20 a_n1756_n1288# 0.040131f
C75 minus.n21 a_n1756_n1288# 0.026518f
C76 minus.n22 a_n1756_n1288# 0.014597f
C77 minus.n23 a_n1756_n1288# 0.026518f
C78 minus.n24 a_n1756_n1288# 0.014597f
C79 minus.n25 a_n1756_n1288# 0.034408f
C80 minus.n26 a_n1756_n1288# 0.034408f
C81 minus.n27 a_n1756_n1288# 0.034408f
C82 minus.n28 a_n1756_n1288# 0.014597f
C83 minus.n29 a_n1756_n1288# 0.026518f
C84 minus.n30 a_n1756_n1288# 0.014597f
C85 minus.n31 a_n1756_n1288# 0.026518f
C86 minus.t11 a_n1756_n1288# 0.033534f
C87 minus.n32 a_n1756_n1288# 0.040077f
C88 minus.n33 a_n1756_n1288# 0.230656f
C89 minus.n34 a_n1756_n1288# 0.997758f
C90 drain_left.t10 a_n1756_n1288# 0.323858f
C91 drain_left.t9 a_n1756_n1288# 0.054698f
C92 drain_left.t13 a_n1756_n1288# 0.054698f
C93 drain_left.n0 a_n1756_n1288# 0.26399f
C94 drain_left.n1 a_n1756_n1288# 0.508243f
C95 drain_left.t8 a_n1756_n1288# 0.054698f
C96 drain_left.t5 a_n1756_n1288# 0.054698f
C97 drain_left.n2 a_n1756_n1288# 0.265464f
C98 drain_left.t12 a_n1756_n1288# 0.054698f
C99 drain_left.t11 a_n1756_n1288# 0.054698f
C100 drain_left.n3 a_n1756_n1288# 0.26399f
C101 drain_left.n4 a_n1756_n1288# 0.4936f
C102 drain_left.n5 a_n1756_n1288# 0.629692f
C103 drain_left.t7 a_n1756_n1288# 0.323859f
C104 drain_left.t1 a_n1756_n1288# 0.054698f
C105 drain_left.t3 a_n1756_n1288# 0.054698f
C106 drain_left.n6 a_n1756_n1288# 0.263991f
C107 drain_left.n7 a_n1756_n1288# 0.521174f
C108 drain_left.t6 a_n1756_n1288# 0.054698f
C109 drain_left.t0 a_n1756_n1288# 0.054698f
C110 drain_left.n8 a_n1756_n1288# 0.263991f
C111 drain_left.n9 a_n1756_n1288# 0.257314f
C112 drain_left.t2 a_n1756_n1288# 0.054698f
C113 drain_left.t4 a_n1756_n1288# 0.054698f
C114 drain_left.n10 a_n1756_n1288# 0.263991f
C115 drain_left.n11 a_n1756_n1288# 0.448067f
C116 source.t19 a_n1756_n1288# 0.347201f
C117 source.n0 a_n1756_n1288# 0.661757f
C118 source.t20 a_n1756_n1288# 0.066129f
C119 source.t22 a_n1756_n1288# 0.066129f
C120 source.n1 a_n1756_n1288# 0.278292f
C121 source.n2 a_n1756_n1288# 0.314418f
C122 source.t25 a_n1756_n1288# 0.066129f
C123 source.t24 a_n1756_n1288# 0.066129f
C124 source.n3 a_n1756_n1288# 0.278292f
C125 source.n4 a_n1756_n1288# 0.314418f
C126 source.t18 a_n1756_n1288# 0.066129f
C127 source.t26 a_n1756_n1288# 0.066129f
C128 source.n5 a_n1756_n1288# 0.278292f
C129 source.n6 a_n1756_n1288# 0.331294f
C130 source.t8 a_n1756_n1288# 0.347201f
C131 source.n7 a_n1756_n1288# 0.381417f
C132 source.t3 a_n1756_n1288# 0.066129f
C133 source.t7 a_n1756_n1288# 0.066129f
C134 source.n8 a_n1756_n1288# 0.278292f
C135 source.n9 a_n1756_n1288# 0.314418f
C136 source.t4 a_n1756_n1288# 0.066129f
C137 source.t6 a_n1756_n1288# 0.066129f
C138 source.n10 a_n1756_n1288# 0.278292f
C139 source.n11 a_n1756_n1288# 0.314418f
C140 source.t12 a_n1756_n1288# 0.066129f
C141 source.t2 a_n1756_n1288# 0.066129f
C142 source.n12 a_n1756_n1288# 0.278292f
C143 source.n13 a_n1756_n1288# 0.919296f
C144 source.t14 a_n1756_n1288# 0.066129f
C145 source.t15 a_n1756_n1288# 0.066129f
C146 source.n14 a_n1756_n1288# 0.278291f
C147 source.n15 a_n1756_n1288# 0.919298f
C148 source.t23 a_n1756_n1288# 0.066129f
C149 source.t17 a_n1756_n1288# 0.066129f
C150 source.n16 a_n1756_n1288# 0.278291f
C151 source.n17 a_n1756_n1288# 0.31442f
C152 source.t16 a_n1756_n1288# 0.066129f
C153 source.t27 a_n1756_n1288# 0.066129f
C154 source.n18 a_n1756_n1288# 0.278291f
C155 source.n19 a_n1756_n1288# 0.31442f
C156 source.t21 a_n1756_n1288# 0.3472f
C157 source.n20 a_n1756_n1288# 0.381418f
C158 source.t1 a_n1756_n1288# 0.066129f
C159 source.t9 a_n1756_n1288# 0.066129f
C160 source.n21 a_n1756_n1288# 0.278291f
C161 source.n22 a_n1756_n1288# 0.331296f
C162 source.t0 a_n1756_n1288# 0.066129f
C163 source.t5 a_n1756_n1288# 0.066129f
C164 source.n23 a_n1756_n1288# 0.278291f
C165 source.n24 a_n1756_n1288# 0.31442f
C166 source.t11 a_n1756_n1288# 0.066129f
C167 source.t10 a_n1756_n1288# 0.066129f
C168 source.n25 a_n1756_n1288# 0.278291f
C169 source.n26 a_n1756_n1288# 0.31442f
C170 source.t13 a_n1756_n1288# 0.3472f
C171 source.n27 a_n1756_n1288# 0.513601f
C172 source.n28 a_n1756_n1288# 0.683401f
C173 plus.n0 a_n1756_n1288# 0.035106f
C174 plus.t11 a_n1756_n1288# 0.030991f
C175 plus.t13 a_n1756_n1288# 0.030991f
C176 plus.t7 a_n1756_n1288# 0.030991f
C177 plus.n1 a_n1756_n1288# 0.038702f
C178 plus.n2 a_n1756_n1288# 0.082062f
C179 plus.t10 a_n1756_n1288# 0.030991f
C180 plus.t12 a_n1756_n1288# 0.030991f
C181 plus.t6 a_n1756_n1288# 0.034214f
C182 plus.n3 a_n1756_n1288# 0.040945f
C183 plus.n4 a_n1756_n1288# 0.027056f
C184 plus.n5 a_n1756_n1288# 0.014893f
C185 plus.n6 a_n1756_n1288# 0.027056f
C186 plus.n7 a_n1756_n1288# 0.014893f
C187 plus.n8 a_n1756_n1288# 0.035106f
C188 plus.n9 a_n1756_n1288# 0.035106f
C189 plus.n10 a_n1756_n1288# 0.035106f
C190 plus.n11 a_n1756_n1288# 0.014893f
C191 plus.n12 a_n1756_n1288# 0.027056f
C192 plus.n13 a_n1756_n1288# 0.014893f
C193 plus.n14 a_n1756_n1288# 0.027056f
C194 plus.t9 a_n1756_n1288# 0.034214f
C195 plus.n15 a_n1756_n1288# 0.04089f
C196 plus.n16 a_n1756_n1288# 0.257106f
C197 plus.n17 a_n1756_n1288# 0.035106f
C198 plus.t3 a_n1756_n1288# 0.034214f
C199 plus.t4 a_n1756_n1288# 0.030991f
C200 plus.t0 a_n1756_n1288# 0.030991f
C201 plus.t1 a_n1756_n1288# 0.030991f
C202 plus.n18 a_n1756_n1288# 0.038702f
C203 plus.n19 a_n1756_n1288# 0.082062f
C204 plus.t2 a_n1756_n1288# 0.030991f
C205 plus.t5 a_n1756_n1288# 0.030991f
C206 plus.t8 a_n1756_n1288# 0.034214f
C207 plus.n20 a_n1756_n1288# 0.040945f
C208 plus.n21 a_n1756_n1288# 0.027056f
C209 plus.n22 a_n1756_n1288# 0.014893f
C210 plus.n23 a_n1756_n1288# 0.027056f
C211 plus.n24 a_n1756_n1288# 0.014893f
C212 plus.n25 a_n1756_n1288# 0.035106f
C213 plus.n26 a_n1756_n1288# 0.035106f
C214 plus.n27 a_n1756_n1288# 0.035106f
C215 plus.n28 a_n1756_n1288# 0.014893f
C216 plus.n29 a_n1756_n1288# 0.027056f
C217 plus.n30 a_n1756_n1288# 0.014893f
C218 plus.n31 a_n1756_n1288# 0.027056f
C219 plus.n32 a_n1756_n1288# 0.04089f
C220 plus.n33 a_n1756_n1288# 0.789636f
.ends

