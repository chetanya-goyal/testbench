* NGSPICE file created from diffpair189.ext - technology: sky130A

.subckt diffpair189 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t25 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X1 drain_left.t22 plus.t1 source.t32 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X2 drain_right.t23 minus.t0 source.t0 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X3 source.t4 minus.t1 drain_right.t22 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X4 a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X5 drain_left.t21 plus.t2 source.t26 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X6 drain_left.t20 plus.t3 source.t28 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X7 source.t8 minus.t2 drain_right.t21 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X8 drain_right.t20 minus.t3 source.t12 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X9 drain_left.t19 plus.t4 source.t22 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X10 source.t42 minus.t4 drain_right.t19 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X11 drain_right.t18 minus.t5 source.t9 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X12 drain_right.t17 minus.t6 source.t6 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X13 source.t23 plus.t5 drain_left.t18 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X14 drain_right.t16 minus.t7 source.t43 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X15 source.t20 plus.t6 drain_left.t17 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X16 drain_left.t16 plus.t7 source.t35 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X17 source.t47 minus.t8 drain_right.t15 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X18 drain_left.t15 plus.t8 source.t29 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X19 source.t13 minus.t9 drain_right.t14 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X20 source.t1 minus.t10 drain_right.t13 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X21 drain_left.t14 plus.t9 source.t24 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X22 a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X23 source.t3 minus.t11 drain_right.t12 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X24 drain_left.t13 plus.t10 source.t27 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X25 source.t21 plus.t11 drain_left.t12 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X26 source.t18 plus.t12 drain_left.t11 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X27 source.t19 plus.t13 drain_left.t10 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X28 source.t34 plus.t14 drain_left.t9 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X29 source.t41 plus.t15 drain_left.t8 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X30 source.t36 plus.t16 drain_left.t7 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X31 drain_left.t6 plus.t17 source.t30 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X32 a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X33 source.t31 plus.t18 drain_left.t5 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X34 source.t37 plus.t19 drain_left.t4 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X35 drain_right.t11 minus.t12 source.t5 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X36 source.t39 plus.t20 drain_left.t3 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X37 drain_right.t10 minus.t13 source.t14 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X38 drain_right.t9 minus.t14 source.t45 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X39 source.t40 plus.t21 drain_left.t2 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X40 source.t2 minus.t15 drain_right.t8 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X41 a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X42 drain_left.t1 plus.t22 source.t38 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X43 drain_right.t7 minus.t16 source.t7 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X44 source.t11 minus.t17 drain_right.t6 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X45 drain_right.t5 minus.t18 source.t15 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X46 drain_right.t4 minus.t19 source.t44 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X47 drain_right.t3 minus.t20 source.t10 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X48 source.t16 minus.t21 drain_right.t2 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X49 drain_left.t0 plus.t23 source.t33 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X50 source.t17 minus.t22 drain_right.t1 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X51 source.t46 minus.t23 drain_right.t0 a_n2224_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n6 plus.t5 442.272
R1 plus.n33 plus.t2 442.272
R2 plus.n42 plus.t8 442.272
R3 plus.n68 plus.t15 442.272
R4 plus.n7 plus.t1 414.521
R5 plus.n8 plus.t14 414.521
R6 plus.n14 plus.t0 414.521
R7 plus.n16 plus.t13 414.521
R8 plus.n3 plus.t23 414.521
R9 plus.n21 plus.t12 414.521
R10 plus.n23 plus.t4 414.521
R11 plus.n24 plus.t20 414.521
R12 plus.n30 plus.t3 414.521
R13 plus.n32 plus.t19 414.521
R14 plus.n44 plus.t6 414.521
R15 plus.n43 plus.t10 414.521
R16 plus.n50 plus.t18 414.521
R17 plus.n52 plus.t7 414.521
R18 plus.n39 plus.t11 414.521
R19 plus.n57 plus.t9 414.521
R20 plus.n59 plus.t16 414.521
R21 plus.n38 plus.t22 414.521
R22 plus.n65 plus.t21 414.521
R23 plus.n67 plus.t17 414.521
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus.n17 plus.n3 30.6732
R75 plus.n22 plus.n21 30.6732
R76 plus.n58 plus.n57 30.6732
R77 plus.n53 plus.n39 30.6732
R78 plus plus.n69 27.9498
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 8.66717
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n0 source.t26 69.6943
R119 source.n11 source.t23 69.6943
R120 source.n12 source.t14 69.6943
R121 source.n23 source.t2 69.6943
R122 source.n47 source.t43 69.6942
R123 source.n36 source.t46 69.6942
R124 source.n35 source.t29 69.6942
R125 source.n24 source.t41 69.6942
R126 source.n2 source.n1 63.0943
R127 source.n4 source.n3 63.0943
R128 source.n6 source.n5 63.0943
R129 source.n8 source.n7 63.0943
R130 source.n10 source.n9 63.0943
R131 source.n14 source.n13 63.0943
R132 source.n16 source.n15 63.0943
R133 source.n18 source.n17 63.0943
R134 source.n20 source.n19 63.0943
R135 source.n22 source.n21 63.0943
R136 source.n46 source.n45 63.0942
R137 source.n44 source.n43 63.0942
R138 source.n42 source.n41 63.0942
R139 source.n40 source.n39 63.0942
R140 source.n38 source.n37 63.0942
R141 source.n34 source.n33 63.0942
R142 source.n32 source.n31 63.0942
R143 source.n30 source.n29 63.0942
R144 source.n28 source.n27 63.0942
R145 source.n26 source.n25 63.0942
R146 source.n24 source.n23 14.9695
R147 source.n48 source.n0 9.45661
R148 source.n45 source.t6 6.6005
R149 source.n45 source.t47 6.6005
R150 source.n43 source.t0 6.6005
R151 source.n43 source.t17 6.6005
R152 source.n41 source.t12 6.6005
R153 source.n41 source.t4 6.6005
R154 source.n39 source.t7 6.6005
R155 source.n39 source.t16 6.6005
R156 source.n37 source.t45 6.6005
R157 source.n37 source.t11 6.6005
R158 source.n33 source.t27 6.6005
R159 source.n33 source.t20 6.6005
R160 source.n31 source.t35 6.6005
R161 source.n31 source.t31 6.6005
R162 source.n29 source.t24 6.6005
R163 source.n29 source.t21 6.6005
R164 source.n27 source.t38 6.6005
R165 source.n27 source.t36 6.6005
R166 source.n25 source.t30 6.6005
R167 source.n25 source.t40 6.6005
R168 source.n1 source.t28 6.6005
R169 source.n1 source.t37 6.6005
R170 source.n3 source.t22 6.6005
R171 source.n3 source.t39 6.6005
R172 source.n5 source.t33 6.6005
R173 source.n5 source.t18 6.6005
R174 source.n7 source.t25 6.6005
R175 source.n7 source.t19 6.6005
R176 source.n9 source.t32 6.6005
R177 source.n9 source.t34 6.6005
R178 source.n13 source.t5 6.6005
R179 source.n13 source.t42 6.6005
R180 source.n15 source.t15 6.6005
R181 source.n15 source.t8 6.6005
R182 source.n17 source.t44 6.6005
R183 source.n17 source.t1 6.6005
R184 source.n19 source.t10 6.6005
R185 source.n19 source.t13 6.6005
R186 source.n21 source.t9 6.6005
R187 source.n21 source.t3 6.6005
R188 source.n48 source.n47 5.51343
R189 source.n23 source.n22 0.5005
R190 source.n22 source.n20 0.5005
R191 source.n20 source.n18 0.5005
R192 source.n18 source.n16 0.5005
R193 source.n16 source.n14 0.5005
R194 source.n14 source.n12 0.5005
R195 source.n11 source.n10 0.5005
R196 source.n10 source.n8 0.5005
R197 source.n8 source.n6 0.5005
R198 source.n6 source.n4 0.5005
R199 source.n4 source.n2 0.5005
R200 source.n2 source.n0 0.5005
R201 source.n26 source.n24 0.5005
R202 source.n28 source.n26 0.5005
R203 source.n30 source.n28 0.5005
R204 source.n32 source.n30 0.5005
R205 source.n34 source.n32 0.5005
R206 source.n35 source.n34 0.5005
R207 source.n38 source.n36 0.5005
R208 source.n40 source.n38 0.5005
R209 source.n42 source.n40 0.5005
R210 source.n44 source.n42 0.5005
R211 source.n46 source.n44 0.5005
R212 source.n47 source.n46 0.5005
R213 source.n12 source.n11 0.470328
R214 source.n36 source.n35 0.470328
R215 source source.n48 0.188
R216 drain_left.n13 drain_left.n11 80.2731
R217 drain_left.n7 drain_left.n5 80.273
R218 drain_left.n2 drain_left.n0 80.273
R219 drain_left.n21 drain_left.n20 79.7731
R220 drain_left.n19 drain_left.n18 79.7731
R221 drain_left.n17 drain_left.n16 79.7731
R222 drain_left.n15 drain_left.n14 79.7731
R223 drain_left.n13 drain_left.n12 79.7731
R224 drain_left.n7 drain_left.n6 79.773
R225 drain_left.n9 drain_left.n8 79.773
R226 drain_left.n4 drain_left.n3 79.773
R227 drain_left.n2 drain_left.n1 79.773
R228 drain_left drain_left.n10 25.2989
R229 drain_left.n5 drain_left.t17 6.6005
R230 drain_left.n5 drain_left.t15 6.6005
R231 drain_left.n6 drain_left.t5 6.6005
R232 drain_left.n6 drain_left.t13 6.6005
R233 drain_left.n8 drain_left.t12 6.6005
R234 drain_left.n8 drain_left.t16 6.6005
R235 drain_left.n3 drain_left.t7 6.6005
R236 drain_left.n3 drain_left.t14 6.6005
R237 drain_left.n1 drain_left.t2 6.6005
R238 drain_left.n1 drain_left.t1 6.6005
R239 drain_left.n0 drain_left.t8 6.6005
R240 drain_left.n0 drain_left.t6 6.6005
R241 drain_left.n20 drain_left.t4 6.6005
R242 drain_left.n20 drain_left.t21 6.6005
R243 drain_left.n18 drain_left.t3 6.6005
R244 drain_left.n18 drain_left.t20 6.6005
R245 drain_left.n16 drain_left.t11 6.6005
R246 drain_left.n16 drain_left.t19 6.6005
R247 drain_left.n14 drain_left.t10 6.6005
R248 drain_left.n14 drain_left.t0 6.6005
R249 drain_left.n12 drain_left.t9 6.6005
R250 drain_left.n12 drain_left.t23 6.6005
R251 drain_left.n11 drain_left.t18 6.6005
R252 drain_left.n11 drain_left.t22 6.6005
R253 drain_left drain_left.n21 6.15322
R254 drain_left.n9 drain_left.n7 0.5005
R255 drain_left.n4 drain_left.n2 0.5005
R256 drain_left.n15 drain_left.n13 0.5005
R257 drain_left.n17 drain_left.n15 0.5005
R258 drain_left.n19 drain_left.n17 0.5005
R259 drain_left.n21 drain_left.n19 0.5005
R260 drain_left.n10 drain_left.n9 0.195154
R261 drain_left.n10 drain_left.n4 0.195154
R262 minus.n33 minus.t15 442.272
R263 minus.n7 minus.t13 442.272
R264 minus.n68 minus.t7 442.272
R265 minus.n41 minus.t23 442.272
R266 minus.n32 minus.t5 414.521
R267 minus.n30 minus.t11 414.521
R268 minus.n3 minus.t20 414.521
R269 minus.n24 minus.t9 414.521
R270 minus.n22 minus.t19 414.521
R271 minus.n4 minus.t10 414.521
R272 minus.n17 minus.t18 414.521
R273 minus.n15 minus.t2 414.521
R274 minus.n8 minus.t12 414.521
R275 minus.n9 minus.t4 414.521
R276 minus.n67 minus.t8 414.521
R277 minus.n65 minus.t6 414.521
R278 minus.n59 minus.t22 414.521
R279 minus.n58 minus.t0 414.521
R280 minus.n56 minus.t1 414.521
R281 minus.n38 minus.t3 414.521
R282 minus.n51 minus.t21 414.521
R283 minus.n49 minus.t16 414.521
R284 minus.n43 minus.t17 414.521
R285 minus.n42 minus.t14 414.521
R286 minus.n11 minus.n7 161.489
R287 minus.n45 minus.n41 161.489
R288 minus.n34 minus.n33 161.3
R289 minus.n31 minus.n0 161.3
R290 minus.n29 minus.n28 161.3
R291 minus.n27 minus.n1 161.3
R292 minus.n26 minus.n25 161.3
R293 minus.n23 minus.n2 161.3
R294 minus.n21 minus.n20 161.3
R295 minus.n19 minus.n18 161.3
R296 minus.n16 minus.n5 161.3
R297 minus.n14 minus.n13 161.3
R298 minus.n12 minus.n6 161.3
R299 minus.n11 minus.n10 161.3
R300 minus.n69 minus.n68 161.3
R301 minus.n66 minus.n35 161.3
R302 minus.n64 minus.n63 161.3
R303 minus.n62 minus.n36 161.3
R304 minus.n61 minus.n60 161.3
R305 minus.n57 minus.n37 161.3
R306 minus.n55 minus.n54 161.3
R307 minus.n53 minus.n52 161.3
R308 minus.n50 minus.n39 161.3
R309 minus.n48 minus.n47 161.3
R310 minus.n46 minus.n40 161.3
R311 minus.n45 minus.n44 161.3
R312 minus.n29 minus.n1 73.0308
R313 minus.n14 minus.n6 73.0308
R314 minus.n48 minus.n40 73.0308
R315 minus.n64 minus.n36 73.0308
R316 minus.n31 minus.n30 68.649
R317 minus.n10 minus.n8 68.649
R318 minus.n44 minus.n43 68.649
R319 minus.n66 minus.n65 68.649
R320 minus.n25 minus.n3 65.7278
R321 minus.n16 minus.n15 65.7278
R322 minus.n50 minus.n49 65.7278
R323 minus.n60 minus.n59 65.7278
R324 minus.n33 minus.n32 56.9641
R325 minus.n9 minus.n7 56.9641
R326 minus.n42 minus.n41 56.9641
R327 minus.n68 minus.n67 56.9641
R328 minus.n24 minus.n23 54.0429
R329 minus.n18 minus.n17 54.0429
R330 minus.n52 minus.n51 54.0429
R331 minus.n58 minus.n57 54.0429
R332 minus.n22 minus.n21 42.3581
R333 minus.n21 minus.n4 42.3581
R334 minus.n55 minus.n38 42.3581
R335 minus.n56 minus.n55 42.3581
R336 minus.n23 minus.n22 30.6732
R337 minus.n18 minus.n4 30.6732
R338 minus.n52 minus.n38 30.6732
R339 minus.n57 minus.n56 30.6732
R340 minus.n70 minus.n34 30.6596
R341 minus.n25 minus.n24 18.9884
R342 minus.n17 minus.n16 18.9884
R343 minus.n51 minus.n50 18.9884
R344 minus.n60 minus.n58 18.9884
R345 minus.n32 minus.n31 16.0672
R346 minus.n10 minus.n9 16.0672
R347 minus.n44 minus.n42 16.0672
R348 minus.n67 minus.n66 16.0672
R349 minus.n3 minus.n1 7.30353
R350 minus.n15 minus.n14 7.30353
R351 minus.n49 minus.n48 7.30353
R352 minus.n59 minus.n36 7.30353
R353 minus.n70 minus.n69 6.43232
R354 minus.n30 minus.n29 4.38232
R355 minus.n8 minus.n6 4.38232
R356 minus.n43 minus.n40 4.38232
R357 minus.n65 minus.n64 4.38232
R358 minus.n34 minus.n0 0.189894
R359 minus.n28 minus.n0 0.189894
R360 minus.n28 minus.n27 0.189894
R361 minus.n27 minus.n26 0.189894
R362 minus.n26 minus.n2 0.189894
R363 minus.n20 minus.n2 0.189894
R364 minus.n20 minus.n19 0.189894
R365 minus.n19 minus.n5 0.189894
R366 minus.n13 minus.n5 0.189894
R367 minus.n13 minus.n12 0.189894
R368 minus.n12 minus.n11 0.189894
R369 minus.n46 minus.n45 0.189894
R370 minus.n47 minus.n46 0.189894
R371 minus.n47 minus.n39 0.189894
R372 minus.n53 minus.n39 0.189894
R373 minus.n54 minus.n53 0.189894
R374 minus.n54 minus.n37 0.189894
R375 minus.n61 minus.n37 0.189894
R376 minus.n62 minus.n61 0.189894
R377 minus.n63 minus.n62 0.189894
R378 minus.n63 minus.n35 0.189894
R379 minus.n69 minus.n35 0.189894
R380 minus minus.n70 0.188
R381 drain_right.n13 drain_right.n11 80.2731
R382 drain_right.n7 drain_right.n5 80.273
R383 drain_right.n2 drain_right.n0 80.273
R384 drain_right.n13 drain_right.n12 79.7731
R385 drain_right.n15 drain_right.n14 79.7731
R386 drain_right.n17 drain_right.n16 79.7731
R387 drain_right.n19 drain_right.n18 79.7731
R388 drain_right.n21 drain_right.n20 79.7731
R389 drain_right.n7 drain_right.n6 79.773
R390 drain_right.n9 drain_right.n8 79.773
R391 drain_right.n4 drain_right.n3 79.773
R392 drain_right.n2 drain_right.n1 79.773
R393 drain_right drain_right.n10 24.7457
R394 drain_right.n5 drain_right.t15 6.6005
R395 drain_right.n5 drain_right.t16 6.6005
R396 drain_right.n6 drain_right.t1 6.6005
R397 drain_right.n6 drain_right.t17 6.6005
R398 drain_right.n8 drain_right.t22 6.6005
R399 drain_right.n8 drain_right.t23 6.6005
R400 drain_right.n3 drain_right.t2 6.6005
R401 drain_right.n3 drain_right.t20 6.6005
R402 drain_right.n1 drain_right.t6 6.6005
R403 drain_right.n1 drain_right.t7 6.6005
R404 drain_right.n0 drain_right.t0 6.6005
R405 drain_right.n0 drain_right.t9 6.6005
R406 drain_right.n11 drain_right.t19 6.6005
R407 drain_right.n11 drain_right.t10 6.6005
R408 drain_right.n12 drain_right.t21 6.6005
R409 drain_right.n12 drain_right.t11 6.6005
R410 drain_right.n14 drain_right.t13 6.6005
R411 drain_right.n14 drain_right.t5 6.6005
R412 drain_right.n16 drain_right.t14 6.6005
R413 drain_right.n16 drain_right.t4 6.6005
R414 drain_right.n18 drain_right.t12 6.6005
R415 drain_right.n18 drain_right.t3 6.6005
R416 drain_right.n20 drain_right.t8 6.6005
R417 drain_right.n20 drain_right.t18 6.6005
R418 drain_right drain_right.n21 6.15322
R419 drain_right.n9 drain_right.n7 0.5005
R420 drain_right.n4 drain_right.n2 0.5005
R421 drain_right.n21 drain_right.n19 0.5005
R422 drain_right.n19 drain_right.n17 0.5005
R423 drain_right.n17 drain_right.n15 0.5005
R424 drain_right.n15 drain_right.n13 0.5005
R425 drain_right.n10 drain_right.n9 0.195154
R426 drain_right.n10 drain_right.n4 0.195154
C0 drain_right plus 0.379713f
C1 drain_right source 14.934099f
C2 drain_left plus 2.55195f
C3 drain_left source 14.933701f
C4 drain_right minus 2.3333f
C5 source plus 2.5621f
C6 drain_left minus 0.177436f
C7 minus plus 4.27439f
C8 drain_right drain_left 1.19771f
C9 source minus 2.54811f
C10 drain_right a_n2224_n1488# 5.207651f
C11 drain_left a_n2224_n1488# 5.5636f
C12 source a_n2224_n1488# 3.872678f
C13 minus a_n2224_n1488# 8.005445f
C14 plus a_n2224_n1488# 9.493441f
C15 drain_right.t0 a_n2224_n1488# 0.081718f
C16 drain_right.t9 a_n2224_n1488# 0.081718f
C17 drain_right.n0 a_n2224_n1488# 0.591841f
C18 drain_right.t6 a_n2224_n1488# 0.081718f
C19 drain_right.t7 a_n2224_n1488# 0.081718f
C20 drain_right.n1 a_n2224_n1488# 0.589344f
C21 drain_right.n2 a_n2224_n1488# 0.785386f
C22 drain_right.t2 a_n2224_n1488# 0.081718f
C23 drain_right.t20 a_n2224_n1488# 0.081718f
C24 drain_right.n3 a_n2224_n1488# 0.589344f
C25 drain_right.n4 a_n2224_n1488# 0.35719f
C26 drain_right.t15 a_n2224_n1488# 0.081718f
C27 drain_right.t16 a_n2224_n1488# 0.081718f
C28 drain_right.n5 a_n2224_n1488# 0.591841f
C29 drain_right.t1 a_n2224_n1488# 0.081718f
C30 drain_right.t17 a_n2224_n1488# 0.081718f
C31 drain_right.n6 a_n2224_n1488# 0.589344f
C32 drain_right.n7 a_n2224_n1488# 0.785386f
C33 drain_right.t22 a_n2224_n1488# 0.081718f
C34 drain_right.t23 a_n2224_n1488# 0.081718f
C35 drain_right.n8 a_n2224_n1488# 0.589344f
C36 drain_right.n9 a_n2224_n1488# 0.35719f
C37 drain_right.n10 a_n2224_n1488# 1.10049f
C38 drain_right.t19 a_n2224_n1488# 0.081718f
C39 drain_right.t10 a_n2224_n1488# 0.081718f
C40 drain_right.n11 a_n2224_n1488# 0.591844f
C41 drain_right.t21 a_n2224_n1488# 0.081718f
C42 drain_right.t11 a_n2224_n1488# 0.081718f
C43 drain_right.n12 a_n2224_n1488# 0.589347f
C44 drain_right.n13 a_n2224_n1488# 0.785381f
C45 drain_right.t13 a_n2224_n1488# 0.081718f
C46 drain_right.t5 a_n2224_n1488# 0.081718f
C47 drain_right.n14 a_n2224_n1488# 0.589347f
C48 drain_right.n15 a_n2224_n1488# 0.386997f
C49 drain_right.t14 a_n2224_n1488# 0.081718f
C50 drain_right.t4 a_n2224_n1488# 0.081718f
C51 drain_right.n16 a_n2224_n1488# 0.589347f
C52 drain_right.n17 a_n2224_n1488# 0.386997f
C53 drain_right.t12 a_n2224_n1488# 0.081718f
C54 drain_right.t3 a_n2224_n1488# 0.081718f
C55 drain_right.n18 a_n2224_n1488# 0.589347f
C56 drain_right.n19 a_n2224_n1488# 0.386997f
C57 drain_right.t8 a_n2224_n1488# 0.081718f
C58 drain_right.t18 a_n2224_n1488# 0.081718f
C59 drain_right.n20 a_n2224_n1488# 0.589347f
C60 drain_right.n21 a_n2224_n1488# 0.671525f
C61 minus.n0 a_n2224_n1488# 0.049302f
C62 minus.t15 a_n2224_n1488# 0.111025f
C63 minus.t5 a_n2224_n1488# 0.10708f
C64 minus.t11 a_n2224_n1488# 0.10708f
C65 minus.n1 a_n2224_n1488# 0.017875f
C66 minus.n2 a_n2224_n1488# 0.049302f
C67 minus.t20 a_n2224_n1488# 0.10708f
C68 minus.n3 a_n2224_n1488# 0.064708f
C69 minus.t9 a_n2224_n1488# 0.10708f
C70 minus.t19 a_n2224_n1488# 0.10708f
C71 minus.t10 a_n2224_n1488# 0.10708f
C72 minus.n4 a_n2224_n1488# 0.064708f
C73 minus.n5 a_n2224_n1488# 0.049302f
C74 minus.t18 a_n2224_n1488# 0.10708f
C75 minus.t2 a_n2224_n1488# 0.10708f
C76 minus.n6 a_n2224_n1488# 0.017267f
C77 minus.t13 a_n2224_n1488# 0.111025f
C78 minus.n7 a_n2224_n1488# 0.077788f
C79 minus.t12 a_n2224_n1488# 0.10708f
C80 minus.n8 a_n2224_n1488# 0.064708f
C81 minus.t4 a_n2224_n1488# 0.10708f
C82 minus.n9 a_n2224_n1488# 0.064708f
C83 minus.n10 a_n2224_n1488# 0.018787f
C84 minus.n11 a_n2224_n1488# 0.102493f
C85 minus.n12 a_n2224_n1488# 0.049302f
C86 minus.n13 a_n2224_n1488# 0.049302f
C87 minus.n14 a_n2224_n1488# 0.017875f
C88 minus.n15 a_n2224_n1488# 0.064708f
C89 minus.n16 a_n2224_n1488# 0.018787f
C90 minus.n17 a_n2224_n1488# 0.064708f
C91 minus.n18 a_n2224_n1488# 0.018787f
C92 minus.n19 a_n2224_n1488# 0.049302f
C93 minus.n20 a_n2224_n1488# 0.049302f
C94 minus.n21 a_n2224_n1488# 0.018787f
C95 minus.n22 a_n2224_n1488# 0.064708f
C96 minus.n23 a_n2224_n1488# 0.018787f
C97 minus.n24 a_n2224_n1488# 0.064708f
C98 minus.n25 a_n2224_n1488# 0.018787f
C99 minus.n26 a_n2224_n1488# 0.049302f
C100 minus.n27 a_n2224_n1488# 0.049302f
C101 minus.n28 a_n2224_n1488# 0.049302f
C102 minus.n29 a_n2224_n1488# 0.017267f
C103 minus.n30 a_n2224_n1488# 0.064708f
C104 minus.n31 a_n2224_n1488# 0.018787f
C105 minus.n32 a_n2224_n1488# 0.064708f
C106 minus.n33 a_n2224_n1488# 0.077725f
C107 minus.n34 a_n2224_n1488# 1.32777f
C108 minus.n35 a_n2224_n1488# 0.049302f
C109 minus.t8 a_n2224_n1488# 0.10708f
C110 minus.t6 a_n2224_n1488# 0.10708f
C111 minus.n36 a_n2224_n1488# 0.017875f
C112 minus.n37 a_n2224_n1488# 0.049302f
C113 minus.t0 a_n2224_n1488# 0.10708f
C114 minus.t1 a_n2224_n1488# 0.10708f
C115 minus.t3 a_n2224_n1488# 0.10708f
C116 minus.n38 a_n2224_n1488# 0.064708f
C117 minus.n39 a_n2224_n1488# 0.049302f
C118 minus.t21 a_n2224_n1488# 0.10708f
C119 minus.t16 a_n2224_n1488# 0.10708f
C120 minus.n40 a_n2224_n1488# 0.017267f
C121 minus.t23 a_n2224_n1488# 0.111025f
C122 minus.n41 a_n2224_n1488# 0.077788f
C123 minus.t14 a_n2224_n1488# 0.10708f
C124 minus.n42 a_n2224_n1488# 0.064708f
C125 minus.t17 a_n2224_n1488# 0.10708f
C126 minus.n43 a_n2224_n1488# 0.064708f
C127 minus.n44 a_n2224_n1488# 0.018787f
C128 minus.n45 a_n2224_n1488# 0.102493f
C129 minus.n46 a_n2224_n1488# 0.049302f
C130 minus.n47 a_n2224_n1488# 0.049302f
C131 minus.n48 a_n2224_n1488# 0.017875f
C132 minus.n49 a_n2224_n1488# 0.064708f
C133 minus.n50 a_n2224_n1488# 0.018787f
C134 minus.n51 a_n2224_n1488# 0.064708f
C135 minus.n52 a_n2224_n1488# 0.018787f
C136 minus.n53 a_n2224_n1488# 0.049302f
C137 minus.n54 a_n2224_n1488# 0.049302f
C138 minus.n55 a_n2224_n1488# 0.018787f
C139 minus.n56 a_n2224_n1488# 0.064708f
C140 minus.n57 a_n2224_n1488# 0.018787f
C141 minus.n58 a_n2224_n1488# 0.064708f
C142 minus.t22 a_n2224_n1488# 0.10708f
C143 minus.n59 a_n2224_n1488# 0.064708f
C144 minus.n60 a_n2224_n1488# 0.018787f
C145 minus.n61 a_n2224_n1488# 0.049302f
C146 minus.n62 a_n2224_n1488# 0.049302f
C147 minus.n63 a_n2224_n1488# 0.049302f
C148 minus.n64 a_n2224_n1488# 0.017267f
C149 minus.n65 a_n2224_n1488# 0.064708f
C150 minus.n66 a_n2224_n1488# 0.018787f
C151 minus.n67 a_n2224_n1488# 0.064708f
C152 minus.t7 a_n2224_n1488# 0.111025f
C153 minus.n68 a_n2224_n1488# 0.077725f
C154 minus.n69 a_n2224_n1488# 0.314437f
C155 minus.n70 a_n2224_n1488# 1.63993f
C156 drain_left.t8 a_n2224_n1488# 0.082497f
C157 drain_left.t6 a_n2224_n1488# 0.082497f
C158 drain_left.n0 a_n2224_n1488# 0.59748f
C159 drain_left.t2 a_n2224_n1488# 0.082497f
C160 drain_left.t1 a_n2224_n1488# 0.082497f
C161 drain_left.n1 a_n2224_n1488# 0.594959f
C162 drain_left.n2 a_n2224_n1488# 0.792869f
C163 drain_left.t7 a_n2224_n1488# 0.082497f
C164 drain_left.t14 a_n2224_n1488# 0.082497f
C165 drain_left.n3 a_n2224_n1488# 0.594959f
C166 drain_left.n4 a_n2224_n1488# 0.360593f
C167 drain_left.t17 a_n2224_n1488# 0.082497f
C168 drain_left.t15 a_n2224_n1488# 0.082497f
C169 drain_left.n5 a_n2224_n1488# 0.59748f
C170 drain_left.t5 a_n2224_n1488# 0.082497f
C171 drain_left.t13 a_n2224_n1488# 0.082497f
C172 drain_left.n6 a_n2224_n1488# 0.594959f
C173 drain_left.n7 a_n2224_n1488# 0.792869f
C174 drain_left.t12 a_n2224_n1488# 0.082497f
C175 drain_left.t16 a_n2224_n1488# 0.082497f
C176 drain_left.n8 a_n2224_n1488# 0.594959f
C177 drain_left.n9 a_n2224_n1488# 0.360593f
C178 drain_left.n10 a_n2224_n1488# 1.1796f
C179 drain_left.t18 a_n2224_n1488# 0.082497f
C180 drain_left.t22 a_n2224_n1488# 0.082497f
C181 drain_left.n11 a_n2224_n1488# 0.597483f
C182 drain_left.t9 a_n2224_n1488# 0.082497f
C183 drain_left.t23 a_n2224_n1488# 0.082497f
C184 drain_left.n12 a_n2224_n1488# 0.594962f
C185 drain_left.n13 a_n2224_n1488# 0.792863f
C186 drain_left.t10 a_n2224_n1488# 0.082497f
C187 drain_left.t0 a_n2224_n1488# 0.082497f
C188 drain_left.n14 a_n2224_n1488# 0.594962f
C189 drain_left.n15 a_n2224_n1488# 0.390684f
C190 drain_left.t11 a_n2224_n1488# 0.082497f
C191 drain_left.t19 a_n2224_n1488# 0.082497f
C192 drain_left.n16 a_n2224_n1488# 0.594962f
C193 drain_left.n17 a_n2224_n1488# 0.390684f
C194 drain_left.t3 a_n2224_n1488# 0.082497f
C195 drain_left.t20 a_n2224_n1488# 0.082497f
C196 drain_left.n18 a_n2224_n1488# 0.594962f
C197 drain_left.n19 a_n2224_n1488# 0.390684f
C198 drain_left.t4 a_n2224_n1488# 0.082497f
C199 drain_left.t21 a_n2224_n1488# 0.082497f
C200 drain_left.n20 a_n2224_n1488# 0.594962f
C201 drain_left.n21 a_n2224_n1488# 0.677923f
C202 source.t26 a_n2224_n1488# 0.689367f
C203 source.n0 a_n2224_n1488# 0.931959f
C204 source.t28 a_n2224_n1488# 0.083018f
C205 source.t37 a_n2224_n1488# 0.083018f
C206 source.n1 a_n2224_n1488# 0.526382f
C207 source.n2 a_n2224_n1488# 0.417894f
C208 source.t22 a_n2224_n1488# 0.083018f
C209 source.t39 a_n2224_n1488# 0.083018f
C210 source.n3 a_n2224_n1488# 0.526382f
C211 source.n4 a_n2224_n1488# 0.417894f
C212 source.t33 a_n2224_n1488# 0.083018f
C213 source.t18 a_n2224_n1488# 0.083018f
C214 source.n5 a_n2224_n1488# 0.526382f
C215 source.n6 a_n2224_n1488# 0.417894f
C216 source.t25 a_n2224_n1488# 0.083018f
C217 source.t19 a_n2224_n1488# 0.083018f
C218 source.n7 a_n2224_n1488# 0.526382f
C219 source.n8 a_n2224_n1488# 0.417894f
C220 source.t32 a_n2224_n1488# 0.083018f
C221 source.t34 a_n2224_n1488# 0.083018f
C222 source.n9 a_n2224_n1488# 0.526382f
C223 source.n10 a_n2224_n1488# 0.417894f
C224 source.t23 a_n2224_n1488# 0.689367f
C225 source.n11 a_n2224_n1488# 0.477917f
C226 source.t14 a_n2224_n1488# 0.689367f
C227 source.n12 a_n2224_n1488# 0.477917f
C228 source.t5 a_n2224_n1488# 0.083018f
C229 source.t42 a_n2224_n1488# 0.083018f
C230 source.n13 a_n2224_n1488# 0.526382f
C231 source.n14 a_n2224_n1488# 0.417894f
C232 source.t15 a_n2224_n1488# 0.083018f
C233 source.t8 a_n2224_n1488# 0.083018f
C234 source.n15 a_n2224_n1488# 0.526382f
C235 source.n16 a_n2224_n1488# 0.417894f
C236 source.t44 a_n2224_n1488# 0.083018f
C237 source.t1 a_n2224_n1488# 0.083018f
C238 source.n17 a_n2224_n1488# 0.526382f
C239 source.n18 a_n2224_n1488# 0.417894f
C240 source.t10 a_n2224_n1488# 0.083018f
C241 source.t13 a_n2224_n1488# 0.083018f
C242 source.n19 a_n2224_n1488# 0.526382f
C243 source.n20 a_n2224_n1488# 0.417894f
C244 source.t9 a_n2224_n1488# 0.083018f
C245 source.t3 a_n2224_n1488# 0.083018f
C246 source.n21 a_n2224_n1488# 0.526382f
C247 source.n22 a_n2224_n1488# 0.417894f
C248 source.t2 a_n2224_n1488# 0.689367f
C249 source.n23 a_n2224_n1488# 1.29582f
C250 source.t41 a_n2224_n1488# 0.689364f
C251 source.n24 a_n2224_n1488# 1.29583f
C252 source.t30 a_n2224_n1488# 0.083018f
C253 source.t40 a_n2224_n1488# 0.083018f
C254 source.n25 a_n2224_n1488# 0.526378f
C255 source.n26 a_n2224_n1488# 0.417898f
C256 source.t38 a_n2224_n1488# 0.083018f
C257 source.t36 a_n2224_n1488# 0.083018f
C258 source.n27 a_n2224_n1488# 0.526378f
C259 source.n28 a_n2224_n1488# 0.417898f
C260 source.t24 a_n2224_n1488# 0.083018f
C261 source.t21 a_n2224_n1488# 0.083018f
C262 source.n29 a_n2224_n1488# 0.526378f
C263 source.n30 a_n2224_n1488# 0.417898f
C264 source.t35 a_n2224_n1488# 0.083018f
C265 source.t31 a_n2224_n1488# 0.083018f
C266 source.n31 a_n2224_n1488# 0.526378f
C267 source.n32 a_n2224_n1488# 0.417898f
C268 source.t27 a_n2224_n1488# 0.083018f
C269 source.t20 a_n2224_n1488# 0.083018f
C270 source.n33 a_n2224_n1488# 0.526378f
C271 source.n34 a_n2224_n1488# 0.417898f
C272 source.t29 a_n2224_n1488# 0.689364f
C273 source.n35 a_n2224_n1488# 0.477921f
C274 source.t46 a_n2224_n1488# 0.689364f
C275 source.n36 a_n2224_n1488# 0.477921f
C276 source.t45 a_n2224_n1488# 0.083018f
C277 source.t11 a_n2224_n1488# 0.083018f
C278 source.n37 a_n2224_n1488# 0.526378f
C279 source.n38 a_n2224_n1488# 0.417898f
C280 source.t7 a_n2224_n1488# 0.083018f
C281 source.t16 a_n2224_n1488# 0.083018f
C282 source.n39 a_n2224_n1488# 0.526378f
C283 source.n40 a_n2224_n1488# 0.417898f
C284 source.t12 a_n2224_n1488# 0.083018f
C285 source.t4 a_n2224_n1488# 0.083018f
C286 source.n41 a_n2224_n1488# 0.526378f
C287 source.n42 a_n2224_n1488# 0.417898f
C288 source.t0 a_n2224_n1488# 0.083018f
C289 source.t17 a_n2224_n1488# 0.083018f
C290 source.n43 a_n2224_n1488# 0.526378f
C291 source.n44 a_n2224_n1488# 0.417898f
C292 source.t6 a_n2224_n1488# 0.083018f
C293 source.t47 a_n2224_n1488# 0.083018f
C294 source.n45 a_n2224_n1488# 0.526378f
C295 source.n46 a_n2224_n1488# 0.417898f
C296 source.t43 a_n2224_n1488# 0.689364f
C297 source.n47 a_n2224_n1488# 0.671707f
C298 source.n48 a_n2224_n1488# 1.01289f
C299 plus.n0 a_n2224_n1488# 0.052039f
C300 plus.t19 a_n2224_n1488# 0.113025f
C301 plus.t3 a_n2224_n1488# 0.113025f
C302 plus.n1 a_n2224_n1488# 0.018867f
C303 plus.n2 a_n2224_n1488# 0.052039f
C304 plus.t4 a_n2224_n1488# 0.113025f
C305 plus.t12 a_n2224_n1488# 0.113025f
C306 plus.t23 a_n2224_n1488# 0.113025f
C307 plus.n3 a_n2224_n1488# 0.068301f
C308 plus.n4 a_n2224_n1488# 0.052039f
C309 plus.t13 a_n2224_n1488# 0.113025f
C310 plus.t0 a_n2224_n1488# 0.113025f
C311 plus.n5 a_n2224_n1488# 0.018226f
C312 plus.t5 a_n2224_n1488# 0.11719f
C313 plus.n6 a_n2224_n1488# 0.082107f
C314 plus.t1 a_n2224_n1488# 0.113025f
C315 plus.n7 a_n2224_n1488# 0.068301f
C316 plus.t14 a_n2224_n1488# 0.113025f
C317 plus.n8 a_n2224_n1488# 0.068301f
C318 plus.n9 a_n2224_n1488# 0.01983f
C319 plus.n10 a_n2224_n1488# 0.108183f
C320 plus.n11 a_n2224_n1488# 0.052039f
C321 plus.n12 a_n2224_n1488# 0.052039f
C322 plus.n13 a_n2224_n1488# 0.018867f
C323 plus.n14 a_n2224_n1488# 0.068301f
C324 plus.n15 a_n2224_n1488# 0.01983f
C325 plus.n16 a_n2224_n1488# 0.068301f
C326 plus.n17 a_n2224_n1488# 0.01983f
C327 plus.n18 a_n2224_n1488# 0.052039f
C328 plus.n19 a_n2224_n1488# 0.052039f
C329 plus.n20 a_n2224_n1488# 0.01983f
C330 plus.n21 a_n2224_n1488# 0.068301f
C331 plus.n22 a_n2224_n1488# 0.01983f
C332 plus.n23 a_n2224_n1488# 0.068301f
C333 plus.t20 a_n2224_n1488# 0.113025f
C334 plus.n24 a_n2224_n1488# 0.068301f
C335 plus.n25 a_n2224_n1488# 0.01983f
C336 plus.n26 a_n2224_n1488# 0.052039f
C337 plus.n27 a_n2224_n1488# 0.052039f
C338 plus.n28 a_n2224_n1488# 0.052039f
C339 plus.n29 a_n2224_n1488# 0.018226f
C340 plus.n30 a_n2224_n1488# 0.068301f
C341 plus.n31 a_n2224_n1488# 0.01983f
C342 plus.n32 a_n2224_n1488# 0.068301f
C343 plus.t2 a_n2224_n1488# 0.11719f
C344 plus.n33 a_n2224_n1488# 0.082041f
C345 plus.n34 a_n2224_n1488# 0.379971f
C346 plus.n35 a_n2224_n1488# 0.052039f
C347 plus.t15 a_n2224_n1488# 0.11719f
C348 plus.t17 a_n2224_n1488# 0.113025f
C349 plus.t21 a_n2224_n1488# 0.113025f
C350 plus.n36 a_n2224_n1488# 0.018867f
C351 plus.n37 a_n2224_n1488# 0.052039f
C352 plus.t22 a_n2224_n1488# 0.113025f
C353 plus.n38 a_n2224_n1488# 0.068301f
C354 plus.t16 a_n2224_n1488# 0.113025f
C355 plus.t9 a_n2224_n1488# 0.113025f
C356 plus.t11 a_n2224_n1488# 0.113025f
C357 plus.n39 a_n2224_n1488# 0.068301f
C358 plus.n40 a_n2224_n1488# 0.052039f
C359 plus.t7 a_n2224_n1488# 0.113025f
C360 plus.t18 a_n2224_n1488# 0.113025f
C361 plus.n41 a_n2224_n1488# 0.018226f
C362 plus.t8 a_n2224_n1488# 0.11719f
C363 plus.n42 a_n2224_n1488# 0.082107f
C364 plus.t10 a_n2224_n1488# 0.113025f
C365 plus.n43 a_n2224_n1488# 0.068301f
C366 plus.t6 a_n2224_n1488# 0.113025f
C367 plus.n44 a_n2224_n1488# 0.068301f
C368 plus.n45 a_n2224_n1488# 0.01983f
C369 plus.n46 a_n2224_n1488# 0.108183f
C370 plus.n47 a_n2224_n1488# 0.052039f
C371 plus.n48 a_n2224_n1488# 0.052039f
C372 plus.n49 a_n2224_n1488# 0.018867f
C373 plus.n50 a_n2224_n1488# 0.068301f
C374 plus.n51 a_n2224_n1488# 0.01983f
C375 plus.n52 a_n2224_n1488# 0.068301f
C376 plus.n53 a_n2224_n1488# 0.01983f
C377 plus.n54 a_n2224_n1488# 0.052039f
C378 plus.n55 a_n2224_n1488# 0.052039f
C379 plus.n56 a_n2224_n1488# 0.01983f
C380 plus.n57 a_n2224_n1488# 0.068301f
C381 plus.n58 a_n2224_n1488# 0.01983f
C382 plus.n59 a_n2224_n1488# 0.068301f
C383 plus.n60 a_n2224_n1488# 0.01983f
C384 plus.n61 a_n2224_n1488# 0.052039f
C385 plus.n62 a_n2224_n1488# 0.052039f
C386 plus.n63 a_n2224_n1488# 0.052039f
C387 plus.n64 a_n2224_n1488# 0.018226f
C388 plus.n65 a_n2224_n1488# 0.068301f
C389 plus.n66 a_n2224_n1488# 0.01983f
C390 plus.n67 a_n2224_n1488# 0.068301f
C391 plus.n68 a_n2224_n1488# 0.082041f
C392 plus.n69 a_n2224_n1488# 1.31557f
.ends

