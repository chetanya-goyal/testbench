* NGSPICE file created from diffpair427.ext - technology: sky130A

.subckt diffpair427 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t31 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 drain_left.t14 plus.t1 source.t30 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 source.t7 minus.t0 drain_right.t15 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X3 drain_left.t13 plus.t2 source.t23 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X4 source.t10 minus.t1 drain_right.t14 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X5 drain_right.t13 minus.t2 source.t9 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X7 drain_left.t12 plus.t3 source.t16 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X8 source.t26 plus.t4 drain_left.t11 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X9 source.t11 minus.t3 drain_right.t12 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 source.t18 plus.t5 drain_left.t10 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X11 source.t2 minus.t4 drain_right.t11 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X12 source.t0 minus.t5 drain_right.t10 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X13 drain_left.t9 plus.t6 source.t27 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X14 source.t19 plus.t7 drain_left.t8 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X15 source.t24 plus.t8 drain_left.t7 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X16 source.t22 plus.t9 drain_left.t6 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X17 a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X18 a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X19 drain_right.t9 minus.t6 source.t1 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X20 drain_right.t8 minus.t7 source.t4 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X21 drain_right.t7 minus.t8 source.t8 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X22 drain_left.t5 plus.t10 source.t28 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X23 drain_right.t6 minus.t9 source.t5 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X24 source.t17 plus.t11 drain_left.t4 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X25 source.t14 minus.t10 drain_right.t5 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X26 source.t15 minus.t11 drain_right.t4 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X27 source.t20 plus.t12 drain_left.t3 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X28 drain_right.t3 minus.t12 source.t6 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X29 drain_right.t2 minus.t13 source.t12 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X30 drain_left.t2 plus.t13 source.t21 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X31 drain_right.t1 minus.t14 source.t13 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X32 a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X33 drain_left.t1 plus.t14 source.t25 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X34 source.t3 minus.t15 drain_right.t0 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X35 source.t29 plus.t15 drain_left.t0 a_n1760_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n4 plus.t4 1323.02
R1 plus.n19 plus.t2 1323.02
R2 plus.n25 plus.t13 1323.02
R3 plus.n40 plus.t5 1323.02
R4 plus.n5 plus.t1 1282.12
R5 plus.n3 plus.t9 1282.12
R6 plus.n10 plus.t0 1282.12
R7 plus.n1 plus.t8 1282.12
R8 plus.n16 plus.t14 1282.12
R9 plus.n18 plus.t7 1282.12
R10 plus.n26 plus.t11 1282.12
R11 plus.n24 plus.t6 1282.12
R12 plus.n31 plus.t15 1282.12
R13 plus.n22 plus.t3 1282.12
R14 plus.n37 plus.t12 1282.12
R15 plus.n39 plus.t10 1282.12
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus plus.n41 29.6354
R47 plus.n6 plus.n5 29.2126
R48 plus.n18 plus.n17 29.2126
R49 plus.n39 plus.n38 29.2126
R50 plus.n27 plus.n26 29.2126
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 12.1103
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n546 source.n486 289.615
R73 source.n474 source.n414 289.615
R74 source.n408 source.n348 289.615
R75 source.n336 source.n276 289.615
R76 source.n60 source.n0 289.615
R77 source.n132 source.n72 289.615
R78 source.n198 source.n138 289.615
R79 source.n270 source.n210 289.615
R80 source.n506 source.n505 185
R81 source.n511 source.n510 185
R82 source.n513 source.n512 185
R83 source.n502 source.n501 185
R84 source.n519 source.n518 185
R85 source.n521 source.n520 185
R86 source.n498 source.n497 185
R87 source.n528 source.n527 185
R88 source.n529 source.n496 185
R89 source.n531 source.n530 185
R90 source.n494 source.n493 185
R91 source.n537 source.n536 185
R92 source.n539 source.n538 185
R93 source.n490 source.n489 185
R94 source.n545 source.n544 185
R95 source.n547 source.n546 185
R96 source.n434 source.n433 185
R97 source.n439 source.n438 185
R98 source.n441 source.n440 185
R99 source.n430 source.n429 185
R100 source.n447 source.n446 185
R101 source.n449 source.n448 185
R102 source.n426 source.n425 185
R103 source.n456 source.n455 185
R104 source.n457 source.n424 185
R105 source.n459 source.n458 185
R106 source.n422 source.n421 185
R107 source.n465 source.n464 185
R108 source.n467 source.n466 185
R109 source.n418 source.n417 185
R110 source.n473 source.n472 185
R111 source.n475 source.n474 185
R112 source.n368 source.n367 185
R113 source.n373 source.n372 185
R114 source.n375 source.n374 185
R115 source.n364 source.n363 185
R116 source.n381 source.n380 185
R117 source.n383 source.n382 185
R118 source.n360 source.n359 185
R119 source.n390 source.n389 185
R120 source.n391 source.n358 185
R121 source.n393 source.n392 185
R122 source.n356 source.n355 185
R123 source.n399 source.n398 185
R124 source.n401 source.n400 185
R125 source.n352 source.n351 185
R126 source.n407 source.n406 185
R127 source.n409 source.n408 185
R128 source.n296 source.n295 185
R129 source.n301 source.n300 185
R130 source.n303 source.n302 185
R131 source.n292 source.n291 185
R132 source.n309 source.n308 185
R133 source.n311 source.n310 185
R134 source.n288 source.n287 185
R135 source.n318 source.n317 185
R136 source.n319 source.n286 185
R137 source.n321 source.n320 185
R138 source.n284 source.n283 185
R139 source.n327 source.n326 185
R140 source.n329 source.n328 185
R141 source.n280 source.n279 185
R142 source.n335 source.n334 185
R143 source.n337 source.n336 185
R144 source.n61 source.n60 185
R145 source.n59 source.n58 185
R146 source.n4 source.n3 185
R147 source.n53 source.n52 185
R148 source.n51 source.n50 185
R149 source.n8 source.n7 185
R150 source.n45 source.n44 185
R151 source.n43 source.n10 185
R152 source.n42 source.n41 185
R153 source.n13 source.n11 185
R154 source.n36 source.n35 185
R155 source.n34 source.n33 185
R156 source.n17 source.n16 185
R157 source.n28 source.n27 185
R158 source.n26 source.n25 185
R159 source.n21 source.n20 185
R160 source.n133 source.n132 185
R161 source.n131 source.n130 185
R162 source.n76 source.n75 185
R163 source.n125 source.n124 185
R164 source.n123 source.n122 185
R165 source.n80 source.n79 185
R166 source.n117 source.n116 185
R167 source.n115 source.n82 185
R168 source.n114 source.n113 185
R169 source.n85 source.n83 185
R170 source.n108 source.n107 185
R171 source.n106 source.n105 185
R172 source.n89 source.n88 185
R173 source.n100 source.n99 185
R174 source.n98 source.n97 185
R175 source.n93 source.n92 185
R176 source.n199 source.n198 185
R177 source.n197 source.n196 185
R178 source.n142 source.n141 185
R179 source.n191 source.n190 185
R180 source.n189 source.n188 185
R181 source.n146 source.n145 185
R182 source.n183 source.n182 185
R183 source.n181 source.n148 185
R184 source.n180 source.n179 185
R185 source.n151 source.n149 185
R186 source.n174 source.n173 185
R187 source.n172 source.n171 185
R188 source.n155 source.n154 185
R189 source.n166 source.n165 185
R190 source.n164 source.n163 185
R191 source.n159 source.n158 185
R192 source.n271 source.n270 185
R193 source.n269 source.n268 185
R194 source.n214 source.n213 185
R195 source.n263 source.n262 185
R196 source.n261 source.n260 185
R197 source.n218 source.n217 185
R198 source.n255 source.n254 185
R199 source.n253 source.n220 185
R200 source.n252 source.n251 185
R201 source.n223 source.n221 185
R202 source.n246 source.n245 185
R203 source.n244 source.n243 185
R204 source.n227 source.n226 185
R205 source.n238 source.n237 185
R206 source.n236 source.n235 185
R207 source.n231 source.n230 185
R208 source.n507 source.t5 149.524
R209 source.n435 source.t3 149.524
R210 source.n369 source.t21 149.524
R211 source.n297 source.t18 149.524
R212 source.n22 source.t23 149.524
R213 source.n94 source.t26 149.524
R214 source.n160 source.t4 149.524
R215 source.n232 source.t2 149.524
R216 source.n511 source.n505 104.615
R217 source.n512 source.n511 104.615
R218 source.n512 source.n501 104.615
R219 source.n519 source.n501 104.615
R220 source.n520 source.n519 104.615
R221 source.n520 source.n497 104.615
R222 source.n528 source.n497 104.615
R223 source.n529 source.n528 104.615
R224 source.n530 source.n529 104.615
R225 source.n530 source.n493 104.615
R226 source.n537 source.n493 104.615
R227 source.n538 source.n537 104.615
R228 source.n538 source.n489 104.615
R229 source.n545 source.n489 104.615
R230 source.n546 source.n545 104.615
R231 source.n439 source.n433 104.615
R232 source.n440 source.n439 104.615
R233 source.n440 source.n429 104.615
R234 source.n447 source.n429 104.615
R235 source.n448 source.n447 104.615
R236 source.n448 source.n425 104.615
R237 source.n456 source.n425 104.615
R238 source.n457 source.n456 104.615
R239 source.n458 source.n457 104.615
R240 source.n458 source.n421 104.615
R241 source.n465 source.n421 104.615
R242 source.n466 source.n465 104.615
R243 source.n466 source.n417 104.615
R244 source.n473 source.n417 104.615
R245 source.n474 source.n473 104.615
R246 source.n373 source.n367 104.615
R247 source.n374 source.n373 104.615
R248 source.n374 source.n363 104.615
R249 source.n381 source.n363 104.615
R250 source.n382 source.n381 104.615
R251 source.n382 source.n359 104.615
R252 source.n390 source.n359 104.615
R253 source.n391 source.n390 104.615
R254 source.n392 source.n391 104.615
R255 source.n392 source.n355 104.615
R256 source.n399 source.n355 104.615
R257 source.n400 source.n399 104.615
R258 source.n400 source.n351 104.615
R259 source.n407 source.n351 104.615
R260 source.n408 source.n407 104.615
R261 source.n301 source.n295 104.615
R262 source.n302 source.n301 104.615
R263 source.n302 source.n291 104.615
R264 source.n309 source.n291 104.615
R265 source.n310 source.n309 104.615
R266 source.n310 source.n287 104.615
R267 source.n318 source.n287 104.615
R268 source.n319 source.n318 104.615
R269 source.n320 source.n319 104.615
R270 source.n320 source.n283 104.615
R271 source.n327 source.n283 104.615
R272 source.n328 source.n327 104.615
R273 source.n328 source.n279 104.615
R274 source.n335 source.n279 104.615
R275 source.n336 source.n335 104.615
R276 source.n60 source.n59 104.615
R277 source.n59 source.n3 104.615
R278 source.n52 source.n3 104.615
R279 source.n52 source.n51 104.615
R280 source.n51 source.n7 104.615
R281 source.n44 source.n7 104.615
R282 source.n44 source.n43 104.615
R283 source.n43 source.n42 104.615
R284 source.n42 source.n11 104.615
R285 source.n35 source.n11 104.615
R286 source.n35 source.n34 104.615
R287 source.n34 source.n16 104.615
R288 source.n27 source.n16 104.615
R289 source.n27 source.n26 104.615
R290 source.n26 source.n20 104.615
R291 source.n132 source.n131 104.615
R292 source.n131 source.n75 104.615
R293 source.n124 source.n75 104.615
R294 source.n124 source.n123 104.615
R295 source.n123 source.n79 104.615
R296 source.n116 source.n79 104.615
R297 source.n116 source.n115 104.615
R298 source.n115 source.n114 104.615
R299 source.n114 source.n83 104.615
R300 source.n107 source.n83 104.615
R301 source.n107 source.n106 104.615
R302 source.n106 source.n88 104.615
R303 source.n99 source.n88 104.615
R304 source.n99 source.n98 104.615
R305 source.n98 source.n92 104.615
R306 source.n198 source.n197 104.615
R307 source.n197 source.n141 104.615
R308 source.n190 source.n141 104.615
R309 source.n190 source.n189 104.615
R310 source.n189 source.n145 104.615
R311 source.n182 source.n145 104.615
R312 source.n182 source.n181 104.615
R313 source.n181 source.n180 104.615
R314 source.n180 source.n149 104.615
R315 source.n173 source.n149 104.615
R316 source.n173 source.n172 104.615
R317 source.n172 source.n154 104.615
R318 source.n165 source.n154 104.615
R319 source.n165 source.n164 104.615
R320 source.n164 source.n158 104.615
R321 source.n270 source.n269 104.615
R322 source.n269 source.n213 104.615
R323 source.n262 source.n213 104.615
R324 source.n262 source.n261 104.615
R325 source.n261 source.n217 104.615
R326 source.n254 source.n217 104.615
R327 source.n254 source.n253 104.615
R328 source.n253 source.n252 104.615
R329 source.n252 source.n221 104.615
R330 source.n245 source.n221 104.615
R331 source.n245 source.n244 104.615
R332 source.n244 source.n226 104.615
R333 source.n237 source.n226 104.615
R334 source.n237 source.n236 104.615
R335 source.n236 source.n230 104.615
R336 source.t5 source.n505 52.3082
R337 source.t3 source.n433 52.3082
R338 source.t21 source.n367 52.3082
R339 source.t18 source.n295 52.3082
R340 source.t23 source.n20 52.3082
R341 source.t26 source.n92 52.3082
R342 source.t4 source.n158 52.3082
R343 source.t2 source.n230 52.3082
R344 source.n67 source.n66 42.8739
R345 source.n69 source.n68 42.8739
R346 source.n71 source.n70 42.8739
R347 source.n205 source.n204 42.8739
R348 source.n207 source.n206 42.8739
R349 source.n209 source.n208 42.8739
R350 source.n485 source.n484 42.8737
R351 source.n483 source.n482 42.8737
R352 source.n481 source.n480 42.8737
R353 source.n347 source.n346 42.8737
R354 source.n345 source.n344 42.8737
R355 source.n343 source.n342 42.8737
R356 source.n551 source.n550 29.8581
R357 source.n479 source.n478 29.8581
R358 source.n413 source.n412 29.8581
R359 source.n341 source.n340 29.8581
R360 source.n65 source.n64 29.8581
R361 source.n137 source.n136 29.8581
R362 source.n203 source.n202 29.8581
R363 source.n275 source.n274 29.8581
R364 source.n341 source.n275 21.7877
R365 source.n552 source.n65 16.2748
R366 source.n531 source.n496 13.1884
R367 source.n459 source.n424 13.1884
R368 source.n393 source.n358 13.1884
R369 source.n321 source.n286 13.1884
R370 source.n45 source.n10 13.1884
R371 source.n117 source.n82 13.1884
R372 source.n183 source.n148 13.1884
R373 source.n255 source.n220 13.1884
R374 source.n527 source.n526 12.8005
R375 source.n532 source.n494 12.8005
R376 source.n455 source.n454 12.8005
R377 source.n460 source.n422 12.8005
R378 source.n389 source.n388 12.8005
R379 source.n394 source.n356 12.8005
R380 source.n317 source.n316 12.8005
R381 source.n322 source.n284 12.8005
R382 source.n46 source.n8 12.8005
R383 source.n41 source.n12 12.8005
R384 source.n118 source.n80 12.8005
R385 source.n113 source.n84 12.8005
R386 source.n184 source.n146 12.8005
R387 source.n179 source.n150 12.8005
R388 source.n256 source.n218 12.8005
R389 source.n251 source.n222 12.8005
R390 source.n525 source.n498 12.0247
R391 source.n536 source.n535 12.0247
R392 source.n453 source.n426 12.0247
R393 source.n464 source.n463 12.0247
R394 source.n387 source.n360 12.0247
R395 source.n398 source.n397 12.0247
R396 source.n315 source.n288 12.0247
R397 source.n326 source.n325 12.0247
R398 source.n50 source.n49 12.0247
R399 source.n40 source.n13 12.0247
R400 source.n122 source.n121 12.0247
R401 source.n112 source.n85 12.0247
R402 source.n188 source.n187 12.0247
R403 source.n178 source.n151 12.0247
R404 source.n260 source.n259 12.0247
R405 source.n250 source.n223 12.0247
R406 source.n522 source.n521 11.249
R407 source.n539 source.n492 11.249
R408 source.n450 source.n449 11.249
R409 source.n467 source.n420 11.249
R410 source.n384 source.n383 11.249
R411 source.n401 source.n354 11.249
R412 source.n312 source.n311 11.249
R413 source.n329 source.n282 11.249
R414 source.n53 source.n6 11.249
R415 source.n37 source.n36 11.249
R416 source.n125 source.n78 11.249
R417 source.n109 source.n108 11.249
R418 source.n191 source.n144 11.249
R419 source.n175 source.n174 11.249
R420 source.n263 source.n216 11.249
R421 source.n247 source.n246 11.249
R422 source.n518 source.n500 10.4732
R423 source.n540 source.n490 10.4732
R424 source.n446 source.n428 10.4732
R425 source.n468 source.n418 10.4732
R426 source.n380 source.n362 10.4732
R427 source.n402 source.n352 10.4732
R428 source.n308 source.n290 10.4732
R429 source.n330 source.n280 10.4732
R430 source.n54 source.n4 10.4732
R431 source.n33 source.n15 10.4732
R432 source.n126 source.n76 10.4732
R433 source.n105 source.n87 10.4732
R434 source.n192 source.n142 10.4732
R435 source.n171 source.n153 10.4732
R436 source.n264 source.n214 10.4732
R437 source.n243 source.n225 10.4732
R438 source.n507 source.n506 10.2747
R439 source.n435 source.n434 10.2747
R440 source.n369 source.n368 10.2747
R441 source.n297 source.n296 10.2747
R442 source.n22 source.n21 10.2747
R443 source.n94 source.n93 10.2747
R444 source.n160 source.n159 10.2747
R445 source.n232 source.n231 10.2747
R446 source.n517 source.n502 9.69747
R447 source.n544 source.n543 9.69747
R448 source.n445 source.n430 9.69747
R449 source.n472 source.n471 9.69747
R450 source.n379 source.n364 9.69747
R451 source.n406 source.n405 9.69747
R452 source.n307 source.n292 9.69747
R453 source.n334 source.n333 9.69747
R454 source.n58 source.n57 9.69747
R455 source.n32 source.n17 9.69747
R456 source.n130 source.n129 9.69747
R457 source.n104 source.n89 9.69747
R458 source.n196 source.n195 9.69747
R459 source.n170 source.n155 9.69747
R460 source.n268 source.n267 9.69747
R461 source.n242 source.n227 9.69747
R462 source.n550 source.n549 9.45567
R463 source.n478 source.n477 9.45567
R464 source.n412 source.n411 9.45567
R465 source.n340 source.n339 9.45567
R466 source.n64 source.n63 9.45567
R467 source.n136 source.n135 9.45567
R468 source.n202 source.n201 9.45567
R469 source.n274 source.n273 9.45567
R470 source.n549 source.n548 9.3005
R471 source.n488 source.n487 9.3005
R472 source.n543 source.n542 9.3005
R473 source.n541 source.n540 9.3005
R474 source.n492 source.n491 9.3005
R475 source.n535 source.n534 9.3005
R476 source.n533 source.n532 9.3005
R477 source.n509 source.n508 9.3005
R478 source.n504 source.n503 9.3005
R479 source.n515 source.n514 9.3005
R480 source.n517 source.n516 9.3005
R481 source.n500 source.n499 9.3005
R482 source.n523 source.n522 9.3005
R483 source.n525 source.n524 9.3005
R484 source.n526 source.n495 9.3005
R485 source.n477 source.n476 9.3005
R486 source.n416 source.n415 9.3005
R487 source.n471 source.n470 9.3005
R488 source.n469 source.n468 9.3005
R489 source.n420 source.n419 9.3005
R490 source.n463 source.n462 9.3005
R491 source.n461 source.n460 9.3005
R492 source.n437 source.n436 9.3005
R493 source.n432 source.n431 9.3005
R494 source.n443 source.n442 9.3005
R495 source.n445 source.n444 9.3005
R496 source.n428 source.n427 9.3005
R497 source.n451 source.n450 9.3005
R498 source.n453 source.n452 9.3005
R499 source.n454 source.n423 9.3005
R500 source.n411 source.n410 9.3005
R501 source.n350 source.n349 9.3005
R502 source.n405 source.n404 9.3005
R503 source.n403 source.n402 9.3005
R504 source.n354 source.n353 9.3005
R505 source.n397 source.n396 9.3005
R506 source.n395 source.n394 9.3005
R507 source.n371 source.n370 9.3005
R508 source.n366 source.n365 9.3005
R509 source.n377 source.n376 9.3005
R510 source.n379 source.n378 9.3005
R511 source.n362 source.n361 9.3005
R512 source.n385 source.n384 9.3005
R513 source.n387 source.n386 9.3005
R514 source.n388 source.n357 9.3005
R515 source.n339 source.n338 9.3005
R516 source.n278 source.n277 9.3005
R517 source.n333 source.n332 9.3005
R518 source.n331 source.n330 9.3005
R519 source.n282 source.n281 9.3005
R520 source.n325 source.n324 9.3005
R521 source.n323 source.n322 9.3005
R522 source.n299 source.n298 9.3005
R523 source.n294 source.n293 9.3005
R524 source.n305 source.n304 9.3005
R525 source.n307 source.n306 9.3005
R526 source.n290 source.n289 9.3005
R527 source.n313 source.n312 9.3005
R528 source.n315 source.n314 9.3005
R529 source.n316 source.n285 9.3005
R530 source.n24 source.n23 9.3005
R531 source.n19 source.n18 9.3005
R532 source.n30 source.n29 9.3005
R533 source.n32 source.n31 9.3005
R534 source.n15 source.n14 9.3005
R535 source.n38 source.n37 9.3005
R536 source.n40 source.n39 9.3005
R537 source.n12 source.n9 9.3005
R538 source.n63 source.n62 9.3005
R539 source.n2 source.n1 9.3005
R540 source.n57 source.n56 9.3005
R541 source.n55 source.n54 9.3005
R542 source.n6 source.n5 9.3005
R543 source.n49 source.n48 9.3005
R544 source.n47 source.n46 9.3005
R545 source.n96 source.n95 9.3005
R546 source.n91 source.n90 9.3005
R547 source.n102 source.n101 9.3005
R548 source.n104 source.n103 9.3005
R549 source.n87 source.n86 9.3005
R550 source.n110 source.n109 9.3005
R551 source.n112 source.n111 9.3005
R552 source.n84 source.n81 9.3005
R553 source.n135 source.n134 9.3005
R554 source.n74 source.n73 9.3005
R555 source.n129 source.n128 9.3005
R556 source.n127 source.n126 9.3005
R557 source.n78 source.n77 9.3005
R558 source.n121 source.n120 9.3005
R559 source.n119 source.n118 9.3005
R560 source.n162 source.n161 9.3005
R561 source.n157 source.n156 9.3005
R562 source.n168 source.n167 9.3005
R563 source.n170 source.n169 9.3005
R564 source.n153 source.n152 9.3005
R565 source.n176 source.n175 9.3005
R566 source.n178 source.n177 9.3005
R567 source.n150 source.n147 9.3005
R568 source.n201 source.n200 9.3005
R569 source.n140 source.n139 9.3005
R570 source.n195 source.n194 9.3005
R571 source.n193 source.n192 9.3005
R572 source.n144 source.n143 9.3005
R573 source.n187 source.n186 9.3005
R574 source.n185 source.n184 9.3005
R575 source.n234 source.n233 9.3005
R576 source.n229 source.n228 9.3005
R577 source.n240 source.n239 9.3005
R578 source.n242 source.n241 9.3005
R579 source.n225 source.n224 9.3005
R580 source.n248 source.n247 9.3005
R581 source.n250 source.n249 9.3005
R582 source.n222 source.n219 9.3005
R583 source.n273 source.n272 9.3005
R584 source.n212 source.n211 9.3005
R585 source.n267 source.n266 9.3005
R586 source.n265 source.n264 9.3005
R587 source.n216 source.n215 9.3005
R588 source.n259 source.n258 9.3005
R589 source.n257 source.n256 9.3005
R590 source.n514 source.n513 8.92171
R591 source.n547 source.n488 8.92171
R592 source.n442 source.n441 8.92171
R593 source.n475 source.n416 8.92171
R594 source.n376 source.n375 8.92171
R595 source.n409 source.n350 8.92171
R596 source.n304 source.n303 8.92171
R597 source.n337 source.n278 8.92171
R598 source.n61 source.n2 8.92171
R599 source.n29 source.n28 8.92171
R600 source.n133 source.n74 8.92171
R601 source.n101 source.n100 8.92171
R602 source.n199 source.n140 8.92171
R603 source.n167 source.n166 8.92171
R604 source.n271 source.n212 8.92171
R605 source.n239 source.n238 8.92171
R606 source.n510 source.n504 8.14595
R607 source.n548 source.n486 8.14595
R608 source.n438 source.n432 8.14595
R609 source.n476 source.n414 8.14595
R610 source.n372 source.n366 8.14595
R611 source.n410 source.n348 8.14595
R612 source.n300 source.n294 8.14595
R613 source.n338 source.n276 8.14595
R614 source.n62 source.n0 8.14595
R615 source.n25 source.n19 8.14595
R616 source.n134 source.n72 8.14595
R617 source.n97 source.n91 8.14595
R618 source.n200 source.n138 8.14595
R619 source.n163 source.n157 8.14595
R620 source.n272 source.n210 8.14595
R621 source.n235 source.n229 8.14595
R622 source.n509 source.n506 7.3702
R623 source.n437 source.n434 7.3702
R624 source.n371 source.n368 7.3702
R625 source.n299 source.n296 7.3702
R626 source.n24 source.n21 7.3702
R627 source.n96 source.n93 7.3702
R628 source.n162 source.n159 7.3702
R629 source.n234 source.n231 7.3702
R630 source.n510 source.n509 5.81868
R631 source.n550 source.n486 5.81868
R632 source.n438 source.n437 5.81868
R633 source.n478 source.n414 5.81868
R634 source.n372 source.n371 5.81868
R635 source.n412 source.n348 5.81868
R636 source.n300 source.n299 5.81868
R637 source.n340 source.n276 5.81868
R638 source.n64 source.n0 5.81868
R639 source.n25 source.n24 5.81868
R640 source.n136 source.n72 5.81868
R641 source.n97 source.n96 5.81868
R642 source.n202 source.n138 5.81868
R643 source.n163 source.n162 5.81868
R644 source.n274 source.n210 5.81868
R645 source.n235 source.n234 5.81868
R646 source.n552 source.n551 5.51343
R647 source.n513 source.n504 5.04292
R648 source.n548 source.n547 5.04292
R649 source.n441 source.n432 5.04292
R650 source.n476 source.n475 5.04292
R651 source.n375 source.n366 5.04292
R652 source.n410 source.n409 5.04292
R653 source.n303 source.n294 5.04292
R654 source.n338 source.n337 5.04292
R655 source.n62 source.n61 5.04292
R656 source.n28 source.n19 5.04292
R657 source.n134 source.n133 5.04292
R658 source.n100 source.n91 5.04292
R659 source.n200 source.n199 5.04292
R660 source.n166 source.n157 5.04292
R661 source.n272 source.n271 5.04292
R662 source.n238 source.n229 5.04292
R663 source.n514 source.n502 4.26717
R664 source.n544 source.n488 4.26717
R665 source.n442 source.n430 4.26717
R666 source.n472 source.n416 4.26717
R667 source.n376 source.n364 4.26717
R668 source.n406 source.n350 4.26717
R669 source.n304 source.n292 4.26717
R670 source.n334 source.n278 4.26717
R671 source.n58 source.n2 4.26717
R672 source.n29 source.n17 4.26717
R673 source.n130 source.n74 4.26717
R674 source.n101 source.n89 4.26717
R675 source.n196 source.n140 4.26717
R676 source.n167 source.n155 4.26717
R677 source.n268 source.n212 4.26717
R678 source.n239 source.n227 4.26717
R679 source.n518 source.n517 3.49141
R680 source.n543 source.n490 3.49141
R681 source.n446 source.n445 3.49141
R682 source.n471 source.n418 3.49141
R683 source.n380 source.n379 3.49141
R684 source.n405 source.n352 3.49141
R685 source.n308 source.n307 3.49141
R686 source.n333 source.n280 3.49141
R687 source.n57 source.n4 3.49141
R688 source.n33 source.n32 3.49141
R689 source.n129 source.n76 3.49141
R690 source.n105 source.n104 3.49141
R691 source.n195 source.n142 3.49141
R692 source.n171 source.n170 3.49141
R693 source.n267 source.n214 3.49141
R694 source.n243 source.n242 3.49141
R695 source.n508 source.n507 2.84303
R696 source.n436 source.n435 2.84303
R697 source.n370 source.n369 2.84303
R698 source.n298 source.n297 2.84303
R699 source.n23 source.n22 2.84303
R700 source.n95 source.n94 2.84303
R701 source.n161 source.n160 2.84303
R702 source.n233 source.n232 2.84303
R703 source.n521 source.n500 2.71565
R704 source.n540 source.n539 2.71565
R705 source.n449 source.n428 2.71565
R706 source.n468 source.n467 2.71565
R707 source.n383 source.n362 2.71565
R708 source.n402 source.n401 2.71565
R709 source.n311 source.n290 2.71565
R710 source.n330 source.n329 2.71565
R711 source.n54 source.n53 2.71565
R712 source.n36 source.n15 2.71565
R713 source.n126 source.n125 2.71565
R714 source.n108 source.n87 2.71565
R715 source.n192 source.n191 2.71565
R716 source.n174 source.n153 2.71565
R717 source.n264 source.n263 2.71565
R718 source.n246 source.n225 2.71565
R719 source.n522 source.n498 1.93989
R720 source.n536 source.n492 1.93989
R721 source.n450 source.n426 1.93989
R722 source.n464 source.n420 1.93989
R723 source.n384 source.n360 1.93989
R724 source.n398 source.n354 1.93989
R725 source.n312 source.n288 1.93989
R726 source.n326 source.n282 1.93989
R727 source.n50 source.n6 1.93989
R728 source.n37 source.n13 1.93989
R729 source.n122 source.n78 1.93989
R730 source.n109 source.n85 1.93989
R731 source.n188 source.n144 1.93989
R732 source.n175 source.n151 1.93989
R733 source.n260 source.n216 1.93989
R734 source.n247 source.n223 1.93989
R735 source.n484 source.t13 1.6505
R736 source.n484 source.t14 1.6505
R737 source.n482 source.t8 1.6505
R738 source.n482 source.t11 1.6505
R739 source.n480 source.t9 1.6505
R740 source.n480 source.t15 1.6505
R741 source.n346 source.t27 1.6505
R742 source.n346 source.t17 1.6505
R743 source.n344 source.t16 1.6505
R744 source.n344 source.t29 1.6505
R745 source.n342 source.t28 1.6505
R746 source.n342 source.t20 1.6505
R747 source.n66 source.t25 1.6505
R748 source.n66 source.t19 1.6505
R749 source.n68 source.t31 1.6505
R750 source.n68 source.t24 1.6505
R751 source.n70 source.t30 1.6505
R752 source.n70 source.t22 1.6505
R753 source.n204 source.t1 1.6505
R754 source.n204 source.t10 1.6505
R755 source.n206 source.t6 1.6505
R756 source.n206 source.t7 1.6505
R757 source.n208 source.t12 1.6505
R758 source.n208 source.t0 1.6505
R759 source.n527 source.n525 1.16414
R760 source.n535 source.n494 1.16414
R761 source.n455 source.n453 1.16414
R762 source.n463 source.n422 1.16414
R763 source.n389 source.n387 1.16414
R764 source.n397 source.n356 1.16414
R765 source.n317 source.n315 1.16414
R766 source.n325 source.n284 1.16414
R767 source.n49 source.n8 1.16414
R768 source.n41 source.n40 1.16414
R769 source.n121 source.n80 1.16414
R770 source.n113 source.n112 1.16414
R771 source.n187 source.n146 1.16414
R772 source.n179 source.n178 1.16414
R773 source.n259 source.n218 1.16414
R774 source.n251 source.n250 1.16414
R775 source.n275 source.n209 0.5005
R776 source.n209 source.n207 0.5005
R777 source.n207 source.n205 0.5005
R778 source.n205 source.n203 0.5005
R779 source.n137 source.n71 0.5005
R780 source.n71 source.n69 0.5005
R781 source.n69 source.n67 0.5005
R782 source.n67 source.n65 0.5005
R783 source.n343 source.n341 0.5005
R784 source.n345 source.n343 0.5005
R785 source.n347 source.n345 0.5005
R786 source.n413 source.n347 0.5005
R787 source.n481 source.n479 0.5005
R788 source.n483 source.n481 0.5005
R789 source.n485 source.n483 0.5005
R790 source.n551 source.n485 0.5005
R791 source.n203 source.n137 0.470328
R792 source.n479 source.n413 0.470328
R793 source.n526 source.n496 0.388379
R794 source.n532 source.n531 0.388379
R795 source.n454 source.n424 0.388379
R796 source.n460 source.n459 0.388379
R797 source.n388 source.n358 0.388379
R798 source.n394 source.n393 0.388379
R799 source.n316 source.n286 0.388379
R800 source.n322 source.n321 0.388379
R801 source.n46 source.n45 0.388379
R802 source.n12 source.n10 0.388379
R803 source.n118 source.n117 0.388379
R804 source.n84 source.n82 0.388379
R805 source.n184 source.n183 0.388379
R806 source.n150 source.n148 0.388379
R807 source.n256 source.n255 0.388379
R808 source.n222 source.n220 0.388379
R809 source source.n552 0.188
R810 source.n508 source.n503 0.155672
R811 source.n515 source.n503 0.155672
R812 source.n516 source.n515 0.155672
R813 source.n516 source.n499 0.155672
R814 source.n523 source.n499 0.155672
R815 source.n524 source.n523 0.155672
R816 source.n524 source.n495 0.155672
R817 source.n533 source.n495 0.155672
R818 source.n534 source.n533 0.155672
R819 source.n534 source.n491 0.155672
R820 source.n541 source.n491 0.155672
R821 source.n542 source.n541 0.155672
R822 source.n542 source.n487 0.155672
R823 source.n549 source.n487 0.155672
R824 source.n436 source.n431 0.155672
R825 source.n443 source.n431 0.155672
R826 source.n444 source.n443 0.155672
R827 source.n444 source.n427 0.155672
R828 source.n451 source.n427 0.155672
R829 source.n452 source.n451 0.155672
R830 source.n452 source.n423 0.155672
R831 source.n461 source.n423 0.155672
R832 source.n462 source.n461 0.155672
R833 source.n462 source.n419 0.155672
R834 source.n469 source.n419 0.155672
R835 source.n470 source.n469 0.155672
R836 source.n470 source.n415 0.155672
R837 source.n477 source.n415 0.155672
R838 source.n370 source.n365 0.155672
R839 source.n377 source.n365 0.155672
R840 source.n378 source.n377 0.155672
R841 source.n378 source.n361 0.155672
R842 source.n385 source.n361 0.155672
R843 source.n386 source.n385 0.155672
R844 source.n386 source.n357 0.155672
R845 source.n395 source.n357 0.155672
R846 source.n396 source.n395 0.155672
R847 source.n396 source.n353 0.155672
R848 source.n403 source.n353 0.155672
R849 source.n404 source.n403 0.155672
R850 source.n404 source.n349 0.155672
R851 source.n411 source.n349 0.155672
R852 source.n298 source.n293 0.155672
R853 source.n305 source.n293 0.155672
R854 source.n306 source.n305 0.155672
R855 source.n306 source.n289 0.155672
R856 source.n313 source.n289 0.155672
R857 source.n314 source.n313 0.155672
R858 source.n314 source.n285 0.155672
R859 source.n323 source.n285 0.155672
R860 source.n324 source.n323 0.155672
R861 source.n324 source.n281 0.155672
R862 source.n331 source.n281 0.155672
R863 source.n332 source.n331 0.155672
R864 source.n332 source.n277 0.155672
R865 source.n339 source.n277 0.155672
R866 source.n63 source.n1 0.155672
R867 source.n56 source.n1 0.155672
R868 source.n56 source.n55 0.155672
R869 source.n55 source.n5 0.155672
R870 source.n48 source.n5 0.155672
R871 source.n48 source.n47 0.155672
R872 source.n47 source.n9 0.155672
R873 source.n39 source.n9 0.155672
R874 source.n39 source.n38 0.155672
R875 source.n38 source.n14 0.155672
R876 source.n31 source.n14 0.155672
R877 source.n31 source.n30 0.155672
R878 source.n30 source.n18 0.155672
R879 source.n23 source.n18 0.155672
R880 source.n135 source.n73 0.155672
R881 source.n128 source.n73 0.155672
R882 source.n128 source.n127 0.155672
R883 source.n127 source.n77 0.155672
R884 source.n120 source.n77 0.155672
R885 source.n120 source.n119 0.155672
R886 source.n119 source.n81 0.155672
R887 source.n111 source.n81 0.155672
R888 source.n111 source.n110 0.155672
R889 source.n110 source.n86 0.155672
R890 source.n103 source.n86 0.155672
R891 source.n103 source.n102 0.155672
R892 source.n102 source.n90 0.155672
R893 source.n95 source.n90 0.155672
R894 source.n201 source.n139 0.155672
R895 source.n194 source.n139 0.155672
R896 source.n194 source.n193 0.155672
R897 source.n193 source.n143 0.155672
R898 source.n186 source.n143 0.155672
R899 source.n186 source.n185 0.155672
R900 source.n185 source.n147 0.155672
R901 source.n177 source.n147 0.155672
R902 source.n177 source.n176 0.155672
R903 source.n176 source.n152 0.155672
R904 source.n169 source.n152 0.155672
R905 source.n169 source.n168 0.155672
R906 source.n168 source.n156 0.155672
R907 source.n161 source.n156 0.155672
R908 source.n273 source.n211 0.155672
R909 source.n266 source.n211 0.155672
R910 source.n266 source.n265 0.155672
R911 source.n265 source.n215 0.155672
R912 source.n258 source.n215 0.155672
R913 source.n258 source.n257 0.155672
R914 source.n257 source.n219 0.155672
R915 source.n249 source.n219 0.155672
R916 source.n249 source.n248 0.155672
R917 source.n248 source.n224 0.155672
R918 source.n241 source.n224 0.155672
R919 source.n241 source.n240 0.155672
R920 source.n240 source.n228 0.155672
R921 source.n233 source.n228 0.155672
R922 drain_left.n9 drain_left.n7 60.0527
R923 drain_left.n5 drain_left.n3 60.0525
R924 drain_left.n2 drain_left.n0 60.0525
R925 drain_left.n11 drain_left.n10 59.5527
R926 drain_left.n9 drain_left.n8 59.5527
R927 drain_left.n5 drain_left.n4 59.5525
R928 drain_left.n2 drain_left.n1 59.5525
R929 drain_left.n13 drain_left.n12 59.5525
R930 drain_left drain_left.n6 30.6171
R931 drain_left drain_left.n13 6.15322
R932 drain_left.n3 drain_left.t4 1.6505
R933 drain_left.n3 drain_left.t2 1.6505
R934 drain_left.n4 drain_left.t0 1.6505
R935 drain_left.n4 drain_left.t9 1.6505
R936 drain_left.n1 drain_left.t3 1.6505
R937 drain_left.n1 drain_left.t12 1.6505
R938 drain_left.n0 drain_left.t10 1.6505
R939 drain_left.n0 drain_left.t5 1.6505
R940 drain_left.n12 drain_left.t8 1.6505
R941 drain_left.n12 drain_left.t13 1.6505
R942 drain_left.n10 drain_left.t7 1.6505
R943 drain_left.n10 drain_left.t1 1.6505
R944 drain_left.n8 drain_left.t6 1.6505
R945 drain_left.n8 drain_left.t15 1.6505
R946 drain_left.n7 drain_left.t11 1.6505
R947 drain_left.n7 drain_left.t14 1.6505
R948 drain_left.n11 drain_left.n9 0.5005
R949 drain_left.n13 drain_left.n11 0.5005
R950 drain_left.n6 drain_left.n5 0.195154
R951 drain_left.n6 drain_left.n2 0.195154
R952 minus.n19 minus.t4 1323.02
R953 minus.n4 minus.t7 1323.02
R954 minus.n40 minus.t9 1323.02
R955 minus.n25 minus.t15 1323.02
R956 minus.n18 minus.t13 1282.12
R957 minus.n16 minus.t5 1282.12
R958 minus.n1 minus.t12 1282.12
R959 minus.n10 minus.t0 1282.12
R960 minus.n3 minus.t6 1282.12
R961 minus.n5 minus.t1 1282.12
R962 minus.n39 minus.t10 1282.12
R963 minus.n37 minus.t14 1282.12
R964 minus.n22 minus.t3 1282.12
R965 minus.n31 minus.t8 1282.12
R966 minus.n24 minus.t11 1282.12
R967 minus.n26 minus.t2 1282.12
R968 minus.n7 minus.n4 161.489
R969 minus.n28 minus.n25 161.489
R970 minus.n20 minus.n19 161.3
R971 minus.n17 minus.n0 161.3
R972 minus.n15 minus.n14 161.3
R973 minus.n13 minus.n12 161.3
R974 minus.n11 minus.n2 161.3
R975 minus.n9 minus.n8 161.3
R976 minus.n7 minus.n6 161.3
R977 minus.n41 minus.n40 161.3
R978 minus.n38 minus.n21 161.3
R979 minus.n36 minus.n35 161.3
R980 minus.n34 minus.n33 161.3
R981 minus.n32 minus.n23 161.3
R982 minus.n30 minus.n29 161.3
R983 minus.n28 minus.n27 161.3
R984 minus.n12 minus.n11 73.0308
R985 minus.n33 minus.n32 73.0308
R986 minus.n15 minus.n1 67.1884
R987 minus.n10 minus.n9 67.1884
R988 minus.n31 minus.n30 67.1884
R989 minus.n36 minus.n22 67.1884
R990 minus.n17 minus.n16 55.5035
R991 minus.n6 minus.n3 55.5035
R992 minus.n27 minus.n24 55.5035
R993 minus.n38 minus.n37 55.5035
R994 minus.n19 minus.n18 43.8187
R995 minus.n5 minus.n4 43.8187
R996 minus.n26 minus.n25 43.8187
R997 minus.n40 minus.n39 43.8187
R998 minus.n42 minus.n20 35.7543
R999 minus.n18 minus.n17 29.2126
R1000 minus.n6 minus.n5 29.2126
R1001 minus.n27 minus.n26 29.2126
R1002 minus.n39 minus.n38 29.2126
R1003 minus.n16 minus.n15 17.5278
R1004 minus.n9 minus.n3 17.5278
R1005 minus.n30 minus.n24 17.5278
R1006 minus.n37 minus.n36 17.5278
R1007 minus.n42 minus.n41 6.46641
R1008 minus.n12 minus.n1 5.84292
R1009 minus.n11 minus.n10 5.84292
R1010 minus.n32 minus.n31 5.84292
R1011 minus.n33 minus.n22 5.84292
R1012 minus.n20 minus.n0 0.189894
R1013 minus.n14 minus.n0 0.189894
R1014 minus.n14 minus.n13 0.189894
R1015 minus.n13 minus.n2 0.189894
R1016 minus.n8 minus.n2 0.189894
R1017 minus.n8 minus.n7 0.189894
R1018 minus.n29 minus.n28 0.189894
R1019 minus.n29 minus.n23 0.189894
R1020 minus.n34 minus.n23 0.189894
R1021 minus.n35 minus.n34 0.189894
R1022 minus.n35 minus.n21 0.189894
R1023 minus.n41 minus.n21 0.189894
R1024 minus minus.n42 0.188
R1025 drain_right.n5 drain_right.n3 60.0525
R1026 drain_right.n2 drain_right.n0 60.0525
R1027 drain_right.n9 drain_right.n7 60.0525
R1028 drain_right.n9 drain_right.n8 59.5527
R1029 drain_right.n11 drain_right.n10 59.5527
R1030 drain_right.n13 drain_right.n12 59.5527
R1031 drain_right.n5 drain_right.n4 59.5525
R1032 drain_right.n2 drain_right.n1 59.5525
R1033 drain_right drain_right.n6 30.0638
R1034 drain_right drain_right.n13 6.15322
R1035 drain_right.n3 drain_right.t5 1.6505
R1036 drain_right.n3 drain_right.t6 1.6505
R1037 drain_right.n4 drain_right.t12 1.6505
R1038 drain_right.n4 drain_right.t1 1.6505
R1039 drain_right.n1 drain_right.t4 1.6505
R1040 drain_right.n1 drain_right.t7 1.6505
R1041 drain_right.n0 drain_right.t0 1.6505
R1042 drain_right.n0 drain_right.t13 1.6505
R1043 drain_right.n7 drain_right.t14 1.6505
R1044 drain_right.n7 drain_right.t8 1.6505
R1045 drain_right.n8 drain_right.t15 1.6505
R1046 drain_right.n8 drain_right.t9 1.6505
R1047 drain_right.n10 drain_right.t10 1.6505
R1048 drain_right.n10 drain_right.t3 1.6505
R1049 drain_right.n12 drain_right.t11 1.6505
R1050 drain_right.n12 drain_right.t2 1.6505
R1051 drain_right.n13 drain_right.n11 0.5005
R1052 drain_right.n11 drain_right.n9 0.5005
R1053 drain_right.n6 drain_right.n5 0.195154
R1054 drain_right.n6 drain_right.n2 0.195154
C0 source plus 4.83397f
C1 drain_left drain_right 0.897273f
C2 drain_left minus 0.171252f
C3 drain_left source 33.242f
C4 drain_left plus 5.35235f
C5 drain_right minus 5.18201f
C6 source drain_right 33.242f
C7 source minus 4.81993f
C8 drain_right plus 0.324551f
C9 plus minus 5.35017f
C10 drain_right a_n1760_n3288# 6.65055f
C11 drain_left a_n1760_n3288# 6.93179f
C12 source a_n1760_n3288# 8.642376f
C13 minus a_n1760_n3288# 6.850471f
C14 plus a_n1760_n3288# 8.88233f
C15 drain_right.t0 a_n1760_n3288# 0.340596f
C16 drain_right.t13 a_n1760_n3288# 0.340596f
C17 drain_right.n0 a_n1760_n3288# 3.03437f
C18 drain_right.t4 a_n1760_n3288# 0.340596f
C19 drain_right.t7 a_n1760_n3288# 0.340596f
C20 drain_right.n1 a_n1760_n3288# 3.03078f
C21 drain_right.n2 a_n1760_n3288# 0.814156f
C22 drain_right.t5 a_n1760_n3288# 0.340596f
C23 drain_right.t6 a_n1760_n3288# 0.340596f
C24 drain_right.n3 a_n1760_n3288# 3.03437f
C25 drain_right.t12 a_n1760_n3288# 0.340596f
C26 drain_right.t1 a_n1760_n3288# 0.340596f
C27 drain_right.n4 a_n1760_n3288# 3.03078f
C28 drain_right.n5 a_n1760_n3288# 0.814156f
C29 drain_right.n6 a_n1760_n3288# 1.64774f
C30 drain_right.t14 a_n1760_n3288# 0.340596f
C31 drain_right.t8 a_n1760_n3288# 0.340596f
C32 drain_right.n7 a_n1760_n3288# 3.03437f
C33 drain_right.t15 a_n1760_n3288# 0.340596f
C34 drain_right.t9 a_n1760_n3288# 0.340596f
C35 drain_right.n8 a_n1760_n3288# 3.03079f
C36 drain_right.n9 a_n1760_n3288# 0.845205f
C37 drain_right.t10 a_n1760_n3288# 0.340596f
C38 drain_right.t3 a_n1760_n3288# 0.340596f
C39 drain_right.n10 a_n1760_n3288# 3.03079f
C40 drain_right.n11 a_n1760_n3288# 0.41716f
C41 drain_right.t11 a_n1760_n3288# 0.340596f
C42 drain_right.t2 a_n1760_n3288# 0.340596f
C43 drain_right.n12 a_n1760_n3288# 3.03079f
C44 drain_right.n13 a_n1760_n3288# 0.713633f
C45 minus.n0 a_n1760_n3288# 0.052266f
C46 minus.t4 a_n1760_n3288# 0.448627f
C47 minus.t13 a_n1760_n3288# 0.443081f
C48 minus.t5 a_n1760_n3288# 0.443081f
C49 minus.t12 a_n1760_n3288# 0.443081f
C50 minus.n1 a_n1760_n3288# 0.178453f
C51 minus.n2 a_n1760_n3288# 0.052266f
C52 minus.t0 a_n1760_n3288# 0.443081f
C53 minus.t6 a_n1760_n3288# 0.443081f
C54 minus.n3 a_n1760_n3288# 0.178453f
C55 minus.t7 a_n1760_n3288# 0.448627f
C56 minus.n4 a_n1760_n3288# 0.193863f
C57 minus.t1 a_n1760_n3288# 0.443081f
C58 minus.n5 a_n1760_n3288# 0.178453f
C59 minus.n6 a_n1760_n3288# 0.019916f
C60 minus.n7 a_n1760_n3288# 0.114448f
C61 minus.n8 a_n1760_n3288# 0.052266f
C62 minus.n9 a_n1760_n3288# 0.019916f
C63 minus.n10 a_n1760_n3288# 0.178453f
C64 minus.n11 a_n1760_n3288# 0.018627f
C65 minus.n12 a_n1760_n3288# 0.018627f
C66 minus.n13 a_n1760_n3288# 0.052266f
C67 minus.n14 a_n1760_n3288# 0.052266f
C68 minus.n15 a_n1760_n3288# 0.019916f
C69 minus.n16 a_n1760_n3288# 0.178453f
C70 minus.n17 a_n1760_n3288# 0.019916f
C71 minus.n18 a_n1760_n3288# 0.178453f
C72 minus.n19 a_n1760_n3288# 0.19379f
C73 minus.n20 a_n1760_n3288# 1.81072f
C74 minus.n21 a_n1760_n3288# 0.052266f
C75 minus.t10 a_n1760_n3288# 0.443081f
C76 minus.t14 a_n1760_n3288# 0.443081f
C77 minus.t3 a_n1760_n3288# 0.443081f
C78 minus.n22 a_n1760_n3288# 0.178453f
C79 minus.n23 a_n1760_n3288# 0.052266f
C80 minus.t8 a_n1760_n3288# 0.443081f
C81 minus.t11 a_n1760_n3288# 0.443081f
C82 minus.n24 a_n1760_n3288# 0.178453f
C83 minus.t15 a_n1760_n3288# 0.448627f
C84 minus.n25 a_n1760_n3288# 0.193863f
C85 minus.t2 a_n1760_n3288# 0.443081f
C86 minus.n26 a_n1760_n3288# 0.178453f
C87 minus.n27 a_n1760_n3288# 0.019916f
C88 minus.n28 a_n1760_n3288# 0.114448f
C89 minus.n29 a_n1760_n3288# 0.052266f
C90 minus.n30 a_n1760_n3288# 0.019916f
C91 minus.n31 a_n1760_n3288# 0.178453f
C92 minus.n32 a_n1760_n3288# 0.018627f
C93 minus.n33 a_n1760_n3288# 0.018627f
C94 minus.n34 a_n1760_n3288# 0.052266f
C95 minus.n35 a_n1760_n3288# 0.052266f
C96 minus.n36 a_n1760_n3288# 0.019916f
C97 minus.n37 a_n1760_n3288# 0.178453f
C98 minus.n38 a_n1760_n3288# 0.019916f
C99 minus.n39 a_n1760_n3288# 0.178453f
C100 minus.t9 a_n1760_n3288# 0.448627f
C101 minus.n40 a_n1760_n3288# 0.19379f
C102 minus.n41 a_n1760_n3288# 0.337557f
C103 minus.n42 a_n1760_n3288# 2.20379f
C104 drain_left.t10 a_n1760_n3288# 0.341122f
C105 drain_left.t5 a_n1760_n3288# 0.341122f
C106 drain_left.n0 a_n1760_n3288# 3.03905f
C107 drain_left.t3 a_n1760_n3288# 0.341122f
C108 drain_left.t12 a_n1760_n3288# 0.341122f
C109 drain_left.n1 a_n1760_n3288# 3.03545f
C110 drain_left.n2 a_n1760_n3288# 0.815413f
C111 drain_left.t4 a_n1760_n3288# 0.341122f
C112 drain_left.t2 a_n1760_n3288# 0.341122f
C113 drain_left.n3 a_n1760_n3288# 3.03905f
C114 drain_left.t0 a_n1760_n3288# 0.341122f
C115 drain_left.t9 a_n1760_n3288# 0.341122f
C116 drain_left.n4 a_n1760_n3288# 3.03545f
C117 drain_left.n5 a_n1760_n3288# 0.815413f
C118 drain_left.n6 a_n1760_n3288# 1.725f
C119 drain_left.t11 a_n1760_n3288# 0.341122f
C120 drain_left.t14 a_n1760_n3288# 0.341122f
C121 drain_left.n7 a_n1760_n3288# 3.03907f
C122 drain_left.t6 a_n1760_n3288# 0.341122f
C123 drain_left.t15 a_n1760_n3288# 0.341122f
C124 drain_left.n8 a_n1760_n3288# 3.03547f
C125 drain_left.n9 a_n1760_n3288# 0.846497f
C126 drain_left.t7 a_n1760_n3288# 0.341122f
C127 drain_left.t1 a_n1760_n3288# 0.341122f
C128 drain_left.n10 a_n1760_n3288# 3.03547f
C129 drain_left.n11 a_n1760_n3288# 0.417804f
C130 drain_left.t8 a_n1760_n3288# 0.341122f
C131 drain_left.t13 a_n1760_n3288# 0.341122f
C132 drain_left.n12 a_n1760_n3288# 3.03545f
C133 drain_left.n13 a_n1760_n3288# 0.714747f
C134 source.n0 a_n1760_n3288# 0.039696f
C135 source.n1 a_n1760_n3288# 0.029968f
C136 source.n2 a_n1760_n3288# 0.016103f
C137 source.n3 a_n1760_n3288# 0.038062f
C138 source.n4 a_n1760_n3288# 0.017051f
C139 source.n5 a_n1760_n3288# 0.029968f
C140 source.n6 a_n1760_n3288# 0.016103f
C141 source.n7 a_n1760_n3288# 0.038062f
C142 source.n8 a_n1760_n3288# 0.017051f
C143 source.n9 a_n1760_n3288# 0.029968f
C144 source.n10 a_n1760_n3288# 0.016577f
C145 source.n11 a_n1760_n3288# 0.038062f
C146 source.n12 a_n1760_n3288# 0.016103f
C147 source.n13 a_n1760_n3288# 0.017051f
C148 source.n14 a_n1760_n3288# 0.029968f
C149 source.n15 a_n1760_n3288# 0.016103f
C150 source.n16 a_n1760_n3288# 0.038062f
C151 source.n17 a_n1760_n3288# 0.017051f
C152 source.n18 a_n1760_n3288# 0.029968f
C153 source.n19 a_n1760_n3288# 0.016103f
C154 source.n20 a_n1760_n3288# 0.028547f
C155 source.n21 a_n1760_n3288# 0.026907f
C156 source.t23 a_n1760_n3288# 0.064285f
C157 source.n22 a_n1760_n3288# 0.216063f
C158 source.n23 a_n1760_n3288# 1.51182f
C159 source.n24 a_n1760_n3288# 0.016103f
C160 source.n25 a_n1760_n3288# 0.017051f
C161 source.n26 a_n1760_n3288# 0.038062f
C162 source.n27 a_n1760_n3288# 0.038062f
C163 source.n28 a_n1760_n3288# 0.017051f
C164 source.n29 a_n1760_n3288# 0.016103f
C165 source.n30 a_n1760_n3288# 0.029968f
C166 source.n31 a_n1760_n3288# 0.029968f
C167 source.n32 a_n1760_n3288# 0.016103f
C168 source.n33 a_n1760_n3288# 0.017051f
C169 source.n34 a_n1760_n3288# 0.038062f
C170 source.n35 a_n1760_n3288# 0.038062f
C171 source.n36 a_n1760_n3288# 0.017051f
C172 source.n37 a_n1760_n3288# 0.016103f
C173 source.n38 a_n1760_n3288# 0.029968f
C174 source.n39 a_n1760_n3288# 0.029968f
C175 source.n40 a_n1760_n3288# 0.016103f
C176 source.n41 a_n1760_n3288# 0.017051f
C177 source.n42 a_n1760_n3288# 0.038062f
C178 source.n43 a_n1760_n3288# 0.038062f
C179 source.n44 a_n1760_n3288# 0.038062f
C180 source.n45 a_n1760_n3288# 0.016577f
C181 source.n46 a_n1760_n3288# 0.016103f
C182 source.n47 a_n1760_n3288# 0.029968f
C183 source.n48 a_n1760_n3288# 0.029968f
C184 source.n49 a_n1760_n3288# 0.016103f
C185 source.n50 a_n1760_n3288# 0.017051f
C186 source.n51 a_n1760_n3288# 0.038062f
C187 source.n52 a_n1760_n3288# 0.038062f
C188 source.n53 a_n1760_n3288# 0.017051f
C189 source.n54 a_n1760_n3288# 0.016103f
C190 source.n55 a_n1760_n3288# 0.029968f
C191 source.n56 a_n1760_n3288# 0.029968f
C192 source.n57 a_n1760_n3288# 0.016103f
C193 source.n58 a_n1760_n3288# 0.017051f
C194 source.n59 a_n1760_n3288# 0.038062f
C195 source.n60 a_n1760_n3288# 0.078108f
C196 source.n61 a_n1760_n3288# 0.017051f
C197 source.n62 a_n1760_n3288# 0.016103f
C198 source.n63 a_n1760_n3288# 0.064356f
C199 source.n64 a_n1760_n3288# 0.043107f
C200 source.n65 a_n1760_n3288# 1.19922f
C201 source.t25 a_n1760_n3288# 0.284176f
C202 source.t19 a_n1760_n3288# 0.284176f
C203 source.n66 a_n1760_n3288# 2.43312f
C204 source.n67 a_n1760_n3288# 0.402943f
C205 source.t31 a_n1760_n3288# 0.284176f
C206 source.t24 a_n1760_n3288# 0.284176f
C207 source.n68 a_n1760_n3288# 2.43312f
C208 source.n69 a_n1760_n3288# 0.402943f
C209 source.t30 a_n1760_n3288# 0.284176f
C210 source.t22 a_n1760_n3288# 0.284176f
C211 source.n70 a_n1760_n3288# 2.43312f
C212 source.n71 a_n1760_n3288# 0.402943f
C213 source.n72 a_n1760_n3288# 0.039696f
C214 source.n73 a_n1760_n3288# 0.029968f
C215 source.n74 a_n1760_n3288# 0.016103f
C216 source.n75 a_n1760_n3288# 0.038062f
C217 source.n76 a_n1760_n3288# 0.017051f
C218 source.n77 a_n1760_n3288# 0.029968f
C219 source.n78 a_n1760_n3288# 0.016103f
C220 source.n79 a_n1760_n3288# 0.038062f
C221 source.n80 a_n1760_n3288# 0.017051f
C222 source.n81 a_n1760_n3288# 0.029968f
C223 source.n82 a_n1760_n3288# 0.016577f
C224 source.n83 a_n1760_n3288# 0.038062f
C225 source.n84 a_n1760_n3288# 0.016103f
C226 source.n85 a_n1760_n3288# 0.017051f
C227 source.n86 a_n1760_n3288# 0.029968f
C228 source.n87 a_n1760_n3288# 0.016103f
C229 source.n88 a_n1760_n3288# 0.038062f
C230 source.n89 a_n1760_n3288# 0.017051f
C231 source.n90 a_n1760_n3288# 0.029968f
C232 source.n91 a_n1760_n3288# 0.016103f
C233 source.n92 a_n1760_n3288# 0.028547f
C234 source.n93 a_n1760_n3288# 0.026907f
C235 source.t26 a_n1760_n3288# 0.064285f
C236 source.n94 a_n1760_n3288# 0.216063f
C237 source.n95 a_n1760_n3288# 1.51182f
C238 source.n96 a_n1760_n3288# 0.016103f
C239 source.n97 a_n1760_n3288# 0.017051f
C240 source.n98 a_n1760_n3288# 0.038062f
C241 source.n99 a_n1760_n3288# 0.038062f
C242 source.n100 a_n1760_n3288# 0.017051f
C243 source.n101 a_n1760_n3288# 0.016103f
C244 source.n102 a_n1760_n3288# 0.029968f
C245 source.n103 a_n1760_n3288# 0.029968f
C246 source.n104 a_n1760_n3288# 0.016103f
C247 source.n105 a_n1760_n3288# 0.017051f
C248 source.n106 a_n1760_n3288# 0.038062f
C249 source.n107 a_n1760_n3288# 0.038062f
C250 source.n108 a_n1760_n3288# 0.017051f
C251 source.n109 a_n1760_n3288# 0.016103f
C252 source.n110 a_n1760_n3288# 0.029968f
C253 source.n111 a_n1760_n3288# 0.029968f
C254 source.n112 a_n1760_n3288# 0.016103f
C255 source.n113 a_n1760_n3288# 0.017051f
C256 source.n114 a_n1760_n3288# 0.038062f
C257 source.n115 a_n1760_n3288# 0.038062f
C258 source.n116 a_n1760_n3288# 0.038062f
C259 source.n117 a_n1760_n3288# 0.016577f
C260 source.n118 a_n1760_n3288# 0.016103f
C261 source.n119 a_n1760_n3288# 0.029968f
C262 source.n120 a_n1760_n3288# 0.029968f
C263 source.n121 a_n1760_n3288# 0.016103f
C264 source.n122 a_n1760_n3288# 0.017051f
C265 source.n123 a_n1760_n3288# 0.038062f
C266 source.n124 a_n1760_n3288# 0.038062f
C267 source.n125 a_n1760_n3288# 0.017051f
C268 source.n126 a_n1760_n3288# 0.016103f
C269 source.n127 a_n1760_n3288# 0.029968f
C270 source.n128 a_n1760_n3288# 0.029968f
C271 source.n129 a_n1760_n3288# 0.016103f
C272 source.n130 a_n1760_n3288# 0.017051f
C273 source.n131 a_n1760_n3288# 0.038062f
C274 source.n132 a_n1760_n3288# 0.078108f
C275 source.n133 a_n1760_n3288# 0.017051f
C276 source.n134 a_n1760_n3288# 0.016103f
C277 source.n135 a_n1760_n3288# 0.064356f
C278 source.n136 a_n1760_n3288# 0.043107f
C279 source.n137 a_n1760_n3288# 0.116476f
C280 source.n138 a_n1760_n3288# 0.039696f
C281 source.n139 a_n1760_n3288# 0.029968f
C282 source.n140 a_n1760_n3288# 0.016103f
C283 source.n141 a_n1760_n3288# 0.038062f
C284 source.n142 a_n1760_n3288# 0.017051f
C285 source.n143 a_n1760_n3288# 0.029968f
C286 source.n144 a_n1760_n3288# 0.016103f
C287 source.n145 a_n1760_n3288# 0.038062f
C288 source.n146 a_n1760_n3288# 0.017051f
C289 source.n147 a_n1760_n3288# 0.029968f
C290 source.n148 a_n1760_n3288# 0.016577f
C291 source.n149 a_n1760_n3288# 0.038062f
C292 source.n150 a_n1760_n3288# 0.016103f
C293 source.n151 a_n1760_n3288# 0.017051f
C294 source.n152 a_n1760_n3288# 0.029968f
C295 source.n153 a_n1760_n3288# 0.016103f
C296 source.n154 a_n1760_n3288# 0.038062f
C297 source.n155 a_n1760_n3288# 0.017051f
C298 source.n156 a_n1760_n3288# 0.029968f
C299 source.n157 a_n1760_n3288# 0.016103f
C300 source.n158 a_n1760_n3288# 0.028547f
C301 source.n159 a_n1760_n3288# 0.026907f
C302 source.t4 a_n1760_n3288# 0.064285f
C303 source.n160 a_n1760_n3288# 0.216063f
C304 source.n161 a_n1760_n3288# 1.51182f
C305 source.n162 a_n1760_n3288# 0.016103f
C306 source.n163 a_n1760_n3288# 0.017051f
C307 source.n164 a_n1760_n3288# 0.038062f
C308 source.n165 a_n1760_n3288# 0.038062f
C309 source.n166 a_n1760_n3288# 0.017051f
C310 source.n167 a_n1760_n3288# 0.016103f
C311 source.n168 a_n1760_n3288# 0.029968f
C312 source.n169 a_n1760_n3288# 0.029968f
C313 source.n170 a_n1760_n3288# 0.016103f
C314 source.n171 a_n1760_n3288# 0.017051f
C315 source.n172 a_n1760_n3288# 0.038062f
C316 source.n173 a_n1760_n3288# 0.038062f
C317 source.n174 a_n1760_n3288# 0.017051f
C318 source.n175 a_n1760_n3288# 0.016103f
C319 source.n176 a_n1760_n3288# 0.029968f
C320 source.n177 a_n1760_n3288# 0.029968f
C321 source.n178 a_n1760_n3288# 0.016103f
C322 source.n179 a_n1760_n3288# 0.017051f
C323 source.n180 a_n1760_n3288# 0.038062f
C324 source.n181 a_n1760_n3288# 0.038062f
C325 source.n182 a_n1760_n3288# 0.038062f
C326 source.n183 a_n1760_n3288# 0.016577f
C327 source.n184 a_n1760_n3288# 0.016103f
C328 source.n185 a_n1760_n3288# 0.029968f
C329 source.n186 a_n1760_n3288# 0.029968f
C330 source.n187 a_n1760_n3288# 0.016103f
C331 source.n188 a_n1760_n3288# 0.017051f
C332 source.n189 a_n1760_n3288# 0.038062f
C333 source.n190 a_n1760_n3288# 0.038062f
C334 source.n191 a_n1760_n3288# 0.017051f
C335 source.n192 a_n1760_n3288# 0.016103f
C336 source.n193 a_n1760_n3288# 0.029968f
C337 source.n194 a_n1760_n3288# 0.029968f
C338 source.n195 a_n1760_n3288# 0.016103f
C339 source.n196 a_n1760_n3288# 0.017051f
C340 source.n197 a_n1760_n3288# 0.038062f
C341 source.n198 a_n1760_n3288# 0.078108f
C342 source.n199 a_n1760_n3288# 0.017051f
C343 source.n200 a_n1760_n3288# 0.016103f
C344 source.n201 a_n1760_n3288# 0.064356f
C345 source.n202 a_n1760_n3288# 0.043107f
C346 source.n203 a_n1760_n3288# 0.116476f
C347 source.t1 a_n1760_n3288# 0.284176f
C348 source.t10 a_n1760_n3288# 0.284176f
C349 source.n204 a_n1760_n3288# 2.43312f
C350 source.n205 a_n1760_n3288# 0.402943f
C351 source.t6 a_n1760_n3288# 0.284176f
C352 source.t7 a_n1760_n3288# 0.284176f
C353 source.n206 a_n1760_n3288# 2.43312f
C354 source.n207 a_n1760_n3288# 0.402943f
C355 source.t12 a_n1760_n3288# 0.284176f
C356 source.t0 a_n1760_n3288# 0.284176f
C357 source.n208 a_n1760_n3288# 2.43312f
C358 source.n209 a_n1760_n3288# 0.402943f
C359 source.n210 a_n1760_n3288# 0.039696f
C360 source.n211 a_n1760_n3288# 0.029968f
C361 source.n212 a_n1760_n3288# 0.016103f
C362 source.n213 a_n1760_n3288# 0.038062f
C363 source.n214 a_n1760_n3288# 0.017051f
C364 source.n215 a_n1760_n3288# 0.029968f
C365 source.n216 a_n1760_n3288# 0.016103f
C366 source.n217 a_n1760_n3288# 0.038062f
C367 source.n218 a_n1760_n3288# 0.017051f
C368 source.n219 a_n1760_n3288# 0.029968f
C369 source.n220 a_n1760_n3288# 0.016577f
C370 source.n221 a_n1760_n3288# 0.038062f
C371 source.n222 a_n1760_n3288# 0.016103f
C372 source.n223 a_n1760_n3288# 0.017051f
C373 source.n224 a_n1760_n3288# 0.029968f
C374 source.n225 a_n1760_n3288# 0.016103f
C375 source.n226 a_n1760_n3288# 0.038062f
C376 source.n227 a_n1760_n3288# 0.017051f
C377 source.n228 a_n1760_n3288# 0.029968f
C378 source.n229 a_n1760_n3288# 0.016103f
C379 source.n230 a_n1760_n3288# 0.028547f
C380 source.n231 a_n1760_n3288# 0.026907f
C381 source.t2 a_n1760_n3288# 0.064285f
C382 source.n232 a_n1760_n3288# 0.216063f
C383 source.n233 a_n1760_n3288# 1.51182f
C384 source.n234 a_n1760_n3288# 0.016103f
C385 source.n235 a_n1760_n3288# 0.017051f
C386 source.n236 a_n1760_n3288# 0.038062f
C387 source.n237 a_n1760_n3288# 0.038062f
C388 source.n238 a_n1760_n3288# 0.017051f
C389 source.n239 a_n1760_n3288# 0.016103f
C390 source.n240 a_n1760_n3288# 0.029968f
C391 source.n241 a_n1760_n3288# 0.029968f
C392 source.n242 a_n1760_n3288# 0.016103f
C393 source.n243 a_n1760_n3288# 0.017051f
C394 source.n244 a_n1760_n3288# 0.038062f
C395 source.n245 a_n1760_n3288# 0.038062f
C396 source.n246 a_n1760_n3288# 0.017051f
C397 source.n247 a_n1760_n3288# 0.016103f
C398 source.n248 a_n1760_n3288# 0.029968f
C399 source.n249 a_n1760_n3288# 0.029968f
C400 source.n250 a_n1760_n3288# 0.016103f
C401 source.n251 a_n1760_n3288# 0.017051f
C402 source.n252 a_n1760_n3288# 0.038062f
C403 source.n253 a_n1760_n3288# 0.038062f
C404 source.n254 a_n1760_n3288# 0.038062f
C405 source.n255 a_n1760_n3288# 0.016577f
C406 source.n256 a_n1760_n3288# 0.016103f
C407 source.n257 a_n1760_n3288# 0.029968f
C408 source.n258 a_n1760_n3288# 0.029968f
C409 source.n259 a_n1760_n3288# 0.016103f
C410 source.n260 a_n1760_n3288# 0.017051f
C411 source.n261 a_n1760_n3288# 0.038062f
C412 source.n262 a_n1760_n3288# 0.038062f
C413 source.n263 a_n1760_n3288# 0.017051f
C414 source.n264 a_n1760_n3288# 0.016103f
C415 source.n265 a_n1760_n3288# 0.029968f
C416 source.n266 a_n1760_n3288# 0.029968f
C417 source.n267 a_n1760_n3288# 0.016103f
C418 source.n268 a_n1760_n3288# 0.017051f
C419 source.n269 a_n1760_n3288# 0.038062f
C420 source.n270 a_n1760_n3288# 0.078108f
C421 source.n271 a_n1760_n3288# 0.017051f
C422 source.n272 a_n1760_n3288# 0.016103f
C423 source.n273 a_n1760_n3288# 0.064356f
C424 source.n274 a_n1760_n3288# 0.043107f
C425 source.n275 a_n1760_n3288# 1.66894f
C426 source.n276 a_n1760_n3288# 0.039696f
C427 source.n277 a_n1760_n3288# 0.029968f
C428 source.n278 a_n1760_n3288# 0.016103f
C429 source.n279 a_n1760_n3288# 0.038062f
C430 source.n280 a_n1760_n3288# 0.017051f
C431 source.n281 a_n1760_n3288# 0.029968f
C432 source.n282 a_n1760_n3288# 0.016103f
C433 source.n283 a_n1760_n3288# 0.038062f
C434 source.n284 a_n1760_n3288# 0.017051f
C435 source.n285 a_n1760_n3288# 0.029968f
C436 source.n286 a_n1760_n3288# 0.016577f
C437 source.n287 a_n1760_n3288# 0.038062f
C438 source.n288 a_n1760_n3288# 0.017051f
C439 source.n289 a_n1760_n3288# 0.029968f
C440 source.n290 a_n1760_n3288# 0.016103f
C441 source.n291 a_n1760_n3288# 0.038062f
C442 source.n292 a_n1760_n3288# 0.017051f
C443 source.n293 a_n1760_n3288# 0.029968f
C444 source.n294 a_n1760_n3288# 0.016103f
C445 source.n295 a_n1760_n3288# 0.028547f
C446 source.n296 a_n1760_n3288# 0.026907f
C447 source.t18 a_n1760_n3288# 0.064285f
C448 source.n297 a_n1760_n3288# 0.216063f
C449 source.n298 a_n1760_n3288# 1.51182f
C450 source.n299 a_n1760_n3288# 0.016103f
C451 source.n300 a_n1760_n3288# 0.017051f
C452 source.n301 a_n1760_n3288# 0.038062f
C453 source.n302 a_n1760_n3288# 0.038062f
C454 source.n303 a_n1760_n3288# 0.017051f
C455 source.n304 a_n1760_n3288# 0.016103f
C456 source.n305 a_n1760_n3288# 0.029968f
C457 source.n306 a_n1760_n3288# 0.029968f
C458 source.n307 a_n1760_n3288# 0.016103f
C459 source.n308 a_n1760_n3288# 0.017051f
C460 source.n309 a_n1760_n3288# 0.038062f
C461 source.n310 a_n1760_n3288# 0.038062f
C462 source.n311 a_n1760_n3288# 0.017051f
C463 source.n312 a_n1760_n3288# 0.016103f
C464 source.n313 a_n1760_n3288# 0.029968f
C465 source.n314 a_n1760_n3288# 0.029968f
C466 source.n315 a_n1760_n3288# 0.016103f
C467 source.n316 a_n1760_n3288# 0.016103f
C468 source.n317 a_n1760_n3288# 0.017051f
C469 source.n318 a_n1760_n3288# 0.038062f
C470 source.n319 a_n1760_n3288# 0.038062f
C471 source.n320 a_n1760_n3288# 0.038062f
C472 source.n321 a_n1760_n3288# 0.016577f
C473 source.n322 a_n1760_n3288# 0.016103f
C474 source.n323 a_n1760_n3288# 0.029968f
C475 source.n324 a_n1760_n3288# 0.029968f
C476 source.n325 a_n1760_n3288# 0.016103f
C477 source.n326 a_n1760_n3288# 0.017051f
C478 source.n327 a_n1760_n3288# 0.038062f
C479 source.n328 a_n1760_n3288# 0.038062f
C480 source.n329 a_n1760_n3288# 0.017051f
C481 source.n330 a_n1760_n3288# 0.016103f
C482 source.n331 a_n1760_n3288# 0.029968f
C483 source.n332 a_n1760_n3288# 0.029968f
C484 source.n333 a_n1760_n3288# 0.016103f
C485 source.n334 a_n1760_n3288# 0.017051f
C486 source.n335 a_n1760_n3288# 0.038062f
C487 source.n336 a_n1760_n3288# 0.078108f
C488 source.n337 a_n1760_n3288# 0.017051f
C489 source.n338 a_n1760_n3288# 0.016103f
C490 source.n339 a_n1760_n3288# 0.064356f
C491 source.n340 a_n1760_n3288# 0.043107f
C492 source.n341 a_n1760_n3288# 1.66894f
C493 source.t28 a_n1760_n3288# 0.284176f
C494 source.t20 a_n1760_n3288# 0.284176f
C495 source.n342 a_n1760_n3288# 2.43311f
C496 source.n343 a_n1760_n3288# 0.402958f
C497 source.t16 a_n1760_n3288# 0.284176f
C498 source.t29 a_n1760_n3288# 0.284176f
C499 source.n344 a_n1760_n3288# 2.43311f
C500 source.n345 a_n1760_n3288# 0.402958f
C501 source.t27 a_n1760_n3288# 0.284176f
C502 source.t17 a_n1760_n3288# 0.284176f
C503 source.n346 a_n1760_n3288# 2.43311f
C504 source.n347 a_n1760_n3288# 0.402958f
C505 source.n348 a_n1760_n3288# 0.039696f
C506 source.n349 a_n1760_n3288# 0.029968f
C507 source.n350 a_n1760_n3288# 0.016103f
C508 source.n351 a_n1760_n3288# 0.038062f
C509 source.n352 a_n1760_n3288# 0.017051f
C510 source.n353 a_n1760_n3288# 0.029968f
C511 source.n354 a_n1760_n3288# 0.016103f
C512 source.n355 a_n1760_n3288# 0.038062f
C513 source.n356 a_n1760_n3288# 0.017051f
C514 source.n357 a_n1760_n3288# 0.029968f
C515 source.n358 a_n1760_n3288# 0.016577f
C516 source.n359 a_n1760_n3288# 0.038062f
C517 source.n360 a_n1760_n3288# 0.017051f
C518 source.n361 a_n1760_n3288# 0.029968f
C519 source.n362 a_n1760_n3288# 0.016103f
C520 source.n363 a_n1760_n3288# 0.038062f
C521 source.n364 a_n1760_n3288# 0.017051f
C522 source.n365 a_n1760_n3288# 0.029968f
C523 source.n366 a_n1760_n3288# 0.016103f
C524 source.n367 a_n1760_n3288# 0.028547f
C525 source.n368 a_n1760_n3288# 0.026907f
C526 source.t21 a_n1760_n3288# 0.064285f
C527 source.n369 a_n1760_n3288# 0.216063f
C528 source.n370 a_n1760_n3288# 1.51182f
C529 source.n371 a_n1760_n3288# 0.016103f
C530 source.n372 a_n1760_n3288# 0.017051f
C531 source.n373 a_n1760_n3288# 0.038062f
C532 source.n374 a_n1760_n3288# 0.038062f
C533 source.n375 a_n1760_n3288# 0.017051f
C534 source.n376 a_n1760_n3288# 0.016103f
C535 source.n377 a_n1760_n3288# 0.029968f
C536 source.n378 a_n1760_n3288# 0.029968f
C537 source.n379 a_n1760_n3288# 0.016103f
C538 source.n380 a_n1760_n3288# 0.017051f
C539 source.n381 a_n1760_n3288# 0.038062f
C540 source.n382 a_n1760_n3288# 0.038062f
C541 source.n383 a_n1760_n3288# 0.017051f
C542 source.n384 a_n1760_n3288# 0.016103f
C543 source.n385 a_n1760_n3288# 0.029968f
C544 source.n386 a_n1760_n3288# 0.029968f
C545 source.n387 a_n1760_n3288# 0.016103f
C546 source.n388 a_n1760_n3288# 0.016103f
C547 source.n389 a_n1760_n3288# 0.017051f
C548 source.n390 a_n1760_n3288# 0.038062f
C549 source.n391 a_n1760_n3288# 0.038062f
C550 source.n392 a_n1760_n3288# 0.038062f
C551 source.n393 a_n1760_n3288# 0.016577f
C552 source.n394 a_n1760_n3288# 0.016103f
C553 source.n395 a_n1760_n3288# 0.029968f
C554 source.n396 a_n1760_n3288# 0.029968f
C555 source.n397 a_n1760_n3288# 0.016103f
C556 source.n398 a_n1760_n3288# 0.017051f
C557 source.n399 a_n1760_n3288# 0.038062f
C558 source.n400 a_n1760_n3288# 0.038062f
C559 source.n401 a_n1760_n3288# 0.017051f
C560 source.n402 a_n1760_n3288# 0.016103f
C561 source.n403 a_n1760_n3288# 0.029968f
C562 source.n404 a_n1760_n3288# 0.029968f
C563 source.n405 a_n1760_n3288# 0.016103f
C564 source.n406 a_n1760_n3288# 0.017051f
C565 source.n407 a_n1760_n3288# 0.038062f
C566 source.n408 a_n1760_n3288# 0.078108f
C567 source.n409 a_n1760_n3288# 0.017051f
C568 source.n410 a_n1760_n3288# 0.016103f
C569 source.n411 a_n1760_n3288# 0.064356f
C570 source.n412 a_n1760_n3288# 0.043107f
C571 source.n413 a_n1760_n3288# 0.116476f
C572 source.n414 a_n1760_n3288# 0.039696f
C573 source.n415 a_n1760_n3288# 0.029968f
C574 source.n416 a_n1760_n3288# 0.016103f
C575 source.n417 a_n1760_n3288# 0.038062f
C576 source.n418 a_n1760_n3288# 0.017051f
C577 source.n419 a_n1760_n3288# 0.029968f
C578 source.n420 a_n1760_n3288# 0.016103f
C579 source.n421 a_n1760_n3288# 0.038062f
C580 source.n422 a_n1760_n3288# 0.017051f
C581 source.n423 a_n1760_n3288# 0.029968f
C582 source.n424 a_n1760_n3288# 0.016577f
C583 source.n425 a_n1760_n3288# 0.038062f
C584 source.n426 a_n1760_n3288# 0.017051f
C585 source.n427 a_n1760_n3288# 0.029968f
C586 source.n428 a_n1760_n3288# 0.016103f
C587 source.n429 a_n1760_n3288# 0.038062f
C588 source.n430 a_n1760_n3288# 0.017051f
C589 source.n431 a_n1760_n3288# 0.029968f
C590 source.n432 a_n1760_n3288# 0.016103f
C591 source.n433 a_n1760_n3288# 0.028547f
C592 source.n434 a_n1760_n3288# 0.026907f
C593 source.t3 a_n1760_n3288# 0.064285f
C594 source.n435 a_n1760_n3288# 0.216063f
C595 source.n436 a_n1760_n3288# 1.51182f
C596 source.n437 a_n1760_n3288# 0.016103f
C597 source.n438 a_n1760_n3288# 0.017051f
C598 source.n439 a_n1760_n3288# 0.038062f
C599 source.n440 a_n1760_n3288# 0.038062f
C600 source.n441 a_n1760_n3288# 0.017051f
C601 source.n442 a_n1760_n3288# 0.016103f
C602 source.n443 a_n1760_n3288# 0.029968f
C603 source.n444 a_n1760_n3288# 0.029968f
C604 source.n445 a_n1760_n3288# 0.016103f
C605 source.n446 a_n1760_n3288# 0.017051f
C606 source.n447 a_n1760_n3288# 0.038062f
C607 source.n448 a_n1760_n3288# 0.038062f
C608 source.n449 a_n1760_n3288# 0.017051f
C609 source.n450 a_n1760_n3288# 0.016103f
C610 source.n451 a_n1760_n3288# 0.029968f
C611 source.n452 a_n1760_n3288# 0.029968f
C612 source.n453 a_n1760_n3288# 0.016103f
C613 source.n454 a_n1760_n3288# 0.016103f
C614 source.n455 a_n1760_n3288# 0.017051f
C615 source.n456 a_n1760_n3288# 0.038062f
C616 source.n457 a_n1760_n3288# 0.038062f
C617 source.n458 a_n1760_n3288# 0.038062f
C618 source.n459 a_n1760_n3288# 0.016577f
C619 source.n460 a_n1760_n3288# 0.016103f
C620 source.n461 a_n1760_n3288# 0.029968f
C621 source.n462 a_n1760_n3288# 0.029968f
C622 source.n463 a_n1760_n3288# 0.016103f
C623 source.n464 a_n1760_n3288# 0.017051f
C624 source.n465 a_n1760_n3288# 0.038062f
C625 source.n466 a_n1760_n3288# 0.038062f
C626 source.n467 a_n1760_n3288# 0.017051f
C627 source.n468 a_n1760_n3288# 0.016103f
C628 source.n469 a_n1760_n3288# 0.029968f
C629 source.n470 a_n1760_n3288# 0.029968f
C630 source.n471 a_n1760_n3288# 0.016103f
C631 source.n472 a_n1760_n3288# 0.017051f
C632 source.n473 a_n1760_n3288# 0.038062f
C633 source.n474 a_n1760_n3288# 0.078108f
C634 source.n475 a_n1760_n3288# 0.017051f
C635 source.n476 a_n1760_n3288# 0.016103f
C636 source.n477 a_n1760_n3288# 0.064356f
C637 source.n478 a_n1760_n3288# 0.043107f
C638 source.n479 a_n1760_n3288# 0.116476f
C639 source.t9 a_n1760_n3288# 0.284176f
C640 source.t15 a_n1760_n3288# 0.284176f
C641 source.n480 a_n1760_n3288# 2.43311f
C642 source.n481 a_n1760_n3288# 0.402958f
C643 source.t8 a_n1760_n3288# 0.284176f
C644 source.t11 a_n1760_n3288# 0.284176f
C645 source.n482 a_n1760_n3288# 2.43311f
C646 source.n483 a_n1760_n3288# 0.402958f
C647 source.t13 a_n1760_n3288# 0.284176f
C648 source.t14 a_n1760_n3288# 0.284176f
C649 source.n484 a_n1760_n3288# 2.43311f
C650 source.n485 a_n1760_n3288# 0.402958f
C651 source.n486 a_n1760_n3288# 0.039696f
C652 source.n487 a_n1760_n3288# 0.029968f
C653 source.n488 a_n1760_n3288# 0.016103f
C654 source.n489 a_n1760_n3288# 0.038062f
C655 source.n490 a_n1760_n3288# 0.017051f
C656 source.n491 a_n1760_n3288# 0.029968f
C657 source.n492 a_n1760_n3288# 0.016103f
C658 source.n493 a_n1760_n3288# 0.038062f
C659 source.n494 a_n1760_n3288# 0.017051f
C660 source.n495 a_n1760_n3288# 0.029968f
C661 source.n496 a_n1760_n3288# 0.016577f
C662 source.n497 a_n1760_n3288# 0.038062f
C663 source.n498 a_n1760_n3288# 0.017051f
C664 source.n499 a_n1760_n3288# 0.029968f
C665 source.n500 a_n1760_n3288# 0.016103f
C666 source.n501 a_n1760_n3288# 0.038062f
C667 source.n502 a_n1760_n3288# 0.017051f
C668 source.n503 a_n1760_n3288# 0.029968f
C669 source.n504 a_n1760_n3288# 0.016103f
C670 source.n505 a_n1760_n3288# 0.028547f
C671 source.n506 a_n1760_n3288# 0.026907f
C672 source.t5 a_n1760_n3288# 0.064285f
C673 source.n507 a_n1760_n3288# 0.216063f
C674 source.n508 a_n1760_n3288# 1.51182f
C675 source.n509 a_n1760_n3288# 0.016103f
C676 source.n510 a_n1760_n3288# 0.017051f
C677 source.n511 a_n1760_n3288# 0.038062f
C678 source.n512 a_n1760_n3288# 0.038062f
C679 source.n513 a_n1760_n3288# 0.017051f
C680 source.n514 a_n1760_n3288# 0.016103f
C681 source.n515 a_n1760_n3288# 0.029968f
C682 source.n516 a_n1760_n3288# 0.029968f
C683 source.n517 a_n1760_n3288# 0.016103f
C684 source.n518 a_n1760_n3288# 0.017051f
C685 source.n519 a_n1760_n3288# 0.038062f
C686 source.n520 a_n1760_n3288# 0.038062f
C687 source.n521 a_n1760_n3288# 0.017051f
C688 source.n522 a_n1760_n3288# 0.016103f
C689 source.n523 a_n1760_n3288# 0.029968f
C690 source.n524 a_n1760_n3288# 0.029968f
C691 source.n525 a_n1760_n3288# 0.016103f
C692 source.n526 a_n1760_n3288# 0.016103f
C693 source.n527 a_n1760_n3288# 0.017051f
C694 source.n528 a_n1760_n3288# 0.038062f
C695 source.n529 a_n1760_n3288# 0.038062f
C696 source.n530 a_n1760_n3288# 0.038062f
C697 source.n531 a_n1760_n3288# 0.016577f
C698 source.n532 a_n1760_n3288# 0.016103f
C699 source.n533 a_n1760_n3288# 0.029968f
C700 source.n534 a_n1760_n3288# 0.029968f
C701 source.n535 a_n1760_n3288# 0.016103f
C702 source.n536 a_n1760_n3288# 0.017051f
C703 source.n537 a_n1760_n3288# 0.038062f
C704 source.n538 a_n1760_n3288# 0.038062f
C705 source.n539 a_n1760_n3288# 0.017051f
C706 source.n540 a_n1760_n3288# 0.016103f
C707 source.n541 a_n1760_n3288# 0.029968f
C708 source.n542 a_n1760_n3288# 0.029968f
C709 source.n543 a_n1760_n3288# 0.016103f
C710 source.n544 a_n1760_n3288# 0.017051f
C711 source.n545 a_n1760_n3288# 0.038062f
C712 source.n546 a_n1760_n3288# 0.078108f
C713 source.n547 a_n1760_n3288# 0.017051f
C714 source.n548 a_n1760_n3288# 0.016103f
C715 source.n549 a_n1760_n3288# 0.064356f
C716 source.n550 a_n1760_n3288# 0.043107f
C717 source.n551 a_n1760_n3288# 0.282312f
C718 source.n552 a_n1760_n3288# 1.87766f
C719 plus.n0 a_n1760_n3288# 0.05331f
C720 plus.t7 a_n1760_n3288# 0.451937f
C721 plus.t14 a_n1760_n3288# 0.451937f
C722 plus.t8 a_n1760_n3288# 0.451937f
C723 plus.n1 a_n1760_n3288# 0.18202f
C724 plus.n2 a_n1760_n3288# 0.05331f
C725 plus.t0 a_n1760_n3288# 0.451937f
C726 plus.t9 a_n1760_n3288# 0.451937f
C727 plus.n3 a_n1760_n3288# 0.18202f
C728 plus.t4 a_n1760_n3288# 0.457594f
C729 plus.n4 a_n1760_n3288# 0.197737f
C730 plus.t1 a_n1760_n3288# 0.451937f
C731 plus.n5 a_n1760_n3288# 0.18202f
C732 plus.n6 a_n1760_n3288# 0.020314f
C733 plus.n7 a_n1760_n3288# 0.116735f
C734 plus.n8 a_n1760_n3288# 0.05331f
C735 plus.n9 a_n1760_n3288# 0.020314f
C736 plus.n10 a_n1760_n3288# 0.18202f
C737 plus.n11 a_n1760_n3288# 0.019f
C738 plus.n12 a_n1760_n3288# 0.019f
C739 plus.n13 a_n1760_n3288# 0.05331f
C740 plus.n14 a_n1760_n3288# 0.05331f
C741 plus.n15 a_n1760_n3288# 0.020314f
C742 plus.n16 a_n1760_n3288# 0.18202f
C743 plus.n17 a_n1760_n3288# 0.020314f
C744 plus.n18 a_n1760_n3288# 0.18202f
C745 plus.t2 a_n1760_n3288# 0.457594f
C746 plus.n19 a_n1760_n3288# 0.197663f
C747 plus.n20 a_n1760_n3288# 0.592177f
C748 plus.n21 a_n1760_n3288# 0.05331f
C749 plus.t5 a_n1760_n3288# 0.457594f
C750 plus.t10 a_n1760_n3288# 0.451937f
C751 plus.t12 a_n1760_n3288# 0.451937f
C752 plus.t3 a_n1760_n3288# 0.451937f
C753 plus.n22 a_n1760_n3288# 0.18202f
C754 plus.n23 a_n1760_n3288# 0.05331f
C755 plus.t15 a_n1760_n3288# 0.451937f
C756 plus.t6 a_n1760_n3288# 0.451937f
C757 plus.n24 a_n1760_n3288# 0.18202f
C758 plus.t13 a_n1760_n3288# 0.457594f
C759 plus.n25 a_n1760_n3288# 0.197737f
C760 plus.t11 a_n1760_n3288# 0.451937f
C761 plus.n26 a_n1760_n3288# 0.18202f
C762 plus.n27 a_n1760_n3288# 0.020314f
C763 plus.n28 a_n1760_n3288# 0.116735f
C764 plus.n29 a_n1760_n3288# 0.05331f
C765 plus.n30 a_n1760_n3288# 0.020314f
C766 plus.n31 a_n1760_n3288# 0.18202f
C767 plus.n32 a_n1760_n3288# 0.019f
C768 plus.n33 a_n1760_n3288# 0.019f
C769 plus.n34 a_n1760_n3288# 0.05331f
C770 plus.n35 a_n1760_n3288# 0.05331f
C771 plus.n36 a_n1760_n3288# 0.020314f
C772 plus.n37 a_n1760_n3288# 0.18202f
C773 plus.n38 a_n1760_n3288# 0.020314f
C774 plus.n39 a_n1760_n3288# 0.18202f
C775 plus.n40 a_n1760_n3288# 0.197663f
C776 plus.n41 a_n1760_n3288# 1.56001f
.ends

