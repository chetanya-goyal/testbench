* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t19 minus.t0 drain_right.t4 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 drain_right.t9 minus.t1 source.t18 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 source.t6 plus.t0 drain_left.t9 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X3 source.t17 minus.t2 drain_right.t8 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X5 a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X6 drain_left.t8 plus.t1 source.t9 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X7 source.t16 minus.t3 drain_right.t3 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X8 drain_right.t1 minus.t4 source.t15 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X9 drain_right.t0 minus.t5 source.t14 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X10 drain_right.t2 minus.t6 source.t13 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X11 drain_left.t7 plus.t2 source.t7 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X12 a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X13 source.t12 minus.t7 drain_right.t6 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X14 drain_right.t7 minus.t8 source.t11 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X15 drain_left.t6 plus.t3 source.t8 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X16 drain_right.t5 minus.t9 source.t10 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X17 source.t5 plus.t4 drain_left.t5 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X18 source.t0 plus.t5 drain_left.t4 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X19 drain_left.t3 plus.t6 source.t4 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X20 source.t1 plus.t7 drain_left.t2 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X21 drain_left.t1 plus.t8 source.t2 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X22 drain_left.t0 plus.t9 source.t3 a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X23 a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# a_n1496_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
R0 minus.n9 minus.t5 413.353
R1 minus.n3 minus.t4 413.353
R2 minus.n20 minus.t6 413.353
R3 minus.n14 minus.t8 413.353
R4 minus.n6 minus.t9 369.534
R5 minus.n8 minus.t7 369.534
R6 minus.n2 minus.t3 369.534
R7 minus.n17 minus.t1 369.534
R8 minus.n19 minus.t0 369.534
R9 minus.n13 minus.t2 369.534
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 26.4683
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t7 270.692
R42 drain_right.n7 drain_right.t0 270.132
R43 drain_right.n6 drain_right.n4 240.694
R44 drain_right.n3 drain_right.n2 240.496
R45 drain_right.n6 drain_right.n5 240.132
R46 drain_right.n1 drain_right.n0 240.131
R47 drain_right.n2 drain_right.t4 30.0005
R48 drain_right.n2 drain_right.t2 30.0005
R49 drain_right.n0 drain_right.t8 30.0005
R50 drain_right.n0 drain_right.t9 30.0005
R51 drain_right.n4 drain_right.t3 30.0005
R52 drain_right.n4 drain_right.t1 30.0005
R53 drain_right.n5 drain_right.t6 30.0005
R54 drain_right.n5 drain_right.t5 30.0005
R55 drain_right drain_right.n3 20.862
R56 drain_right drain_right.n7 5.93339
R57 drain_right.n7 drain_right.n6 0.560845
R58 drain_right.n3 drain_right.n1 0.0852402
R59 source.n0 source.t3 253.454
R60 source.n5 source.t15 253.454
R61 source.n19 source.t13 253.453
R62 source.n14 source.t9 253.453
R63 source.n2 source.n1 223.454
R64 source.n4 source.n3 223.454
R65 source.n7 source.n6 223.454
R66 source.n9 source.n8 223.454
R67 source.n18 source.n17 223.453
R68 source.n16 source.n15 223.453
R69 source.n13 source.n12 223.453
R70 source.n11 source.n10 223.453
R71 source.n17 source.t18 30.0005
R72 source.n17 source.t19 30.0005
R73 source.n15 source.t11 30.0005
R74 source.n15 source.t17 30.0005
R75 source.n12 source.t2 30.0005
R76 source.n12 source.t6 30.0005
R77 source.n10 source.t7 30.0005
R78 source.n10 source.t5 30.0005
R79 source.n1 source.t4 30.0005
R80 source.n1 source.t0 30.0005
R81 source.n3 source.t8 30.0005
R82 source.n3 source.t1 30.0005
R83 source.n6 source.t10 30.0005
R84 source.n6 source.t16 30.0005
R85 source.n8 source.t14 30.0005
R86 source.n8 source.t12 30.0005
R87 source.n11 source.n9 14.0751
R88 source.n20 source.n0 7.97163
R89 source.n20 source.n19 5.5436
R90 source.n5 source.n4 0.7505
R91 source.n16 source.n14 0.7505
R92 source.n9 source.n7 0.560845
R93 source.n7 source.n5 0.560845
R94 source.n4 source.n2 0.560845
R95 source.n2 source.n0 0.560845
R96 source.n13 source.n11 0.560845
R97 source.n14 source.n13 0.560845
R98 source.n18 source.n16 0.560845
R99 source.n19 source.n18 0.560845
R100 source source.n20 0.188
R101 plus.n3 plus.t3 413.353
R102 plus.n9 plus.t9 413.353
R103 plus.n14 plus.t1 413.353
R104 plus.n20 plus.t2 413.353
R105 plus.n6 plus.t6 369.534
R106 plus.n2 plus.t7 369.534
R107 plus.n8 plus.t5 369.534
R108 plus.n17 plus.t8 369.534
R109 plus.n13 plus.t0 369.534
R110 plus.n19 plus.t4 369.534
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 24.5161
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 7.99103
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t6 270.693
R142 drain_left.n1 drain_left.t7 270.692
R143 drain_left.n3 drain_left.n2 240.496
R144 drain_left.n7 drain_left.n6 240.132
R145 drain_left.n5 drain_left.n4 240.132
R146 drain_left.n1 drain_left.n0 240.131
R147 drain_left.n2 drain_left.t9 30.0005
R148 drain_left.n2 drain_left.t8 30.0005
R149 drain_left.n0 drain_left.t5 30.0005
R150 drain_left.n0 drain_left.t1 30.0005
R151 drain_left.n6 drain_left.t4 30.0005
R152 drain_left.n6 drain_left.t0 30.0005
R153 drain_left.n4 drain_left.t2 30.0005
R154 drain_left.n4 drain_left.t3 30.0005
R155 drain_left drain_left.n3 21.4152
R156 drain_left drain_left.n7 6.21356
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 minus drain_left 0.17838f
C1 drain_right drain_left 0.732337f
C2 source minus 0.706589f
C3 drain_right source 3.7799f
C4 plus drain_left 0.698885f
C5 drain_right minus 0.556194f
C6 source plus 0.720507f
C7 plus minus 2.97595f
C8 drain_right plus 0.305269f
C9 source drain_left 3.78189f
C10 drain_right a_n1496_n1088# 3.189083f
C11 drain_left a_n1496_n1088# 3.39626f
C12 source a_n1496_n1088# 2.099247f
C13 minus a_n1496_n1088# 4.610388f
C14 plus a_n1496_n1088# 5.408668f
C15 drain_left.t7 a_n1496_n1088# 0.1195f
C16 drain_left.t5 a_n1496_n1088# 0.02591f
C17 drain_left.t1 a_n1496_n1088# 0.02591f
C18 drain_left.n0 a_n1496_n1088# 0.084065f
C19 drain_left.n1 a_n1496_n1088# 0.412545f
C20 drain_left.t9 a_n1496_n1088# 0.02591f
C21 drain_left.t8 a_n1496_n1088# 0.02591f
C22 drain_left.n2 a_n1496_n1088# 0.084408f
C23 drain_left.n3 a_n1496_n1088# 0.732835f
C24 drain_left.t6 a_n1496_n1088# 0.119501f
C25 drain_left.t2 a_n1496_n1088# 0.02591f
C26 drain_left.t3 a_n1496_n1088# 0.02591f
C27 drain_left.n4 a_n1496_n1088# 0.084065f
C28 drain_left.n5 a_n1496_n1088# 0.439788f
C29 drain_left.t4 a_n1496_n1088# 0.02591f
C30 drain_left.t0 a_n1496_n1088# 0.02591f
C31 drain_left.n6 a_n1496_n1088# 0.084065f
C32 drain_left.n7 a_n1496_n1088# 0.410184f
C33 plus.n0 a_n1496_n1088# 0.04f
C34 plus.t5 a_n1496_n1088# 0.018497f
C35 plus.t6 a_n1496_n1088# 0.018497f
C36 plus.n1 a_n1496_n1088# 0.016969f
C37 plus.t3 a_n1496_n1088# 0.021039f
C38 plus.t7 a_n1496_n1088# 0.018497f
C39 plus.n2 a_n1496_n1088# 0.025223f
C40 plus.n3 a_n1496_n1088# 0.038469f
C41 plus.n4 a_n1496_n1088# 0.086112f
C42 plus.n5 a_n1496_n1088# 0.04f
C43 plus.n6 a_n1496_n1088# 0.038492f
C44 plus.n7 a_n1496_n1088# 0.016969f
C45 plus.n8 a_n1496_n1088# 0.025223f
C46 plus.t9 a_n1496_n1088# 0.021039f
C47 plus.n9 a_n1496_n1088# 0.038415f
C48 plus.n10 a_n1496_n1088# 0.275608f
C49 plus.n11 a_n1496_n1088# 0.04f
C50 plus.t2 a_n1496_n1088# 0.021039f
C51 plus.t4 a_n1496_n1088# 0.018497f
C52 plus.t8 a_n1496_n1088# 0.018497f
C53 plus.n12 a_n1496_n1088# 0.016969f
C54 plus.t0 a_n1496_n1088# 0.018497f
C55 plus.n13 a_n1496_n1088# 0.025223f
C56 plus.t1 a_n1496_n1088# 0.021039f
C57 plus.n14 a_n1496_n1088# 0.038469f
C58 plus.n15 a_n1496_n1088# 0.086112f
C59 plus.n16 a_n1496_n1088# 0.04f
C60 plus.n17 a_n1496_n1088# 0.038492f
C61 plus.n18 a_n1496_n1088# 0.016969f
C62 plus.n19 a_n1496_n1088# 0.025223f
C63 plus.n20 a_n1496_n1088# 0.038415f
C64 plus.n21 a_n1496_n1088# 0.813404f
C65 source.t3 a_n1496_n1088# 0.145851f
C66 source.n0 a_n1496_n1088# 0.557315f
C67 source.t4 a_n1496_n1088# 0.034793f
C68 source.t0 a_n1496_n1088# 0.034793f
C69 source.n1 a_n1496_n1088# 0.098134f
C70 source.n2 a_n1496_n1088# 0.283408f
C71 source.t8 a_n1496_n1088# 0.034793f
C72 source.t1 a_n1496_n1088# 0.034793f
C73 source.n3 a_n1496_n1088# 0.098134f
C74 source.n4 a_n1496_n1088# 0.301167f
C75 source.t15 a_n1496_n1088# 0.145851f
C76 source.n5 a_n1496_n1088# 0.316077f
C77 source.t10 a_n1496_n1088# 0.034793f
C78 source.t16 a_n1496_n1088# 0.034793f
C79 source.n6 a_n1496_n1088# 0.098134f
C80 source.n7 a_n1496_n1088# 0.283408f
C81 source.t14 a_n1496_n1088# 0.034793f
C82 source.t12 a_n1496_n1088# 0.034793f
C83 source.n8 a_n1496_n1088# 0.098134f
C84 source.n9 a_n1496_n1088# 0.828061f
C85 source.t7 a_n1496_n1088# 0.034793f
C86 source.t5 a_n1496_n1088# 0.034793f
C87 source.n10 a_n1496_n1088# 0.098133f
C88 source.n11 a_n1496_n1088# 0.828061f
C89 source.t2 a_n1496_n1088# 0.034793f
C90 source.t6 a_n1496_n1088# 0.034793f
C91 source.n12 a_n1496_n1088# 0.098133f
C92 source.n13 a_n1496_n1088# 0.283408f
C93 source.t9 a_n1496_n1088# 0.145851f
C94 source.n14 a_n1496_n1088# 0.316077f
C95 source.t11 a_n1496_n1088# 0.034793f
C96 source.t17 a_n1496_n1088# 0.034793f
C97 source.n15 a_n1496_n1088# 0.098133f
C98 source.n16 a_n1496_n1088# 0.301167f
C99 source.t18 a_n1496_n1088# 0.034793f
C100 source.t19 a_n1496_n1088# 0.034793f
C101 source.n17 a_n1496_n1088# 0.098133f
C102 source.n18 a_n1496_n1088# 0.283408f
C103 source.t13 a_n1496_n1088# 0.145851f
C104 source.n19 a_n1496_n1088# 0.455172f
C105 source.n20 a_n1496_n1088# 0.589189f
C106 drain_right.t7 a_n1496_n1088# 0.122223f
C107 drain_right.t8 a_n1496_n1088# 0.0265f
C108 drain_right.t9 a_n1496_n1088# 0.0265f
C109 drain_right.n0 a_n1496_n1088# 0.08598f
C110 drain_right.n1 a_n1496_n1088# 0.421945f
C111 drain_right.t4 a_n1496_n1088# 0.0265f
C112 drain_right.t2 a_n1496_n1088# 0.0265f
C113 drain_right.n2 a_n1496_n1088# 0.086331f
C114 drain_right.n3 a_n1496_n1088# 0.706655f
C115 drain_right.t3 a_n1496_n1088# 0.0265f
C116 drain_right.t1 a_n1496_n1088# 0.0265f
C117 drain_right.n4 a_n1496_n1088# 0.086548f
C118 drain_right.t6 a_n1496_n1088# 0.0265f
C119 drain_right.t5 a_n1496_n1088# 0.0265f
C120 drain_right.n5 a_n1496_n1088# 0.08598f
C121 drain_right.n6 a_n1496_n1088# 0.477746f
C122 drain_right.t0 a_n1496_n1088# 0.121777f
C123 drain_right.n7 a_n1496_n1088# 0.401143f
C124 minus.n0 a_n1496_n1088# 0.03895f
C125 minus.t5 a_n1496_n1088# 0.020487f
C126 minus.t7 a_n1496_n1088# 0.018011f
C127 minus.t9 a_n1496_n1088# 0.018011f
C128 minus.n1 a_n1496_n1088# 0.016523f
C129 minus.t3 a_n1496_n1088# 0.018011f
C130 minus.n2 a_n1496_n1088# 0.02456f
C131 minus.t4 a_n1496_n1088# 0.020487f
C132 minus.n3 a_n1496_n1088# 0.037459f
C133 minus.n4 a_n1496_n1088# 0.083851f
C134 minus.n5 a_n1496_n1088# 0.03895f
C135 minus.n6 a_n1496_n1088# 0.037481f
C136 minus.n7 a_n1496_n1088# 0.016523f
C137 minus.n8 a_n1496_n1088# 0.02456f
C138 minus.n9 a_n1496_n1088# 0.037406f
C139 minus.n10 a_n1496_n1088# 0.812837f
C140 minus.n11 a_n1496_n1088# 0.03895f
C141 minus.t0 a_n1496_n1088# 0.018011f
C142 minus.t1 a_n1496_n1088# 0.018011f
C143 minus.n12 a_n1496_n1088# 0.016523f
C144 minus.t8 a_n1496_n1088# 0.020487f
C145 minus.t2 a_n1496_n1088# 0.018011f
C146 minus.n13 a_n1496_n1088# 0.02456f
C147 minus.n14 a_n1496_n1088# 0.037459f
C148 minus.n15 a_n1496_n1088# 0.083851f
C149 minus.n16 a_n1496_n1088# 0.03895f
C150 minus.n17 a_n1496_n1088# 0.037481f
C151 minus.n18 a_n1496_n1088# 0.016523f
C152 minus.n19 a_n1496_n1088# 0.02456f
C153 minus.t6 a_n1496_n1088# 0.020487f
C154 minus.n20 a_n1496_n1088# 0.037406f
C155 minus.n21 a_n1496_n1088# 0.255908f
C156 minus.n22 a_n1496_n1088# 1.00313f
.ends

