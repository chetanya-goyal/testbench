* NGSPICE file created from diffpair583.ext - technology: sky130A

.subckt diffpair583 minus drain_right drain_left source plus
X0 a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X1 drain_left.t7 plus.t0 source.t4 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X2 drain_left.t6 plus.t1 source.t3 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X3 drain_left.t5 plus.t2 source.t8 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X4 source.t11 minus.t0 drain_right.t7 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X5 source.t12 minus.t1 drain_right.t6 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X6 source.t13 minus.t2 drain_right.t5 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X7 source.t5 plus.t3 drain_left.t4 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X8 source.t7 plus.t4 drain_left.t3 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X9 a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X10 drain_right.t4 minus.t3 source.t14 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X11 a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X12 a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X13 source.t6 plus.t5 drain_left.t2 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X14 drain_left.t1 plus.t6 source.t9 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X15 drain_right.t3 minus.t4 source.t0 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X16 drain_right.t2 minus.t5 source.t15 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X17 drain_right.t1 minus.t6 source.t1 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X18 source.t10 plus.t7 drain_left.t0 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X19 source.t2 minus.t7 drain_right.t0 a_n1296_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
R0 plus.n1 plus.t4 2107.36
R1 plus.n5 plus.t0 2107.36
R2 plus.n8 plus.t2 2107.36
R3 plus.n12 plus.t3 2107.36
R4 plus.n2 plus.t1 2053.32
R5 plus.n4 plus.t5 2053.32
R6 plus.n9 plus.t7 2053.32
R7 plus.n11 plus.t6 2053.32
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus plus.n13 30.9422
R19 plus.n2 plus.n1 30.6732
R20 plus.n5 plus.n4 30.6732
R21 plus.n12 plus.n11 30.6732
R22 plus.n9 plus.n8 30.6732
R23 plus plus.n6 15.1747
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n0 source.t4 44.1297
R27 source.n3 source.t7 44.1296
R28 source.n4 source.t15 44.1296
R29 source.n7 source.t11 44.1296
R30 source.n15 source.t1 44.1295
R31 source.n12 source.t12 44.1295
R32 source.n11 source.t8 44.1295
R33 source.n8 source.t5 44.1295
R34 source.n2 source.n1 43.1397
R35 source.n6 source.n5 43.1397
R36 source.n14 source.n13 43.1396
R37 source.n10 source.n9 43.1396
R38 source.n8 source.n7 27.8483
R39 source.n16 source.n0 22.3354
R40 source.n16 source.n15 5.51343
R41 source.n13 source.t14 0.9905
R42 source.n13 source.t2 0.9905
R43 source.n9 source.t9 0.9905
R44 source.n9 source.t10 0.9905
R45 source.n1 source.t3 0.9905
R46 source.n1 source.t6 0.9905
R47 source.n5 source.t0 0.9905
R48 source.n5 source.t13 0.9905
R49 source.n7 source.n6 0.5005
R50 source.n6 source.n4 0.5005
R51 source.n3 source.n2 0.5005
R52 source.n2 source.n0 0.5005
R53 source.n10 source.n8 0.5005
R54 source.n11 source.n10 0.5005
R55 source.n14 source.n12 0.5005
R56 source.n15 source.n14 0.5005
R57 source.n4 source.n3 0.470328
R58 source.n12 source.n11 0.470328
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 60.3185
R61 drain_left.n2 drain_left.n1 60.0131
R62 drain_left.n2 drain_left.n0 60.0131
R63 drain_left.n5 drain_left.n4 59.8185
R64 drain_left drain_left.n2 35.1777
R65 drain_left drain_left.n5 6.15322
R66 drain_left.n1 drain_left.t0 0.9905
R67 drain_left.n1 drain_left.t5 0.9905
R68 drain_left.n0 drain_left.t4 0.9905
R69 drain_left.n0 drain_left.t1 0.9905
R70 drain_left.n4 drain_left.t2 0.9905
R71 drain_left.n4 drain_left.t7 0.9905
R72 drain_left.n3 drain_left.t3 0.9905
R73 drain_left.n3 drain_left.t6 0.9905
R74 minus.n5 minus.t0 2107.36
R75 minus.n1 minus.t5 2107.36
R76 minus.n12 minus.t6 2107.36
R77 minus.n8 minus.t1 2107.36
R78 minus.n4 minus.t4 2053.32
R79 minus.n2 minus.t2 2053.32
R80 minus.n11 minus.t7 2053.32
R81 minus.n9 minus.t3 2053.32
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 42.3581
R89 minus.n3 minus.n2 42.3581
R90 minus.n10 minus.n9 42.3581
R91 minus.n11 minus.n10 42.3581
R92 minus.n14 minus.n6 40.0914
R93 minus.n5 minus.n4 30.6732
R94 minus.n2 minus.n1 30.6732
R95 minus.n9 minus.n8 30.6732
R96 minus.n12 minus.n11 30.6732
R97 minus.n14 minus.n13 6.5005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 60.3185
R102 drain_right.n2 drain_right.n1 60.0131
R103 drain_right.n2 drain_right.n0 60.0131
R104 drain_right.n5 drain_right.n4 59.8185
R105 drain_right drain_right.n2 34.6245
R106 drain_right drain_right.n5 6.15322
R107 drain_right.n1 drain_right.t0 0.9905
R108 drain_right.n1 drain_right.t1 0.9905
R109 drain_right.n0 drain_right.t6 0.9905
R110 drain_right.n0 drain_right.t4 0.9905
R111 drain_right.n3 drain_right.t5 0.9905
R112 drain_right.n3 drain_right.t2 0.9905
R113 drain_right.n4 drain_right.t7 0.9905
R114 drain_right.n4 drain_right.t3 0.9905
C0 source minus 3.96744f
C1 minus plus 6.24761f
C2 drain_right drain_left 0.605638f
C3 drain_right source 28.695501f
C4 drain_right plus 0.275273f
C5 drain_right minus 4.77533f
C6 source drain_left 28.696598f
C7 drain_left plus 4.89733f
C8 drain_left minus 0.170438f
C9 source plus 3.98148f
C10 drain_right a_n1296_n4888# 7.650031f
C11 drain_left a_n1296_n4888# 7.8456f
C12 source a_n1296_n4888# 12.798121f
C13 minus a_n1296_n4888# 5.518497f
C14 plus a_n1296_n4888# 8.184f
C15 drain_right.t6 a_n1296_n4888# 0.562431f
C16 drain_right.t4 a_n1296_n4888# 0.562431f
C17 drain_right.n0 a_n1296_n4888# 5.14316f
C18 drain_right.t0 a_n1296_n4888# 0.562431f
C19 drain_right.t1 a_n1296_n4888# 0.562431f
C20 drain_right.n1 a_n1296_n4888# 5.14316f
C21 drain_right.n2 a_n1296_n4888# 2.95416f
C22 drain_right.t5 a_n1296_n4888# 0.562431f
C23 drain_right.t2 a_n1296_n4888# 0.562431f
C24 drain_right.n3 a_n1296_n4888# 5.14542f
C25 drain_right.t7 a_n1296_n4888# 0.562431f
C26 drain_right.t3 a_n1296_n4888# 0.562431f
C27 drain_right.n4 a_n1296_n4888# 5.14186f
C28 drain_right.n5 a_n1296_n4888# 1.13447f
C29 minus.n0 a_n1296_n4888# 0.132592f
C30 minus.t0 a_n1296_n4888# 0.819547f
C31 minus.t4 a_n1296_n4888# 0.81163f
C32 minus.t2 a_n1296_n4888# 0.81163f
C33 minus.t5 a_n1296_n4888# 0.819547f
C34 minus.n1 a_n1296_n4888# 0.322859f
C35 minus.n2 a_n1296_n4888# 0.304462f
C36 minus.n3 a_n1296_n4888# 0.021962f
C37 minus.n4 a_n1296_n4888# 0.304462f
C38 minus.n5 a_n1296_n4888# 0.322771f
C39 minus.n6 a_n1296_n4888# 2.38204f
C40 minus.n7 a_n1296_n4888# 0.132592f
C41 minus.t7 a_n1296_n4888# 0.81163f
C42 minus.t3 a_n1296_n4888# 0.81163f
C43 minus.t1 a_n1296_n4888# 0.819547f
C44 minus.n8 a_n1296_n4888# 0.322859f
C45 minus.n9 a_n1296_n4888# 0.304462f
C46 minus.n10 a_n1296_n4888# 0.021962f
C47 minus.n11 a_n1296_n4888# 0.304462f
C48 minus.t6 a_n1296_n4888# 0.819547f
C49 minus.n12 a_n1296_n4888# 0.322771f
C50 minus.n13 a_n1296_n4888# 0.376866f
C51 minus.n14 a_n1296_n4888# 2.86032f
C52 drain_left.t4 a_n1296_n4888# 0.561775f
C53 drain_left.t1 a_n1296_n4888# 0.561775f
C54 drain_left.n0 a_n1296_n4888# 5.13716f
C55 drain_left.t0 a_n1296_n4888# 0.561775f
C56 drain_left.t5 a_n1296_n4888# 0.561775f
C57 drain_left.n1 a_n1296_n4888# 5.13716f
C58 drain_left.n2 a_n1296_n4888# 3.02534f
C59 drain_left.t3 a_n1296_n4888# 0.561775f
C60 drain_left.t6 a_n1296_n4888# 0.561775f
C61 drain_left.n3 a_n1296_n4888# 5.13942f
C62 drain_left.t2 a_n1296_n4888# 0.561775f
C63 drain_left.t7 a_n1296_n4888# 0.561775f
C64 drain_left.n4 a_n1296_n4888# 5.13586f
C65 drain_left.n5 a_n1296_n4888# 1.13314f
C66 source.t4 a_n1296_n4888# 4.47661f
C67 source.n0 a_n1296_n4888# 1.89863f
C68 source.t3 a_n1296_n4888# 0.39171f
C69 source.t6 a_n1296_n4888# 0.39171f
C70 source.n1 a_n1296_n4888# 3.50206f
C71 source.n2 a_n1296_n4888# 0.334365f
C72 source.t7 a_n1296_n4888# 4.47662f
C73 source.n3 a_n1296_n4888# 0.42569f
C74 source.t15 a_n1296_n4888# 4.47662f
C75 source.n4 a_n1296_n4888# 0.42569f
C76 source.t0 a_n1296_n4888# 0.39171f
C77 source.t13 a_n1296_n4888# 0.39171f
C78 source.n5 a_n1296_n4888# 3.50206f
C79 source.n6 a_n1296_n4888# 0.334365f
C80 source.t11 a_n1296_n4888# 4.47662f
C81 source.n7 a_n1296_n4888# 2.33638f
C82 source.t5 a_n1296_n4888# 4.4766f
C83 source.n8 a_n1296_n4888# 2.33641f
C84 source.t9 a_n1296_n4888# 0.39171f
C85 source.t10 a_n1296_n4888# 0.39171f
C86 source.n9 a_n1296_n4888# 3.50206f
C87 source.n10 a_n1296_n4888# 0.334358f
C88 source.t8 a_n1296_n4888# 4.4766f
C89 source.n11 a_n1296_n4888# 0.425715f
C90 source.t12 a_n1296_n4888# 4.4766f
C91 source.n12 a_n1296_n4888# 0.425715f
C92 source.t14 a_n1296_n4888# 0.39171f
C93 source.t2 a_n1296_n4888# 0.39171f
C94 source.n13 a_n1296_n4888# 3.50206f
C95 source.n14 a_n1296_n4888# 0.334358f
C96 source.t1 a_n1296_n4888# 4.4766f
C97 source.n15 a_n1296_n4888# 0.562868f
C98 source.n16 a_n1296_n4888# 2.22893f
C99 plus.n0 a_n1296_n4888# 0.134522f
C100 plus.t5 a_n1296_n4888# 0.823439f
C101 plus.t1 a_n1296_n4888# 0.823439f
C102 plus.t4 a_n1296_n4888# 0.831471f
C103 plus.n1 a_n1296_n4888# 0.327557f
C104 plus.n2 a_n1296_n4888# 0.308892f
C105 plus.n3 a_n1296_n4888# 0.022281f
C106 plus.n4 a_n1296_n4888# 0.308892f
C107 plus.t0 a_n1296_n4888# 0.831471f
C108 plus.n5 a_n1296_n4888# 0.327467f
C109 plus.n6 a_n1296_n4888# 0.887939f
C110 plus.n7 a_n1296_n4888# 0.134522f
C111 plus.t3 a_n1296_n4888# 0.831471f
C112 plus.t6 a_n1296_n4888# 0.823439f
C113 plus.t7 a_n1296_n4888# 0.823439f
C114 plus.t2 a_n1296_n4888# 0.831471f
C115 plus.n8 a_n1296_n4888# 0.327557f
C116 plus.n9 a_n1296_n4888# 0.308892f
C117 plus.n10 a_n1296_n4888# 0.022281f
C118 plus.n11 a_n1296_n4888# 0.308892f
C119 plus.n12 a_n1296_n4888# 0.327467f
C120 plus.n13 a_n1296_n4888# 1.89681f
.ends

