* NGSPICE file created from diffpair224.ext - technology: sky130A

.subckt diffpair224 minus drain_right drain_left source plus
X0 source.t17 minus.t0 drain_right.t5 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 drain_right.t0 minus.t1 source.t16 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 drain_left.t9 plus.t0 source.t1 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X3 source.t15 minus.t2 drain_right.t1 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X4 a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X5 drain_left.t8 plus.t1 source.t18 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X6 drain_left.t7 plus.t2 source.t5 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X7 source.t14 minus.t3 drain_right.t8 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X8 drain_right.t6 minus.t4 source.t13 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X9 drain_right.t2 minus.t5 source.t12 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X10 drain_left.t6 plus.t3 source.t0 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X11 source.t19 plus.t4 drain_left.t5 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X12 a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X13 drain_right.t4 minus.t6 source.t11 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X14 a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X15 drain_left.t4 plus.t5 source.t2 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 drain_right.t9 minus.t7 source.t10 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X17 source.t3 plus.t6 drain_left.t3 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X18 drain_right.t3 minus.t8 source.t9 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X19 source.t7 plus.t7 drain_left.t2 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X20 a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X21 drain_left.t1 plus.t8 source.t4 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X22 source.t6 plus.t9 drain_left.t0 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 source.t8 minus.t9 drain_right.t7 a_n1952_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n3 minus.t8 182.153
R1 minus.n17 minus.t1 182.153
R2 minus.n13 minus.n12 161.3
R3 minus.n11 minus.n0 161.3
R4 minus.n10 minus.n9 161.3
R5 minus.n8 minus.n1 161.3
R6 minus.n7 minus.n6 161.3
R7 minus.n5 minus.n2 161.3
R8 minus.n27 minus.n26 161.3
R9 minus.n25 minus.n14 161.3
R10 minus.n24 minus.n23 161.3
R11 minus.n22 minus.n15 161.3
R12 minus.n21 minus.n20 161.3
R13 minus.n19 minus.n16 161.3
R14 minus.n4 minus.t2 159.405
R15 minus.n6 minus.t7 159.405
R16 minus.n10 minus.t9 159.405
R17 minus.n12 minus.t6 159.405
R18 minus.n18 minus.t0 159.405
R19 minus.n20 minus.t4 159.405
R20 minus.n24 minus.t3 159.405
R21 minus.n26 minus.t5 159.405
R22 minus.n3 minus.n2 44.8741
R23 minus.n17 minus.n16 44.8741
R24 minus.n12 minus.n11 30.6732
R25 minus.n26 minus.n25 30.6732
R26 minus.n28 minus.n13 29.8357
R27 minus.n5 minus.n4 26.2914
R28 minus.n10 minus.n1 26.2914
R29 minus.n19 minus.n18 26.2914
R30 minus.n24 minus.n15 26.2914
R31 minus.n6 minus.n5 21.9096
R32 minus.n6 minus.n1 21.9096
R33 minus.n20 minus.n19 21.9096
R34 minus.n20 minus.n15 21.9096
R35 minus.n4 minus.n3 19.0667
R36 minus.n18 minus.n17 19.0667
R37 minus.n11 minus.n10 17.5278
R38 minus.n25 minus.n24 17.5278
R39 minus.n28 minus.n27 6.63876
R40 minus.n13 minus.n0 0.189894
R41 minus.n9 minus.n0 0.189894
R42 minus.n9 minus.n8 0.189894
R43 minus.n8 minus.n7 0.189894
R44 minus.n7 minus.n2 0.189894
R45 minus.n21 minus.n16 0.189894
R46 minus.n22 minus.n21 0.189894
R47 minus.n23 minus.n22 0.189894
R48 minus.n23 minus.n14 0.189894
R49 minus.n27 minus.n14 0.189894
R50 minus minus.n28 0.188
R51 drain_right.n1 drain_right.t0 87.2609
R52 drain_right.n7 drain_right.t4 86.3731
R53 drain_right.n6 drain_right.n4 80.661
R54 drain_right.n3 drain_right.n2 80.3836
R55 drain_right.n6 drain_right.n5 79.7731
R56 drain_right.n1 drain_right.n0 79.773
R57 drain_right drain_right.n3 23.7694
R58 drain_right.n2 drain_right.t8 6.6005
R59 drain_right.n2 drain_right.t2 6.6005
R60 drain_right.n0 drain_right.t5 6.6005
R61 drain_right.n0 drain_right.t6 6.6005
R62 drain_right.n4 drain_right.t1 6.6005
R63 drain_right.n4 drain_right.t3 6.6005
R64 drain_right.n5 drain_right.t7 6.6005
R65 drain_right.n5 drain_right.t9 6.6005
R66 drain_right drain_right.n7 6.09718
R67 drain_right.n7 drain_right.n6 0.888431
R68 drain_right.n3 drain_right.n1 0.167137
R69 source.n0 source.t18 69.6943
R70 source.n5 source.t9 69.6943
R71 source.n19 source.t12 69.6942
R72 source.n14 source.t0 69.6942
R73 source.n2 source.n1 63.0943
R74 source.n4 source.n3 63.0943
R75 source.n7 source.n6 63.0943
R76 source.n9 source.n8 63.0943
R77 source.n18 source.n17 63.0942
R78 source.n16 source.n15 63.0942
R79 source.n13 source.n12 63.0942
R80 source.n11 source.n10 63.0942
R81 source.n11 source.n9 16.2454
R82 source.n20 source.n0 9.65058
R83 source.n17 source.t13 6.6005
R84 source.n17 source.t14 6.6005
R85 source.n15 source.t16 6.6005
R86 source.n15 source.t17 6.6005
R87 source.n12 source.t2 6.6005
R88 source.n12 source.t19 6.6005
R89 source.n10 source.t4 6.6005
R90 source.n10 source.t6 6.6005
R91 source.n1 source.t1 6.6005
R92 source.n1 source.t3 6.6005
R93 source.n3 source.t5 6.6005
R94 source.n3 source.t7 6.6005
R95 source.n6 source.t10 6.6005
R96 source.n6 source.t15 6.6005
R97 source.n8 source.t11 6.6005
R98 source.n8 source.t8 6.6005
R99 source.n20 source.n19 5.7074
R100 source.n5 source.n4 0.914293
R101 source.n16 source.n14 0.914293
R102 source.n9 source.n7 0.888431
R103 source.n7 source.n5 0.888431
R104 source.n4 source.n2 0.888431
R105 source.n2 source.n0 0.888431
R106 source.n13 source.n11 0.888431
R107 source.n14 source.n13 0.888431
R108 source.n18 source.n16 0.888431
R109 source.n19 source.n18 0.888431
R110 source source.n20 0.188
R111 plus.n3 plus.t2 182.153
R112 plus.n17 plus.t3 182.153
R113 plus.n6 plus.n5 161.3
R114 plus.n7 plus.n2 161.3
R115 plus.n9 plus.n8 161.3
R116 plus.n10 plus.n1 161.3
R117 plus.n11 plus.n0 161.3
R118 plus.n13 plus.n12 161.3
R119 plus.n20 plus.n19 161.3
R120 plus.n21 plus.n16 161.3
R121 plus.n23 plus.n22 161.3
R122 plus.n24 plus.n15 161.3
R123 plus.n25 plus.n14 161.3
R124 plus.n27 plus.n26 161.3
R125 plus.n12 plus.t1 159.405
R126 plus.n10 plus.t6 159.405
R127 plus.n2 plus.t0 159.405
R128 plus.n4 plus.t7 159.405
R129 plus.n26 plus.t8 159.405
R130 plus.n24 plus.t9 159.405
R131 plus.n16 plus.t5 159.405
R132 plus.n18 plus.t4 159.405
R133 plus.n6 plus.n3 44.8741
R134 plus.n20 plus.n17 44.8741
R135 plus.n12 plus.n11 30.6732
R136 plus.n26 plus.n25 30.6732
R137 plus plus.n27 27.1259
R138 plus.n10 plus.n9 26.2914
R139 plus.n5 plus.n4 26.2914
R140 plus.n24 plus.n23 26.2914
R141 plus.n19 plus.n18 26.2914
R142 plus.n9 plus.n2 21.9096
R143 plus.n5 plus.n2 21.9096
R144 plus.n23 plus.n16 21.9096
R145 plus.n19 plus.n16 21.9096
R146 plus.n4 plus.n3 19.0667
R147 plus.n18 plus.n17 19.0667
R148 plus.n11 plus.n10 17.5278
R149 plus.n25 plus.n24 17.5278
R150 plus plus.n13 8.87361
R151 plus.n7 plus.n6 0.189894
R152 plus.n8 plus.n7 0.189894
R153 plus.n8 plus.n1 0.189894
R154 plus.n1 plus.n0 0.189894
R155 plus.n13 plus.n0 0.189894
R156 plus.n27 plus.n14 0.189894
R157 plus.n15 plus.n14 0.189894
R158 plus.n22 plus.n15 0.189894
R159 plus.n22 plus.n21 0.189894
R160 plus.n21 plus.n20 0.189894
R161 drain_left.n5 drain_left.t7 87.261
R162 drain_left.n1 drain_left.t1 87.2609
R163 drain_left.n3 drain_left.n2 80.3836
R164 drain_left.n7 drain_left.n6 79.7731
R165 drain_left.n5 drain_left.n4 79.7731
R166 drain_left.n1 drain_left.n0 79.773
R167 drain_left drain_left.n3 24.3226
R168 drain_left.n2 drain_left.t5 6.6005
R169 drain_left.n2 drain_left.t6 6.6005
R170 drain_left.n0 drain_left.t0 6.6005
R171 drain_left.n0 drain_left.t4 6.6005
R172 drain_left.n6 drain_left.t3 6.6005
R173 drain_left.n6 drain_left.t8 6.6005
R174 drain_left.n4 drain_left.t2 6.6005
R175 drain_left.n4 drain_left.t9 6.6005
R176 drain_left drain_left.n7 6.54115
R177 drain_left.n7 drain_left.n5 0.888431
R178 drain_left.n3 drain_left.n1 0.167137
C0 source minus 2.30466f
C1 minus plus 3.91697f
C2 drain_left minus 0.177062f
C3 source plus 2.31878f
C4 source drain_left 5.5191f
C5 drain_left plus 2.2015f
C6 drain_right minus 2.01185f
C7 source drain_right 5.51828f
C8 drain_right plus 0.35148f
C9 drain_right drain_left 0.966289f
C10 drain_right a_n1952_n1488# 4.39814f
C11 drain_left a_n1952_n1488# 4.70891f
C12 source a_n1952_n1488# 3.020271f
C13 minus a_n1952_n1488# 6.907189f
C14 plus a_n1952_n1488# 8.15008f
C15 drain_left.t1 a_n1952_n1488# 0.544467f
C16 drain_left.t0 a_n1952_n1488# 0.058473f
C17 drain_left.t4 a_n1952_n1488# 0.058473f
C18 drain_left.n0 a_n1952_n1488# 0.421701f
C19 drain_left.n1 a_n1952_n1488# 0.599333f
C20 drain_left.t5 a_n1952_n1488# 0.058473f
C21 drain_left.t6 a_n1952_n1488# 0.058473f
C22 drain_left.n2 a_n1952_n1488# 0.424188f
C23 drain_left.n3 a_n1952_n1488# 1.11907f
C24 drain_left.t7 a_n1952_n1488# 0.544469f
C25 drain_left.t2 a_n1952_n1488# 0.058473f
C26 drain_left.t9 a_n1952_n1488# 0.058473f
C27 drain_left.n4 a_n1952_n1488# 0.421703f
C28 drain_left.n5 a_n1952_n1488# 0.653223f
C29 drain_left.t3 a_n1952_n1488# 0.058473f
C30 drain_left.t8 a_n1952_n1488# 0.058473f
C31 drain_left.n6 a_n1952_n1488# 0.421703f
C32 drain_left.n7 a_n1952_n1488# 0.556739f
C33 plus.n0 a_n1952_n1488# 0.046452f
C34 plus.t1 a_n1952_n1488# 0.292515f
C35 plus.t6 a_n1952_n1488# 0.292515f
C36 plus.n1 a_n1952_n1488# 0.046452f
C37 plus.t0 a_n1952_n1488# 0.292515f
C38 plus.n2 a_n1952_n1488# 0.170367f
C39 plus.t2 a_n1952_n1488# 0.313771f
C40 plus.n3 a_n1952_n1488# 0.153347f
C41 plus.t7 a_n1952_n1488# 0.292515f
C42 plus.n4 a_n1952_n1488# 0.175048f
C43 plus.n5 a_n1952_n1488# 0.010541f
C44 plus.n6 a_n1952_n1488# 0.19402f
C45 plus.n7 a_n1952_n1488# 0.046452f
C46 plus.n8 a_n1952_n1488# 0.046452f
C47 plus.n9 a_n1952_n1488# 0.010541f
C48 plus.n10 a_n1952_n1488# 0.170367f
C49 plus.n11 a_n1952_n1488# 0.010541f
C50 plus.n12 a_n1952_n1488# 0.16779f
C51 plus.n13 a_n1952_n1488# 0.362885f
C52 plus.n14 a_n1952_n1488# 0.046452f
C53 plus.t8 a_n1952_n1488# 0.292515f
C54 plus.n15 a_n1952_n1488# 0.046452f
C55 plus.t9 a_n1952_n1488# 0.292515f
C56 plus.t5 a_n1952_n1488# 0.292515f
C57 plus.n16 a_n1952_n1488# 0.170367f
C58 plus.t3 a_n1952_n1488# 0.313771f
C59 plus.n17 a_n1952_n1488# 0.153347f
C60 plus.t4 a_n1952_n1488# 0.292515f
C61 plus.n18 a_n1952_n1488# 0.175048f
C62 plus.n19 a_n1952_n1488# 0.010541f
C63 plus.n20 a_n1952_n1488# 0.19402f
C64 plus.n21 a_n1952_n1488# 0.046452f
C65 plus.n22 a_n1952_n1488# 0.046452f
C66 plus.n23 a_n1952_n1488# 0.010541f
C67 plus.n24 a_n1952_n1488# 0.170367f
C68 plus.n25 a_n1952_n1488# 0.010541f
C69 plus.n26 a_n1952_n1488# 0.16779f
C70 plus.n27 a_n1952_n1488# 1.13179f
C71 source.t18 a_n1952_n1488# 0.591871f
C72 source.n0 a_n1952_n1488# 0.86619f
C73 source.t1 a_n1952_n1488# 0.071277f
C74 source.t3 a_n1952_n1488# 0.071277f
C75 source.n1 a_n1952_n1488# 0.451937f
C76 source.n2 a_n1952_n1488# 0.433956f
C77 source.t5 a_n1952_n1488# 0.071277f
C78 source.t7 a_n1952_n1488# 0.071277f
C79 source.n3 a_n1952_n1488# 0.451937f
C80 source.n4 a_n1952_n1488# 0.436462f
C81 source.t9 a_n1952_n1488# 0.591871f
C82 source.n5 a_n1952_n1488# 0.490919f
C83 source.t10 a_n1952_n1488# 0.071277f
C84 source.t15 a_n1952_n1488# 0.071277f
C85 source.n6 a_n1952_n1488# 0.451937f
C86 source.n7 a_n1952_n1488# 0.433956f
C87 source.t11 a_n1952_n1488# 0.071277f
C88 source.t8 a_n1952_n1488# 0.071277f
C89 source.n8 a_n1952_n1488# 0.451937f
C90 source.n9 a_n1952_n1488# 1.21928f
C91 source.t4 a_n1952_n1488# 0.071277f
C92 source.t6 a_n1952_n1488# 0.071277f
C93 source.n10 a_n1952_n1488# 0.451933f
C94 source.n11 a_n1952_n1488# 1.21929f
C95 source.t2 a_n1952_n1488# 0.071277f
C96 source.t19 a_n1952_n1488# 0.071277f
C97 source.n12 a_n1952_n1488# 0.451933f
C98 source.n13 a_n1952_n1488# 0.43396f
C99 source.t0 a_n1952_n1488# 0.591868f
C100 source.n14 a_n1952_n1488# 0.490922f
C101 source.t16 a_n1952_n1488# 0.071277f
C102 source.t17 a_n1952_n1488# 0.071277f
C103 source.n15 a_n1952_n1488# 0.451933f
C104 source.n16 a_n1952_n1488# 0.436465f
C105 source.t13 a_n1952_n1488# 0.071277f
C106 source.t14 a_n1952_n1488# 0.071277f
C107 source.n17 a_n1952_n1488# 0.451933f
C108 source.n18 a_n1952_n1488# 0.43396f
C109 source.t12 a_n1952_n1488# 0.591868f
C110 source.n19 a_n1952_n1488# 0.644032f
C111 source.n20 a_n1952_n1488# 0.886605f
C112 drain_right.t0 a_n1952_n1488# 0.537054f
C113 drain_right.t5 a_n1952_n1488# 0.057677f
C114 drain_right.t6 a_n1952_n1488# 0.057677f
C115 drain_right.n0 a_n1952_n1488# 0.41596f
C116 drain_right.n1 a_n1952_n1488# 0.591174f
C117 drain_right.t8 a_n1952_n1488# 0.057677f
C118 drain_right.t2 a_n1952_n1488# 0.057677f
C119 drain_right.n2 a_n1952_n1488# 0.418414f
C120 drain_right.n3 a_n1952_n1488# 1.05568f
C121 drain_right.t1 a_n1952_n1488# 0.057677f
C122 drain_right.t3 a_n1952_n1488# 0.057677f
C123 drain_right.n4 a_n1952_n1488# 0.419747f
C124 drain_right.t7 a_n1952_n1488# 0.057677f
C125 drain_right.t9 a_n1952_n1488# 0.057677f
C126 drain_right.n5 a_n1952_n1488# 0.415962f
C127 drain_right.n6 a_n1952_n1488# 0.673948f
C128 drain_right.t4 a_n1952_n1488# 0.533866f
C129 drain_right.n7 a_n1952_n1488# 0.537154f
C130 minus.n0 a_n1952_n1488# 0.044844f
C131 minus.n1 a_n1952_n1488# 0.010176f
C132 minus.t9 a_n1952_n1488# 0.282392f
C133 minus.n2 a_n1952_n1488# 0.187306f
C134 minus.t8 a_n1952_n1488# 0.302912f
C135 minus.n3 a_n1952_n1488# 0.14804f
C136 minus.t2 a_n1952_n1488# 0.282392f
C137 minus.n4 a_n1952_n1488# 0.16899f
C138 minus.n5 a_n1952_n1488# 0.010176f
C139 minus.t7 a_n1952_n1488# 0.282392f
C140 minus.n6 a_n1952_n1488# 0.164472f
C141 minus.n7 a_n1952_n1488# 0.044844f
C142 minus.n8 a_n1952_n1488# 0.044844f
C143 minus.n9 a_n1952_n1488# 0.044844f
C144 minus.n10 a_n1952_n1488# 0.164472f
C145 minus.n11 a_n1952_n1488# 0.010176f
C146 minus.t6 a_n1952_n1488# 0.282392f
C147 minus.n12 a_n1952_n1488# 0.161983f
C148 minus.n13 a_n1952_n1488# 1.16151f
C149 minus.n14 a_n1952_n1488# 0.044844f
C150 minus.n15 a_n1952_n1488# 0.010176f
C151 minus.n16 a_n1952_n1488# 0.187306f
C152 minus.t1 a_n1952_n1488# 0.302912f
C153 minus.n17 a_n1952_n1488# 0.14804f
C154 minus.t0 a_n1952_n1488# 0.282392f
C155 minus.n18 a_n1952_n1488# 0.16899f
C156 minus.n19 a_n1952_n1488# 0.010176f
C157 minus.t4 a_n1952_n1488# 0.282392f
C158 minus.n20 a_n1952_n1488# 0.164472f
C159 minus.n21 a_n1952_n1488# 0.044844f
C160 minus.n22 a_n1952_n1488# 0.044844f
C161 minus.n23 a_n1952_n1488# 0.044844f
C162 minus.t3 a_n1952_n1488# 0.282392f
C163 minus.n24 a_n1952_n1488# 0.164472f
C164 minus.n25 a_n1952_n1488# 0.010176f
C165 minus.t5 a_n1952_n1488# 0.282392f
C166 minus.n26 a_n1952_n1488# 0.161983f
C167 minus.n27 a_n1952_n1488# 0.307746f
C168 minus.n28 a_n1952_n1488# 1.42599f
.ends

