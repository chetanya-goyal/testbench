* NGSPICE file created from diffpair211.ext - technology: sky130A

.subckt diffpair211 minus drain_right drain_left source plus
X0 a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X1 a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X2 a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X3 drain_right.t3 minus.t0 source.t6 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X4 drain_left.t3 plus.t0 source.t0 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X5 a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X6 source.t5 minus.t1 drain_right.t2 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X7 drain_right.t1 minus.t2 source.t7 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X8 source.t4 minus.t3 drain_right.t0 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X9 drain_left.t2 plus.t1 source.t1 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X10 source.t3 plus.t2 drain_left.t1 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X11 source.t2 plus.t3 drain_left.t0 a_n1274_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n0 minus.t2 206.953
R1 minus.n1 minus.t3 206.953
R2 minus.n0 minus.t1 206.929
R3 minus.n1 minus.t0 206.929
R4 minus.n2 minus.n0 97.4828
R5 minus.n2 minus.n1 76.854
R6 minus minus.n2 0.188
R7 source.n0 source.t1 69.6943
R8 source.n1 source.t3 69.6943
R9 source.n2 source.t7 69.6943
R10 source.n3 source.t5 69.6943
R11 source.n7 source.t6 69.6942
R12 source.n6 source.t4 69.6942
R13 source.n5 source.t0 69.6942
R14 source.n4 source.t2 69.6942
R15 source.n4 source.n3 15.2713
R16 source.n8 source.n0 9.60747
R17 source.n8 source.n7 5.66429
R18 source.n3 source.n2 0.802224
R19 source.n1 source.n0 0.802224
R20 source.n5 source.n4 0.802224
R21 source.n7 source.n6 0.802224
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 101.371
R26 drain_right drain_right.n1 86.2276
R27 drain_right.n0 drain_right.t0 6.6005
R28 drain_right.n0 drain_right.t3 6.6005
R29 drain_right.n1 drain_right.t2 6.6005
R30 drain_right.n1 drain_right.t1 6.6005
R31 plus.n0 plus.t2 206.953
R32 plus.n1 plus.t0 206.953
R33 plus.n0 plus.t1 206.929
R34 plus.n1 plus.t3 206.929
R35 plus plus.n1 94.773
R36 plus plus.n0 79.0889
R37 drain_left drain_left.n0 101.924
R38 drain_left drain_left.n1 86.2276
R39 drain_left.n0 drain_left.t0 6.6005
R40 drain_left.n0 drain_left.t3 6.6005
R41 drain_left.n1 drain_left.t1 6.6005
R42 drain_left.n1 drain_left.t2 6.6005
C0 plus drain_right 0.278426f
C1 plus source 0.992459f
C2 plus minus 3.06677f
C3 drain_left drain_right 0.544764f
C4 drain_left source 2.93289f
C5 drain_left minus 0.175416f
C6 source drain_right 2.93326f
C7 minus drain_right 0.951666f
C8 source minus 0.978461f
C9 plus drain_left 1.07136f
C10 drain_right a_n1274_n1488# 3.73111f
C11 drain_left a_n1274_n1488# 3.87356f
C12 source a_n1274_n1488# 3.482985f
C13 minus a_n1274_n1488# 4.072623f
C14 plus a_n1274_n1488# 5.61492f
C15 drain_left.t0 a_n1274_n1488# 0.046685f
C16 drain_left.t3 a_n1274_n1488# 0.046685f
C17 drain_left.n0 a_n1274_n1488# 0.451926f
C18 drain_left.t1 a_n1274_n1488# 0.046685f
C19 drain_left.t2 a_n1274_n1488# 0.046685f
C20 drain_left.n1 a_n1274_n1488# 0.36955f
C21 plus.t1 a_n1274_n1488# 0.193061f
C22 plus.t2 a_n1274_n1488# 0.193077f
C23 plus.n0 a_n1274_n1488# 0.228273f
C24 plus.t3 a_n1274_n1488# 0.193061f
C25 plus.t0 a_n1274_n1488# 0.193077f
C26 plus.n1 a_n1274_n1488# 0.388602f
C27 drain_right.t0 a_n1274_n1488# 0.047959f
C28 drain_right.t3 a_n1274_n1488# 0.047959f
C29 drain_right.n0 a_n1274_n1488# 0.453325f
C30 drain_right.t2 a_n1274_n1488# 0.047959f
C31 drain_right.t1 a_n1274_n1488# 0.047959f
C32 drain_right.n1 a_n1274_n1488# 0.379635f
C33 source.t1 a_n1274_n1488# 0.305163f
C34 source.n0 a_n1274_n1488# 0.43905f
C35 source.t3 a_n1274_n1488# 0.305163f
C36 source.n1 a_n1274_n1488# 0.226631f
C37 source.t7 a_n1274_n1488# 0.305163f
C38 source.n2 a_n1274_n1488# 0.226631f
C39 source.t5 a_n1274_n1488# 0.305163f
C40 source.n3 a_n1274_n1488# 0.603764f
C41 source.t2 a_n1274_n1488# 0.305161f
C42 source.n4 a_n1274_n1488# 0.603766f
C43 source.t0 a_n1274_n1488# 0.305161f
C44 source.n5 a_n1274_n1488# 0.226632f
C45 source.t4 a_n1274_n1488# 0.305161f
C46 source.n6 a_n1274_n1488# 0.226632f
C47 source.t6 a_n1274_n1488# 0.305161f
C48 source.n7 a_n1274_n1488# 0.324376f
C49 source.n8 a_n1274_n1488# 0.455129f
C50 minus.t2 a_n1274_n1488# 0.188918f
C51 minus.t1 a_n1274_n1488# 0.188902f
C52 minus.n0 a_n1274_n1488# 0.406366f
C53 minus.t3 a_n1274_n1488# 0.188918f
C54 minus.t0 a_n1274_n1488# 0.188902f
C55 minus.n1 a_n1274_n1488# 0.212854f
C56 minus.n2 a_n1274_n1488# 1.70346f
.ends

