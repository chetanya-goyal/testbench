* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t11 minus.t0 drain_right.t3 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 source.t5 plus.t0 drain_left.t5 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X2 source.t10 minus.t1 drain_right.t2 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 drain_left.t4 plus.t1 source.t0 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X4 a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X5 drain_right.t1 minus.t2 source.t9 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X6 a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X7 a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X8 drain_right.t4 minus.t3 source.t8 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X9 source.t4 plus.t2 drain_left.t3 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X10 drain_right.t0 minus.t4 source.t7 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X11 drain_left.t2 plus.t3 source.t2 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X12 drain_right.t5 minus.t5 source.t6 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X13 drain_left.t1 plus.t4 source.t1 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X14 drain_left.t0 plus.t5 source.t3 a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X15 a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# a_n1380_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
R0 minus.n0 minus.t3 201.787
R1 minus.n4 minus.t5 201.787
R2 minus.n1 minus.t1 174.966
R3 minus.n2 minus.t2 174.966
R4 minus.n5 minus.t0 174.966
R5 minus.n6 minus.t4 174.966
R6 minus.n3 minus.n2 161.3
R7 minus.n7 minus.n6 161.3
R8 minus.n2 minus.n1 48.2005
R9 minus.n6 minus.n5 48.2005
R10 minus.n3 minus.n0 45.1367
R11 minus.n7 minus.n4 45.1367
R12 minus.n8 minus.n3 26.8054
R13 minus.n1 minus.n0 13.3799
R14 minus.n5 minus.n4 13.3799
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 drain_right.n2 drain_right.n0 289.615
R18 drain_right.n12 drain_right.n10 289.615
R19 drain_right.n3 drain_right.n2 185
R20 drain_right.n13 drain_right.n12 185
R21 drain_right.t5 drain_right.n1 167.117
R22 drain_right.t1 drain_right.n11 167.117
R23 drain_right.n17 drain_right.n9 101.511
R24 drain_right.n8 drain_right.n7 100.919
R25 drain_right.n2 drain_right.t5 52.3082
R26 drain_right.n12 drain_right.t1 52.3082
R27 drain_right.n8 drain_right.n6 48.5697
R28 drain_right.n17 drain_right.n16 48.0884
R29 drain_right drain_right.n8 21.2058
R30 drain_right.n7 drain_right.t3 9.9005
R31 drain_right.n7 drain_right.t0 9.9005
R32 drain_right.n9 drain_right.t2 9.9005
R33 drain_right.n9 drain_right.t4 9.9005
R34 drain_right.n3 drain_right.n1 9.71174
R35 drain_right.n13 drain_right.n11 9.71174
R36 drain_right.n6 drain_right.n5 9.45567
R37 drain_right.n16 drain_right.n15 9.45567
R38 drain_right.n5 drain_right.n4 9.3005
R39 drain_right.n15 drain_right.n14 9.3005
R40 drain_right.n6 drain_right.n0 8.14595
R41 drain_right.n16 drain_right.n10 8.14595
R42 drain_right.n4 drain_right.n3 7.3702
R43 drain_right.n14 drain_right.n13 7.3702
R44 drain_right drain_right.n17 6.01097
R45 drain_right.n4 drain_right.n0 5.81868
R46 drain_right.n14 drain_right.n10 5.81868
R47 drain_right.n5 drain_right.n1 3.44771
R48 drain_right.n15 drain_right.n11 3.44771
R49 source.n34 source.n32 289.615
R50 source.n24 source.n22 289.615
R51 source.n2 source.n0 289.615
R52 source.n12 source.n10 289.615
R53 source.n35 source.n34 185
R54 source.n25 source.n24 185
R55 source.n3 source.n2 185
R56 source.n13 source.n12 185
R57 source.t7 source.n33 167.117
R58 source.t3 source.n23 167.117
R59 source.t1 source.n1 167.117
R60 source.t8 source.n11 167.117
R61 source.n9 source.n8 84.1169
R62 source.n19 source.n18 84.1169
R63 source.n31 source.n30 84.1168
R64 source.n21 source.n20 84.1168
R65 source.n34 source.t7 52.3082
R66 source.n24 source.t3 52.3082
R67 source.n2 source.t1 52.3082
R68 source.n12 source.t8 52.3082
R69 source.n39 source.n38 31.4096
R70 source.n29 source.n28 31.4096
R71 source.n7 source.n6 31.4096
R72 source.n17 source.n16 31.4096
R73 source.n21 source.n19 15.143
R74 source.n30 source.t6 9.9005
R75 source.n30 source.t11 9.9005
R76 source.n20 source.t2 9.9005
R77 source.n20 source.t5 9.9005
R78 source.n8 source.t0 9.9005
R79 source.n8 source.t4 9.9005
R80 source.n18 source.t9 9.9005
R81 source.n18 source.t10 9.9005
R82 source.n35 source.n33 9.71174
R83 source.n25 source.n23 9.71174
R84 source.n3 source.n1 9.71174
R85 source.n13 source.n11 9.71174
R86 source.n38 source.n37 9.45567
R87 source.n28 source.n27 9.45567
R88 source.n6 source.n5 9.45567
R89 source.n16 source.n15 9.45567
R90 source.n37 source.n36 9.3005
R91 source.n27 source.n26 9.3005
R92 source.n5 source.n4 9.3005
R93 source.n15 source.n14 9.3005
R94 source.n40 source.n7 8.8068
R95 source.n38 source.n32 8.14595
R96 source.n28 source.n22 8.14595
R97 source.n6 source.n0 8.14595
R98 source.n16 source.n10 8.14595
R99 source.n36 source.n35 7.3702
R100 source.n26 source.n25 7.3702
R101 source.n4 source.n3 7.3702
R102 source.n14 source.n13 7.3702
R103 source.n36 source.n32 5.81868
R104 source.n26 source.n22 5.81868
R105 source.n4 source.n0 5.81868
R106 source.n14 source.n10 5.81868
R107 source.n40 source.n39 5.62119
R108 source.n37 source.n33 3.44771
R109 source.n27 source.n23 3.44771
R110 source.n5 source.n1 3.44771
R111 source.n15 source.n11 3.44771
R112 source.n17 source.n9 0.828086
R113 source.n31 source.n29 0.828086
R114 source.n19 source.n17 0.716017
R115 source.n9 source.n7 0.716017
R116 source.n29 source.n21 0.716017
R117 source.n39 source.n31 0.716017
R118 source source.n40 0.188
R119 plus.n0 plus.t1 201.787
R120 plus.n4 plus.t5 201.787
R121 plus.n2 plus.t4 174.966
R122 plus.n1 plus.t2 174.966
R123 plus.n6 plus.t3 174.966
R124 plus.n5 plus.t0 174.966
R125 plus.n3 plus.n2 161.3
R126 plus.n7 plus.n6 161.3
R127 plus.n2 plus.n1 48.2005
R128 plus.n6 plus.n5 48.2005
R129 plus.n3 plus.n0 45.1367
R130 plus.n7 plus.n4 45.1367
R131 plus plus.n7 24.4744
R132 plus.n1 plus.n0 13.3799
R133 plus.n5 plus.n4 13.3799
R134 plus plus.n3 8.38876
R135 drain_left.n2 drain_left.n0 289.615
R136 drain_left.n11 drain_left.n9 289.615
R137 drain_left.n3 drain_left.n2 185
R138 drain_left.n12 drain_left.n11 185
R139 drain_left.t2 drain_left.n1 167.117
R140 drain_left.t4 drain_left.n10 167.117
R141 drain_left.n8 drain_left.n7 100.919
R142 drain_left.n17 drain_left.n16 100.796
R143 drain_left.n2 drain_left.t2 52.3082
R144 drain_left.n11 drain_left.t4 52.3082
R145 drain_left.n17 drain_left.n15 48.8039
R146 drain_left.n8 drain_left.n6 48.5697
R147 drain_left drain_left.n8 21.759
R148 drain_left.n7 drain_left.t5 9.9005
R149 drain_left.n7 drain_left.t0 9.9005
R150 drain_left.n16 drain_left.t3 9.9005
R151 drain_left.n16 drain_left.t1 9.9005
R152 drain_left.n3 drain_left.n1 9.71174
R153 drain_left.n12 drain_left.n10 9.71174
R154 drain_left.n6 drain_left.n5 9.45567
R155 drain_left.n15 drain_left.n14 9.45567
R156 drain_left.n5 drain_left.n4 9.3005
R157 drain_left.n14 drain_left.n13 9.3005
R158 drain_left.n6 drain_left.n0 8.14595
R159 drain_left.n15 drain_left.n9 8.14595
R160 drain_left.n4 drain_left.n3 7.3702
R161 drain_left.n13 drain_left.n12 7.3702
R162 drain_left drain_left.n17 6.36873
R163 drain_left.n4 drain_left.n0 5.81868
R164 drain_left.n13 drain_left.n9 5.81868
R165 drain_left.n5 drain_left.n1 3.44771
R166 drain_left.n14 drain_left.n10 3.44771
C0 drain_right minus 0.879687f
C1 drain_right source 3.39246f
C2 drain_left drain_right 0.635665f
C3 minus source 1.00765f
C4 drain_left minus 0.177479f
C5 drain_left source 3.39459f
C6 plus drain_right 0.292135f
C7 plus minus 3.02475f
C8 plus source 1.0217f
C9 plus drain_left 1.00992f
C10 drain_right a_n1380_n1288# 3.121646f
C11 drain_left a_n1380_n1288# 3.291576f
C12 source a_n1380_n1288# 2.406267f
C13 minus a_n1380_n1288# 4.485902f
C14 plus a_n1380_n1288# 5.131541f
C15 drain_left.n0 a_n1380_n1288# 0.027318f
C16 drain_left.n1 a_n1380_n1288# 0.060445f
C17 drain_left.t2 a_n1380_n1288# 0.045361f
C18 drain_left.n2 a_n1380_n1288# 0.047307f
C19 drain_left.n3 a_n1380_n1288# 0.01525f
C20 drain_left.n4 a_n1380_n1288# 0.010058f
C21 drain_left.n5 a_n1380_n1288# 0.133236f
C22 drain_left.n6 a_n1380_n1288# 0.043527f
C23 drain_left.t5 a_n1380_n1288# 0.029581f
C24 drain_left.t0 a_n1380_n1288# 0.029581f
C25 drain_left.n7 a_n1380_n1288# 0.186089f
C26 drain_left.n8 a_n1380_n1288# 0.7256f
C27 drain_left.n9 a_n1380_n1288# 0.027318f
C28 drain_left.n10 a_n1380_n1288# 0.060445f
C29 drain_left.t4 a_n1380_n1288# 0.045361f
C30 drain_left.n11 a_n1380_n1288# 0.047307f
C31 drain_left.n12 a_n1380_n1288# 0.01525f
C32 drain_left.n13 a_n1380_n1288# 0.010058f
C33 drain_left.n14 a_n1380_n1288# 0.133236f
C34 drain_left.n15 a_n1380_n1288# 0.044032f
C35 drain_left.t3 a_n1380_n1288# 0.029581f
C36 drain_left.t1 a_n1380_n1288# 0.029581f
C37 drain_left.n16 a_n1380_n1288# 0.185839f
C38 drain_left.n17 a_n1380_n1288# 0.467821f
C39 plus.t1 a_n1380_n1288# 0.11114f
C40 plus.n0 a_n1380_n1288# 0.063987f
C41 plus.t4 a_n1380_n1288# 0.101419f
C42 plus.t2 a_n1380_n1288# 0.101419f
C43 plus.n1 a_n1380_n1288# 0.080487f
C44 plus.n2 a_n1380_n1288# 0.073056f
C45 plus.n3 a_n1380_n1288# 0.337612f
C46 plus.t5 a_n1380_n1288# 0.11114f
C47 plus.n4 a_n1380_n1288# 0.063987f
C48 plus.t3 a_n1380_n1288# 0.101419f
C49 plus.t0 a_n1380_n1288# 0.101419f
C50 plus.n5 a_n1380_n1288# 0.080487f
C51 plus.n6 a_n1380_n1288# 0.073056f
C52 plus.n7 a_n1380_n1288# 0.772792f
C53 source.n0 a_n1380_n1288# 0.034775f
C54 source.n1 a_n1380_n1288# 0.076944f
C55 source.t1 a_n1380_n1288# 0.057743f
C56 source.n2 a_n1380_n1288# 0.06022f
C57 source.n3 a_n1380_n1288# 0.019412f
C58 source.n4 a_n1380_n1288# 0.012803f
C59 source.n5 a_n1380_n1288# 0.169604f
C60 source.n6 a_n1380_n1288# 0.038122f
C61 source.n7 a_n1380_n1288# 0.383217f
C62 source.t0 a_n1380_n1288# 0.037656f
C63 source.t4 a_n1380_n1288# 0.037656f
C64 source.n8 a_n1380_n1288# 0.201306f
C65 source.n9 a_n1380_n1288# 0.303701f
C66 source.n10 a_n1380_n1288# 0.034775f
C67 source.n11 a_n1380_n1288# 0.076944f
C68 source.t8 a_n1380_n1288# 0.057743f
C69 source.n12 a_n1380_n1288# 0.06022f
C70 source.n13 a_n1380_n1288# 0.019412f
C71 source.n14 a_n1380_n1288# 0.012803f
C72 source.n15 a_n1380_n1288# 0.169604f
C73 source.n16 a_n1380_n1288# 0.038122f
C74 source.n17 a_n1380_n1288# 0.138081f
C75 source.t9 a_n1380_n1288# 0.037656f
C76 source.t10 a_n1380_n1288# 0.037656f
C77 source.n18 a_n1380_n1288# 0.201306f
C78 source.n19 a_n1380_n1288# 0.828882f
C79 source.t2 a_n1380_n1288# 0.037656f
C80 source.t5 a_n1380_n1288# 0.037656f
C81 source.n20 a_n1380_n1288# 0.201305f
C82 source.n21 a_n1380_n1288# 0.828883f
C83 source.n22 a_n1380_n1288# 0.034775f
C84 source.n23 a_n1380_n1288# 0.076944f
C85 source.t3 a_n1380_n1288# 0.057743f
C86 source.n24 a_n1380_n1288# 0.06022f
C87 source.n25 a_n1380_n1288# 0.019412f
C88 source.n26 a_n1380_n1288# 0.012803f
C89 source.n27 a_n1380_n1288# 0.169604f
C90 source.n28 a_n1380_n1288# 0.038122f
C91 source.n29 a_n1380_n1288# 0.138081f
C92 source.t6 a_n1380_n1288# 0.037656f
C93 source.t11 a_n1380_n1288# 0.037656f
C94 source.n30 a_n1380_n1288# 0.201305f
C95 source.n31 a_n1380_n1288# 0.303702f
C96 source.n32 a_n1380_n1288# 0.034775f
C97 source.n33 a_n1380_n1288# 0.076944f
C98 source.t7 a_n1380_n1288# 0.057743f
C99 source.n34 a_n1380_n1288# 0.06022f
C100 source.n35 a_n1380_n1288# 0.019412f
C101 source.n36 a_n1380_n1288# 0.012803f
C102 source.n37 a_n1380_n1288# 0.169604f
C103 source.n38 a_n1380_n1288# 0.038122f
C104 source.n39 a_n1380_n1288# 0.25563f
C105 source.n40 a_n1380_n1288# 0.594761f
C106 drain_right.n0 a_n1380_n1288# 0.02792f
C107 drain_right.n1 a_n1380_n1288# 0.061776f
C108 drain_right.t5 a_n1380_n1288# 0.046359f
C109 drain_right.n2 a_n1380_n1288# 0.048348f
C110 drain_right.n3 a_n1380_n1288# 0.015586f
C111 drain_right.n4 a_n1380_n1288# 0.010279f
C112 drain_right.n5 a_n1380_n1288# 0.136169f
C113 drain_right.n6 a_n1380_n1288# 0.044485f
C114 drain_right.t3 a_n1380_n1288# 0.030232f
C115 drain_right.t0 a_n1380_n1288# 0.030232f
C116 drain_right.n7 a_n1380_n1288# 0.190185f
C117 drain_right.n8 a_n1380_n1288# 0.703912f
C118 drain_right.t2 a_n1380_n1288# 0.030232f
C119 drain_right.t4 a_n1380_n1288# 0.030232f
C120 drain_right.n9 a_n1380_n1288# 0.191637f
C121 drain_right.n10 a_n1380_n1288# 0.02792f
C122 drain_right.n11 a_n1380_n1288# 0.061776f
C123 drain_right.t1 a_n1380_n1288# 0.046359f
C124 drain_right.n12 a_n1380_n1288# 0.048348f
C125 drain_right.n13 a_n1380_n1288# 0.015586f
C126 drain_right.n14 a_n1380_n1288# 0.010279f
C127 drain_right.n15 a_n1380_n1288# 0.136169f
C128 drain_right.n16 a_n1380_n1288# 0.043823f
C129 drain_right.n17 a_n1380_n1288# 0.488681f
C130 minus.t3 a_n1380_n1288# 0.10874f
C131 minus.n0 a_n1380_n1288# 0.062605f
C132 minus.t1 a_n1380_n1288# 0.099228f
C133 minus.n1 a_n1380_n1288# 0.078749f
C134 minus.t2 a_n1380_n1288# 0.099228f
C135 minus.n2 a_n1380_n1288# 0.071478f
C136 minus.n3 a_n1380_n1288# 0.783538f
C137 minus.t5 a_n1380_n1288# 0.10874f
C138 minus.n4 a_n1380_n1288# 0.062605f
C139 minus.t0 a_n1380_n1288# 0.099228f
C140 minus.n5 a_n1380_n1288# 0.078749f
C141 minus.t4 a_n1380_n1288# 0.099228f
C142 minus.n6 a_n1380_n1288# 0.071478f
C143 minus.n7 a_n1380_n1288# 0.310604f
C144 minus.n8 a_n1380_n1288# 0.844763f
.ends

