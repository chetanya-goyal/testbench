* NGSPICE file created from diffpair55.ext - technology: sky130A

.subckt diffpair55 minus drain_right drain_left source plus
X0 source.t21 plus.t0 drain_left.t11 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X1 drain_left.t3 plus.t1 source.t20 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X2 drain_right.t11 minus.t0 source.t22 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X3 source.t23 minus.t1 drain_right.t10 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X4 source.t4 minus.t2 drain_right.t9 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 drain_right.t8 minus.t3 source.t0 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X6 source.t19 plus.t2 drain_left.t4 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X7 a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X8 source.t18 plus.t3 drain_left.t2 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X9 source.t3 minus.t4 drain_right.t7 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X10 drain_right.t6 minus.t5 source.t8 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 drain_left.t7 plus.t4 source.t17 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X12 drain_left.t0 plus.t5 source.t16 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 source.t7 minus.t6 drain_right.t5 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 drain_left.t8 plus.t6 source.t15 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 source.t14 plus.t7 drain_left.t9 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X16 drain_right.t4 minus.t7 source.t9 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X17 a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X18 drain_left.t6 plus.t8 source.t13 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X19 source.t12 plus.t9 drain_left.t1 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X20 source.t2 minus.t8 drain_right.t3 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X22 source.t11 plus.t10 drain_left.t10 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X23 a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X24 drain_right.t2 minus.t9 source.t6 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X25 drain_right.t1 minus.t10 source.t1 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X26 source.t5 minus.t11 drain_right.t0 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X27 drain_left.t5 plus.t11 source.t10 a_n2018_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n8 plus.n1 161.3
R1 plus.n9 plus.n0 161.3
R2 plus.n11 plus.n10 161.3
R3 plus.n20 plus.n13 161.3
R4 plus.n21 plus.n12 161.3
R5 plus.n23 plus.n22 161.3
R6 plus.n4 plus.t9 130.698
R7 plus.n16 plus.t4 130.698
R8 plus.n10 plus.t1 105.638
R9 plus.n8 plus.t3 105.638
R10 plus.n7 plus.t5 105.638
R11 plus.n6 plus.t7 105.638
R12 plus.n5 plus.t8 105.638
R13 plus.n22 plus.t2 105.638
R14 plus.n20 plus.t6 105.638
R15 plus.n19 plus.t10 105.638
R16 plus.n18 plus.t11 105.638
R17 plus.n17 plus.t0 105.638
R18 plus.n6 plus.n3 80.6037
R19 plus.n7 plus.n2 80.6037
R20 plus.n18 plus.n15 80.6037
R21 plus.n19 plus.n14 80.6037
R22 plus.n8 plus.n7 48.2005
R23 plus.n7 plus.n6 48.2005
R24 plus.n6 plus.n5 48.2005
R25 plus.n20 plus.n19 48.2005
R26 plus.n19 plus.n18 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n4 plus.n3 45.0744
R29 plus.n16 plus.n15 45.0744
R30 plus.n10 plus.n9 40.1672
R31 plus.n22 plus.n21 40.1672
R32 plus plus.n23 26.5672
R33 plus.n5 plus.n4 16.1124
R34 plus.n17 plus.n16 16.1124
R35 plus plus.n11 8.06489
R36 plus.n9 plus.n8 8.03383
R37 plus.n21 plus.n20 8.03383
R38 plus.n3 plus.n2 0.380177
R39 plus.n15 plus.n14 0.380177
R40 plus.n2 plus.n1 0.285035
R41 plus.n14 plus.n13 0.285035
R42 plus.n1 plus.n0 0.189894
R43 plus.n11 plus.n0 0.189894
R44 plus.n23 plus.n12 0.189894
R45 plus.n13 plus.n12 0.189894
R46 drain_left.n6 drain_left.n4 240.935
R47 drain_left.n3 drain_left.n2 240.879
R48 drain_left.n3 drain_left.n0 240.879
R49 drain_left.n8 drain_left.n7 240.132
R50 drain_left.n6 drain_left.n5 240.132
R51 drain_left.n3 drain_left.n1 240.131
R52 drain_left drain_left.n3 23.0424
R53 drain_left.n1 drain_left.t10 19.8005
R54 drain_left.n1 drain_left.t5 19.8005
R55 drain_left.n2 drain_left.t11 19.8005
R56 drain_left.n2 drain_left.t7 19.8005
R57 drain_left.n0 drain_left.t4 19.8005
R58 drain_left.n0 drain_left.t8 19.8005
R59 drain_left.n7 drain_left.t2 19.8005
R60 drain_left.n7 drain_left.t3 19.8005
R61 drain_left.n5 drain_left.t9 19.8005
R62 drain_left.n5 drain_left.t0 19.8005
R63 drain_left.n4 drain_left.t1 19.8005
R64 drain_left.n4 drain_left.t6 19.8005
R65 drain_left drain_left.n8 6.45494
R66 drain_left.n8 drain_left.n6 0.802224
R67 source.n0 source.t20 243.255
R68 source.n5 source.t12 243.255
R69 source.n6 source.t9 243.255
R70 source.n11 source.t23 243.255
R71 source.n23 source.t6 243.254
R72 source.n18 source.t5 243.254
R73 source.n17 source.t17 243.254
R74 source.n12 source.t19 243.254
R75 source.n2 source.n1 223.454
R76 source.n4 source.n3 223.454
R77 source.n8 source.n7 223.454
R78 source.n10 source.n9 223.454
R79 source.n22 source.n21 223.453
R80 source.n20 source.n19 223.453
R81 source.n16 source.n15 223.453
R82 source.n14 source.n13 223.453
R83 source.n21 source.t1 19.8005
R84 source.n21 source.t2 19.8005
R85 source.n19 source.t0 19.8005
R86 source.n19 source.t4 19.8005
R87 source.n15 source.t10 19.8005
R88 source.n15 source.t21 19.8005
R89 source.n13 source.t15 19.8005
R90 source.n13 source.t11 19.8005
R91 source.n1 source.t16 19.8005
R92 source.n1 source.t18 19.8005
R93 source.n3 source.t13 19.8005
R94 source.n3 source.t14 19.8005
R95 source.n7 source.t8 19.8005
R96 source.n7 source.t7 19.8005
R97 source.n9 source.t22 19.8005
R98 source.n9 source.t3 19.8005
R99 source.n12 source.n11 13.7561
R100 source.n24 source.n0 8.09232
R101 source.n24 source.n23 5.66429
R102 source.n11 source.n10 0.802224
R103 source.n10 source.n8 0.802224
R104 source.n8 source.n6 0.802224
R105 source.n5 source.n4 0.802224
R106 source.n4 source.n2 0.802224
R107 source.n2 source.n0 0.802224
R108 source.n14 source.n12 0.802224
R109 source.n16 source.n14 0.802224
R110 source.n17 source.n16 0.802224
R111 source.n20 source.n18 0.802224
R112 source.n22 source.n20 0.802224
R113 source.n23 source.n22 0.802224
R114 source.n6 source.n5 0.470328
R115 source.n18 source.n17 0.470328
R116 source source.n24 0.188
R117 minus.n11 minus.n10 161.3
R118 minus.n9 minus.n0 161.3
R119 minus.n8 minus.n7 161.3
R120 minus.n23 minus.n22 161.3
R121 minus.n21 minus.n12 161.3
R122 minus.n20 minus.n19 161.3
R123 minus.n2 minus.t7 130.698
R124 minus.n14 minus.t11 130.698
R125 minus.n3 minus.t6 105.638
R126 minus.n4 minus.t5 105.638
R127 minus.n1 minus.t4 105.638
R128 minus.n8 minus.t0 105.638
R129 minus.n10 minus.t1 105.638
R130 minus.n15 minus.t3 105.638
R131 minus.n16 minus.t2 105.638
R132 minus.n13 minus.t10 105.638
R133 minus.n20 minus.t8 105.638
R134 minus.n22 minus.t9 105.638
R135 minus.n6 minus.n1 80.6037
R136 minus.n5 minus.n4 80.6037
R137 minus.n18 minus.n13 80.6037
R138 minus.n17 minus.n16 80.6037
R139 minus.n4 minus.n3 48.2005
R140 minus.n4 minus.n1 48.2005
R141 minus.n8 minus.n1 48.2005
R142 minus.n16 minus.n15 48.2005
R143 minus.n16 minus.n13 48.2005
R144 minus.n20 minus.n13 48.2005
R145 minus.n5 minus.n2 45.0744
R146 minus.n17 minus.n14 45.0744
R147 minus.n10 minus.n9 40.1672
R148 minus.n22 minus.n21 40.1672
R149 minus.n24 minus.n11 28.5194
R150 minus.n3 minus.n2 16.1124
R151 minus.n15 minus.n14 16.1124
R152 minus.n9 minus.n8 8.03383
R153 minus.n21 minus.n20 8.03383
R154 minus.n24 minus.n23 6.58762
R155 minus.n6 minus.n5 0.380177
R156 minus.n18 minus.n17 0.380177
R157 minus.n7 minus.n6 0.285035
R158 minus.n19 minus.n18 0.285035
R159 minus.n11 minus.n0 0.189894
R160 minus.n7 minus.n0 0.189894
R161 minus.n19 minus.n12 0.189894
R162 minus.n23 minus.n12 0.189894
R163 minus minus.n24 0.188
R164 drain_right.n6 drain_right.n4 240.935
R165 drain_right.n3 drain_right.n2 240.879
R166 drain_right.n3 drain_right.n0 240.879
R167 drain_right.n6 drain_right.n5 240.132
R168 drain_right.n8 drain_right.n7 240.132
R169 drain_right.n3 drain_right.n1 240.131
R170 drain_right drain_right.n3 22.4891
R171 drain_right.n1 drain_right.t9 19.8005
R172 drain_right.n1 drain_right.t1 19.8005
R173 drain_right.n2 drain_right.t3 19.8005
R174 drain_right.n2 drain_right.t2 19.8005
R175 drain_right.n0 drain_right.t0 19.8005
R176 drain_right.n0 drain_right.t8 19.8005
R177 drain_right.n4 drain_right.t5 19.8005
R178 drain_right.n4 drain_right.t4 19.8005
R179 drain_right.n5 drain_right.t7 19.8005
R180 drain_right.n5 drain_right.t6 19.8005
R181 drain_right.n7 drain_right.t10 19.8005
R182 drain_right.n7 drain_right.t11 19.8005
R183 drain_right drain_right.n8 6.45494
R184 drain_right.n8 drain_right.n6 0.802224
C0 plus drain_right 0.360795f
C1 drain_left drain_right 1.01302f
C2 source drain_right 3.8463f
C3 minus plus 3.63638f
C4 minus drain_left 0.179185f
C5 minus source 1.48739f
C6 plus drain_left 1.23685f
C7 source plus 1.50125f
C8 minus drain_right 1.03985f
C9 source drain_left 3.8448f
C10 drain_right a_n2018_n1088# 3.55673f
C11 drain_left a_n2018_n1088# 3.80964f
C12 source a_n2018_n1088# 2.54919f
C13 minus a_n2018_n1088# 7.021203f
C14 plus a_n2018_n1088# 7.627316f
C15 drain_right.t0 a_n2018_n1088# 0.016092f
C16 drain_right.t8 a_n2018_n1088# 0.016092f
C17 drain_right.n0 a_n2018_n1088# 0.063311f
C18 drain_right.t9 a_n2018_n1088# 0.016092f
C19 drain_right.t1 a_n2018_n1088# 0.016092f
C20 drain_right.n1 a_n2018_n1088# 0.062528f
C21 drain_right.t3 a_n2018_n1088# 0.016092f
C22 drain_right.t2 a_n2018_n1088# 0.016092f
C23 drain_right.n2 a_n2018_n1088# 0.063311f
C24 drain_right.n3 a_n2018_n1088# 1.25766f
C25 drain_right.t5 a_n2018_n1088# 0.016092f
C26 drain_right.t4 a_n2018_n1088# 0.016092f
C27 drain_right.n4 a_n2018_n1088# 0.063379f
C28 drain_right.t7 a_n2018_n1088# 0.016092f
C29 drain_right.t6 a_n2018_n1088# 0.016092f
C30 drain_right.n5 a_n2018_n1088# 0.062528f
C31 drain_right.n6 a_n2018_n1088# 0.502579f
C32 drain_right.t10 a_n2018_n1088# 0.016092f
C33 drain_right.t11 a_n2018_n1088# 0.016092f
C34 drain_right.n7 a_n2018_n1088# 0.062528f
C35 drain_right.n8 a_n2018_n1088# 0.425182f
C36 minus.n0 a_n2018_n1088# 0.027659f
C37 minus.t4 a_n2018_n1088# 0.056274f
C38 minus.n1 a_n2018_n1088# 0.063556f
C39 minus.t0 a_n2018_n1088# 0.056274f
C40 minus.t7 a_n2018_n1088# 0.0672f
C41 minus.n2 a_n2018_n1088# 0.048166f
C42 minus.t6 a_n2018_n1088# 0.056274f
C43 minus.n3 a_n2018_n1088# 0.062546f
C44 minus.t5 a_n2018_n1088# 0.056274f
C45 minus.n4 a_n2018_n1088# 0.063556f
C46 minus.n5 a_n2018_n1088# 0.141755f
C47 minus.n6 a_n2018_n1088# 0.046069f
C48 minus.n7 a_n2018_n1088# 0.036907f
C49 minus.n8 a_n2018_n1088# 0.058218f
C50 minus.n9 a_n2018_n1088# 0.006276f
C51 minus.t1 a_n2018_n1088# 0.056274f
C52 minus.n10 a_n2018_n1088# 0.056342f
C53 minus.n11 a_n2018_n1088# 0.661572f
C54 minus.n12 a_n2018_n1088# 0.027659f
C55 minus.t10 a_n2018_n1088# 0.056274f
C56 minus.n13 a_n2018_n1088# 0.063556f
C57 minus.t11 a_n2018_n1088# 0.0672f
C58 minus.n14 a_n2018_n1088# 0.048166f
C59 minus.t3 a_n2018_n1088# 0.056274f
C60 minus.n15 a_n2018_n1088# 0.062546f
C61 minus.t2 a_n2018_n1088# 0.056274f
C62 minus.n16 a_n2018_n1088# 0.063556f
C63 minus.n17 a_n2018_n1088# 0.141755f
C64 minus.n18 a_n2018_n1088# 0.046069f
C65 minus.n19 a_n2018_n1088# 0.036907f
C66 minus.t8 a_n2018_n1088# 0.056274f
C67 minus.n20 a_n2018_n1088# 0.058218f
C68 minus.n21 a_n2018_n1088# 0.006276f
C69 minus.t9 a_n2018_n1088# 0.056274f
C70 minus.n22 a_n2018_n1088# 0.056342f
C71 minus.n23 a_n2018_n1088# 0.186512f
C72 minus.n24 a_n2018_n1088# 0.814506f
C73 source.t20 a_n2018_n1088# 0.105219f
C74 source.n0 a_n2018_n1088# 0.487427f
C75 source.t16 a_n2018_n1088# 0.018904f
C76 source.t18 a_n2018_n1088# 0.018904f
C77 source.n1 a_n2018_n1088# 0.06131f
C78 source.n2 a_n2018_n1088# 0.270526f
C79 source.t13 a_n2018_n1088# 0.018904f
C80 source.t14 a_n2018_n1088# 0.018904f
C81 source.n3 a_n2018_n1088# 0.06131f
C82 source.n4 a_n2018_n1088# 0.270526f
C83 source.t12 a_n2018_n1088# 0.105219f
C84 source.n5 a_n2018_n1088# 0.25259f
C85 source.t9 a_n2018_n1088# 0.105219f
C86 source.n6 a_n2018_n1088# 0.25259f
C87 source.t8 a_n2018_n1088# 0.018904f
C88 source.t7 a_n2018_n1088# 0.018904f
C89 source.n7 a_n2018_n1088# 0.06131f
C90 source.n8 a_n2018_n1088# 0.270526f
C91 source.t22 a_n2018_n1088# 0.018904f
C92 source.t3 a_n2018_n1088# 0.018904f
C93 source.n9 a_n2018_n1088# 0.06131f
C94 source.n10 a_n2018_n1088# 0.270526f
C95 source.t23 a_n2018_n1088# 0.105219f
C96 source.n11 a_n2018_n1088# 0.683359f
C97 source.t19 a_n2018_n1088# 0.105219f
C98 source.n12 a_n2018_n1088# 0.68336f
C99 source.t15 a_n2018_n1088# 0.018904f
C100 source.t11 a_n2018_n1088# 0.018904f
C101 source.n13 a_n2018_n1088# 0.06131f
C102 source.n14 a_n2018_n1088# 0.270526f
C103 source.t10 a_n2018_n1088# 0.018904f
C104 source.t21 a_n2018_n1088# 0.018904f
C105 source.n15 a_n2018_n1088# 0.06131f
C106 source.n16 a_n2018_n1088# 0.270526f
C107 source.t17 a_n2018_n1088# 0.105219f
C108 source.n17 a_n2018_n1088# 0.25259f
C109 source.t5 a_n2018_n1088# 0.105219f
C110 source.n18 a_n2018_n1088# 0.25259f
C111 source.t0 a_n2018_n1088# 0.018904f
C112 source.t4 a_n2018_n1088# 0.018904f
C113 source.n19 a_n2018_n1088# 0.06131f
C114 source.n20 a_n2018_n1088# 0.270526f
C115 source.t1 a_n2018_n1088# 0.018904f
C116 source.t2 a_n2018_n1088# 0.018904f
C117 source.n21 a_n2018_n1088# 0.06131f
C118 source.n22 a_n2018_n1088# 0.270526f
C119 source.t6 a_n2018_n1088# 0.105219f
C120 source.n23 a_n2018_n1088# 0.403432f
C121 source.n24 a_n2018_n1088# 0.492876f
C122 drain_left.t4 a_n2018_n1088# 0.015761f
C123 drain_left.t8 a_n2018_n1088# 0.015761f
C124 drain_left.n0 a_n2018_n1088# 0.062011f
C125 drain_left.t10 a_n2018_n1088# 0.015761f
C126 drain_left.t5 a_n2018_n1088# 0.015761f
C127 drain_left.n1 a_n2018_n1088# 0.061244f
C128 drain_left.t11 a_n2018_n1088# 0.015761f
C129 drain_left.t7 a_n2018_n1088# 0.015761f
C130 drain_left.n2 a_n2018_n1088# 0.062011f
C131 drain_left.n3 a_n2018_n1088# 1.27035f
C132 drain_left.t1 a_n2018_n1088# 0.015761f
C133 drain_left.t6 a_n2018_n1088# 0.015761f
C134 drain_left.n4 a_n2018_n1088# 0.062078f
C135 drain_left.t9 a_n2018_n1088# 0.015761f
C136 drain_left.t0 a_n2018_n1088# 0.015761f
C137 drain_left.n5 a_n2018_n1088# 0.061244f
C138 drain_left.n6 a_n2018_n1088# 0.49226f
C139 drain_left.t2 a_n2018_n1088# 0.015761f
C140 drain_left.t3 a_n2018_n1088# 0.015761f
C141 drain_left.n7 a_n2018_n1088# 0.061244f
C142 drain_left.n8 a_n2018_n1088# 0.416451f
C143 plus.n0 a_n2018_n1088# 0.028095f
C144 plus.t1 a_n2018_n1088# 0.057163f
C145 plus.t3 a_n2018_n1088# 0.057163f
C146 plus.n1 a_n2018_n1088# 0.03749f
C147 plus.t5 a_n2018_n1088# 0.057163f
C148 plus.n2 a_n2018_n1088# 0.046796f
C149 plus.t7 a_n2018_n1088# 0.057163f
C150 plus.n3 a_n2018_n1088# 0.143992f
C151 plus.t8 a_n2018_n1088# 0.057163f
C152 plus.t9 a_n2018_n1088# 0.068261f
C153 plus.n4 a_n2018_n1088# 0.048926f
C154 plus.n5 a_n2018_n1088# 0.063533f
C155 plus.n6 a_n2018_n1088# 0.064559f
C156 plus.n7 a_n2018_n1088# 0.064559f
C157 plus.n8 a_n2018_n1088# 0.059137f
C158 plus.n9 a_n2018_n1088# 0.006375f
C159 plus.n10 a_n2018_n1088# 0.057231f
C160 plus.n11 a_n2018_n1088# 0.19871f
C161 plus.n12 a_n2018_n1088# 0.028095f
C162 plus.t2 a_n2018_n1088# 0.057163f
C163 plus.n13 a_n2018_n1088# 0.03749f
C164 plus.t6 a_n2018_n1088# 0.057163f
C165 plus.n14 a_n2018_n1088# 0.046796f
C166 plus.t10 a_n2018_n1088# 0.057163f
C167 plus.n15 a_n2018_n1088# 0.143992f
C168 plus.t11 a_n2018_n1088# 0.057163f
C169 plus.t4 a_n2018_n1088# 0.068261f
C170 plus.n16 a_n2018_n1088# 0.048926f
C171 plus.t0 a_n2018_n1088# 0.057163f
C172 plus.n17 a_n2018_n1088# 0.063533f
C173 plus.n18 a_n2018_n1088# 0.064559f
C174 plus.n19 a_n2018_n1088# 0.064559f
C175 plus.n20 a_n2018_n1088# 0.059137f
C176 plus.n21 a_n2018_n1088# 0.006375f
C177 plus.n22 a_n2018_n1088# 0.057231f
C178 plus.n23 a_n2018_n1088# 0.650688f
.ends

