* NGSPICE file created from diffpair559.ext - technology: sky130A

.subckt diffpair559 minus drain_right drain_left source plus
X0 source.t42 plus.t0 drain_left.t19 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X1 drain_right.t23 minus.t0 source.t3 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X2 drain_left.t2 plus.t1 source.t41 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X3 source.t0 minus.t1 drain_right.t22 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X4 source.t11 minus.t2 drain_right.t21 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X5 source.t40 plus.t2 drain_left.t1 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X6 source.t39 plus.t3 drain_left.t16 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X7 drain_right.t20 minus.t3 source.t46 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X8 drain_right.t19 minus.t4 source.t4 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X9 source.t38 plus.t4 drain_left.t15 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X11 drain_right.t18 minus.t5 source.t45 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X12 source.t17 minus.t6 drain_right.t17 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X13 drain_left.t6 plus.t5 source.t37 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X14 source.t36 plus.t6 drain_left.t5 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X15 drain_right.t16 minus.t7 source.t15 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X16 a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X17 drain_right.t15 minus.t8 source.t6 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X18 source.t35 plus.t7 drain_left.t10 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X19 source.t5 minus.t9 drain_right.t14 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X20 drain_left.t9 plus.t8 source.t34 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X21 source.t9 minus.t10 drain_right.t13 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X22 source.t2 minus.t11 drain_right.t12 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X23 drain_right.t11 minus.t12 source.t8 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X24 drain_right.t10 minus.t13 source.t10 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X25 source.t33 plus.t9 drain_left.t12 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X26 drain_left.t11 plus.t10 source.t32 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X27 drain_right.t9 minus.t14 source.t43 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X28 drain_left.t4 plus.t11 source.t31 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X29 source.t30 plus.t12 drain_left.t3 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X30 source.t16 minus.t15 drain_right.t8 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X31 drain_right.t7 minus.t16 source.t18 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X32 drain_left.t14 plus.t13 source.t29 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X33 drain_left.t13 plus.t14 source.t28 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X34 source.t44 minus.t17 drain_right.t6 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X35 drain_right.t5 minus.t18 source.t7 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X36 drain_right.t4 minus.t19 source.t13 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X37 source.t27 plus.t15 drain_left.t21 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X38 a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X39 drain_left.t20 plus.t16 source.t26 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X40 drain_left.t8 plus.t17 source.t25 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X41 source.t47 minus.t20 drain_right.t3 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X42 source.t24 plus.t18 drain_left.t7 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X43 drain_left.t18 plus.t19 source.t23 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X44 source.t22 plus.t20 drain_left.t17 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X45 drain_left.t23 plus.t21 source.t21 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X46 drain_left.t22 plus.t22 source.t20 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X47 a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X48 source.t12 minus.t21 drain_right.t2 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X49 source.t19 plus.t23 drain_left.t0 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X50 source.t14 minus.t22 drain_right.t1 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X51 source.t1 minus.t23 drain_right.t0 a_n3654_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n10 plus.t23 522.415
R1 plus.n46 plus.t1 522.415
R2 plus.n34 plus.t5 500.979
R3 plus.n32 plus.t6 500.979
R4 plus.n31 plus.t8 500.979
R5 plus.n3 plus.t12 500.979
R6 plus.n25 plus.t14 500.979
R7 plus.n5 plus.t15 500.979
R8 plus.n20 plus.t16 500.979
R9 plus.n18 plus.t20 500.979
R10 plus.n8 plus.t17 500.979
R11 plus.n12 plus.t18 500.979
R12 plus.n11 plus.t21 500.979
R13 plus.n70 plus.t3 500.979
R14 plus.n68 plus.t11 500.979
R15 plus.n67 plus.t0 500.979
R16 plus.n39 plus.t10 500.979
R17 plus.n61 plus.t4 500.979
R18 plus.n41 plus.t13 500.979
R19 plus.n56 plus.t2 500.979
R20 plus.n54 plus.t19 500.979
R21 plus.n44 plus.t7 500.979
R22 plus.n48 plus.t22 500.979
R23 plus.n47 plus.t9 500.979
R24 plus.n14 plus.n13 161.3
R25 plus.n15 plus.n8 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n18 plus.n7 161.3
R28 plus.n19 plus.n6 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n25 plus.n4 161.3
R31 plus.n27 plus.n26 161.3
R32 plus.n28 plus.n3 161.3
R33 plus.n30 plus.n29 161.3
R34 plus.n33 plus.n0 161.3
R35 plus.n35 plus.n34 161.3
R36 plus.n50 plus.n49 161.3
R37 plus.n51 plus.n44 161.3
R38 plus.n53 plus.n52 161.3
R39 plus.n54 plus.n43 161.3
R40 plus.n55 plus.n42 161.3
R41 plus.n60 plus.n59 161.3
R42 plus.n61 plus.n40 161.3
R43 plus.n63 plus.n62 161.3
R44 plus.n64 plus.n39 161.3
R45 plus.n66 plus.n65 161.3
R46 plus.n69 plus.n36 161.3
R47 plus.n71 plus.n70 161.3
R48 plus.n12 plus.n9 80.6037
R49 plus.n21 plus.n20 80.6037
R50 plus.n22 plus.n5 80.6037
R51 plus.n31 plus.n2 80.6037
R52 plus.n32 plus.n1 80.6037
R53 plus.n48 plus.n45 80.6037
R54 plus.n57 plus.n56 80.6037
R55 plus.n58 plus.n41 80.6037
R56 plus.n67 plus.n38 80.6037
R57 plus.n68 plus.n37 80.6037
R58 plus.n32 plus.n31 48.2005
R59 plus.n20 plus.n5 48.2005
R60 plus.n12 plus.n11 48.2005
R61 plus.n68 plus.n67 48.2005
R62 plus.n56 plus.n41 48.2005
R63 plus.n48 plus.n47 48.2005
R64 plus.n31 plus.n30 44.549
R65 plus.n13 plus.n12 44.549
R66 plus.n67 plus.n66 44.549
R67 plus.n49 plus.n48 44.549
R68 plus.n24 plus.n5 41.6278
R69 plus.n20 plus.n19 41.6278
R70 plus.n60 plus.n41 41.6278
R71 plus.n56 plus.n55 41.6278
R72 plus.n33 plus.n32 38.7066
R73 plus.n69 plus.n68 38.7066
R74 plus plus.n71 38.1392
R75 plus.n10 plus.n9 31.6825
R76 plus.n46 plus.n45 31.6825
R77 plus.n26 plus.n3 25.5611
R78 plus.n17 plus.n8 25.5611
R79 plus.n62 plus.n39 25.5611
R80 plus.n53 plus.n44 25.5611
R81 plus.n26 plus.n25 22.6399
R82 plus.n18 plus.n17 22.6399
R83 plus.n62 plus.n61 22.6399
R84 plus.n54 plus.n53 22.6399
R85 plus.n11 plus.n10 17.2341
R86 plus.n47 plus.n46 17.2341
R87 plus plus.n35 13.4399
R88 plus.n34 plus.n33 9.49444
R89 plus.n70 plus.n69 9.49444
R90 plus.n25 plus.n24 6.57323
R91 plus.n19 plus.n18 6.57323
R92 plus.n61 plus.n60 6.57323
R93 plus.n55 plus.n54 6.57323
R94 plus.n30 plus.n3 3.65202
R95 plus.n13 plus.n8 3.65202
R96 plus.n66 plus.n39 3.65202
R97 plus.n49 plus.n44 3.65202
R98 plus.n22 plus.n21 0.380177
R99 plus.n2 plus.n1 0.380177
R100 plus.n38 plus.n37 0.380177
R101 plus.n58 plus.n57 0.380177
R102 plus.n14 plus.n9 0.285035
R103 plus.n21 plus.n6 0.285035
R104 plus.n23 plus.n22 0.285035
R105 plus.n29 plus.n2 0.285035
R106 plus.n1 plus.n0 0.285035
R107 plus.n37 plus.n36 0.285035
R108 plus.n65 plus.n38 0.285035
R109 plus.n59 plus.n58 0.285035
R110 plus.n57 plus.n42 0.285035
R111 plus.n50 plus.n45 0.285035
R112 plus.n15 plus.n14 0.189894
R113 plus.n16 plus.n15 0.189894
R114 plus.n16 plus.n7 0.189894
R115 plus.n7 plus.n6 0.189894
R116 plus.n23 plus.n4 0.189894
R117 plus.n27 plus.n4 0.189894
R118 plus.n28 plus.n27 0.189894
R119 plus.n29 plus.n28 0.189894
R120 plus.n35 plus.n0 0.189894
R121 plus.n71 plus.n36 0.189894
R122 plus.n65 plus.n64 0.189894
R123 plus.n64 plus.n63 0.189894
R124 plus.n63 plus.n40 0.189894
R125 plus.n59 plus.n40 0.189894
R126 plus.n43 plus.n42 0.189894
R127 plus.n52 plus.n43 0.189894
R128 plus.n52 plus.n51 0.189894
R129 plus.n51 plus.n50 0.189894
R130 drain_left.n13 drain_left.n11 61.8539
R131 drain_left.n7 drain_left.n5 61.8537
R132 drain_left.n2 drain_left.n0 61.8537
R133 drain_left.n19 drain_left.n18 60.8798
R134 drain_left.n17 drain_left.n16 60.8798
R135 drain_left.n15 drain_left.n14 60.8798
R136 drain_left.n13 drain_left.n12 60.8798
R137 drain_left.n21 drain_left.n20 60.8796
R138 drain_left.n7 drain_left.n6 60.8796
R139 drain_left.n9 drain_left.n8 60.8796
R140 drain_left.n4 drain_left.n3 60.8796
R141 drain_left.n2 drain_left.n1 60.8796
R142 drain_left drain_left.n10 38.8941
R143 drain_left drain_left.n21 6.62735
R144 drain_left.n5 drain_left.t12 1.3205
R145 drain_left.n5 drain_left.t2 1.3205
R146 drain_left.n6 drain_left.t10 1.3205
R147 drain_left.n6 drain_left.t22 1.3205
R148 drain_left.n8 drain_left.t1 1.3205
R149 drain_left.n8 drain_left.t18 1.3205
R150 drain_left.n3 drain_left.t15 1.3205
R151 drain_left.n3 drain_left.t14 1.3205
R152 drain_left.n1 drain_left.t19 1.3205
R153 drain_left.n1 drain_left.t11 1.3205
R154 drain_left.n0 drain_left.t16 1.3205
R155 drain_left.n0 drain_left.t4 1.3205
R156 drain_left.n20 drain_left.t5 1.3205
R157 drain_left.n20 drain_left.t6 1.3205
R158 drain_left.n18 drain_left.t3 1.3205
R159 drain_left.n18 drain_left.t9 1.3205
R160 drain_left.n16 drain_left.t21 1.3205
R161 drain_left.n16 drain_left.t13 1.3205
R162 drain_left.n14 drain_left.t17 1.3205
R163 drain_left.n14 drain_left.t20 1.3205
R164 drain_left.n12 drain_left.t7 1.3205
R165 drain_left.n12 drain_left.t8 1.3205
R166 drain_left.n11 drain_left.t0 1.3205
R167 drain_left.n11 drain_left.t23 1.3205
R168 drain_left.n9 drain_left.n7 0.974638
R169 drain_left.n4 drain_left.n2 0.974638
R170 drain_left.n15 drain_left.n13 0.974638
R171 drain_left.n17 drain_left.n15 0.974638
R172 drain_left.n19 drain_left.n17 0.974638
R173 drain_left.n21 drain_left.n19 0.974638
R174 drain_left.n10 drain_left.n9 0.432223
R175 drain_left.n10 drain_left.n4 0.432223
R176 source.n11 source.t19 45.521
R177 source.n12 source.t43 45.521
R178 source.n23 source.t2 45.521
R179 source.n47 source.t3 45.5208
R180 source.n36 source.t11 45.5208
R181 source.n35 source.t41 45.5208
R182 source.n24 source.t39 45.5208
R183 source.n0 source.t37 45.5208
R184 source.n2 source.n1 44.201
R185 source.n4 source.n3 44.201
R186 source.n6 source.n5 44.201
R187 source.n8 source.n7 44.201
R188 source.n10 source.n9 44.201
R189 source.n14 source.n13 44.201
R190 source.n16 source.n15 44.201
R191 source.n18 source.n17 44.201
R192 source.n20 source.n19 44.201
R193 source.n22 source.n21 44.201
R194 source.n46 source.n45 44.2008
R195 source.n44 source.n43 44.2008
R196 source.n42 source.n41 44.2008
R197 source.n40 source.n39 44.2008
R198 source.n38 source.n37 44.2008
R199 source.n34 source.n33 44.2008
R200 source.n32 source.n31 44.2008
R201 source.n30 source.n29 44.2008
R202 source.n28 source.n27 44.2008
R203 source.n26 source.n25 44.2008
R204 source.n24 source.n23 24.5346
R205 source.n48 source.n0 18.7846
R206 source.n48 source.n47 5.7505
R207 source.n45 source.t4 1.3205
R208 source.n45 source.t5 1.3205
R209 source.n43 source.t46 1.3205
R210 source.n43 source.t1 1.3205
R211 source.n41 source.t45 1.3205
R212 source.n41 source.t12 1.3205
R213 source.n39 source.t6 1.3205
R214 source.n39 source.t0 1.3205
R215 source.n37 source.t18 1.3205
R216 source.n37 source.t14 1.3205
R217 source.n33 source.t20 1.3205
R218 source.n33 source.t33 1.3205
R219 source.n31 source.t23 1.3205
R220 source.n31 source.t35 1.3205
R221 source.n29 source.t29 1.3205
R222 source.n29 source.t40 1.3205
R223 source.n27 source.t32 1.3205
R224 source.n27 source.t38 1.3205
R225 source.n25 source.t31 1.3205
R226 source.n25 source.t42 1.3205
R227 source.n1 source.t34 1.3205
R228 source.n1 source.t36 1.3205
R229 source.n3 source.t28 1.3205
R230 source.n3 source.t30 1.3205
R231 source.n5 source.t26 1.3205
R232 source.n5 source.t27 1.3205
R233 source.n7 source.t25 1.3205
R234 source.n7 source.t22 1.3205
R235 source.n9 source.t21 1.3205
R236 source.n9 source.t24 1.3205
R237 source.n13 source.t15 1.3205
R238 source.n13 source.t9 1.3205
R239 source.n15 source.t13 1.3205
R240 source.n15 source.t44 1.3205
R241 source.n17 source.t8 1.3205
R242 source.n17 source.t16 1.3205
R243 source.n19 source.t7 1.3205
R244 source.n19 source.t47 1.3205
R245 source.n21 source.t10 1.3205
R246 source.n21 source.t17 1.3205
R247 source.n23 source.n22 0.974638
R248 source.n22 source.n20 0.974638
R249 source.n20 source.n18 0.974638
R250 source.n18 source.n16 0.974638
R251 source.n16 source.n14 0.974638
R252 source.n14 source.n12 0.974638
R253 source.n11 source.n10 0.974638
R254 source.n10 source.n8 0.974638
R255 source.n8 source.n6 0.974638
R256 source.n6 source.n4 0.974638
R257 source.n4 source.n2 0.974638
R258 source.n2 source.n0 0.974638
R259 source.n26 source.n24 0.974638
R260 source.n28 source.n26 0.974638
R261 source.n30 source.n28 0.974638
R262 source.n32 source.n30 0.974638
R263 source.n34 source.n32 0.974638
R264 source.n35 source.n34 0.974638
R265 source.n38 source.n36 0.974638
R266 source.n40 source.n38 0.974638
R267 source.n42 source.n40 0.974638
R268 source.n44 source.n42 0.974638
R269 source.n46 source.n44 0.974638
R270 source.n47 source.n46 0.974638
R271 source.n12 source.n11 0.470328
R272 source.n36 source.n35 0.470328
R273 source source.n48 0.188
R274 minus.n8 minus.t14 522.415
R275 minus.n44 minus.t2 522.415
R276 minus.n9 minus.t10 500.979
R277 minus.n10 minus.t7 500.979
R278 minus.n14 minus.t17 500.979
R279 minus.n16 minus.t19 500.979
R280 minus.n20 minus.t15 500.979
R281 minus.n21 minus.t12 500.979
R282 minus.n3 minus.t20 500.979
R283 minus.n27 minus.t18 500.979
R284 minus.n1 minus.t6 500.979
R285 minus.n32 minus.t13 500.979
R286 minus.n34 minus.t11 500.979
R287 minus.n45 minus.t16 500.979
R288 minus.n46 minus.t22 500.979
R289 minus.n50 minus.t8 500.979
R290 minus.n52 minus.t1 500.979
R291 minus.n56 minus.t5 500.979
R292 minus.n57 minus.t21 500.979
R293 minus.n39 minus.t3 500.979
R294 minus.n63 minus.t23 500.979
R295 minus.n37 minus.t4 500.979
R296 minus.n68 minus.t9 500.979
R297 minus.n70 minus.t0 500.979
R298 minus.n35 minus.n34 161.3
R299 minus.n33 minus.n0 161.3
R300 minus.n29 minus.n28 161.3
R301 minus.n27 minus.n2 161.3
R302 minus.n26 minus.n25 161.3
R303 minus.n24 minus.n3 161.3
R304 minus.n23 minus.n22 161.3
R305 minus.n18 minus.n5 161.3
R306 minus.n17 minus.n16 161.3
R307 minus.n15 minus.n6 161.3
R308 minus.n14 minus.n13 161.3
R309 minus.n12 minus.n7 161.3
R310 minus.n71 minus.n70 161.3
R311 minus.n69 minus.n36 161.3
R312 minus.n65 minus.n64 161.3
R313 minus.n63 minus.n38 161.3
R314 minus.n62 minus.n61 161.3
R315 minus.n60 minus.n39 161.3
R316 minus.n59 minus.n58 161.3
R317 minus.n54 minus.n41 161.3
R318 minus.n53 minus.n52 161.3
R319 minus.n51 minus.n42 161.3
R320 minus.n50 minus.n49 161.3
R321 minus.n48 minus.n43 161.3
R322 minus.n32 minus.n31 80.6037
R323 minus.n30 minus.n1 80.6037
R324 minus.n21 minus.n4 80.6037
R325 minus.n20 minus.n19 80.6037
R326 minus.n11 minus.n10 80.6037
R327 minus.n68 minus.n67 80.6037
R328 minus.n66 minus.n37 80.6037
R329 minus.n57 minus.n40 80.6037
R330 minus.n56 minus.n55 80.6037
R331 minus.n47 minus.n46 80.6037
R332 minus.n10 minus.n9 48.2005
R333 minus.n21 minus.n20 48.2005
R334 minus.n32 minus.n1 48.2005
R335 minus.n46 minus.n45 48.2005
R336 minus.n57 minus.n56 48.2005
R337 minus.n68 minus.n37 48.2005
R338 minus.n72 minus.n35 45.3944
R339 minus.n10 minus.n7 44.549
R340 minus.n28 minus.n1 44.549
R341 minus.n46 minus.n43 44.549
R342 minus.n64 minus.n37 44.549
R343 minus.n20 minus.n5 41.6278
R344 minus.n22 minus.n21 41.6278
R345 minus.n56 minus.n41 41.6278
R346 minus.n58 minus.n57 41.6278
R347 minus.n33 minus.n32 38.7066
R348 minus.n69 minus.n68 38.7066
R349 minus.n11 minus.n8 31.6825
R350 minus.n47 minus.n44 31.6825
R351 minus.n15 minus.n14 25.5611
R352 minus.n27 minus.n26 25.5611
R353 minus.n51 minus.n50 25.5611
R354 minus.n63 minus.n62 25.5611
R355 minus.n16 minus.n15 22.6399
R356 minus.n26 minus.n3 22.6399
R357 minus.n52 minus.n51 22.6399
R358 minus.n62 minus.n39 22.6399
R359 minus.n9 minus.n8 17.2341
R360 minus.n45 minus.n44 17.2341
R361 minus.n34 minus.n33 9.49444
R362 minus.n70 minus.n69 9.49444
R363 minus.n72 minus.n71 6.65959
R364 minus.n16 minus.n5 6.57323
R365 minus.n22 minus.n3 6.57323
R366 minus.n52 minus.n41 6.57323
R367 minus.n58 minus.n39 6.57323
R368 minus.n14 minus.n7 3.65202
R369 minus.n28 minus.n27 3.65202
R370 minus.n50 minus.n43 3.65202
R371 minus.n64 minus.n63 3.65202
R372 minus.n31 minus.n30 0.380177
R373 minus.n19 minus.n4 0.380177
R374 minus.n55 minus.n40 0.380177
R375 minus.n67 minus.n66 0.380177
R376 minus.n31 minus.n0 0.285035
R377 minus.n30 minus.n29 0.285035
R378 minus.n23 minus.n4 0.285035
R379 minus.n19 minus.n18 0.285035
R380 minus.n12 minus.n11 0.285035
R381 minus.n48 minus.n47 0.285035
R382 minus.n55 minus.n54 0.285035
R383 minus.n59 minus.n40 0.285035
R384 minus.n66 minus.n65 0.285035
R385 minus.n67 minus.n36 0.285035
R386 minus.n35 minus.n0 0.189894
R387 minus.n29 minus.n2 0.189894
R388 minus.n25 minus.n2 0.189894
R389 minus.n25 minus.n24 0.189894
R390 minus.n24 minus.n23 0.189894
R391 minus.n18 minus.n17 0.189894
R392 minus.n17 minus.n6 0.189894
R393 minus.n13 minus.n6 0.189894
R394 minus.n13 minus.n12 0.189894
R395 minus.n49 minus.n48 0.189894
R396 minus.n49 minus.n42 0.189894
R397 minus.n53 minus.n42 0.189894
R398 minus.n54 minus.n53 0.189894
R399 minus.n60 minus.n59 0.189894
R400 minus.n61 minus.n60 0.189894
R401 minus.n61 minus.n38 0.189894
R402 minus.n65 minus.n38 0.189894
R403 minus.n71 minus.n36 0.189894
R404 minus minus.n72 0.188
R405 drain_right.n13 drain_right.n11 61.8538
R406 drain_right.n7 drain_right.n5 61.8537
R407 drain_right.n2 drain_right.n0 61.8537
R408 drain_right.n13 drain_right.n12 60.8798
R409 drain_right.n15 drain_right.n14 60.8798
R410 drain_right.n17 drain_right.n16 60.8798
R411 drain_right.n19 drain_right.n18 60.8798
R412 drain_right.n21 drain_right.n20 60.8798
R413 drain_right.n7 drain_right.n6 60.8796
R414 drain_right.n9 drain_right.n8 60.8796
R415 drain_right.n4 drain_right.n3 60.8796
R416 drain_right.n2 drain_right.n1 60.8796
R417 drain_right drain_right.n10 38.3409
R418 drain_right drain_right.n21 6.62735
R419 drain_right.n5 drain_right.t14 1.3205
R420 drain_right.n5 drain_right.t23 1.3205
R421 drain_right.n6 drain_right.t0 1.3205
R422 drain_right.n6 drain_right.t19 1.3205
R423 drain_right.n8 drain_right.t2 1.3205
R424 drain_right.n8 drain_right.t20 1.3205
R425 drain_right.n3 drain_right.t22 1.3205
R426 drain_right.n3 drain_right.t18 1.3205
R427 drain_right.n1 drain_right.t1 1.3205
R428 drain_right.n1 drain_right.t15 1.3205
R429 drain_right.n0 drain_right.t21 1.3205
R430 drain_right.n0 drain_right.t7 1.3205
R431 drain_right.n11 drain_right.t13 1.3205
R432 drain_right.n11 drain_right.t9 1.3205
R433 drain_right.n12 drain_right.t6 1.3205
R434 drain_right.n12 drain_right.t16 1.3205
R435 drain_right.n14 drain_right.t8 1.3205
R436 drain_right.n14 drain_right.t4 1.3205
R437 drain_right.n16 drain_right.t3 1.3205
R438 drain_right.n16 drain_right.t11 1.3205
R439 drain_right.n18 drain_right.t17 1.3205
R440 drain_right.n18 drain_right.t5 1.3205
R441 drain_right.n20 drain_right.t12 1.3205
R442 drain_right.n20 drain_right.t10 1.3205
R443 drain_right.n9 drain_right.n7 0.974638
R444 drain_right.n4 drain_right.n2 0.974638
R445 drain_right.n21 drain_right.n19 0.974638
R446 drain_right.n19 drain_right.n17 0.974638
R447 drain_right.n17 drain_right.n15 0.974638
R448 drain_right.n15 drain_right.n13 0.974638
R449 drain_right.n10 drain_right.n9 0.432223
R450 drain_right.n10 drain_right.n4 0.432223
C0 drain_right plus 0.526806f
C1 drain_right minus 19.8877f
C2 drain_left plus 20.2552f
C3 drain_left minus 0.175388f
C4 drain_right source 31.8265f
C5 minus plus 8.26435f
C6 drain_left source 31.8234f
C7 source plus 20.189499f
C8 drain_left drain_right 2.02887f
C9 minus source 20.1754f
C10 drain_right a_n3654_n3888# 8.78523f
C11 drain_left a_n3654_n3888# 9.28933f
C12 source a_n3654_n3888# 11.418134f
C13 minus a_n3654_n3888# 15.076556f
C14 plus a_n3654_n3888# 17.05676f
C15 drain_right.t21 a_n3654_n3888# 0.326023f
C16 drain_right.t7 a_n3654_n3888# 0.326023f
C17 drain_right.n0 a_n3654_n3888# 2.95331f
C18 drain_right.t1 a_n3654_n3888# 0.326023f
C19 drain_right.t15 a_n3654_n3888# 0.326023f
C20 drain_right.n1 a_n3654_n3888# 2.94686f
C21 drain_right.n2 a_n3654_n3888# 0.800526f
C22 drain_right.t22 a_n3654_n3888# 0.326023f
C23 drain_right.t18 a_n3654_n3888# 0.326023f
C24 drain_right.n3 a_n3654_n3888# 2.94686f
C25 drain_right.n4 a_n3654_n3888# 0.35135f
C26 drain_right.t14 a_n3654_n3888# 0.326023f
C27 drain_right.t23 a_n3654_n3888# 0.326023f
C28 drain_right.n5 a_n3654_n3888# 2.95331f
C29 drain_right.t0 a_n3654_n3888# 0.326023f
C30 drain_right.t19 a_n3654_n3888# 0.326023f
C31 drain_right.n6 a_n3654_n3888# 2.94686f
C32 drain_right.n7 a_n3654_n3888# 0.800526f
C33 drain_right.t2 a_n3654_n3888# 0.326023f
C34 drain_right.t20 a_n3654_n3888# 0.326023f
C35 drain_right.n8 a_n3654_n3888# 2.94686f
C36 drain_right.n9 a_n3654_n3888# 0.35135f
C37 drain_right.n10 a_n3654_n3888# 2.03663f
C38 drain_right.t13 a_n3654_n3888# 0.326023f
C39 drain_right.t9 a_n3654_n3888# 0.326023f
C40 drain_right.n11 a_n3654_n3888# 2.9533f
C41 drain_right.t6 a_n3654_n3888# 0.326023f
C42 drain_right.t16 a_n3654_n3888# 0.326023f
C43 drain_right.n12 a_n3654_n3888# 2.94687f
C44 drain_right.n13 a_n3654_n3888# 0.800532f
C45 drain_right.t8 a_n3654_n3888# 0.326023f
C46 drain_right.t4 a_n3654_n3888# 0.326023f
C47 drain_right.n14 a_n3654_n3888# 2.94687f
C48 drain_right.n15 a_n3654_n3888# 0.397943f
C49 drain_right.t3 a_n3654_n3888# 0.326023f
C50 drain_right.t11 a_n3654_n3888# 0.326023f
C51 drain_right.n16 a_n3654_n3888# 2.94687f
C52 drain_right.n17 a_n3654_n3888# 0.397943f
C53 drain_right.t17 a_n3654_n3888# 0.326023f
C54 drain_right.t5 a_n3654_n3888# 0.326023f
C55 drain_right.n18 a_n3654_n3888# 2.94687f
C56 drain_right.n19 a_n3654_n3888# 0.397943f
C57 drain_right.t12 a_n3654_n3888# 0.326023f
C58 drain_right.t10 a_n3654_n3888# 0.326023f
C59 drain_right.n20 a_n3654_n3888# 2.94687f
C60 drain_right.n21 a_n3654_n3888# 0.644573f
C61 minus.n0 a_n3654_n3888# 0.049493f
C62 minus.t6 a_n3654_n3888# 1.26481f
C63 minus.n1 a_n3654_n3888# 0.495519f
C64 minus.t13 a_n3654_n3888# 1.26481f
C65 minus.n2 a_n3654_n3888# 0.037091f
C66 minus.t20 a_n3654_n3888# 1.26481f
C67 minus.n3 a_n3654_n3888# 0.484701f
C68 minus.n4 a_n3654_n3888# 0.061779f
C69 minus.n5 a_n3654_n3888# 0.008417f
C70 minus.t15 a_n3654_n3888# 1.26481f
C71 minus.n6 a_n3654_n3888# 0.037091f
C72 minus.n7 a_n3654_n3888# 0.008417f
C73 minus.t17 a_n3654_n3888# 1.26481f
C74 minus.t14 a_n3654_n3888# 1.28482f
C75 minus.n8 a_n3654_n3888# 0.471336f
C76 minus.t10 a_n3654_n3888# 1.26481f
C77 minus.n9 a_n3654_n3888# 0.4955f
C78 minus.t7 a_n3654_n3888# 1.26481f
C79 minus.n10 a_n3654_n3888# 0.495519f
C80 minus.n11 a_n3654_n3888# 0.213183f
C81 minus.n12 a_n3654_n3888# 0.049493f
C82 minus.n13 a_n3654_n3888# 0.037091f
C83 minus.n14 a_n3654_n3888# 0.484701f
C84 minus.n15 a_n3654_n3888# 0.008417f
C85 minus.t19 a_n3654_n3888# 1.26481f
C86 minus.n16 a_n3654_n3888# 0.484701f
C87 minus.n17 a_n3654_n3888# 0.037091f
C88 minus.n18 a_n3654_n3888# 0.049493f
C89 minus.n19 a_n3654_n3888# 0.061779f
C90 minus.n20 a_n3654_n3888# 0.495061f
C91 minus.t12 a_n3654_n3888# 1.26481f
C92 minus.n21 a_n3654_n3888# 0.495061f
C93 minus.n22 a_n3654_n3888# 0.008417f
C94 minus.n23 a_n3654_n3888# 0.049493f
C95 minus.n24 a_n3654_n3888# 0.037091f
C96 minus.n25 a_n3654_n3888# 0.037091f
C97 minus.n26 a_n3654_n3888# 0.008417f
C98 minus.t18 a_n3654_n3888# 1.26481f
C99 minus.n27 a_n3654_n3888# 0.484701f
C100 minus.n28 a_n3654_n3888# 0.008417f
C101 minus.n29 a_n3654_n3888# 0.049493f
C102 minus.n30 a_n3654_n3888# 0.061779f
C103 minus.n31 a_n3654_n3888# 0.061779f
C104 minus.n32 a_n3654_n3888# 0.494604f
C105 minus.n33 a_n3654_n3888# 0.008417f
C106 minus.t11 a_n3654_n3888# 1.26481f
C107 minus.n34 a_n3654_n3888# 0.481614f
C108 minus.n35 a_n3654_n3888# 1.84244f
C109 minus.n36 a_n3654_n3888# 0.049493f
C110 minus.t4 a_n3654_n3888# 1.26481f
C111 minus.n37 a_n3654_n3888# 0.495519f
C112 minus.n38 a_n3654_n3888# 0.037091f
C113 minus.t3 a_n3654_n3888# 1.26481f
C114 minus.n39 a_n3654_n3888# 0.484701f
C115 minus.n40 a_n3654_n3888# 0.061779f
C116 minus.n41 a_n3654_n3888# 0.008417f
C117 minus.n42 a_n3654_n3888# 0.037091f
C118 minus.n43 a_n3654_n3888# 0.008417f
C119 minus.t2 a_n3654_n3888# 1.28482f
C120 minus.n44 a_n3654_n3888# 0.471336f
C121 minus.t16 a_n3654_n3888# 1.26481f
C122 minus.n45 a_n3654_n3888# 0.4955f
C123 minus.t22 a_n3654_n3888# 1.26481f
C124 minus.n46 a_n3654_n3888# 0.495519f
C125 minus.n47 a_n3654_n3888# 0.213183f
C126 minus.n48 a_n3654_n3888# 0.049493f
C127 minus.n49 a_n3654_n3888# 0.037091f
C128 minus.t8 a_n3654_n3888# 1.26481f
C129 minus.n50 a_n3654_n3888# 0.484701f
C130 minus.n51 a_n3654_n3888# 0.008417f
C131 minus.t1 a_n3654_n3888# 1.26481f
C132 minus.n52 a_n3654_n3888# 0.484701f
C133 minus.n53 a_n3654_n3888# 0.037091f
C134 minus.n54 a_n3654_n3888# 0.049493f
C135 minus.n55 a_n3654_n3888# 0.061779f
C136 minus.t5 a_n3654_n3888# 1.26481f
C137 minus.n56 a_n3654_n3888# 0.495061f
C138 minus.t21 a_n3654_n3888# 1.26481f
C139 minus.n57 a_n3654_n3888# 0.495061f
C140 minus.n58 a_n3654_n3888# 0.008417f
C141 minus.n59 a_n3654_n3888# 0.049493f
C142 minus.n60 a_n3654_n3888# 0.037091f
C143 minus.n61 a_n3654_n3888# 0.037091f
C144 minus.n62 a_n3654_n3888# 0.008417f
C145 minus.t23 a_n3654_n3888# 1.26481f
C146 minus.n63 a_n3654_n3888# 0.484701f
C147 minus.n64 a_n3654_n3888# 0.008417f
C148 minus.n65 a_n3654_n3888# 0.049493f
C149 minus.n66 a_n3654_n3888# 0.061779f
C150 minus.n67 a_n3654_n3888# 0.061779f
C151 minus.t9 a_n3654_n3888# 1.26481f
C152 minus.n68 a_n3654_n3888# 0.494604f
C153 minus.n69 a_n3654_n3888# 0.008417f
C154 minus.t0 a_n3654_n3888# 1.26481f
C155 minus.n70 a_n3654_n3888# 0.481614f
C156 minus.n71 a_n3654_n3888# 0.256331f
C157 minus.n72 a_n3654_n3888# 2.17699f
C158 source.t37 a_n3654_n3888# 3.18288f
C159 source.n0 a_n3654_n3888# 1.52788f
C160 source.t34 a_n3654_n3888# 0.284018f
C161 source.t36 a_n3654_n3888# 0.284018f
C162 source.n1 a_n3654_n3888# 2.49486f
C163 source.n2 a_n3654_n3888# 0.386437f
C164 source.t28 a_n3654_n3888# 0.284018f
C165 source.t30 a_n3654_n3888# 0.284018f
C166 source.n3 a_n3654_n3888# 2.49486f
C167 source.n4 a_n3654_n3888# 0.386437f
C168 source.t26 a_n3654_n3888# 0.284018f
C169 source.t27 a_n3654_n3888# 0.284018f
C170 source.n5 a_n3654_n3888# 2.49486f
C171 source.n6 a_n3654_n3888# 0.386437f
C172 source.t25 a_n3654_n3888# 0.284018f
C173 source.t22 a_n3654_n3888# 0.284018f
C174 source.n7 a_n3654_n3888# 2.49486f
C175 source.n8 a_n3654_n3888# 0.386437f
C176 source.t21 a_n3654_n3888# 0.284018f
C177 source.t24 a_n3654_n3888# 0.284018f
C178 source.n9 a_n3654_n3888# 2.49486f
C179 source.n10 a_n3654_n3888# 0.386437f
C180 source.t19 a_n3654_n3888# 3.18288f
C181 source.n11 a_n3654_n3888# 0.434072f
C182 source.t43 a_n3654_n3888# 3.18288f
C183 source.n12 a_n3654_n3888# 0.434072f
C184 source.t15 a_n3654_n3888# 0.284018f
C185 source.t9 a_n3654_n3888# 0.284018f
C186 source.n13 a_n3654_n3888# 2.49486f
C187 source.n14 a_n3654_n3888# 0.386437f
C188 source.t13 a_n3654_n3888# 0.284018f
C189 source.t44 a_n3654_n3888# 0.284018f
C190 source.n15 a_n3654_n3888# 2.49486f
C191 source.n16 a_n3654_n3888# 0.386437f
C192 source.t8 a_n3654_n3888# 0.284018f
C193 source.t16 a_n3654_n3888# 0.284018f
C194 source.n17 a_n3654_n3888# 2.49486f
C195 source.n18 a_n3654_n3888# 0.386437f
C196 source.t7 a_n3654_n3888# 0.284018f
C197 source.t47 a_n3654_n3888# 0.284018f
C198 source.n19 a_n3654_n3888# 2.49486f
C199 source.n20 a_n3654_n3888# 0.386437f
C200 source.t10 a_n3654_n3888# 0.284018f
C201 source.t17 a_n3654_n3888# 0.284018f
C202 source.n21 a_n3654_n3888# 2.49486f
C203 source.n22 a_n3654_n3888# 0.386437f
C204 source.t2 a_n3654_n3888# 3.18288f
C205 source.n23 a_n3654_n3888# 1.93917f
C206 source.t39 a_n3654_n3888# 3.18288f
C207 source.n24 a_n3654_n3888# 1.93917f
C208 source.t31 a_n3654_n3888# 0.284018f
C209 source.t42 a_n3654_n3888# 0.284018f
C210 source.n25 a_n3654_n3888# 2.49485f
C211 source.n26 a_n3654_n3888# 0.38644f
C212 source.t32 a_n3654_n3888# 0.284018f
C213 source.t38 a_n3654_n3888# 0.284018f
C214 source.n27 a_n3654_n3888# 2.49485f
C215 source.n28 a_n3654_n3888# 0.38644f
C216 source.t29 a_n3654_n3888# 0.284018f
C217 source.t40 a_n3654_n3888# 0.284018f
C218 source.n29 a_n3654_n3888# 2.49485f
C219 source.n30 a_n3654_n3888# 0.38644f
C220 source.t23 a_n3654_n3888# 0.284018f
C221 source.t35 a_n3654_n3888# 0.284018f
C222 source.n31 a_n3654_n3888# 2.49485f
C223 source.n32 a_n3654_n3888# 0.38644f
C224 source.t20 a_n3654_n3888# 0.284018f
C225 source.t33 a_n3654_n3888# 0.284018f
C226 source.n33 a_n3654_n3888# 2.49485f
C227 source.n34 a_n3654_n3888# 0.38644f
C228 source.t41 a_n3654_n3888# 3.18288f
C229 source.n35 a_n3654_n3888# 0.434076f
C230 source.t11 a_n3654_n3888# 3.18288f
C231 source.n36 a_n3654_n3888# 0.434076f
C232 source.t18 a_n3654_n3888# 0.284018f
C233 source.t14 a_n3654_n3888# 0.284018f
C234 source.n37 a_n3654_n3888# 2.49485f
C235 source.n38 a_n3654_n3888# 0.38644f
C236 source.t6 a_n3654_n3888# 0.284018f
C237 source.t0 a_n3654_n3888# 0.284018f
C238 source.n39 a_n3654_n3888# 2.49485f
C239 source.n40 a_n3654_n3888# 0.38644f
C240 source.t45 a_n3654_n3888# 0.284018f
C241 source.t12 a_n3654_n3888# 0.284018f
C242 source.n41 a_n3654_n3888# 2.49485f
C243 source.n42 a_n3654_n3888# 0.38644f
C244 source.t46 a_n3654_n3888# 0.284018f
C245 source.t1 a_n3654_n3888# 0.284018f
C246 source.n43 a_n3654_n3888# 2.49485f
C247 source.n44 a_n3654_n3888# 0.38644f
C248 source.t4 a_n3654_n3888# 0.284018f
C249 source.t5 a_n3654_n3888# 0.284018f
C250 source.n45 a_n3654_n3888# 2.49485f
C251 source.n46 a_n3654_n3888# 0.38644f
C252 source.t3 a_n3654_n3888# 3.18288f
C253 source.n47 a_n3654_n3888# 0.59556f
C254 source.n48 a_n3654_n3888# 1.77195f
C255 drain_left.t16 a_n3654_n3888# 0.327795f
C256 drain_left.t4 a_n3654_n3888# 0.327795f
C257 drain_left.n0 a_n3654_n3888# 2.96936f
C258 drain_left.t19 a_n3654_n3888# 0.327795f
C259 drain_left.t11 a_n3654_n3888# 0.327795f
C260 drain_left.n1 a_n3654_n3888# 2.96288f
C261 drain_left.n2 a_n3654_n3888# 0.804877f
C262 drain_left.t15 a_n3654_n3888# 0.327795f
C263 drain_left.t14 a_n3654_n3888# 0.327795f
C264 drain_left.n3 a_n3654_n3888# 2.96288f
C265 drain_left.n4 a_n3654_n3888# 0.35326f
C266 drain_left.t12 a_n3654_n3888# 0.327795f
C267 drain_left.t2 a_n3654_n3888# 0.327795f
C268 drain_left.n5 a_n3654_n3888# 2.96936f
C269 drain_left.t10 a_n3654_n3888# 0.327795f
C270 drain_left.t22 a_n3654_n3888# 0.327795f
C271 drain_left.n6 a_n3654_n3888# 2.96288f
C272 drain_left.n7 a_n3654_n3888# 0.804877f
C273 drain_left.t1 a_n3654_n3888# 0.327795f
C274 drain_left.t18 a_n3654_n3888# 0.327795f
C275 drain_left.n8 a_n3654_n3888# 2.96288f
C276 drain_left.n9 a_n3654_n3888# 0.35326f
C277 drain_left.n10 a_n3654_n3888# 2.10375f
C278 drain_left.t0 a_n3654_n3888# 0.327795f
C279 drain_left.t23 a_n3654_n3888# 0.327795f
C280 drain_left.n11 a_n3654_n3888# 2.96936f
C281 drain_left.t7 a_n3654_n3888# 0.327795f
C282 drain_left.t8 a_n3654_n3888# 0.327795f
C283 drain_left.n12 a_n3654_n3888# 2.96288f
C284 drain_left.n13 a_n3654_n3888# 0.804872f
C285 drain_left.t17 a_n3654_n3888# 0.327795f
C286 drain_left.t20 a_n3654_n3888# 0.327795f
C287 drain_left.n14 a_n3654_n3888# 2.96288f
C288 drain_left.n15 a_n3654_n3888# 0.400105f
C289 drain_left.t21 a_n3654_n3888# 0.327795f
C290 drain_left.t13 a_n3654_n3888# 0.327795f
C291 drain_left.n16 a_n3654_n3888# 2.96288f
C292 drain_left.n17 a_n3654_n3888# 0.400105f
C293 drain_left.t3 a_n3654_n3888# 0.327795f
C294 drain_left.t9 a_n3654_n3888# 0.327795f
C295 drain_left.n18 a_n3654_n3888# 2.96288f
C296 drain_left.n19 a_n3654_n3888# 0.400105f
C297 drain_left.t5 a_n3654_n3888# 0.327795f
C298 drain_left.t6 a_n3654_n3888# 0.327795f
C299 drain_left.n20 a_n3654_n3888# 2.96287f
C300 drain_left.n21 a_n3654_n3888# 0.648087f
C301 plus.n0 a_n3654_n3888# 0.049979f
C302 plus.t5 a_n3654_n3888# 1.27724f
C303 plus.t6 a_n3654_n3888# 1.27724f
C304 plus.n1 a_n3654_n3888# 0.062386f
C305 plus.t8 a_n3654_n3888# 1.27724f
C306 plus.n2 a_n3654_n3888# 0.062386f
C307 plus.t12 a_n3654_n3888# 1.27724f
C308 plus.n3 a_n3654_n3888# 0.489465f
C309 plus.n4 a_n3654_n3888# 0.037455f
C310 plus.t14 a_n3654_n3888# 1.27724f
C311 plus.t15 a_n3654_n3888# 1.27724f
C312 plus.n5 a_n3654_n3888# 0.499928f
C313 plus.n6 a_n3654_n3888# 0.049979f
C314 plus.t16 a_n3654_n3888# 1.27724f
C315 plus.t20 a_n3654_n3888# 1.27724f
C316 plus.n7 a_n3654_n3888# 0.037455f
C317 plus.t17 a_n3654_n3888# 1.27724f
C318 plus.n8 a_n3654_n3888# 0.489465f
C319 plus.n9 a_n3654_n3888# 0.215279f
C320 plus.t18 a_n3654_n3888# 1.27724f
C321 plus.t21 a_n3654_n3888# 1.27724f
C322 plus.t23 a_n3654_n3888# 1.29745f
C323 plus.n10 a_n3654_n3888# 0.475969f
C324 plus.n11 a_n3654_n3888# 0.50037f
C325 plus.n12 a_n3654_n3888# 0.500389f
C326 plus.n13 a_n3654_n3888# 0.008499f
C327 plus.n14 a_n3654_n3888# 0.049979f
C328 plus.n15 a_n3654_n3888# 0.037455f
C329 plus.n16 a_n3654_n3888# 0.037455f
C330 plus.n17 a_n3654_n3888# 0.008499f
C331 plus.n18 a_n3654_n3888# 0.489465f
C332 plus.n19 a_n3654_n3888# 0.008499f
C333 plus.n20 a_n3654_n3888# 0.499928f
C334 plus.n21 a_n3654_n3888# 0.062386f
C335 plus.n22 a_n3654_n3888# 0.062386f
C336 plus.n23 a_n3654_n3888# 0.049979f
C337 plus.n24 a_n3654_n3888# 0.008499f
C338 plus.n25 a_n3654_n3888# 0.489465f
C339 plus.n26 a_n3654_n3888# 0.008499f
C340 plus.n27 a_n3654_n3888# 0.037455f
C341 plus.n28 a_n3654_n3888# 0.037455f
C342 plus.n29 a_n3654_n3888# 0.049979f
C343 plus.n30 a_n3654_n3888# 0.008499f
C344 plus.n31 a_n3654_n3888# 0.500389f
C345 plus.n32 a_n3654_n3888# 0.499466f
C346 plus.n33 a_n3654_n3888# 0.008499f
C347 plus.n34 a_n3654_n3888# 0.486348f
C348 plus.n35 a_n3654_n3888# 0.487346f
C349 plus.n36 a_n3654_n3888# 0.049979f
C350 plus.t3 a_n3654_n3888# 1.27724f
C351 plus.n37 a_n3654_n3888# 0.062386f
C352 plus.t11 a_n3654_n3888# 1.27724f
C353 plus.n38 a_n3654_n3888# 0.062386f
C354 plus.t0 a_n3654_n3888# 1.27724f
C355 plus.t10 a_n3654_n3888# 1.27724f
C356 plus.n39 a_n3654_n3888# 0.489465f
C357 plus.n40 a_n3654_n3888# 0.037455f
C358 plus.t4 a_n3654_n3888# 1.27724f
C359 plus.t13 a_n3654_n3888# 1.27724f
C360 plus.n41 a_n3654_n3888# 0.499928f
C361 plus.n42 a_n3654_n3888# 0.049979f
C362 plus.t2 a_n3654_n3888# 1.27724f
C363 plus.n43 a_n3654_n3888# 0.037455f
C364 plus.t19 a_n3654_n3888# 1.27724f
C365 plus.t7 a_n3654_n3888# 1.27724f
C366 plus.n44 a_n3654_n3888# 0.489465f
C367 plus.n45 a_n3654_n3888# 0.215279f
C368 plus.t22 a_n3654_n3888# 1.27724f
C369 plus.t1 a_n3654_n3888# 1.29745f
C370 plus.n46 a_n3654_n3888# 0.475969f
C371 plus.t9 a_n3654_n3888# 1.27724f
C372 plus.n47 a_n3654_n3888# 0.50037f
C373 plus.n48 a_n3654_n3888# 0.500389f
C374 plus.n49 a_n3654_n3888# 0.008499f
C375 plus.n50 a_n3654_n3888# 0.049979f
C376 plus.n51 a_n3654_n3888# 0.037455f
C377 plus.n52 a_n3654_n3888# 0.037455f
C378 plus.n53 a_n3654_n3888# 0.008499f
C379 plus.n54 a_n3654_n3888# 0.489465f
C380 plus.n55 a_n3654_n3888# 0.008499f
C381 plus.n56 a_n3654_n3888# 0.499928f
C382 plus.n57 a_n3654_n3888# 0.062386f
C383 plus.n58 a_n3654_n3888# 0.062386f
C384 plus.n59 a_n3654_n3888# 0.049979f
C385 plus.n60 a_n3654_n3888# 0.008499f
C386 plus.n61 a_n3654_n3888# 0.489465f
C387 plus.n62 a_n3654_n3888# 0.008499f
C388 plus.n63 a_n3654_n3888# 0.037455f
C389 plus.n64 a_n3654_n3888# 0.037455f
C390 plus.n65 a_n3654_n3888# 0.049979f
C391 plus.n66 a_n3654_n3888# 0.008499f
C392 plus.n67 a_n3654_n3888# 0.500389f
C393 plus.n68 a_n3654_n3888# 0.499466f
C394 plus.n69 a_n3654_n3888# 0.008499f
C395 plus.n70 a_n3654_n3888# 0.486348f
C396 plus.n71 a_n3654_n3888# 1.56644f
.ends

