* NGSPICE file created from diffpair385.ext - technology: sky130A

.subckt diffpair385 minus drain_right drain_left source plus
X0 source.t17 plus.t0 drain_left.t5 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X1 source.t19 minus.t0 drain_right.t11 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X2 source.t16 plus.t1 drain_left.t10 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X3 source.t15 plus.t2 drain_left.t2 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X4 source.t14 plus.t3 drain_left.t7 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X5 drain_left.t11 plus.t4 source.t13 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X6 drain_right.t10 minus.t1 source.t20 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X7 drain_left.t3 plus.t5 source.t12 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X8 drain_right.t9 minus.t2 source.t21 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X9 drain_left.t0 plus.t6 source.t11 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X10 a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X11 drain_left.t6 plus.t7 source.t10 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X12 drain_right.t8 minus.t3 source.t22 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X13 a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X14 drain_right.t7 minus.t4 source.t1 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X15 drain_left.t4 plus.t8 source.t9 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X16 drain_left.t1 plus.t9 source.t8 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X17 source.t23 minus.t5 drain_right.t6 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X18 source.t7 plus.t10 drain_left.t9 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X19 drain_right.t5 minus.t6 source.t3 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X20 a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X21 source.t18 minus.t7 drain_right.t4 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X22 source.t6 plus.t11 drain_left.t8 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X23 source.t2 minus.t8 drain_right.t3 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X24 source.t0 minus.t9 drain_right.t2 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X25 a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X26 drain_right.t1 minus.t10 source.t4 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X27 source.t5 minus.t11 drain_right.t0 a_n2158_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
R0 plus.n5 plus.t2 389.281
R1 plus.n23 plus.t9 389.281
R2 plus.n16 plus.t7 365.976
R3 plus.n14 plus.t1 365.976
R4 plus.n2 plus.t6 365.976
R5 plus.n8 plus.t0 365.976
R6 plus.n4 plus.t8 365.976
R7 plus.n34 plus.t11 365.976
R8 plus.n32 plus.t4 365.976
R9 plus.n20 plus.t3 365.976
R10 plus.n26 plus.t5 365.976
R11 plus.n22 plus.t10 365.976
R12 plus.n7 plus.n6 161.3
R13 plus.n8 plus.n3 161.3
R14 plus.n10 plus.n9 161.3
R15 plus.n11 plus.n2 161.3
R16 plus.n13 plus.n12 161.3
R17 plus.n14 plus.n1 161.3
R18 plus.n15 plus.n0 161.3
R19 plus.n17 plus.n16 161.3
R20 plus.n25 plus.n24 161.3
R21 plus.n26 plus.n21 161.3
R22 plus.n28 plus.n27 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus.n16 plus.n15 32.8641
R31 plus.n34 plus.n33 32.8641
R32 plus plus.n35 30.1846
R33 plus.n14 plus.n13 28.4823
R34 plus.n7 plus.n4 28.4823
R35 plus.n32 plus.n31 28.4823
R36 plus.n25 plus.n22 28.4823
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 11.152
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 drain_left.n6 drain_left.n4 66.4255
R65 drain_left.n3 drain_left.n2 66.3699
R66 drain_left.n3 drain_left.n0 66.3699
R67 drain_left.n6 drain_left.n5 65.5376
R68 drain_left.n8 drain_left.n7 65.5374
R69 drain_left.n3 drain_left.n1 65.5373
R70 drain_left drain_left.n3 29.534
R71 drain_left drain_left.n8 6.54115
R72 drain_left.n1 drain_left.t7 2.2005
R73 drain_left.n1 drain_left.t3 2.2005
R74 drain_left.n2 drain_left.t9 2.2005
R75 drain_left.n2 drain_left.t1 2.2005
R76 drain_left.n0 drain_left.t8 2.2005
R77 drain_left.n0 drain_left.t11 2.2005
R78 drain_left.n7 drain_left.t10 2.2005
R79 drain_left.n7 drain_left.t6 2.2005
R80 drain_left.n5 drain_left.t5 2.2005
R81 drain_left.n5 drain_left.t0 2.2005
R82 drain_left.n4 drain_left.t2 2.2005
R83 drain_left.n4 drain_left.t4 2.2005
R84 drain_left.n8 drain_left.n6 0.888431
R85 source.n5 source.t15 51.0588
R86 source.n6 source.t1 51.0588
R87 source.n11 source.t0 51.0588
R88 source.n23 source.t22 51.0586
R89 source.n18 source.t5 51.0586
R90 source.n17 source.t8 51.0586
R91 source.n12 source.t6 51.0586
R92 source.n0 source.t10 51.0586
R93 source.n2 source.n1 48.8588
R94 source.n4 source.n3 48.8588
R95 source.n8 source.n7 48.8588
R96 source.n10 source.n9 48.8588
R97 source.n22 source.n21 48.8586
R98 source.n20 source.n19 48.8586
R99 source.n16 source.n15 48.8586
R100 source.n14 source.n13 48.8586
R101 source.n12 source.n11 19.9029
R102 source.n24 source.n0 14.196
R103 source.n24 source.n23 5.7074
R104 source.n21 source.t3 2.2005
R105 source.n21 source.t18 2.2005
R106 source.n19 source.t4 2.2005
R107 source.n19 source.t23 2.2005
R108 source.n15 source.t12 2.2005
R109 source.n15 source.t7 2.2005
R110 source.n13 source.t13 2.2005
R111 source.n13 source.t14 2.2005
R112 source.n1 source.t11 2.2005
R113 source.n1 source.t16 2.2005
R114 source.n3 source.t9 2.2005
R115 source.n3 source.t17 2.2005
R116 source.n7 source.t21 2.2005
R117 source.n7 source.t19 2.2005
R118 source.n9 source.t20 2.2005
R119 source.n9 source.t2 2.2005
R120 source.n11 source.n10 0.888431
R121 source.n10 source.n8 0.888431
R122 source.n8 source.n6 0.888431
R123 source.n5 source.n4 0.888431
R124 source.n4 source.n2 0.888431
R125 source.n2 source.n0 0.888431
R126 source.n14 source.n12 0.888431
R127 source.n16 source.n14 0.888431
R128 source.n17 source.n16 0.888431
R129 source.n20 source.n18 0.888431
R130 source.n22 source.n20 0.888431
R131 source.n23 source.n22 0.888431
R132 source.n6 source.n5 0.470328
R133 source.n18 source.n17 0.470328
R134 source source.n24 0.188
R135 minus.n5 minus.t4 389.281
R136 minus.n23 minus.t11 389.281
R137 minus.n4 minus.t0 365.976
R138 minus.n8 minus.t2 365.976
R139 minus.n10 minus.t8 365.976
R140 minus.n14 minus.t1 365.976
R141 minus.n16 minus.t9 365.976
R142 minus.n22 minus.t10 365.976
R143 minus.n26 minus.t5 365.976
R144 minus.n28 minus.t6 365.976
R145 minus.n32 minus.t7 365.976
R146 minus.n34 minus.t3 365.976
R147 minus.n17 minus.n16 161.3
R148 minus.n15 minus.n0 161.3
R149 minus.n14 minus.n13 161.3
R150 minus.n12 minus.n1 161.3
R151 minus.n11 minus.n10 161.3
R152 minus.n9 minus.n2 161.3
R153 minus.n8 minus.n7 161.3
R154 minus.n6 minus.n3 161.3
R155 minus.n35 minus.n34 161.3
R156 minus.n33 minus.n18 161.3
R157 minus.n32 minus.n31 161.3
R158 minus.n30 minus.n19 161.3
R159 minus.n29 minus.n28 161.3
R160 minus.n27 minus.n20 161.3
R161 minus.n26 minus.n25 161.3
R162 minus.n24 minus.n21 161.3
R163 minus.n6 minus.n5 44.8907
R164 minus.n24 minus.n23 44.8907
R165 minus.n36 minus.n17 35.1672
R166 minus.n16 minus.n15 32.8641
R167 minus.n34 minus.n33 32.8641
R168 minus.n4 minus.n3 28.4823
R169 minus.n14 minus.n1 28.4823
R170 minus.n22 minus.n21 28.4823
R171 minus.n32 minus.n19 28.4823
R172 minus.n10 minus.n9 24.1005
R173 minus.n9 minus.n8 24.1005
R174 minus.n27 minus.n26 24.1005
R175 minus.n28 minus.n27 24.1005
R176 minus.n8 minus.n3 19.7187
R177 minus.n10 minus.n1 19.7187
R178 minus.n26 minus.n21 19.7187
R179 minus.n28 minus.n19 19.7187
R180 minus.n5 minus.n4 18.4104
R181 minus.n23 minus.n22 18.4104
R182 minus.n15 minus.n14 15.3369
R183 minus.n33 minus.n32 15.3369
R184 minus.n36 minus.n35 6.64444
R185 minus.n17 minus.n0 0.189894
R186 minus.n13 minus.n0 0.189894
R187 minus.n13 minus.n12 0.189894
R188 minus.n12 minus.n11 0.189894
R189 minus.n11 minus.n2 0.189894
R190 minus.n7 minus.n2 0.189894
R191 minus.n7 minus.n6 0.189894
R192 minus.n25 minus.n24 0.189894
R193 minus.n25 minus.n20 0.189894
R194 minus.n29 minus.n20 0.189894
R195 minus.n30 minus.n29 0.189894
R196 minus.n31 minus.n30 0.189894
R197 minus.n31 minus.n18 0.189894
R198 minus.n35 minus.n18 0.189894
R199 minus minus.n36 0.188
R200 drain_right.n6 drain_right.n4 66.4254
R201 drain_right.n3 drain_right.n2 66.3699
R202 drain_right.n3 drain_right.n0 66.3699
R203 drain_right.n6 drain_right.n5 65.5376
R204 drain_right.n8 drain_right.n7 65.5376
R205 drain_right.n3 drain_right.n1 65.5373
R206 drain_right drain_right.n3 28.9808
R207 drain_right drain_right.n8 6.54115
R208 drain_right.n1 drain_right.t6 2.2005
R209 drain_right.n1 drain_right.t5 2.2005
R210 drain_right.n2 drain_right.t4 2.2005
R211 drain_right.n2 drain_right.t8 2.2005
R212 drain_right.n0 drain_right.t0 2.2005
R213 drain_right.n0 drain_right.t1 2.2005
R214 drain_right.n4 drain_right.t11 2.2005
R215 drain_right.n4 drain_right.t7 2.2005
R216 drain_right.n5 drain_right.t3 2.2005
R217 drain_right.n5 drain_right.t9 2.2005
R218 drain_right.n7 drain_right.t2 2.2005
R219 drain_right.n7 drain_right.t10 2.2005
R220 drain_right.n8 drain_right.n6 0.888431
C0 source drain_right 12.3341f
C1 minus plus 5.27923f
C2 drain_left drain_right 1.08491f
C3 source plus 6.0616f
C4 drain_left plus 6.24949f
C5 minus source 6.04756f
C6 minus drain_left 0.17184f
C7 drain_right plus 0.366822f
C8 minus drain_right 6.03775f
C9 source drain_left 12.332f
C10 drain_right a_n2158_n2688# 5.627861f
C11 drain_left a_n2158_n2688# 5.9396f
C12 source a_n2158_n2688# 7.411844f
C13 minus a_n2158_n2688# 8.307476f
C14 plus a_n2158_n2688# 9.864679f
C15 drain_right.t0 a_n2158_n2688# 0.191299f
C16 drain_right.t1 a_n2158_n2688# 0.191299f
C17 drain_right.n0 a_n2158_n2688# 1.67794f
C18 drain_right.t6 a_n2158_n2688# 0.191299f
C19 drain_right.t5 a_n2158_n2688# 0.191299f
C20 drain_right.n1 a_n2158_n2688# 1.67322f
C21 drain_right.t4 a_n2158_n2688# 0.191299f
C22 drain_right.t8 a_n2158_n2688# 0.191299f
C23 drain_right.n2 a_n2158_n2688# 1.67794f
C24 drain_right.n3 a_n2158_n2688# 2.22924f
C25 drain_right.t11 a_n2158_n2688# 0.191299f
C26 drain_right.t7 a_n2158_n2688# 0.191299f
C27 drain_right.n4 a_n2158_n2688# 1.6783f
C28 drain_right.t3 a_n2158_n2688# 0.191299f
C29 drain_right.t9 a_n2158_n2688# 0.191299f
C30 drain_right.n5 a_n2158_n2688# 1.67323f
C31 drain_right.n6 a_n2158_n2688# 0.744489f
C32 drain_right.t2 a_n2158_n2688# 0.191299f
C33 drain_right.t10 a_n2158_n2688# 0.191299f
C34 drain_right.n7 a_n2158_n2688# 1.67323f
C35 drain_right.n8 a_n2158_n2688# 0.607277f
C36 minus.n0 a_n2158_n2688# 0.041887f
C37 minus.n1 a_n2158_n2688# 0.009505f
C38 minus.t1 a_n2158_n2688# 0.756802f
C39 minus.n2 a_n2158_n2688# 0.041887f
C40 minus.n3 a_n2158_n2688# 0.009505f
C41 minus.t2 a_n2158_n2688# 0.756802f
C42 minus.t4 a_n2158_n2688# 0.775833f
C43 minus.t0 a_n2158_n2688# 0.756802f
C44 minus.n4 a_n2158_n2688# 0.322655f
C45 minus.n5 a_n2158_n2688# 0.302688f
C46 minus.n6 a_n2158_n2688# 0.175723f
C47 minus.n7 a_n2158_n2688# 0.041887f
C48 minus.n8 a_n2158_n2688# 0.31797f
C49 minus.n9 a_n2158_n2688# 0.009505f
C50 minus.t8 a_n2158_n2688# 0.756802f
C51 minus.n10 a_n2158_n2688# 0.31797f
C52 minus.n11 a_n2158_n2688# 0.041887f
C53 minus.n12 a_n2158_n2688# 0.041887f
C54 minus.n13 a_n2158_n2688# 0.041887f
C55 minus.n14 a_n2158_n2688# 0.31797f
C56 minus.n15 a_n2158_n2688# 0.009505f
C57 minus.t9 a_n2158_n2688# 0.756802f
C58 minus.n16 a_n2158_n2688# 0.316033f
C59 minus.n17 a_n2158_n2688# 1.41963f
C60 minus.n18 a_n2158_n2688# 0.041887f
C61 minus.n19 a_n2158_n2688# 0.009505f
C62 minus.n20 a_n2158_n2688# 0.041887f
C63 minus.n21 a_n2158_n2688# 0.009505f
C64 minus.t11 a_n2158_n2688# 0.775833f
C65 minus.t10 a_n2158_n2688# 0.756802f
C66 minus.n22 a_n2158_n2688# 0.322655f
C67 minus.n23 a_n2158_n2688# 0.302688f
C68 minus.n24 a_n2158_n2688# 0.175723f
C69 minus.n25 a_n2158_n2688# 0.041887f
C70 minus.t5 a_n2158_n2688# 0.756802f
C71 minus.n26 a_n2158_n2688# 0.31797f
C72 minus.n27 a_n2158_n2688# 0.009505f
C73 minus.t6 a_n2158_n2688# 0.756802f
C74 minus.n28 a_n2158_n2688# 0.31797f
C75 minus.n29 a_n2158_n2688# 0.041887f
C76 minus.n30 a_n2158_n2688# 0.041887f
C77 minus.n31 a_n2158_n2688# 0.041887f
C78 minus.t7 a_n2158_n2688# 0.756802f
C79 minus.n32 a_n2158_n2688# 0.31797f
C80 minus.n33 a_n2158_n2688# 0.009505f
C81 minus.t3 a_n2158_n2688# 0.756802f
C82 minus.n34 a_n2158_n2688# 0.316033f
C83 minus.n35 a_n2158_n2688# 0.288007f
C84 minus.n36 a_n2158_n2688# 1.72447f
C85 source.t10 a_n2158_n2688# 1.70949f
C86 source.n0 a_n2158_n2688# 1.02488f
C87 source.t11 a_n2158_n2688# 0.160313f
C88 source.t16 a_n2158_n2688# 0.160313f
C89 source.n1 a_n2158_n2688# 1.34203f
C90 source.n2 a_n2158_n2688# 0.339069f
C91 source.t9 a_n2158_n2688# 0.160313f
C92 source.t17 a_n2158_n2688# 0.160313f
C93 source.n3 a_n2158_n2688# 1.34203f
C94 source.n4 a_n2158_n2688# 0.339069f
C95 source.t15 a_n2158_n2688# 1.70949f
C96 source.n5 a_n2158_n2688# 0.378458f
C97 source.t1 a_n2158_n2688# 1.70949f
C98 source.n6 a_n2158_n2688# 0.378458f
C99 source.t21 a_n2158_n2688# 0.160313f
C100 source.t19 a_n2158_n2688# 0.160313f
C101 source.n7 a_n2158_n2688# 1.34203f
C102 source.n8 a_n2158_n2688# 0.339069f
C103 source.t20 a_n2158_n2688# 0.160313f
C104 source.t2 a_n2158_n2688# 0.160313f
C105 source.n9 a_n2158_n2688# 1.34203f
C106 source.n10 a_n2158_n2688# 0.339069f
C107 source.t0 a_n2158_n2688# 1.70949f
C108 source.n11 a_n2158_n2688# 1.36061f
C109 source.t6 a_n2158_n2688# 1.70949f
C110 source.n12 a_n2158_n2688# 1.36061f
C111 source.t13 a_n2158_n2688# 0.160313f
C112 source.t14 a_n2158_n2688# 0.160313f
C113 source.n13 a_n2158_n2688# 1.34203f
C114 source.n14 a_n2158_n2688# 0.339073f
C115 source.t12 a_n2158_n2688# 0.160313f
C116 source.t7 a_n2158_n2688# 0.160313f
C117 source.n15 a_n2158_n2688# 1.34203f
C118 source.n16 a_n2158_n2688# 0.339073f
C119 source.t8 a_n2158_n2688# 1.70949f
C120 source.n17 a_n2158_n2688# 0.378463f
C121 source.t5 a_n2158_n2688# 1.70949f
C122 source.n18 a_n2158_n2688# 0.378463f
C123 source.t4 a_n2158_n2688# 0.160313f
C124 source.t23 a_n2158_n2688# 0.160313f
C125 source.n19 a_n2158_n2688# 1.34203f
C126 source.n20 a_n2158_n2688# 0.339073f
C127 source.t3 a_n2158_n2688# 0.160313f
C128 source.t18 a_n2158_n2688# 0.160313f
C129 source.n21 a_n2158_n2688# 1.34203f
C130 source.n22 a_n2158_n2688# 0.339073f
C131 source.t22 a_n2158_n2688# 1.70949f
C132 source.n23 a_n2158_n2688# 0.525498f
C133 source.n24 a_n2158_n2688# 1.18688f
C134 drain_left.t8 a_n2158_n2688# 0.192284f
C135 drain_left.t11 a_n2158_n2688# 0.192284f
C136 drain_left.n0 a_n2158_n2688# 1.68658f
C137 drain_left.t7 a_n2158_n2688# 0.192284f
C138 drain_left.t3 a_n2158_n2688# 0.192284f
C139 drain_left.n1 a_n2158_n2688# 1.68184f
C140 drain_left.t9 a_n2158_n2688# 0.192284f
C141 drain_left.t1 a_n2158_n2688# 0.192284f
C142 drain_left.n2 a_n2158_n2688# 1.68658f
C143 drain_left.n3 a_n2158_n2688# 2.29609f
C144 drain_left.t2 a_n2158_n2688# 0.192284f
C145 drain_left.t4 a_n2158_n2688# 0.192284f
C146 drain_left.n4 a_n2158_n2688# 1.68695f
C147 drain_left.t5 a_n2158_n2688# 0.192284f
C148 drain_left.t0 a_n2158_n2688# 0.192284f
C149 drain_left.n5 a_n2158_n2688# 1.68184f
C150 drain_left.n6 a_n2158_n2688# 0.748316f
C151 drain_left.t10 a_n2158_n2688# 0.192284f
C152 drain_left.t6 a_n2158_n2688# 0.192284f
C153 drain_left.n7 a_n2158_n2688# 1.68184f
C154 drain_left.n8 a_n2158_n2688# 0.610412f
C155 plus.n0 a_n2158_n2688# 0.042824f
C156 plus.t7 a_n2158_n2688# 0.773714f
C157 plus.t1 a_n2158_n2688# 0.773714f
C158 plus.n1 a_n2158_n2688# 0.042824f
C159 plus.t6 a_n2158_n2688# 0.773714f
C160 plus.n2 a_n2158_n2688# 0.325076f
C161 plus.n3 a_n2158_n2688# 0.042824f
C162 plus.t0 a_n2158_n2688# 0.773714f
C163 plus.t8 a_n2158_n2688# 0.773714f
C164 plus.n4 a_n2158_n2688# 0.329865f
C165 plus.t2 a_n2158_n2688# 0.793171f
C166 plus.n5 a_n2158_n2688# 0.309452f
C167 plus.n6 a_n2158_n2688# 0.179649f
C168 plus.n7 a_n2158_n2688# 0.009718f
C169 plus.n8 a_n2158_n2688# 0.325076f
C170 plus.n9 a_n2158_n2688# 0.009718f
C171 plus.n10 a_n2158_n2688# 0.042824f
C172 plus.n11 a_n2158_n2688# 0.042824f
C173 plus.n12 a_n2158_n2688# 0.042824f
C174 plus.n13 a_n2158_n2688# 0.009718f
C175 plus.n14 a_n2158_n2688# 0.325076f
C176 plus.n15 a_n2158_n2688# 0.009718f
C177 plus.n16 a_n2158_n2688# 0.323095f
C178 plus.n17 a_n2158_n2688# 0.435594f
C179 plus.n18 a_n2158_n2688# 0.042824f
C180 plus.t11 a_n2158_n2688# 0.773714f
C181 plus.n19 a_n2158_n2688# 0.042824f
C182 plus.t4 a_n2158_n2688# 0.773714f
C183 plus.t3 a_n2158_n2688# 0.773714f
C184 plus.n20 a_n2158_n2688# 0.325076f
C185 plus.n21 a_n2158_n2688# 0.042824f
C186 plus.t5 a_n2158_n2688# 0.773714f
C187 plus.t10 a_n2158_n2688# 0.773714f
C188 plus.n22 a_n2158_n2688# 0.329865f
C189 plus.t9 a_n2158_n2688# 0.793171f
C190 plus.n23 a_n2158_n2688# 0.309452f
C191 plus.n24 a_n2158_n2688# 0.179649f
C192 plus.n25 a_n2158_n2688# 0.009718f
C193 plus.n26 a_n2158_n2688# 0.325076f
C194 plus.n27 a_n2158_n2688# 0.009718f
C195 plus.n28 a_n2158_n2688# 0.042824f
C196 plus.n29 a_n2158_n2688# 0.042824f
C197 plus.n30 a_n2158_n2688# 0.042824f
C198 plus.n31 a_n2158_n2688# 0.009718f
C199 plus.n32 a_n2158_n2688# 0.325076f
C200 plus.n33 a_n2158_n2688# 0.009718f
C201 plus.n34 a_n2158_n2688# 0.323095f
C202 plus.n35 a_n2158_n2688# 1.26954f
.ends

