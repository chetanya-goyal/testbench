* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t11 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 drain_left.t13 plus.t0 source.t6 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X2 drain_right.t12 minus.t1 source.t26 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X3 source.t5 plus.t1 drain_left.t12 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X5 source.t13 plus.t2 drain_left.t11 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X6 source.t25 minus.t2 drain_right.t9 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X7 drain_right.t3 minus.t3 source.t24 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X8 a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X9 a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X10 drain_left.t10 plus.t3 source.t3 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X11 a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X12 source.t23 minus.t4 drain_right.t0 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 source.t22 minus.t5 drain_right.t7 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X14 drain_right.t6 minus.t6 source.t21 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X15 drain_right.t8 minus.t7 source.t20 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 drain_right.t10 minus.t8 source.t19 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X17 drain_left.t9 plus.t4 source.t2 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X18 source.t18 minus.t9 drain_right.t13 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X19 drain_right.t4 minus.t10 source.t17 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X20 drain_left.t8 plus.t5 source.t7 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X21 drain_right.t5 minus.t11 source.t16 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X22 drain_right.t1 minus.t12 source.t15 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X23 source.t1 plus.t6 drain_left.t7 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X24 source.t4 plus.t7 drain_left.t6 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X25 source.t14 minus.t13 drain_right.t2 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X26 drain_left.t5 plus.t8 source.t10 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X27 drain_left.t4 plus.t9 source.t11 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 source.t12 plus.t10 drain_left.t3 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X29 source.t0 plus.t11 drain_left.t2 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X30 drain_left.t1 plus.t12 source.t8 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 drain_left.t0 plus.t13 source.t9 a_n1756_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
R0 minus.n15 minus.t12 435.262
R1 minus.n3 minus.t6 435.262
R2 minus.n32 minus.t3 435.262
R3 minus.n20 minus.t10 435.262
R4 minus.n1 minus.t9 369.534
R5 minus.n14 minus.t13 369.534
R6 minus.n12 minus.t7 369.534
R7 minus.n6 minus.t11 369.534
R8 minus.n4 minus.t5 369.534
R9 minus.n18 minus.t0 369.534
R10 minus.n31 minus.t4 369.534
R11 minus.n29 minus.t8 369.534
R12 minus.n23 minus.t1 369.534
R13 minus.n21 minus.t2 369.534
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 51.1217
R33 minus.n6 minus.n5 51.1217
R34 minus.n23 minus.n22 51.1217
R35 minus.n30 minus.n29 51.1217
R36 minus.n14 minus.n13 43.8187
R37 minus.n5 minus.n4 43.8187
R38 minus.n22 minus.n21 43.8187
R39 minus.n31 minus.n30 43.8187
R40 minus.n15 minus.n14 29.2126
R41 minus.n4 minus.n3 29.2126
R42 minus.n21 minus.n20 29.2126
R43 minus.n32 minus.n31 29.2126
R44 minus.n34 minus.n16 27.51
R45 minus.n12 minus.n11 21.9096
R46 minus.n7 minus.n6 21.9096
R47 minus.n24 minus.n23 21.9096
R48 minus.n29 minus.n28 21.9096
R49 minus.n34 minus.n33 6.57058
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n1 drain_right.t4 270.692
R62 drain_right.n11 drain_right.t1 270.132
R63 drain_right.n8 drain_right.n6 240.694
R64 drain_right.n4 drain_right.n2 240.692
R65 drain_right.n8 drain_right.n7 240.132
R66 drain_right.n10 drain_right.n9 240.132
R67 drain_right.n4 drain_right.n3 240.131
R68 drain_right.n1 drain_right.n0 240.131
R69 drain_right.n2 drain_right.t0 30.0005
R70 drain_right.n2 drain_right.t3 30.0005
R71 drain_right.n3 drain_right.t11 30.0005
R72 drain_right.n3 drain_right.t10 30.0005
R73 drain_right.n0 drain_right.t9 30.0005
R74 drain_right.n0 drain_right.t12 30.0005
R75 drain_right.n6 drain_right.t7 30.0005
R76 drain_right.n6 drain_right.t6 30.0005
R77 drain_right.n7 drain_right.t13 30.0005
R78 drain_right.n7 drain_right.t5 30.0005
R79 drain_right.n9 drain_right.t2 30.0005
R80 drain_right.n9 drain_right.t8 30.0005
R81 drain_right drain_right.n5 21.7025
R82 drain_right drain_right.n11 5.93339
R83 drain_right.n11 drain_right.n10 0.560845
R84 drain_right.n10 drain_right.n8 0.560845
R85 drain_right.n5 drain_right.n1 0.365413
R86 drain_right.n5 drain_right.n4 0.0852402
R87 source.n0 source.t10 253.454
R88 source.n7 source.t21 253.454
R89 source.n27 source.t24 253.453
R90 source.n20 source.t3 253.453
R91 source.n2 source.n1 223.454
R92 source.n4 source.n3 223.454
R93 source.n6 source.n5 223.454
R94 source.n9 source.n8 223.454
R95 source.n11 source.n10 223.454
R96 source.n13 source.n12 223.454
R97 source.n26 source.n25 223.453
R98 source.n24 source.n23 223.453
R99 source.n22 source.n21 223.453
R100 source.n19 source.n18 223.453
R101 source.n17 source.n16 223.453
R102 source.n15 source.n14 223.453
R103 source.n25 source.t19 30.0005
R104 source.n25 source.t23 30.0005
R105 source.n23 source.t26 30.0005
R106 source.n23 source.t27 30.0005
R107 source.n21 source.t17 30.0005
R108 source.n21 source.t25 30.0005
R109 source.n18 source.t8 30.0005
R110 source.n18 source.t13 30.0005
R111 source.n16 source.t2 30.0005
R112 source.n16 source.t1 30.0005
R113 source.n14 source.t6 30.0005
R114 source.n14 source.t5 30.0005
R115 source.n1 source.t9 30.0005
R116 source.n1 source.t12 30.0005
R117 source.n3 source.t11 30.0005
R118 source.n3 source.t4 30.0005
R119 source.n5 source.t7 30.0005
R120 source.n5 source.t0 30.0005
R121 source.n8 source.t16 30.0005
R122 source.n8 source.t22 30.0005
R123 source.n10 source.t20 30.0005
R124 source.n10 source.t18 30.0005
R125 source.n12 source.t15 30.0005
R126 source.n12 source.t14 30.0005
R127 source.n15 source.n13 14.0751
R128 source.n28 source.n0 7.97163
R129 source.n28 source.n27 5.5436
R130 source.n7 source.n6 0.7505
R131 source.n22 source.n20 0.7505
R132 source.n13 source.n11 0.560845
R133 source.n11 source.n9 0.560845
R134 source.n9 source.n7 0.560845
R135 source.n6 source.n4 0.560845
R136 source.n4 source.n2 0.560845
R137 source.n2 source.n0 0.560845
R138 source.n17 source.n15 0.560845
R139 source.n19 source.n17 0.560845
R140 source.n20 source.n19 0.560845
R141 source.n24 source.n22 0.560845
R142 source.n26 source.n24 0.560845
R143 source.n27 source.n26 0.560845
R144 source source.n28 0.188
R145 plus.n3 plus.t5 435.262
R146 plus.n15 plus.t8 435.262
R147 plus.n20 plus.t3 435.262
R148 plus.n32 plus.t0 435.262
R149 plus.n1 plus.t7 369.534
R150 plus.n4 plus.t11 369.534
R151 plus.n6 plus.t9 369.534
R152 plus.n12 plus.t13 369.534
R153 plus.n14 plus.t10 369.534
R154 plus.n18 plus.t6 369.534
R155 plus.n21 plus.t2 369.534
R156 plus.n23 plus.t12 369.534
R157 plus.n29 plus.t4 369.534
R158 plus.n31 plus.t1 369.534
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 51.1217
R178 plus.n13 plus.n12 51.1217
R179 plus.n30 plus.n29 51.1217
R180 plus.n23 plus.n22 51.1217
R181 plus.n5 plus.n4 43.8187
R182 plus.n14 plus.n13 43.8187
R183 plus.n31 plus.n30 43.8187
R184 plus.n22 plus.n21 43.8187
R185 plus.n4 plus.n3 29.2126
R186 plus.n15 plus.n14 29.2126
R187 plus.n32 plus.n31 29.2126
R188 plus.n21 plus.n20 29.2126
R189 plus plus.n33 25.5577
R190 plus.n7 plus.n6 21.9096
R191 plus.n12 plus.n11 21.9096
R192 plus.n29 plus.n28 21.9096
R193 plus.n24 plus.n23 21.9096
R194 plus plus.n16 8.04785
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t8 270.693
R206 drain_left.n1 drain_left.t13 270.692
R207 drain_left.n4 drain_left.n2 240.692
R208 drain_left.n11 drain_left.n10 240.132
R209 drain_left.n9 drain_left.n8 240.132
R210 drain_left.n7 drain_left.n6 240.132
R211 drain_left.n4 drain_left.n3 240.131
R212 drain_left.n1 drain_left.n0 240.131
R213 drain_left.n2 drain_left.t11 30.0005
R214 drain_left.n2 drain_left.t10 30.0005
R215 drain_left.n3 drain_left.t7 30.0005
R216 drain_left.n3 drain_left.t1 30.0005
R217 drain_left.n0 drain_left.t12 30.0005
R218 drain_left.n0 drain_left.t9 30.0005
R219 drain_left.n10 drain_left.t3 30.0005
R220 drain_left.n10 drain_left.t5 30.0005
R221 drain_left.n8 drain_left.t6 30.0005
R222 drain_left.n8 drain_left.t0 30.0005
R223 drain_left.n6 drain_left.t2 30.0005
R224 drain_left.n6 drain_left.t4 30.0005
R225 drain_left drain_left.n5 22.2557
R226 drain_left drain_left.n11 6.21356
R227 drain_left.n9 drain_left.n7 0.560845
R228 drain_left.n11 drain_left.n9 0.560845
R229 drain_left.n5 drain_left.n1 0.365413
R230 drain_left.n5 drain_left.n4 0.0852402
C0 drain_right drain_left 0.89725f
C1 drain_right source 4.83891f
C2 minus drain_left 0.1789f
C3 plus drain_left 0.850994f
C4 minus source 0.884496f
C5 plus source 0.898414f
C6 source drain_left 4.84038f
C7 drain_right minus 0.681224f
C8 drain_right plus 0.332956f
C9 plus minus 3.29676f
C10 drain_right a_n1756_n1088# 3.58998f
C11 drain_left a_n1756_n1088# 3.83347f
C12 source a_n1756_n1088# 2.244264f
C13 minus a_n1756_n1088# 5.566708f
C14 plus a_n1756_n1088# 6.356206f
C15 drain_left.t13 a_n1756_n1088# 0.12341f
C16 drain_left.t12 a_n1756_n1088# 0.026757f
C17 drain_left.t9 a_n1756_n1088# 0.026757f
C18 drain_left.n0 a_n1756_n1088# 0.086816f
C19 drain_left.n1 a_n1756_n1088# 0.441524f
C20 drain_left.t11 a_n1756_n1088# 0.026757f
C21 drain_left.t10 a_n1756_n1088# 0.026757f
C22 drain_left.n2 a_n1756_n1088# 0.087388f
C23 drain_left.t7 a_n1756_n1088# 0.026757f
C24 drain_left.t1 a_n1756_n1088# 0.026757f
C25 drain_left.n3 a_n1756_n1088# 0.086816f
C26 drain_left.n4 a_n1756_n1088# 0.454253f
C27 drain_left.n5 a_n1756_n1088# 0.579885f
C28 drain_left.t8 a_n1756_n1088# 0.12341f
C29 drain_left.t2 a_n1756_n1088# 0.026757f
C30 drain_left.t4 a_n1756_n1088# 0.026757f
C31 drain_left.n6 a_n1756_n1088# 0.086816f
C32 drain_left.n7 a_n1756_n1088# 0.454177f
C33 drain_left.t6 a_n1756_n1088# 0.026757f
C34 drain_left.t0 a_n1756_n1088# 0.026757f
C35 drain_left.n8 a_n1756_n1088# 0.086816f
C36 drain_left.n9 a_n1756_n1088# 0.236979f
C37 drain_left.t3 a_n1756_n1088# 0.026757f
C38 drain_left.t5 a_n1756_n1088# 0.026757f
C39 drain_left.n10 a_n1756_n1088# 0.086816f
C40 drain_left.n11 a_n1756_n1088# 0.423605f
C41 plus.n0 a_n1756_n1088# 0.036919f
C42 plus.t10 a_n1756_n1088# 0.017072f
C43 plus.t13 a_n1756_n1088# 0.017072f
C44 plus.t7 a_n1756_n1088# 0.017072f
C45 plus.n1 a_n1756_n1088# 0.035527f
C46 plus.n2 a_n1756_n1088# 0.0863f
C47 plus.t9 a_n1756_n1088# 0.017072f
C48 plus.t11 a_n1756_n1088# 0.017072f
C49 plus.t5 a_n1756_n1088# 0.020931f
C50 plus.n3 a_n1756_n1088# 0.037417f
C51 plus.n4 a_n1756_n1088# 0.02328f
C52 plus.n5 a_n1756_n1088# 0.015662f
C53 plus.n6 a_n1756_n1088# 0.02328f
C54 plus.n7 a_n1756_n1088# 0.015662f
C55 plus.n8 a_n1756_n1088# 0.036919f
C56 plus.n9 a_n1756_n1088# 0.036919f
C57 plus.n10 a_n1756_n1088# 0.036919f
C58 plus.n11 a_n1756_n1088# 0.015662f
C59 plus.n12 a_n1756_n1088# 0.02328f
C60 plus.n13 a_n1756_n1088# 0.015662f
C61 plus.n14 a_n1756_n1088# 0.02328f
C62 plus.t8 a_n1756_n1088# 0.020931f
C63 plus.n15 a_n1756_n1088# 0.037359f
C64 plus.n16 a_n1756_n1088# 0.259569f
C65 plus.n17 a_n1756_n1088# 0.036919f
C66 plus.t0 a_n1756_n1088# 0.020931f
C67 plus.t1 a_n1756_n1088# 0.017072f
C68 plus.t4 a_n1756_n1088# 0.017072f
C69 plus.t6 a_n1756_n1088# 0.017072f
C70 plus.n18 a_n1756_n1088# 0.035527f
C71 plus.n19 a_n1756_n1088# 0.0863f
C72 plus.t12 a_n1756_n1088# 0.017072f
C73 plus.t2 a_n1756_n1088# 0.017072f
C74 plus.t3 a_n1756_n1088# 0.020931f
C75 plus.n20 a_n1756_n1088# 0.037417f
C76 plus.n21 a_n1756_n1088# 0.02328f
C77 plus.n22 a_n1756_n1088# 0.015662f
C78 plus.n23 a_n1756_n1088# 0.02328f
C79 plus.n24 a_n1756_n1088# 0.015662f
C80 plus.n25 a_n1756_n1088# 0.036919f
C81 plus.n26 a_n1756_n1088# 0.036919f
C82 plus.n27 a_n1756_n1088# 0.036919f
C83 plus.n28 a_n1756_n1088# 0.015662f
C84 plus.n29 a_n1756_n1088# 0.02328f
C85 plus.n30 a_n1756_n1088# 0.015662f
C86 plus.n31 a_n1756_n1088# 0.02328f
C87 plus.n32 a_n1756_n1088# 0.037359f
C88 plus.n33 a_n1756_n1088# 0.804121f
C89 source.t10 a_n1756_n1088# 0.148883f
C90 source.n0 a_n1756_n1088# 0.568899f
C91 source.t9 a_n1756_n1088# 0.035516f
C92 source.t12 a_n1756_n1088# 0.035516f
C93 source.n1 a_n1756_n1088# 0.100174f
C94 source.n2 a_n1756_n1088# 0.289299f
C95 source.t11 a_n1756_n1088# 0.035516f
C96 source.t4 a_n1756_n1088# 0.035516f
C97 source.n3 a_n1756_n1088# 0.100174f
C98 source.n4 a_n1756_n1088# 0.289299f
C99 source.t7 a_n1756_n1088# 0.035516f
C100 source.t0 a_n1756_n1088# 0.035516f
C101 source.n5 a_n1756_n1088# 0.100174f
C102 source.n6 a_n1756_n1088# 0.307427f
C103 source.t21 a_n1756_n1088# 0.148883f
C104 source.n7 a_n1756_n1088# 0.322647f
C105 source.t16 a_n1756_n1088# 0.035516f
C106 source.t22 a_n1756_n1088# 0.035516f
C107 source.n8 a_n1756_n1088# 0.100174f
C108 source.n9 a_n1756_n1088# 0.289299f
C109 source.t20 a_n1756_n1088# 0.035516f
C110 source.t18 a_n1756_n1088# 0.035516f
C111 source.n10 a_n1756_n1088# 0.100174f
C112 source.n11 a_n1756_n1088# 0.289299f
C113 source.t15 a_n1756_n1088# 0.035516f
C114 source.t14 a_n1756_n1088# 0.035516f
C115 source.n12 a_n1756_n1088# 0.100174f
C116 source.n13 a_n1756_n1088# 0.845273f
C117 source.t6 a_n1756_n1088# 0.035516f
C118 source.t5 a_n1756_n1088# 0.035516f
C119 source.n14 a_n1756_n1088# 0.100173f
C120 source.n15 a_n1756_n1088# 0.845273f
C121 source.t2 a_n1756_n1088# 0.035516f
C122 source.t1 a_n1756_n1088# 0.035516f
C123 source.n16 a_n1756_n1088# 0.100173f
C124 source.n17 a_n1756_n1088# 0.289299f
C125 source.t8 a_n1756_n1088# 0.035516f
C126 source.t13 a_n1756_n1088# 0.035516f
C127 source.n18 a_n1756_n1088# 0.100173f
C128 source.n19 a_n1756_n1088# 0.289299f
C129 source.t3 a_n1756_n1088# 0.148883f
C130 source.n20 a_n1756_n1088# 0.322647f
C131 source.t17 a_n1756_n1088# 0.035516f
C132 source.t25 a_n1756_n1088# 0.035516f
C133 source.n21 a_n1756_n1088# 0.100173f
C134 source.n22 a_n1756_n1088# 0.307427f
C135 source.t26 a_n1756_n1088# 0.035516f
C136 source.t27 a_n1756_n1088# 0.035516f
C137 source.n23 a_n1756_n1088# 0.100173f
C138 source.n24 a_n1756_n1088# 0.289299f
C139 source.t19 a_n1756_n1088# 0.035516f
C140 source.t23 a_n1756_n1088# 0.035516f
C141 source.n25 a_n1756_n1088# 0.100173f
C142 source.n26 a_n1756_n1088# 0.289299f
C143 source.t24 a_n1756_n1088# 0.148883f
C144 source.n27 a_n1756_n1088# 0.464633f
C145 source.n28 a_n1756_n1088# 0.601436f
C146 drain_right.t4 a_n1756_n1088# 0.1257f
C147 drain_right.t9 a_n1756_n1088# 0.027254f
C148 drain_right.t12 a_n1756_n1088# 0.027254f
C149 drain_right.n0 a_n1756_n1088# 0.088426f
C150 drain_right.n1 a_n1756_n1088# 0.449715f
C151 drain_right.t0 a_n1756_n1088# 0.027254f
C152 drain_right.t3 a_n1756_n1088# 0.027254f
C153 drain_right.n2 a_n1756_n1088# 0.089009f
C154 drain_right.t11 a_n1756_n1088# 0.027254f
C155 drain_right.t10 a_n1756_n1088# 0.027254f
C156 drain_right.n3 a_n1756_n1088# 0.088426f
C157 drain_right.n4 a_n1756_n1088# 0.462679f
C158 drain_right.n5 a_n1756_n1088# 0.546622f
C159 drain_right.t7 a_n1756_n1088# 0.027254f
C160 drain_right.t6 a_n1756_n1088# 0.027254f
C161 drain_right.n6 a_n1756_n1088# 0.089009f
C162 drain_right.t13 a_n1756_n1088# 0.027254f
C163 drain_right.t5 a_n1756_n1088# 0.027254f
C164 drain_right.n7 a_n1756_n1088# 0.088426f
C165 drain_right.n8 a_n1756_n1088# 0.491335f
C166 drain_right.t2 a_n1756_n1088# 0.027254f
C167 drain_right.t8 a_n1756_n1088# 0.027254f
C168 drain_right.n9 a_n1756_n1088# 0.088426f
C169 drain_right.n10 a_n1756_n1088# 0.241375f
C170 drain_right.t1 a_n1756_n1088# 0.125241f
C171 drain_right.n11 a_n1756_n1088# 0.412554f
C172 minus.n0 a_n1756_n1088# 0.036103f
C173 minus.t12 a_n1756_n1088# 0.020468f
C174 minus.t13 a_n1756_n1088# 0.016694f
C175 minus.t7 a_n1756_n1088# 0.016694f
C176 minus.t9 a_n1756_n1088# 0.016694f
C177 minus.n1 a_n1756_n1088# 0.034741f
C178 minus.n2 a_n1756_n1088# 0.084391f
C179 minus.t11 a_n1756_n1088# 0.016694f
C180 minus.t5 a_n1756_n1088# 0.016694f
C181 minus.t6 a_n1756_n1088# 0.020468f
C182 minus.n3 a_n1756_n1088# 0.036589f
C183 minus.n4 a_n1756_n1088# 0.022765f
C184 minus.n5 a_n1756_n1088# 0.015315f
C185 minus.n6 a_n1756_n1088# 0.022765f
C186 minus.n7 a_n1756_n1088# 0.015315f
C187 minus.n8 a_n1756_n1088# 0.036103f
C188 minus.n9 a_n1756_n1088# 0.036103f
C189 minus.n10 a_n1756_n1088# 0.036103f
C190 minus.n11 a_n1756_n1088# 0.015315f
C191 minus.n12 a_n1756_n1088# 0.022765f
C192 minus.n13 a_n1756_n1088# 0.015315f
C193 minus.n14 a_n1756_n1088# 0.022765f
C194 minus.n15 a_n1756_n1088# 0.036532f
C195 minus.n16 a_n1756_n1088# 0.809855f
C196 minus.n17 a_n1756_n1088# 0.036103f
C197 minus.t4 a_n1756_n1088# 0.016694f
C198 minus.t8 a_n1756_n1088# 0.016694f
C199 minus.t0 a_n1756_n1088# 0.016694f
C200 minus.n18 a_n1756_n1088# 0.034741f
C201 minus.n19 a_n1756_n1088# 0.084391f
C202 minus.t1 a_n1756_n1088# 0.016694f
C203 minus.t2 a_n1756_n1088# 0.016694f
C204 minus.t10 a_n1756_n1088# 0.020468f
C205 minus.n20 a_n1756_n1088# 0.036589f
C206 minus.n21 a_n1756_n1088# 0.022765f
C207 minus.n22 a_n1756_n1088# 0.015315f
C208 minus.n23 a_n1756_n1088# 0.022765f
C209 minus.n24 a_n1756_n1088# 0.015315f
C210 minus.n25 a_n1756_n1088# 0.036103f
C211 minus.n26 a_n1756_n1088# 0.036103f
C212 minus.n27 a_n1756_n1088# 0.036103f
C213 minus.n28 a_n1756_n1088# 0.015315f
C214 minus.n29 a_n1756_n1088# 0.022765f
C215 minus.n30 a_n1756_n1088# 0.015315f
C216 minus.n31 a_n1756_n1088# 0.022765f
C217 minus.t3 a_n1756_n1088# 0.020468f
C218 minus.n32 a_n1756_n1088# 0.036532f
C219 minus.n33 a_n1756_n1088# 0.242013f
C220 minus.n34 a_n1756_n1088# 0.997646f
.ends

