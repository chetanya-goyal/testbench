* NGSPICE file created from diffpair463.ext - technology: sky130A

.subckt diffpair463 minus drain_right drain_left source plus
X0 a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X1 source.t15 minus.t0 drain_right.t5 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X2 source.t7 plus.t0 drain_left.t7 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X3 source.t14 minus.t1 drain_right.t6 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X4 drain_right.t1 minus.t2 source.t13 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X5 source.t6 plus.t1 drain_left.t6 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X6 a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X7 source.t3 plus.t2 drain_left.t5 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X8 drain_right.t2 minus.t3 source.t12 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X9 drain_left.t4 plus.t3 source.t5 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X10 drain_right.t0 minus.t4 source.t11 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X11 drain_left.t3 plus.t4 source.t4 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X12 drain_left.t2 plus.t5 source.t1 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X13 a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X14 drain_left.t1 plus.t6 source.t2 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X15 source.t10 minus.t5 drain_right.t7 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X16 source.t0 plus.t7 drain_left.t0 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X17 a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X18 drain_right.t4 minus.t6 source.t9 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X19 source.t8 minus.t7 drain_right.t3 a_n1746_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
R0 minus.n3 minus.t4 491.44
R1 minus.n13 minus.t0 491.44
R2 minus.n2 minus.t1 469.262
R3 minus.n6 minus.t3 469.262
R4 minus.n8 minus.t7 469.262
R5 minus.n12 minus.t2 469.262
R6 minus.n16 minus.t5 469.262
R7 minus.n18 minus.t6 469.262
R8 minus.n9 minus.n8 161.3
R9 minus.n7 minus.n0 161.3
R10 minus.n6 minus.n5 161.3
R11 minus.n4 minus.n1 161.3
R12 minus.n19 minus.n18 161.3
R13 minus.n17 minus.n10 161.3
R14 minus.n16 minus.n15 161.3
R15 minus.n14 minus.n11 161.3
R16 minus.n4 minus.n3 44.862
R17 minus.n14 minus.n13 44.862
R18 minus.n20 minus.n9 35.8679
R19 minus.n8 minus.n7 28.4823
R20 minus.n18 minus.n17 28.4823
R21 minus.n6 minus.n1 24.1005
R22 minus.n2 minus.n1 24.1005
R23 minus.n12 minus.n11 24.1005
R24 minus.n16 minus.n11 24.1005
R25 minus.n7 minus.n6 19.7187
R26 minus.n17 minus.n16 19.7187
R27 minus.n3 minus.n2 19.7081
R28 minus.n13 minus.n12 19.7081
R29 minus.n20 minus.n19 6.63308
R30 minus.n9 minus.n0 0.189894
R31 minus.n5 minus.n0 0.189894
R32 minus.n5 minus.n4 0.189894
R33 minus.n15 minus.n14 0.189894
R34 minus.n15 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 drain_right.n5 drain_right.n3 60.4404
R38 drain_right.n2 drain_right.n1 59.9411
R39 drain_right.n2 drain_right.n0 59.9411
R40 drain_right.n5 drain_right.n4 59.5527
R41 drain_right drain_right.n2 29.9216
R42 drain_right drain_right.n5 6.54115
R43 drain_right.n1 drain_right.t7 1.6505
R44 drain_right.n1 drain_right.t4 1.6505
R45 drain_right.n0 drain_right.t5 1.6505
R46 drain_right.n0 drain_right.t1 1.6505
R47 drain_right.n3 drain_right.t6 1.6505
R48 drain_right.n3 drain_right.t0 1.6505
R49 drain_right.n4 drain_right.t3 1.6505
R50 drain_right.n4 drain_right.t2 1.6505
R51 source.n530 source.n470 289.615
R52 source.n462 source.n402 289.615
R53 source.n396 source.n336 289.615
R54 source.n328 source.n268 289.615
R55 source.n60 source.n0 289.615
R56 source.n128 source.n68 289.615
R57 source.n194 source.n134 289.615
R58 source.n262 source.n202 289.615
R59 source.n490 source.n489 185
R60 source.n495 source.n494 185
R61 source.n497 source.n496 185
R62 source.n486 source.n485 185
R63 source.n503 source.n502 185
R64 source.n505 source.n504 185
R65 source.n482 source.n481 185
R66 source.n512 source.n511 185
R67 source.n513 source.n480 185
R68 source.n515 source.n514 185
R69 source.n478 source.n477 185
R70 source.n521 source.n520 185
R71 source.n523 source.n522 185
R72 source.n474 source.n473 185
R73 source.n529 source.n528 185
R74 source.n531 source.n530 185
R75 source.n422 source.n421 185
R76 source.n427 source.n426 185
R77 source.n429 source.n428 185
R78 source.n418 source.n417 185
R79 source.n435 source.n434 185
R80 source.n437 source.n436 185
R81 source.n414 source.n413 185
R82 source.n444 source.n443 185
R83 source.n445 source.n412 185
R84 source.n447 source.n446 185
R85 source.n410 source.n409 185
R86 source.n453 source.n452 185
R87 source.n455 source.n454 185
R88 source.n406 source.n405 185
R89 source.n461 source.n460 185
R90 source.n463 source.n462 185
R91 source.n356 source.n355 185
R92 source.n361 source.n360 185
R93 source.n363 source.n362 185
R94 source.n352 source.n351 185
R95 source.n369 source.n368 185
R96 source.n371 source.n370 185
R97 source.n348 source.n347 185
R98 source.n378 source.n377 185
R99 source.n379 source.n346 185
R100 source.n381 source.n380 185
R101 source.n344 source.n343 185
R102 source.n387 source.n386 185
R103 source.n389 source.n388 185
R104 source.n340 source.n339 185
R105 source.n395 source.n394 185
R106 source.n397 source.n396 185
R107 source.n288 source.n287 185
R108 source.n293 source.n292 185
R109 source.n295 source.n294 185
R110 source.n284 source.n283 185
R111 source.n301 source.n300 185
R112 source.n303 source.n302 185
R113 source.n280 source.n279 185
R114 source.n310 source.n309 185
R115 source.n311 source.n278 185
R116 source.n313 source.n312 185
R117 source.n276 source.n275 185
R118 source.n319 source.n318 185
R119 source.n321 source.n320 185
R120 source.n272 source.n271 185
R121 source.n327 source.n326 185
R122 source.n329 source.n328 185
R123 source.n61 source.n60 185
R124 source.n59 source.n58 185
R125 source.n4 source.n3 185
R126 source.n53 source.n52 185
R127 source.n51 source.n50 185
R128 source.n8 source.n7 185
R129 source.n45 source.n44 185
R130 source.n43 source.n10 185
R131 source.n42 source.n41 185
R132 source.n13 source.n11 185
R133 source.n36 source.n35 185
R134 source.n34 source.n33 185
R135 source.n17 source.n16 185
R136 source.n28 source.n27 185
R137 source.n26 source.n25 185
R138 source.n21 source.n20 185
R139 source.n129 source.n128 185
R140 source.n127 source.n126 185
R141 source.n72 source.n71 185
R142 source.n121 source.n120 185
R143 source.n119 source.n118 185
R144 source.n76 source.n75 185
R145 source.n113 source.n112 185
R146 source.n111 source.n78 185
R147 source.n110 source.n109 185
R148 source.n81 source.n79 185
R149 source.n104 source.n103 185
R150 source.n102 source.n101 185
R151 source.n85 source.n84 185
R152 source.n96 source.n95 185
R153 source.n94 source.n93 185
R154 source.n89 source.n88 185
R155 source.n195 source.n194 185
R156 source.n193 source.n192 185
R157 source.n138 source.n137 185
R158 source.n187 source.n186 185
R159 source.n185 source.n184 185
R160 source.n142 source.n141 185
R161 source.n179 source.n178 185
R162 source.n177 source.n144 185
R163 source.n176 source.n175 185
R164 source.n147 source.n145 185
R165 source.n170 source.n169 185
R166 source.n168 source.n167 185
R167 source.n151 source.n150 185
R168 source.n162 source.n161 185
R169 source.n160 source.n159 185
R170 source.n155 source.n154 185
R171 source.n263 source.n262 185
R172 source.n261 source.n260 185
R173 source.n206 source.n205 185
R174 source.n255 source.n254 185
R175 source.n253 source.n252 185
R176 source.n210 source.n209 185
R177 source.n247 source.n246 185
R178 source.n245 source.n212 185
R179 source.n244 source.n243 185
R180 source.n215 source.n213 185
R181 source.n238 source.n237 185
R182 source.n236 source.n235 185
R183 source.n219 source.n218 185
R184 source.n230 source.n229 185
R185 source.n228 source.n227 185
R186 source.n223 source.n222 185
R187 source.n491 source.t9 149.524
R188 source.n423 source.t15 149.524
R189 source.n357 source.t2 149.524
R190 source.n289 source.t3 149.524
R191 source.n22 source.t5 149.524
R192 source.n90 source.t6 149.524
R193 source.n156 source.t11 149.524
R194 source.n224 source.t8 149.524
R195 source.n495 source.n489 104.615
R196 source.n496 source.n495 104.615
R197 source.n496 source.n485 104.615
R198 source.n503 source.n485 104.615
R199 source.n504 source.n503 104.615
R200 source.n504 source.n481 104.615
R201 source.n512 source.n481 104.615
R202 source.n513 source.n512 104.615
R203 source.n514 source.n513 104.615
R204 source.n514 source.n477 104.615
R205 source.n521 source.n477 104.615
R206 source.n522 source.n521 104.615
R207 source.n522 source.n473 104.615
R208 source.n529 source.n473 104.615
R209 source.n530 source.n529 104.615
R210 source.n427 source.n421 104.615
R211 source.n428 source.n427 104.615
R212 source.n428 source.n417 104.615
R213 source.n435 source.n417 104.615
R214 source.n436 source.n435 104.615
R215 source.n436 source.n413 104.615
R216 source.n444 source.n413 104.615
R217 source.n445 source.n444 104.615
R218 source.n446 source.n445 104.615
R219 source.n446 source.n409 104.615
R220 source.n453 source.n409 104.615
R221 source.n454 source.n453 104.615
R222 source.n454 source.n405 104.615
R223 source.n461 source.n405 104.615
R224 source.n462 source.n461 104.615
R225 source.n361 source.n355 104.615
R226 source.n362 source.n361 104.615
R227 source.n362 source.n351 104.615
R228 source.n369 source.n351 104.615
R229 source.n370 source.n369 104.615
R230 source.n370 source.n347 104.615
R231 source.n378 source.n347 104.615
R232 source.n379 source.n378 104.615
R233 source.n380 source.n379 104.615
R234 source.n380 source.n343 104.615
R235 source.n387 source.n343 104.615
R236 source.n388 source.n387 104.615
R237 source.n388 source.n339 104.615
R238 source.n395 source.n339 104.615
R239 source.n396 source.n395 104.615
R240 source.n293 source.n287 104.615
R241 source.n294 source.n293 104.615
R242 source.n294 source.n283 104.615
R243 source.n301 source.n283 104.615
R244 source.n302 source.n301 104.615
R245 source.n302 source.n279 104.615
R246 source.n310 source.n279 104.615
R247 source.n311 source.n310 104.615
R248 source.n312 source.n311 104.615
R249 source.n312 source.n275 104.615
R250 source.n319 source.n275 104.615
R251 source.n320 source.n319 104.615
R252 source.n320 source.n271 104.615
R253 source.n327 source.n271 104.615
R254 source.n328 source.n327 104.615
R255 source.n60 source.n59 104.615
R256 source.n59 source.n3 104.615
R257 source.n52 source.n3 104.615
R258 source.n52 source.n51 104.615
R259 source.n51 source.n7 104.615
R260 source.n44 source.n7 104.615
R261 source.n44 source.n43 104.615
R262 source.n43 source.n42 104.615
R263 source.n42 source.n11 104.615
R264 source.n35 source.n11 104.615
R265 source.n35 source.n34 104.615
R266 source.n34 source.n16 104.615
R267 source.n27 source.n16 104.615
R268 source.n27 source.n26 104.615
R269 source.n26 source.n20 104.615
R270 source.n128 source.n127 104.615
R271 source.n127 source.n71 104.615
R272 source.n120 source.n71 104.615
R273 source.n120 source.n119 104.615
R274 source.n119 source.n75 104.615
R275 source.n112 source.n75 104.615
R276 source.n112 source.n111 104.615
R277 source.n111 source.n110 104.615
R278 source.n110 source.n79 104.615
R279 source.n103 source.n79 104.615
R280 source.n103 source.n102 104.615
R281 source.n102 source.n84 104.615
R282 source.n95 source.n84 104.615
R283 source.n95 source.n94 104.615
R284 source.n94 source.n88 104.615
R285 source.n194 source.n193 104.615
R286 source.n193 source.n137 104.615
R287 source.n186 source.n137 104.615
R288 source.n186 source.n185 104.615
R289 source.n185 source.n141 104.615
R290 source.n178 source.n141 104.615
R291 source.n178 source.n177 104.615
R292 source.n177 source.n176 104.615
R293 source.n176 source.n145 104.615
R294 source.n169 source.n145 104.615
R295 source.n169 source.n168 104.615
R296 source.n168 source.n150 104.615
R297 source.n161 source.n150 104.615
R298 source.n161 source.n160 104.615
R299 source.n160 source.n154 104.615
R300 source.n262 source.n261 104.615
R301 source.n261 source.n205 104.615
R302 source.n254 source.n205 104.615
R303 source.n254 source.n253 104.615
R304 source.n253 source.n209 104.615
R305 source.n246 source.n209 104.615
R306 source.n246 source.n245 104.615
R307 source.n245 source.n244 104.615
R308 source.n244 source.n213 104.615
R309 source.n237 source.n213 104.615
R310 source.n237 source.n236 104.615
R311 source.n236 source.n218 104.615
R312 source.n229 source.n218 104.615
R313 source.n229 source.n228 104.615
R314 source.n228 source.n222 104.615
R315 source.t9 source.n489 52.3082
R316 source.t15 source.n421 52.3082
R317 source.t2 source.n355 52.3082
R318 source.t3 source.n287 52.3082
R319 source.t5 source.n20 52.3082
R320 source.t6 source.n88 52.3082
R321 source.t11 source.n154 52.3082
R322 source.t8 source.n222 52.3082
R323 source.n67 source.n66 42.8739
R324 source.n201 source.n200 42.8739
R325 source.n469 source.n468 42.8737
R326 source.n335 source.n334 42.8737
R327 source.n535 source.n534 29.8581
R328 source.n467 source.n466 29.8581
R329 source.n401 source.n400 29.8581
R330 source.n333 source.n332 29.8581
R331 source.n65 source.n64 29.8581
R332 source.n133 source.n132 29.8581
R333 source.n199 source.n198 29.8581
R334 source.n267 source.n266 29.8581
R335 source.n333 source.n267 22.1757
R336 source.n536 source.n65 16.4688
R337 source.n515 source.n480 13.1884
R338 source.n447 source.n412 13.1884
R339 source.n381 source.n346 13.1884
R340 source.n313 source.n278 13.1884
R341 source.n45 source.n10 13.1884
R342 source.n113 source.n78 13.1884
R343 source.n179 source.n144 13.1884
R344 source.n247 source.n212 13.1884
R345 source.n511 source.n510 12.8005
R346 source.n516 source.n478 12.8005
R347 source.n443 source.n442 12.8005
R348 source.n448 source.n410 12.8005
R349 source.n377 source.n376 12.8005
R350 source.n382 source.n344 12.8005
R351 source.n309 source.n308 12.8005
R352 source.n314 source.n276 12.8005
R353 source.n46 source.n8 12.8005
R354 source.n41 source.n12 12.8005
R355 source.n114 source.n76 12.8005
R356 source.n109 source.n80 12.8005
R357 source.n180 source.n142 12.8005
R358 source.n175 source.n146 12.8005
R359 source.n248 source.n210 12.8005
R360 source.n243 source.n214 12.8005
R361 source.n509 source.n482 12.0247
R362 source.n520 source.n519 12.0247
R363 source.n441 source.n414 12.0247
R364 source.n452 source.n451 12.0247
R365 source.n375 source.n348 12.0247
R366 source.n386 source.n385 12.0247
R367 source.n307 source.n280 12.0247
R368 source.n318 source.n317 12.0247
R369 source.n50 source.n49 12.0247
R370 source.n40 source.n13 12.0247
R371 source.n118 source.n117 12.0247
R372 source.n108 source.n81 12.0247
R373 source.n184 source.n183 12.0247
R374 source.n174 source.n147 12.0247
R375 source.n252 source.n251 12.0247
R376 source.n242 source.n215 12.0247
R377 source.n506 source.n505 11.249
R378 source.n523 source.n476 11.249
R379 source.n438 source.n437 11.249
R380 source.n455 source.n408 11.249
R381 source.n372 source.n371 11.249
R382 source.n389 source.n342 11.249
R383 source.n304 source.n303 11.249
R384 source.n321 source.n274 11.249
R385 source.n53 source.n6 11.249
R386 source.n37 source.n36 11.249
R387 source.n121 source.n74 11.249
R388 source.n105 source.n104 11.249
R389 source.n187 source.n140 11.249
R390 source.n171 source.n170 11.249
R391 source.n255 source.n208 11.249
R392 source.n239 source.n238 11.249
R393 source.n502 source.n484 10.4732
R394 source.n524 source.n474 10.4732
R395 source.n434 source.n416 10.4732
R396 source.n456 source.n406 10.4732
R397 source.n368 source.n350 10.4732
R398 source.n390 source.n340 10.4732
R399 source.n300 source.n282 10.4732
R400 source.n322 source.n272 10.4732
R401 source.n54 source.n4 10.4732
R402 source.n33 source.n15 10.4732
R403 source.n122 source.n72 10.4732
R404 source.n101 source.n83 10.4732
R405 source.n188 source.n138 10.4732
R406 source.n167 source.n149 10.4732
R407 source.n256 source.n206 10.4732
R408 source.n235 source.n217 10.4732
R409 source.n491 source.n490 10.2747
R410 source.n423 source.n422 10.2747
R411 source.n357 source.n356 10.2747
R412 source.n289 source.n288 10.2747
R413 source.n22 source.n21 10.2747
R414 source.n90 source.n89 10.2747
R415 source.n156 source.n155 10.2747
R416 source.n224 source.n223 10.2747
R417 source.n501 source.n486 9.69747
R418 source.n528 source.n527 9.69747
R419 source.n433 source.n418 9.69747
R420 source.n460 source.n459 9.69747
R421 source.n367 source.n352 9.69747
R422 source.n394 source.n393 9.69747
R423 source.n299 source.n284 9.69747
R424 source.n326 source.n325 9.69747
R425 source.n58 source.n57 9.69747
R426 source.n32 source.n17 9.69747
R427 source.n126 source.n125 9.69747
R428 source.n100 source.n85 9.69747
R429 source.n192 source.n191 9.69747
R430 source.n166 source.n151 9.69747
R431 source.n260 source.n259 9.69747
R432 source.n234 source.n219 9.69747
R433 source.n534 source.n533 9.45567
R434 source.n466 source.n465 9.45567
R435 source.n400 source.n399 9.45567
R436 source.n332 source.n331 9.45567
R437 source.n64 source.n63 9.45567
R438 source.n132 source.n131 9.45567
R439 source.n198 source.n197 9.45567
R440 source.n266 source.n265 9.45567
R441 source.n533 source.n532 9.3005
R442 source.n472 source.n471 9.3005
R443 source.n527 source.n526 9.3005
R444 source.n525 source.n524 9.3005
R445 source.n476 source.n475 9.3005
R446 source.n519 source.n518 9.3005
R447 source.n517 source.n516 9.3005
R448 source.n493 source.n492 9.3005
R449 source.n488 source.n487 9.3005
R450 source.n499 source.n498 9.3005
R451 source.n501 source.n500 9.3005
R452 source.n484 source.n483 9.3005
R453 source.n507 source.n506 9.3005
R454 source.n509 source.n508 9.3005
R455 source.n510 source.n479 9.3005
R456 source.n465 source.n464 9.3005
R457 source.n404 source.n403 9.3005
R458 source.n459 source.n458 9.3005
R459 source.n457 source.n456 9.3005
R460 source.n408 source.n407 9.3005
R461 source.n451 source.n450 9.3005
R462 source.n449 source.n448 9.3005
R463 source.n425 source.n424 9.3005
R464 source.n420 source.n419 9.3005
R465 source.n431 source.n430 9.3005
R466 source.n433 source.n432 9.3005
R467 source.n416 source.n415 9.3005
R468 source.n439 source.n438 9.3005
R469 source.n441 source.n440 9.3005
R470 source.n442 source.n411 9.3005
R471 source.n399 source.n398 9.3005
R472 source.n338 source.n337 9.3005
R473 source.n393 source.n392 9.3005
R474 source.n391 source.n390 9.3005
R475 source.n342 source.n341 9.3005
R476 source.n385 source.n384 9.3005
R477 source.n383 source.n382 9.3005
R478 source.n359 source.n358 9.3005
R479 source.n354 source.n353 9.3005
R480 source.n365 source.n364 9.3005
R481 source.n367 source.n366 9.3005
R482 source.n350 source.n349 9.3005
R483 source.n373 source.n372 9.3005
R484 source.n375 source.n374 9.3005
R485 source.n376 source.n345 9.3005
R486 source.n331 source.n330 9.3005
R487 source.n270 source.n269 9.3005
R488 source.n325 source.n324 9.3005
R489 source.n323 source.n322 9.3005
R490 source.n274 source.n273 9.3005
R491 source.n317 source.n316 9.3005
R492 source.n315 source.n314 9.3005
R493 source.n291 source.n290 9.3005
R494 source.n286 source.n285 9.3005
R495 source.n297 source.n296 9.3005
R496 source.n299 source.n298 9.3005
R497 source.n282 source.n281 9.3005
R498 source.n305 source.n304 9.3005
R499 source.n307 source.n306 9.3005
R500 source.n308 source.n277 9.3005
R501 source.n24 source.n23 9.3005
R502 source.n19 source.n18 9.3005
R503 source.n30 source.n29 9.3005
R504 source.n32 source.n31 9.3005
R505 source.n15 source.n14 9.3005
R506 source.n38 source.n37 9.3005
R507 source.n40 source.n39 9.3005
R508 source.n12 source.n9 9.3005
R509 source.n63 source.n62 9.3005
R510 source.n2 source.n1 9.3005
R511 source.n57 source.n56 9.3005
R512 source.n55 source.n54 9.3005
R513 source.n6 source.n5 9.3005
R514 source.n49 source.n48 9.3005
R515 source.n47 source.n46 9.3005
R516 source.n92 source.n91 9.3005
R517 source.n87 source.n86 9.3005
R518 source.n98 source.n97 9.3005
R519 source.n100 source.n99 9.3005
R520 source.n83 source.n82 9.3005
R521 source.n106 source.n105 9.3005
R522 source.n108 source.n107 9.3005
R523 source.n80 source.n77 9.3005
R524 source.n131 source.n130 9.3005
R525 source.n70 source.n69 9.3005
R526 source.n125 source.n124 9.3005
R527 source.n123 source.n122 9.3005
R528 source.n74 source.n73 9.3005
R529 source.n117 source.n116 9.3005
R530 source.n115 source.n114 9.3005
R531 source.n158 source.n157 9.3005
R532 source.n153 source.n152 9.3005
R533 source.n164 source.n163 9.3005
R534 source.n166 source.n165 9.3005
R535 source.n149 source.n148 9.3005
R536 source.n172 source.n171 9.3005
R537 source.n174 source.n173 9.3005
R538 source.n146 source.n143 9.3005
R539 source.n197 source.n196 9.3005
R540 source.n136 source.n135 9.3005
R541 source.n191 source.n190 9.3005
R542 source.n189 source.n188 9.3005
R543 source.n140 source.n139 9.3005
R544 source.n183 source.n182 9.3005
R545 source.n181 source.n180 9.3005
R546 source.n226 source.n225 9.3005
R547 source.n221 source.n220 9.3005
R548 source.n232 source.n231 9.3005
R549 source.n234 source.n233 9.3005
R550 source.n217 source.n216 9.3005
R551 source.n240 source.n239 9.3005
R552 source.n242 source.n241 9.3005
R553 source.n214 source.n211 9.3005
R554 source.n265 source.n264 9.3005
R555 source.n204 source.n203 9.3005
R556 source.n259 source.n258 9.3005
R557 source.n257 source.n256 9.3005
R558 source.n208 source.n207 9.3005
R559 source.n251 source.n250 9.3005
R560 source.n249 source.n248 9.3005
R561 source.n498 source.n497 8.92171
R562 source.n531 source.n472 8.92171
R563 source.n430 source.n429 8.92171
R564 source.n463 source.n404 8.92171
R565 source.n364 source.n363 8.92171
R566 source.n397 source.n338 8.92171
R567 source.n296 source.n295 8.92171
R568 source.n329 source.n270 8.92171
R569 source.n61 source.n2 8.92171
R570 source.n29 source.n28 8.92171
R571 source.n129 source.n70 8.92171
R572 source.n97 source.n96 8.92171
R573 source.n195 source.n136 8.92171
R574 source.n163 source.n162 8.92171
R575 source.n263 source.n204 8.92171
R576 source.n231 source.n230 8.92171
R577 source.n494 source.n488 8.14595
R578 source.n532 source.n470 8.14595
R579 source.n426 source.n420 8.14595
R580 source.n464 source.n402 8.14595
R581 source.n360 source.n354 8.14595
R582 source.n398 source.n336 8.14595
R583 source.n292 source.n286 8.14595
R584 source.n330 source.n268 8.14595
R585 source.n62 source.n0 8.14595
R586 source.n25 source.n19 8.14595
R587 source.n130 source.n68 8.14595
R588 source.n93 source.n87 8.14595
R589 source.n196 source.n134 8.14595
R590 source.n159 source.n153 8.14595
R591 source.n264 source.n202 8.14595
R592 source.n227 source.n221 8.14595
R593 source.n493 source.n490 7.3702
R594 source.n425 source.n422 7.3702
R595 source.n359 source.n356 7.3702
R596 source.n291 source.n288 7.3702
R597 source.n24 source.n21 7.3702
R598 source.n92 source.n89 7.3702
R599 source.n158 source.n155 7.3702
R600 source.n226 source.n223 7.3702
R601 source.n494 source.n493 5.81868
R602 source.n534 source.n470 5.81868
R603 source.n426 source.n425 5.81868
R604 source.n466 source.n402 5.81868
R605 source.n360 source.n359 5.81868
R606 source.n400 source.n336 5.81868
R607 source.n292 source.n291 5.81868
R608 source.n332 source.n268 5.81868
R609 source.n64 source.n0 5.81868
R610 source.n25 source.n24 5.81868
R611 source.n132 source.n68 5.81868
R612 source.n93 source.n92 5.81868
R613 source.n198 source.n134 5.81868
R614 source.n159 source.n158 5.81868
R615 source.n266 source.n202 5.81868
R616 source.n227 source.n226 5.81868
R617 source.n536 source.n535 5.7074
R618 source.n497 source.n488 5.04292
R619 source.n532 source.n531 5.04292
R620 source.n429 source.n420 5.04292
R621 source.n464 source.n463 5.04292
R622 source.n363 source.n354 5.04292
R623 source.n398 source.n397 5.04292
R624 source.n295 source.n286 5.04292
R625 source.n330 source.n329 5.04292
R626 source.n62 source.n61 5.04292
R627 source.n28 source.n19 5.04292
R628 source.n130 source.n129 5.04292
R629 source.n96 source.n87 5.04292
R630 source.n196 source.n195 5.04292
R631 source.n162 source.n153 5.04292
R632 source.n264 source.n263 5.04292
R633 source.n230 source.n221 5.04292
R634 source.n498 source.n486 4.26717
R635 source.n528 source.n472 4.26717
R636 source.n430 source.n418 4.26717
R637 source.n460 source.n404 4.26717
R638 source.n364 source.n352 4.26717
R639 source.n394 source.n338 4.26717
R640 source.n296 source.n284 4.26717
R641 source.n326 source.n270 4.26717
R642 source.n58 source.n2 4.26717
R643 source.n29 source.n17 4.26717
R644 source.n126 source.n70 4.26717
R645 source.n97 source.n85 4.26717
R646 source.n192 source.n136 4.26717
R647 source.n163 source.n151 4.26717
R648 source.n260 source.n204 4.26717
R649 source.n231 source.n219 4.26717
R650 source.n502 source.n501 3.49141
R651 source.n527 source.n474 3.49141
R652 source.n434 source.n433 3.49141
R653 source.n459 source.n406 3.49141
R654 source.n368 source.n367 3.49141
R655 source.n393 source.n340 3.49141
R656 source.n300 source.n299 3.49141
R657 source.n325 source.n272 3.49141
R658 source.n57 source.n4 3.49141
R659 source.n33 source.n32 3.49141
R660 source.n125 source.n72 3.49141
R661 source.n101 source.n100 3.49141
R662 source.n191 source.n138 3.49141
R663 source.n167 source.n166 3.49141
R664 source.n259 source.n206 3.49141
R665 source.n235 source.n234 3.49141
R666 source.n492 source.n491 2.84303
R667 source.n424 source.n423 2.84303
R668 source.n358 source.n357 2.84303
R669 source.n290 source.n289 2.84303
R670 source.n23 source.n22 2.84303
R671 source.n91 source.n90 2.84303
R672 source.n157 source.n156 2.84303
R673 source.n225 source.n224 2.84303
R674 source.n505 source.n484 2.71565
R675 source.n524 source.n523 2.71565
R676 source.n437 source.n416 2.71565
R677 source.n456 source.n455 2.71565
R678 source.n371 source.n350 2.71565
R679 source.n390 source.n389 2.71565
R680 source.n303 source.n282 2.71565
R681 source.n322 source.n321 2.71565
R682 source.n54 source.n53 2.71565
R683 source.n36 source.n15 2.71565
R684 source.n122 source.n121 2.71565
R685 source.n104 source.n83 2.71565
R686 source.n188 source.n187 2.71565
R687 source.n170 source.n149 2.71565
R688 source.n256 source.n255 2.71565
R689 source.n238 source.n217 2.71565
R690 source.n506 source.n482 1.93989
R691 source.n520 source.n476 1.93989
R692 source.n438 source.n414 1.93989
R693 source.n452 source.n408 1.93989
R694 source.n372 source.n348 1.93989
R695 source.n386 source.n342 1.93989
R696 source.n304 source.n280 1.93989
R697 source.n318 source.n274 1.93989
R698 source.n50 source.n6 1.93989
R699 source.n37 source.n13 1.93989
R700 source.n118 source.n74 1.93989
R701 source.n105 source.n81 1.93989
R702 source.n184 source.n140 1.93989
R703 source.n171 source.n147 1.93989
R704 source.n252 source.n208 1.93989
R705 source.n239 source.n215 1.93989
R706 source.n468 source.t13 1.6505
R707 source.n468 source.t10 1.6505
R708 source.n334 source.t1 1.6505
R709 source.n334 source.t0 1.6505
R710 source.n66 source.t4 1.6505
R711 source.n66 source.t7 1.6505
R712 source.n200 source.t12 1.6505
R713 source.n200 source.t14 1.6505
R714 source.n511 source.n509 1.16414
R715 source.n519 source.n478 1.16414
R716 source.n443 source.n441 1.16414
R717 source.n451 source.n410 1.16414
R718 source.n377 source.n375 1.16414
R719 source.n385 source.n344 1.16414
R720 source.n309 source.n307 1.16414
R721 source.n317 source.n276 1.16414
R722 source.n49 source.n8 1.16414
R723 source.n41 source.n40 1.16414
R724 source.n117 source.n76 1.16414
R725 source.n109 source.n108 1.16414
R726 source.n183 source.n142 1.16414
R727 source.n175 source.n174 1.16414
R728 source.n251 source.n210 1.16414
R729 source.n243 source.n242 1.16414
R730 source.n267 source.n201 0.888431
R731 source.n201 source.n199 0.888431
R732 source.n133 source.n67 0.888431
R733 source.n67 source.n65 0.888431
R734 source.n335 source.n333 0.888431
R735 source.n401 source.n335 0.888431
R736 source.n469 source.n467 0.888431
R737 source.n535 source.n469 0.888431
R738 source.n199 source.n133 0.470328
R739 source.n467 source.n401 0.470328
R740 source.n510 source.n480 0.388379
R741 source.n516 source.n515 0.388379
R742 source.n442 source.n412 0.388379
R743 source.n448 source.n447 0.388379
R744 source.n376 source.n346 0.388379
R745 source.n382 source.n381 0.388379
R746 source.n308 source.n278 0.388379
R747 source.n314 source.n313 0.388379
R748 source.n46 source.n45 0.388379
R749 source.n12 source.n10 0.388379
R750 source.n114 source.n113 0.388379
R751 source.n80 source.n78 0.388379
R752 source.n180 source.n179 0.388379
R753 source.n146 source.n144 0.388379
R754 source.n248 source.n247 0.388379
R755 source.n214 source.n212 0.388379
R756 source source.n536 0.188
R757 source.n492 source.n487 0.155672
R758 source.n499 source.n487 0.155672
R759 source.n500 source.n499 0.155672
R760 source.n500 source.n483 0.155672
R761 source.n507 source.n483 0.155672
R762 source.n508 source.n507 0.155672
R763 source.n508 source.n479 0.155672
R764 source.n517 source.n479 0.155672
R765 source.n518 source.n517 0.155672
R766 source.n518 source.n475 0.155672
R767 source.n525 source.n475 0.155672
R768 source.n526 source.n525 0.155672
R769 source.n526 source.n471 0.155672
R770 source.n533 source.n471 0.155672
R771 source.n424 source.n419 0.155672
R772 source.n431 source.n419 0.155672
R773 source.n432 source.n431 0.155672
R774 source.n432 source.n415 0.155672
R775 source.n439 source.n415 0.155672
R776 source.n440 source.n439 0.155672
R777 source.n440 source.n411 0.155672
R778 source.n449 source.n411 0.155672
R779 source.n450 source.n449 0.155672
R780 source.n450 source.n407 0.155672
R781 source.n457 source.n407 0.155672
R782 source.n458 source.n457 0.155672
R783 source.n458 source.n403 0.155672
R784 source.n465 source.n403 0.155672
R785 source.n358 source.n353 0.155672
R786 source.n365 source.n353 0.155672
R787 source.n366 source.n365 0.155672
R788 source.n366 source.n349 0.155672
R789 source.n373 source.n349 0.155672
R790 source.n374 source.n373 0.155672
R791 source.n374 source.n345 0.155672
R792 source.n383 source.n345 0.155672
R793 source.n384 source.n383 0.155672
R794 source.n384 source.n341 0.155672
R795 source.n391 source.n341 0.155672
R796 source.n392 source.n391 0.155672
R797 source.n392 source.n337 0.155672
R798 source.n399 source.n337 0.155672
R799 source.n290 source.n285 0.155672
R800 source.n297 source.n285 0.155672
R801 source.n298 source.n297 0.155672
R802 source.n298 source.n281 0.155672
R803 source.n305 source.n281 0.155672
R804 source.n306 source.n305 0.155672
R805 source.n306 source.n277 0.155672
R806 source.n315 source.n277 0.155672
R807 source.n316 source.n315 0.155672
R808 source.n316 source.n273 0.155672
R809 source.n323 source.n273 0.155672
R810 source.n324 source.n323 0.155672
R811 source.n324 source.n269 0.155672
R812 source.n331 source.n269 0.155672
R813 source.n63 source.n1 0.155672
R814 source.n56 source.n1 0.155672
R815 source.n56 source.n55 0.155672
R816 source.n55 source.n5 0.155672
R817 source.n48 source.n5 0.155672
R818 source.n48 source.n47 0.155672
R819 source.n47 source.n9 0.155672
R820 source.n39 source.n9 0.155672
R821 source.n39 source.n38 0.155672
R822 source.n38 source.n14 0.155672
R823 source.n31 source.n14 0.155672
R824 source.n31 source.n30 0.155672
R825 source.n30 source.n18 0.155672
R826 source.n23 source.n18 0.155672
R827 source.n131 source.n69 0.155672
R828 source.n124 source.n69 0.155672
R829 source.n124 source.n123 0.155672
R830 source.n123 source.n73 0.155672
R831 source.n116 source.n73 0.155672
R832 source.n116 source.n115 0.155672
R833 source.n115 source.n77 0.155672
R834 source.n107 source.n77 0.155672
R835 source.n107 source.n106 0.155672
R836 source.n106 source.n82 0.155672
R837 source.n99 source.n82 0.155672
R838 source.n99 source.n98 0.155672
R839 source.n98 source.n86 0.155672
R840 source.n91 source.n86 0.155672
R841 source.n197 source.n135 0.155672
R842 source.n190 source.n135 0.155672
R843 source.n190 source.n189 0.155672
R844 source.n189 source.n139 0.155672
R845 source.n182 source.n139 0.155672
R846 source.n182 source.n181 0.155672
R847 source.n181 source.n143 0.155672
R848 source.n173 source.n143 0.155672
R849 source.n173 source.n172 0.155672
R850 source.n172 source.n148 0.155672
R851 source.n165 source.n148 0.155672
R852 source.n165 source.n164 0.155672
R853 source.n164 source.n152 0.155672
R854 source.n157 source.n152 0.155672
R855 source.n265 source.n203 0.155672
R856 source.n258 source.n203 0.155672
R857 source.n258 source.n257 0.155672
R858 source.n257 source.n207 0.155672
R859 source.n250 source.n207 0.155672
R860 source.n250 source.n249 0.155672
R861 source.n249 source.n211 0.155672
R862 source.n241 source.n211 0.155672
R863 source.n241 source.n240 0.155672
R864 source.n240 source.n216 0.155672
R865 source.n233 source.n216 0.155672
R866 source.n233 source.n232 0.155672
R867 source.n232 source.n220 0.155672
R868 source.n225 source.n220 0.155672
R869 plus.n3 plus.t1 491.44
R870 plus.n13 plus.t6 491.44
R871 plus.n8 plus.t3 469.262
R872 plus.n6 plus.t0 469.262
R873 plus.n2 plus.t4 469.262
R874 plus.n18 plus.t2 469.262
R875 plus.n16 plus.t5 469.262
R876 plus.n12 plus.t7 469.262
R877 plus.n5 plus.n4 161.3
R878 plus.n6 plus.n1 161.3
R879 plus.n7 plus.n0 161.3
R880 plus.n9 plus.n8 161.3
R881 plus.n15 plus.n14 161.3
R882 plus.n16 plus.n11 161.3
R883 plus.n17 plus.n10 161.3
R884 plus.n19 plus.n18 161.3
R885 plus.n4 plus.n3 44.862
R886 plus.n14 plus.n13 44.862
R887 plus plus.n19 29.749
R888 plus.n8 plus.n7 28.4823
R889 plus.n18 plus.n17 28.4823
R890 plus.n5 plus.n2 24.1005
R891 plus.n6 plus.n5 24.1005
R892 plus.n16 plus.n15 24.1005
R893 plus.n15 plus.n12 24.1005
R894 plus.n7 plus.n6 19.7187
R895 plus.n17 plus.n16 19.7187
R896 plus.n3 plus.n2 19.7081
R897 plus.n13 plus.n12 19.7081
R898 plus plus.n9 12.277
R899 plus.n4 plus.n1 0.189894
R900 plus.n1 plus.n0 0.189894
R901 plus.n9 plus.n0 0.189894
R902 plus.n19 plus.n10 0.189894
R903 plus.n11 plus.n10 0.189894
R904 plus.n14 plus.n11 0.189894
R905 drain_left.n5 drain_left.n3 60.4406
R906 drain_left.n2 drain_left.n1 59.9411
R907 drain_left.n2 drain_left.n0 59.9411
R908 drain_left.n5 drain_left.n4 59.5525
R909 drain_left drain_left.n2 30.4748
R910 drain_left drain_left.n5 6.54115
R911 drain_left.n1 drain_left.t0 1.6505
R912 drain_left.n1 drain_left.t1 1.6505
R913 drain_left.n0 drain_left.t5 1.6505
R914 drain_left.n0 drain_left.t2 1.6505
R915 drain_left.n4 drain_left.t7 1.6505
R916 drain_left.n4 drain_left.t4 1.6505
R917 drain_left.n3 drain_left.t6 1.6505
R918 drain_left.n3 drain_left.t3 1.6505
C0 drain_right plus 0.322995f
C1 drain_left drain_right 0.821811f
C2 plus minus 5.31941f
C3 drain_left minus 0.171089f
C4 drain_right minus 5.53266f
C5 source plus 5.29229f
C6 drain_left source 11.2293f
C7 source drain_right 11.231099f
C8 drain_left plus 5.7015f
C9 source minus 5.27825f
C10 drain_right a_n1746_n3288# 5.664559f
C11 drain_left a_n1746_n3288# 5.9269f
C12 source a_n1746_n3288# 8.956371f
C13 minus a_n1746_n3288# 6.76313f
C14 plus a_n1746_n3288# 8.454321f
C15 drain_left.t5 a_n1746_n3288# 0.257023f
C16 drain_left.t2 a_n1746_n3288# 0.257023f
C17 drain_left.n0 a_n1746_n3288# 2.28939f
C18 drain_left.t0 a_n1746_n3288# 0.257023f
C19 drain_left.t1 a_n1746_n3288# 0.257023f
C20 drain_left.n1 a_n1746_n3288# 2.28939f
C21 drain_left.n2 a_n1746_n3288# 2.02288f
C22 drain_left.t6 a_n1746_n3288# 0.257023f
C23 drain_left.t3 a_n1746_n3288# 0.257023f
C24 drain_left.n3 a_n1746_n3288# 2.2929f
C25 drain_left.t7 a_n1746_n3288# 0.257023f
C26 drain_left.t4 a_n1746_n3288# 0.257023f
C27 drain_left.n4 a_n1746_n3288# 2.28711f
C28 drain_left.n5 a_n1746_n3288# 1.01001f
C29 plus.n0 a_n1746_n3288# 0.044741f
C30 plus.t3 a_n1746_n3288# 1.07167f
C31 plus.t0 a_n1746_n3288# 1.07167f
C32 plus.n1 a_n1746_n3288# 0.044741f
C33 plus.t4 a_n1746_n3288# 1.07167f
C34 plus.n2 a_n1746_n3288# 0.43145f
C35 plus.t1 a_n1746_n3288# 1.09095f
C36 plus.n3 a_n1746_n3288# 0.412241f
C37 plus.n4 a_n1746_n3288# 0.186054f
C38 plus.n5 a_n1746_n3288# 0.010153f
C39 plus.n6 a_n1746_n3288# 0.427401f
C40 plus.n7 a_n1746_n3288# 0.010153f
C41 plus.n8 a_n1746_n3288# 0.424505f
C42 plus.n9 a_n1746_n3288# 0.51477f
C43 plus.n10 a_n1746_n3288# 0.044741f
C44 plus.t2 a_n1746_n3288# 1.07167f
C45 plus.n11 a_n1746_n3288# 0.044741f
C46 plus.t5 a_n1746_n3288# 1.07167f
C47 plus.t7 a_n1746_n3288# 1.07167f
C48 plus.n12 a_n1746_n3288# 0.43145f
C49 plus.t6 a_n1746_n3288# 1.09095f
C50 plus.n13 a_n1746_n3288# 0.412241f
C51 plus.n14 a_n1746_n3288# 0.186054f
C52 plus.n15 a_n1746_n3288# 0.010153f
C53 plus.n16 a_n1746_n3288# 0.427401f
C54 plus.n17 a_n1746_n3288# 0.010153f
C55 plus.n18 a_n1746_n3288# 0.424505f
C56 plus.n19 a_n1746_n3288# 1.32311f
C57 source.n0 a_n1746_n3288# 0.026456f
C58 source.n1 a_n1746_n3288# 0.019973f
C59 source.n2 a_n1746_n3288# 0.010732f
C60 source.n3 a_n1746_n3288# 0.025368f
C61 source.n4 a_n1746_n3288# 0.011364f
C62 source.n5 a_n1746_n3288# 0.019973f
C63 source.n6 a_n1746_n3288# 0.010732f
C64 source.n7 a_n1746_n3288# 0.025368f
C65 source.n8 a_n1746_n3288# 0.011364f
C66 source.n9 a_n1746_n3288# 0.019973f
C67 source.n10 a_n1746_n3288# 0.011048f
C68 source.n11 a_n1746_n3288# 0.025368f
C69 source.n12 a_n1746_n3288# 0.010732f
C70 source.n13 a_n1746_n3288# 0.011364f
C71 source.n14 a_n1746_n3288# 0.019973f
C72 source.n15 a_n1746_n3288# 0.010732f
C73 source.n16 a_n1746_n3288# 0.025368f
C74 source.n17 a_n1746_n3288# 0.011364f
C75 source.n18 a_n1746_n3288# 0.019973f
C76 source.n19 a_n1746_n3288# 0.010732f
C77 source.n20 a_n1746_n3288# 0.019026f
C78 source.n21 a_n1746_n3288# 0.017933f
C79 source.t5 a_n1746_n3288# 0.042845f
C80 source.n22 a_n1746_n3288# 0.144002f
C81 source.n23 a_n1746_n3288# 1.0076f
C82 source.n24 a_n1746_n3288# 0.010732f
C83 source.n25 a_n1746_n3288# 0.011364f
C84 source.n26 a_n1746_n3288# 0.025368f
C85 source.n27 a_n1746_n3288# 0.025368f
C86 source.n28 a_n1746_n3288# 0.011364f
C87 source.n29 a_n1746_n3288# 0.010732f
C88 source.n30 a_n1746_n3288# 0.019973f
C89 source.n31 a_n1746_n3288# 0.019973f
C90 source.n32 a_n1746_n3288# 0.010732f
C91 source.n33 a_n1746_n3288# 0.011364f
C92 source.n34 a_n1746_n3288# 0.025368f
C93 source.n35 a_n1746_n3288# 0.025368f
C94 source.n36 a_n1746_n3288# 0.011364f
C95 source.n37 a_n1746_n3288# 0.010732f
C96 source.n38 a_n1746_n3288# 0.019973f
C97 source.n39 a_n1746_n3288# 0.019973f
C98 source.n40 a_n1746_n3288# 0.010732f
C99 source.n41 a_n1746_n3288# 0.011364f
C100 source.n42 a_n1746_n3288# 0.025368f
C101 source.n43 a_n1746_n3288# 0.025368f
C102 source.n44 a_n1746_n3288# 0.025368f
C103 source.n45 a_n1746_n3288# 0.011048f
C104 source.n46 a_n1746_n3288# 0.010732f
C105 source.n47 a_n1746_n3288# 0.019973f
C106 source.n48 a_n1746_n3288# 0.019973f
C107 source.n49 a_n1746_n3288# 0.010732f
C108 source.n50 a_n1746_n3288# 0.011364f
C109 source.n51 a_n1746_n3288# 0.025368f
C110 source.n52 a_n1746_n3288# 0.025368f
C111 source.n53 a_n1746_n3288# 0.011364f
C112 source.n54 a_n1746_n3288# 0.010732f
C113 source.n55 a_n1746_n3288# 0.019973f
C114 source.n56 a_n1746_n3288# 0.019973f
C115 source.n57 a_n1746_n3288# 0.010732f
C116 source.n58 a_n1746_n3288# 0.011364f
C117 source.n59 a_n1746_n3288# 0.025368f
C118 source.n60 a_n1746_n3288# 0.052057f
C119 source.n61 a_n1746_n3288# 0.011364f
C120 source.n62 a_n1746_n3288# 0.010732f
C121 source.n63 a_n1746_n3288# 0.042892f
C122 source.n64 a_n1746_n3288# 0.02873f
C123 source.n65 a_n1746_n3288# 0.840184f
C124 source.t4 a_n1746_n3288# 0.189398f
C125 source.t7 a_n1746_n3288# 0.189398f
C126 source.n66 a_n1746_n3288# 1.62163f
C127 source.n67 a_n1746_n3288# 0.318486f
C128 source.n68 a_n1746_n3288# 0.026456f
C129 source.n69 a_n1746_n3288# 0.019973f
C130 source.n70 a_n1746_n3288# 0.010732f
C131 source.n71 a_n1746_n3288# 0.025368f
C132 source.n72 a_n1746_n3288# 0.011364f
C133 source.n73 a_n1746_n3288# 0.019973f
C134 source.n74 a_n1746_n3288# 0.010732f
C135 source.n75 a_n1746_n3288# 0.025368f
C136 source.n76 a_n1746_n3288# 0.011364f
C137 source.n77 a_n1746_n3288# 0.019973f
C138 source.n78 a_n1746_n3288# 0.011048f
C139 source.n79 a_n1746_n3288# 0.025368f
C140 source.n80 a_n1746_n3288# 0.010732f
C141 source.n81 a_n1746_n3288# 0.011364f
C142 source.n82 a_n1746_n3288# 0.019973f
C143 source.n83 a_n1746_n3288# 0.010732f
C144 source.n84 a_n1746_n3288# 0.025368f
C145 source.n85 a_n1746_n3288# 0.011364f
C146 source.n86 a_n1746_n3288# 0.019973f
C147 source.n87 a_n1746_n3288# 0.010732f
C148 source.n88 a_n1746_n3288# 0.019026f
C149 source.n89 a_n1746_n3288# 0.017933f
C150 source.t6 a_n1746_n3288# 0.042845f
C151 source.n90 a_n1746_n3288# 0.144002f
C152 source.n91 a_n1746_n3288# 1.0076f
C153 source.n92 a_n1746_n3288# 0.010732f
C154 source.n93 a_n1746_n3288# 0.011364f
C155 source.n94 a_n1746_n3288# 0.025368f
C156 source.n95 a_n1746_n3288# 0.025368f
C157 source.n96 a_n1746_n3288# 0.011364f
C158 source.n97 a_n1746_n3288# 0.010732f
C159 source.n98 a_n1746_n3288# 0.019973f
C160 source.n99 a_n1746_n3288# 0.019973f
C161 source.n100 a_n1746_n3288# 0.010732f
C162 source.n101 a_n1746_n3288# 0.011364f
C163 source.n102 a_n1746_n3288# 0.025368f
C164 source.n103 a_n1746_n3288# 0.025368f
C165 source.n104 a_n1746_n3288# 0.011364f
C166 source.n105 a_n1746_n3288# 0.010732f
C167 source.n106 a_n1746_n3288# 0.019973f
C168 source.n107 a_n1746_n3288# 0.019973f
C169 source.n108 a_n1746_n3288# 0.010732f
C170 source.n109 a_n1746_n3288# 0.011364f
C171 source.n110 a_n1746_n3288# 0.025368f
C172 source.n111 a_n1746_n3288# 0.025368f
C173 source.n112 a_n1746_n3288# 0.025368f
C174 source.n113 a_n1746_n3288# 0.011048f
C175 source.n114 a_n1746_n3288# 0.010732f
C176 source.n115 a_n1746_n3288# 0.019973f
C177 source.n116 a_n1746_n3288# 0.019973f
C178 source.n117 a_n1746_n3288# 0.010732f
C179 source.n118 a_n1746_n3288# 0.011364f
C180 source.n119 a_n1746_n3288# 0.025368f
C181 source.n120 a_n1746_n3288# 0.025368f
C182 source.n121 a_n1746_n3288# 0.011364f
C183 source.n122 a_n1746_n3288# 0.010732f
C184 source.n123 a_n1746_n3288# 0.019973f
C185 source.n124 a_n1746_n3288# 0.019973f
C186 source.n125 a_n1746_n3288# 0.010732f
C187 source.n126 a_n1746_n3288# 0.011364f
C188 source.n127 a_n1746_n3288# 0.025368f
C189 source.n128 a_n1746_n3288# 0.052057f
C190 source.n129 a_n1746_n3288# 0.011364f
C191 source.n130 a_n1746_n3288# 0.010732f
C192 source.n131 a_n1746_n3288# 0.042892f
C193 source.n132 a_n1746_n3288# 0.02873f
C194 source.n133 a_n1746_n3288# 0.102595f
C195 source.n134 a_n1746_n3288# 0.026456f
C196 source.n135 a_n1746_n3288# 0.019973f
C197 source.n136 a_n1746_n3288# 0.010732f
C198 source.n137 a_n1746_n3288# 0.025368f
C199 source.n138 a_n1746_n3288# 0.011364f
C200 source.n139 a_n1746_n3288# 0.019973f
C201 source.n140 a_n1746_n3288# 0.010732f
C202 source.n141 a_n1746_n3288# 0.025368f
C203 source.n142 a_n1746_n3288# 0.011364f
C204 source.n143 a_n1746_n3288# 0.019973f
C205 source.n144 a_n1746_n3288# 0.011048f
C206 source.n145 a_n1746_n3288# 0.025368f
C207 source.n146 a_n1746_n3288# 0.010732f
C208 source.n147 a_n1746_n3288# 0.011364f
C209 source.n148 a_n1746_n3288# 0.019973f
C210 source.n149 a_n1746_n3288# 0.010732f
C211 source.n150 a_n1746_n3288# 0.025368f
C212 source.n151 a_n1746_n3288# 0.011364f
C213 source.n152 a_n1746_n3288# 0.019973f
C214 source.n153 a_n1746_n3288# 0.010732f
C215 source.n154 a_n1746_n3288# 0.019026f
C216 source.n155 a_n1746_n3288# 0.017933f
C217 source.t11 a_n1746_n3288# 0.042845f
C218 source.n156 a_n1746_n3288# 0.144002f
C219 source.n157 a_n1746_n3288# 1.0076f
C220 source.n158 a_n1746_n3288# 0.010732f
C221 source.n159 a_n1746_n3288# 0.011364f
C222 source.n160 a_n1746_n3288# 0.025368f
C223 source.n161 a_n1746_n3288# 0.025368f
C224 source.n162 a_n1746_n3288# 0.011364f
C225 source.n163 a_n1746_n3288# 0.010732f
C226 source.n164 a_n1746_n3288# 0.019973f
C227 source.n165 a_n1746_n3288# 0.019973f
C228 source.n166 a_n1746_n3288# 0.010732f
C229 source.n167 a_n1746_n3288# 0.011364f
C230 source.n168 a_n1746_n3288# 0.025368f
C231 source.n169 a_n1746_n3288# 0.025368f
C232 source.n170 a_n1746_n3288# 0.011364f
C233 source.n171 a_n1746_n3288# 0.010732f
C234 source.n172 a_n1746_n3288# 0.019973f
C235 source.n173 a_n1746_n3288# 0.019973f
C236 source.n174 a_n1746_n3288# 0.010732f
C237 source.n175 a_n1746_n3288# 0.011364f
C238 source.n176 a_n1746_n3288# 0.025368f
C239 source.n177 a_n1746_n3288# 0.025368f
C240 source.n178 a_n1746_n3288# 0.025368f
C241 source.n179 a_n1746_n3288# 0.011048f
C242 source.n180 a_n1746_n3288# 0.010732f
C243 source.n181 a_n1746_n3288# 0.019973f
C244 source.n182 a_n1746_n3288# 0.019973f
C245 source.n183 a_n1746_n3288# 0.010732f
C246 source.n184 a_n1746_n3288# 0.011364f
C247 source.n185 a_n1746_n3288# 0.025368f
C248 source.n186 a_n1746_n3288# 0.025368f
C249 source.n187 a_n1746_n3288# 0.011364f
C250 source.n188 a_n1746_n3288# 0.010732f
C251 source.n189 a_n1746_n3288# 0.019973f
C252 source.n190 a_n1746_n3288# 0.019973f
C253 source.n191 a_n1746_n3288# 0.010732f
C254 source.n192 a_n1746_n3288# 0.011364f
C255 source.n193 a_n1746_n3288# 0.025368f
C256 source.n194 a_n1746_n3288# 0.052057f
C257 source.n195 a_n1746_n3288# 0.011364f
C258 source.n196 a_n1746_n3288# 0.010732f
C259 source.n197 a_n1746_n3288# 0.042892f
C260 source.n198 a_n1746_n3288# 0.02873f
C261 source.n199 a_n1746_n3288# 0.102595f
C262 source.t12 a_n1746_n3288# 0.189398f
C263 source.t14 a_n1746_n3288# 0.189398f
C264 source.n200 a_n1746_n3288# 1.62163f
C265 source.n201 a_n1746_n3288# 0.318486f
C266 source.n202 a_n1746_n3288# 0.026456f
C267 source.n203 a_n1746_n3288# 0.019973f
C268 source.n204 a_n1746_n3288# 0.010732f
C269 source.n205 a_n1746_n3288# 0.025368f
C270 source.n206 a_n1746_n3288# 0.011364f
C271 source.n207 a_n1746_n3288# 0.019973f
C272 source.n208 a_n1746_n3288# 0.010732f
C273 source.n209 a_n1746_n3288# 0.025368f
C274 source.n210 a_n1746_n3288# 0.011364f
C275 source.n211 a_n1746_n3288# 0.019973f
C276 source.n212 a_n1746_n3288# 0.011048f
C277 source.n213 a_n1746_n3288# 0.025368f
C278 source.n214 a_n1746_n3288# 0.010732f
C279 source.n215 a_n1746_n3288# 0.011364f
C280 source.n216 a_n1746_n3288# 0.019973f
C281 source.n217 a_n1746_n3288# 0.010732f
C282 source.n218 a_n1746_n3288# 0.025368f
C283 source.n219 a_n1746_n3288# 0.011364f
C284 source.n220 a_n1746_n3288# 0.019973f
C285 source.n221 a_n1746_n3288# 0.010732f
C286 source.n222 a_n1746_n3288# 0.019026f
C287 source.n223 a_n1746_n3288# 0.017933f
C288 source.t8 a_n1746_n3288# 0.042845f
C289 source.n224 a_n1746_n3288# 0.144002f
C290 source.n225 a_n1746_n3288# 1.0076f
C291 source.n226 a_n1746_n3288# 0.010732f
C292 source.n227 a_n1746_n3288# 0.011364f
C293 source.n228 a_n1746_n3288# 0.025368f
C294 source.n229 a_n1746_n3288# 0.025368f
C295 source.n230 a_n1746_n3288# 0.011364f
C296 source.n231 a_n1746_n3288# 0.010732f
C297 source.n232 a_n1746_n3288# 0.019973f
C298 source.n233 a_n1746_n3288# 0.019973f
C299 source.n234 a_n1746_n3288# 0.010732f
C300 source.n235 a_n1746_n3288# 0.011364f
C301 source.n236 a_n1746_n3288# 0.025368f
C302 source.n237 a_n1746_n3288# 0.025368f
C303 source.n238 a_n1746_n3288# 0.011364f
C304 source.n239 a_n1746_n3288# 0.010732f
C305 source.n240 a_n1746_n3288# 0.019973f
C306 source.n241 a_n1746_n3288# 0.019973f
C307 source.n242 a_n1746_n3288# 0.010732f
C308 source.n243 a_n1746_n3288# 0.011364f
C309 source.n244 a_n1746_n3288# 0.025368f
C310 source.n245 a_n1746_n3288# 0.025368f
C311 source.n246 a_n1746_n3288# 0.025368f
C312 source.n247 a_n1746_n3288# 0.011048f
C313 source.n248 a_n1746_n3288# 0.010732f
C314 source.n249 a_n1746_n3288# 0.019973f
C315 source.n250 a_n1746_n3288# 0.019973f
C316 source.n251 a_n1746_n3288# 0.010732f
C317 source.n252 a_n1746_n3288# 0.011364f
C318 source.n253 a_n1746_n3288# 0.025368f
C319 source.n254 a_n1746_n3288# 0.025368f
C320 source.n255 a_n1746_n3288# 0.011364f
C321 source.n256 a_n1746_n3288# 0.010732f
C322 source.n257 a_n1746_n3288# 0.019973f
C323 source.n258 a_n1746_n3288# 0.019973f
C324 source.n259 a_n1746_n3288# 0.010732f
C325 source.n260 a_n1746_n3288# 0.011364f
C326 source.n261 a_n1746_n3288# 0.025368f
C327 source.n262 a_n1746_n3288# 0.052057f
C328 source.n263 a_n1746_n3288# 0.011364f
C329 source.n264 a_n1746_n3288# 0.010732f
C330 source.n265 a_n1746_n3288# 0.042892f
C331 source.n266 a_n1746_n3288# 0.02873f
C332 source.n267 a_n1746_n3288# 1.16225f
C333 source.n268 a_n1746_n3288# 0.026456f
C334 source.n269 a_n1746_n3288# 0.019973f
C335 source.n270 a_n1746_n3288# 0.010732f
C336 source.n271 a_n1746_n3288# 0.025368f
C337 source.n272 a_n1746_n3288# 0.011364f
C338 source.n273 a_n1746_n3288# 0.019973f
C339 source.n274 a_n1746_n3288# 0.010732f
C340 source.n275 a_n1746_n3288# 0.025368f
C341 source.n276 a_n1746_n3288# 0.011364f
C342 source.n277 a_n1746_n3288# 0.019973f
C343 source.n278 a_n1746_n3288# 0.011048f
C344 source.n279 a_n1746_n3288# 0.025368f
C345 source.n280 a_n1746_n3288# 0.011364f
C346 source.n281 a_n1746_n3288# 0.019973f
C347 source.n282 a_n1746_n3288# 0.010732f
C348 source.n283 a_n1746_n3288# 0.025368f
C349 source.n284 a_n1746_n3288# 0.011364f
C350 source.n285 a_n1746_n3288# 0.019973f
C351 source.n286 a_n1746_n3288# 0.010732f
C352 source.n287 a_n1746_n3288# 0.019026f
C353 source.n288 a_n1746_n3288# 0.017933f
C354 source.t3 a_n1746_n3288# 0.042845f
C355 source.n289 a_n1746_n3288# 0.144002f
C356 source.n290 a_n1746_n3288# 1.0076f
C357 source.n291 a_n1746_n3288# 0.010732f
C358 source.n292 a_n1746_n3288# 0.011364f
C359 source.n293 a_n1746_n3288# 0.025368f
C360 source.n294 a_n1746_n3288# 0.025368f
C361 source.n295 a_n1746_n3288# 0.011364f
C362 source.n296 a_n1746_n3288# 0.010732f
C363 source.n297 a_n1746_n3288# 0.019973f
C364 source.n298 a_n1746_n3288# 0.019973f
C365 source.n299 a_n1746_n3288# 0.010732f
C366 source.n300 a_n1746_n3288# 0.011364f
C367 source.n301 a_n1746_n3288# 0.025368f
C368 source.n302 a_n1746_n3288# 0.025368f
C369 source.n303 a_n1746_n3288# 0.011364f
C370 source.n304 a_n1746_n3288# 0.010732f
C371 source.n305 a_n1746_n3288# 0.019973f
C372 source.n306 a_n1746_n3288# 0.019973f
C373 source.n307 a_n1746_n3288# 0.010732f
C374 source.n308 a_n1746_n3288# 0.010732f
C375 source.n309 a_n1746_n3288# 0.011364f
C376 source.n310 a_n1746_n3288# 0.025368f
C377 source.n311 a_n1746_n3288# 0.025368f
C378 source.n312 a_n1746_n3288# 0.025368f
C379 source.n313 a_n1746_n3288# 0.011048f
C380 source.n314 a_n1746_n3288# 0.010732f
C381 source.n315 a_n1746_n3288# 0.019973f
C382 source.n316 a_n1746_n3288# 0.019973f
C383 source.n317 a_n1746_n3288# 0.010732f
C384 source.n318 a_n1746_n3288# 0.011364f
C385 source.n319 a_n1746_n3288# 0.025368f
C386 source.n320 a_n1746_n3288# 0.025368f
C387 source.n321 a_n1746_n3288# 0.011364f
C388 source.n322 a_n1746_n3288# 0.010732f
C389 source.n323 a_n1746_n3288# 0.019973f
C390 source.n324 a_n1746_n3288# 0.019973f
C391 source.n325 a_n1746_n3288# 0.010732f
C392 source.n326 a_n1746_n3288# 0.011364f
C393 source.n327 a_n1746_n3288# 0.025368f
C394 source.n328 a_n1746_n3288# 0.052057f
C395 source.n329 a_n1746_n3288# 0.011364f
C396 source.n330 a_n1746_n3288# 0.010732f
C397 source.n331 a_n1746_n3288# 0.042892f
C398 source.n332 a_n1746_n3288# 0.02873f
C399 source.n333 a_n1746_n3288# 1.16225f
C400 source.t1 a_n1746_n3288# 0.189398f
C401 source.t0 a_n1746_n3288# 0.189398f
C402 source.n334 a_n1746_n3288# 1.62162f
C403 source.n335 a_n1746_n3288# 0.318496f
C404 source.n336 a_n1746_n3288# 0.026456f
C405 source.n337 a_n1746_n3288# 0.019973f
C406 source.n338 a_n1746_n3288# 0.010732f
C407 source.n339 a_n1746_n3288# 0.025368f
C408 source.n340 a_n1746_n3288# 0.011364f
C409 source.n341 a_n1746_n3288# 0.019973f
C410 source.n342 a_n1746_n3288# 0.010732f
C411 source.n343 a_n1746_n3288# 0.025368f
C412 source.n344 a_n1746_n3288# 0.011364f
C413 source.n345 a_n1746_n3288# 0.019973f
C414 source.n346 a_n1746_n3288# 0.011048f
C415 source.n347 a_n1746_n3288# 0.025368f
C416 source.n348 a_n1746_n3288# 0.011364f
C417 source.n349 a_n1746_n3288# 0.019973f
C418 source.n350 a_n1746_n3288# 0.010732f
C419 source.n351 a_n1746_n3288# 0.025368f
C420 source.n352 a_n1746_n3288# 0.011364f
C421 source.n353 a_n1746_n3288# 0.019973f
C422 source.n354 a_n1746_n3288# 0.010732f
C423 source.n355 a_n1746_n3288# 0.019026f
C424 source.n356 a_n1746_n3288# 0.017933f
C425 source.t2 a_n1746_n3288# 0.042845f
C426 source.n357 a_n1746_n3288# 0.144002f
C427 source.n358 a_n1746_n3288# 1.0076f
C428 source.n359 a_n1746_n3288# 0.010732f
C429 source.n360 a_n1746_n3288# 0.011364f
C430 source.n361 a_n1746_n3288# 0.025368f
C431 source.n362 a_n1746_n3288# 0.025368f
C432 source.n363 a_n1746_n3288# 0.011364f
C433 source.n364 a_n1746_n3288# 0.010732f
C434 source.n365 a_n1746_n3288# 0.019973f
C435 source.n366 a_n1746_n3288# 0.019973f
C436 source.n367 a_n1746_n3288# 0.010732f
C437 source.n368 a_n1746_n3288# 0.011364f
C438 source.n369 a_n1746_n3288# 0.025368f
C439 source.n370 a_n1746_n3288# 0.025368f
C440 source.n371 a_n1746_n3288# 0.011364f
C441 source.n372 a_n1746_n3288# 0.010732f
C442 source.n373 a_n1746_n3288# 0.019973f
C443 source.n374 a_n1746_n3288# 0.019973f
C444 source.n375 a_n1746_n3288# 0.010732f
C445 source.n376 a_n1746_n3288# 0.010732f
C446 source.n377 a_n1746_n3288# 0.011364f
C447 source.n378 a_n1746_n3288# 0.025368f
C448 source.n379 a_n1746_n3288# 0.025368f
C449 source.n380 a_n1746_n3288# 0.025368f
C450 source.n381 a_n1746_n3288# 0.011048f
C451 source.n382 a_n1746_n3288# 0.010732f
C452 source.n383 a_n1746_n3288# 0.019973f
C453 source.n384 a_n1746_n3288# 0.019973f
C454 source.n385 a_n1746_n3288# 0.010732f
C455 source.n386 a_n1746_n3288# 0.011364f
C456 source.n387 a_n1746_n3288# 0.025368f
C457 source.n388 a_n1746_n3288# 0.025368f
C458 source.n389 a_n1746_n3288# 0.011364f
C459 source.n390 a_n1746_n3288# 0.010732f
C460 source.n391 a_n1746_n3288# 0.019973f
C461 source.n392 a_n1746_n3288# 0.019973f
C462 source.n393 a_n1746_n3288# 0.010732f
C463 source.n394 a_n1746_n3288# 0.011364f
C464 source.n395 a_n1746_n3288# 0.025368f
C465 source.n396 a_n1746_n3288# 0.052057f
C466 source.n397 a_n1746_n3288# 0.011364f
C467 source.n398 a_n1746_n3288# 0.010732f
C468 source.n399 a_n1746_n3288# 0.042892f
C469 source.n400 a_n1746_n3288# 0.02873f
C470 source.n401 a_n1746_n3288# 0.102595f
C471 source.n402 a_n1746_n3288# 0.026456f
C472 source.n403 a_n1746_n3288# 0.019973f
C473 source.n404 a_n1746_n3288# 0.010732f
C474 source.n405 a_n1746_n3288# 0.025368f
C475 source.n406 a_n1746_n3288# 0.011364f
C476 source.n407 a_n1746_n3288# 0.019973f
C477 source.n408 a_n1746_n3288# 0.010732f
C478 source.n409 a_n1746_n3288# 0.025368f
C479 source.n410 a_n1746_n3288# 0.011364f
C480 source.n411 a_n1746_n3288# 0.019973f
C481 source.n412 a_n1746_n3288# 0.011048f
C482 source.n413 a_n1746_n3288# 0.025368f
C483 source.n414 a_n1746_n3288# 0.011364f
C484 source.n415 a_n1746_n3288# 0.019973f
C485 source.n416 a_n1746_n3288# 0.010732f
C486 source.n417 a_n1746_n3288# 0.025368f
C487 source.n418 a_n1746_n3288# 0.011364f
C488 source.n419 a_n1746_n3288# 0.019973f
C489 source.n420 a_n1746_n3288# 0.010732f
C490 source.n421 a_n1746_n3288# 0.019026f
C491 source.n422 a_n1746_n3288# 0.017933f
C492 source.t15 a_n1746_n3288# 0.042845f
C493 source.n423 a_n1746_n3288# 0.144002f
C494 source.n424 a_n1746_n3288# 1.0076f
C495 source.n425 a_n1746_n3288# 0.010732f
C496 source.n426 a_n1746_n3288# 0.011364f
C497 source.n427 a_n1746_n3288# 0.025368f
C498 source.n428 a_n1746_n3288# 0.025368f
C499 source.n429 a_n1746_n3288# 0.011364f
C500 source.n430 a_n1746_n3288# 0.010732f
C501 source.n431 a_n1746_n3288# 0.019973f
C502 source.n432 a_n1746_n3288# 0.019973f
C503 source.n433 a_n1746_n3288# 0.010732f
C504 source.n434 a_n1746_n3288# 0.011364f
C505 source.n435 a_n1746_n3288# 0.025368f
C506 source.n436 a_n1746_n3288# 0.025368f
C507 source.n437 a_n1746_n3288# 0.011364f
C508 source.n438 a_n1746_n3288# 0.010732f
C509 source.n439 a_n1746_n3288# 0.019973f
C510 source.n440 a_n1746_n3288# 0.019973f
C511 source.n441 a_n1746_n3288# 0.010732f
C512 source.n442 a_n1746_n3288# 0.010732f
C513 source.n443 a_n1746_n3288# 0.011364f
C514 source.n444 a_n1746_n3288# 0.025368f
C515 source.n445 a_n1746_n3288# 0.025368f
C516 source.n446 a_n1746_n3288# 0.025368f
C517 source.n447 a_n1746_n3288# 0.011048f
C518 source.n448 a_n1746_n3288# 0.010732f
C519 source.n449 a_n1746_n3288# 0.019973f
C520 source.n450 a_n1746_n3288# 0.019973f
C521 source.n451 a_n1746_n3288# 0.010732f
C522 source.n452 a_n1746_n3288# 0.011364f
C523 source.n453 a_n1746_n3288# 0.025368f
C524 source.n454 a_n1746_n3288# 0.025368f
C525 source.n455 a_n1746_n3288# 0.011364f
C526 source.n456 a_n1746_n3288# 0.010732f
C527 source.n457 a_n1746_n3288# 0.019973f
C528 source.n458 a_n1746_n3288# 0.019973f
C529 source.n459 a_n1746_n3288# 0.010732f
C530 source.n460 a_n1746_n3288# 0.011364f
C531 source.n461 a_n1746_n3288# 0.025368f
C532 source.n462 a_n1746_n3288# 0.052057f
C533 source.n463 a_n1746_n3288# 0.011364f
C534 source.n464 a_n1746_n3288# 0.010732f
C535 source.n465 a_n1746_n3288# 0.042892f
C536 source.n466 a_n1746_n3288# 0.02873f
C537 source.n467 a_n1746_n3288# 0.102595f
C538 source.t13 a_n1746_n3288# 0.189398f
C539 source.t10 a_n1746_n3288# 0.189398f
C540 source.n468 a_n1746_n3288# 1.62162f
C541 source.n469 a_n1746_n3288# 0.318496f
C542 source.n470 a_n1746_n3288# 0.026456f
C543 source.n471 a_n1746_n3288# 0.019973f
C544 source.n472 a_n1746_n3288# 0.010732f
C545 source.n473 a_n1746_n3288# 0.025368f
C546 source.n474 a_n1746_n3288# 0.011364f
C547 source.n475 a_n1746_n3288# 0.019973f
C548 source.n476 a_n1746_n3288# 0.010732f
C549 source.n477 a_n1746_n3288# 0.025368f
C550 source.n478 a_n1746_n3288# 0.011364f
C551 source.n479 a_n1746_n3288# 0.019973f
C552 source.n480 a_n1746_n3288# 0.011048f
C553 source.n481 a_n1746_n3288# 0.025368f
C554 source.n482 a_n1746_n3288# 0.011364f
C555 source.n483 a_n1746_n3288# 0.019973f
C556 source.n484 a_n1746_n3288# 0.010732f
C557 source.n485 a_n1746_n3288# 0.025368f
C558 source.n486 a_n1746_n3288# 0.011364f
C559 source.n487 a_n1746_n3288# 0.019973f
C560 source.n488 a_n1746_n3288# 0.010732f
C561 source.n489 a_n1746_n3288# 0.019026f
C562 source.n490 a_n1746_n3288# 0.017933f
C563 source.t9 a_n1746_n3288# 0.042845f
C564 source.n491 a_n1746_n3288# 0.144002f
C565 source.n492 a_n1746_n3288# 1.0076f
C566 source.n493 a_n1746_n3288# 0.010732f
C567 source.n494 a_n1746_n3288# 0.011364f
C568 source.n495 a_n1746_n3288# 0.025368f
C569 source.n496 a_n1746_n3288# 0.025368f
C570 source.n497 a_n1746_n3288# 0.011364f
C571 source.n498 a_n1746_n3288# 0.010732f
C572 source.n499 a_n1746_n3288# 0.019973f
C573 source.n500 a_n1746_n3288# 0.019973f
C574 source.n501 a_n1746_n3288# 0.010732f
C575 source.n502 a_n1746_n3288# 0.011364f
C576 source.n503 a_n1746_n3288# 0.025368f
C577 source.n504 a_n1746_n3288# 0.025368f
C578 source.n505 a_n1746_n3288# 0.011364f
C579 source.n506 a_n1746_n3288# 0.010732f
C580 source.n507 a_n1746_n3288# 0.019973f
C581 source.n508 a_n1746_n3288# 0.019973f
C582 source.n509 a_n1746_n3288# 0.010732f
C583 source.n510 a_n1746_n3288# 0.010732f
C584 source.n511 a_n1746_n3288# 0.011364f
C585 source.n512 a_n1746_n3288# 0.025368f
C586 source.n513 a_n1746_n3288# 0.025368f
C587 source.n514 a_n1746_n3288# 0.025368f
C588 source.n515 a_n1746_n3288# 0.011048f
C589 source.n516 a_n1746_n3288# 0.010732f
C590 source.n517 a_n1746_n3288# 0.019973f
C591 source.n518 a_n1746_n3288# 0.019973f
C592 source.n519 a_n1746_n3288# 0.010732f
C593 source.n520 a_n1746_n3288# 0.011364f
C594 source.n521 a_n1746_n3288# 0.025368f
C595 source.n522 a_n1746_n3288# 0.025368f
C596 source.n523 a_n1746_n3288# 0.011364f
C597 source.n524 a_n1746_n3288# 0.010732f
C598 source.n525 a_n1746_n3288# 0.019973f
C599 source.n526 a_n1746_n3288# 0.019973f
C600 source.n527 a_n1746_n3288# 0.010732f
C601 source.n528 a_n1746_n3288# 0.011364f
C602 source.n529 a_n1746_n3288# 0.025368f
C603 source.n530 a_n1746_n3288# 0.052057f
C604 source.n531 a_n1746_n3288# 0.011364f
C605 source.n532 a_n1746_n3288# 0.010732f
C606 source.n533 a_n1746_n3288# 0.042892f
C607 source.n534 a_n1746_n3288# 0.02873f
C608 source.n535 a_n1746_n3288# 0.232879f
C609 source.n536 a_n1746_n3288# 1.26564f
C610 drain_right.t5 a_n1746_n3288# 0.255585f
C611 drain_right.t1 a_n1746_n3288# 0.255585f
C612 drain_right.n0 a_n1746_n3288# 2.27658f
C613 drain_right.t7 a_n1746_n3288# 0.255585f
C614 drain_right.t4 a_n1746_n3288# 0.255585f
C615 drain_right.n1 a_n1746_n3288# 2.27658f
C616 drain_right.n2 a_n1746_n3288# 1.95553f
C617 drain_right.t6 a_n1746_n3288# 0.255585f
C618 drain_right.t0 a_n1746_n3288# 0.255585f
C619 drain_right.n3 a_n1746_n3288# 2.28006f
C620 drain_right.t3 a_n1746_n3288# 0.255585f
C621 drain_right.t2 a_n1746_n3288# 0.255585f
C622 drain_right.n4 a_n1746_n3288# 2.27432f
C623 drain_right.n5 a_n1746_n3288# 1.00436f
C624 minus.n0 a_n1746_n3288# 0.043948f
C625 minus.n1 a_n1746_n3288# 0.009973f
C626 minus.t3 a_n1746_n3288# 1.05268f
C627 minus.t4 a_n1746_n3288# 1.07161f
C628 minus.t1 a_n1746_n3288# 1.05268f
C629 minus.n2 a_n1746_n3288# 0.423804f
C630 minus.n3 a_n1746_n3288# 0.404935f
C631 minus.n4 a_n1746_n3288# 0.182757f
C632 minus.n5 a_n1746_n3288# 0.043948f
C633 minus.n6 a_n1746_n3288# 0.419827f
C634 minus.n7 a_n1746_n3288# 0.009973f
C635 minus.t7 a_n1746_n3288# 1.05268f
C636 minus.n8 a_n1746_n3288# 0.416982f
C637 minus.n9 a_n1746_n3288# 1.53587f
C638 minus.n10 a_n1746_n3288# 0.043948f
C639 minus.n11 a_n1746_n3288# 0.009973f
C640 minus.t0 a_n1746_n3288# 1.07161f
C641 minus.t2 a_n1746_n3288# 1.05268f
C642 minus.n12 a_n1746_n3288# 0.423804f
C643 minus.n13 a_n1746_n3288# 0.404935f
C644 minus.n14 a_n1746_n3288# 0.182757f
C645 minus.n15 a_n1746_n3288# 0.043948f
C646 minus.t5 a_n1746_n3288# 1.05268f
C647 minus.n16 a_n1746_n3288# 0.419827f
C648 minus.n17 a_n1746_n3288# 0.009973f
C649 minus.t6 a_n1746_n3288# 1.05268f
C650 minus.n18 a_n1746_n3288# 0.416982f
C651 minus.n19 a_n1746_n3288# 0.301014f
C652 minus.n20 a_n1746_n3288# 1.86269f
.ends

