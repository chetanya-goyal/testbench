* NGSPICE file created from diffpair599.ext - technology: sky130A

.subckt diffpair599 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t47 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 source.t45 plus.t1 drain_left.t22 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X2 drain_left.t21 plus.t2 source.t32 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X3 drain_left.t20 plus.t3 source.t31 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X4 source.t12 minus.t0 drain_right.t23 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X5 drain_right.t22 minus.t1 source.t5 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X6 drain_right.t21 minus.t2 source.t14 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X7 source.t6 minus.t3 drain_right.t20 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X8 source.t19 minus.t4 drain_right.t19 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X9 source.t23 minus.t5 drain_right.t18 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X10 source.t42 plus.t4 drain_left.t19 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X11 drain_right.t17 minus.t6 source.t13 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X12 drain_right.t16 minus.t7 source.t0 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X13 source.t43 plus.t5 drain_left.t18 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X14 drain_left.t17 plus.t6 source.t44 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X15 drain_left.t16 plus.t7 source.t46 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X16 a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X17 drain_right.t15 minus.t8 source.t4 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X18 source.t9 minus.t9 drain_right.t14 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X19 drain_left.t15 plus.t8 source.t30 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X20 drain_left.t14 plus.t9 source.t29 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X21 source.t39 plus.t10 drain_left.t13 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X22 drain_left.t12 plus.t11 source.t38 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X23 source.t16 minus.t10 drain_right.t13 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X24 source.t21 minus.t11 drain_right.t12 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X25 source.t1 minus.t12 drain_right.t11 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X26 a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X27 source.t37 plus.t12 drain_left.t11 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X28 drain_right.t10 minus.t13 source.t8 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X29 source.t10 minus.t14 drain_right.t9 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X30 drain_left.t10 plus.t13 source.t25 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X31 drain_left.t9 plus.t14 source.t36 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X32 source.t35 plus.t15 drain_left.t8 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X33 source.t34 plus.t16 drain_left.t7 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X34 source.t33 plus.t17 drain_left.t6 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X35 source.t40 plus.t18 drain_left.t5 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X36 drain_left.t4 plus.t19 source.t28 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X37 drain_right.t8 minus.t15 source.t15 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X38 drain_right.t7 minus.t16 source.t20 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X39 drain_right.t6 minus.t17 source.t11 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X40 drain_right.t5 minus.t18 source.t18 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X41 a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X42 source.t17 minus.t19 drain_right.t4 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X43 source.t22 minus.t20 drain_right.t3 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X44 source.t3 minus.t21 drain_right.t2 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X45 a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X46 drain_right.t1 minus.t22 source.t7 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X47 drain_right.t0 minus.t23 source.t2 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X48 source.t24 plus.t20 drain_left.t3 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X49 source.t27 plus.t21 drain_left.t2 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X50 source.t26 plus.t22 drain_left.t1 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X51 drain_left.t0 plus.t23 source.t41 a_n2354_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
R0 plus.n9 plus.t4 1742.5
R1 plus.n35 plus.t6 1742.5
R2 plus.n46 plus.t0 1742.5
R3 plus.n72 plus.t5 1742.5
R4 plus.n8 plus.t11 1711.1
R5 plus.n13 plus.t16 1711.1
R6 plus.n15 plus.t23 1711.1
R7 plus.n5 plus.t10 1711.1
R8 plus.n20 plus.t14 1711.1
R9 plus.n3 plus.t22 1711.1
R10 plus.n26 plus.t3 1711.1
R11 plus.n28 plus.t12 1711.1
R12 plus.n1 plus.t19 1711.1
R13 plus.n34 plus.t1 1711.1
R14 plus.n45 plus.t15 1711.1
R15 plus.n50 plus.t2 1711.1
R16 plus.n52 plus.t17 1711.1
R17 plus.n42 plus.t8 1711.1
R18 plus.n57 plus.t18 1711.1
R19 plus.n40 plus.t9 1711.1
R20 plus.n63 plus.t20 1711.1
R21 plus.n65 plus.t7 1711.1
R22 plus.n38 plus.t21 1711.1
R23 plus.n71 plus.t13 1711.1
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 34.9195
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus plus.n36 15.1444
R88 plus.n8 plus.n7 12.4157
R89 plus.n34 plus.n33 12.4157
R90 plus.n71 plus.n70 12.4157
R91 plus.n45 plus.n44 12.4157
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 source.n0 source.t44 44.1297
R125 source.n11 source.t42 44.1296
R126 source.n12 source.t8 44.1296
R127 source.n23 source.t6 44.1296
R128 source.n47 source.t13 44.1295
R129 source.n36 source.t23 44.1295
R130 source.n35 source.t47 44.1295
R131 source.n24 source.t43 44.1295
R132 source.n2 source.n1 43.1397
R133 source.n4 source.n3 43.1397
R134 source.n6 source.n5 43.1397
R135 source.n8 source.n7 43.1397
R136 source.n10 source.n9 43.1397
R137 source.n14 source.n13 43.1397
R138 source.n16 source.n15 43.1397
R139 source.n18 source.n17 43.1397
R140 source.n20 source.n19 43.1397
R141 source.n22 source.n21 43.1397
R142 source.n46 source.n45 43.1396
R143 source.n44 source.n43 43.1396
R144 source.n42 source.n41 43.1396
R145 source.n40 source.n39 43.1396
R146 source.n38 source.n37 43.1396
R147 source.n34 source.n33 43.1396
R148 source.n32 source.n31 43.1396
R149 source.n30 source.n29 43.1396
R150 source.n28 source.n27 43.1396
R151 source.n26 source.n25 43.1396
R152 source.n24 source.n23 27.8914
R153 source.n48 source.n0 22.357
R154 source.n48 source.n47 5.53498
R155 source.n45 source.t0 0.9905
R156 source.n45 source.t10 0.9905
R157 source.n43 source.t7 0.9905
R158 source.n43 source.t17 0.9905
R159 source.n41 source.t2 0.9905
R160 source.n41 source.t16 0.9905
R161 source.n39 source.t15 0.9905
R162 source.n39 source.t21 0.9905
R163 source.n37 source.t20 0.9905
R164 source.n37 source.t19 0.9905
R165 source.n33 source.t32 0.9905
R166 source.n33 source.t35 0.9905
R167 source.n31 source.t30 0.9905
R168 source.n31 source.t33 0.9905
R169 source.n29 source.t29 0.9905
R170 source.n29 source.t40 0.9905
R171 source.n27 source.t46 0.9905
R172 source.n27 source.t24 0.9905
R173 source.n25 source.t25 0.9905
R174 source.n25 source.t27 0.9905
R175 source.n1 source.t28 0.9905
R176 source.n1 source.t45 0.9905
R177 source.n3 source.t31 0.9905
R178 source.n3 source.t37 0.9905
R179 source.n5 source.t36 0.9905
R180 source.n5 source.t26 0.9905
R181 source.n7 source.t41 0.9905
R182 source.n7 source.t39 0.9905
R183 source.n9 source.t38 0.9905
R184 source.n9 source.t34 0.9905
R185 source.n13 source.t5 0.9905
R186 source.n13 source.t22 0.9905
R187 source.n15 source.t11 0.9905
R188 source.n15 source.t1 0.9905
R189 source.n17 source.t4 0.9905
R190 source.n17 source.t12 0.9905
R191 source.n19 source.t14 0.9905
R192 source.n19 source.t3 0.9905
R193 source.n21 source.t18 0.9905
R194 source.n21 source.t9 0.9905
R195 source.n23 source.n22 0.543603
R196 source.n22 source.n20 0.543603
R197 source.n20 source.n18 0.543603
R198 source.n18 source.n16 0.543603
R199 source.n16 source.n14 0.543603
R200 source.n14 source.n12 0.543603
R201 source.n11 source.n10 0.543603
R202 source.n10 source.n8 0.543603
R203 source.n8 source.n6 0.543603
R204 source.n6 source.n4 0.543603
R205 source.n4 source.n2 0.543603
R206 source.n2 source.n0 0.543603
R207 source.n26 source.n24 0.543603
R208 source.n28 source.n26 0.543603
R209 source.n30 source.n28 0.543603
R210 source.n32 source.n30 0.543603
R211 source.n34 source.n32 0.543603
R212 source.n35 source.n34 0.543603
R213 source.n38 source.n36 0.543603
R214 source.n40 source.n38 0.543603
R215 source.n42 source.n40 0.543603
R216 source.n44 source.n42 0.543603
R217 source.n46 source.n44 0.543603
R218 source.n47 source.n46 0.543603
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 60.3616
R223 drain_left.n7 drain_left.n5 60.3615
R224 drain_left.n2 drain_left.n0 60.3615
R225 drain_left.n21 drain_left.n20 59.8185
R226 drain_left.n19 drain_left.n18 59.8185
R227 drain_left.n17 drain_left.n16 59.8185
R228 drain_left.n15 drain_left.n14 59.8185
R229 drain_left.n13 drain_left.n12 59.8185
R230 drain_left.n7 drain_left.n6 59.8184
R231 drain_left.n9 drain_left.n8 59.8184
R232 drain_left.n4 drain_left.n3 59.8184
R233 drain_left.n2 drain_left.n1 59.8184
R234 drain_left drain_left.n10 38.5872
R235 drain_left drain_left.n21 6.19632
R236 drain_left.n5 drain_left.t8 0.9905
R237 drain_left.n5 drain_left.t23 0.9905
R238 drain_left.n6 drain_left.t6 0.9905
R239 drain_left.n6 drain_left.t21 0.9905
R240 drain_left.n8 drain_left.t5 0.9905
R241 drain_left.n8 drain_left.t15 0.9905
R242 drain_left.n3 drain_left.t3 0.9905
R243 drain_left.n3 drain_left.t14 0.9905
R244 drain_left.n1 drain_left.t2 0.9905
R245 drain_left.n1 drain_left.t16 0.9905
R246 drain_left.n0 drain_left.t18 0.9905
R247 drain_left.n0 drain_left.t10 0.9905
R248 drain_left.n20 drain_left.t22 0.9905
R249 drain_left.n20 drain_left.t17 0.9905
R250 drain_left.n18 drain_left.t11 0.9905
R251 drain_left.n18 drain_left.t4 0.9905
R252 drain_left.n16 drain_left.t1 0.9905
R253 drain_left.n16 drain_left.t20 0.9905
R254 drain_left.n14 drain_left.t13 0.9905
R255 drain_left.n14 drain_left.t9 0.9905
R256 drain_left.n12 drain_left.t7 0.9905
R257 drain_left.n12 drain_left.t0 0.9905
R258 drain_left.n11 drain_left.t19 0.9905
R259 drain_left.n11 drain_left.t12 0.9905
R260 drain_left.n9 drain_left.n7 0.543603
R261 drain_left.n4 drain_left.n2 0.543603
R262 drain_left.n15 drain_left.n13 0.543603
R263 drain_left.n17 drain_left.n15 0.543603
R264 drain_left.n19 drain_left.n17 0.543603
R265 drain_left.n21 drain_left.n19 0.543603
R266 drain_left.n10 drain_left.n9 0.216706
R267 drain_left.n10 drain_left.n4 0.216706
R268 minus.n35 minus.t3 1742.5
R269 minus.n9 minus.t13 1742.5
R270 minus.n72 minus.t6 1742.5
R271 minus.n46 minus.t5 1742.5
R272 minus.n34 minus.t18 1711.1
R273 minus.n1 minus.t9 1711.1
R274 minus.n28 minus.t2 1711.1
R275 minus.n26 minus.t21 1711.1
R276 minus.n3 minus.t8 1711.1
R277 minus.n20 minus.t0 1711.1
R278 minus.n5 minus.t17 1711.1
R279 minus.n15 minus.t12 1711.1
R280 minus.n13 minus.t1 1711.1
R281 minus.n8 minus.t20 1711.1
R282 minus.n71 minus.t14 1711.1
R283 minus.n38 minus.t7 1711.1
R284 minus.n65 minus.t19 1711.1
R285 minus.n63 minus.t22 1711.1
R286 minus.n40 minus.t10 1711.1
R287 minus.n57 minus.t23 1711.1
R288 minus.n42 minus.t11 1711.1
R289 minus.n52 minus.t15 1711.1
R290 minus.n50 minus.t4 1711.1
R291 minus.n45 minus.t16 1711.1
R292 minus.n10 minus.n9 161.489
R293 minus.n47 minus.n46 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n32 minus.n31 161.3
R297 minus.n30 minus.n29 161.3
R298 minus.n27 minus.n2 161.3
R299 minus.n25 minus.n24 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n19 minus.n18 161.3
R303 minus.n17 minus.n16 161.3
R304 minus.n14 minus.n6 161.3
R305 minus.n12 minus.n11 161.3
R306 minus.n10 minus.n7 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n69 minus.n68 161.3
R310 minus.n67 minus.n66 161.3
R311 minus.n64 minus.n39 161.3
R312 minus.n62 minus.n61 161.3
R313 minus.n60 minus.n59 161.3
R314 minus.n58 minus.n41 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n54 minus.n53 161.3
R317 minus.n51 minus.n43 161.3
R318 minus.n49 minus.n48 161.3
R319 minus.n47 minus.n44 161.3
R320 minus.n33 minus.n32 73.0308
R321 minus.n22 minus.n21 73.0308
R322 minus.n12 minus.n7 73.0308
R323 minus.n49 minus.n44 73.0308
R324 minus.n59 minus.n58 73.0308
R325 minus.n70 minus.n69 73.0308
R326 minus.n29 minus.n1 66.4581
R327 minus.n14 minus.n13 66.4581
R328 minus.n51 minus.n50 66.4581
R329 minus.n66 minus.n38 66.4581
R330 minus.n25 minus.n3 63.5369
R331 minus.n20 minus.n19 63.5369
R332 minus.n57 minus.n56 63.5369
R333 minus.n62 minus.n40 63.5369
R334 minus.n35 minus.n34 60.6157
R335 minus.n9 minus.n8 60.6157
R336 minus.n46 minus.n45 60.6157
R337 minus.n72 minus.n71 60.6157
R338 minus.n28 minus.n27 47.4702
R339 minus.n16 minus.n15 47.4702
R340 minus.n53 minus.n52 47.4702
R341 minus.n65 minus.n64 47.4702
R342 minus.n27 minus.n26 44.549
R343 minus.n16 minus.n5 44.549
R344 minus.n53 minus.n42 44.549
R345 minus.n64 minus.n63 44.549
R346 minus.n74 minus.n36 44.0687
R347 minus.n26 minus.n25 28.4823
R348 minus.n19 minus.n5 28.4823
R349 minus.n56 minus.n42 28.4823
R350 minus.n63 minus.n62 28.4823
R351 minus.n29 minus.n28 25.5611
R352 minus.n15 minus.n14 25.5611
R353 minus.n52 minus.n51 25.5611
R354 minus.n66 minus.n65 25.5611
R355 minus.n34 minus.n33 12.4157
R356 minus.n8 minus.n7 12.4157
R357 minus.n45 minus.n44 12.4157
R358 minus.n71 minus.n70 12.4157
R359 minus.n22 minus.n3 9.49444
R360 minus.n21 minus.n20 9.49444
R361 minus.n58 minus.n57 9.49444
R362 minus.n59 minus.n40 9.49444
R363 minus.n32 minus.n1 6.57323
R364 minus.n13 minus.n12 6.57323
R365 minus.n50 minus.n49 6.57323
R366 minus.n69 minus.n38 6.57323
R367 minus.n74 minus.n73 6.4702
R368 minus.n36 minus.n0 0.189894
R369 minus.n31 minus.n0 0.189894
R370 minus.n31 minus.n30 0.189894
R371 minus.n30 minus.n2 0.189894
R372 minus.n24 minus.n2 0.189894
R373 minus.n24 minus.n23 0.189894
R374 minus.n23 minus.n4 0.189894
R375 minus.n18 minus.n4 0.189894
R376 minus.n18 minus.n17 0.189894
R377 minus.n17 minus.n6 0.189894
R378 minus.n11 minus.n6 0.189894
R379 minus.n11 minus.n10 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n48 minus.n43 0.189894
R382 minus.n54 minus.n43 0.189894
R383 minus.n55 minus.n54 0.189894
R384 minus.n55 minus.n41 0.189894
R385 minus.n60 minus.n41 0.189894
R386 minus.n61 minus.n60 0.189894
R387 minus.n61 minus.n39 0.189894
R388 minus.n67 minus.n39 0.189894
R389 minus.n68 minus.n67 0.189894
R390 minus.n68 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 60.3616
R394 drain_right.n7 drain_right.n5 60.3615
R395 drain_right.n2 drain_right.n0 60.3615
R396 drain_right.n13 drain_right.n12 59.8185
R397 drain_right.n15 drain_right.n14 59.8185
R398 drain_right.n17 drain_right.n16 59.8185
R399 drain_right.n19 drain_right.n18 59.8185
R400 drain_right.n21 drain_right.n20 59.8185
R401 drain_right.n7 drain_right.n6 59.8184
R402 drain_right.n9 drain_right.n8 59.8184
R403 drain_right.n4 drain_right.n3 59.8184
R404 drain_right.n2 drain_right.n1 59.8184
R405 drain_right drain_right.n10 38.0339
R406 drain_right drain_right.n21 6.19632
R407 drain_right.n5 drain_right.t9 0.9905
R408 drain_right.n5 drain_right.t17 0.9905
R409 drain_right.n6 drain_right.t4 0.9905
R410 drain_right.n6 drain_right.t16 0.9905
R411 drain_right.n8 drain_right.t13 0.9905
R412 drain_right.n8 drain_right.t1 0.9905
R413 drain_right.n3 drain_right.t12 0.9905
R414 drain_right.n3 drain_right.t0 0.9905
R415 drain_right.n1 drain_right.t19 0.9905
R416 drain_right.n1 drain_right.t8 0.9905
R417 drain_right.n0 drain_right.t18 0.9905
R418 drain_right.n0 drain_right.t7 0.9905
R419 drain_right.n11 drain_right.t3 0.9905
R420 drain_right.n11 drain_right.t10 0.9905
R421 drain_right.n12 drain_right.t11 0.9905
R422 drain_right.n12 drain_right.t22 0.9905
R423 drain_right.n14 drain_right.t23 0.9905
R424 drain_right.n14 drain_right.t6 0.9905
R425 drain_right.n16 drain_right.t2 0.9905
R426 drain_right.n16 drain_right.t15 0.9905
R427 drain_right.n18 drain_right.t14 0.9905
R428 drain_right.n18 drain_right.t21 0.9905
R429 drain_right.n20 drain_right.t20 0.9905
R430 drain_right.n20 drain_right.t5 0.9905
R431 drain_right.n9 drain_right.n7 0.543603
R432 drain_right.n4 drain_right.n2 0.543603
R433 drain_right.n21 drain_right.n19 0.543603
R434 drain_right.n19 drain_right.n17 0.543603
R435 drain_right.n17 drain_right.n15 0.543603
R436 drain_right.n15 drain_right.n13 0.543603
R437 drain_right.n10 drain_right.n9 0.216706
R438 drain_right.n10 drain_right.n4 0.216706
C0 drain_left minus 0.172624f
C1 plus source 13.117599f
C2 drain_left drain_right 1.26597f
C3 minus plus 7.57549f
C4 plus drain_right 0.387992f
C5 minus source 13.103499f
C6 drain_right source 71.50671f
C7 minus drain_right 13.6137f
C8 drain_left plus 13.845901f
C9 drain_left source 71.506f
C10 drain_right a_n2354_n4888# 9.04497f
C11 drain_left a_n2354_n4888# 9.394731f
C12 source a_n2354_n4888# 13.191905f
C13 minus a_n2354_n4888# 9.817587f
C14 plus a_n2354_n4888# 12.37036f
C15 drain_right.t18 a_n2354_n4888# 0.544769f
C16 drain_right.t7 a_n2354_n4888# 0.544769f
C17 drain_right.n0 a_n2354_n4888# 4.98422f
C18 drain_right.t19 a_n2354_n4888# 0.544769f
C19 drain_right.t8 a_n2354_n4888# 0.544769f
C20 drain_right.n1 a_n2354_n4888# 4.98039f
C21 drain_right.n2 a_n2354_n4888# 0.833076f
C22 drain_right.t12 a_n2354_n4888# 0.544769f
C23 drain_right.t0 a_n2354_n4888# 0.544769f
C24 drain_right.n3 a_n2354_n4888# 4.98039f
C25 drain_right.n4 a_n2354_n4888# 0.378899f
C26 drain_right.t9 a_n2354_n4888# 0.544769f
C27 drain_right.t17 a_n2354_n4888# 0.544769f
C28 drain_right.n5 a_n2354_n4888# 4.98422f
C29 drain_right.t4 a_n2354_n4888# 0.544769f
C30 drain_right.t16 a_n2354_n4888# 0.544769f
C31 drain_right.n6 a_n2354_n4888# 4.98039f
C32 drain_right.n7 a_n2354_n4888# 0.833076f
C33 drain_right.t13 a_n2354_n4888# 0.544769f
C34 drain_right.t1 a_n2354_n4888# 0.544769f
C35 drain_right.n8 a_n2354_n4888# 4.98039f
C36 drain_right.n9 a_n2354_n4888# 0.378899f
C37 drain_right.n10 a_n2354_n4888# 2.47608f
C38 drain_right.t3 a_n2354_n4888# 0.544769f
C39 drain_right.t10 a_n2354_n4888# 0.544769f
C40 drain_right.n11 a_n2354_n4888# 4.98422f
C41 drain_right.t11 a_n2354_n4888# 0.544769f
C42 drain_right.t22 a_n2354_n4888# 0.544769f
C43 drain_right.n12 a_n2354_n4888# 4.98039f
C44 drain_right.n13 a_n2354_n4888# 0.83309f
C45 drain_right.t23 a_n2354_n4888# 0.544769f
C46 drain_right.t6 a_n2354_n4888# 0.544769f
C47 drain_right.n14 a_n2354_n4888# 4.98039f
C48 drain_right.n15 a_n2354_n4888# 0.411517f
C49 drain_right.t2 a_n2354_n4888# 0.544769f
C50 drain_right.t15 a_n2354_n4888# 0.544769f
C51 drain_right.n16 a_n2354_n4888# 4.98039f
C52 drain_right.n17 a_n2354_n4888# 0.411517f
C53 drain_right.t14 a_n2354_n4888# 0.544769f
C54 drain_right.t21 a_n2354_n4888# 0.544769f
C55 drain_right.n18 a_n2354_n4888# 4.98039f
C56 drain_right.n19 a_n2354_n4888# 0.411517f
C57 drain_right.t20 a_n2354_n4888# 0.544769f
C58 drain_right.t5 a_n2354_n4888# 0.544769f
C59 drain_right.n20 a_n2354_n4888# 4.98039f
C60 drain_right.n21 a_n2354_n4888# 0.698424f
C61 minus.n0 a_n2354_n4888# 0.048679f
C62 minus.t3 a_n2354_n4888# 0.828143f
C63 minus.t18 a_n2354_n4888# 0.822628f
C64 minus.t9 a_n2354_n4888# 0.822628f
C65 minus.n1 a_n2354_n4888# 0.305587f
C66 minus.n2 a_n2354_n4888# 0.048679f
C67 minus.t2 a_n2354_n4888# 0.822628f
C68 minus.t21 a_n2354_n4888# 0.822628f
C69 minus.t8 a_n2354_n4888# 0.822628f
C70 minus.n3 a_n2354_n4888# 0.305587f
C71 minus.n4 a_n2354_n4888# 0.048679f
C72 minus.t0 a_n2354_n4888# 0.822628f
C73 minus.t17 a_n2354_n4888# 0.822628f
C74 minus.n5 a_n2354_n4888# 0.305587f
C75 minus.n6 a_n2354_n4888# 0.048679f
C76 minus.t12 a_n2354_n4888# 0.822628f
C77 minus.t1 a_n2354_n4888# 0.822628f
C78 minus.n7 a_n2354_n4888# 0.0187f
C79 minus.t20 a_n2354_n4888# 0.822628f
C80 minus.n8 a_n2354_n4888# 0.305587f
C81 minus.t13 a_n2354_n4888# 0.828143f
C82 minus.n9 a_n2354_n4888# 0.320637f
C83 minus.n10 a_n2354_n4888# 0.104197f
C84 minus.n11 a_n2354_n4888# 0.048679f
C85 minus.n12 a_n2354_n4888# 0.017499f
C86 minus.n13 a_n2354_n4888# 0.305587f
C87 minus.n14 a_n2354_n4888# 0.02005f
C88 minus.n15 a_n2354_n4888# 0.305587f
C89 minus.n16 a_n2354_n4888# 0.02005f
C90 minus.n17 a_n2354_n4888# 0.048679f
C91 minus.n18 a_n2354_n4888# 0.048679f
C92 minus.n19 a_n2354_n4888# 0.02005f
C93 minus.n20 a_n2354_n4888# 0.305587f
C94 minus.n21 a_n2354_n4888# 0.018099f
C95 minus.n22 a_n2354_n4888# 0.018099f
C96 minus.n23 a_n2354_n4888# 0.048679f
C97 minus.n24 a_n2354_n4888# 0.048679f
C98 minus.n25 a_n2354_n4888# 0.02005f
C99 minus.n26 a_n2354_n4888# 0.305587f
C100 minus.n27 a_n2354_n4888# 0.02005f
C101 minus.n28 a_n2354_n4888# 0.305587f
C102 minus.n29 a_n2354_n4888# 0.02005f
C103 minus.n30 a_n2354_n4888# 0.048679f
C104 minus.n31 a_n2354_n4888# 0.048679f
C105 minus.n32 a_n2354_n4888# 0.017499f
C106 minus.n33 a_n2354_n4888# 0.0187f
C107 minus.n34 a_n2354_n4888# 0.305587f
C108 minus.n35 a_n2354_n4888# 0.320572f
C109 minus.n36 a_n2354_n4888# 2.31163f
C110 minus.n37 a_n2354_n4888# 0.048679f
C111 minus.t14 a_n2354_n4888# 0.822628f
C112 minus.t7 a_n2354_n4888# 0.822628f
C113 minus.n38 a_n2354_n4888# 0.305587f
C114 minus.n39 a_n2354_n4888# 0.048679f
C115 minus.t19 a_n2354_n4888# 0.822628f
C116 minus.t22 a_n2354_n4888# 0.822628f
C117 minus.t10 a_n2354_n4888# 0.822628f
C118 minus.n40 a_n2354_n4888# 0.305587f
C119 minus.n41 a_n2354_n4888# 0.048679f
C120 minus.t23 a_n2354_n4888# 0.822628f
C121 minus.t11 a_n2354_n4888# 0.822628f
C122 minus.n42 a_n2354_n4888# 0.305587f
C123 minus.n43 a_n2354_n4888# 0.048679f
C124 minus.t15 a_n2354_n4888# 0.822628f
C125 minus.t4 a_n2354_n4888# 0.822628f
C126 minus.n44 a_n2354_n4888# 0.0187f
C127 minus.t5 a_n2354_n4888# 0.828143f
C128 minus.t16 a_n2354_n4888# 0.822628f
C129 minus.n45 a_n2354_n4888# 0.305587f
C130 minus.n46 a_n2354_n4888# 0.320637f
C131 minus.n47 a_n2354_n4888# 0.104197f
C132 minus.n48 a_n2354_n4888# 0.048679f
C133 minus.n49 a_n2354_n4888# 0.017499f
C134 minus.n50 a_n2354_n4888# 0.305587f
C135 minus.n51 a_n2354_n4888# 0.02005f
C136 minus.n52 a_n2354_n4888# 0.305587f
C137 minus.n53 a_n2354_n4888# 0.02005f
C138 minus.n54 a_n2354_n4888# 0.048679f
C139 minus.n55 a_n2354_n4888# 0.048679f
C140 minus.n56 a_n2354_n4888# 0.02005f
C141 minus.n57 a_n2354_n4888# 0.305587f
C142 minus.n58 a_n2354_n4888# 0.018099f
C143 minus.n59 a_n2354_n4888# 0.018099f
C144 minus.n60 a_n2354_n4888# 0.048679f
C145 minus.n61 a_n2354_n4888# 0.048679f
C146 minus.n62 a_n2354_n4888# 0.02005f
C147 minus.n63 a_n2354_n4888# 0.305587f
C148 minus.n64 a_n2354_n4888# 0.02005f
C149 minus.n65 a_n2354_n4888# 0.305587f
C150 minus.n66 a_n2354_n4888# 0.02005f
C151 minus.n67 a_n2354_n4888# 0.048679f
C152 minus.n68 a_n2354_n4888# 0.048679f
C153 minus.n69 a_n2354_n4888# 0.017499f
C154 minus.n70 a_n2354_n4888# 0.0187f
C155 minus.n71 a_n2354_n4888# 0.305587f
C156 minus.t6 a_n2354_n4888# 0.828143f
C157 minus.n72 a_n2354_n4888# 0.320572f
C158 minus.n73 a_n2354_n4888# 0.314831f
C159 minus.n74 a_n2354_n4888# 2.74515f
C160 drain_left.t18 a_n2354_n4888# 0.545185f
C161 drain_left.t10 a_n2354_n4888# 0.545185f
C162 drain_left.n0 a_n2354_n4888# 4.988029f
C163 drain_left.t2 a_n2354_n4888# 0.545185f
C164 drain_left.t16 a_n2354_n4888# 0.545185f
C165 drain_left.n1 a_n2354_n4888# 4.9842f
C166 drain_left.n2 a_n2354_n4888# 0.833713f
C167 drain_left.t3 a_n2354_n4888# 0.545185f
C168 drain_left.t14 a_n2354_n4888# 0.545185f
C169 drain_left.n3 a_n2354_n4888# 4.9842f
C170 drain_left.n4 a_n2354_n4888# 0.379189f
C171 drain_left.t8 a_n2354_n4888# 0.545185f
C172 drain_left.t23 a_n2354_n4888# 0.545185f
C173 drain_left.n5 a_n2354_n4888# 4.988029f
C174 drain_left.t6 a_n2354_n4888# 0.545185f
C175 drain_left.t21 a_n2354_n4888# 0.545185f
C176 drain_left.n6 a_n2354_n4888# 4.9842f
C177 drain_left.n7 a_n2354_n4888# 0.833713f
C178 drain_left.t5 a_n2354_n4888# 0.545185f
C179 drain_left.t15 a_n2354_n4888# 0.545185f
C180 drain_left.n8 a_n2354_n4888# 4.9842f
C181 drain_left.n9 a_n2354_n4888# 0.379189f
C182 drain_left.n10 a_n2354_n4888# 2.54924f
C183 drain_left.t19 a_n2354_n4888# 0.545185f
C184 drain_left.t12 a_n2354_n4888# 0.545185f
C185 drain_left.n11 a_n2354_n4888# 4.988029f
C186 drain_left.t7 a_n2354_n4888# 0.545185f
C187 drain_left.t0 a_n2354_n4888# 0.545185f
C188 drain_left.n12 a_n2354_n4888# 4.9842f
C189 drain_left.n13 a_n2354_n4888# 0.833727f
C190 drain_left.t13 a_n2354_n4888# 0.545185f
C191 drain_left.t9 a_n2354_n4888# 0.545185f
C192 drain_left.n14 a_n2354_n4888# 4.9842f
C193 drain_left.n15 a_n2354_n4888# 0.411832f
C194 drain_left.t1 a_n2354_n4888# 0.545185f
C195 drain_left.t20 a_n2354_n4888# 0.545185f
C196 drain_left.n16 a_n2354_n4888# 4.9842f
C197 drain_left.n17 a_n2354_n4888# 0.411832f
C198 drain_left.t11 a_n2354_n4888# 0.545185f
C199 drain_left.t4 a_n2354_n4888# 0.545185f
C200 drain_left.n18 a_n2354_n4888# 4.9842f
C201 drain_left.n19 a_n2354_n4888# 0.411832f
C202 drain_left.t22 a_n2354_n4888# 0.545185f
C203 drain_left.t17 a_n2354_n4888# 0.545185f
C204 drain_left.n20 a_n2354_n4888# 4.9842f
C205 drain_left.n21 a_n2354_n4888# 0.698958f
C206 source.t44 a_n2354_n4888# 5.42984f
C207 source.n0 a_n2354_n4888# 2.30949f
C208 source.t28 a_n2354_n4888# 0.475119f
C209 source.t45 a_n2354_n4888# 0.475119f
C210 source.n1 a_n2354_n4888# 4.24776f
C211 source.n2 a_n2354_n4888# 0.413913f
C212 source.t31 a_n2354_n4888# 0.475119f
C213 source.t37 a_n2354_n4888# 0.475119f
C214 source.n3 a_n2354_n4888# 4.24776f
C215 source.n4 a_n2354_n4888# 0.413913f
C216 source.t36 a_n2354_n4888# 0.475119f
C217 source.t26 a_n2354_n4888# 0.475119f
C218 source.n5 a_n2354_n4888# 4.24776f
C219 source.n6 a_n2354_n4888# 0.413913f
C220 source.t41 a_n2354_n4888# 0.475119f
C221 source.t39 a_n2354_n4888# 0.475119f
C222 source.n7 a_n2354_n4888# 4.24776f
C223 source.n8 a_n2354_n4888# 0.413913f
C224 source.t38 a_n2354_n4888# 0.475119f
C225 source.t34 a_n2354_n4888# 0.475119f
C226 source.n9 a_n2354_n4888# 4.24776f
C227 source.n10 a_n2354_n4888# 0.413913f
C228 source.t42 a_n2354_n4888# 5.42985f
C229 source.n11 a_n2354_n4888# 0.520509f
C230 source.t8 a_n2354_n4888# 5.42985f
C231 source.n12 a_n2354_n4888# 0.520509f
C232 source.t5 a_n2354_n4888# 0.475119f
C233 source.t22 a_n2354_n4888# 0.475119f
C234 source.n13 a_n2354_n4888# 4.24776f
C235 source.n14 a_n2354_n4888# 0.413913f
C236 source.t11 a_n2354_n4888# 0.475119f
C237 source.t1 a_n2354_n4888# 0.475119f
C238 source.n15 a_n2354_n4888# 4.24776f
C239 source.n16 a_n2354_n4888# 0.413913f
C240 source.t4 a_n2354_n4888# 0.475119f
C241 source.t12 a_n2354_n4888# 0.475119f
C242 source.n17 a_n2354_n4888# 4.24776f
C243 source.n18 a_n2354_n4888# 0.413913f
C244 source.t14 a_n2354_n4888# 0.475119f
C245 source.t3 a_n2354_n4888# 0.475119f
C246 source.n19 a_n2354_n4888# 4.24776f
C247 source.n20 a_n2354_n4888# 0.413913f
C248 source.t18 a_n2354_n4888# 0.475119f
C249 source.t9 a_n2354_n4888# 0.475119f
C250 source.n21 a_n2354_n4888# 4.24776f
C251 source.n22 a_n2354_n4888# 0.413913f
C252 source.t6 a_n2354_n4888# 5.42985f
C253 source.n23 a_n2354_n4888# 2.84223f
C254 source.t43 a_n2354_n4888# 5.42982f
C255 source.n24 a_n2354_n4888# 2.84226f
C256 source.t25 a_n2354_n4888# 0.475119f
C257 source.t27 a_n2354_n4888# 0.475119f
C258 source.n25 a_n2354_n4888# 4.24777f
C259 source.n26 a_n2354_n4888# 0.413904f
C260 source.t46 a_n2354_n4888# 0.475119f
C261 source.t24 a_n2354_n4888# 0.475119f
C262 source.n27 a_n2354_n4888# 4.24777f
C263 source.n28 a_n2354_n4888# 0.413904f
C264 source.t29 a_n2354_n4888# 0.475119f
C265 source.t40 a_n2354_n4888# 0.475119f
C266 source.n29 a_n2354_n4888# 4.24777f
C267 source.n30 a_n2354_n4888# 0.413904f
C268 source.t30 a_n2354_n4888# 0.475119f
C269 source.t33 a_n2354_n4888# 0.475119f
C270 source.n31 a_n2354_n4888# 4.24777f
C271 source.n32 a_n2354_n4888# 0.413904f
C272 source.t32 a_n2354_n4888# 0.475119f
C273 source.t35 a_n2354_n4888# 0.475119f
C274 source.n33 a_n2354_n4888# 4.24777f
C275 source.n34 a_n2354_n4888# 0.413904f
C276 source.t47 a_n2354_n4888# 5.42982f
C277 source.n35 a_n2354_n4888# 0.520539f
C278 source.t23 a_n2354_n4888# 5.42982f
C279 source.n36 a_n2354_n4888# 0.520539f
C280 source.t20 a_n2354_n4888# 0.475119f
C281 source.t19 a_n2354_n4888# 0.475119f
C282 source.n37 a_n2354_n4888# 4.24777f
C283 source.n38 a_n2354_n4888# 0.413904f
C284 source.t15 a_n2354_n4888# 0.475119f
C285 source.t21 a_n2354_n4888# 0.475119f
C286 source.n39 a_n2354_n4888# 4.24777f
C287 source.n40 a_n2354_n4888# 0.413904f
C288 source.t2 a_n2354_n4888# 0.475119f
C289 source.t16 a_n2354_n4888# 0.475119f
C290 source.n41 a_n2354_n4888# 4.24777f
C291 source.n42 a_n2354_n4888# 0.413904f
C292 source.t7 a_n2354_n4888# 0.475119f
C293 source.t17 a_n2354_n4888# 0.475119f
C294 source.n43 a_n2354_n4888# 4.24777f
C295 source.n44 a_n2354_n4888# 0.413904f
C296 source.t0 a_n2354_n4888# 0.475119f
C297 source.t10 a_n2354_n4888# 0.475119f
C298 source.n45 a_n2354_n4888# 4.24777f
C299 source.n46 a_n2354_n4888# 0.413904f
C300 source.t13 a_n2354_n4888# 5.42982f
C301 source.n47 a_n2354_n4888# 0.690239f
C302 source.n48 a_n2354_n4888# 2.70615f
C303 plus.n0 a_n2354_n4888# 0.049104f
C304 plus.t1 a_n2354_n4888# 0.829806f
C305 plus.t19 a_n2354_n4888# 0.829806f
C306 plus.n1 a_n2354_n4888# 0.308253f
C307 plus.n2 a_n2354_n4888# 0.049104f
C308 plus.t12 a_n2354_n4888# 0.829806f
C309 plus.t3 a_n2354_n4888# 0.829806f
C310 plus.t22 a_n2354_n4888# 0.829806f
C311 plus.n3 a_n2354_n4888# 0.308253f
C312 plus.n4 a_n2354_n4888# 0.049104f
C313 plus.t14 a_n2354_n4888# 0.829806f
C314 plus.t10 a_n2354_n4888# 0.829806f
C315 plus.n5 a_n2354_n4888# 0.308253f
C316 plus.n6 a_n2354_n4888# 0.049104f
C317 plus.t23 a_n2354_n4888# 0.829806f
C318 plus.t16 a_n2354_n4888# 0.829806f
C319 plus.n7 a_n2354_n4888# 0.018863f
C320 plus.t4 a_n2354_n4888# 0.83537f
C321 plus.t11 a_n2354_n4888# 0.829806f
C322 plus.n8 a_n2354_n4888# 0.308253f
C323 plus.n9 a_n2354_n4888# 0.323435f
C324 plus.n10 a_n2354_n4888# 0.105106f
C325 plus.n11 a_n2354_n4888# 0.049104f
C326 plus.n12 a_n2354_n4888# 0.017652f
C327 plus.n13 a_n2354_n4888# 0.308253f
C328 plus.n14 a_n2354_n4888# 0.020225f
C329 plus.n15 a_n2354_n4888# 0.308253f
C330 plus.n16 a_n2354_n4888# 0.020225f
C331 plus.n17 a_n2354_n4888# 0.049104f
C332 plus.n18 a_n2354_n4888# 0.049104f
C333 plus.n19 a_n2354_n4888# 0.020225f
C334 plus.n20 a_n2354_n4888# 0.308253f
C335 plus.n21 a_n2354_n4888# 0.018257f
C336 plus.n22 a_n2354_n4888# 0.018257f
C337 plus.n23 a_n2354_n4888# 0.049104f
C338 plus.n24 a_n2354_n4888# 0.049104f
C339 plus.n25 a_n2354_n4888# 0.020225f
C340 plus.n26 a_n2354_n4888# 0.308253f
C341 plus.n27 a_n2354_n4888# 0.020225f
C342 plus.n28 a_n2354_n4888# 0.308253f
C343 plus.n29 a_n2354_n4888# 0.020225f
C344 plus.n30 a_n2354_n4888# 0.049104f
C345 plus.n31 a_n2354_n4888# 0.049104f
C346 plus.n32 a_n2354_n4888# 0.017652f
C347 plus.n33 a_n2354_n4888# 0.018863f
C348 plus.n34 a_n2354_n4888# 0.308253f
C349 plus.t6 a_n2354_n4888# 0.83537f
C350 plus.n35 a_n2354_n4888# 0.323369f
C351 plus.n36 a_n2354_n4888# 0.742246f
C352 plus.n37 a_n2354_n4888# 0.049104f
C353 plus.t5 a_n2354_n4888# 0.83537f
C354 plus.t13 a_n2354_n4888# 0.829806f
C355 plus.t21 a_n2354_n4888# 0.829806f
C356 plus.n38 a_n2354_n4888# 0.308253f
C357 plus.n39 a_n2354_n4888# 0.049104f
C358 plus.t7 a_n2354_n4888# 0.829806f
C359 plus.t20 a_n2354_n4888# 0.829806f
C360 plus.t9 a_n2354_n4888# 0.829806f
C361 plus.n40 a_n2354_n4888# 0.308253f
C362 plus.n41 a_n2354_n4888# 0.049104f
C363 plus.t18 a_n2354_n4888# 0.829806f
C364 plus.t8 a_n2354_n4888# 0.829806f
C365 plus.n42 a_n2354_n4888# 0.308253f
C366 plus.n43 a_n2354_n4888# 0.049104f
C367 plus.t17 a_n2354_n4888# 0.829806f
C368 plus.t2 a_n2354_n4888# 0.829806f
C369 plus.n44 a_n2354_n4888# 0.018863f
C370 plus.t15 a_n2354_n4888# 0.829806f
C371 plus.n45 a_n2354_n4888# 0.308253f
C372 plus.t0 a_n2354_n4888# 0.83537f
C373 plus.n46 a_n2354_n4888# 0.323435f
C374 plus.n47 a_n2354_n4888# 0.105106f
C375 plus.n48 a_n2354_n4888# 0.049104f
C376 plus.n49 a_n2354_n4888# 0.017652f
C377 plus.n50 a_n2354_n4888# 0.308253f
C378 plus.n51 a_n2354_n4888# 0.020225f
C379 plus.n52 a_n2354_n4888# 0.308253f
C380 plus.n53 a_n2354_n4888# 0.020225f
C381 plus.n54 a_n2354_n4888# 0.049104f
C382 plus.n55 a_n2354_n4888# 0.049104f
C383 plus.n56 a_n2354_n4888# 0.020225f
C384 plus.n57 a_n2354_n4888# 0.308253f
C385 plus.n58 a_n2354_n4888# 0.018257f
C386 plus.n59 a_n2354_n4888# 0.018257f
C387 plus.n60 a_n2354_n4888# 0.049104f
C388 plus.n61 a_n2354_n4888# 0.049104f
C389 plus.n62 a_n2354_n4888# 0.020225f
C390 plus.n63 a_n2354_n4888# 0.308253f
C391 plus.n64 a_n2354_n4888# 0.020225f
C392 plus.n65 a_n2354_n4888# 0.308253f
C393 plus.n66 a_n2354_n4888# 0.020225f
C394 plus.n67 a_n2354_n4888# 0.049104f
C395 plus.n68 a_n2354_n4888# 0.049104f
C396 plus.n69 a_n2354_n4888# 0.017652f
C397 plus.n70 a_n2354_n4888# 0.018863f
C398 plus.n71 a_n2354_n4888# 0.308253f
C399 plus.n72 a_n2354_n4888# 0.323369f
C400 plus.n73 a_n2354_n4888# 1.85758f
.ends

