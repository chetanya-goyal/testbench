* NGSPICE file created from diffpair43.ext - technology: sky130A

.subckt diffpair43 minus drain_right drain_left source plus
X0 source.t15 minus.t0 drain_right.t6 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X1 source.t2 plus.t0 drain_left.t7 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 drain_right.t0 minus.t1 source.t14 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 source.t13 minus.t2 drain_right.t5 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X5 drain_left.t6 plus.t1 source.t3 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X6 drain_left.t5 plus.t2 source.t5 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X8 a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X9 source.t12 minus.t3 drain_right.t4 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X10 drain_right.t2 minus.t4 source.t11 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X11 drain_left.t4 plus.t3 source.t6 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X12 drain_right.t1 minus.t5 source.t10 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X13 drain_right.t3 minus.t6 source.t9 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 drain_left.t3 plus.t4 source.t0 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X15 source.t7 plus.t5 drain_left.t2 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 source.t8 minus.t7 drain_right.t7 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X17 source.t1 plus.t6 drain_left.t1 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X18 a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X19 source.t4 plus.t7 drain_left.t0 a_n1546_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
R0 minus.n7 minus.n6 161.3
R1 minus.n5 minus.n0 161.3
R2 minus.n4 minus.n3 161.3
R3 minus.n15 minus.n14 161.3
R4 minus.n13 minus.n8 161.3
R5 minus.n12 minus.n11 161.3
R6 minus.n2 minus.t5 147.749
R7 minus.n10 minus.t3 147.749
R8 minus.n1 minus.t0 126.766
R9 minus.n5 minus.t1 126.766
R10 minus.n6 minus.t7 126.766
R11 minus.n9 minus.t6 126.766
R12 minus.n13 minus.t2 126.766
R13 minus.n14 minus.t4 126.766
R14 minus.n3 minus.n2 70.4033
R15 minus.n11 minus.n10 70.4033
R16 minus.n6 minus.n5 48.2005
R17 minus.n14 minus.n13 48.2005
R18 minus.n16 minus.n7 26.7391
R19 minus.n5 minus.n4 24.1005
R20 minus.n4 minus.n1 24.1005
R21 minus.n12 minus.n9 24.1005
R22 minus.n13 minus.n12 24.1005
R23 minus.n2 minus.n1 20.9576
R24 minus.n10 minus.n9 20.9576
R25 minus.n16 minus.n15 6.5952
R26 minus.n7 minus.n0 0.189894
R27 minus.n3 minus.n0 0.189894
R28 minus.n11 minus.n8 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 drain_right.n5 drain_right.n3 240.849
R32 drain_right.n2 drain_right.n1 240.435
R33 drain_right.n2 drain_right.n0 240.435
R34 drain_right.n5 drain_right.n4 240.132
R35 drain_right drain_right.n2 20.9848
R36 drain_right.n1 drain_right.t5 19.8005
R37 drain_right.n1 drain_right.t2 19.8005
R38 drain_right.n0 drain_right.t4 19.8005
R39 drain_right.n0 drain_right.t3 19.8005
R40 drain_right.n3 drain_right.t6 19.8005
R41 drain_right.n3 drain_right.t1 19.8005
R42 drain_right.n4 drain_right.t7 19.8005
R43 drain_right.n4 drain_right.t0 19.8005
R44 drain_right drain_right.n5 6.36873
R45 source.n0 source.t3 243.255
R46 source.n3 source.t2 243.255
R47 source.n4 source.t10 243.255
R48 source.n7 source.t8 243.255
R49 source.n15 source.t11 243.254
R50 source.n12 source.t12 243.254
R51 source.n11 source.t6 243.254
R52 source.n8 source.t1 243.254
R53 source.n2 source.n1 223.454
R54 source.n6 source.n5 223.454
R55 source.n14 source.n13 223.453
R56 source.n10 source.n9 223.453
R57 source.n13 source.t9 19.8005
R58 source.n13 source.t13 19.8005
R59 source.n9 source.t5 19.8005
R60 source.n9 source.t7 19.8005
R61 source.n1 source.t0 19.8005
R62 source.n1 source.t4 19.8005
R63 source.n5 source.t14 19.8005
R64 source.n5 source.t15 19.8005
R65 source.n8 source.n7 13.6699
R66 source.n16 source.n0 8.04922
R67 source.n16 source.n15 5.62119
R68 source.n7 source.n6 0.716017
R69 source.n6 source.n4 0.716017
R70 source.n3 source.n2 0.716017
R71 source.n2 source.n0 0.716017
R72 source.n10 source.n8 0.716017
R73 source.n11 source.n10 0.716017
R74 source.n14 source.n12 0.716017
R75 source.n15 source.n14 0.716017
R76 source.n4 source.n3 0.470328
R77 source.n12 source.n11 0.470328
R78 source source.n16 0.188
R79 plus.n4 plus.n3 161.3
R80 plus.n5 plus.n0 161.3
R81 plus.n7 plus.n6 161.3
R82 plus.n12 plus.n11 161.3
R83 plus.n13 plus.n8 161.3
R84 plus.n15 plus.n14 161.3
R85 plus.n2 plus.t0 147.749
R86 plus.n10 plus.t3 147.749
R87 plus.n6 plus.t1 126.766
R88 plus.n5 plus.t7 126.766
R89 plus.n1 plus.t4 126.766
R90 plus.n14 plus.t6 126.766
R91 plus.n13 plus.t2 126.766
R92 plus.n9 plus.t5 126.766
R93 plus.n3 plus.n2 70.4033
R94 plus.n11 plus.n10 70.4033
R95 plus.n6 plus.n5 48.2005
R96 plus.n14 plus.n13 48.2005
R97 plus plus.n15 24.7869
R98 plus.n4 plus.n1 24.1005
R99 plus.n5 plus.n4 24.1005
R100 plus.n13 plus.n12 24.1005
R101 plus.n12 plus.n9 24.1005
R102 plus.n2 plus.n1 20.9576
R103 plus.n10 plus.n9 20.9576
R104 plus plus.n7 8.07247
R105 plus.n3 plus.n0 0.189894
R106 plus.n7 plus.n0 0.189894
R107 plus.n15 plus.n8 0.189894
R108 plus.n11 plus.n8 0.189894
R109 drain_left.n5 drain_left.n3 240.849
R110 drain_left.n2 drain_left.n1 240.435
R111 drain_left.n2 drain_left.n0 240.435
R112 drain_left.n5 drain_left.n4 240.132
R113 drain_left drain_left.n2 21.538
R114 drain_left.n1 drain_left.t2 19.8005
R115 drain_left.n1 drain_left.t4 19.8005
R116 drain_left.n0 drain_left.t1 19.8005
R117 drain_left.n0 drain_left.t5 19.8005
R118 drain_left.n4 drain_left.t0 19.8005
R119 drain_left.n4 drain_left.t6 19.8005
R120 drain_left.n3 drain_left.t7 19.8005
R121 drain_left.n3 drain_left.t3 19.8005
R122 drain_left drain_left.n5 6.36873
C0 minus plus 3.04382f
C1 source minus 0.99267f
C2 drain_right plus 0.310324f
C3 source drain_right 2.90989f
C4 source plus 1.00653f
C5 minus drain_left 0.178253f
C6 drain_right drain_left 0.727179f
C7 drain_left plus 0.870722f
C8 source drain_left 2.90941f
C9 minus drain_right 0.722741f
C10 drain_right a_n1546_n1088# 2.97287f
C11 drain_left a_n1546_n1088# 3.165308f
C12 source a_n1546_n1088# 2.355083f
C13 minus a_n1546_n1088# 5.057362f
C14 plus a_n1546_n1088# 5.709867f
C15 drain_left.t1 a_n1546_n1088# 0.015837f
C16 drain_left.t5 a_n1546_n1088# 0.015837f
C17 drain_left.n0 a_n1546_n1088# 0.061808f
C18 drain_left.t2 a_n1546_n1088# 0.015837f
C19 drain_left.t4 a_n1546_n1088# 0.015837f
C20 drain_left.n1 a_n1546_n1088# 0.061808f
C21 drain_left.n2 a_n1546_n1088# 0.921232f
C22 drain_left.t7 a_n1546_n1088# 0.015837f
C23 drain_left.t3 a_n1546_n1088# 0.015837f
C24 drain_left.n3 a_n1546_n1088# 0.062252f
C25 drain_left.t0 a_n1546_n1088# 0.015837f
C26 drain_left.t6 a_n1546_n1088# 0.015837f
C27 drain_left.n4 a_n1546_n1088# 0.061537f
C28 drain_left.n5 a_n1546_n1088# 0.64465f
C29 plus.n0 a_n1546_n1088# 0.033292f
C30 plus.t1 a_n1546_n1088# 0.056446f
C31 plus.t7 a_n1546_n1088# 0.056446f
C32 plus.t4 a_n1546_n1088# 0.056446f
C33 plus.n1 a_n1546_n1088# 0.062101f
C34 plus.t0 a_n1546_n1088# 0.064791f
C35 plus.n2 a_n1546_n1088# 0.050625f
C36 plus.n3 a_n1546_n1088# 0.109676f
C37 plus.n4 a_n1546_n1088# 0.007555f
C38 plus.n5 a_n1546_n1088# 0.062101f
C39 plus.n6 a_n1546_n1088# 0.058714f
C40 plus.n7 a_n1546_n1088# 0.236085f
C41 plus.n8 a_n1546_n1088# 0.033292f
C42 plus.t6 a_n1546_n1088# 0.056446f
C43 plus.t2 a_n1546_n1088# 0.056446f
C44 plus.t5 a_n1546_n1088# 0.056446f
C45 plus.n9 a_n1546_n1088# 0.062101f
C46 plus.t3 a_n1546_n1088# 0.064791f
C47 plus.n10 a_n1546_n1088# 0.050625f
C48 plus.n11 a_n1546_n1088# 0.109676f
C49 plus.n12 a_n1546_n1088# 0.007555f
C50 plus.n13 a_n1546_n1088# 0.062101f
C51 plus.n14 a_n1546_n1088# 0.058714f
C52 plus.n15 a_n1546_n1088# 0.691932f
C53 source.t3 a_n1546_n1088# 0.101907f
C54 source.n0 a_n1546_n1088# 0.460599f
C55 source.t0 a_n1546_n1088# 0.018309f
C56 source.t4 a_n1546_n1088# 0.018309f
C57 source.n1 a_n1546_n1088# 0.05938f
C58 source.n2 a_n1546_n1088# 0.249138f
C59 source.t2 a_n1546_n1088# 0.101907f
C60 source.n3 a_n1546_n1088# 0.238203f
C61 source.t10 a_n1546_n1088# 0.101907f
C62 source.n4 a_n1546_n1088# 0.238203f
C63 source.t14 a_n1546_n1088# 0.018309f
C64 source.t15 a_n1546_n1088# 0.018309f
C65 source.n5 a_n1546_n1088# 0.05938f
C66 source.n6 a_n1546_n1088# 0.249138f
C67 source.t8 a_n1546_n1088# 0.101907f
C68 source.n7 a_n1546_n1088# 0.648976f
C69 source.t1 a_n1546_n1088# 0.101907f
C70 source.n8 a_n1546_n1088# 0.648976f
C71 source.t5 a_n1546_n1088# 0.018309f
C72 source.t7 a_n1546_n1088# 0.018309f
C73 source.n9 a_n1546_n1088# 0.05938f
C74 source.n10 a_n1546_n1088# 0.249138f
C75 source.t6 a_n1546_n1088# 0.101907f
C76 source.n11 a_n1546_n1088# 0.238203f
C77 source.t12 a_n1546_n1088# 0.101907f
C78 source.n12 a_n1546_n1088# 0.238203f
C79 source.t9 a_n1546_n1088# 0.018309f
C80 source.t13 a_n1546_n1088# 0.018309f
C81 source.n13 a_n1546_n1088# 0.05938f
C82 source.n14 a_n1546_n1088# 0.249138f
C83 source.t11 a_n1546_n1088# 0.101907f
C84 source.n15 a_n1546_n1088# 0.379224f
C85 source.n16 a_n1546_n1088# 0.474608f
C86 drain_right.t4 a_n1546_n1088# 0.016277f
C87 drain_right.t3 a_n1546_n1088# 0.016277f
C88 drain_right.n0 a_n1546_n1088# 0.063526f
C89 drain_right.t5 a_n1546_n1088# 0.016277f
C90 drain_right.t2 a_n1546_n1088# 0.016277f
C91 drain_right.n1 a_n1546_n1088# 0.063526f
C92 drain_right.n2 a_n1546_n1088# 0.906935f
C93 drain_right.t6 a_n1546_n1088# 0.016277f
C94 drain_right.t1 a_n1546_n1088# 0.016277f
C95 drain_right.n3 a_n1546_n1088# 0.063982f
C96 drain_right.t7 a_n1546_n1088# 0.016277f
C97 drain_right.t0 a_n1546_n1088# 0.016277f
C98 drain_right.n4 a_n1546_n1088# 0.063247f
C99 drain_right.n5 a_n1546_n1088# 0.662561f
C100 minus.n0 a_n1546_n1088# 0.032561f
C101 minus.t0 a_n1546_n1088# 0.055207f
C102 minus.n1 a_n1546_n1088# 0.060737f
C103 minus.t5 a_n1546_n1088# 0.063369f
C104 minus.n2 a_n1546_n1088# 0.049514f
C105 minus.n3 a_n1546_n1088# 0.107269f
C106 minus.n4 a_n1546_n1088# 0.007389f
C107 minus.t1 a_n1546_n1088# 0.055207f
C108 minus.n5 a_n1546_n1088# 0.060737f
C109 minus.t7 a_n1546_n1088# 0.055207f
C110 minus.n6 a_n1546_n1088# 0.057425f
C111 minus.n7 a_n1546_n1088# 0.694977f
C112 minus.n8 a_n1546_n1088# 0.032561f
C113 minus.t6 a_n1546_n1088# 0.055207f
C114 minus.n9 a_n1546_n1088# 0.060737f
C115 minus.t3 a_n1546_n1088# 0.063369f
C116 minus.n10 a_n1546_n1088# 0.049514f
C117 minus.n11 a_n1546_n1088# 0.107269f
C118 minus.n12 a_n1546_n1088# 0.007389f
C119 minus.t2 a_n1546_n1088# 0.055207f
C120 minus.n13 a_n1546_n1088# 0.060737f
C121 minus.t4 a_n1546_n1088# 0.055207f
C122 minus.n14 a_n1546_n1088# 0.057425f
C123 minus.n15 a_n1546_n1088# 0.220146f
C124 minus.n16 a_n1546_n1088# 0.854246f
.ends

