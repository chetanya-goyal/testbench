* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right minus source a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X1 drain_right minus source a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X2 drain_left plus source a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X3 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X4 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5 drain_left plus source a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X6 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7 a_n976_n1092# a_n976_n1092# a_n976_n1092# a_n976_n1092# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
.ends

