* NGSPICE file created from diffpair467.ext - technology: sky130A

.subckt diffpair467 minus drain_right drain_left source plus
X0 a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X1 source.t31 plus.t0 drain_left.t6 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X2 drain_left.t5 plus.t1 source.t30 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X3 source.t29 plus.t2 drain_left.t0 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X4 source.t7 minus.t0 drain_right.t15 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X5 source.t28 plus.t3 drain_left.t9 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X6 source.t8 minus.t1 drain_right.t14 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X7 drain_right.t13 minus.t2 source.t10 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X8 source.t27 plus.t4 drain_left.t1 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X9 source.t26 plus.t5 drain_left.t10 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X10 a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X11 drain_right.t12 minus.t3 source.t6 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X12 a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X13 source.t25 plus.t6 drain_left.t2 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X14 drain_right.t11 minus.t4 source.t15 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X15 drain_left.t11 plus.t7 source.t24 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X16 drain_left.t4 plus.t8 source.t23 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X17 drain_right.t10 minus.t5 source.t2 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X18 drain_left.t7 plus.t9 source.t22 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X19 drain_right.t9 minus.t6 source.t1 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X20 drain_left.t15 plus.t10 source.t21 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X21 drain_right.t8 minus.t7 source.t3 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X22 drain_left.t3 plus.t11 source.t20 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X23 drain_left.t14 plus.t12 source.t19 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X24 drain_right.t7 minus.t8 source.t4 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X25 source.t9 minus.t9 drain_right.t6 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X26 source.t18 plus.t13 drain_left.t12 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X27 source.t11 minus.t10 drain_right.t5 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X28 a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X29 drain_left.t13 plus.t14 source.t17 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X30 source.t0 minus.t11 drain_right.t4 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X31 source.t16 plus.t15 drain_left.t8 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X32 drain_right.t3 minus.t12 source.t13 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X33 source.t12 minus.t13 drain_right.t2 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X34 source.t14 minus.t14 drain_right.t1 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X35 source.t5 minus.t15 drain_right.t0 a_n2570_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
R0 plus.n7 plus.t5 493.637
R1 plus.n33 plus.t14 493.637
R2 plus.n24 plus.t8 469.262
R3 plus.n22 plus.t2 469.262
R4 plus.n2 plus.t10 469.262
R5 plus.n16 plus.t4 469.262
R6 plus.n4 plus.t9 469.262
R7 plus.n10 plus.t3 469.262
R8 plus.n6 plus.t11 469.262
R9 plus.n50 plus.t13 469.262
R10 plus.n48 plus.t1 469.262
R11 plus.n28 plus.t0 469.262
R12 plus.n42 plus.t7 469.262
R13 plus.n30 plus.t6 469.262
R14 plus.n36 plus.t12 469.262
R15 plus.n32 plus.t15 469.262
R16 plus.n9 plus.n8 161.3
R17 plus.n10 plus.n5 161.3
R18 plus.n12 plus.n11 161.3
R19 plus.n13 plus.n4 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n16 plus.n3 161.3
R22 plus.n18 plus.n17 161.3
R23 plus.n19 plus.n2 161.3
R24 plus.n21 plus.n20 161.3
R25 plus.n22 plus.n1 161.3
R26 plus.n23 plus.n0 161.3
R27 plus.n25 plus.n24 161.3
R28 plus.n35 plus.n34 161.3
R29 plus.n36 plus.n31 161.3
R30 plus.n38 plus.n37 161.3
R31 plus.n39 plus.n30 161.3
R32 plus.n41 plus.n40 161.3
R33 plus.n42 plus.n29 161.3
R34 plus.n44 plus.n43 161.3
R35 plus.n45 plus.n28 161.3
R36 plus.n47 plus.n46 161.3
R37 plus.n48 plus.n27 161.3
R38 plus.n49 plus.n26 161.3
R39 plus.n51 plus.n50 161.3
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus plus.n51 32.893
R45 plus.n22 plus.n21 32.8641
R46 plus.n9 plus.n6 32.8641
R47 plus.n48 plus.n47 32.8641
R48 plus.n35 plus.n32 32.8641
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus plus.n25 12.2997
R68 plus.n23 plus.n22 10.955
R69 plus.n49 plus.n48 10.955
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 drain_left.n9 drain_left.n7 60.4406
R93 drain_left.n5 drain_left.n3 60.4404
R94 drain_left.n2 drain_left.n0 60.4404
R95 drain_left.n11 drain_left.n10 59.5527
R96 drain_left.n9 drain_left.n8 59.5527
R97 drain_left.n5 drain_left.n4 59.5525
R98 drain_left.n2 drain_left.n1 59.5525
R99 drain_left.n13 drain_left.n12 59.5525
R100 drain_left drain_left.n6 33.1386
R101 drain_left drain_left.n13 6.54115
R102 drain_left.n3 drain_left.t8 1.6505
R103 drain_left.n3 drain_left.t13 1.6505
R104 drain_left.n4 drain_left.t2 1.6505
R105 drain_left.n4 drain_left.t14 1.6505
R106 drain_left.n1 drain_left.t6 1.6505
R107 drain_left.n1 drain_left.t11 1.6505
R108 drain_left.n0 drain_left.t12 1.6505
R109 drain_left.n0 drain_left.t5 1.6505
R110 drain_left.n12 drain_left.t0 1.6505
R111 drain_left.n12 drain_left.t4 1.6505
R112 drain_left.n10 drain_left.t1 1.6505
R113 drain_left.n10 drain_left.t15 1.6505
R114 drain_left.n8 drain_left.t9 1.6505
R115 drain_left.n8 drain_left.t7 1.6505
R116 drain_left.n7 drain_left.t10 1.6505
R117 drain_left.n7 drain_left.t3 1.6505
R118 drain_left.n11 drain_left.n9 0.888431
R119 drain_left.n13 drain_left.n11 0.888431
R120 drain_left.n6 drain_left.n5 0.389119
R121 drain_left.n6 drain_left.n2 0.389119
R122 source.n546 source.n486 289.615
R123 source.n474 source.n414 289.615
R124 source.n408 source.n348 289.615
R125 source.n336 source.n276 289.615
R126 source.n60 source.n0 289.615
R127 source.n132 source.n72 289.615
R128 source.n198 source.n138 289.615
R129 source.n270 source.n210 289.615
R130 source.n506 source.n505 185
R131 source.n511 source.n510 185
R132 source.n513 source.n512 185
R133 source.n502 source.n501 185
R134 source.n519 source.n518 185
R135 source.n521 source.n520 185
R136 source.n498 source.n497 185
R137 source.n528 source.n527 185
R138 source.n529 source.n496 185
R139 source.n531 source.n530 185
R140 source.n494 source.n493 185
R141 source.n537 source.n536 185
R142 source.n539 source.n538 185
R143 source.n490 source.n489 185
R144 source.n545 source.n544 185
R145 source.n547 source.n546 185
R146 source.n434 source.n433 185
R147 source.n439 source.n438 185
R148 source.n441 source.n440 185
R149 source.n430 source.n429 185
R150 source.n447 source.n446 185
R151 source.n449 source.n448 185
R152 source.n426 source.n425 185
R153 source.n456 source.n455 185
R154 source.n457 source.n424 185
R155 source.n459 source.n458 185
R156 source.n422 source.n421 185
R157 source.n465 source.n464 185
R158 source.n467 source.n466 185
R159 source.n418 source.n417 185
R160 source.n473 source.n472 185
R161 source.n475 source.n474 185
R162 source.n368 source.n367 185
R163 source.n373 source.n372 185
R164 source.n375 source.n374 185
R165 source.n364 source.n363 185
R166 source.n381 source.n380 185
R167 source.n383 source.n382 185
R168 source.n360 source.n359 185
R169 source.n390 source.n389 185
R170 source.n391 source.n358 185
R171 source.n393 source.n392 185
R172 source.n356 source.n355 185
R173 source.n399 source.n398 185
R174 source.n401 source.n400 185
R175 source.n352 source.n351 185
R176 source.n407 source.n406 185
R177 source.n409 source.n408 185
R178 source.n296 source.n295 185
R179 source.n301 source.n300 185
R180 source.n303 source.n302 185
R181 source.n292 source.n291 185
R182 source.n309 source.n308 185
R183 source.n311 source.n310 185
R184 source.n288 source.n287 185
R185 source.n318 source.n317 185
R186 source.n319 source.n286 185
R187 source.n321 source.n320 185
R188 source.n284 source.n283 185
R189 source.n327 source.n326 185
R190 source.n329 source.n328 185
R191 source.n280 source.n279 185
R192 source.n335 source.n334 185
R193 source.n337 source.n336 185
R194 source.n61 source.n60 185
R195 source.n59 source.n58 185
R196 source.n4 source.n3 185
R197 source.n53 source.n52 185
R198 source.n51 source.n50 185
R199 source.n8 source.n7 185
R200 source.n45 source.n44 185
R201 source.n43 source.n10 185
R202 source.n42 source.n41 185
R203 source.n13 source.n11 185
R204 source.n36 source.n35 185
R205 source.n34 source.n33 185
R206 source.n17 source.n16 185
R207 source.n28 source.n27 185
R208 source.n26 source.n25 185
R209 source.n21 source.n20 185
R210 source.n133 source.n132 185
R211 source.n131 source.n130 185
R212 source.n76 source.n75 185
R213 source.n125 source.n124 185
R214 source.n123 source.n122 185
R215 source.n80 source.n79 185
R216 source.n117 source.n116 185
R217 source.n115 source.n82 185
R218 source.n114 source.n113 185
R219 source.n85 source.n83 185
R220 source.n108 source.n107 185
R221 source.n106 source.n105 185
R222 source.n89 source.n88 185
R223 source.n100 source.n99 185
R224 source.n98 source.n97 185
R225 source.n93 source.n92 185
R226 source.n199 source.n198 185
R227 source.n197 source.n196 185
R228 source.n142 source.n141 185
R229 source.n191 source.n190 185
R230 source.n189 source.n188 185
R231 source.n146 source.n145 185
R232 source.n183 source.n182 185
R233 source.n181 source.n148 185
R234 source.n180 source.n179 185
R235 source.n151 source.n149 185
R236 source.n174 source.n173 185
R237 source.n172 source.n171 185
R238 source.n155 source.n154 185
R239 source.n166 source.n165 185
R240 source.n164 source.n163 185
R241 source.n159 source.n158 185
R242 source.n271 source.n270 185
R243 source.n269 source.n268 185
R244 source.n214 source.n213 185
R245 source.n263 source.n262 185
R246 source.n261 source.n260 185
R247 source.n218 source.n217 185
R248 source.n255 source.n254 185
R249 source.n253 source.n220 185
R250 source.n252 source.n251 185
R251 source.n223 source.n221 185
R252 source.n246 source.n245 185
R253 source.n244 source.n243 185
R254 source.n227 source.n226 185
R255 source.n238 source.n237 185
R256 source.n236 source.n235 185
R257 source.n231 source.n230 185
R258 source.n507 source.t1 149.524
R259 source.n435 source.t7 149.524
R260 source.n369 source.t17 149.524
R261 source.n297 source.t18 149.524
R262 source.n22 source.t23 149.524
R263 source.n94 source.t26 149.524
R264 source.n160 source.t3 149.524
R265 source.n232 source.t11 149.524
R266 source.n511 source.n505 104.615
R267 source.n512 source.n511 104.615
R268 source.n512 source.n501 104.615
R269 source.n519 source.n501 104.615
R270 source.n520 source.n519 104.615
R271 source.n520 source.n497 104.615
R272 source.n528 source.n497 104.615
R273 source.n529 source.n528 104.615
R274 source.n530 source.n529 104.615
R275 source.n530 source.n493 104.615
R276 source.n537 source.n493 104.615
R277 source.n538 source.n537 104.615
R278 source.n538 source.n489 104.615
R279 source.n545 source.n489 104.615
R280 source.n546 source.n545 104.615
R281 source.n439 source.n433 104.615
R282 source.n440 source.n439 104.615
R283 source.n440 source.n429 104.615
R284 source.n447 source.n429 104.615
R285 source.n448 source.n447 104.615
R286 source.n448 source.n425 104.615
R287 source.n456 source.n425 104.615
R288 source.n457 source.n456 104.615
R289 source.n458 source.n457 104.615
R290 source.n458 source.n421 104.615
R291 source.n465 source.n421 104.615
R292 source.n466 source.n465 104.615
R293 source.n466 source.n417 104.615
R294 source.n473 source.n417 104.615
R295 source.n474 source.n473 104.615
R296 source.n373 source.n367 104.615
R297 source.n374 source.n373 104.615
R298 source.n374 source.n363 104.615
R299 source.n381 source.n363 104.615
R300 source.n382 source.n381 104.615
R301 source.n382 source.n359 104.615
R302 source.n390 source.n359 104.615
R303 source.n391 source.n390 104.615
R304 source.n392 source.n391 104.615
R305 source.n392 source.n355 104.615
R306 source.n399 source.n355 104.615
R307 source.n400 source.n399 104.615
R308 source.n400 source.n351 104.615
R309 source.n407 source.n351 104.615
R310 source.n408 source.n407 104.615
R311 source.n301 source.n295 104.615
R312 source.n302 source.n301 104.615
R313 source.n302 source.n291 104.615
R314 source.n309 source.n291 104.615
R315 source.n310 source.n309 104.615
R316 source.n310 source.n287 104.615
R317 source.n318 source.n287 104.615
R318 source.n319 source.n318 104.615
R319 source.n320 source.n319 104.615
R320 source.n320 source.n283 104.615
R321 source.n327 source.n283 104.615
R322 source.n328 source.n327 104.615
R323 source.n328 source.n279 104.615
R324 source.n335 source.n279 104.615
R325 source.n336 source.n335 104.615
R326 source.n60 source.n59 104.615
R327 source.n59 source.n3 104.615
R328 source.n52 source.n3 104.615
R329 source.n52 source.n51 104.615
R330 source.n51 source.n7 104.615
R331 source.n44 source.n7 104.615
R332 source.n44 source.n43 104.615
R333 source.n43 source.n42 104.615
R334 source.n42 source.n11 104.615
R335 source.n35 source.n11 104.615
R336 source.n35 source.n34 104.615
R337 source.n34 source.n16 104.615
R338 source.n27 source.n16 104.615
R339 source.n27 source.n26 104.615
R340 source.n26 source.n20 104.615
R341 source.n132 source.n131 104.615
R342 source.n131 source.n75 104.615
R343 source.n124 source.n75 104.615
R344 source.n124 source.n123 104.615
R345 source.n123 source.n79 104.615
R346 source.n116 source.n79 104.615
R347 source.n116 source.n115 104.615
R348 source.n115 source.n114 104.615
R349 source.n114 source.n83 104.615
R350 source.n107 source.n83 104.615
R351 source.n107 source.n106 104.615
R352 source.n106 source.n88 104.615
R353 source.n99 source.n88 104.615
R354 source.n99 source.n98 104.615
R355 source.n98 source.n92 104.615
R356 source.n198 source.n197 104.615
R357 source.n197 source.n141 104.615
R358 source.n190 source.n141 104.615
R359 source.n190 source.n189 104.615
R360 source.n189 source.n145 104.615
R361 source.n182 source.n145 104.615
R362 source.n182 source.n181 104.615
R363 source.n181 source.n180 104.615
R364 source.n180 source.n149 104.615
R365 source.n173 source.n149 104.615
R366 source.n173 source.n172 104.615
R367 source.n172 source.n154 104.615
R368 source.n165 source.n154 104.615
R369 source.n165 source.n164 104.615
R370 source.n164 source.n158 104.615
R371 source.n270 source.n269 104.615
R372 source.n269 source.n213 104.615
R373 source.n262 source.n213 104.615
R374 source.n262 source.n261 104.615
R375 source.n261 source.n217 104.615
R376 source.n254 source.n217 104.615
R377 source.n254 source.n253 104.615
R378 source.n253 source.n252 104.615
R379 source.n252 source.n221 104.615
R380 source.n245 source.n221 104.615
R381 source.n245 source.n244 104.615
R382 source.n244 source.n226 104.615
R383 source.n237 source.n226 104.615
R384 source.n237 source.n236 104.615
R385 source.n236 source.n230 104.615
R386 source.t1 source.n505 52.3082
R387 source.t7 source.n433 52.3082
R388 source.t17 source.n367 52.3082
R389 source.t18 source.n295 52.3082
R390 source.t23 source.n20 52.3082
R391 source.t26 source.n92 52.3082
R392 source.t3 source.n158 52.3082
R393 source.t11 source.n230 52.3082
R394 source.n67 source.n66 42.8739
R395 source.n69 source.n68 42.8739
R396 source.n71 source.n70 42.8739
R397 source.n205 source.n204 42.8739
R398 source.n207 source.n206 42.8739
R399 source.n209 source.n208 42.8739
R400 source.n485 source.n484 42.8737
R401 source.n483 source.n482 42.8737
R402 source.n481 source.n480 42.8737
R403 source.n347 source.n346 42.8737
R404 source.n345 source.n344 42.8737
R405 source.n343 source.n342 42.8737
R406 source.n551 source.n550 29.8581
R407 source.n479 source.n478 29.8581
R408 source.n413 source.n412 29.8581
R409 source.n341 source.n340 29.8581
R410 source.n65 source.n64 29.8581
R411 source.n137 source.n136 29.8581
R412 source.n203 source.n202 29.8581
R413 source.n275 source.n274 29.8581
R414 source.n341 source.n275 22.1757
R415 source.n552 source.n65 16.4688
R416 source.n531 source.n496 13.1884
R417 source.n459 source.n424 13.1884
R418 source.n393 source.n358 13.1884
R419 source.n321 source.n286 13.1884
R420 source.n45 source.n10 13.1884
R421 source.n117 source.n82 13.1884
R422 source.n183 source.n148 13.1884
R423 source.n255 source.n220 13.1884
R424 source.n527 source.n526 12.8005
R425 source.n532 source.n494 12.8005
R426 source.n455 source.n454 12.8005
R427 source.n460 source.n422 12.8005
R428 source.n389 source.n388 12.8005
R429 source.n394 source.n356 12.8005
R430 source.n317 source.n316 12.8005
R431 source.n322 source.n284 12.8005
R432 source.n46 source.n8 12.8005
R433 source.n41 source.n12 12.8005
R434 source.n118 source.n80 12.8005
R435 source.n113 source.n84 12.8005
R436 source.n184 source.n146 12.8005
R437 source.n179 source.n150 12.8005
R438 source.n256 source.n218 12.8005
R439 source.n251 source.n222 12.8005
R440 source.n525 source.n498 12.0247
R441 source.n536 source.n535 12.0247
R442 source.n453 source.n426 12.0247
R443 source.n464 source.n463 12.0247
R444 source.n387 source.n360 12.0247
R445 source.n398 source.n397 12.0247
R446 source.n315 source.n288 12.0247
R447 source.n326 source.n325 12.0247
R448 source.n50 source.n49 12.0247
R449 source.n40 source.n13 12.0247
R450 source.n122 source.n121 12.0247
R451 source.n112 source.n85 12.0247
R452 source.n188 source.n187 12.0247
R453 source.n178 source.n151 12.0247
R454 source.n260 source.n259 12.0247
R455 source.n250 source.n223 12.0247
R456 source.n522 source.n521 11.249
R457 source.n539 source.n492 11.249
R458 source.n450 source.n449 11.249
R459 source.n467 source.n420 11.249
R460 source.n384 source.n383 11.249
R461 source.n401 source.n354 11.249
R462 source.n312 source.n311 11.249
R463 source.n329 source.n282 11.249
R464 source.n53 source.n6 11.249
R465 source.n37 source.n36 11.249
R466 source.n125 source.n78 11.249
R467 source.n109 source.n108 11.249
R468 source.n191 source.n144 11.249
R469 source.n175 source.n174 11.249
R470 source.n263 source.n216 11.249
R471 source.n247 source.n246 11.249
R472 source.n518 source.n500 10.4732
R473 source.n540 source.n490 10.4732
R474 source.n446 source.n428 10.4732
R475 source.n468 source.n418 10.4732
R476 source.n380 source.n362 10.4732
R477 source.n402 source.n352 10.4732
R478 source.n308 source.n290 10.4732
R479 source.n330 source.n280 10.4732
R480 source.n54 source.n4 10.4732
R481 source.n33 source.n15 10.4732
R482 source.n126 source.n76 10.4732
R483 source.n105 source.n87 10.4732
R484 source.n192 source.n142 10.4732
R485 source.n171 source.n153 10.4732
R486 source.n264 source.n214 10.4732
R487 source.n243 source.n225 10.4732
R488 source.n507 source.n506 10.2747
R489 source.n435 source.n434 10.2747
R490 source.n369 source.n368 10.2747
R491 source.n297 source.n296 10.2747
R492 source.n22 source.n21 10.2747
R493 source.n94 source.n93 10.2747
R494 source.n160 source.n159 10.2747
R495 source.n232 source.n231 10.2747
R496 source.n517 source.n502 9.69747
R497 source.n544 source.n543 9.69747
R498 source.n445 source.n430 9.69747
R499 source.n472 source.n471 9.69747
R500 source.n379 source.n364 9.69747
R501 source.n406 source.n405 9.69747
R502 source.n307 source.n292 9.69747
R503 source.n334 source.n333 9.69747
R504 source.n58 source.n57 9.69747
R505 source.n32 source.n17 9.69747
R506 source.n130 source.n129 9.69747
R507 source.n104 source.n89 9.69747
R508 source.n196 source.n195 9.69747
R509 source.n170 source.n155 9.69747
R510 source.n268 source.n267 9.69747
R511 source.n242 source.n227 9.69747
R512 source.n550 source.n549 9.45567
R513 source.n478 source.n477 9.45567
R514 source.n412 source.n411 9.45567
R515 source.n340 source.n339 9.45567
R516 source.n64 source.n63 9.45567
R517 source.n136 source.n135 9.45567
R518 source.n202 source.n201 9.45567
R519 source.n274 source.n273 9.45567
R520 source.n549 source.n548 9.3005
R521 source.n488 source.n487 9.3005
R522 source.n543 source.n542 9.3005
R523 source.n541 source.n540 9.3005
R524 source.n492 source.n491 9.3005
R525 source.n535 source.n534 9.3005
R526 source.n533 source.n532 9.3005
R527 source.n509 source.n508 9.3005
R528 source.n504 source.n503 9.3005
R529 source.n515 source.n514 9.3005
R530 source.n517 source.n516 9.3005
R531 source.n500 source.n499 9.3005
R532 source.n523 source.n522 9.3005
R533 source.n525 source.n524 9.3005
R534 source.n526 source.n495 9.3005
R535 source.n477 source.n476 9.3005
R536 source.n416 source.n415 9.3005
R537 source.n471 source.n470 9.3005
R538 source.n469 source.n468 9.3005
R539 source.n420 source.n419 9.3005
R540 source.n463 source.n462 9.3005
R541 source.n461 source.n460 9.3005
R542 source.n437 source.n436 9.3005
R543 source.n432 source.n431 9.3005
R544 source.n443 source.n442 9.3005
R545 source.n445 source.n444 9.3005
R546 source.n428 source.n427 9.3005
R547 source.n451 source.n450 9.3005
R548 source.n453 source.n452 9.3005
R549 source.n454 source.n423 9.3005
R550 source.n411 source.n410 9.3005
R551 source.n350 source.n349 9.3005
R552 source.n405 source.n404 9.3005
R553 source.n403 source.n402 9.3005
R554 source.n354 source.n353 9.3005
R555 source.n397 source.n396 9.3005
R556 source.n395 source.n394 9.3005
R557 source.n371 source.n370 9.3005
R558 source.n366 source.n365 9.3005
R559 source.n377 source.n376 9.3005
R560 source.n379 source.n378 9.3005
R561 source.n362 source.n361 9.3005
R562 source.n385 source.n384 9.3005
R563 source.n387 source.n386 9.3005
R564 source.n388 source.n357 9.3005
R565 source.n339 source.n338 9.3005
R566 source.n278 source.n277 9.3005
R567 source.n333 source.n332 9.3005
R568 source.n331 source.n330 9.3005
R569 source.n282 source.n281 9.3005
R570 source.n325 source.n324 9.3005
R571 source.n323 source.n322 9.3005
R572 source.n299 source.n298 9.3005
R573 source.n294 source.n293 9.3005
R574 source.n305 source.n304 9.3005
R575 source.n307 source.n306 9.3005
R576 source.n290 source.n289 9.3005
R577 source.n313 source.n312 9.3005
R578 source.n315 source.n314 9.3005
R579 source.n316 source.n285 9.3005
R580 source.n24 source.n23 9.3005
R581 source.n19 source.n18 9.3005
R582 source.n30 source.n29 9.3005
R583 source.n32 source.n31 9.3005
R584 source.n15 source.n14 9.3005
R585 source.n38 source.n37 9.3005
R586 source.n40 source.n39 9.3005
R587 source.n12 source.n9 9.3005
R588 source.n63 source.n62 9.3005
R589 source.n2 source.n1 9.3005
R590 source.n57 source.n56 9.3005
R591 source.n55 source.n54 9.3005
R592 source.n6 source.n5 9.3005
R593 source.n49 source.n48 9.3005
R594 source.n47 source.n46 9.3005
R595 source.n96 source.n95 9.3005
R596 source.n91 source.n90 9.3005
R597 source.n102 source.n101 9.3005
R598 source.n104 source.n103 9.3005
R599 source.n87 source.n86 9.3005
R600 source.n110 source.n109 9.3005
R601 source.n112 source.n111 9.3005
R602 source.n84 source.n81 9.3005
R603 source.n135 source.n134 9.3005
R604 source.n74 source.n73 9.3005
R605 source.n129 source.n128 9.3005
R606 source.n127 source.n126 9.3005
R607 source.n78 source.n77 9.3005
R608 source.n121 source.n120 9.3005
R609 source.n119 source.n118 9.3005
R610 source.n162 source.n161 9.3005
R611 source.n157 source.n156 9.3005
R612 source.n168 source.n167 9.3005
R613 source.n170 source.n169 9.3005
R614 source.n153 source.n152 9.3005
R615 source.n176 source.n175 9.3005
R616 source.n178 source.n177 9.3005
R617 source.n150 source.n147 9.3005
R618 source.n201 source.n200 9.3005
R619 source.n140 source.n139 9.3005
R620 source.n195 source.n194 9.3005
R621 source.n193 source.n192 9.3005
R622 source.n144 source.n143 9.3005
R623 source.n187 source.n186 9.3005
R624 source.n185 source.n184 9.3005
R625 source.n234 source.n233 9.3005
R626 source.n229 source.n228 9.3005
R627 source.n240 source.n239 9.3005
R628 source.n242 source.n241 9.3005
R629 source.n225 source.n224 9.3005
R630 source.n248 source.n247 9.3005
R631 source.n250 source.n249 9.3005
R632 source.n222 source.n219 9.3005
R633 source.n273 source.n272 9.3005
R634 source.n212 source.n211 9.3005
R635 source.n267 source.n266 9.3005
R636 source.n265 source.n264 9.3005
R637 source.n216 source.n215 9.3005
R638 source.n259 source.n258 9.3005
R639 source.n257 source.n256 9.3005
R640 source.n514 source.n513 8.92171
R641 source.n547 source.n488 8.92171
R642 source.n442 source.n441 8.92171
R643 source.n475 source.n416 8.92171
R644 source.n376 source.n375 8.92171
R645 source.n409 source.n350 8.92171
R646 source.n304 source.n303 8.92171
R647 source.n337 source.n278 8.92171
R648 source.n61 source.n2 8.92171
R649 source.n29 source.n28 8.92171
R650 source.n133 source.n74 8.92171
R651 source.n101 source.n100 8.92171
R652 source.n199 source.n140 8.92171
R653 source.n167 source.n166 8.92171
R654 source.n271 source.n212 8.92171
R655 source.n239 source.n238 8.92171
R656 source.n510 source.n504 8.14595
R657 source.n548 source.n486 8.14595
R658 source.n438 source.n432 8.14595
R659 source.n476 source.n414 8.14595
R660 source.n372 source.n366 8.14595
R661 source.n410 source.n348 8.14595
R662 source.n300 source.n294 8.14595
R663 source.n338 source.n276 8.14595
R664 source.n62 source.n0 8.14595
R665 source.n25 source.n19 8.14595
R666 source.n134 source.n72 8.14595
R667 source.n97 source.n91 8.14595
R668 source.n200 source.n138 8.14595
R669 source.n163 source.n157 8.14595
R670 source.n272 source.n210 8.14595
R671 source.n235 source.n229 8.14595
R672 source.n509 source.n506 7.3702
R673 source.n437 source.n434 7.3702
R674 source.n371 source.n368 7.3702
R675 source.n299 source.n296 7.3702
R676 source.n24 source.n21 7.3702
R677 source.n96 source.n93 7.3702
R678 source.n162 source.n159 7.3702
R679 source.n234 source.n231 7.3702
R680 source.n510 source.n509 5.81868
R681 source.n550 source.n486 5.81868
R682 source.n438 source.n437 5.81868
R683 source.n478 source.n414 5.81868
R684 source.n372 source.n371 5.81868
R685 source.n412 source.n348 5.81868
R686 source.n300 source.n299 5.81868
R687 source.n340 source.n276 5.81868
R688 source.n64 source.n0 5.81868
R689 source.n25 source.n24 5.81868
R690 source.n136 source.n72 5.81868
R691 source.n97 source.n96 5.81868
R692 source.n202 source.n138 5.81868
R693 source.n163 source.n162 5.81868
R694 source.n274 source.n210 5.81868
R695 source.n235 source.n234 5.81868
R696 source.n552 source.n551 5.7074
R697 source.n513 source.n504 5.04292
R698 source.n548 source.n547 5.04292
R699 source.n441 source.n432 5.04292
R700 source.n476 source.n475 5.04292
R701 source.n375 source.n366 5.04292
R702 source.n410 source.n409 5.04292
R703 source.n303 source.n294 5.04292
R704 source.n338 source.n337 5.04292
R705 source.n62 source.n61 5.04292
R706 source.n28 source.n19 5.04292
R707 source.n134 source.n133 5.04292
R708 source.n100 source.n91 5.04292
R709 source.n200 source.n199 5.04292
R710 source.n166 source.n157 5.04292
R711 source.n272 source.n271 5.04292
R712 source.n238 source.n229 5.04292
R713 source.n514 source.n502 4.26717
R714 source.n544 source.n488 4.26717
R715 source.n442 source.n430 4.26717
R716 source.n472 source.n416 4.26717
R717 source.n376 source.n364 4.26717
R718 source.n406 source.n350 4.26717
R719 source.n304 source.n292 4.26717
R720 source.n334 source.n278 4.26717
R721 source.n58 source.n2 4.26717
R722 source.n29 source.n17 4.26717
R723 source.n130 source.n74 4.26717
R724 source.n101 source.n89 4.26717
R725 source.n196 source.n140 4.26717
R726 source.n167 source.n155 4.26717
R727 source.n268 source.n212 4.26717
R728 source.n239 source.n227 4.26717
R729 source.n518 source.n517 3.49141
R730 source.n543 source.n490 3.49141
R731 source.n446 source.n445 3.49141
R732 source.n471 source.n418 3.49141
R733 source.n380 source.n379 3.49141
R734 source.n405 source.n352 3.49141
R735 source.n308 source.n307 3.49141
R736 source.n333 source.n280 3.49141
R737 source.n57 source.n4 3.49141
R738 source.n33 source.n32 3.49141
R739 source.n129 source.n76 3.49141
R740 source.n105 source.n104 3.49141
R741 source.n195 source.n142 3.49141
R742 source.n171 source.n170 3.49141
R743 source.n267 source.n214 3.49141
R744 source.n243 source.n242 3.49141
R745 source.n508 source.n507 2.84303
R746 source.n436 source.n435 2.84303
R747 source.n370 source.n369 2.84303
R748 source.n298 source.n297 2.84303
R749 source.n23 source.n22 2.84303
R750 source.n95 source.n94 2.84303
R751 source.n161 source.n160 2.84303
R752 source.n233 source.n232 2.84303
R753 source.n521 source.n500 2.71565
R754 source.n540 source.n539 2.71565
R755 source.n449 source.n428 2.71565
R756 source.n468 source.n467 2.71565
R757 source.n383 source.n362 2.71565
R758 source.n402 source.n401 2.71565
R759 source.n311 source.n290 2.71565
R760 source.n330 source.n329 2.71565
R761 source.n54 source.n53 2.71565
R762 source.n36 source.n15 2.71565
R763 source.n126 source.n125 2.71565
R764 source.n108 source.n87 2.71565
R765 source.n192 source.n191 2.71565
R766 source.n174 source.n153 2.71565
R767 source.n264 source.n263 2.71565
R768 source.n246 source.n225 2.71565
R769 source.n522 source.n498 1.93989
R770 source.n536 source.n492 1.93989
R771 source.n450 source.n426 1.93989
R772 source.n464 source.n420 1.93989
R773 source.n384 source.n360 1.93989
R774 source.n398 source.n354 1.93989
R775 source.n312 source.n288 1.93989
R776 source.n326 source.n282 1.93989
R777 source.n50 source.n6 1.93989
R778 source.n37 source.n13 1.93989
R779 source.n122 source.n78 1.93989
R780 source.n109 source.n85 1.93989
R781 source.n188 source.n144 1.93989
R782 source.n175 source.n151 1.93989
R783 source.n260 source.n216 1.93989
R784 source.n247 source.n223 1.93989
R785 source.n484 source.t4 1.6505
R786 source.n484 source.t9 1.6505
R787 source.n482 source.t13 1.6505
R788 source.n482 source.t5 1.6505
R789 source.n480 source.t10 1.6505
R790 source.n480 source.t0 1.6505
R791 source.n346 source.t19 1.6505
R792 source.n346 source.t16 1.6505
R793 source.n344 source.t24 1.6505
R794 source.n344 source.t25 1.6505
R795 source.n342 source.t30 1.6505
R796 source.n342 source.t31 1.6505
R797 source.n66 source.t21 1.6505
R798 source.n66 source.t29 1.6505
R799 source.n68 source.t22 1.6505
R800 source.n68 source.t27 1.6505
R801 source.n70 source.t20 1.6505
R802 source.n70 source.t28 1.6505
R803 source.n204 source.t2 1.6505
R804 source.n204 source.t8 1.6505
R805 source.n206 source.t15 1.6505
R806 source.n206 source.t12 1.6505
R807 source.n208 source.t6 1.6505
R808 source.n208 source.t14 1.6505
R809 source.n527 source.n525 1.16414
R810 source.n535 source.n494 1.16414
R811 source.n455 source.n453 1.16414
R812 source.n463 source.n422 1.16414
R813 source.n389 source.n387 1.16414
R814 source.n397 source.n356 1.16414
R815 source.n317 source.n315 1.16414
R816 source.n325 source.n284 1.16414
R817 source.n49 source.n8 1.16414
R818 source.n41 source.n40 1.16414
R819 source.n121 source.n80 1.16414
R820 source.n113 source.n112 1.16414
R821 source.n187 source.n146 1.16414
R822 source.n179 source.n178 1.16414
R823 source.n259 source.n218 1.16414
R824 source.n251 source.n250 1.16414
R825 source.n275 source.n209 0.888431
R826 source.n209 source.n207 0.888431
R827 source.n207 source.n205 0.888431
R828 source.n205 source.n203 0.888431
R829 source.n137 source.n71 0.888431
R830 source.n71 source.n69 0.888431
R831 source.n69 source.n67 0.888431
R832 source.n67 source.n65 0.888431
R833 source.n343 source.n341 0.888431
R834 source.n345 source.n343 0.888431
R835 source.n347 source.n345 0.888431
R836 source.n413 source.n347 0.888431
R837 source.n481 source.n479 0.888431
R838 source.n483 source.n481 0.888431
R839 source.n485 source.n483 0.888431
R840 source.n551 source.n485 0.888431
R841 source.n203 source.n137 0.470328
R842 source.n479 source.n413 0.470328
R843 source.n526 source.n496 0.388379
R844 source.n532 source.n531 0.388379
R845 source.n454 source.n424 0.388379
R846 source.n460 source.n459 0.388379
R847 source.n388 source.n358 0.388379
R848 source.n394 source.n393 0.388379
R849 source.n316 source.n286 0.388379
R850 source.n322 source.n321 0.388379
R851 source.n46 source.n45 0.388379
R852 source.n12 source.n10 0.388379
R853 source.n118 source.n117 0.388379
R854 source.n84 source.n82 0.388379
R855 source.n184 source.n183 0.388379
R856 source.n150 source.n148 0.388379
R857 source.n256 source.n255 0.388379
R858 source.n222 source.n220 0.388379
R859 source source.n552 0.188
R860 source.n508 source.n503 0.155672
R861 source.n515 source.n503 0.155672
R862 source.n516 source.n515 0.155672
R863 source.n516 source.n499 0.155672
R864 source.n523 source.n499 0.155672
R865 source.n524 source.n523 0.155672
R866 source.n524 source.n495 0.155672
R867 source.n533 source.n495 0.155672
R868 source.n534 source.n533 0.155672
R869 source.n534 source.n491 0.155672
R870 source.n541 source.n491 0.155672
R871 source.n542 source.n541 0.155672
R872 source.n542 source.n487 0.155672
R873 source.n549 source.n487 0.155672
R874 source.n436 source.n431 0.155672
R875 source.n443 source.n431 0.155672
R876 source.n444 source.n443 0.155672
R877 source.n444 source.n427 0.155672
R878 source.n451 source.n427 0.155672
R879 source.n452 source.n451 0.155672
R880 source.n452 source.n423 0.155672
R881 source.n461 source.n423 0.155672
R882 source.n462 source.n461 0.155672
R883 source.n462 source.n419 0.155672
R884 source.n469 source.n419 0.155672
R885 source.n470 source.n469 0.155672
R886 source.n470 source.n415 0.155672
R887 source.n477 source.n415 0.155672
R888 source.n370 source.n365 0.155672
R889 source.n377 source.n365 0.155672
R890 source.n378 source.n377 0.155672
R891 source.n378 source.n361 0.155672
R892 source.n385 source.n361 0.155672
R893 source.n386 source.n385 0.155672
R894 source.n386 source.n357 0.155672
R895 source.n395 source.n357 0.155672
R896 source.n396 source.n395 0.155672
R897 source.n396 source.n353 0.155672
R898 source.n403 source.n353 0.155672
R899 source.n404 source.n403 0.155672
R900 source.n404 source.n349 0.155672
R901 source.n411 source.n349 0.155672
R902 source.n298 source.n293 0.155672
R903 source.n305 source.n293 0.155672
R904 source.n306 source.n305 0.155672
R905 source.n306 source.n289 0.155672
R906 source.n313 source.n289 0.155672
R907 source.n314 source.n313 0.155672
R908 source.n314 source.n285 0.155672
R909 source.n323 source.n285 0.155672
R910 source.n324 source.n323 0.155672
R911 source.n324 source.n281 0.155672
R912 source.n331 source.n281 0.155672
R913 source.n332 source.n331 0.155672
R914 source.n332 source.n277 0.155672
R915 source.n339 source.n277 0.155672
R916 source.n63 source.n1 0.155672
R917 source.n56 source.n1 0.155672
R918 source.n56 source.n55 0.155672
R919 source.n55 source.n5 0.155672
R920 source.n48 source.n5 0.155672
R921 source.n48 source.n47 0.155672
R922 source.n47 source.n9 0.155672
R923 source.n39 source.n9 0.155672
R924 source.n39 source.n38 0.155672
R925 source.n38 source.n14 0.155672
R926 source.n31 source.n14 0.155672
R927 source.n31 source.n30 0.155672
R928 source.n30 source.n18 0.155672
R929 source.n23 source.n18 0.155672
R930 source.n135 source.n73 0.155672
R931 source.n128 source.n73 0.155672
R932 source.n128 source.n127 0.155672
R933 source.n127 source.n77 0.155672
R934 source.n120 source.n77 0.155672
R935 source.n120 source.n119 0.155672
R936 source.n119 source.n81 0.155672
R937 source.n111 source.n81 0.155672
R938 source.n111 source.n110 0.155672
R939 source.n110 source.n86 0.155672
R940 source.n103 source.n86 0.155672
R941 source.n103 source.n102 0.155672
R942 source.n102 source.n90 0.155672
R943 source.n95 source.n90 0.155672
R944 source.n201 source.n139 0.155672
R945 source.n194 source.n139 0.155672
R946 source.n194 source.n193 0.155672
R947 source.n193 source.n143 0.155672
R948 source.n186 source.n143 0.155672
R949 source.n186 source.n185 0.155672
R950 source.n185 source.n147 0.155672
R951 source.n177 source.n147 0.155672
R952 source.n177 source.n176 0.155672
R953 source.n176 source.n152 0.155672
R954 source.n169 source.n152 0.155672
R955 source.n169 source.n168 0.155672
R956 source.n168 source.n156 0.155672
R957 source.n161 source.n156 0.155672
R958 source.n273 source.n211 0.155672
R959 source.n266 source.n211 0.155672
R960 source.n266 source.n265 0.155672
R961 source.n265 source.n215 0.155672
R962 source.n258 source.n215 0.155672
R963 source.n258 source.n257 0.155672
R964 source.n257 source.n219 0.155672
R965 source.n249 source.n219 0.155672
R966 source.n249 source.n248 0.155672
R967 source.n248 source.n224 0.155672
R968 source.n241 source.n224 0.155672
R969 source.n241 source.n240 0.155672
R970 source.n240 source.n228 0.155672
R971 source.n233 source.n228 0.155672
R972 minus.n7 minus.t7 493.637
R973 minus.n33 minus.t0 493.637
R974 minus.n6 minus.t1 469.262
R975 minus.n10 minus.t5 469.262
R976 minus.n12 minus.t13 469.262
R977 minus.n16 minus.t4 469.262
R978 minus.n18 minus.t14 469.262
R979 minus.n22 minus.t3 469.262
R980 minus.n24 minus.t10 469.262
R981 minus.n32 minus.t2 469.262
R982 minus.n36 minus.t11 469.262
R983 minus.n38 minus.t12 469.262
R984 minus.n42 minus.t15 469.262
R985 minus.n44 minus.t8 469.262
R986 minus.n48 minus.t9 469.262
R987 minus.n50 minus.t6 469.262
R988 minus.n25 minus.n24 161.3
R989 minus.n23 minus.n0 161.3
R990 minus.n22 minus.n21 161.3
R991 minus.n20 minus.n1 161.3
R992 minus.n19 minus.n18 161.3
R993 minus.n17 minus.n2 161.3
R994 minus.n16 minus.n15 161.3
R995 minus.n14 minus.n3 161.3
R996 minus.n13 minus.n12 161.3
R997 minus.n11 minus.n4 161.3
R998 minus.n10 minus.n9 161.3
R999 minus.n8 minus.n5 161.3
R1000 minus.n51 minus.n50 161.3
R1001 minus.n49 minus.n26 161.3
R1002 minus.n48 minus.n47 161.3
R1003 minus.n46 minus.n27 161.3
R1004 minus.n45 minus.n44 161.3
R1005 minus.n43 minus.n28 161.3
R1006 minus.n42 minus.n41 161.3
R1007 minus.n40 minus.n29 161.3
R1008 minus.n39 minus.n38 161.3
R1009 minus.n37 minus.n30 161.3
R1010 minus.n36 minus.n35 161.3
R1011 minus.n34 minus.n31 161.3
R1012 minus.n8 minus.n7 44.9377
R1013 minus.n34 minus.n33 44.9377
R1014 minus.n52 minus.n25 39.0119
R1015 minus.n24 minus.n23 37.246
R1016 minus.n50 minus.n49 37.246
R1017 minus.n6 minus.n5 32.8641
R1018 minus.n22 minus.n1 32.8641
R1019 minus.n32 minus.n31 32.8641
R1020 minus.n48 minus.n27 32.8641
R1021 minus.n11 minus.n10 28.4823
R1022 minus.n18 minus.n17 28.4823
R1023 minus.n37 minus.n36 28.4823
R1024 minus.n44 minus.n43 28.4823
R1025 minus.n16 minus.n3 24.1005
R1026 minus.n12 minus.n3 24.1005
R1027 minus.n38 minus.n29 24.1005
R1028 minus.n42 minus.n29 24.1005
R1029 minus.n12 minus.n11 19.7187
R1030 minus.n17 minus.n16 19.7187
R1031 minus.n38 minus.n37 19.7187
R1032 minus.n43 minus.n42 19.7187
R1033 minus.n7 minus.n6 17.0522
R1034 minus.n33 minus.n32 17.0522
R1035 minus.n10 minus.n5 15.3369
R1036 minus.n18 minus.n1 15.3369
R1037 minus.n36 minus.n31 15.3369
R1038 minus.n44 minus.n27 15.3369
R1039 minus.n23 minus.n22 10.955
R1040 minus.n49 minus.n48 10.955
R1041 minus.n52 minus.n51 6.6558
R1042 minus.n25 minus.n0 0.189894
R1043 minus.n21 minus.n0 0.189894
R1044 minus.n21 minus.n20 0.189894
R1045 minus.n20 minus.n19 0.189894
R1046 minus.n19 minus.n2 0.189894
R1047 minus.n15 minus.n2 0.189894
R1048 minus.n15 minus.n14 0.189894
R1049 minus.n14 minus.n13 0.189894
R1050 minus.n13 minus.n4 0.189894
R1051 minus.n9 minus.n4 0.189894
R1052 minus.n9 minus.n8 0.189894
R1053 minus.n35 minus.n34 0.189894
R1054 minus.n35 minus.n30 0.189894
R1055 minus.n39 minus.n30 0.189894
R1056 minus.n40 minus.n39 0.189894
R1057 minus.n41 minus.n40 0.189894
R1058 minus.n41 minus.n28 0.189894
R1059 minus.n45 minus.n28 0.189894
R1060 minus.n46 minus.n45 0.189894
R1061 minus.n47 minus.n46 0.189894
R1062 minus.n47 minus.n26 0.189894
R1063 minus.n51 minus.n26 0.189894
R1064 minus minus.n52 0.188
R1065 drain_right.n5 drain_right.n3 60.4404
R1066 drain_right.n2 drain_right.n0 60.4404
R1067 drain_right.n9 drain_right.n7 60.4404
R1068 drain_right.n9 drain_right.n8 59.5527
R1069 drain_right.n11 drain_right.n10 59.5527
R1070 drain_right.n13 drain_right.n12 59.5527
R1071 drain_right.n5 drain_right.n4 59.5525
R1072 drain_right.n2 drain_right.n1 59.5525
R1073 drain_right drain_right.n6 32.5854
R1074 drain_right drain_right.n13 6.54115
R1075 drain_right.n3 drain_right.t6 1.6505
R1076 drain_right.n3 drain_right.t9 1.6505
R1077 drain_right.n4 drain_right.t0 1.6505
R1078 drain_right.n4 drain_right.t7 1.6505
R1079 drain_right.n1 drain_right.t4 1.6505
R1080 drain_right.n1 drain_right.t3 1.6505
R1081 drain_right.n0 drain_right.t15 1.6505
R1082 drain_right.n0 drain_right.t13 1.6505
R1083 drain_right.n7 drain_right.t14 1.6505
R1084 drain_right.n7 drain_right.t8 1.6505
R1085 drain_right.n8 drain_right.t2 1.6505
R1086 drain_right.n8 drain_right.t10 1.6505
R1087 drain_right.n10 drain_right.t1 1.6505
R1088 drain_right.n10 drain_right.t11 1.6505
R1089 drain_right.n12 drain_right.t5 1.6505
R1090 drain_right.n12 drain_right.t12 1.6505
R1091 drain_right.n13 drain_right.n11 0.888431
R1092 drain_right.n11 drain_right.n9 0.888431
R1093 drain_right.n6 drain_right.n5 0.389119
R1094 drain_right.n6 drain_right.n2 0.389119
C0 drain_left source 19.7937f
C1 minus source 10.265f
C2 plus drain_left 10.4935f
C3 drain_right source 19.7959f
C4 minus plus 6.35016f
C5 drain_right plus 0.410755f
C6 minus drain_left 0.172697f
C7 plus source 10.279099f
C8 drain_right drain_left 1.34352f
C9 drain_right minus 10.2388f
C10 drain_right a_n2570_n3288# 6.78093f
C11 drain_left a_n2570_n3288# 7.15042f
C12 source a_n2570_n3288# 9.260922f
C13 minus a_n2570_n3288# 10.255851f
C14 plus a_n2570_n3288# 12.01726f
C15 drain_right.t15 a_n2570_n3288# 0.257073f
C16 drain_right.t13 a_n2570_n3288# 0.257073f
C17 drain_right.n0 a_n2570_n3288# 2.29334f
C18 drain_right.t4 a_n2570_n3288# 0.257073f
C19 drain_right.t3 a_n2570_n3288# 0.257073f
C20 drain_right.n1 a_n2570_n3288# 2.28756f
C21 drain_right.n2 a_n2570_n3288# 0.728429f
C22 drain_right.t6 a_n2570_n3288# 0.257073f
C23 drain_right.t9 a_n2570_n3288# 0.257073f
C24 drain_right.n3 a_n2570_n3288# 2.29334f
C25 drain_right.t0 a_n2570_n3288# 0.257073f
C26 drain_right.t7 a_n2570_n3288# 0.257073f
C27 drain_right.n4 a_n2570_n3288# 2.28756f
C28 drain_right.n5 a_n2570_n3288# 0.728429f
C29 drain_right.n6 a_n2570_n3288# 1.50124f
C30 drain_right.t14 a_n2570_n3288# 0.257073f
C31 drain_right.t8 a_n2570_n3288# 0.257073f
C32 drain_right.n7 a_n2570_n3288# 2.29334f
C33 drain_right.t2 a_n2570_n3288# 0.257073f
C34 drain_right.t10 a_n2570_n3288# 0.257073f
C35 drain_right.n8 a_n2570_n3288# 2.28756f
C36 drain_right.n9 a_n2570_n3288# 0.770418f
C37 drain_right.t1 a_n2570_n3288# 0.257073f
C38 drain_right.t11 a_n2570_n3288# 0.257073f
C39 drain_right.n10 a_n2570_n3288# 2.28756f
C40 drain_right.n11 a_n2570_n3288# 0.382636f
C41 drain_right.t5 a_n2570_n3288# 0.257073f
C42 drain_right.t12 a_n2570_n3288# 0.257073f
C43 drain_right.n12 a_n2570_n3288# 2.28756f
C44 drain_right.n13 a_n2570_n3288# 0.622421f
C45 minus.n0 a_n2570_n3288# 0.040585f
C46 minus.n1 a_n2570_n3288# 0.00921f
C47 minus.t3 a_n2570_n3288# 0.972123f
C48 minus.n2 a_n2570_n3288# 0.040585f
C49 minus.n3 a_n2570_n3288# 0.00921f
C50 minus.t4 a_n2570_n3288# 0.972123f
C51 minus.n4 a_n2570_n3288# 0.040585f
C52 minus.n5 a_n2570_n3288# 0.00921f
C53 minus.t5 a_n2570_n3288# 0.972123f
C54 minus.t7 a_n2570_n3288# 0.991274f
C55 minus.t1 a_n2570_n3288# 0.972123f
C56 minus.n6 a_n2570_n3288# 0.393261f
C57 minus.n7 a_n2570_n3288# 0.371926f
C58 minus.n8 a_n2570_n3288# 0.171746f
C59 minus.n9 a_n2570_n3288# 0.040585f
C60 minus.n10 a_n2570_n3288# 0.387701f
C61 minus.n11 a_n2570_n3288# 0.00921f
C62 minus.t13 a_n2570_n3288# 0.972123f
C63 minus.n12 a_n2570_n3288# 0.387701f
C64 minus.n13 a_n2570_n3288# 0.040585f
C65 minus.n14 a_n2570_n3288# 0.040585f
C66 minus.n15 a_n2570_n3288# 0.040585f
C67 minus.n16 a_n2570_n3288# 0.387701f
C68 minus.n17 a_n2570_n3288# 0.00921f
C69 minus.t14 a_n2570_n3288# 0.972123f
C70 minus.n18 a_n2570_n3288# 0.387701f
C71 minus.n19 a_n2570_n3288# 0.040585f
C72 minus.n20 a_n2570_n3288# 0.040585f
C73 minus.n21 a_n2570_n3288# 0.040585f
C74 minus.n22 a_n2570_n3288# 0.387701f
C75 minus.n23 a_n2570_n3288# 0.00921f
C76 minus.t10 a_n2570_n3288# 0.972123f
C77 minus.n24 a_n2570_n3288# 0.386575f
C78 minus.n25 a_n2570_n3288# 1.61429f
C79 minus.n26 a_n2570_n3288# 0.040585f
C80 minus.n27 a_n2570_n3288# 0.00921f
C81 minus.n28 a_n2570_n3288# 0.040585f
C82 minus.n29 a_n2570_n3288# 0.00921f
C83 minus.n30 a_n2570_n3288# 0.040585f
C84 minus.n31 a_n2570_n3288# 0.00921f
C85 minus.t0 a_n2570_n3288# 0.991274f
C86 minus.t2 a_n2570_n3288# 0.972123f
C87 minus.n32 a_n2570_n3288# 0.393261f
C88 minus.n33 a_n2570_n3288# 0.371926f
C89 minus.n34 a_n2570_n3288# 0.171746f
C90 minus.n35 a_n2570_n3288# 0.040585f
C91 minus.t11 a_n2570_n3288# 0.972123f
C92 minus.n36 a_n2570_n3288# 0.387701f
C93 minus.n37 a_n2570_n3288# 0.00921f
C94 minus.t12 a_n2570_n3288# 0.972123f
C95 minus.n38 a_n2570_n3288# 0.387701f
C96 minus.n39 a_n2570_n3288# 0.040585f
C97 minus.n40 a_n2570_n3288# 0.040585f
C98 minus.n41 a_n2570_n3288# 0.040585f
C99 minus.t15 a_n2570_n3288# 0.972123f
C100 minus.n42 a_n2570_n3288# 0.387701f
C101 minus.n43 a_n2570_n3288# 0.00921f
C102 minus.t8 a_n2570_n3288# 0.972123f
C103 minus.n44 a_n2570_n3288# 0.387701f
C104 minus.n45 a_n2570_n3288# 0.040585f
C105 minus.n46 a_n2570_n3288# 0.040585f
C106 minus.n47 a_n2570_n3288# 0.040585f
C107 minus.t9 a_n2570_n3288# 0.972123f
C108 minus.n48 a_n2570_n3288# 0.387701f
C109 minus.n49 a_n2570_n3288# 0.00921f
C110 minus.t6 a_n2570_n3288# 0.972123f
C111 minus.n50 a_n2570_n3288# 0.386575f
C112 minus.n51 a_n2570_n3288# 0.280124f
C113 minus.n52 a_n2570_n3288# 1.94044f
C114 source.n0 a_n2570_n3288# 0.030895f
C115 source.n1 a_n2570_n3288# 0.023324f
C116 source.n2 a_n2570_n3288# 0.012533f
C117 source.n3 a_n2570_n3288# 0.029624f
C118 source.n4 a_n2570_n3288# 0.01327f
C119 source.n5 a_n2570_n3288# 0.023324f
C120 source.n6 a_n2570_n3288# 0.012533f
C121 source.n7 a_n2570_n3288# 0.029624f
C122 source.n8 a_n2570_n3288# 0.01327f
C123 source.n9 a_n2570_n3288# 0.023324f
C124 source.n10 a_n2570_n3288# 0.012902f
C125 source.n11 a_n2570_n3288# 0.029624f
C126 source.n12 a_n2570_n3288# 0.012533f
C127 source.n13 a_n2570_n3288# 0.01327f
C128 source.n14 a_n2570_n3288# 0.023324f
C129 source.n15 a_n2570_n3288# 0.012533f
C130 source.n16 a_n2570_n3288# 0.029624f
C131 source.n17 a_n2570_n3288# 0.01327f
C132 source.n18 a_n2570_n3288# 0.023324f
C133 source.n19 a_n2570_n3288# 0.012533f
C134 source.n20 a_n2570_n3288# 0.022218f
C135 source.n21 a_n2570_n3288# 0.020942f
C136 source.t23 a_n2570_n3288# 0.050033f
C137 source.n22 a_n2570_n3288# 0.168161f
C138 source.n23 a_n2570_n3288# 1.17664f
C139 source.n24 a_n2570_n3288# 0.012533f
C140 source.n25 a_n2570_n3288# 0.01327f
C141 source.n26 a_n2570_n3288# 0.029624f
C142 source.n27 a_n2570_n3288# 0.029624f
C143 source.n28 a_n2570_n3288# 0.01327f
C144 source.n29 a_n2570_n3288# 0.012533f
C145 source.n30 a_n2570_n3288# 0.023324f
C146 source.n31 a_n2570_n3288# 0.023324f
C147 source.n32 a_n2570_n3288# 0.012533f
C148 source.n33 a_n2570_n3288# 0.01327f
C149 source.n34 a_n2570_n3288# 0.029624f
C150 source.n35 a_n2570_n3288# 0.029624f
C151 source.n36 a_n2570_n3288# 0.01327f
C152 source.n37 a_n2570_n3288# 0.012533f
C153 source.n38 a_n2570_n3288# 0.023324f
C154 source.n39 a_n2570_n3288# 0.023324f
C155 source.n40 a_n2570_n3288# 0.012533f
C156 source.n41 a_n2570_n3288# 0.01327f
C157 source.n42 a_n2570_n3288# 0.029624f
C158 source.n43 a_n2570_n3288# 0.029624f
C159 source.n44 a_n2570_n3288# 0.029624f
C160 source.n45 a_n2570_n3288# 0.012902f
C161 source.n46 a_n2570_n3288# 0.012533f
C162 source.n47 a_n2570_n3288# 0.023324f
C163 source.n48 a_n2570_n3288# 0.023324f
C164 source.n49 a_n2570_n3288# 0.012533f
C165 source.n50 a_n2570_n3288# 0.01327f
C166 source.n51 a_n2570_n3288# 0.029624f
C167 source.n52 a_n2570_n3288# 0.029624f
C168 source.n53 a_n2570_n3288# 0.01327f
C169 source.n54 a_n2570_n3288# 0.012533f
C170 source.n55 a_n2570_n3288# 0.023324f
C171 source.n56 a_n2570_n3288# 0.023324f
C172 source.n57 a_n2570_n3288# 0.012533f
C173 source.n58 a_n2570_n3288# 0.01327f
C174 source.n59 a_n2570_n3288# 0.029624f
C175 source.n60 a_n2570_n3288# 0.060791f
C176 source.n61 a_n2570_n3288# 0.01327f
C177 source.n62 a_n2570_n3288# 0.012533f
C178 source.n63 a_n2570_n3288# 0.050088f
C179 source.n64 a_n2570_n3288# 0.03355f
C180 source.n65 a_n2570_n3288# 0.981142f
C181 source.t21 a_n2570_n3288# 0.221173f
C182 source.t29 a_n2570_n3288# 0.221173f
C183 source.n66 a_n2570_n3288# 1.89369f
C184 source.n67 a_n2570_n3288# 0.371918f
C185 source.t22 a_n2570_n3288# 0.221173f
C186 source.t27 a_n2570_n3288# 0.221173f
C187 source.n68 a_n2570_n3288# 1.89369f
C188 source.n69 a_n2570_n3288# 0.371918f
C189 source.t20 a_n2570_n3288# 0.221173f
C190 source.t28 a_n2570_n3288# 0.221173f
C191 source.n70 a_n2570_n3288# 1.89369f
C192 source.n71 a_n2570_n3288# 0.371918f
C193 source.n72 a_n2570_n3288# 0.030895f
C194 source.n73 a_n2570_n3288# 0.023324f
C195 source.n74 a_n2570_n3288# 0.012533f
C196 source.n75 a_n2570_n3288# 0.029624f
C197 source.n76 a_n2570_n3288# 0.01327f
C198 source.n77 a_n2570_n3288# 0.023324f
C199 source.n78 a_n2570_n3288# 0.012533f
C200 source.n79 a_n2570_n3288# 0.029624f
C201 source.n80 a_n2570_n3288# 0.01327f
C202 source.n81 a_n2570_n3288# 0.023324f
C203 source.n82 a_n2570_n3288# 0.012902f
C204 source.n83 a_n2570_n3288# 0.029624f
C205 source.n84 a_n2570_n3288# 0.012533f
C206 source.n85 a_n2570_n3288# 0.01327f
C207 source.n86 a_n2570_n3288# 0.023324f
C208 source.n87 a_n2570_n3288# 0.012533f
C209 source.n88 a_n2570_n3288# 0.029624f
C210 source.n89 a_n2570_n3288# 0.01327f
C211 source.n90 a_n2570_n3288# 0.023324f
C212 source.n91 a_n2570_n3288# 0.012533f
C213 source.n92 a_n2570_n3288# 0.022218f
C214 source.n93 a_n2570_n3288# 0.020942f
C215 source.t26 a_n2570_n3288# 0.050033f
C216 source.n94 a_n2570_n3288# 0.168161f
C217 source.n95 a_n2570_n3288# 1.17664f
C218 source.n96 a_n2570_n3288# 0.012533f
C219 source.n97 a_n2570_n3288# 0.01327f
C220 source.n98 a_n2570_n3288# 0.029624f
C221 source.n99 a_n2570_n3288# 0.029624f
C222 source.n100 a_n2570_n3288# 0.01327f
C223 source.n101 a_n2570_n3288# 0.012533f
C224 source.n102 a_n2570_n3288# 0.023324f
C225 source.n103 a_n2570_n3288# 0.023324f
C226 source.n104 a_n2570_n3288# 0.012533f
C227 source.n105 a_n2570_n3288# 0.01327f
C228 source.n106 a_n2570_n3288# 0.029624f
C229 source.n107 a_n2570_n3288# 0.029624f
C230 source.n108 a_n2570_n3288# 0.01327f
C231 source.n109 a_n2570_n3288# 0.012533f
C232 source.n110 a_n2570_n3288# 0.023324f
C233 source.n111 a_n2570_n3288# 0.023324f
C234 source.n112 a_n2570_n3288# 0.012533f
C235 source.n113 a_n2570_n3288# 0.01327f
C236 source.n114 a_n2570_n3288# 0.029624f
C237 source.n115 a_n2570_n3288# 0.029624f
C238 source.n116 a_n2570_n3288# 0.029624f
C239 source.n117 a_n2570_n3288# 0.012902f
C240 source.n118 a_n2570_n3288# 0.012533f
C241 source.n119 a_n2570_n3288# 0.023324f
C242 source.n120 a_n2570_n3288# 0.023324f
C243 source.n121 a_n2570_n3288# 0.012533f
C244 source.n122 a_n2570_n3288# 0.01327f
C245 source.n123 a_n2570_n3288# 0.029624f
C246 source.n124 a_n2570_n3288# 0.029624f
C247 source.n125 a_n2570_n3288# 0.01327f
C248 source.n126 a_n2570_n3288# 0.012533f
C249 source.n127 a_n2570_n3288# 0.023324f
C250 source.n128 a_n2570_n3288# 0.023324f
C251 source.n129 a_n2570_n3288# 0.012533f
C252 source.n130 a_n2570_n3288# 0.01327f
C253 source.n131 a_n2570_n3288# 0.029624f
C254 source.n132 a_n2570_n3288# 0.060791f
C255 source.n133 a_n2570_n3288# 0.01327f
C256 source.n134 a_n2570_n3288# 0.012533f
C257 source.n135 a_n2570_n3288# 0.050088f
C258 source.n136 a_n2570_n3288# 0.03355f
C259 source.n137 a_n2570_n3288# 0.119807f
C260 source.n138 a_n2570_n3288# 0.030895f
C261 source.n139 a_n2570_n3288# 0.023324f
C262 source.n140 a_n2570_n3288# 0.012533f
C263 source.n141 a_n2570_n3288# 0.029624f
C264 source.n142 a_n2570_n3288# 0.01327f
C265 source.n143 a_n2570_n3288# 0.023324f
C266 source.n144 a_n2570_n3288# 0.012533f
C267 source.n145 a_n2570_n3288# 0.029624f
C268 source.n146 a_n2570_n3288# 0.01327f
C269 source.n147 a_n2570_n3288# 0.023324f
C270 source.n148 a_n2570_n3288# 0.012902f
C271 source.n149 a_n2570_n3288# 0.029624f
C272 source.n150 a_n2570_n3288# 0.012533f
C273 source.n151 a_n2570_n3288# 0.01327f
C274 source.n152 a_n2570_n3288# 0.023324f
C275 source.n153 a_n2570_n3288# 0.012533f
C276 source.n154 a_n2570_n3288# 0.029624f
C277 source.n155 a_n2570_n3288# 0.01327f
C278 source.n156 a_n2570_n3288# 0.023324f
C279 source.n157 a_n2570_n3288# 0.012533f
C280 source.n158 a_n2570_n3288# 0.022218f
C281 source.n159 a_n2570_n3288# 0.020942f
C282 source.t3 a_n2570_n3288# 0.050033f
C283 source.n160 a_n2570_n3288# 0.168161f
C284 source.n161 a_n2570_n3288# 1.17664f
C285 source.n162 a_n2570_n3288# 0.012533f
C286 source.n163 a_n2570_n3288# 0.01327f
C287 source.n164 a_n2570_n3288# 0.029624f
C288 source.n165 a_n2570_n3288# 0.029624f
C289 source.n166 a_n2570_n3288# 0.01327f
C290 source.n167 a_n2570_n3288# 0.012533f
C291 source.n168 a_n2570_n3288# 0.023324f
C292 source.n169 a_n2570_n3288# 0.023324f
C293 source.n170 a_n2570_n3288# 0.012533f
C294 source.n171 a_n2570_n3288# 0.01327f
C295 source.n172 a_n2570_n3288# 0.029624f
C296 source.n173 a_n2570_n3288# 0.029624f
C297 source.n174 a_n2570_n3288# 0.01327f
C298 source.n175 a_n2570_n3288# 0.012533f
C299 source.n176 a_n2570_n3288# 0.023324f
C300 source.n177 a_n2570_n3288# 0.023324f
C301 source.n178 a_n2570_n3288# 0.012533f
C302 source.n179 a_n2570_n3288# 0.01327f
C303 source.n180 a_n2570_n3288# 0.029624f
C304 source.n181 a_n2570_n3288# 0.029624f
C305 source.n182 a_n2570_n3288# 0.029624f
C306 source.n183 a_n2570_n3288# 0.012902f
C307 source.n184 a_n2570_n3288# 0.012533f
C308 source.n185 a_n2570_n3288# 0.023324f
C309 source.n186 a_n2570_n3288# 0.023324f
C310 source.n187 a_n2570_n3288# 0.012533f
C311 source.n188 a_n2570_n3288# 0.01327f
C312 source.n189 a_n2570_n3288# 0.029624f
C313 source.n190 a_n2570_n3288# 0.029624f
C314 source.n191 a_n2570_n3288# 0.01327f
C315 source.n192 a_n2570_n3288# 0.012533f
C316 source.n193 a_n2570_n3288# 0.023324f
C317 source.n194 a_n2570_n3288# 0.023324f
C318 source.n195 a_n2570_n3288# 0.012533f
C319 source.n196 a_n2570_n3288# 0.01327f
C320 source.n197 a_n2570_n3288# 0.029624f
C321 source.n198 a_n2570_n3288# 0.060791f
C322 source.n199 a_n2570_n3288# 0.01327f
C323 source.n200 a_n2570_n3288# 0.012533f
C324 source.n201 a_n2570_n3288# 0.050088f
C325 source.n202 a_n2570_n3288# 0.03355f
C326 source.n203 a_n2570_n3288# 0.119807f
C327 source.t2 a_n2570_n3288# 0.221173f
C328 source.t8 a_n2570_n3288# 0.221173f
C329 source.n204 a_n2570_n3288# 1.89369f
C330 source.n205 a_n2570_n3288# 0.371918f
C331 source.t15 a_n2570_n3288# 0.221173f
C332 source.t12 a_n2570_n3288# 0.221173f
C333 source.n206 a_n2570_n3288# 1.89369f
C334 source.n207 a_n2570_n3288# 0.371918f
C335 source.t6 a_n2570_n3288# 0.221173f
C336 source.t14 a_n2570_n3288# 0.221173f
C337 source.n208 a_n2570_n3288# 1.89369f
C338 source.n209 a_n2570_n3288# 0.371918f
C339 source.n210 a_n2570_n3288# 0.030895f
C340 source.n211 a_n2570_n3288# 0.023324f
C341 source.n212 a_n2570_n3288# 0.012533f
C342 source.n213 a_n2570_n3288# 0.029624f
C343 source.n214 a_n2570_n3288# 0.01327f
C344 source.n215 a_n2570_n3288# 0.023324f
C345 source.n216 a_n2570_n3288# 0.012533f
C346 source.n217 a_n2570_n3288# 0.029624f
C347 source.n218 a_n2570_n3288# 0.01327f
C348 source.n219 a_n2570_n3288# 0.023324f
C349 source.n220 a_n2570_n3288# 0.012902f
C350 source.n221 a_n2570_n3288# 0.029624f
C351 source.n222 a_n2570_n3288# 0.012533f
C352 source.n223 a_n2570_n3288# 0.01327f
C353 source.n224 a_n2570_n3288# 0.023324f
C354 source.n225 a_n2570_n3288# 0.012533f
C355 source.n226 a_n2570_n3288# 0.029624f
C356 source.n227 a_n2570_n3288# 0.01327f
C357 source.n228 a_n2570_n3288# 0.023324f
C358 source.n229 a_n2570_n3288# 0.012533f
C359 source.n230 a_n2570_n3288# 0.022218f
C360 source.n231 a_n2570_n3288# 0.020942f
C361 source.t11 a_n2570_n3288# 0.050033f
C362 source.n232 a_n2570_n3288# 0.168161f
C363 source.n233 a_n2570_n3288# 1.17664f
C364 source.n234 a_n2570_n3288# 0.012533f
C365 source.n235 a_n2570_n3288# 0.01327f
C366 source.n236 a_n2570_n3288# 0.029624f
C367 source.n237 a_n2570_n3288# 0.029624f
C368 source.n238 a_n2570_n3288# 0.01327f
C369 source.n239 a_n2570_n3288# 0.012533f
C370 source.n240 a_n2570_n3288# 0.023324f
C371 source.n241 a_n2570_n3288# 0.023324f
C372 source.n242 a_n2570_n3288# 0.012533f
C373 source.n243 a_n2570_n3288# 0.01327f
C374 source.n244 a_n2570_n3288# 0.029624f
C375 source.n245 a_n2570_n3288# 0.029624f
C376 source.n246 a_n2570_n3288# 0.01327f
C377 source.n247 a_n2570_n3288# 0.012533f
C378 source.n248 a_n2570_n3288# 0.023324f
C379 source.n249 a_n2570_n3288# 0.023324f
C380 source.n250 a_n2570_n3288# 0.012533f
C381 source.n251 a_n2570_n3288# 0.01327f
C382 source.n252 a_n2570_n3288# 0.029624f
C383 source.n253 a_n2570_n3288# 0.029624f
C384 source.n254 a_n2570_n3288# 0.029624f
C385 source.n255 a_n2570_n3288# 0.012902f
C386 source.n256 a_n2570_n3288# 0.012533f
C387 source.n257 a_n2570_n3288# 0.023324f
C388 source.n258 a_n2570_n3288# 0.023324f
C389 source.n259 a_n2570_n3288# 0.012533f
C390 source.n260 a_n2570_n3288# 0.01327f
C391 source.n261 a_n2570_n3288# 0.029624f
C392 source.n262 a_n2570_n3288# 0.029624f
C393 source.n263 a_n2570_n3288# 0.01327f
C394 source.n264 a_n2570_n3288# 0.012533f
C395 source.n265 a_n2570_n3288# 0.023324f
C396 source.n266 a_n2570_n3288# 0.023324f
C397 source.n267 a_n2570_n3288# 0.012533f
C398 source.n268 a_n2570_n3288# 0.01327f
C399 source.n269 a_n2570_n3288# 0.029624f
C400 source.n270 a_n2570_n3288# 0.060791f
C401 source.n271 a_n2570_n3288# 0.01327f
C402 source.n272 a_n2570_n3288# 0.012533f
C403 source.n273 a_n2570_n3288# 0.050088f
C404 source.n274 a_n2570_n3288# 0.03355f
C405 source.n275 a_n2570_n3288# 1.35724f
C406 source.n276 a_n2570_n3288# 0.030895f
C407 source.n277 a_n2570_n3288# 0.023324f
C408 source.n278 a_n2570_n3288# 0.012533f
C409 source.n279 a_n2570_n3288# 0.029624f
C410 source.n280 a_n2570_n3288# 0.01327f
C411 source.n281 a_n2570_n3288# 0.023324f
C412 source.n282 a_n2570_n3288# 0.012533f
C413 source.n283 a_n2570_n3288# 0.029624f
C414 source.n284 a_n2570_n3288# 0.01327f
C415 source.n285 a_n2570_n3288# 0.023324f
C416 source.n286 a_n2570_n3288# 0.012902f
C417 source.n287 a_n2570_n3288# 0.029624f
C418 source.n288 a_n2570_n3288# 0.01327f
C419 source.n289 a_n2570_n3288# 0.023324f
C420 source.n290 a_n2570_n3288# 0.012533f
C421 source.n291 a_n2570_n3288# 0.029624f
C422 source.n292 a_n2570_n3288# 0.01327f
C423 source.n293 a_n2570_n3288# 0.023324f
C424 source.n294 a_n2570_n3288# 0.012533f
C425 source.n295 a_n2570_n3288# 0.022218f
C426 source.n296 a_n2570_n3288# 0.020942f
C427 source.t18 a_n2570_n3288# 0.050033f
C428 source.n297 a_n2570_n3288# 0.168161f
C429 source.n298 a_n2570_n3288# 1.17664f
C430 source.n299 a_n2570_n3288# 0.012533f
C431 source.n300 a_n2570_n3288# 0.01327f
C432 source.n301 a_n2570_n3288# 0.029624f
C433 source.n302 a_n2570_n3288# 0.029624f
C434 source.n303 a_n2570_n3288# 0.01327f
C435 source.n304 a_n2570_n3288# 0.012533f
C436 source.n305 a_n2570_n3288# 0.023324f
C437 source.n306 a_n2570_n3288# 0.023324f
C438 source.n307 a_n2570_n3288# 0.012533f
C439 source.n308 a_n2570_n3288# 0.01327f
C440 source.n309 a_n2570_n3288# 0.029624f
C441 source.n310 a_n2570_n3288# 0.029624f
C442 source.n311 a_n2570_n3288# 0.01327f
C443 source.n312 a_n2570_n3288# 0.012533f
C444 source.n313 a_n2570_n3288# 0.023324f
C445 source.n314 a_n2570_n3288# 0.023324f
C446 source.n315 a_n2570_n3288# 0.012533f
C447 source.n316 a_n2570_n3288# 0.012533f
C448 source.n317 a_n2570_n3288# 0.01327f
C449 source.n318 a_n2570_n3288# 0.029624f
C450 source.n319 a_n2570_n3288# 0.029624f
C451 source.n320 a_n2570_n3288# 0.029624f
C452 source.n321 a_n2570_n3288# 0.012902f
C453 source.n322 a_n2570_n3288# 0.012533f
C454 source.n323 a_n2570_n3288# 0.023324f
C455 source.n324 a_n2570_n3288# 0.023324f
C456 source.n325 a_n2570_n3288# 0.012533f
C457 source.n326 a_n2570_n3288# 0.01327f
C458 source.n327 a_n2570_n3288# 0.029624f
C459 source.n328 a_n2570_n3288# 0.029624f
C460 source.n329 a_n2570_n3288# 0.01327f
C461 source.n330 a_n2570_n3288# 0.012533f
C462 source.n331 a_n2570_n3288# 0.023324f
C463 source.n332 a_n2570_n3288# 0.023324f
C464 source.n333 a_n2570_n3288# 0.012533f
C465 source.n334 a_n2570_n3288# 0.01327f
C466 source.n335 a_n2570_n3288# 0.029624f
C467 source.n336 a_n2570_n3288# 0.060791f
C468 source.n337 a_n2570_n3288# 0.01327f
C469 source.n338 a_n2570_n3288# 0.012533f
C470 source.n339 a_n2570_n3288# 0.050088f
C471 source.n340 a_n2570_n3288# 0.03355f
C472 source.n341 a_n2570_n3288# 1.35724f
C473 source.t30 a_n2570_n3288# 0.221173f
C474 source.t31 a_n2570_n3288# 0.221173f
C475 source.n342 a_n2570_n3288# 1.89367f
C476 source.n343 a_n2570_n3288# 0.37193f
C477 source.t24 a_n2570_n3288# 0.221173f
C478 source.t25 a_n2570_n3288# 0.221173f
C479 source.n344 a_n2570_n3288# 1.89367f
C480 source.n345 a_n2570_n3288# 0.37193f
C481 source.t19 a_n2570_n3288# 0.221173f
C482 source.t16 a_n2570_n3288# 0.221173f
C483 source.n346 a_n2570_n3288# 1.89367f
C484 source.n347 a_n2570_n3288# 0.37193f
C485 source.n348 a_n2570_n3288# 0.030895f
C486 source.n349 a_n2570_n3288# 0.023324f
C487 source.n350 a_n2570_n3288# 0.012533f
C488 source.n351 a_n2570_n3288# 0.029624f
C489 source.n352 a_n2570_n3288# 0.01327f
C490 source.n353 a_n2570_n3288# 0.023324f
C491 source.n354 a_n2570_n3288# 0.012533f
C492 source.n355 a_n2570_n3288# 0.029624f
C493 source.n356 a_n2570_n3288# 0.01327f
C494 source.n357 a_n2570_n3288# 0.023324f
C495 source.n358 a_n2570_n3288# 0.012902f
C496 source.n359 a_n2570_n3288# 0.029624f
C497 source.n360 a_n2570_n3288# 0.01327f
C498 source.n361 a_n2570_n3288# 0.023324f
C499 source.n362 a_n2570_n3288# 0.012533f
C500 source.n363 a_n2570_n3288# 0.029624f
C501 source.n364 a_n2570_n3288# 0.01327f
C502 source.n365 a_n2570_n3288# 0.023324f
C503 source.n366 a_n2570_n3288# 0.012533f
C504 source.n367 a_n2570_n3288# 0.022218f
C505 source.n368 a_n2570_n3288# 0.020942f
C506 source.t17 a_n2570_n3288# 0.050033f
C507 source.n369 a_n2570_n3288# 0.168161f
C508 source.n370 a_n2570_n3288# 1.17664f
C509 source.n371 a_n2570_n3288# 0.012533f
C510 source.n372 a_n2570_n3288# 0.01327f
C511 source.n373 a_n2570_n3288# 0.029624f
C512 source.n374 a_n2570_n3288# 0.029624f
C513 source.n375 a_n2570_n3288# 0.01327f
C514 source.n376 a_n2570_n3288# 0.012533f
C515 source.n377 a_n2570_n3288# 0.023324f
C516 source.n378 a_n2570_n3288# 0.023324f
C517 source.n379 a_n2570_n3288# 0.012533f
C518 source.n380 a_n2570_n3288# 0.01327f
C519 source.n381 a_n2570_n3288# 0.029624f
C520 source.n382 a_n2570_n3288# 0.029624f
C521 source.n383 a_n2570_n3288# 0.01327f
C522 source.n384 a_n2570_n3288# 0.012533f
C523 source.n385 a_n2570_n3288# 0.023324f
C524 source.n386 a_n2570_n3288# 0.023324f
C525 source.n387 a_n2570_n3288# 0.012533f
C526 source.n388 a_n2570_n3288# 0.012533f
C527 source.n389 a_n2570_n3288# 0.01327f
C528 source.n390 a_n2570_n3288# 0.029624f
C529 source.n391 a_n2570_n3288# 0.029624f
C530 source.n392 a_n2570_n3288# 0.029624f
C531 source.n393 a_n2570_n3288# 0.012902f
C532 source.n394 a_n2570_n3288# 0.012533f
C533 source.n395 a_n2570_n3288# 0.023324f
C534 source.n396 a_n2570_n3288# 0.023324f
C535 source.n397 a_n2570_n3288# 0.012533f
C536 source.n398 a_n2570_n3288# 0.01327f
C537 source.n399 a_n2570_n3288# 0.029624f
C538 source.n400 a_n2570_n3288# 0.029624f
C539 source.n401 a_n2570_n3288# 0.01327f
C540 source.n402 a_n2570_n3288# 0.012533f
C541 source.n403 a_n2570_n3288# 0.023324f
C542 source.n404 a_n2570_n3288# 0.023324f
C543 source.n405 a_n2570_n3288# 0.012533f
C544 source.n406 a_n2570_n3288# 0.01327f
C545 source.n407 a_n2570_n3288# 0.029624f
C546 source.n408 a_n2570_n3288# 0.060791f
C547 source.n409 a_n2570_n3288# 0.01327f
C548 source.n410 a_n2570_n3288# 0.012533f
C549 source.n411 a_n2570_n3288# 0.050088f
C550 source.n412 a_n2570_n3288# 0.03355f
C551 source.n413 a_n2570_n3288# 0.119807f
C552 source.n414 a_n2570_n3288# 0.030895f
C553 source.n415 a_n2570_n3288# 0.023324f
C554 source.n416 a_n2570_n3288# 0.012533f
C555 source.n417 a_n2570_n3288# 0.029624f
C556 source.n418 a_n2570_n3288# 0.01327f
C557 source.n419 a_n2570_n3288# 0.023324f
C558 source.n420 a_n2570_n3288# 0.012533f
C559 source.n421 a_n2570_n3288# 0.029624f
C560 source.n422 a_n2570_n3288# 0.01327f
C561 source.n423 a_n2570_n3288# 0.023324f
C562 source.n424 a_n2570_n3288# 0.012902f
C563 source.n425 a_n2570_n3288# 0.029624f
C564 source.n426 a_n2570_n3288# 0.01327f
C565 source.n427 a_n2570_n3288# 0.023324f
C566 source.n428 a_n2570_n3288# 0.012533f
C567 source.n429 a_n2570_n3288# 0.029624f
C568 source.n430 a_n2570_n3288# 0.01327f
C569 source.n431 a_n2570_n3288# 0.023324f
C570 source.n432 a_n2570_n3288# 0.012533f
C571 source.n433 a_n2570_n3288# 0.022218f
C572 source.n434 a_n2570_n3288# 0.020942f
C573 source.t7 a_n2570_n3288# 0.050033f
C574 source.n435 a_n2570_n3288# 0.168161f
C575 source.n436 a_n2570_n3288# 1.17664f
C576 source.n437 a_n2570_n3288# 0.012533f
C577 source.n438 a_n2570_n3288# 0.01327f
C578 source.n439 a_n2570_n3288# 0.029624f
C579 source.n440 a_n2570_n3288# 0.029624f
C580 source.n441 a_n2570_n3288# 0.01327f
C581 source.n442 a_n2570_n3288# 0.012533f
C582 source.n443 a_n2570_n3288# 0.023324f
C583 source.n444 a_n2570_n3288# 0.023324f
C584 source.n445 a_n2570_n3288# 0.012533f
C585 source.n446 a_n2570_n3288# 0.01327f
C586 source.n447 a_n2570_n3288# 0.029624f
C587 source.n448 a_n2570_n3288# 0.029624f
C588 source.n449 a_n2570_n3288# 0.01327f
C589 source.n450 a_n2570_n3288# 0.012533f
C590 source.n451 a_n2570_n3288# 0.023324f
C591 source.n452 a_n2570_n3288# 0.023324f
C592 source.n453 a_n2570_n3288# 0.012533f
C593 source.n454 a_n2570_n3288# 0.012533f
C594 source.n455 a_n2570_n3288# 0.01327f
C595 source.n456 a_n2570_n3288# 0.029624f
C596 source.n457 a_n2570_n3288# 0.029624f
C597 source.n458 a_n2570_n3288# 0.029624f
C598 source.n459 a_n2570_n3288# 0.012902f
C599 source.n460 a_n2570_n3288# 0.012533f
C600 source.n461 a_n2570_n3288# 0.023324f
C601 source.n462 a_n2570_n3288# 0.023324f
C602 source.n463 a_n2570_n3288# 0.012533f
C603 source.n464 a_n2570_n3288# 0.01327f
C604 source.n465 a_n2570_n3288# 0.029624f
C605 source.n466 a_n2570_n3288# 0.029624f
C606 source.n467 a_n2570_n3288# 0.01327f
C607 source.n468 a_n2570_n3288# 0.012533f
C608 source.n469 a_n2570_n3288# 0.023324f
C609 source.n470 a_n2570_n3288# 0.023324f
C610 source.n471 a_n2570_n3288# 0.012533f
C611 source.n472 a_n2570_n3288# 0.01327f
C612 source.n473 a_n2570_n3288# 0.029624f
C613 source.n474 a_n2570_n3288# 0.060791f
C614 source.n475 a_n2570_n3288# 0.01327f
C615 source.n476 a_n2570_n3288# 0.012533f
C616 source.n477 a_n2570_n3288# 0.050088f
C617 source.n478 a_n2570_n3288# 0.03355f
C618 source.n479 a_n2570_n3288# 0.119807f
C619 source.t10 a_n2570_n3288# 0.221173f
C620 source.t0 a_n2570_n3288# 0.221173f
C621 source.n480 a_n2570_n3288# 1.89367f
C622 source.n481 a_n2570_n3288# 0.37193f
C623 source.t13 a_n2570_n3288# 0.221173f
C624 source.t5 a_n2570_n3288# 0.221173f
C625 source.n482 a_n2570_n3288# 1.89367f
C626 source.n483 a_n2570_n3288# 0.37193f
C627 source.t4 a_n2570_n3288# 0.221173f
C628 source.t9 a_n2570_n3288# 0.221173f
C629 source.n484 a_n2570_n3288# 1.89367f
C630 source.n485 a_n2570_n3288# 0.37193f
C631 source.n486 a_n2570_n3288# 0.030895f
C632 source.n487 a_n2570_n3288# 0.023324f
C633 source.n488 a_n2570_n3288# 0.012533f
C634 source.n489 a_n2570_n3288# 0.029624f
C635 source.n490 a_n2570_n3288# 0.01327f
C636 source.n491 a_n2570_n3288# 0.023324f
C637 source.n492 a_n2570_n3288# 0.012533f
C638 source.n493 a_n2570_n3288# 0.029624f
C639 source.n494 a_n2570_n3288# 0.01327f
C640 source.n495 a_n2570_n3288# 0.023324f
C641 source.n496 a_n2570_n3288# 0.012902f
C642 source.n497 a_n2570_n3288# 0.029624f
C643 source.n498 a_n2570_n3288# 0.01327f
C644 source.n499 a_n2570_n3288# 0.023324f
C645 source.n500 a_n2570_n3288# 0.012533f
C646 source.n501 a_n2570_n3288# 0.029624f
C647 source.n502 a_n2570_n3288# 0.01327f
C648 source.n503 a_n2570_n3288# 0.023324f
C649 source.n504 a_n2570_n3288# 0.012533f
C650 source.n505 a_n2570_n3288# 0.022218f
C651 source.n506 a_n2570_n3288# 0.020942f
C652 source.t1 a_n2570_n3288# 0.050033f
C653 source.n507 a_n2570_n3288# 0.168161f
C654 source.n508 a_n2570_n3288# 1.17664f
C655 source.n509 a_n2570_n3288# 0.012533f
C656 source.n510 a_n2570_n3288# 0.01327f
C657 source.n511 a_n2570_n3288# 0.029624f
C658 source.n512 a_n2570_n3288# 0.029624f
C659 source.n513 a_n2570_n3288# 0.01327f
C660 source.n514 a_n2570_n3288# 0.012533f
C661 source.n515 a_n2570_n3288# 0.023324f
C662 source.n516 a_n2570_n3288# 0.023324f
C663 source.n517 a_n2570_n3288# 0.012533f
C664 source.n518 a_n2570_n3288# 0.01327f
C665 source.n519 a_n2570_n3288# 0.029624f
C666 source.n520 a_n2570_n3288# 0.029624f
C667 source.n521 a_n2570_n3288# 0.01327f
C668 source.n522 a_n2570_n3288# 0.012533f
C669 source.n523 a_n2570_n3288# 0.023324f
C670 source.n524 a_n2570_n3288# 0.023324f
C671 source.n525 a_n2570_n3288# 0.012533f
C672 source.n526 a_n2570_n3288# 0.012533f
C673 source.n527 a_n2570_n3288# 0.01327f
C674 source.n528 a_n2570_n3288# 0.029624f
C675 source.n529 a_n2570_n3288# 0.029624f
C676 source.n530 a_n2570_n3288# 0.029624f
C677 source.n531 a_n2570_n3288# 0.012902f
C678 source.n532 a_n2570_n3288# 0.012533f
C679 source.n533 a_n2570_n3288# 0.023324f
C680 source.n534 a_n2570_n3288# 0.023324f
C681 source.n535 a_n2570_n3288# 0.012533f
C682 source.n536 a_n2570_n3288# 0.01327f
C683 source.n537 a_n2570_n3288# 0.029624f
C684 source.n538 a_n2570_n3288# 0.029624f
C685 source.n539 a_n2570_n3288# 0.01327f
C686 source.n540 a_n2570_n3288# 0.012533f
C687 source.n541 a_n2570_n3288# 0.023324f
C688 source.n542 a_n2570_n3288# 0.023324f
C689 source.n543 a_n2570_n3288# 0.012533f
C690 source.n544 a_n2570_n3288# 0.01327f
C691 source.n545 a_n2570_n3288# 0.029624f
C692 source.n546 a_n2570_n3288# 0.060791f
C693 source.n547 a_n2570_n3288# 0.01327f
C694 source.n548 a_n2570_n3288# 0.012533f
C695 source.n549 a_n2570_n3288# 0.050088f
C696 source.n550 a_n2570_n3288# 0.03355f
C697 source.n551 a_n2570_n3288# 0.271949f
C698 source.n552 a_n2570_n3288# 1.47797f
C699 drain_left.t12 a_n2570_n3288# 0.258729f
C700 drain_left.t5 a_n2570_n3288# 0.258729f
C701 drain_left.n0 a_n2570_n3288# 2.30811f
C702 drain_left.t6 a_n2570_n3288# 0.258729f
C703 drain_left.t11 a_n2570_n3288# 0.258729f
C704 drain_left.n1 a_n2570_n3288# 2.30229f
C705 drain_left.n2 a_n2570_n3288# 0.733121f
C706 drain_left.t8 a_n2570_n3288# 0.258729f
C707 drain_left.t13 a_n2570_n3288# 0.258729f
C708 drain_left.n3 a_n2570_n3288# 2.30811f
C709 drain_left.t2 a_n2570_n3288# 0.258729f
C710 drain_left.t14 a_n2570_n3288# 0.258729f
C711 drain_left.n4 a_n2570_n3288# 2.30229f
C712 drain_left.n5 a_n2570_n3288# 0.733121f
C713 drain_left.n6 a_n2570_n3288# 1.56684f
C714 drain_left.t10 a_n2570_n3288# 0.258729f
C715 drain_left.t3 a_n2570_n3288# 0.258729f
C716 drain_left.n7 a_n2570_n3288# 2.30812f
C717 drain_left.t9 a_n2570_n3288# 0.258729f
C718 drain_left.t7 a_n2570_n3288# 0.258729f
C719 drain_left.n8 a_n2570_n3288# 2.3023f
C720 drain_left.n9 a_n2570_n3288# 0.775372f
C721 drain_left.t1 a_n2570_n3288# 0.258729f
C722 drain_left.t15 a_n2570_n3288# 0.258729f
C723 drain_left.n10 a_n2570_n3288# 2.3023f
C724 drain_left.n11 a_n2570_n3288# 0.385101f
C725 drain_left.t0 a_n2570_n3288# 0.258729f
C726 drain_left.t4 a_n2570_n3288# 0.258729f
C727 drain_left.n12 a_n2570_n3288# 2.30229f
C728 drain_left.n13 a_n2570_n3288# 0.62644f
C729 plus.n0 a_n2570_n3288# 0.041163f
C730 plus.t8 a_n2570_n3288# 0.985972f
C731 plus.t2 a_n2570_n3288# 0.985972f
C732 plus.n1 a_n2570_n3288# 0.041163f
C733 plus.t10 a_n2570_n3288# 0.985972f
C734 plus.n2 a_n2570_n3288# 0.393224f
C735 plus.n3 a_n2570_n3288# 0.041163f
C736 plus.t4 a_n2570_n3288# 0.985972f
C737 plus.t9 a_n2570_n3288# 0.985972f
C738 plus.n4 a_n2570_n3288# 0.393224f
C739 plus.n5 a_n2570_n3288# 0.041163f
C740 plus.t3 a_n2570_n3288# 0.985972f
C741 plus.t11 a_n2570_n3288# 0.985972f
C742 plus.n6 a_n2570_n3288# 0.398863f
C743 plus.t5 a_n2570_n3288# 1.0054f
C744 plus.n7 a_n2570_n3288# 0.377225f
C745 plus.n8 a_n2570_n3288# 0.174193f
C746 plus.n9 a_n2570_n3288# 0.009341f
C747 plus.n10 a_n2570_n3288# 0.393224f
C748 plus.n11 a_n2570_n3288# 0.009341f
C749 plus.n12 a_n2570_n3288# 0.041163f
C750 plus.n13 a_n2570_n3288# 0.041163f
C751 plus.n14 a_n2570_n3288# 0.041163f
C752 plus.n15 a_n2570_n3288# 0.009341f
C753 plus.n16 a_n2570_n3288# 0.393224f
C754 plus.n17 a_n2570_n3288# 0.009341f
C755 plus.n18 a_n2570_n3288# 0.041163f
C756 plus.n19 a_n2570_n3288# 0.041163f
C757 plus.n20 a_n2570_n3288# 0.041163f
C758 plus.n21 a_n2570_n3288# 0.009341f
C759 plus.n22 a_n2570_n3288# 0.393224f
C760 plus.n23 a_n2570_n3288# 0.009341f
C761 plus.n24 a_n2570_n3288# 0.392082f
C762 plus.n25 a_n2570_n3288# 0.475827f
C763 plus.n26 a_n2570_n3288# 0.041163f
C764 plus.t13 a_n2570_n3288# 0.985972f
C765 plus.n27 a_n2570_n3288# 0.041163f
C766 plus.t1 a_n2570_n3288# 0.985972f
C767 plus.t0 a_n2570_n3288# 0.985972f
C768 plus.n28 a_n2570_n3288# 0.393224f
C769 plus.n29 a_n2570_n3288# 0.041163f
C770 plus.t7 a_n2570_n3288# 0.985972f
C771 plus.t6 a_n2570_n3288# 0.985972f
C772 plus.n30 a_n2570_n3288# 0.393224f
C773 plus.n31 a_n2570_n3288# 0.041163f
C774 plus.t12 a_n2570_n3288# 0.985972f
C775 plus.t15 a_n2570_n3288# 0.985972f
C776 plus.n32 a_n2570_n3288# 0.398863f
C777 plus.t14 a_n2570_n3288# 1.0054f
C778 plus.n33 a_n2570_n3288# 0.377225f
C779 plus.n34 a_n2570_n3288# 0.174193f
C780 plus.n35 a_n2570_n3288# 0.009341f
C781 plus.n36 a_n2570_n3288# 0.393224f
C782 plus.n37 a_n2570_n3288# 0.009341f
C783 plus.n38 a_n2570_n3288# 0.041163f
C784 plus.n39 a_n2570_n3288# 0.041163f
C785 plus.n40 a_n2570_n3288# 0.041163f
C786 plus.n41 a_n2570_n3288# 0.009341f
C787 plus.n42 a_n2570_n3288# 0.393224f
C788 plus.n43 a_n2570_n3288# 0.009341f
C789 plus.n44 a_n2570_n3288# 0.041163f
C790 plus.n45 a_n2570_n3288# 0.041163f
C791 plus.n46 a_n2570_n3288# 0.041163f
C792 plus.n47 a_n2570_n3288# 0.009341f
C793 plus.n48 a_n2570_n3288# 0.393224f
C794 plus.n49 a_n2570_n3288# 0.009341f
C795 plus.n50 a_n2570_n3288# 0.392082f
C796 plus.n51 a_n2570_n3288# 1.39579f
.ends

