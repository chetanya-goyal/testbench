* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t8 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 drain_right.t4 minus.t1 source.t6 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X2 a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X3 drain_left.t5 plus.t0 source.t2 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X4 a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X5 drain_left.t4 plus.t1 source.t1 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X6 a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X7 source.t5 plus.t2 drain_left.t3 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X8 drain_right.t3 minus.t2 source.t9 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X9 source.t4 plus.t3 drain_left.t2 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X10 a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X11 drain_right.t2 minus.t3 source.t7 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X12 source.t11 minus.t4 drain_right.t1 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X13 drain_left.t1 plus.t4 source.t0 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X14 source.t10 minus.t5 drain_right.t0 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 drain_left.t0 plus.t5 source.t3 a_n1220_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
R0 minus.n2 minus.t1 320.603
R1 minus.n0 minus.t3 320.603
R2 minus.n6 minus.t2 320.603
R3 minus.n4 minus.t0 320.603
R4 minus.n1 minus.t5 265.101
R5 minus.n5 minus.t4 265.101
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 26.1994
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 source.n34 source.n32 289.615
R18 source.n24 source.n22 289.615
R19 source.n2 source.n0 289.615
R20 source.n12 source.n10 289.615
R21 source.n35 source.n34 185
R22 source.n25 source.n24 185
R23 source.n3 source.n2 185
R24 source.n13 source.n12 185
R25 source.t9 source.n33 167.117
R26 source.t3 source.n23 167.117
R27 source.t0 source.n1 167.117
R28 source.t7 source.n11 167.117
R29 source.n9 source.n8 84.1169
R30 source.n19 source.n18 84.1169
R31 source.n31 source.n30 84.1168
R32 source.n21 source.n20 84.1168
R33 source.n34 source.t9 52.3082
R34 source.n24 source.t3 52.3082
R35 source.n2 source.t0 52.3082
R36 source.n12 source.t7 52.3082
R37 source.n39 source.n38 31.4096
R38 source.n29 source.n28 31.4096
R39 source.n7 source.n6 31.4096
R40 source.n17 source.n16 31.4096
R41 source.n21 source.n19 14.7982
R42 source.n30 source.t8 9.9005
R43 source.n30 source.t11 9.9005
R44 source.n20 source.t1 9.9005
R45 source.n20 source.t4 9.9005
R46 source.n8 source.t2 9.9005
R47 source.n8 source.t5 9.9005
R48 source.n18 source.t6 9.9005
R49 source.n18 source.t10 9.9005
R50 source.n35 source.n33 9.71174
R51 source.n25 source.n23 9.71174
R52 source.n3 source.n1 9.71174
R53 source.n13 source.n11 9.71174
R54 source.n38 source.n37 9.45567
R55 source.n28 source.n27 9.45567
R56 source.n6 source.n5 9.45567
R57 source.n16 source.n15 9.45567
R58 source.n37 source.n36 9.3005
R59 source.n27 source.n26 9.3005
R60 source.n5 source.n4 9.3005
R61 source.n15 source.n14 9.3005
R62 source.n40 source.n7 8.72059
R63 source.n38 source.n32 8.14595
R64 source.n28 source.n22 8.14595
R65 source.n6 source.n0 8.14595
R66 source.n16 source.n10 8.14595
R67 source.n36 source.n35 7.3702
R68 source.n26 source.n25 7.3702
R69 source.n4 source.n3 7.3702
R70 source.n14 source.n13 7.3702
R71 source.n36 source.n32 5.81868
R72 source.n26 source.n22 5.81868
R73 source.n4 source.n0 5.81868
R74 source.n14 source.n10 5.81868
R75 source.n40 source.n39 5.53498
R76 source.n37 source.n33 3.44771
R77 source.n27 source.n23 3.44771
R78 source.n5 source.n1 3.44771
R79 source.n15 source.n11 3.44771
R80 source.n17 source.n9 0.741879
R81 source.n31 source.n29 0.741879
R82 source.n19 source.n17 0.543603
R83 source.n9 source.n7 0.543603
R84 source.n29 source.n21 0.543603
R85 source.n39 source.n31 0.543603
R86 source source.n40 0.188
R87 drain_right.n2 drain_right.n0 289.615
R88 drain_right.n12 drain_right.n10 289.615
R89 drain_right.n3 drain_right.n2 185
R90 drain_right.n13 drain_right.n12 185
R91 drain_right.t5 drain_right.n1 167.117
R92 drain_right.t4 drain_right.n11 167.117
R93 drain_right.n17 drain_right.n9 101.338
R94 drain_right.n8 drain_right.n7 100.876
R95 drain_right.n2 drain_right.t5 52.3082
R96 drain_right.n12 drain_right.t4 52.3082
R97 drain_right.n8 drain_right.n6 48.4404
R98 drain_right.n17 drain_right.n16 48.0884
R99 drain_right drain_right.n8 20.7316
R100 drain_right.n7 drain_right.t1 9.9005
R101 drain_right.n7 drain_right.t3 9.9005
R102 drain_right.n9 drain_right.t0 9.9005
R103 drain_right.n9 drain_right.t2 9.9005
R104 drain_right.n3 drain_right.n1 9.71174
R105 drain_right.n13 drain_right.n11 9.71174
R106 drain_right.n6 drain_right.n5 9.45567
R107 drain_right.n16 drain_right.n15 9.45567
R108 drain_right.n5 drain_right.n4 9.3005
R109 drain_right.n15 drain_right.n14 9.3005
R110 drain_right.n6 drain_right.n0 8.14595
R111 drain_right.n16 drain_right.n10 8.14595
R112 drain_right.n4 drain_right.n3 7.3702
R113 drain_right.n14 drain_right.n13 7.3702
R114 drain_right drain_right.n17 5.92477
R115 drain_right.n4 drain_right.n0 5.81868
R116 drain_right.n14 drain_right.n10 5.81868
R117 drain_right.n5 drain_right.n1 3.44771
R118 drain_right.n15 drain_right.n11 3.44771
R119 plus.n0 plus.t0 320.603
R120 plus.n2 plus.t4 320.603
R121 plus.n4 plus.t5 320.603
R122 plus.n6 plus.t1 320.603
R123 plus.n1 plus.t2 265.101
R124 plus.n5 plus.t3 265.101
R125 plus.n3 plus.n0 161.489
R126 plus.n7 plus.n4 161.489
R127 plus.n3 plus.n2 161.3
R128 plus.n7 plus.n6 161.3
R129 plus.n1 plus.n0 36.5157
R130 plus.n2 plus.n1 36.5157
R131 plus.n6 plus.n5 36.5157
R132 plus.n5 plus.n4 36.5157
R133 plus plus.n7 23.8683
R134 plus plus.n3 8.38876
R135 drain_left.n2 drain_left.n0 289.615
R136 drain_left.n11 drain_left.n9 289.615
R137 drain_left.n3 drain_left.n2 185
R138 drain_left.n12 drain_left.n11 185
R139 drain_left.t4 drain_left.n1 167.117
R140 drain_left.t5 drain_left.n10 167.117
R141 drain_left.n8 drain_left.n7 100.876
R142 drain_left.n17 drain_left.n16 100.796
R143 drain_left.n2 drain_left.t4 52.3082
R144 drain_left.n11 drain_left.t5 52.3082
R145 drain_left.n17 drain_left.n15 48.6315
R146 drain_left.n8 drain_left.n6 48.4404
R147 drain_left drain_left.n8 21.2849
R148 drain_left.n7 drain_left.t2 9.9005
R149 drain_left.n7 drain_left.t0 9.9005
R150 drain_left.n16 drain_left.t3 9.9005
R151 drain_left.n16 drain_left.t1 9.9005
R152 drain_left.n3 drain_left.n1 9.71174
R153 drain_left.n12 drain_left.n10 9.71174
R154 drain_left.n6 drain_left.n5 9.45567
R155 drain_left.n15 drain_left.n14 9.45567
R156 drain_left.n5 drain_left.n4 9.3005
R157 drain_left.n14 drain_left.n13 9.3005
R158 drain_left.n6 drain_left.n0 8.14595
R159 drain_left.n15 drain_left.n9 8.14595
R160 drain_left.n4 drain_left.n3 7.3702
R161 drain_left.n13 drain_left.n12 7.3702
R162 drain_left drain_left.n17 6.19632
R163 drain_left.n4 drain_left.n0 5.81868
R164 drain_left.n13 drain_left.n9 5.81868
R165 drain_left.n5 drain_left.n1 3.44771
R166 drain_left.n14 drain_left.n10 3.44771
C0 plus drain_left 0.829965f
C1 drain_right minus 0.716298f
C2 drain_right source 3.71842f
C3 drain_left drain_right 0.564935f
C4 minus source 0.76729f
C5 drain_left minus 0.176975f
C6 drain_left source 3.72197f
C7 plus drain_right 0.274854f
C8 plus minus 2.82396f
C9 plus source 0.781362f
C10 drain_right a_n1220_n1288# 3.05876f
C11 drain_left a_n1220_n1288# 3.21266f
C12 source a_n1220_n1288# 2.325339f
C13 minus a_n1220_n1288# 3.868054f
C14 plus a_n1220_n1288# 4.601633f
C15 drain_left.n0 a_n1220_n1288# 0.03091f
C16 drain_left.n1 a_n1220_n1288# 0.068393f
C17 drain_left.t4 a_n1220_n1288# 0.051326f
C18 drain_left.n2 a_n1220_n1288# 0.053527f
C19 drain_left.n3 a_n1220_n1288# 0.017255f
C20 drain_left.n4 a_n1220_n1288# 0.01138f
C21 drain_left.n5 a_n1220_n1288# 0.150756f
C22 drain_left.n6 a_n1220_n1288# 0.048994f
C23 drain_left.t2 a_n1220_n1288# 0.033471f
C24 drain_left.t0 a_n1220_n1288# 0.033471f
C25 drain_left.n7 a_n1220_n1288# 0.210449f
C26 drain_left.n8 a_n1220_n1288# 0.755862f
C27 drain_left.n9 a_n1220_n1288# 0.03091f
C28 drain_left.n10 a_n1220_n1288# 0.068393f
C29 drain_left.t5 a_n1220_n1288# 0.051326f
C30 drain_left.n11 a_n1220_n1288# 0.053527f
C31 drain_left.n12 a_n1220_n1288# 0.017255f
C32 drain_left.n13 a_n1220_n1288# 0.01138f
C33 drain_left.n14 a_n1220_n1288# 0.150756f
C34 drain_left.n15 a_n1220_n1288# 0.049379f
C35 drain_left.t3 a_n1220_n1288# 0.033471f
C36 drain_left.t1 a_n1220_n1288# 0.033471f
C37 drain_left.n16 a_n1220_n1288# 0.210275f
C38 drain_left.n17 a_n1220_n1288# 0.488809f
C39 plus.t0 a_n1220_n1288# 0.075827f
C40 plus.n0 a_n1220_n1288# 0.057863f
C41 plus.t2 a_n1220_n1288# 0.066997f
C42 plus.n1 a_n1220_n1288# 0.046792f
C43 plus.t4 a_n1220_n1288# 0.075827f
C44 plus.n2 a_n1220_n1288# 0.057803f
C45 plus.n3 a_n1220_n1288# 0.325343f
C46 plus.t5 a_n1220_n1288# 0.075827f
C47 plus.n4 a_n1220_n1288# 0.057863f
C48 plus.t1 a_n1220_n1288# 0.075827f
C49 plus.t3 a_n1220_n1288# 0.066997f
C50 plus.n5 a_n1220_n1288# 0.046792f
C51 plus.n6 a_n1220_n1288# 0.057803f
C52 plus.n7 a_n1220_n1288# 0.799758f
C53 drain_right.n0 a_n1220_n1288# 0.031618f
C54 drain_right.n1 a_n1220_n1288# 0.06996f
C55 drain_right.t5 a_n1220_n1288# 0.052501f
C56 drain_right.n2 a_n1220_n1288# 0.054753f
C57 drain_right.n3 a_n1220_n1288# 0.01765f
C58 drain_right.n4 a_n1220_n1288# 0.011641f
C59 drain_right.n5 a_n1220_n1288# 0.154208f
C60 drain_right.n6 a_n1220_n1288# 0.050116f
C61 drain_right.t1 a_n1220_n1288# 0.034237f
C62 drain_right.t3 a_n1220_n1288# 0.034237f
C63 drain_right.n7 a_n1220_n1288# 0.215269f
C64 drain_right.n8 a_n1220_n1288# 0.730463f
C65 drain_right.t0 a_n1220_n1288# 0.034237f
C66 drain_right.t2 a_n1220_n1288# 0.034237f
C67 drain_right.n9 a_n1220_n1288# 0.216433f
C68 drain_right.n10 a_n1220_n1288# 0.031618f
C69 drain_right.n11 a_n1220_n1288# 0.06996f
C70 drain_right.t4 a_n1220_n1288# 0.052501f
C71 drain_right.n12 a_n1220_n1288# 0.054753f
C72 drain_right.n13 a_n1220_n1288# 0.01765f
C73 drain_right.n14 a_n1220_n1288# 0.011641f
C74 drain_right.n15 a_n1220_n1288# 0.154208f
C75 drain_right.n16 a_n1220_n1288# 0.049629f
C76 drain_right.n17 a_n1220_n1288# 0.508679f
C77 source.n0 a_n1220_n1288# 0.03906f
C78 source.n1 a_n1220_n1288# 0.086425f
C79 source.t0 a_n1220_n1288# 0.064858f
C80 source.n2 a_n1220_n1288# 0.06764f
C81 source.n3 a_n1220_n1288# 0.021805f
C82 source.n4 a_n1220_n1288# 0.01438f
C83 source.n5 a_n1220_n1288# 0.190502f
C84 source.n6 a_n1220_n1288# 0.042819f
C85 source.n7 a_n1220_n1288# 0.404055f
C86 source.t2 a_n1220_n1288# 0.042295f
C87 source.t5 a_n1220_n1288# 0.042295f
C88 source.n8 a_n1220_n1288# 0.22611f
C89 source.n9 a_n1220_n1288# 0.318821f
C90 source.n10 a_n1220_n1288# 0.03906f
C91 source.n11 a_n1220_n1288# 0.086425f
C92 source.t7 a_n1220_n1288# 0.064858f
C93 source.n12 a_n1220_n1288# 0.06764f
C94 source.n13 a_n1220_n1288# 0.021805f
C95 source.n14 a_n1220_n1288# 0.01438f
C96 source.n15 a_n1220_n1288# 0.190502f
C97 source.n16 a_n1220_n1288# 0.042819f
C98 source.n17 a_n1220_n1288# 0.132794f
C99 source.t6 a_n1220_n1288# 0.042295f
C100 source.t10 a_n1220_n1288# 0.042295f
C101 source.n18 a_n1220_n1288# 0.22611f
C102 source.n19 a_n1220_n1288# 0.886412f
C103 source.t1 a_n1220_n1288# 0.042295f
C104 source.t4 a_n1220_n1288# 0.042295f
C105 source.n20 a_n1220_n1288# 0.226109f
C106 source.n21 a_n1220_n1288# 0.886413f
C107 source.n22 a_n1220_n1288# 0.03906f
C108 source.n23 a_n1220_n1288# 0.086425f
C109 source.t3 a_n1220_n1288# 0.064858f
C110 source.n24 a_n1220_n1288# 0.06764f
C111 source.n25 a_n1220_n1288# 0.021805f
C112 source.n26 a_n1220_n1288# 0.01438f
C113 source.n27 a_n1220_n1288# 0.190502f
C114 source.n28 a_n1220_n1288# 0.042819f
C115 source.n29 a_n1220_n1288# 0.132794f
C116 source.t8 a_n1220_n1288# 0.042295f
C117 source.t11 a_n1220_n1288# 0.042295f
C118 source.n30 a_n1220_n1288# 0.226109f
C119 source.n31 a_n1220_n1288# 0.318822f
C120 source.n32 a_n1220_n1288# 0.03906f
C121 source.n33 a_n1220_n1288# 0.086425f
C122 source.t9 a_n1220_n1288# 0.064858f
C123 source.n34 a_n1220_n1288# 0.06764f
C124 source.n35 a_n1220_n1288# 0.021805f
C125 source.n36 a_n1220_n1288# 0.01438f
C126 source.n37 a_n1220_n1288# 0.190502f
C127 source.n38 a_n1220_n1288# 0.042819f
C128 source.n39 a_n1220_n1288# 0.260446f
C129 source.n40 a_n1220_n1288# 0.66164f
C130 minus.t3 a_n1220_n1288# 0.073804f
C131 minus.n0 a_n1220_n1288# 0.056319f
C132 minus.t1 a_n1220_n1288# 0.073804f
C133 minus.t5 a_n1220_n1288# 0.06521f
C134 minus.n1 a_n1220_n1288# 0.045543f
C135 minus.n2 a_n1220_n1288# 0.056261f
C136 minus.n3 a_n1220_n1288# 0.80688f
C137 minus.t0 a_n1220_n1288# 0.073804f
C138 minus.n4 a_n1220_n1288# 0.056319f
C139 minus.t4 a_n1220_n1288# 0.06521f
C140 minus.n5 a_n1220_n1288# 0.045543f
C141 minus.t2 a_n1220_n1288# 0.073804f
C142 minus.n6 a_n1220_n1288# 0.056261f
C143 minus.n7 a_n1220_n1288# 0.293938f
C144 minus.n8 a_n1220_n1288# 0.933044f
.ends

