* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X1 drain_left.t13 plus.t0 source.t21 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X2 drain_left.t12 plus.t1 source.t16 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 source.t8 minus.t0 drain_right.t13 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X4 drain_right.t12 minus.t1 source.t0 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X5 source.t11 minus.t2 drain_right.t11 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X6 drain_left.t11 plus.t2 source.t25 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X7 drain_left.t10 plus.t3 source.t27 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X8 drain_left.t9 plus.t4 source.t17 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X9 drain_left.t8 plus.t5 source.t22 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X10 source.t19 plus.t6 drain_left.t7 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X11 drain_right.t10 minus.t3 source.t2 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X12 drain_right.t9 minus.t4 source.t6 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 drain_right.t8 minus.t5 source.t3 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X14 drain_left.t6 plus.t7 source.t18 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X15 source.t23 plus.t8 drain_left.t5 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X16 source.t20 plus.t9 drain_left.t4 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X17 source.t15 plus.t10 drain_left.t3 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X18 source.t10 minus.t6 drain_right.t7 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_right.t6 minus.t7 source.t13 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X20 a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X21 drain_right.t5 minus.t8 source.t12 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X22 source.t26 plus.t11 drain_left.t2 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X24 source.t4 minus.t9 drain_right.t4 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X25 drain_right.t3 minus.t10 source.t7 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X26 drain_right.t2 minus.t11 source.t9 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X27 source.t14 plus.t12 drain_left.t1 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X28 drain_left.t0 plus.t13 source.t24 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X29 source.t1 minus.t12 drain_right.t1 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X30 source.t5 minus.t13 drain_right.t0 a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X31 a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# a_n2364_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
R0 plus.n8 plus.n7 161.3
R1 plus.n9 plus.n4 161.3
R2 plus.n11 plus.n10 161.3
R3 plus.n12 plus.n3 161.3
R4 plus.n14 plus.n13 161.3
R5 plus.n15 plus.n2 161.3
R6 plus.n17 plus.n16 161.3
R7 plus.n18 plus.n1 161.3
R8 plus.n19 plus.n0 161.3
R9 plus.n21 plus.n20 161.3
R10 plus.n30 plus.n29 161.3
R11 plus.n31 plus.n26 161.3
R12 plus.n33 plus.n32 161.3
R13 plus.n34 plus.n25 161.3
R14 plus.n36 plus.n35 161.3
R15 plus.n37 plus.n24 161.3
R16 plus.n39 plus.n38 161.3
R17 plus.n40 plus.n23 161.3
R18 plus.n41 plus.n22 161.3
R19 plus.n43 plus.n42 161.3
R20 plus.n5 plus.t4 148.822
R21 plus.n27 plus.t13 148.822
R22 plus.n20 plus.t0 124.977
R23 plus.n18 plus.t10 124.977
R24 plus.n2 plus.t3 124.977
R25 plus.n12 plus.t8 124.977
R26 plus.n4 plus.t1 124.977
R27 plus.n6 plus.t11 124.977
R28 plus.n42 plus.t7 124.977
R29 plus.n40 plus.t9 124.977
R30 plus.n24 plus.t5 124.977
R31 plus.n34 plus.t6 124.977
R32 plus.n26 plus.t2 124.977
R33 plus.n28 plus.t12 124.977
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus.n18 plus.n17 30.6732
R39 plus.n7 plus.n6 30.6732
R40 plus.n40 plus.n39 30.6732
R41 plus.n29 plus.n28 30.6732
R42 plus plus.n43 28.3191
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus.n19 plus.n18 13.146
R58 plus.n41 plus.n40 13.146
R59 plus plus.n21 8.50618
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n50 source.n48 289.615
R79 source.n36 source.n34 289.615
R80 source.n2 source.n0 289.615
R81 source.n16 source.n14 289.615
R82 source.n51 source.n50 185
R83 source.n37 source.n36 185
R84 source.n3 source.n2 185
R85 source.n17 source.n16 185
R86 source.t0 source.n49 167.117
R87 source.t24 source.n35 167.117
R88 source.t21 source.n1 167.117
R89 source.t13 source.n15 167.117
R90 source.n9 source.n8 84.1169
R91 source.n11 source.n10 84.1169
R92 source.n13 source.n12 84.1169
R93 source.n23 source.n22 84.1169
R94 source.n25 source.n24 84.1169
R95 source.n27 source.n26 84.1169
R96 source.n47 source.n46 84.1168
R97 source.n45 source.n44 84.1168
R98 source.n43 source.n42 84.1168
R99 source.n33 source.n32 84.1168
R100 source.n31 source.n30 84.1168
R101 source.n29 source.n28 84.1168
R102 source.n50 source.t0 52.3082
R103 source.n36 source.t24 52.3082
R104 source.n2 source.t21 52.3082
R105 source.n16 source.t13 52.3082
R106 source.n55 source.n54 31.4096
R107 source.n41 source.n40 31.4096
R108 source.n7 source.n6 31.4096
R109 source.n21 source.n20 31.4096
R110 source.n29 source.n27 15.4878
R111 source.n46 source.t9 9.9005
R112 source.n46 source.t11 9.9005
R113 source.n44 source.t7 9.9005
R114 source.n44 source.t4 9.9005
R115 source.n42 source.t12 9.9005
R116 source.n42 source.t10 9.9005
R117 source.n32 source.t25 9.9005
R118 source.n32 source.t14 9.9005
R119 source.n30 source.t22 9.9005
R120 source.n30 source.t19 9.9005
R121 source.n28 source.t18 9.9005
R122 source.n28 source.t20 9.9005
R123 source.n8 source.t27 9.9005
R124 source.n8 source.t15 9.9005
R125 source.n10 source.t16 9.9005
R126 source.n10 source.t23 9.9005
R127 source.n12 source.t17 9.9005
R128 source.n12 source.t26 9.9005
R129 source.n22 source.t3 9.9005
R130 source.n22 source.t8 9.9005
R131 source.n24 source.t6 9.9005
R132 source.n24 source.t1 9.9005
R133 source.n26 source.t2 9.9005
R134 source.n26 source.t5 9.9005
R135 source.n51 source.n49 9.71174
R136 source.n37 source.n35 9.71174
R137 source.n3 source.n1 9.71174
R138 source.n17 source.n15 9.71174
R139 source.n54 source.n53 9.45567
R140 source.n40 source.n39 9.45567
R141 source.n6 source.n5 9.45567
R142 source.n20 source.n19 9.45567
R143 source.n53 source.n52 9.3005
R144 source.n39 source.n38 9.3005
R145 source.n5 source.n4 9.3005
R146 source.n19 source.n18 9.3005
R147 source.n56 source.n7 8.893
R148 source.n54 source.n48 8.14595
R149 source.n40 source.n34 8.14595
R150 source.n6 source.n0 8.14595
R151 source.n20 source.n14 8.14595
R152 source.n52 source.n51 7.3702
R153 source.n38 source.n37 7.3702
R154 source.n4 source.n3 7.3702
R155 source.n18 source.n17 7.3702
R156 source.n52 source.n48 5.81868
R157 source.n38 source.n34 5.81868
R158 source.n4 source.n0 5.81868
R159 source.n18 source.n14 5.81868
R160 source.n56 source.n55 5.7074
R161 source.n53 source.n49 3.44771
R162 source.n39 source.n35 3.44771
R163 source.n5 source.n1 3.44771
R164 source.n19 source.n15 3.44771
R165 source.n21 source.n13 0.914293
R166 source.n43 source.n41 0.914293
R167 source.n27 source.n25 0.888431
R168 source.n25 source.n23 0.888431
R169 source.n23 source.n21 0.888431
R170 source.n13 source.n11 0.888431
R171 source.n11 source.n9 0.888431
R172 source.n9 source.n7 0.888431
R173 source.n31 source.n29 0.888431
R174 source.n33 source.n31 0.888431
R175 source.n41 source.n33 0.888431
R176 source.n45 source.n43 0.888431
R177 source.n47 source.n45 0.888431
R178 source.n55 source.n47 0.888431
R179 source source.n56 0.188
R180 drain_left.n2 drain_left.n0 289.615
R181 drain_left.n15 drain_left.n13 289.615
R182 drain_left.n3 drain_left.n2 185
R183 drain_left.n16 drain_left.n15 185
R184 drain_left.t6 drain_left.n1 167.117
R185 drain_left.t9 drain_left.n14 167.117
R186 drain_left.n11 drain_left.n9 101.683
R187 drain_left.n25 drain_left.n24 100.796
R188 drain_left.n23 drain_left.n22 100.796
R189 drain_left.n21 drain_left.n20 100.796
R190 drain_left.n11 drain_left.n10 100.796
R191 drain_left.n8 drain_left.n7 100.796
R192 drain_left.n2 drain_left.t6 52.3082
R193 drain_left.n15 drain_left.t9 52.3082
R194 drain_left.n8 drain_left.n6 48.9763
R195 drain_left.n21 drain_left.n19 48.9763
R196 drain_left drain_left.n12 24.8969
R197 drain_left.n9 drain_left.t1 9.9005
R198 drain_left.n9 drain_left.t0 9.9005
R199 drain_left.n10 drain_left.t7 9.9005
R200 drain_left.n10 drain_left.t11 9.9005
R201 drain_left.n7 drain_left.t4 9.9005
R202 drain_left.n7 drain_left.t8 9.9005
R203 drain_left.n24 drain_left.t3 9.9005
R204 drain_left.n24 drain_left.t13 9.9005
R205 drain_left.n22 drain_left.t5 9.9005
R206 drain_left.n22 drain_left.t10 9.9005
R207 drain_left.n20 drain_left.t2 9.9005
R208 drain_left.n20 drain_left.t12 9.9005
R209 drain_left.n3 drain_left.n1 9.71174
R210 drain_left.n16 drain_left.n14 9.71174
R211 drain_left.n6 drain_left.n5 9.45567
R212 drain_left.n19 drain_left.n18 9.45567
R213 drain_left.n5 drain_left.n4 9.3005
R214 drain_left.n18 drain_left.n17 9.3005
R215 drain_left.n6 drain_left.n0 8.14595
R216 drain_left.n19 drain_left.n13 8.14595
R217 drain_left.n4 drain_left.n3 7.3702
R218 drain_left.n17 drain_left.n16 7.3702
R219 drain_left drain_left.n25 6.54115
R220 drain_left.n4 drain_left.n0 5.81868
R221 drain_left.n17 drain_left.n13 5.81868
R222 drain_left.n5 drain_left.n1 3.44771
R223 drain_left.n18 drain_left.n14 3.44771
R224 drain_left.n23 drain_left.n21 0.888431
R225 drain_left.n25 drain_left.n23 0.888431
R226 drain_left.n12 drain_left.n8 0.611102
R227 drain_left.n12 drain_left.n11 0.167137
R228 minus.n21 minus.n20 161.3
R229 minus.n19 minus.n0 161.3
R230 minus.n18 minus.n17 161.3
R231 minus.n16 minus.n1 161.3
R232 minus.n15 minus.n14 161.3
R233 minus.n13 minus.n2 161.3
R234 minus.n12 minus.n11 161.3
R235 minus.n10 minus.n3 161.3
R236 minus.n9 minus.n8 161.3
R237 minus.n7 minus.n4 161.3
R238 minus.n43 minus.n42 161.3
R239 minus.n41 minus.n22 161.3
R240 minus.n40 minus.n39 161.3
R241 minus.n38 minus.n23 161.3
R242 minus.n37 minus.n36 161.3
R243 minus.n35 minus.n24 161.3
R244 minus.n34 minus.n33 161.3
R245 minus.n32 minus.n25 161.3
R246 minus.n31 minus.n30 161.3
R247 minus.n29 minus.n26 161.3
R248 minus.n5 minus.t7 148.822
R249 minus.n27 minus.t8 148.822
R250 minus.n6 minus.t0 124.977
R251 minus.n8 minus.t5 124.977
R252 minus.n12 minus.t12 124.977
R253 minus.n14 minus.t4 124.977
R254 minus.n18 minus.t13 124.977
R255 minus.n20 minus.t3 124.977
R256 minus.n28 minus.t6 124.977
R257 minus.n30 minus.t10 124.977
R258 minus.n34 minus.t9 124.977
R259 minus.n36 minus.t11 124.977
R260 minus.n40 minus.t2 124.977
R261 minus.n42 minus.t1 124.977
R262 minus.n5 minus.n4 44.9119
R263 minus.n27 minus.n26 44.9119
R264 minus.n20 minus.n19 35.055
R265 minus.n42 minus.n41 35.055
R266 minus.n7 minus.n6 30.6732
R267 minus.n18 minus.n1 30.6732
R268 minus.n29 minus.n28 30.6732
R269 minus.n40 minus.n23 30.6732
R270 minus.n44 minus.n21 30.6501
R271 minus.n8 minus.n3 26.2914
R272 minus.n14 minus.n13 26.2914
R273 minus.n30 minus.n25 26.2914
R274 minus.n36 minus.n35 26.2914
R275 minus.n12 minus.n3 21.9096
R276 minus.n13 minus.n12 21.9096
R277 minus.n34 minus.n25 21.9096
R278 minus.n35 minus.n34 21.9096
R279 minus.n6 minus.n5 17.739
R280 minus.n28 minus.n27 17.739
R281 minus.n8 minus.n7 17.5278
R282 minus.n14 minus.n1 17.5278
R283 minus.n30 minus.n29 17.5278
R284 minus.n36 minus.n23 17.5278
R285 minus.n19 minus.n18 13.146
R286 minus.n41 minus.n40 13.146
R287 minus.n44 minus.n43 6.65012
R288 minus.n21 minus.n0 0.189894
R289 minus.n17 minus.n0 0.189894
R290 minus.n17 minus.n16 0.189894
R291 minus.n16 minus.n15 0.189894
R292 minus.n15 minus.n2 0.189894
R293 minus.n11 minus.n2 0.189894
R294 minus.n11 minus.n10 0.189894
R295 minus.n10 minus.n9 0.189894
R296 minus.n9 minus.n4 0.189894
R297 minus.n31 minus.n26 0.189894
R298 minus.n32 minus.n31 0.189894
R299 minus.n33 minus.n32 0.189894
R300 minus.n33 minus.n24 0.189894
R301 minus.n37 minus.n24 0.189894
R302 minus.n38 minus.n37 0.189894
R303 minus.n39 minus.n38 0.189894
R304 minus.n39 minus.n22 0.189894
R305 minus.n43 minus.n22 0.189894
R306 minus minus.n44 0.188
R307 drain_right.n2 drain_right.n0 289.615
R308 drain_right.n20 drain_right.n18 289.615
R309 drain_right.n3 drain_right.n2 185
R310 drain_right.n21 drain_right.n20 185
R311 drain_right.t5 drain_right.n1 167.117
R312 drain_right.t10 drain_right.n19 167.117
R313 drain_right.n15 drain_right.n13 101.683
R314 drain_right.n11 drain_right.n9 101.683
R315 drain_right.n15 drain_right.n14 100.796
R316 drain_right.n17 drain_right.n16 100.796
R317 drain_right.n11 drain_right.n10 100.796
R318 drain_right.n8 drain_right.n7 100.796
R319 drain_right.n2 drain_right.t5 52.3082
R320 drain_right.n20 drain_right.t10 52.3082
R321 drain_right.n8 drain_right.n6 48.9763
R322 drain_right.n25 drain_right.n24 48.0884
R323 drain_right drain_right.n12 24.3437
R324 drain_right.n9 drain_right.t11 9.9005
R325 drain_right.n9 drain_right.t12 9.9005
R326 drain_right.n10 drain_right.t4 9.9005
R327 drain_right.n10 drain_right.t2 9.9005
R328 drain_right.n7 drain_right.t7 9.9005
R329 drain_right.n7 drain_right.t3 9.9005
R330 drain_right.n13 drain_right.t13 9.9005
R331 drain_right.n13 drain_right.t6 9.9005
R332 drain_right.n14 drain_right.t1 9.9005
R333 drain_right.n14 drain_right.t8 9.9005
R334 drain_right.n16 drain_right.t0 9.9005
R335 drain_right.n16 drain_right.t9 9.9005
R336 drain_right.n3 drain_right.n1 9.71174
R337 drain_right.n21 drain_right.n19 9.71174
R338 drain_right.n6 drain_right.n5 9.45567
R339 drain_right.n24 drain_right.n23 9.45567
R340 drain_right.n5 drain_right.n4 9.3005
R341 drain_right.n23 drain_right.n22 9.3005
R342 drain_right.n6 drain_right.n0 8.14595
R343 drain_right.n24 drain_right.n18 8.14595
R344 drain_right.n4 drain_right.n3 7.3702
R345 drain_right.n22 drain_right.n21 7.3702
R346 drain_right drain_right.n25 6.09718
R347 drain_right.n4 drain_right.n0 5.81868
R348 drain_right.n22 drain_right.n18 5.81868
R349 drain_right.n5 drain_right.n1 3.44771
R350 drain_right.n23 drain_right.n19 3.44771
R351 drain_right.n25 drain_right.n17 0.888431
R352 drain_right.n17 drain_right.n15 0.888431
R353 drain_right.n12 drain_right.n8 0.611102
R354 drain_right.n12 drain_right.n11 0.167137
C0 minus drain_right 1.96518f
C1 source minus 2.47625f
C2 drain_left drain_right 1.23072f
C3 source drain_left 5.78739f
C4 drain_left minus 0.179135f
C5 plus drain_right 0.396777f
C6 source plus 2.4903f
C7 plus minus 4.24844f
C8 plus drain_left 2.19788f
C9 source drain_right 5.78742f
C10 drain_right a_n2364_n1288# 4.32841f
C11 drain_left a_n2364_n1288# 5.07707f
C12 source a_n2364_n1288# 2.775385f
C13 minus a_n2364_n1288# 8.552599f
C14 plus a_n2364_n1288# 9.81833f
C15 drain_right.n0 a_n2364_n1288# 0.02751f
C16 drain_right.n1 a_n2364_n1288# 0.06087f
C17 drain_right.t5 a_n2364_n1288# 0.04568f
C18 drain_right.n2 a_n2364_n1288# 0.04764f
C19 drain_right.n3 a_n2364_n1288# 0.015357f
C20 drain_right.n4 a_n2364_n1288# 0.010128f
C21 drain_right.n5 a_n2364_n1288# 0.134173f
C22 drain_right.n6 a_n2364_n1288# 0.044806f
C23 drain_right.t7 a_n2364_n1288# 0.029789f
C24 drain_right.t3 a_n2364_n1288# 0.029789f
C25 drain_right.n7 a_n2364_n1288# 0.187145f
C26 drain_right.n8 a_n2364_n1288# 0.323999f
C27 drain_right.t11 a_n2364_n1288# 0.029789f
C28 drain_right.t12 a_n2364_n1288# 0.029789f
C29 drain_right.n9 a_n2364_n1288# 0.189413f
C30 drain_right.t4 a_n2364_n1288# 0.029789f
C31 drain_right.t2 a_n2364_n1288# 0.029789f
C32 drain_right.n10 a_n2364_n1288# 0.187145f
C33 drain_right.n11 a_n2364_n1288# 0.468378f
C34 drain_right.n12 a_n2364_n1288# 0.61406f
C35 drain_right.t13 a_n2364_n1288# 0.029789f
C36 drain_right.t6 a_n2364_n1288# 0.029789f
C37 drain_right.n13 a_n2364_n1288# 0.189414f
C38 drain_right.t1 a_n2364_n1288# 0.029789f
C39 drain_right.t8 a_n2364_n1288# 0.029789f
C40 drain_right.n14 a_n2364_n1288# 0.187146f
C41 drain_right.n15 a_n2364_n1288# 0.509561f
C42 drain_right.t0 a_n2364_n1288# 0.029789f
C43 drain_right.t9 a_n2364_n1288# 0.029789f
C44 drain_right.n16 a_n2364_n1288# 0.187146f
C45 drain_right.n17 a_n2364_n1288# 0.252118f
C46 drain_right.n18 a_n2364_n1288# 0.02751f
C47 drain_right.n19 a_n2364_n1288# 0.06087f
C48 drain_right.t10 a_n2364_n1288# 0.04568f
C49 drain_right.n20 a_n2364_n1288# 0.04764f
C50 drain_right.n21 a_n2364_n1288# 0.015357f
C51 drain_right.n22 a_n2364_n1288# 0.010128f
C52 drain_right.n23 a_n2364_n1288# 0.134173f
C53 drain_right.n24 a_n2364_n1288# 0.043181f
C54 drain_right.n25 a_n2364_n1288# 0.26286f
C55 minus.n0 a_n2364_n1288# 0.033866f
C56 minus.n1 a_n2364_n1288# 0.007685f
C57 minus.t13 a_n2364_n1288# 0.146824f
C58 minus.n2 a_n2364_n1288# 0.033866f
C59 minus.n3 a_n2364_n1288# 0.007685f
C60 minus.t12 a_n2364_n1288# 0.146824f
C61 minus.n4 a_n2364_n1288# 0.142692f
C62 minus.t7 a_n2364_n1288# 0.163183f
C63 minus.n5 a_n2364_n1288# 0.088645f
C64 minus.t0 a_n2364_n1288# 0.146824f
C65 minus.n6 a_n2364_n1288# 0.106257f
C66 minus.n7 a_n2364_n1288# 0.007685f
C67 minus.t5 a_n2364_n1288# 0.146824f
C68 minus.n8 a_n2364_n1288# 0.102062f
C69 minus.n9 a_n2364_n1288# 0.033866f
C70 minus.n10 a_n2364_n1288# 0.033866f
C71 minus.n11 a_n2364_n1288# 0.033866f
C72 minus.n12 a_n2364_n1288# 0.102062f
C73 minus.n13 a_n2364_n1288# 0.007685f
C74 minus.t4 a_n2364_n1288# 0.146824f
C75 minus.n14 a_n2364_n1288# 0.102062f
C76 minus.n15 a_n2364_n1288# 0.033866f
C77 minus.n16 a_n2364_n1288# 0.033866f
C78 minus.n17 a_n2364_n1288# 0.033866f
C79 minus.n18 a_n2364_n1288# 0.102062f
C80 minus.n19 a_n2364_n1288# 0.007685f
C81 minus.t3 a_n2364_n1288# 0.146824f
C82 minus.n20 a_n2364_n1288# 0.100809f
C83 minus.n21 a_n2364_n1288# 0.918299f
C84 minus.n22 a_n2364_n1288# 0.033866f
C85 minus.n23 a_n2364_n1288# 0.007685f
C86 minus.n24 a_n2364_n1288# 0.033866f
C87 minus.n25 a_n2364_n1288# 0.007685f
C88 minus.n26 a_n2364_n1288# 0.142692f
C89 minus.t8 a_n2364_n1288# 0.163183f
C90 minus.n27 a_n2364_n1288# 0.088645f
C91 minus.t6 a_n2364_n1288# 0.146824f
C92 minus.n28 a_n2364_n1288# 0.106257f
C93 minus.n29 a_n2364_n1288# 0.007685f
C94 minus.t10 a_n2364_n1288# 0.146824f
C95 minus.n30 a_n2364_n1288# 0.102062f
C96 minus.n31 a_n2364_n1288# 0.033866f
C97 minus.n32 a_n2364_n1288# 0.033866f
C98 minus.n33 a_n2364_n1288# 0.033866f
C99 minus.t9 a_n2364_n1288# 0.146824f
C100 minus.n34 a_n2364_n1288# 0.102062f
C101 minus.n35 a_n2364_n1288# 0.007685f
C102 minus.t11 a_n2364_n1288# 0.146824f
C103 minus.n36 a_n2364_n1288# 0.102062f
C104 minus.n37 a_n2364_n1288# 0.033866f
C105 minus.n38 a_n2364_n1288# 0.033866f
C106 minus.n39 a_n2364_n1288# 0.033866f
C107 minus.t2 a_n2364_n1288# 0.146824f
C108 minus.n40 a_n2364_n1288# 0.102062f
C109 minus.n41 a_n2364_n1288# 0.007685f
C110 minus.t1 a_n2364_n1288# 0.146824f
C111 minus.n42 a_n2364_n1288# 0.100809f
C112 minus.n43 a_n2364_n1288# 0.233301f
C113 minus.n44 a_n2364_n1288# 1.1259f
C114 drain_left.n0 a_n2364_n1288# 0.037469f
C115 drain_left.n1 a_n2364_n1288# 0.082905f
C116 drain_left.t6 a_n2364_n1288# 0.062216f
C117 drain_left.n2 a_n2364_n1288# 0.064885f
C118 drain_left.n3 a_n2364_n1288# 0.020916f
C119 drain_left.n4 a_n2364_n1288# 0.013795f
C120 drain_left.n5 a_n2364_n1288# 0.182743f
C121 drain_left.n6 a_n2364_n1288# 0.061025f
C122 drain_left.t4 a_n2364_n1288# 0.040573f
C123 drain_left.t8 a_n2364_n1288# 0.040573f
C124 drain_left.n7 a_n2364_n1288# 0.254891f
C125 drain_left.n8 a_n2364_n1288# 0.441285f
C126 drain_left.t1 a_n2364_n1288# 0.040573f
C127 drain_left.t0 a_n2364_n1288# 0.040573f
C128 drain_left.n9 a_n2364_n1288# 0.257979f
C129 drain_left.t7 a_n2364_n1288# 0.040573f
C130 drain_left.t11 a_n2364_n1288# 0.040573f
C131 drain_left.n10 a_n2364_n1288# 0.254891f
C132 drain_left.n11 a_n2364_n1288# 0.637928f
C133 drain_left.n12 a_n2364_n1288# 0.886392f
C134 drain_left.n13 a_n2364_n1288# 0.037469f
C135 drain_left.n14 a_n2364_n1288# 0.082905f
C136 drain_left.t9 a_n2364_n1288# 0.062216f
C137 drain_left.n15 a_n2364_n1288# 0.064885f
C138 drain_left.n16 a_n2364_n1288# 0.020916f
C139 drain_left.n17 a_n2364_n1288# 0.013795f
C140 drain_left.n18 a_n2364_n1288# 0.182743f
C141 drain_left.n19 a_n2364_n1288# 0.061025f
C142 drain_left.t2 a_n2364_n1288# 0.040573f
C143 drain_left.t12 a_n2364_n1288# 0.040573f
C144 drain_left.n20 a_n2364_n1288# 0.254892f
C145 drain_left.n21 a_n2364_n1288# 0.463249f
C146 drain_left.t5 a_n2364_n1288# 0.040573f
C147 drain_left.t10 a_n2364_n1288# 0.040573f
C148 drain_left.n22 a_n2364_n1288# 0.254892f
C149 drain_left.n23 a_n2364_n1288# 0.343384f
C150 drain_left.t3 a_n2364_n1288# 0.040573f
C151 drain_left.t13 a_n2364_n1288# 0.040573f
C152 drain_left.n24 a_n2364_n1288# 0.254892f
C153 drain_left.n25 a_n2364_n1288# 0.57045f
C154 source.n0 a_n2364_n1288# 0.048932f
C155 source.n1 a_n2364_n1288# 0.108268f
C156 source.t21 a_n2364_n1288# 0.08125f
C157 source.n2 a_n2364_n1288# 0.084735f
C158 source.n3 a_n2364_n1288# 0.027316f
C159 source.n4 a_n2364_n1288# 0.018015f
C160 source.n5 a_n2364_n1288# 0.23865f
C161 source.n6 a_n2364_n1288# 0.053641f
C162 source.n7 a_n2364_n1288# 0.572175f
C163 source.t27 a_n2364_n1288# 0.052985f
C164 source.t15 a_n2364_n1288# 0.052985f
C165 source.n8 a_n2364_n1288# 0.283258f
C166 source.n9 a_n2364_n1288# 0.452482f
C167 source.t16 a_n2364_n1288# 0.052985f
C168 source.t23 a_n2364_n1288# 0.052985f
C169 source.n10 a_n2364_n1288# 0.283258f
C170 source.n11 a_n2364_n1288# 0.452482f
C171 source.t17 a_n2364_n1288# 0.052985f
C172 source.t26 a_n2364_n1288# 0.052985f
C173 source.n12 a_n2364_n1288# 0.283258f
C174 source.n13 a_n2364_n1288# 0.455276f
C175 source.n14 a_n2364_n1288# 0.048932f
C176 source.n15 a_n2364_n1288# 0.108268f
C177 source.t13 a_n2364_n1288# 0.08125f
C178 source.n16 a_n2364_n1288# 0.084735f
C179 source.n17 a_n2364_n1288# 0.027316f
C180 source.n18 a_n2364_n1288# 0.018015f
C181 source.n19 a_n2364_n1288# 0.23865f
C182 source.n20 a_n2364_n1288# 0.053641f
C183 source.n21 a_n2364_n1288# 0.222232f
C184 source.t3 a_n2364_n1288# 0.052985f
C185 source.t8 a_n2364_n1288# 0.052985f
C186 source.n22 a_n2364_n1288# 0.283258f
C187 source.n23 a_n2364_n1288# 0.452482f
C188 source.t6 a_n2364_n1288# 0.052985f
C189 source.t1 a_n2364_n1288# 0.052985f
C190 source.n24 a_n2364_n1288# 0.283258f
C191 source.n25 a_n2364_n1288# 0.452482f
C192 source.t2 a_n2364_n1288# 0.052985f
C193 source.t5 a_n2364_n1288# 0.052985f
C194 source.n26 a_n2364_n1288# 0.283258f
C195 source.n27 a_n2364_n1288# 1.2222f
C196 source.t18 a_n2364_n1288# 0.052985f
C197 source.t20 a_n2364_n1288# 0.052985f
C198 source.n28 a_n2364_n1288# 0.283257f
C199 source.n29 a_n2364_n1288# 1.2222f
C200 source.t22 a_n2364_n1288# 0.052985f
C201 source.t19 a_n2364_n1288# 0.052985f
C202 source.n30 a_n2364_n1288# 0.283257f
C203 source.n31 a_n2364_n1288# 0.452484f
C204 source.t25 a_n2364_n1288# 0.052985f
C205 source.t14 a_n2364_n1288# 0.052985f
C206 source.n32 a_n2364_n1288# 0.283257f
C207 source.n33 a_n2364_n1288# 0.452484f
C208 source.n34 a_n2364_n1288# 0.048932f
C209 source.n35 a_n2364_n1288# 0.108268f
C210 source.t24 a_n2364_n1288# 0.08125f
C211 source.n36 a_n2364_n1288# 0.084735f
C212 source.n37 a_n2364_n1288# 0.027316f
C213 source.n38 a_n2364_n1288# 0.018015f
C214 source.n39 a_n2364_n1288# 0.23865f
C215 source.n40 a_n2364_n1288# 0.053641f
C216 source.n41 a_n2364_n1288# 0.222232f
C217 source.t12 a_n2364_n1288# 0.052985f
C218 source.t10 a_n2364_n1288# 0.052985f
C219 source.n42 a_n2364_n1288# 0.283257f
C220 source.n43 a_n2364_n1288# 0.455278f
C221 source.t7 a_n2364_n1288# 0.052985f
C222 source.t4 a_n2364_n1288# 0.052985f
C223 source.n44 a_n2364_n1288# 0.283257f
C224 source.n45 a_n2364_n1288# 0.452484f
C225 source.t9 a_n2364_n1288# 0.052985f
C226 source.t11 a_n2364_n1288# 0.052985f
C227 source.n46 a_n2364_n1288# 0.283257f
C228 source.n47 a_n2364_n1288# 0.452484f
C229 source.n48 a_n2364_n1288# 0.048932f
C230 source.n49 a_n2364_n1288# 0.108268f
C231 source.t0 a_n2364_n1288# 0.08125f
C232 source.n50 a_n2364_n1288# 0.084735f
C233 source.n51 a_n2364_n1288# 0.027316f
C234 source.n52 a_n2364_n1288# 0.018015f
C235 source.n53 a_n2364_n1288# 0.23865f
C236 source.n54 a_n2364_n1288# 0.053641f
C237 source.n55 a_n2364_n1288# 0.392959f
C238 source.n56 a_n2364_n1288# 0.845181f
C239 plus.n0 a_n2364_n1288# 0.045451f
C240 plus.t0 a_n2364_n1288# 0.197048f
C241 plus.t10 a_n2364_n1288# 0.197048f
C242 plus.n1 a_n2364_n1288# 0.045451f
C243 plus.t3 a_n2364_n1288# 0.197048f
C244 plus.n2 a_n2364_n1288# 0.136975f
C245 plus.n3 a_n2364_n1288# 0.045451f
C246 plus.t8 a_n2364_n1288# 0.197048f
C247 plus.t1 a_n2364_n1288# 0.197048f
C248 plus.n4 a_n2364_n1288# 0.136975f
C249 plus.t4 a_n2364_n1288# 0.219004f
C250 plus.n5 a_n2364_n1288# 0.118969f
C251 plus.t11 a_n2364_n1288# 0.197048f
C252 plus.n6 a_n2364_n1288# 0.142605f
C253 plus.n7 a_n2364_n1288# 0.010314f
C254 plus.n8 a_n2364_n1288# 0.191504f
C255 plus.n9 a_n2364_n1288# 0.045451f
C256 plus.n10 a_n2364_n1288# 0.045451f
C257 plus.n11 a_n2364_n1288# 0.010314f
C258 plus.n12 a_n2364_n1288# 0.136975f
C259 plus.n13 a_n2364_n1288# 0.010314f
C260 plus.n14 a_n2364_n1288# 0.045451f
C261 plus.n15 a_n2364_n1288# 0.045451f
C262 plus.n16 a_n2364_n1288# 0.045451f
C263 plus.n17 a_n2364_n1288# 0.010314f
C264 plus.n18 a_n2364_n1288# 0.136975f
C265 plus.n19 a_n2364_n1288# 0.010314f
C266 plus.n20 a_n2364_n1288# 0.135294f
C267 plus.n21 a_n2364_n1288# 0.34176f
C268 plus.n22 a_n2364_n1288# 0.045451f
C269 plus.t7 a_n2364_n1288# 0.197048f
C270 plus.n23 a_n2364_n1288# 0.045451f
C271 plus.t9 a_n2364_n1288# 0.197048f
C272 plus.t5 a_n2364_n1288# 0.197048f
C273 plus.n24 a_n2364_n1288# 0.136975f
C274 plus.n25 a_n2364_n1288# 0.045451f
C275 plus.t6 a_n2364_n1288# 0.197048f
C276 plus.t2 a_n2364_n1288# 0.197048f
C277 plus.n26 a_n2364_n1288# 0.136975f
C278 plus.t13 a_n2364_n1288# 0.219004f
C279 plus.n27 a_n2364_n1288# 0.118969f
C280 plus.t12 a_n2364_n1288# 0.197048f
C281 plus.n28 a_n2364_n1288# 0.142605f
C282 plus.n29 a_n2364_n1288# 0.010314f
C283 plus.n30 a_n2364_n1288# 0.191504f
C284 plus.n31 a_n2364_n1288# 0.045451f
C285 plus.n32 a_n2364_n1288# 0.045451f
C286 plus.n33 a_n2364_n1288# 0.010314f
C287 plus.n34 a_n2364_n1288# 0.136975f
C288 plus.n35 a_n2364_n1288# 0.010314f
C289 plus.n36 a_n2364_n1288# 0.045451f
C290 plus.n37 a_n2364_n1288# 0.045451f
C291 plus.n38 a_n2364_n1288# 0.045451f
C292 plus.n39 a_n2364_n1288# 0.010314f
C293 plus.n40 a_n2364_n1288# 0.136975f
C294 plus.n41 a_n2364_n1288# 0.010314f
C295 plus.n42 a_n2364_n1288# 0.135294f
C296 plus.n43 a_n2364_n1288# 1.17345f
.ends

