* NGSPICE file created from diffpair253.ext - technology: sky130A

.subckt diffpair253 minus drain_right drain_left source plus
X0 a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X1 drain_right.t7 minus.t0 source.t10 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X3 drain_left.t7 plus.t0 source.t1 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X5 source.t14 plus.t1 drain_left.t6 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X6 source.t11 minus.t1 drain_right.t6 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X8 source.t4 plus.t2 drain_left.t5 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X9 drain_left.t4 plus.t3 source.t0 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X10 drain_left.t3 plus.t4 source.t15 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X11 drain_right.t5 minus.t2 source.t6 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X12 source.t2 plus.t5 drain_left.t2 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X13 drain_left.t1 plus.t6 source.t3 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X14 source.t12 minus.t3 drain_right.t4 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X15 source.t13 minus.t4 drain_right.t3 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X16 source.t7 minus.t5 drain_right.t2 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X17 drain_right.t1 minus.t6 source.t8 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X18 drain_right.t0 minus.t7 source.t9 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X19 source.t5 plus.t7 drain_left.t0 a_n1246_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n5 minus.t5 922.739
R1 minus.n1 minus.t2 922.739
R2 minus.n12 minus.t6 922.739
R3 minus.n8 minus.t4 922.739
R4 minus.n4 minus.t0 879.65
R5 minus.n2 minus.t1 879.65
R6 minus.n11 minus.t3 879.65
R7 minus.n9 minus.t7 879.65
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 38.7066
R15 minus.n3 minus.n2 38.7066
R16 minus.n10 minus.n9 38.7066
R17 minus.n11 minus.n10 38.7066
R18 minus.n5 minus.n4 34.3247
R19 minus.n2 minus.n1 34.3247
R20 minus.n9 minus.n8 34.3247
R21 minus.n12 minus.n11 34.3247
R22 minus.n14 minus.n6 29.2391
R23 minus.n14 minus.n13 6.44368
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n258 source.n232 289.615
R28 source.n224 source.n198 289.615
R29 source.n192 source.n166 289.615
R30 source.n158 source.n132 289.615
R31 source.n26 source.n0 289.615
R32 source.n60 source.n34 289.615
R33 source.n92 source.n66 289.615
R34 source.n126 source.n100 289.615
R35 source.n243 source.n242 185
R36 source.n240 source.n239 185
R37 source.n249 source.n248 185
R38 source.n251 source.n250 185
R39 source.n236 source.n235 185
R40 source.n257 source.n256 185
R41 source.n259 source.n258 185
R42 source.n209 source.n208 185
R43 source.n206 source.n205 185
R44 source.n215 source.n214 185
R45 source.n217 source.n216 185
R46 source.n202 source.n201 185
R47 source.n223 source.n222 185
R48 source.n225 source.n224 185
R49 source.n177 source.n176 185
R50 source.n174 source.n173 185
R51 source.n183 source.n182 185
R52 source.n185 source.n184 185
R53 source.n170 source.n169 185
R54 source.n191 source.n190 185
R55 source.n193 source.n192 185
R56 source.n143 source.n142 185
R57 source.n140 source.n139 185
R58 source.n149 source.n148 185
R59 source.n151 source.n150 185
R60 source.n136 source.n135 185
R61 source.n157 source.n156 185
R62 source.n159 source.n158 185
R63 source.n27 source.n26 185
R64 source.n25 source.n24 185
R65 source.n4 source.n3 185
R66 source.n19 source.n18 185
R67 source.n17 source.n16 185
R68 source.n8 source.n7 185
R69 source.n11 source.n10 185
R70 source.n61 source.n60 185
R71 source.n59 source.n58 185
R72 source.n38 source.n37 185
R73 source.n53 source.n52 185
R74 source.n51 source.n50 185
R75 source.n42 source.n41 185
R76 source.n45 source.n44 185
R77 source.n93 source.n92 185
R78 source.n91 source.n90 185
R79 source.n70 source.n69 185
R80 source.n85 source.n84 185
R81 source.n83 source.n82 185
R82 source.n74 source.n73 185
R83 source.n77 source.n76 185
R84 source.n127 source.n126 185
R85 source.n125 source.n124 185
R86 source.n104 source.n103 185
R87 source.n119 source.n118 185
R88 source.n117 source.n116 185
R89 source.n108 source.n107 185
R90 source.n111 source.n110 185
R91 source.t8 source.n241 147.661
R92 source.t13 source.n207 147.661
R93 source.t15 source.n175 147.661
R94 source.t14 source.n141 147.661
R95 source.t3 source.n9 147.661
R96 source.t4 source.n43 147.661
R97 source.t6 source.n75 147.661
R98 source.t7 source.n109 147.661
R99 source.n242 source.n239 104.615
R100 source.n249 source.n239 104.615
R101 source.n250 source.n249 104.615
R102 source.n250 source.n235 104.615
R103 source.n257 source.n235 104.615
R104 source.n258 source.n257 104.615
R105 source.n208 source.n205 104.615
R106 source.n215 source.n205 104.615
R107 source.n216 source.n215 104.615
R108 source.n216 source.n201 104.615
R109 source.n223 source.n201 104.615
R110 source.n224 source.n223 104.615
R111 source.n176 source.n173 104.615
R112 source.n183 source.n173 104.615
R113 source.n184 source.n183 104.615
R114 source.n184 source.n169 104.615
R115 source.n191 source.n169 104.615
R116 source.n192 source.n191 104.615
R117 source.n142 source.n139 104.615
R118 source.n149 source.n139 104.615
R119 source.n150 source.n149 104.615
R120 source.n150 source.n135 104.615
R121 source.n157 source.n135 104.615
R122 source.n158 source.n157 104.615
R123 source.n26 source.n25 104.615
R124 source.n25 source.n3 104.615
R125 source.n18 source.n3 104.615
R126 source.n18 source.n17 104.615
R127 source.n17 source.n7 104.615
R128 source.n10 source.n7 104.615
R129 source.n60 source.n59 104.615
R130 source.n59 source.n37 104.615
R131 source.n52 source.n37 104.615
R132 source.n52 source.n51 104.615
R133 source.n51 source.n41 104.615
R134 source.n44 source.n41 104.615
R135 source.n92 source.n91 104.615
R136 source.n91 source.n69 104.615
R137 source.n84 source.n69 104.615
R138 source.n84 source.n83 104.615
R139 source.n83 source.n73 104.615
R140 source.n76 source.n73 104.615
R141 source.n126 source.n125 104.615
R142 source.n125 source.n103 104.615
R143 source.n118 source.n103 104.615
R144 source.n118 source.n117 104.615
R145 source.n117 source.n107 104.615
R146 source.n110 source.n107 104.615
R147 source.n242 source.t8 52.3082
R148 source.n208 source.t13 52.3082
R149 source.n176 source.t15 52.3082
R150 source.n142 source.t14 52.3082
R151 source.n10 source.t3 52.3082
R152 source.n44 source.t4 52.3082
R153 source.n76 source.t6 52.3082
R154 source.n110 source.t7 52.3082
R155 source.n33 source.n32 50.512
R156 source.n99 source.n98 50.512
R157 source.n231 source.n230 50.5119
R158 source.n165 source.n164 50.5119
R159 source.n263 source.n262 32.1853
R160 source.n229 source.n228 32.1853
R161 source.n197 source.n196 32.1853
R162 source.n163 source.n162 32.1853
R163 source.n31 source.n30 32.1853
R164 source.n65 source.n64 32.1853
R165 source.n97 source.n96 32.1853
R166 source.n131 source.n130 32.1853
R167 source.n163 source.n131 17.1992
R168 source.n243 source.n241 15.6674
R169 source.n209 source.n207 15.6674
R170 source.n177 source.n175 15.6674
R171 source.n143 source.n141 15.6674
R172 source.n11 source.n9 15.6674
R173 source.n45 source.n43 15.6674
R174 source.n77 source.n75 15.6674
R175 source.n111 source.n109 15.6674
R176 source.n244 source.n240 12.8005
R177 source.n210 source.n206 12.8005
R178 source.n178 source.n174 12.8005
R179 source.n144 source.n140 12.8005
R180 source.n12 source.n8 12.8005
R181 source.n46 source.n42 12.8005
R182 source.n78 source.n74 12.8005
R183 source.n112 source.n108 12.8005
R184 source.n248 source.n247 12.0247
R185 source.n214 source.n213 12.0247
R186 source.n182 source.n181 12.0247
R187 source.n148 source.n147 12.0247
R188 source.n16 source.n15 12.0247
R189 source.n50 source.n49 12.0247
R190 source.n82 source.n81 12.0247
R191 source.n116 source.n115 12.0247
R192 source.n264 source.n31 11.7078
R193 source.n251 source.n238 11.249
R194 source.n217 source.n204 11.249
R195 source.n185 source.n172 11.249
R196 source.n151 source.n138 11.249
R197 source.n19 source.n6 11.249
R198 source.n53 source.n40 11.249
R199 source.n85 source.n72 11.249
R200 source.n119 source.n106 11.249
R201 source.n252 source.n236 10.4732
R202 source.n218 source.n202 10.4732
R203 source.n186 source.n170 10.4732
R204 source.n152 source.n136 10.4732
R205 source.n20 source.n4 10.4732
R206 source.n54 source.n38 10.4732
R207 source.n86 source.n70 10.4732
R208 source.n120 source.n104 10.4732
R209 source.n256 source.n255 9.69747
R210 source.n222 source.n221 9.69747
R211 source.n190 source.n189 9.69747
R212 source.n156 source.n155 9.69747
R213 source.n24 source.n23 9.69747
R214 source.n58 source.n57 9.69747
R215 source.n90 source.n89 9.69747
R216 source.n124 source.n123 9.69747
R217 source.n262 source.n261 9.45567
R218 source.n228 source.n227 9.45567
R219 source.n196 source.n195 9.45567
R220 source.n162 source.n161 9.45567
R221 source.n30 source.n29 9.45567
R222 source.n64 source.n63 9.45567
R223 source.n96 source.n95 9.45567
R224 source.n130 source.n129 9.45567
R225 source.n261 source.n260 9.3005
R226 source.n234 source.n233 9.3005
R227 source.n255 source.n254 9.3005
R228 source.n253 source.n252 9.3005
R229 source.n238 source.n237 9.3005
R230 source.n247 source.n246 9.3005
R231 source.n245 source.n244 9.3005
R232 source.n227 source.n226 9.3005
R233 source.n200 source.n199 9.3005
R234 source.n221 source.n220 9.3005
R235 source.n219 source.n218 9.3005
R236 source.n204 source.n203 9.3005
R237 source.n213 source.n212 9.3005
R238 source.n211 source.n210 9.3005
R239 source.n195 source.n194 9.3005
R240 source.n168 source.n167 9.3005
R241 source.n189 source.n188 9.3005
R242 source.n187 source.n186 9.3005
R243 source.n172 source.n171 9.3005
R244 source.n181 source.n180 9.3005
R245 source.n179 source.n178 9.3005
R246 source.n161 source.n160 9.3005
R247 source.n134 source.n133 9.3005
R248 source.n155 source.n154 9.3005
R249 source.n153 source.n152 9.3005
R250 source.n138 source.n137 9.3005
R251 source.n147 source.n146 9.3005
R252 source.n145 source.n144 9.3005
R253 source.n29 source.n28 9.3005
R254 source.n2 source.n1 9.3005
R255 source.n23 source.n22 9.3005
R256 source.n21 source.n20 9.3005
R257 source.n6 source.n5 9.3005
R258 source.n15 source.n14 9.3005
R259 source.n13 source.n12 9.3005
R260 source.n63 source.n62 9.3005
R261 source.n36 source.n35 9.3005
R262 source.n57 source.n56 9.3005
R263 source.n55 source.n54 9.3005
R264 source.n40 source.n39 9.3005
R265 source.n49 source.n48 9.3005
R266 source.n47 source.n46 9.3005
R267 source.n95 source.n94 9.3005
R268 source.n68 source.n67 9.3005
R269 source.n89 source.n88 9.3005
R270 source.n87 source.n86 9.3005
R271 source.n72 source.n71 9.3005
R272 source.n81 source.n80 9.3005
R273 source.n79 source.n78 9.3005
R274 source.n129 source.n128 9.3005
R275 source.n102 source.n101 9.3005
R276 source.n123 source.n122 9.3005
R277 source.n121 source.n120 9.3005
R278 source.n106 source.n105 9.3005
R279 source.n115 source.n114 9.3005
R280 source.n113 source.n112 9.3005
R281 source.n259 source.n234 8.92171
R282 source.n225 source.n200 8.92171
R283 source.n193 source.n168 8.92171
R284 source.n159 source.n134 8.92171
R285 source.n27 source.n2 8.92171
R286 source.n61 source.n36 8.92171
R287 source.n93 source.n68 8.92171
R288 source.n127 source.n102 8.92171
R289 source.n260 source.n232 8.14595
R290 source.n226 source.n198 8.14595
R291 source.n194 source.n166 8.14595
R292 source.n160 source.n132 8.14595
R293 source.n28 source.n0 8.14595
R294 source.n62 source.n34 8.14595
R295 source.n94 source.n66 8.14595
R296 source.n128 source.n100 8.14595
R297 source.n262 source.n232 5.81868
R298 source.n228 source.n198 5.81868
R299 source.n196 source.n166 5.81868
R300 source.n162 source.n132 5.81868
R301 source.n30 source.n0 5.81868
R302 source.n64 source.n34 5.81868
R303 source.n96 source.n66 5.81868
R304 source.n130 source.n100 5.81868
R305 source.n264 source.n263 5.49188
R306 source.n260 source.n259 5.04292
R307 source.n226 source.n225 5.04292
R308 source.n194 source.n193 5.04292
R309 source.n160 source.n159 5.04292
R310 source.n28 source.n27 5.04292
R311 source.n62 source.n61 5.04292
R312 source.n94 source.n93 5.04292
R313 source.n128 source.n127 5.04292
R314 source.n245 source.n241 4.38594
R315 source.n211 source.n207 4.38594
R316 source.n179 source.n175 4.38594
R317 source.n145 source.n141 4.38594
R318 source.n13 source.n9 4.38594
R319 source.n47 source.n43 4.38594
R320 source.n79 source.n75 4.38594
R321 source.n113 source.n109 4.38594
R322 source.n256 source.n234 4.26717
R323 source.n222 source.n200 4.26717
R324 source.n190 source.n168 4.26717
R325 source.n156 source.n134 4.26717
R326 source.n24 source.n2 4.26717
R327 source.n58 source.n36 4.26717
R328 source.n90 source.n68 4.26717
R329 source.n124 source.n102 4.26717
R330 source.n255 source.n236 3.49141
R331 source.n221 source.n202 3.49141
R332 source.n189 source.n170 3.49141
R333 source.n155 source.n136 3.49141
R334 source.n23 source.n4 3.49141
R335 source.n57 source.n38 3.49141
R336 source.n89 source.n70 3.49141
R337 source.n123 source.n104 3.49141
R338 source.n230 source.t9 3.3005
R339 source.n230 source.t12 3.3005
R340 source.n164 source.t0 3.3005
R341 source.n164 source.t2 3.3005
R342 source.n32 source.t1 3.3005
R343 source.n32 source.t5 3.3005
R344 source.n98 source.t10 3.3005
R345 source.n98 source.t11 3.3005
R346 source.n252 source.n251 2.71565
R347 source.n218 source.n217 2.71565
R348 source.n186 source.n185 2.71565
R349 source.n152 source.n151 2.71565
R350 source.n20 source.n19 2.71565
R351 source.n54 source.n53 2.71565
R352 source.n86 source.n85 2.71565
R353 source.n120 source.n119 2.71565
R354 source.n248 source.n238 1.93989
R355 source.n214 source.n204 1.93989
R356 source.n182 source.n172 1.93989
R357 source.n148 source.n138 1.93989
R358 source.n16 source.n6 1.93989
R359 source.n50 source.n40 1.93989
R360 source.n82 source.n72 1.93989
R361 source.n116 source.n106 1.93989
R362 source.n247 source.n240 1.16414
R363 source.n213 source.n206 1.16414
R364 source.n181 source.n174 1.16414
R365 source.n147 source.n140 1.16414
R366 source.n15 source.n8 1.16414
R367 source.n49 source.n42 1.16414
R368 source.n81 source.n74 1.16414
R369 source.n115 source.n108 1.16414
R370 source.n97 source.n65 0.470328
R371 source.n229 source.n197 0.470328
R372 source.n131 source.n99 0.457397
R373 source.n99 source.n97 0.457397
R374 source.n65 source.n33 0.457397
R375 source.n33 source.n31 0.457397
R376 source.n165 source.n163 0.457397
R377 source.n197 source.n165 0.457397
R378 source.n231 source.n229 0.457397
R379 source.n263 source.n231 0.457397
R380 source.n244 source.n243 0.388379
R381 source.n210 source.n209 0.388379
R382 source.n178 source.n177 0.388379
R383 source.n144 source.n143 0.388379
R384 source.n12 source.n11 0.388379
R385 source.n46 source.n45 0.388379
R386 source.n78 source.n77 0.388379
R387 source.n112 source.n111 0.388379
R388 source source.n264 0.188
R389 source.n246 source.n245 0.155672
R390 source.n246 source.n237 0.155672
R391 source.n253 source.n237 0.155672
R392 source.n254 source.n253 0.155672
R393 source.n254 source.n233 0.155672
R394 source.n261 source.n233 0.155672
R395 source.n212 source.n211 0.155672
R396 source.n212 source.n203 0.155672
R397 source.n219 source.n203 0.155672
R398 source.n220 source.n219 0.155672
R399 source.n220 source.n199 0.155672
R400 source.n227 source.n199 0.155672
R401 source.n180 source.n179 0.155672
R402 source.n180 source.n171 0.155672
R403 source.n187 source.n171 0.155672
R404 source.n188 source.n187 0.155672
R405 source.n188 source.n167 0.155672
R406 source.n195 source.n167 0.155672
R407 source.n146 source.n145 0.155672
R408 source.n146 source.n137 0.155672
R409 source.n153 source.n137 0.155672
R410 source.n154 source.n153 0.155672
R411 source.n154 source.n133 0.155672
R412 source.n161 source.n133 0.155672
R413 source.n29 source.n1 0.155672
R414 source.n22 source.n1 0.155672
R415 source.n22 source.n21 0.155672
R416 source.n21 source.n5 0.155672
R417 source.n14 source.n5 0.155672
R418 source.n14 source.n13 0.155672
R419 source.n63 source.n35 0.155672
R420 source.n56 source.n35 0.155672
R421 source.n56 source.n55 0.155672
R422 source.n55 source.n39 0.155672
R423 source.n48 source.n39 0.155672
R424 source.n48 source.n47 0.155672
R425 source.n95 source.n67 0.155672
R426 source.n88 source.n67 0.155672
R427 source.n88 source.n87 0.155672
R428 source.n87 source.n71 0.155672
R429 source.n80 source.n71 0.155672
R430 source.n80 source.n79 0.155672
R431 source.n129 source.n101 0.155672
R432 source.n122 source.n101 0.155672
R433 source.n122 source.n121 0.155672
R434 source.n121 source.n105 0.155672
R435 source.n114 source.n105 0.155672
R436 source.n114 source.n113 0.155672
R437 drain_right.n5 drain_right.n3 67.6476
R438 drain_right.n2 drain_right.n1 67.3638
R439 drain_right.n2 drain_right.n0 67.3638
R440 drain_right.n5 drain_right.n4 67.1908
R441 drain_right drain_right.n2 23.8675
R442 drain_right drain_right.n5 6.11011
R443 drain_right.n1 drain_right.t4 3.3005
R444 drain_right.n1 drain_right.t1 3.3005
R445 drain_right.n0 drain_right.t3 3.3005
R446 drain_right.n0 drain_right.t0 3.3005
R447 drain_right.n3 drain_right.t6 3.3005
R448 drain_right.n3 drain_right.t5 3.3005
R449 drain_right.n4 drain_right.t2 3.3005
R450 drain_right.n4 drain_right.t7 3.3005
R451 plus.n1 plus.t2 922.739
R452 plus.n5 plus.t6 922.739
R453 plus.n8 plus.t4 922.739
R454 plus.n12 plus.t1 922.739
R455 plus.n2 plus.t0 879.65
R456 plus.n4 plus.t7 879.65
R457 plus.n9 plus.t5 879.65
R458 plus.n11 plus.t3 879.65
R459 plus.n1 plus.n0 161.489
R460 plus.n8 plus.n7 161.489
R461 plus.n3 plus.n0 161.3
R462 plus.n6 plus.n5 161.3
R463 plus.n10 plus.n7 161.3
R464 plus.n13 plus.n12 161.3
R465 plus.n3 plus.n2 38.7066
R466 plus.n4 plus.n3 38.7066
R467 plus.n11 plus.n10 38.7066
R468 plus.n10 plus.n9 38.7066
R469 plus.n2 plus.n1 34.3247
R470 plus.n5 plus.n4 34.3247
R471 plus.n12 plus.n11 34.3247
R472 plus.n9 plus.n8 34.3247
R473 plus plus.n13 25.393
R474 plus plus.n6 9.81489
R475 plus.n6 plus.n0 0.189894
R476 plus.n13 plus.n7 0.189894
R477 drain_left.n5 drain_left.n3 67.6477
R478 drain_left.n2 drain_left.n1 67.3638
R479 drain_left.n2 drain_left.n0 67.3638
R480 drain_left.n5 drain_left.n4 67.1907
R481 drain_left drain_left.n2 24.4208
R482 drain_left drain_left.n5 6.11011
R483 drain_left.n1 drain_left.t2 3.3005
R484 drain_left.n1 drain_left.t3 3.3005
R485 drain_left.n0 drain_left.t6 3.3005
R486 drain_left.n0 drain_left.t4 3.3005
R487 drain_left.n4 drain_left.t0 3.3005
R488 drain_left.n4 drain_left.t1 3.3005
R489 drain_left.n3 drain_left.t5 3.3005
R490 drain_left.n3 drain_left.t7 3.3005
C0 drain_left plus 1.60447f
C1 source minus 1.29278f
C2 source drain_right 10.7096f
C3 source drain_left 10.7111f
C4 source plus 1.30679f
C5 drain_right minus 1.48767f
C6 drain_left minus 0.17017f
C7 minus plus 3.59723f
C8 drain_right drain_left 0.58123f
C9 drain_right plus 0.269775f
C10 drain_right a_n1246_n2088# 4.20884f
C11 drain_left a_n1246_n2088# 4.37423f
C12 source a_n1246_n2088# 5.053015f
C13 minus a_n1246_n2088# 4.321347f
C14 plus a_n1246_n2088# 5.161171f
C15 drain_left.t6 a_n1246_n2088# 0.147063f
C16 drain_left.t4 a_n1246_n2088# 0.147063f
C17 drain_left.n0 a_n1246_n2088# 1.22736f
C18 drain_left.t2 a_n1246_n2088# 0.147063f
C19 drain_left.t3 a_n1246_n2088# 0.147063f
C20 drain_left.n1 a_n1246_n2088# 1.22736f
C21 drain_left.n2 a_n1246_n2088# 1.57827f
C22 drain_left.t5 a_n1246_n2088# 0.147063f
C23 drain_left.t7 a_n1246_n2088# 0.147063f
C24 drain_left.n3 a_n1246_n2088# 1.22891f
C25 drain_left.t0 a_n1246_n2088# 0.147063f
C26 drain_left.t1 a_n1246_n2088# 0.147063f
C27 drain_left.n4 a_n1246_n2088# 1.22651f
C28 drain_left.n5 a_n1246_n2088# 0.950073f
C29 plus.n0 a_n1246_n2088# 0.072718f
C30 plus.t7 a_n1246_n2088# 0.114184f
C31 plus.t0 a_n1246_n2088# 0.114184f
C32 plus.t2 a_n1246_n2088# 0.116786f
C33 plus.n1 a_n1246_n2088# 0.064881f
C34 plus.n2 a_n1246_n2088# 0.055844f
C35 plus.n3 a_n1246_n2088# 0.011696f
C36 plus.n4 a_n1246_n2088# 0.055844f
C37 plus.t6 a_n1246_n2088# 0.116786f
C38 plus.n5 a_n1246_n2088# 0.064835f
C39 plus.n6 a_n1246_n2088# 0.281543f
C40 plus.n7 a_n1246_n2088# 0.072718f
C41 plus.t1 a_n1246_n2088# 0.116786f
C42 plus.t3 a_n1246_n2088# 0.114184f
C43 plus.t5 a_n1246_n2088# 0.114184f
C44 plus.t4 a_n1246_n2088# 0.116786f
C45 plus.n8 a_n1246_n2088# 0.064881f
C46 plus.n9 a_n1246_n2088# 0.055844f
C47 plus.n10 a_n1246_n2088# 0.011696f
C48 plus.n11 a_n1246_n2088# 0.055844f
C49 plus.n12 a_n1246_n2088# 0.064835f
C50 plus.n13 a_n1246_n2088# 0.750151f
C51 drain_right.t3 a_n1246_n2088# 0.14875f
C52 drain_right.t0 a_n1246_n2088# 0.14875f
C53 drain_right.n0 a_n1246_n2088# 1.24143f
C54 drain_right.t4 a_n1246_n2088# 0.14875f
C55 drain_right.t1 a_n1246_n2088# 0.14875f
C56 drain_right.n1 a_n1246_n2088# 1.24143f
C57 drain_right.n2 a_n1246_n2088# 1.53203f
C58 drain_right.t6 a_n1246_n2088# 0.14875f
C59 drain_right.t5 a_n1246_n2088# 0.14875f
C60 drain_right.n3 a_n1246_n2088# 1.243f
C61 drain_right.t2 a_n1246_n2088# 0.14875f
C62 drain_right.t7 a_n1246_n2088# 0.14875f
C63 drain_right.n4 a_n1246_n2088# 1.24058f
C64 drain_right.n5 a_n1246_n2088# 0.96097f
C65 source.n0 a_n1246_n2088# 0.03474f
C66 source.n1 a_n1246_n2088# 0.024716f
C67 source.n2 a_n1246_n2088# 0.013281f
C68 source.n3 a_n1246_n2088# 0.031392f
C69 source.n4 a_n1246_n2088# 0.014062f
C70 source.n5 a_n1246_n2088# 0.024716f
C71 source.n6 a_n1246_n2088# 0.013281f
C72 source.n7 a_n1246_n2088# 0.031392f
C73 source.n8 a_n1246_n2088# 0.014062f
C74 source.n9 a_n1246_n2088# 0.105766f
C75 source.t3 a_n1246_n2088# 0.051165f
C76 source.n10 a_n1246_n2088# 0.023544f
C77 source.n11 a_n1246_n2088# 0.018543f
C78 source.n12 a_n1246_n2088# 0.013281f
C79 source.n13 a_n1246_n2088# 0.588087f
C80 source.n14 a_n1246_n2088# 0.024716f
C81 source.n15 a_n1246_n2088# 0.013281f
C82 source.n16 a_n1246_n2088# 0.014062f
C83 source.n17 a_n1246_n2088# 0.031392f
C84 source.n18 a_n1246_n2088# 0.031392f
C85 source.n19 a_n1246_n2088# 0.014062f
C86 source.n20 a_n1246_n2088# 0.013281f
C87 source.n21 a_n1246_n2088# 0.024716f
C88 source.n22 a_n1246_n2088# 0.024716f
C89 source.n23 a_n1246_n2088# 0.013281f
C90 source.n24 a_n1246_n2088# 0.014062f
C91 source.n25 a_n1246_n2088# 0.031392f
C92 source.n26 a_n1246_n2088# 0.067958f
C93 source.n27 a_n1246_n2088# 0.014062f
C94 source.n28 a_n1246_n2088# 0.013281f
C95 source.n29 a_n1246_n2088# 0.057129f
C96 source.n30 a_n1246_n2088# 0.038025f
C97 source.n31 a_n1246_n2088# 0.586888f
C98 source.t1 a_n1246_n2088# 0.117187f
C99 source.t5 a_n1246_n2088# 0.117187f
C100 source.n32 a_n1246_n2088# 0.91266f
C101 source.n33 a_n1246_n2088# 0.304461f
C102 source.n34 a_n1246_n2088# 0.03474f
C103 source.n35 a_n1246_n2088# 0.024716f
C104 source.n36 a_n1246_n2088# 0.013281f
C105 source.n37 a_n1246_n2088# 0.031392f
C106 source.n38 a_n1246_n2088# 0.014062f
C107 source.n39 a_n1246_n2088# 0.024716f
C108 source.n40 a_n1246_n2088# 0.013281f
C109 source.n41 a_n1246_n2088# 0.031392f
C110 source.n42 a_n1246_n2088# 0.014062f
C111 source.n43 a_n1246_n2088# 0.105766f
C112 source.t4 a_n1246_n2088# 0.051165f
C113 source.n44 a_n1246_n2088# 0.023544f
C114 source.n45 a_n1246_n2088# 0.018543f
C115 source.n46 a_n1246_n2088# 0.013281f
C116 source.n47 a_n1246_n2088# 0.588087f
C117 source.n48 a_n1246_n2088# 0.024716f
C118 source.n49 a_n1246_n2088# 0.013281f
C119 source.n50 a_n1246_n2088# 0.014062f
C120 source.n51 a_n1246_n2088# 0.031392f
C121 source.n52 a_n1246_n2088# 0.031392f
C122 source.n53 a_n1246_n2088# 0.014062f
C123 source.n54 a_n1246_n2088# 0.013281f
C124 source.n55 a_n1246_n2088# 0.024716f
C125 source.n56 a_n1246_n2088# 0.024716f
C126 source.n57 a_n1246_n2088# 0.013281f
C127 source.n58 a_n1246_n2088# 0.014062f
C128 source.n59 a_n1246_n2088# 0.031392f
C129 source.n60 a_n1246_n2088# 0.067958f
C130 source.n61 a_n1246_n2088# 0.014062f
C131 source.n62 a_n1246_n2088# 0.013281f
C132 source.n63 a_n1246_n2088# 0.057129f
C133 source.n64 a_n1246_n2088# 0.038025f
C134 source.n65 a_n1246_n2088# 0.094913f
C135 source.n66 a_n1246_n2088# 0.03474f
C136 source.n67 a_n1246_n2088# 0.024716f
C137 source.n68 a_n1246_n2088# 0.013281f
C138 source.n69 a_n1246_n2088# 0.031392f
C139 source.n70 a_n1246_n2088# 0.014062f
C140 source.n71 a_n1246_n2088# 0.024716f
C141 source.n72 a_n1246_n2088# 0.013281f
C142 source.n73 a_n1246_n2088# 0.031392f
C143 source.n74 a_n1246_n2088# 0.014062f
C144 source.n75 a_n1246_n2088# 0.105766f
C145 source.t6 a_n1246_n2088# 0.051165f
C146 source.n76 a_n1246_n2088# 0.023544f
C147 source.n77 a_n1246_n2088# 0.018543f
C148 source.n78 a_n1246_n2088# 0.013281f
C149 source.n79 a_n1246_n2088# 0.588087f
C150 source.n80 a_n1246_n2088# 0.024716f
C151 source.n81 a_n1246_n2088# 0.013281f
C152 source.n82 a_n1246_n2088# 0.014062f
C153 source.n83 a_n1246_n2088# 0.031392f
C154 source.n84 a_n1246_n2088# 0.031392f
C155 source.n85 a_n1246_n2088# 0.014062f
C156 source.n86 a_n1246_n2088# 0.013281f
C157 source.n87 a_n1246_n2088# 0.024716f
C158 source.n88 a_n1246_n2088# 0.024716f
C159 source.n89 a_n1246_n2088# 0.013281f
C160 source.n90 a_n1246_n2088# 0.014062f
C161 source.n91 a_n1246_n2088# 0.031392f
C162 source.n92 a_n1246_n2088# 0.067958f
C163 source.n93 a_n1246_n2088# 0.014062f
C164 source.n94 a_n1246_n2088# 0.013281f
C165 source.n95 a_n1246_n2088# 0.057129f
C166 source.n96 a_n1246_n2088# 0.038025f
C167 source.n97 a_n1246_n2088# 0.094913f
C168 source.t10 a_n1246_n2088# 0.117187f
C169 source.t11 a_n1246_n2088# 0.117187f
C170 source.n98 a_n1246_n2088# 0.91266f
C171 source.n99 a_n1246_n2088# 0.304461f
C172 source.n100 a_n1246_n2088# 0.03474f
C173 source.n101 a_n1246_n2088# 0.024716f
C174 source.n102 a_n1246_n2088# 0.013281f
C175 source.n103 a_n1246_n2088# 0.031392f
C176 source.n104 a_n1246_n2088# 0.014062f
C177 source.n105 a_n1246_n2088# 0.024716f
C178 source.n106 a_n1246_n2088# 0.013281f
C179 source.n107 a_n1246_n2088# 0.031392f
C180 source.n108 a_n1246_n2088# 0.014062f
C181 source.n109 a_n1246_n2088# 0.105766f
C182 source.t7 a_n1246_n2088# 0.051165f
C183 source.n110 a_n1246_n2088# 0.023544f
C184 source.n111 a_n1246_n2088# 0.018543f
C185 source.n112 a_n1246_n2088# 0.013281f
C186 source.n113 a_n1246_n2088# 0.588087f
C187 source.n114 a_n1246_n2088# 0.024716f
C188 source.n115 a_n1246_n2088# 0.013281f
C189 source.n116 a_n1246_n2088# 0.014062f
C190 source.n117 a_n1246_n2088# 0.031392f
C191 source.n118 a_n1246_n2088# 0.031392f
C192 source.n119 a_n1246_n2088# 0.014062f
C193 source.n120 a_n1246_n2088# 0.013281f
C194 source.n121 a_n1246_n2088# 0.024716f
C195 source.n122 a_n1246_n2088# 0.024716f
C196 source.n123 a_n1246_n2088# 0.013281f
C197 source.n124 a_n1246_n2088# 0.014062f
C198 source.n125 a_n1246_n2088# 0.031392f
C199 source.n126 a_n1246_n2088# 0.067958f
C200 source.n127 a_n1246_n2088# 0.014062f
C201 source.n128 a_n1246_n2088# 0.013281f
C202 source.n129 a_n1246_n2088# 0.057129f
C203 source.n130 a_n1246_n2088# 0.038025f
C204 source.n131 a_n1246_n2088# 0.903123f
C205 source.n132 a_n1246_n2088# 0.03474f
C206 source.n133 a_n1246_n2088# 0.024716f
C207 source.n134 a_n1246_n2088# 0.013281f
C208 source.n135 a_n1246_n2088# 0.031392f
C209 source.n136 a_n1246_n2088# 0.014062f
C210 source.n137 a_n1246_n2088# 0.024716f
C211 source.n138 a_n1246_n2088# 0.013281f
C212 source.n139 a_n1246_n2088# 0.031392f
C213 source.n140 a_n1246_n2088# 0.014062f
C214 source.n141 a_n1246_n2088# 0.105766f
C215 source.t14 a_n1246_n2088# 0.051165f
C216 source.n142 a_n1246_n2088# 0.023544f
C217 source.n143 a_n1246_n2088# 0.018543f
C218 source.n144 a_n1246_n2088# 0.013281f
C219 source.n145 a_n1246_n2088# 0.588087f
C220 source.n146 a_n1246_n2088# 0.024716f
C221 source.n147 a_n1246_n2088# 0.013281f
C222 source.n148 a_n1246_n2088# 0.014062f
C223 source.n149 a_n1246_n2088# 0.031392f
C224 source.n150 a_n1246_n2088# 0.031392f
C225 source.n151 a_n1246_n2088# 0.014062f
C226 source.n152 a_n1246_n2088# 0.013281f
C227 source.n153 a_n1246_n2088# 0.024716f
C228 source.n154 a_n1246_n2088# 0.024716f
C229 source.n155 a_n1246_n2088# 0.013281f
C230 source.n156 a_n1246_n2088# 0.014062f
C231 source.n157 a_n1246_n2088# 0.031392f
C232 source.n158 a_n1246_n2088# 0.067958f
C233 source.n159 a_n1246_n2088# 0.014062f
C234 source.n160 a_n1246_n2088# 0.013281f
C235 source.n161 a_n1246_n2088# 0.057129f
C236 source.n162 a_n1246_n2088# 0.038025f
C237 source.n163 a_n1246_n2088# 0.903123f
C238 source.t0 a_n1246_n2088# 0.117187f
C239 source.t2 a_n1246_n2088# 0.117187f
C240 source.n164 a_n1246_n2088# 0.912654f
C241 source.n165 a_n1246_n2088# 0.304467f
C242 source.n166 a_n1246_n2088# 0.03474f
C243 source.n167 a_n1246_n2088# 0.024716f
C244 source.n168 a_n1246_n2088# 0.013281f
C245 source.n169 a_n1246_n2088# 0.031392f
C246 source.n170 a_n1246_n2088# 0.014062f
C247 source.n171 a_n1246_n2088# 0.024716f
C248 source.n172 a_n1246_n2088# 0.013281f
C249 source.n173 a_n1246_n2088# 0.031392f
C250 source.n174 a_n1246_n2088# 0.014062f
C251 source.n175 a_n1246_n2088# 0.105766f
C252 source.t15 a_n1246_n2088# 0.051165f
C253 source.n176 a_n1246_n2088# 0.023544f
C254 source.n177 a_n1246_n2088# 0.018543f
C255 source.n178 a_n1246_n2088# 0.013281f
C256 source.n179 a_n1246_n2088# 0.588087f
C257 source.n180 a_n1246_n2088# 0.024716f
C258 source.n181 a_n1246_n2088# 0.013281f
C259 source.n182 a_n1246_n2088# 0.014062f
C260 source.n183 a_n1246_n2088# 0.031392f
C261 source.n184 a_n1246_n2088# 0.031392f
C262 source.n185 a_n1246_n2088# 0.014062f
C263 source.n186 a_n1246_n2088# 0.013281f
C264 source.n187 a_n1246_n2088# 0.024716f
C265 source.n188 a_n1246_n2088# 0.024716f
C266 source.n189 a_n1246_n2088# 0.013281f
C267 source.n190 a_n1246_n2088# 0.014062f
C268 source.n191 a_n1246_n2088# 0.031392f
C269 source.n192 a_n1246_n2088# 0.067958f
C270 source.n193 a_n1246_n2088# 0.014062f
C271 source.n194 a_n1246_n2088# 0.013281f
C272 source.n195 a_n1246_n2088# 0.057129f
C273 source.n196 a_n1246_n2088# 0.038025f
C274 source.n197 a_n1246_n2088# 0.094913f
C275 source.n198 a_n1246_n2088# 0.03474f
C276 source.n199 a_n1246_n2088# 0.024716f
C277 source.n200 a_n1246_n2088# 0.013281f
C278 source.n201 a_n1246_n2088# 0.031392f
C279 source.n202 a_n1246_n2088# 0.014062f
C280 source.n203 a_n1246_n2088# 0.024716f
C281 source.n204 a_n1246_n2088# 0.013281f
C282 source.n205 a_n1246_n2088# 0.031392f
C283 source.n206 a_n1246_n2088# 0.014062f
C284 source.n207 a_n1246_n2088# 0.105766f
C285 source.t13 a_n1246_n2088# 0.051165f
C286 source.n208 a_n1246_n2088# 0.023544f
C287 source.n209 a_n1246_n2088# 0.018543f
C288 source.n210 a_n1246_n2088# 0.013281f
C289 source.n211 a_n1246_n2088# 0.588087f
C290 source.n212 a_n1246_n2088# 0.024716f
C291 source.n213 a_n1246_n2088# 0.013281f
C292 source.n214 a_n1246_n2088# 0.014062f
C293 source.n215 a_n1246_n2088# 0.031392f
C294 source.n216 a_n1246_n2088# 0.031392f
C295 source.n217 a_n1246_n2088# 0.014062f
C296 source.n218 a_n1246_n2088# 0.013281f
C297 source.n219 a_n1246_n2088# 0.024716f
C298 source.n220 a_n1246_n2088# 0.024716f
C299 source.n221 a_n1246_n2088# 0.013281f
C300 source.n222 a_n1246_n2088# 0.014062f
C301 source.n223 a_n1246_n2088# 0.031392f
C302 source.n224 a_n1246_n2088# 0.067958f
C303 source.n225 a_n1246_n2088# 0.014062f
C304 source.n226 a_n1246_n2088# 0.013281f
C305 source.n227 a_n1246_n2088# 0.057129f
C306 source.n228 a_n1246_n2088# 0.038025f
C307 source.n229 a_n1246_n2088# 0.094913f
C308 source.t9 a_n1246_n2088# 0.117187f
C309 source.t12 a_n1246_n2088# 0.117187f
C310 source.n230 a_n1246_n2088# 0.912654f
C311 source.n231 a_n1246_n2088# 0.304467f
C312 source.n232 a_n1246_n2088# 0.03474f
C313 source.n233 a_n1246_n2088# 0.024716f
C314 source.n234 a_n1246_n2088# 0.013281f
C315 source.n235 a_n1246_n2088# 0.031392f
C316 source.n236 a_n1246_n2088# 0.014062f
C317 source.n237 a_n1246_n2088# 0.024716f
C318 source.n238 a_n1246_n2088# 0.013281f
C319 source.n239 a_n1246_n2088# 0.031392f
C320 source.n240 a_n1246_n2088# 0.014062f
C321 source.n241 a_n1246_n2088# 0.105766f
C322 source.t8 a_n1246_n2088# 0.051165f
C323 source.n242 a_n1246_n2088# 0.023544f
C324 source.n243 a_n1246_n2088# 0.018543f
C325 source.n244 a_n1246_n2088# 0.013281f
C326 source.n245 a_n1246_n2088# 0.588087f
C327 source.n246 a_n1246_n2088# 0.024716f
C328 source.n247 a_n1246_n2088# 0.013281f
C329 source.n248 a_n1246_n2088# 0.014062f
C330 source.n249 a_n1246_n2088# 0.031392f
C331 source.n250 a_n1246_n2088# 0.031392f
C332 source.n251 a_n1246_n2088# 0.014062f
C333 source.n252 a_n1246_n2088# 0.013281f
C334 source.n253 a_n1246_n2088# 0.024716f
C335 source.n254 a_n1246_n2088# 0.024716f
C336 source.n255 a_n1246_n2088# 0.013281f
C337 source.n256 a_n1246_n2088# 0.014062f
C338 source.n257 a_n1246_n2088# 0.031392f
C339 source.n258 a_n1246_n2088# 0.067958f
C340 source.n259 a_n1246_n2088# 0.014062f
C341 source.n260 a_n1246_n2088# 0.013281f
C342 source.n261 a_n1246_n2088# 0.057129f
C343 source.n262 a_n1246_n2088# 0.038025f
C344 source.n263 a_n1246_n2088# 0.22893f
C345 source.n264 a_n1246_n2088# 1.00801f
C346 minus.n0 a_n1246_n2088# 0.071379f
C347 minus.t5 a_n1246_n2088# 0.114636f
C348 minus.t0 a_n1246_n2088# 0.112081f
C349 minus.t1 a_n1246_n2088# 0.112081f
C350 minus.t2 a_n1246_n2088# 0.114636f
C351 minus.n1 a_n1246_n2088# 0.063686f
C352 minus.n2 a_n1246_n2088# 0.054815f
C353 minus.n3 a_n1246_n2088# 0.011481f
C354 minus.n4 a_n1246_n2088# 0.054815f
C355 minus.n5 a_n1246_n2088# 0.063641f
C356 minus.n6 a_n1246_n2088# 0.81419f
C357 minus.n7 a_n1246_n2088# 0.071379f
C358 minus.t3 a_n1246_n2088# 0.112081f
C359 minus.t7 a_n1246_n2088# 0.112081f
C360 minus.t4 a_n1246_n2088# 0.114636f
C361 minus.n8 a_n1246_n2088# 0.063686f
C362 minus.n9 a_n1246_n2088# 0.054815f
C363 minus.n10 a_n1246_n2088# 0.011481f
C364 minus.n11 a_n1246_n2088# 0.054815f
C365 minus.t6 a_n1246_n2088# 0.114636f
C366 minus.n12 a_n1246_n2088# 0.063641f
C367 minus.n13 a_n1246_n2088# 0.209957f
C368 minus.n14 a_n1246_n2088# 1.00782f
.ends

