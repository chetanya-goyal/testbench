* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t28 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X1 drain_right.t19 minus.t0 source.t14 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X2 a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X3 source.t15 minus.t1 drain_right.t18 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 drain_right.t17 minus.t2 source.t36 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X5 source.t16 plus.t1 drain_left.t18 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X6 source.t17 plus.t2 drain_left.t17 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 source.t26 plus.t3 drain_left.t16 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X8 source.t39 minus.t3 drain_right.t16 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X9 drain_right.t15 minus.t4 source.t37 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 source.t18 plus.t4 drain_left.t15 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 drain_right.t14 minus.t5 source.t12 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 drain_right.t13 minus.t6 source.t10 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 source.t9 minus.t7 drain_right.t12 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X15 a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X16 drain_left.t14 plus.t5 source.t24 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 drain_left.t13 plus.t6 source.t27 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 source.t11 minus.t8 drain_right.t11 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X19 source.t20 plus.t7 drain_left.t12 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X20 source.t38 minus.t9 drain_right.t10 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X21 drain_right.t9 minus.t10 source.t13 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 source.t8 minus.t11 drain_right.t8 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 drain_left.t11 plus.t8 source.t19 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X24 drain_left.t10 plus.t9 source.t21 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X25 drain_right.t7 minus.t12 source.t6 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X26 drain_right.t6 minus.t13 source.t7 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 drain_right.t5 minus.t14 source.t1 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X28 drain_left.t9 plus.t10 source.t31 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 drain_right.t4 minus.t15 source.t3 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 source.t5 minus.t16 drain_right.t3 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 source.t35 plus.t11 drain_left.t8 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X32 source.t30 plus.t12 drain_left.t7 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X33 source.t4 minus.t17 drain_right.t2 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X34 source.t32 plus.t13 drain_left.t6 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X35 source.t25 plus.t14 drain_left.t5 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X36 source.t0 minus.t18 drain_right.t1 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X37 drain_left.t4 plus.t15 source.t34 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X38 drain_left.t3 plus.t16 source.t29 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X39 source.t23 plus.t17 drain_left.t2 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X40 a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X41 source.t2 minus.t19 drain_right.t0 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X42 drain_left.t1 plus.t18 source.t22 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X43 drain_left.t0 plus.t19 source.t33 a_n2542_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
R0 plus.n10 plus.n9 161.3
R1 plus.n11 plus.n6 161.3
R2 plus.n12 plus.n5 161.3
R3 plus.n14 plus.n13 161.3
R4 plus.n15 plus.n4 161.3
R5 plus.n17 plus.n16 161.3
R6 plus.n18 plus.n3 161.3
R7 plus.n19 plus.n2 161.3
R8 plus.n21 plus.n20 161.3
R9 plus.n22 plus.n1 161.3
R10 plus.n24 plus.n23 161.3
R11 plus.n25 plus.n0 161.3
R12 plus.n27 plus.n26 161.3
R13 plus.n38 plus.n37 161.3
R14 plus.n39 plus.n34 161.3
R15 plus.n40 plus.n33 161.3
R16 plus.n42 plus.n41 161.3
R17 plus.n43 plus.n32 161.3
R18 plus.n45 plus.n44 161.3
R19 plus.n46 plus.n31 161.3
R20 plus.n47 plus.n30 161.3
R21 plus.n49 plus.n48 161.3
R22 plus.n50 plus.n29 161.3
R23 plus.n52 plus.n51 161.3
R24 plus.n53 plus.n28 161.3
R25 plus.n55 plus.n54 161.3
R26 plus.n8 plus.t3 147.749
R27 plus.n36 plus.t8 147.749
R28 plus.n26 plus.t9 126.766
R29 plus.n25 plus.t2 126.766
R30 plus.n1 plus.t16 126.766
R31 plus.n19 plus.t7 126.766
R32 plus.n18 plus.t19 126.766
R33 plus.n4 plus.t14 126.766
R34 plus.n13 plus.t5 126.766
R35 plus.n11 plus.t17 126.766
R36 plus.n7 plus.t10 126.766
R37 plus.n54 plus.t1 126.766
R38 plus.n53 plus.t18 126.766
R39 plus.n29 plus.t4 126.766
R40 plus.n47 plus.t15 126.766
R41 plus.n46 plus.t12 126.766
R42 plus.n32 plus.t0 126.766
R43 plus.n41 plus.t13 126.766
R44 plus.n39 plus.t6 126.766
R45 plus.n35 plus.t11 126.766
R46 plus.n9 plus.n8 70.4033
R47 plus.n37 plus.n36 70.4033
R48 plus.n26 plus.n25 48.2005
R49 plus.n19 plus.n18 48.2005
R50 plus.n13 plus.n4 48.2005
R51 plus.n54 plus.n53 48.2005
R52 plus.n47 plus.n46 48.2005
R53 plus.n41 plus.n32 48.2005
R54 plus.n20 plus.n1 47.4702
R55 plus.n12 plus.n11 47.4702
R56 plus.n48 plus.n29 47.4702
R57 plus.n40 plus.n39 47.4702
R58 plus plus.n55 28.5558
R59 plus.n24 plus.n1 25.5611
R60 plus.n11 plus.n10 25.5611
R61 plus.n52 plus.n29 25.5611
R62 plus.n39 plus.n38 25.5611
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n25 plus.n24 22.6399
R68 plus.n10 plus.n7 22.6399
R69 plus.n53 plus.n52 22.6399
R70 plus.n38 plus.n35 22.6399
R71 plus.n8 plus.n7 20.9576
R72 plus.n36 plus.n35 20.9576
R73 plus plus.n27 8.06868
R74 plus.n20 plus.n19 0.730803
R75 plus.n13 plus.n12 0.730803
R76 plus.n48 plus.n47 0.730803
R77 plus.n41 plus.n40 0.730803
R78 plus.n9 plus.n6 0.189894
R79 plus.n6 plus.n5 0.189894
R80 plus.n14 plus.n5 0.189894
R81 plus.n15 plus.n14 0.189894
R82 plus.n16 plus.n15 0.189894
R83 plus.n16 plus.n3 0.189894
R84 plus.n3 plus.n2 0.189894
R85 plus.n21 plus.n2 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n23 plus.n22 0.189894
R88 plus.n23 plus.n0 0.189894
R89 plus.n27 plus.n0 0.189894
R90 plus.n55 plus.n28 0.189894
R91 plus.n51 plus.n28 0.189894
R92 plus.n51 plus.n50 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n30 0.189894
R95 plus.n31 plus.n30 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n34 plus.n33 0.189894
R101 plus.n37 plus.n34 0.189894
R102 source.n0 source.t21 243.255
R103 source.n9 source.t26 243.255
R104 source.n10 source.t6 243.255
R105 source.n19 source.t39 243.255
R106 source.n39 source.t36 243.254
R107 source.n30 source.t11 243.254
R108 source.n29 source.t19 243.254
R109 source.n20 source.t16 243.254
R110 source.n2 source.n1 223.454
R111 source.n4 source.n3 223.454
R112 source.n6 source.n5 223.454
R113 source.n8 source.n7 223.454
R114 source.n12 source.n11 223.454
R115 source.n14 source.n13 223.454
R116 source.n16 source.n15 223.454
R117 source.n18 source.n17 223.454
R118 source.n38 source.n37 223.453
R119 source.n36 source.n35 223.453
R120 source.n34 source.n33 223.453
R121 source.n32 source.n31 223.453
R122 source.n28 source.n27 223.453
R123 source.n26 source.n25 223.453
R124 source.n24 source.n23 223.453
R125 source.n22 source.n21 223.453
R126 source.n37 source.t12 19.8005
R127 source.n37 source.t5 19.8005
R128 source.n35 source.t1 19.8005
R129 source.n35 source.t0 19.8005
R130 source.n33 source.t13 19.8005
R131 source.n33 source.t2 19.8005
R132 source.n31 source.t7 19.8005
R133 source.n31 source.t9 19.8005
R134 source.n27 source.t27 19.8005
R135 source.n27 source.t35 19.8005
R136 source.n25 source.t28 19.8005
R137 source.n25 source.t32 19.8005
R138 source.n23 source.t34 19.8005
R139 source.n23 source.t30 19.8005
R140 source.n21 source.t22 19.8005
R141 source.n21 source.t18 19.8005
R142 source.n1 source.t29 19.8005
R143 source.n1 source.t17 19.8005
R144 source.n3 source.t33 19.8005
R145 source.n3 source.t20 19.8005
R146 source.n5 source.t24 19.8005
R147 source.n5 source.t25 19.8005
R148 source.n7 source.t31 19.8005
R149 source.n7 source.t23 19.8005
R150 source.n11 source.t10 19.8005
R151 source.n11 source.t15 19.8005
R152 source.n13 source.t37 19.8005
R153 source.n13 source.t4 19.8005
R154 source.n15 source.t14 19.8005
R155 source.n15 source.t38 19.8005
R156 source.n17 source.t3 19.8005
R157 source.n17 source.t8 19.8005
R158 source.n20 source.n19 13.6699
R159 source.n40 source.n0 8.04922
R160 source.n40 source.n39 5.62119
R161 source.n19 source.n18 0.716017
R162 source.n18 source.n16 0.716017
R163 source.n16 source.n14 0.716017
R164 source.n14 source.n12 0.716017
R165 source.n12 source.n10 0.716017
R166 source.n9 source.n8 0.716017
R167 source.n8 source.n6 0.716017
R168 source.n6 source.n4 0.716017
R169 source.n4 source.n2 0.716017
R170 source.n2 source.n0 0.716017
R171 source.n22 source.n20 0.716017
R172 source.n24 source.n22 0.716017
R173 source.n26 source.n24 0.716017
R174 source.n28 source.n26 0.716017
R175 source.n29 source.n28 0.716017
R176 source.n32 source.n30 0.716017
R177 source.n34 source.n32 0.716017
R178 source.n36 source.n34 0.716017
R179 source.n38 source.n36 0.716017
R180 source.n39 source.n38 0.716017
R181 source.n10 source.n9 0.470328
R182 source.n30 source.n29 0.470328
R183 source source.n40 0.188
R184 drain_left.n10 drain_left.n8 240.849
R185 drain_left.n6 drain_left.n4 240.847
R186 drain_left.n2 drain_left.n0 240.847
R187 drain_left.n16 drain_left.n15 240.132
R188 drain_left.n14 drain_left.n13 240.132
R189 drain_left.n12 drain_left.n11 240.132
R190 drain_left.n10 drain_left.n9 240.132
R191 drain_left.n7 drain_left.n3 240.131
R192 drain_left.n6 drain_left.n5 240.131
R193 drain_left.n2 drain_left.n1 240.131
R194 drain_left drain_left.n7 24.7579
R195 drain_left.n3 drain_left.t7 19.8005
R196 drain_left.n3 drain_left.t19 19.8005
R197 drain_left.n4 drain_left.t8 19.8005
R198 drain_left.n4 drain_left.t11 19.8005
R199 drain_left.n5 drain_left.t6 19.8005
R200 drain_left.n5 drain_left.t13 19.8005
R201 drain_left.n1 drain_left.t15 19.8005
R202 drain_left.n1 drain_left.t4 19.8005
R203 drain_left.n0 drain_left.t18 19.8005
R204 drain_left.n0 drain_left.t1 19.8005
R205 drain_left.n15 drain_left.t17 19.8005
R206 drain_left.n15 drain_left.t10 19.8005
R207 drain_left.n13 drain_left.t12 19.8005
R208 drain_left.n13 drain_left.t3 19.8005
R209 drain_left.n11 drain_left.t5 19.8005
R210 drain_left.n11 drain_left.t0 19.8005
R211 drain_left.n9 drain_left.t2 19.8005
R212 drain_left.n9 drain_left.t14 19.8005
R213 drain_left.n8 drain_left.t16 19.8005
R214 drain_left.n8 drain_left.t9 19.8005
R215 drain_left drain_left.n16 6.36873
R216 drain_left.n12 drain_left.n10 0.716017
R217 drain_left.n14 drain_left.n12 0.716017
R218 drain_left.n16 drain_left.n14 0.716017
R219 drain_left.n7 drain_left.n6 0.660671
R220 drain_left.n7 drain_left.n2 0.660671
R221 minus.n27 minus.n26 161.3
R222 minus.n25 minus.n0 161.3
R223 minus.n24 minus.n23 161.3
R224 minus.n22 minus.n1 161.3
R225 minus.n21 minus.n20 161.3
R226 minus.n19 minus.n2 161.3
R227 minus.n18 minus.n17 161.3
R228 minus.n16 minus.n3 161.3
R229 minus.n15 minus.n14 161.3
R230 minus.n13 minus.n4 161.3
R231 minus.n12 minus.n11 161.3
R232 minus.n10 minus.n5 161.3
R233 minus.n9 minus.n8 161.3
R234 minus.n55 minus.n54 161.3
R235 minus.n53 minus.n28 161.3
R236 minus.n52 minus.n51 161.3
R237 minus.n50 minus.n29 161.3
R238 minus.n49 minus.n48 161.3
R239 minus.n47 minus.n30 161.3
R240 minus.n46 minus.n45 161.3
R241 minus.n44 minus.n31 161.3
R242 minus.n43 minus.n42 161.3
R243 minus.n41 minus.n32 161.3
R244 minus.n40 minus.n39 161.3
R245 minus.n38 minus.n33 161.3
R246 minus.n37 minus.n36 161.3
R247 minus.n6 minus.t12 147.749
R248 minus.n34 minus.t8 147.749
R249 minus.n7 minus.t1 126.766
R250 minus.n5 minus.t6 126.766
R251 minus.n13 minus.t17 126.766
R252 minus.n14 minus.t4 126.766
R253 minus.n18 minus.t9 126.766
R254 minus.n19 minus.t0 126.766
R255 minus.n1 minus.t11 126.766
R256 minus.n25 minus.t15 126.766
R257 minus.n26 minus.t3 126.766
R258 minus.n35 minus.t13 126.766
R259 minus.n33 minus.t7 126.766
R260 minus.n41 minus.t10 126.766
R261 minus.n42 minus.t19 126.766
R262 minus.n46 minus.t14 126.766
R263 minus.n47 minus.t18 126.766
R264 minus.n29 minus.t5 126.766
R265 minus.n53 minus.t16 126.766
R266 minus.n54 minus.t2 126.766
R267 minus.n9 minus.n6 70.4033
R268 minus.n37 minus.n34 70.4033
R269 minus.n14 minus.n13 48.2005
R270 minus.n19 minus.n18 48.2005
R271 minus.n26 minus.n25 48.2005
R272 minus.n42 minus.n41 48.2005
R273 minus.n47 minus.n46 48.2005
R274 minus.n54 minus.n53 48.2005
R275 minus.n12 minus.n5 47.4702
R276 minus.n20 minus.n1 47.4702
R277 minus.n40 minus.n33 47.4702
R278 minus.n48 minus.n29 47.4702
R279 minus.n56 minus.n27 30.5081
R280 minus.n8 minus.n5 25.5611
R281 minus.n24 minus.n1 25.5611
R282 minus.n36 minus.n33 25.5611
R283 minus.n52 minus.n29 25.5611
R284 minus.n18 minus.n3 24.1005
R285 minus.n14 minus.n3 24.1005
R286 minus.n42 minus.n31 24.1005
R287 minus.n46 minus.n31 24.1005
R288 minus.n8 minus.n7 22.6399
R289 minus.n25 minus.n24 22.6399
R290 minus.n36 minus.n35 22.6399
R291 minus.n53 minus.n52 22.6399
R292 minus.n7 minus.n6 20.9576
R293 minus.n35 minus.n34 20.9576
R294 minus.n56 minus.n55 6.59141
R295 minus.n13 minus.n12 0.730803
R296 minus.n20 minus.n19 0.730803
R297 minus.n41 minus.n40 0.730803
R298 minus.n48 minus.n47 0.730803
R299 minus.n27 minus.n0 0.189894
R300 minus.n23 minus.n0 0.189894
R301 minus.n23 minus.n22 0.189894
R302 minus.n22 minus.n21 0.189894
R303 minus.n21 minus.n2 0.189894
R304 minus.n17 minus.n2 0.189894
R305 minus.n17 minus.n16 0.189894
R306 minus.n16 minus.n15 0.189894
R307 minus.n15 minus.n4 0.189894
R308 minus.n11 minus.n4 0.189894
R309 minus.n11 minus.n10 0.189894
R310 minus.n10 minus.n9 0.189894
R311 minus.n38 minus.n37 0.189894
R312 minus.n39 minus.n38 0.189894
R313 minus.n39 minus.n32 0.189894
R314 minus.n43 minus.n32 0.189894
R315 minus.n44 minus.n43 0.189894
R316 minus.n45 minus.n44 0.189894
R317 minus.n45 minus.n30 0.189894
R318 minus.n49 minus.n30 0.189894
R319 minus.n50 minus.n49 0.189894
R320 minus.n51 minus.n50 0.189894
R321 minus.n51 minus.n28 0.189894
R322 minus.n55 minus.n28 0.189894
R323 minus minus.n56 0.188
R324 drain_right.n10 drain_right.n8 240.849
R325 drain_right.n6 drain_right.n4 240.847
R326 drain_right.n2 drain_right.n0 240.847
R327 drain_right.n10 drain_right.n9 240.132
R328 drain_right.n12 drain_right.n11 240.132
R329 drain_right.n14 drain_right.n13 240.132
R330 drain_right.n16 drain_right.n15 240.132
R331 drain_right.n7 drain_right.n3 240.131
R332 drain_right.n6 drain_right.n5 240.131
R333 drain_right.n2 drain_right.n1 240.131
R334 drain_right drain_right.n7 24.2047
R335 drain_right.n3 drain_right.t0 19.8005
R336 drain_right.n3 drain_right.t5 19.8005
R337 drain_right.n4 drain_right.t3 19.8005
R338 drain_right.n4 drain_right.t17 19.8005
R339 drain_right.n5 drain_right.t1 19.8005
R340 drain_right.n5 drain_right.t14 19.8005
R341 drain_right.n1 drain_right.t12 19.8005
R342 drain_right.n1 drain_right.t9 19.8005
R343 drain_right.n0 drain_right.t11 19.8005
R344 drain_right.n0 drain_right.t6 19.8005
R345 drain_right.n8 drain_right.t18 19.8005
R346 drain_right.n8 drain_right.t7 19.8005
R347 drain_right.n9 drain_right.t2 19.8005
R348 drain_right.n9 drain_right.t13 19.8005
R349 drain_right.n11 drain_right.t10 19.8005
R350 drain_right.n11 drain_right.t15 19.8005
R351 drain_right.n13 drain_right.t8 19.8005
R352 drain_right.n13 drain_right.t19 19.8005
R353 drain_right.n15 drain_right.t16 19.8005
R354 drain_right.n15 drain_right.t4 19.8005
R355 drain_right drain_right.n16 6.36873
R356 drain_right.n16 drain_right.n14 0.716017
R357 drain_right.n14 drain_right.n12 0.716017
R358 drain_right.n12 drain_right.n10 0.716017
R359 drain_right.n7 drain_right.n6 0.660671
R360 drain_right.n7 drain_right.n2 0.660671
C0 drain_right plus 0.416967f
C1 drain_right drain_left 1.35905f
C2 drain_right source 5.76694f
C3 plus minus 4.29277f
C4 minus drain_left 0.180519f
C5 minus source 2.05893f
C6 plus drain_left 1.69542f
C7 plus source 2.0728f
C8 source drain_left 5.76563f
C9 drain_right minus 1.44385f
C10 drain_right a_n2542_n1088# 4.41064f
C11 drain_left a_n2542_n1088# 4.737741f
C12 source a_n2542_n1088# 2.782396f
C13 minus a_n2542_n1088# 9.20787f
C14 plus a_n2542_n1088# 10.228951f
C15 drain_right.t11 a_n2542_n1088# 0.017691f
C16 drain_right.t6 a_n2542_n1088# 0.017691f
C17 drain_right.n0 a_n2542_n1088# 0.069541f
C18 drain_right.t12 a_n2542_n1088# 0.017691f
C19 drain_right.t9 a_n2542_n1088# 0.017691f
C20 drain_right.n1 a_n2542_n1088# 0.068743f
C21 drain_right.n2 a_n2542_n1088# 0.524588f
C22 drain_right.t0 a_n2542_n1088# 0.017691f
C23 drain_right.t5 a_n2542_n1088# 0.017691f
C24 drain_right.n3 a_n2542_n1088# 0.068743f
C25 drain_right.t3 a_n2542_n1088# 0.017691f
C26 drain_right.t17 a_n2542_n1088# 0.017691f
C27 drain_right.n4 a_n2542_n1088# 0.069541f
C28 drain_right.t1 a_n2542_n1088# 0.017691f
C29 drain_right.t14 a_n2542_n1088# 0.017691f
C30 drain_right.n5 a_n2542_n1088# 0.068743f
C31 drain_right.n6 a_n2542_n1088# 0.524588f
C32 drain_right.n7 a_n2542_n1088# 0.932139f
C33 drain_right.t18 a_n2542_n1088# 0.017691f
C34 drain_right.t7 a_n2542_n1088# 0.017691f
C35 drain_right.n8 a_n2542_n1088# 0.069541f
C36 drain_right.t2 a_n2542_n1088# 0.017691f
C37 drain_right.t13 a_n2542_n1088# 0.017691f
C38 drain_right.n9 a_n2542_n1088# 0.068743f
C39 drain_right.n10 a_n2542_n1088# 0.527794f
C40 drain_right.t10 a_n2542_n1088# 0.017691f
C41 drain_right.t15 a_n2542_n1088# 0.017691f
C42 drain_right.n11 a_n2542_n1088# 0.068743f
C43 drain_right.n12 a_n2542_n1088# 0.259788f
C44 drain_right.t8 a_n2542_n1088# 0.017691f
C45 drain_right.t19 a_n2542_n1088# 0.017691f
C46 drain_right.n13 a_n2542_n1088# 0.068743f
C47 drain_right.n14 a_n2542_n1088# 0.259788f
C48 drain_right.t16 a_n2542_n1088# 0.017691f
C49 drain_right.t4 a_n2542_n1088# 0.017691f
C50 drain_right.n15 a_n2542_n1088# 0.068743f
C51 drain_right.n16 a_n2542_n1088# 0.452126f
C52 minus.n0 a_n2542_n1088# 0.037981f
C53 minus.t11 a_n2542_n1088# 0.064397f
C54 minus.n1 a_n2542_n1088# 0.070965f
C55 minus.n2 a_n2542_n1088# 0.037981f
C56 minus.n3 a_n2542_n1088# 0.008619f
C57 minus.t9 a_n2542_n1088# 0.064397f
C58 minus.n4 a_n2542_n1088# 0.037981f
C59 minus.t6 a_n2542_n1088# 0.064397f
C60 minus.n5 a_n2542_n1088# 0.070965f
C61 minus.t12 a_n2542_n1088# 0.073917f
C62 minus.n6 a_n2542_n1088# 0.057754f
C63 minus.t1 a_n2542_n1088# 0.064397f
C64 minus.n7 a_n2542_n1088# 0.070613f
C65 minus.n8 a_n2542_n1088# 0.008619f
C66 minus.n9 a_n2542_n1088# 0.124658f
C67 minus.n10 a_n2542_n1088# 0.037981f
C68 minus.n11 a_n2542_n1088# 0.037981f
C69 minus.n12 a_n2542_n1088# 0.008619f
C70 minus.t17 a_n2542_n1088# 0.064397f
C71 minus.n13 a_n2542_n1088# 0.067101f
C72 minus.t4 a_n2542_n1088# 0.064397f
C73 minus.n14 a_n2542_n1088# 0.070848f
C74 minus.n15 a_n2542_n1088# 0.037981f
C75 minus.n16 a_n2542_n1088# 0.037981f
C76 minus.n17 a_n2542_n1088# 0.037981f
C77 minus.n18 a_n2542_n1088# 0.070848f
C78 minus.t0 a_n2542_n1088# 0.064397f
C79 minus.n19 a_n2542_n1088# 0.067101f
C80 minus.n20 a_n2542_n1088# 0.008619f
C81 minus.n21 a_n2542_n1088# 0.037981f
C82 minus.n22 a_n2542_n1088# 0.037981f
C83 minus.n23 a_n2542_n1088# 0.037981f
C84 minus.n24 a_n2542_n1088# 0.008619f
C85 minus.t15 a_n2542_n1088# 0.064397f
C86 minus.n25 a_n2542_n1088# 0.070613f
C87 minus.t3 a_n2542_n1088# 0.064397f
C88 minus.n26 a_n2542_n1088# 0.066984f
C89 minus.n27 a_n2542_n1088# 1.01985f
C90 minus.n28 a_n2542_n1088# 0.037981f
C91 minus.t5 a_n2542_n1088# 0.064397f
C92 minus.n29 a_n2542_n1088# 0.070965f
C93 minus.n30 a_n2542_n1088# 0.037981f
C94 minus.n31 a_n2542_n1088# 0.008619f
C95 minus.n32 a_n2542_n1088# 0.037981f
C96 minus.t7 a_n2542_n1088# 0.064397f
C97 minus.n33 a_n2542_n1088# 0.070965f
C98 minus.t8 a_n2542_n1088# 0.073917f
C99 minus.n34 a_n2542_n1088# 0.057754f
C100 minus.t13 a_n2542_n1088# 0.064397f
C101 minus.n35 a_n2542_n1088# 0.070613f
C102 minus.n36 a_n2542_n1088# 0.008619f
C103 minus.n37 a_n2542_n1088# 0.124658f
C104 minus.n38 a_n2542_n1088# 0.037981f
C105 minus.n39 a_n2542_n1088# 0.037981f
C106 minus.n40 a_n2542_n1088# 0.008619f
C107 minus.t10 a_n2542_n1088# 0.064397f
C108 minus.n41 a_n2542_n1088# 0.067101f
C109 minus.t19 a_n2542_n1088# 0.064397f
C110 minus.n42 a_n2542_n1088# 0.070848f
C111 minus.n43 a_n2542_n1088# 0.037981f
C112 minus.n44 a_n2542_n1088# 0.037981f
C113 minus.n45 a_n2542_n1088# 0.037981f
C114 minus.t14 a_n2542_n1088# 0.064397f
C115 minus.n46 a_n2542_n1088# 0.070848f
C116 minus.t18 a_n2542_n1088# 0.064397f
C117 minus.n47 a_n2542_n1088# 0.067101f
C118 minus.n48 a_n2542_n1088# 0.008619f
C119 minus.n49 a_n2542_n1088# 0.037981f
C120 minus.n50 a_n2542_n1088# 0.037981f
C121 minus.n51 a_n2542_n1088# 0.037981f
C122 minus.n52 a_n2542_n1088# 0.008619f
C123 minus.t16 a_n2542_n1088# 0.064397f
C124 minus.n53 a_n2542_n1088# 0.070613f
C125 minus.t2 a_n2542_n1088# 0.064397f
C126 minus.n54 a_n2542_n1088# 0.066984f
C127 minus.n55 a_n2542_n1088# 0.256455f
C128 minus.n56 a_n2542_n1088# 1.25312f
C129 drain_left.t18 a_n2542_n1088# 0.017428f
C130 drain_left.t1 a_n2542_n1088# 0.017428f
C131 drain_left.n0 a_n2542_n1088# 0.068507f
C132 drain_left.t15 a_n2542_n1088# 0.017428f
C133 drain_left.t4 a_n2542_n1088# 0.017428f
C134 drain_left.n1 a_n2542_n1088# 0.06772f
C135 drain_left.n2 a_n2542_n1088# 0.516784f
C136 drain_left.t7 a_n2542_n1088# 0.017428f
C137 drain_left.t19 a_n2542_n1088# 0.017428f
C138 drain_left.n3 a_n2542_n1088# 0.06772f
C139 drain_left.t8 a_n2542_n1088# 0.017428f
C140 drain_left.t11 a_n2542_n1088# 0.017428f
C141 drain_left.n4 a_n2542_n1088# 0.068507f
C142 drain_left.t6 a_n2542_n1088# 0.017428f
C143 drain_left.t13 a_n2542_n1088# 0.017428f
C144 drain_left.n5 a_n2542_n1088# 0.06772f
C145 drain_left.n6 a_n2542_n1088# 0.516784f
C146 drain_left.n7 a_n2542_n1088# 0.960695f
C147 drain_left.t16 a_n2542_n1088# 0.017428f
C148 drain_left.t9 a_n2542_n1088# 0.017428f
C149 drain_left.n8 a_n2542_n1088# 0.068507f
C150 drain_left.t2 a_n2542_n1088# 0.017428f
C151 drain_left.t14 a_n2542_n1088# 0.017428f
C152 drain_left.n9 a_n2542_n1088# 0.06772f
C153 drain_left.n10 a_n2542_n1088# 0.519943f
C154 drain_left.t5 a_n2542_n1088# 0.017428f
C155 drain_left.t0 a_n2542_n1088# 0.017428f
C156 drain_left.n11 a_n2542_n1088# 0.06772f
C157 drain_left.n12 a_n2542_n1088# 0.255923f
C158 drain_left.t12 a_n2542_n1088# 0.017428f
C159 drain_left.t3 a_n2542_n1088# 0.017428f
C160 drain_left.n13 a_n2542_n1088# 0.06772f
C161 drain_left.n14 a_n2542_n1088# 0.255923f
C162 drain_left.t17 a_n2542_n1088# 0.017428f
C163 drain_left.t10 a_n2542_n1088# 0.017428f
C164 drain_left.n15 a_n2542_n1088# 0.06772f
C165 drain_left.n16 a_n2542_n1088# 0.445401f
C166 source.t21 a_n2542_n1088# 0.161959f
C167 source.n0 a_n2542_n1088# 0.732019f
C168 source.t29 a_n2542_n1088# 0.029099f
C169 source.t17 a_n2542_n1088# 0.029099f
C170 source.n1 a_n2542_n1088# 0.094371f
C171 source.n2 a_n2542_n1088# 0.395949f
C172 source.t33 a_n2542_n1088# 0.029099f
C173 source.t20 a_n2542_n1088# 0.029099f
C174 source.n3 a_n2542_n1088# 0.094371f
C175 source.n4 a_n2542_n1088# 0.395949f
C176 source.t24 a_n2542_n1088# 0.029099f
C177 source.t25 a_n2542_n1088# 0.029099f
C178 source.n5 a_n2542_n1088# 0.094371f
C179 source.n6 a_n2542_n1088# 0.395949f
C180 source.t31 a_n2542_n1088# 0.029099f
C181 source.t23 a_n2542_n1088# 0.029099f
C182 source.n7 a_n2542_n1088# 0.094371f
C183 source.n8 a_n2542_n1088# 0.395949f
C184 source.t26 a_n2542_n1088# 0.161959f
C185 source.n9 a_n2542_n1088# 0.37857f
C186 source.t6 a_n2542_n1088# 0.161959f
C187 source.n10 a_n2542_n1088# 0.37857f
C188 source.t10 a_n2542_n1088# 0.029099f
C189 source.t15 a_n2542_n1088# 0.029099f
C190 source.n11 a_n2542_n1088# 0.094371f
C191 source.n12 a_n2542_n1088# 0.395949f
C192 source.t37 a_n2542_n1088# 0.029099f
C193 source.t4 a_n2542_n1088# 0.029099f
C194 source.n13 a_n2542_n1088# 0.094371f
C195 source.n14 a_n2542_n1088# 0.395949f
C196 source.t14 a_n2542_n1088# 0.029099f
C197 source.t38 a_n2542_n1088# 0.029099f
C198 source.n15 a_n2542_n1088# 0.094371f
C199 source.n16 a_n2542_n1088# 0.395949f
C200 source.t3 a_n2542_n1088# 0.029099f
C201 source.t8 a_n2542_n1088# 0.029099f
C202 source.n17 a_n2542_n1088# 0.094371f
C203 source.n18 a_n2542_n1088# 0.395949f
C204 source.t39 a_n2542_n1088# 0.161959f
C205 source.n19 a_n2542_n1088# 1.0314f
C206 source.t16 a_n2542_n1088# 0.161958f
C207 source.n20 a_n2542_n1088# 1.0314f
C208 source.t22 a_n2542_n1088# 0.029099f
C209 source.t18 a_n2542_n1088# 0.029099f
C210 source.n21 a_n2542_n1088# 0.094371f
C211 source.n22 a_n2542_n1088# 0.395949f
C212 source.t34 a_n2542_n1088# 0.029099f
C213 source.t30 a_n2542_n1088# 0.029099f
C214 source.n23 a_n2542_n1088# 0.094371f
C215 source.n24 a_n2542_n1088# 0.395949f
C216 source.t28 a_n2542_n1088# 0.029099f
C217 source.t32 a_n2542_n1088# 0.029099f
C218 source.n25 a_n2542_n1088# 0.094371f
C219 source.n26 a_n2542_n1088# 0.395949f
C220 source.t27 a_n2542_n1088# 0.029099f
C221 source.t35 a_n2542_n1088# 0.029099f
C222 source.n27 a_n2542_n1088# 0.094371f
C223 source.n28 a_n2542_n1088# 0.395949f
C224 source.t19 a_n2542_n1088# 0.161958f
C225 source.n29 a_n2542_n1088# 0.37857f
C226 source.t11 a_n2542_n1088# 0.161958f
C227 source.n30 a_n2542_n1088# 0.37857f
C228 source.t7 a_n2542_n1088# 0.029099f
C229 source.t9 a_n2542_n1088# 0.029099f
C230 source.n31 a_n2542_n1088# 0.094371f
C231 source.n32 a_n2542_n1088# 0.395949f
C232 source.t13 a_n2542_n1088# 0.029099f
C233 source.t2 a_n2542_n1088# 0.029099f
C234 source.n33 a_n2542_n1088# 0.094371f
C235 source.n34 a_n2542_n1088# 0.395949f
C236 source.t1 a_n2542_n1088# 0.029099f
C237 source.t0 a_n2542_n1088# 0.029099f
C238 source.n35 a_n2542_n1088# 0.094371f
C239 source.n36 a_n2542_n1088# 0.395949f
C240 source.t12 a_n2542_n1088# 0.029099f
C241 source.t5 a_n2542_n1088# 0.029099f
C242 source.n37 a_n2542_n1088# 0.094371f
C243 source.n38 a_n2542_n1088# 0.395949f
C244 source.t36 a_n2542_n1088# 0.161958f
C245 source.n39 a_n2542_n1088# 0.602692f
C246 source.n40 a_n2542_n1088# 0.754282f
C247 plus.n0 a_n2542_n1088# 0.038442f
C248 plus.t9 a_n2542_n1088# 0.065179f
C249 plus.t2 a_n2542_n1088# 0.065179f
C250 plus.t16 a_n2542_n1088# 0.065179f
C251 plus.n1 a_n2542_n1088# 0.071827f
C252 plus.n2 a_n2542_n1088# 0.038442f
C253 plus.t7 a_n2542_n1088# 0.065179f
C254 plus.t19 a_n2542_n1088# 0.065179f
C255 plus.n3 a_n2542_n1088# 0.038442f
C256 plus.t14 a_n2542_n1088# 0.065179f
C257 plus.n4 a_n2542_n1088# 0.071708f
C258 plus.n5 a_n2542_n1088# 0.038442f
C259 plus.t5 a_n2542_n1088# 0.065179f
C260 plus.t17 a_n2542_n1088# 0.065179f
C261 plus.n6 a_n2542_n1088# 0.038442f
C262 plus.t10 a_n2542_n1088# 0.065179f
C263 plus.n7 a_n2542_n1088# 0.071471f
C264 plus.t3 a_n2542_n1088# 0.074815f
C265 plus.n8 a_n2542_n1088# 0.058456f
C266 plus.n9 a_n2542_n1088# 0.126172f
C267 plus.n10 a_n2542_n1088# 0.008723f
C268 plus.n11 a_n2542_n1088# 0.071827f
C269 plus.n12 a_n2542_n1088# 0.008723f
C270 plus.n13 a_n2542_n1088# 0.067916f
C271 plus.n14 a_n2542_n1088# 0.038442f
C272 plus.n15 a_n2542_n1088# 0.038442f
C273 plus.n16 a_n2542_n1088# 0.038442f
C274 plus.n17 a_n2542_n1088# 0.008723f
C275 plus.n18 a_n2542_n1088# 0.071708f
C276 plus.n19 a_n2542_n1088# 0.067916f
C277 plus.n20 a_n2542_n1088# 0.008723f
C278 plus.n21 a_n2542_n1088# 0.038442f
C279 plus.n22 a_n2542_n1088# 0.038442f
C280 plus.n23 a_n2542_n1088# 0.038442f
C281 plus.n24 a_n2542_n1088# 0.008723f
C282 plus.n25 a_n2542_n1088# 0.071471f
C283 plus.n26 a_n2542_n1088# 0.067797f
C284 plus.n27 a_n2542_n1088# 0.272251f
C285 plus.n28 a_n2542_n1088# 0.038442f
C286 plus.t1 a_n2542_n1088# 0.065179f
C287 plus.t18 a_n2542_n1088# 0.065179f
C288 plus.t4 a_n2542_n1088# 0.065179f
C289 plus.n29 a_n2542_n1088# 0.071827f
C290 plus.n30 a_n2542_n1088# 0.038442f
C291 plus.t15 a_n2542_n1088# 0.065179f
C292 plus.n31 a_n2542_n1088# 0.038442f
C293 plus.t12 a_n2542_n1088# 0.065179f
C294 plus.t0 a_n2542_n1088# 0.065179f
C295 plus.n32 a_n2542_n1088# 0.071708f
C296 plus.n33 a_n2542_n1088# 0.038442f
C297 plus.t13 a_n2542_n1088# 0.065179f
C298 plus.n34 a_n2542_n1088# 0.038442f
C299 plus.t6 a_n2542_n1088# 0.065179f
C300 plus.t11 a_n2542_n1088# 0.065179f
C301 plus.n35 a_n2542_n1088# 0.071471f
C302 plus.t8 a_n2542_n1088# 0.074815f
C303 plus.n36 a_n2542_n1088# 0.058456f
C304 plus.n37 a_n2542_n1088# 0.126172f
C305 plus.n38 a_n2542_n1088# 0.008723f
C306 plus.n39 a_n2542_n1088# 0.071827f
C307 plus.n40 a_n2542_n1088# 0.008723f
C308 plus.n41 a_n2542_n1088# 0.067916f
C309 plus.n42 a_n2542_n1088# 0.038442f
C310 plus.n43 a_n2542_n1088# 0.038442f
C311 plus.n44 a_n2542_n1088# 0.038442f
C312 plus.n45 a_n2542_n1088# 0.008723f
C313 plus.n46 a_n2542_n1088# 0.071708f
C314 plus.n47 a_n2542_n1088# 0.067916f
C315 plus.n48 a_n2542_n1088# 0.008723f
C316 plus.n49 a_n2542_n1088# 0.038442f
C317 plus.n50 a_n2542_n1088# 0.038442f
C318 plus.n51 a_n2542_n1088# 0.038442f
C319 plus.n52 a_n2542_n1088# 0.008723f
C320 plus.n53 a_n2542_n1088# 0.071471f
C321 plus.n54 a_n2542_n1088# 0.067797f
C322 plus.n55 a_n2542_n1088# 0.99578f
.ends

